module SPEEDY_Rounds7_0 ( Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  wire   n2, n3, n4, n5, n7, n10, n11, n12, n13, n17, n19, n21, n25, n26, n28,
         n29, n32, n35, n36, n37, n40, n42, n43, n45, n46, n50, n52, n53, n54,
         n56, n57, n59, n61, n62, n63, n64, n70, n71, n76, n81, n85, n89, n94,
         n98, n99, n104, n105, n106, n109, n110, n113, n114, n118, n119, n121,
         n122, n123, n124, n126, n129, n130, n133, n135, n137, n138, n139,
         n140, n142, n149, n154, n155, n156, n157, n158, n159, n160, n161,
         n164, n167, n170, n171, n178, n180, n182, n183, n184, n187, n190,
         n193, n195, n196, n197, n198, n199, n200, n205, n207, n208, n209,
         n212, n214, n215, n217, n219, n220, n224, n229, n230, n231, n232,
         n233, n237, n238, n242, n248, n250, n251, n252, n253, n254, n257,
         n259, n260, n261, n263, n266, n269, n272, n274, n275, n277, n278,
         n280, n281, n282, n284, n287, n288, n291, n293, n295, n296, n298,
         n299, n301, n302, n305, n306, n307, n309, n310, n311, n314, n317,
         n318, n319, n320, n321, n326, n327, n331, n334, n336, n342, n343,
         n344, n345, n346, n347, n353, n354, n355, n357, n359, n360, n362,
         n364, n365, n367, n370, n371, n372, n378, n379, n382, n383, n384,
         n385, n386, n387, n388, n391, n396, n399, n400, n404, n406, n407,
         n411, n412, n416, n422, n423, n424, n425, n427, n430, n431, n434,
         n436, n437, n438, n439, n440, n441, n442, n443, n445, n446, n447,
         n449, n450, n451, n452, n454, n455, n457, n459, n462, n465, n467,
         n471, n474, n476, n479, n481, n482, n484, n485, n487, n489, n491,
         n494, n495, n496, n502, n505, n507, n509, n514, n515, n517, n518,
         n523, n524, n525, n526, n528, n529, n530, n531, n532, n533, n538,
         n540, n541, n542, n543, n545, n547, n548, n550, n551, n552, n554,
         n556, n557, n560, n562, n566, n576, n579, n580, n583, n584, n585,
         n586, n587, n588, n589, n591, n596, n598, n599, n601, n603, n605,
         n606, n608, n609, n611, n614, n615, n616, n619, n621, n626, n628,
         n629, n632, n633, n635, n636, n637, n638, n639, n640, n642, n644,
         n646, n648, n649, n650, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n672,
         n673, n674, n675, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n688, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n704, n705, n706, n707, n708, n709, n710,
         n711, n713, n714, n718, n719, n720, n721, n722, n723, n724, n727,
         n728, n729, n730, n731, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n754, n755, n756, n759, n760, n761, n762, n763, n764, n765,
         n767, n769, n770, n771, n772, n773, n774, n775, n777, n778, n779,
         n780, n781, n782, n783, n784, n787, n788, n789, n790, n791, n792,
         n794, n798, n800, n801, n802, n807, n808, n810, n812, n813, n814,
         n815, n816, n817, n819, n820, n821, n823, n824, n825, n826, n828,
         n830, n831, n832, n833, n834, n835, n837, n838, n839, n840, n841,
         n844, n845, n846, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n865, n866, n867,
         n869, n870, n871, n873, n875, n876, n877, n878, n879, n881, n882,
         n883, n885, n886, n888, n889, n892, n893, n894, n896, n898, n900,
         n902, n903, n906, n907, n910, n911, n914, n915, n916, n917, n918,
         n919, n920, n921, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n933, n934, n935, n936, n937, n938, n939, n941, n943, n944,
         n945, n946, n948, n949, n950, n951, n952, n953, n954, n955, n957,
         n958, n959, n960, n961, n962, n963, n965, n966, n967, n968, n969,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n997, n998, n999, n1000, n1002, n1003, n1006, n1008,
         n1009, n1010, n1011, n1012, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1024, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1038, n1039, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1065,
         n1066, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1076, n1077,
         n1079, n1080, n1081, n1082, n1084, n1085, n1086, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1112,
         n1113, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1151, n1152, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1165, n1167,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1181, n1182, n1183, n1184, n1186, n1187, n1189, n1190, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1200, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1211, n1212, n1214, n1215, n1217,
         n1218, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1229,
         n1230, n1231, n1232, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1242, n1243, n1244, n1245, n1249, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1265, n1267, n1268,
         n1269, n1270, n1271, n1273, n1274, n1275, n1276, n1279, n1280, n1282,
         n1283, n1284, n1285, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1297, n1298, n1299, n1300, n1301, n1302, n1304, n1306, n1307,
         n1308, n1310, n1312, n1313, n1314, n1315, n1316, n1318, n1319, n1320,
         n1322, n1323, n1324, n1326, n1327, n1328, n1329, n1331, n1332, n1333,
         n1334, n1335, n1337, n1338, n1339, n1340, n1341, n1342, n1344, n1345,
         n1346, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1361, n1362, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1374, n1375, n1377, n1378, n1379, n1380, n1382, n1383,
         n1385, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1424, n1425, n1426, n1427, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1444, n1445, n1446, n1447, n1448, n1450, n1451, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1477, n1478, n1480, n1481, n1483, n1484, n1486, n1487, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1497, n1500, n1502, n1503,
         n1504, n1505, n1506, n1507, n1509, n1510, n1511, n1512, n1514, n1515,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1527, n1528, n1529,
         n1530, n1531, n1532, n1534, n1535, n1536, n1537, n1539, n1541, n1543,
         n1545, n1546, n1547, n1548, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1563, n1564, n1565, n1566, n1567,
         n1570, n1573, n1574, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1586, n1587, n1588, n1589, n1591, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1612, n1613, n1614, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1675, n1676,
         n1678, n1679, n1680, n1681, n1683, n1684, n1686, n1687, n1688, n1689,
         n1690, n1692, n1693, n1694, n1695, n1697, n1698, n1699, n1700, n1702,
         n1703, n1704, n1706, n1707, n1708, n1710, n1711, n1713, n1714, n1717,
         n1718, n1719, n1722, n1723, n1724, n1725, n1726, n1727, n1730, n1733,
         n1734, n1735, n1737, n1738, n1740, n1741, n1742, n1743, n1745, n1746,
         n1752, n1753, n1755, n1757, n1758, n1759, n1760, n1763, n1765, n1766,
         n1769, n1771, n1775, n1777, n1778, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1790, n1791, n1792, n1793, n1794, n1796, n1797,
         n1798, n1799, n1802, n1805, n1807, n1808, n1809, n1812, n1813, n1814,
         n1815, n1816, n1817, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1827, n1829, n1830, n1831, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1842, n1843, n1844, n1845, n1847, n1849, n1850, n1851, n1852,
         n1855, n1859, n1861, n1862, n1864, n1865, n1866, n1867, n1868, n1872,
         n1873, n1874, n1875, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1890, n1891, n1893, n1894, n1895, n1896, n1897,
         n1898, n1902, n1904, n1906, n1907, n1909, n1911, n1912, n1913, n1914,
         n1915, n1917, n1918, n1919, n1921, n1923, n1929, n1930, n1932, n1933,
         n1934, n1936, n1938, n1939, n1940, n1944, n1945, n1946, n1947, n1948,
         n1949, n1951, n1953, n1954, n1956, n1961, n1962, n1965, n1966, n1969,
         n1971, n1978, n1980, n1984, n1986, n1989, n1990, n1991, n1992, n1993,
         n1995, n1996, n1997, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2008, n2009, n2012, n2013, n2016, n2017, n2018, n2022, n2023, n2025,
         n2028, n2029, n2030, n2031, n2032, n2035, n2036, n2041, n2042, n2044,
         n2045, n2046, n2047, n2049, n2050, n2052, n2055, n2057, n2058, n2059,
         n2060, n2062, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2073,
         n2075, n2076, n2077, n2078, n2079, n2081, n2082, n2084, n2085, n2086,
         n2087, n2088, n2089, n2091, n2092, n2094, n2096, n2097, n2100, n2101,
         n2102, n2104, n2105, n2106, n2107, n2110, n2111, n2112, n2113, n2114,
         n2116, n2117, n2119, n2120, n2121, n2122, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2132, n2134, n2135, n2136, n2138, n2139, n2140,
         n2142, n2145, n2147, n2148, n2149, n2150, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2166,
         n2167, n2168, n2170, n2175, n2176, n2177, n2178, n2182, n2184, n2185,
         n2186, n2187, n2189, n2190, n2191, n2192, n2193, n2195, n2196, n2198,
         n2199, n2200, n2202, n2203, n2205, n2207, n2208, n2209, n2211, n2214,
         n2215, n2216, n2217, n2218, n2220, n2221, n2222, n2223, n2226, n2229,
         n2231, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2242, n2243,
         n2246, n2247, n2248, n2250, n2253, n2254, n2257, n2258, n2259, n2260,
         n2262, n2263, n2264, n2268, n2269, n2270, n2272, n2273, n2274, n2276,
         n2277, n2278, n2279, n2280, n2281, n2283, n2284, n2285, n2288, n2292,
         n2294, n2296, n2297, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2309, n2310, n2311, n2316, n2317, n2318, n2319, n2321, n2322, n2326,
         n2327, n2328, n2330, n2331, n2333, n2334, n2335, n2336, n2338, n2339,
         n2340, n2341, n2342, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2354, n2356, n2362, n2363, n2364, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2398, n2400, n2402, n2403, n2404, n2405, n2410, n2413, n2416,
         n2417, n2418, n2421, n2423, n2424, n2428, n2429, n2430, n2431, n2434,
         n2435, n2436, n2437, n2439, n2443, n2445, n2446, n2448, n2449, n2450,
         n2451, n2453, n2454, n2456, n2457, n2458, n2461, n2462, n2464, n2465,
         n2466, n2467, n2469, n2471, n2473, n2474, n2475, n2476, n2478, n2479,
         n2480, n2481, n2482, n2484, n2485, n2487, n2488, n2489, n2490, n2491,
         n2493, n2495, n2496, n2498, n2500, n2502, n2503, n2505, n2506, n2507,
         n2510, n2511, n2512, n2515, n2518, n2519, n2520, n2522, n2524, n2525,
         n2526, n2527, n2529, n2530, n2531, n2532, n2533, n2534, n2537, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2549, n2553, n2554, n2555,
         n2557, n2559, n2560, n2561, n2563, n2566, n2569, n2572, n2573, n2574,
         n2576, n2579, n2580, n2581, n2582, n2585, n2586, n2587, n2588, n2589,
         n2590, n2592, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2603, n2604, n2607, n2608, n2610, n2613, n2614, n2615, n2616, n2618,
         n2621, n2622, n2623, n2625, n2626, n2627, n2628, n2629, n2630, n2632,
         n2633, n2634, n2635, n2637, n2639, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2653, n2654, n2656, n2657, n2658, n2660,
         n2662, n2663, n2664, n2666, n2667, n2668, n2671, n2674, n2675, n2677,
         n2678, n2679, n2681, n2682, n2683, n2684, n2685, n2688, n2690, n2692,
         n2695, n2696, n2697, n2698, n2701, n2703, n2704, n2705, n2707, n2709,
         n2711, n2712, n2713, n2714, n2716, n2717, n2721, n2722, n2725, n2726,
         n2727, n2728, n2730, n2731, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2745, n2746, n2747, n2751, n2752, n2753, n2754,
         n2757, n2758, n2759, n2760, n2761, n2765, n2766, n2767, n2768, n2769,
         n2771, n2772, n2774, n2778, n2780, n2781, n2782, n2784, n2785, n2788,
         n2789, n2790, n2792, n2794, n2795, n2796, n2798, n2799, n2800, n2801,
         n2802, n2803, n2805, n2806, n2808, n2812, n2813, n2814, n2815, n2816,
         n2818, n2819, n2822, n2823, n2824, n2825, n2830, n2832, n2833, n2835,
         n2837, n2838, n2839, n2840, n2841, n2842, n2846, n2847, n2848, n2850,
         n2853, n2856, n2858, n2859, n2860, n2861, n2864, n2865, n2866, n2867,
         n2868, n2870, n2872, n2873, n2874, n2876, n2877, n2878, n2880, n2881,
         n2882, n2883, n2886, n2888, n2889, n2891, n2892, n2895, n2896, n2898,
         n2899, n2900, n2903, n2904, n2905, n2906, n2907, n2909, n2910, n2914,
         n2915, n2919, n2920, n2921, n2922, n2923, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2935, n2937, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2949, n2950, n2953, n2954, n2955, n2957, n2958,
         n2959, n2960, n2961, n2962, n2965, n2966, n2967, n2968, n2969, n2971,
         n2972, n2974, n2975, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2995, n2996, n2997,
         n2998, n3001, n3002, n3003, n3004, n3005, n3006, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3018, n3019, n3021, n3022, n3023, n3024,
         n3025, n3027, n3028, n3029, n3031, n3032, n3035, n3036, n3037, n3039,
         n3040, n3041, n3044, n3045, n3046, n3047, n3048, n3050, n3052, n3053,
         n3055, n3056, n3057, n3058, n3059, n3060, n3065, n3066, n3067, n3069,
         n3070, n3071, n3072, n3076, n3077, n3081, n3082, n3083, n3085, n3086,
         n3088, n3090, n3091, n3092, n3093, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3105, n3106, n3107, n3109, n3110, n3111,
         n3112, n3114, n3116, n3117, n3118, n3119, n3120, n3122, n3124, n3125,
         n3126, n3127, n3128, n3129, n3133, n3134, n3135, n3136, n3137, n3140,
         n3141, n3142, n3145, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3161, n3163, n3164, n3166, n3167, n3169, n3170,
         n3172, n3174, n3175, n3181, n3185, n3186, n3187, n3188, n3190, n3191,
         n3192, n3193, n3194, n3195, n3198, n3199, n3200, n3203, n3206, n3207,
         n3213, n3214, n3215, n3217, n3218, n3219, n3221, n3223, n3224, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3239, n3240, n3241, n3242, n3244, n3245, n3246, n3247, n3248,
         n3250, n3252, n3253, n3255, n3256, n3257, n3258, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3273, n3274,
         n3275, n3276, n3277, n3278, n3280, n3282, n3283, n3284, n3285, n3287,
         n3288, n3289, n3290, n3292, n3293, n3294, n3295, n3297, n3299, n3301,
         n3303, n3304, n3305, n3307, n3309, n3310, n3312, n3313, n3316, n3317,
         n3319, n3320, n3323, n3325, n3326, n3327, n3328, n3330, n3331, n3332,
         n3333, n3336, n3337, n3342, n3343, n3345, n3346, n3348, n3349, n3350,
         n3351, n3352, n3356, n3359, n3360, n3361, n3363, n3364, n3365, n3366,
         n3368, n3369, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3382, n3383, n3386, n3387, n3388, n3389, n3390, n3392, n3393,
         n3395, n3398, n3399, n3402, n3404, n3409, n3410, n3411, n3412, n3413,
         n3415, n3417, n3422, n3424, n3426, n3427, n3429, n3430, n3433, n3434,
         n3435, n3437, n3438, n3441, n3443, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3478, n3480, n3484, n3486,
         n3487, n3488, n3489, n3490, n3493, n3495, n3496, n3497, n3498, n3499,
         n3501, n3503, n3506, n3507, n3509, n3510, n3511, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3521, n3522, n3523, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3538, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3557, n3559, n3560, n3561, n3562,
         n3564, n3568, n3571, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3581, n3583, n3584, n3585, n3589, n3593, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3609, n3610, n3611, n3612, n3614,
         n3616, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3637, n3638, n3639,
         n3641, n3642, n3644, n3645, n3647, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3659, n3662, n3663, n3664, n3665, n3666,
         n3668, n3669, n3670, n3671, n3672, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3685, n3687, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3703,
         n3705, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3722, n3723, n3725, n3726, n3727, n3731, n3732,
         n3733, n3734, n3735, n3736, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3760, n3761, n3769, n3770, n3771, n3773,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3787, n3790, n3791, n3792, n3793, n3794, n3795, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3806, n3807, n3809, n3811, n3813, n3815,
         n3818, n3819, n3820, n3821, n3823, n3824, n3825, n3826, n3827, n3832,
         n3833, n3835, n3837, n3838, n3839, n3840, n3843, n3844, n3845, n3846,
         n3849, n3850, n3851, n3852, n3855, n3857, n3858, n3860, n3861, n3862,
         n3863, n3864, n3865, n3867, n3868, n3869, n3872, n3873, n3874, n3877,
         n3878, n3879, n3884, n3885, n3886, n3887, n3889, n3890, n3891, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3903, n3904, n3906,
         n3907, n3909, n3912, n3913, n3914, n3916, n3917, n3918, n3919, n3920,
         n3921, n3923, n3926, n3927, n3928, n3929, n3930, n3932, n3935, n3937,
         n3938, n3941, n3943, n3944, n3945, n3947, n3949, n3951, n3952, n3953,
         n3954, n3956, n3958, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3969, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3981, n3983, n3985, n3986, n3988, n3989, n3990, n3992, n3993, n3995,
         n3996, n3998, n3999, n4000, n4001, n4002, n4005, n4007, n4008, n4009,
         n4010, n4011, n4013, n4014, n4015, n4016, n4018, n4021, n4022, n4023,
         n4024, n4025, n4028, n4033, n4034, n4037, n4038, n4039, n4041, n4045,
         n4046, n4047, n4048, n4050, n4051, n4053, n4056, n4057, n4058, n4059,
         n4061, n4062, n4063, n4064, n4065, n4066, n4070, n4072, n4073, n4075,
         n4076, n4077, n4079, n4080, n4081, n4083, n4084, n4085, n4086, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4098, n4099, n4100, n4102,
         n4104, n4105, n4107, n4108, n4109, n4110, n4111, n4114, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4126, n4127, n4128, n4129,
         n4131, n4132, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4159, n4160, n4161, n4162, n4163, n4168, n4169, n4171, n4172, n4173,
         n4176, n4177, n4178, n4179, n4182, n4183, n4184, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4204, n4205, n4207, n4209, n4210, n4211, n4214, n4215, n4216,
         n4217, n4218, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4231, n4232, n4235, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4246, n4247, n4248, n4251, n4253, n4254, n4255, n4256,
         n4257, n4258, n4266, n4268, n4269, n4270, n4271, n4272, n4273, n4277,
         n4278, n4279, n4280, n4282, n4283, n4284, n4286, n4287, n4288, n4290,
         n4291, n4292, n4293, n4294, n4296, n4297, n4298, n4300, n4301, n4302,
         n4305, n4306, n4308, n4313, n4314, n4315, n4316, n4317, n4318, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4332,
         n4333, n4334, n4335, n4336, n4337, n4339, n4340, n4341, n4342, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4359, n4360, n4361, n4362, n4364, n4366, n4367, n4368,
         n4369, n4371, n4372, n4373, n4375, n4377, n4378, n4379, n4381, n4382,
         n4384, n4385, n4386, n4387, n4388, n4391, n4392, n4393, n4396, n4397,
         n4398, n4399, n4400, n4401, n4409, n4410, n4411, n4412, n4413, n4415,
         n4416, n4417, n4419, n4423, n4424, n4427, n4428, n4429, n4430, n4431,
         n4433, n4434, n4436, n4438, n4439, n4440, n4441, n4442, n4443, n4445,
         n4447, n4448, n4449, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4472, n4473, n4475, n4476, n4477, n4479, n4483, n4484, n4485,
         n4486, n4489, n4490, n4492, n4493, n4494, n4495, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4506, n4507, n4508, n4511, n4512,
         n4515, n4516, n4518, n4519, n4520, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4531, n4534, n4536, n4538, n4540, n4542, n4543, n4549,
         n4550, n4551, n4552, n4553, n4556, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4568, n4570, n4572, n4573, n4574, n4576,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4587, n4588, n4589,
         n4591, n4592, n4595, n4597, n4599, n4600, n4601, n4602, n4603, n4604,
         n4606, n4608, n4610, n4611, n4612, n4613, n4616, n4618, n4619, n4620,
         n4621, n4622, n4624, n4625, n4627, n4629, n4630, n4631, n4632, n4633,
         n4634, n4636, n4637, n4638, n4640, n4641, n4642, n4644, n4646, n4647,
         n4649, n4651, n4655, n4656, n4658, n4660, n4661, n4662, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4673, n4674, n4677, n4682,
         n4686, n4687, n4688, n4689, n4690, n4694, n4697, n4698, n4699, n4700,
         n4702, n4703, n4704, n4707, n4709, n4713, n4714, n4715, n4716, n4720,
         n4724, n4726, n4729, n4730, n4734, n4736, n4737, n4738, n4739, n4741,
         n4743, n4745, n4746, n4748, n4750, n4752, n4754, n4755, n4756, n4759,
         n4760, n4761, n4765, n4766, n4767, n4768, n4769, n4771, n4772, n4773,
         n4775, n4776, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4788,
         n4790, n4791, n4792, n4794, n4796, n4799, n4800, n4801, n4803, n4805,
         n4807, n4808, n4809, n4815, n4816, n4819, n4821, n4823, n4824, n4825,
         n4827, n4828, n4829, n4832, n4833, n4834, n4840, n4841, n4845, n4846,
         n4847, n4849, n4850, n4851, n4852, n4853, n4854, n4856, n4857, n4858,
         n4859, n4862, n4864, n4865, n4866, n4867, n4868, n4869, n4871, n4874,
         n4875, n4876, n4878, n4879, n4880, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4905, n4908, n4909, n4910, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4924, n4925, n4926, n4927,
         n4929, n4931, n4932, n4934, n4935, n4936, n4937, n4938, n4941, n4945,
         n4946, n4947, n4948, n4949, n4950, n4952, n4956, n4957, n4958, n4959,
         n4960, n4963, n4964, n4967, n4968, n4969, n4970, n4972, n4973, n4975,
         n4976, n4977, n4978, n4980, n4982, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4997, n4999, n5001, n5002, n5003, n5005, n5006,
         n5009, n5010, n5011, n5012, n5014, n5015, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5026, n5027, n5028, n5030, n5031, n5033, n5034,
         n5035, n5037, n5038, n5039, n5041, n5042, n5044, n5047, n5048, n5049,
         n5050, n5051, n5053, n5054, n5055, n5056, n5058, n5059, n5061, n5062,
         n5063, n5065, n5066, n5067, n5070, n5071, n5073, n5075, n5077, n5078,
         n5080, n5082, n5083, n5084, n5085, n5086, n5088, n5089, n5090, n5091,
         n5093, n5094, n5096, n5098, n5100, n5101, n5103, n5104, n5107, n5108,
         n5110, n5111, n5112, n5114, n5115, n5116, n5118, n5119, n5120, n5122,
         n5123, n5124, n5126, n5127, n5129, n5130, n5131, n5132, n5137, n5138,
         n5139, n5140, n5142, n5143, n5144, n5145, n5146, n5147, n5149, n5150,
         n5151, n5152, n5153, n5154, n5156, n5158, n5160, n5161, n5162, n5164,
         n5166, n5167, n5171, n5172, n5174, n5176, n5177, n5179, n5181, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5214, n5215, n5218, n5219, n5220, n5221, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5231, n5232, n5233, n5235, n5236, n5237,
         n5238, n5239, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5251, n5252, n5253, n5254, n5255, n5258, n5261, n5263, n5264,
         n5266, n5270, n5271, n5274, n5276, n5277, n5279, n5282, n5283, n5284,
         n5285, n5286, n5287, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5297, n5299, n5300, n5302, n5303, n5304, n5305, n5306, n5308, n5309,
         n5311, n5312, n5314, n5315, n5316, n5317, n5318, n5320, n5322, n5323,
         n5325, n5326, n5327, n5330, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5342, n5343, n5344, n5345, n5347, n5348, n5350, n5351, n5352,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5363, n5365,
         n5366, n5367, n5369, n5370, n5371, n5374, n5377, n5380, n5381, n5382,
         n5383, n5384, n5385, n5387, n5388, n5389, n5390, n5391, n5392, n5394,
         n5395, n5396, n5397, n5398, n5399, n5401, n5402, n5403, n5405, n5407,
         n5408, n5410, n5412, n5413, n5414, n5415, n5417, n5418, n5422, n5423,
         n5424, n5427, n5430, n5431, n5432, n5433, n5434, n5436, n5437, n5438,
         n5439, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5461, n5462, n5463, n5464, n5465, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5477, n5479, n5480, n5481, n5483, n5484,
         n5486, n5487, n5488, n5490, n5491, n5492, n5494, n5495, n5496, n5497,
         n5498, n5500, n5501, n5503, n5504, n5505, n5508, n5509, n5510, n5511,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5522, n5524, n5525,
         n5527, n5530, n5531, n5533, n5534, n5535, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5569,
         n5570, n5571, n5572, n5576, n5577, n5579, n5580, n5581, n5582, n5583,
         n5584, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5596, n5597,
         n5598, n5599, n5600, n5601, n5603, n5607, n5609, n5610, n5613, n5616,
         n5617, n5618, n5619, n5621, n5622, n5623, n5625, n5628, n5629, n5630,
         n5632, n5634, n5635, n5636, n5637, n5638, n5639, n5641, n5642, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5655, n5656,
         n5657, n5658, n5662, n5664, n5665, n5667, n5669, n5670, n5671, n5672,
         n5674, n5675, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5686, n5687, n5688, n5690, n5691, n5692, n5693, n5694, n5695, n5697,
         n5698, n5699, n5702, n5703, n5705, n5706, n5707, n5709, n5710, n5711,
         n5712, n5713, n5714, n5716, n5717, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5728, n5730, n5731, n5732, n5733, n5734, n5736,
         n5737, n5738, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5753, n5755, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5781, n5782,
         n5785, n5786, n5787, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5798, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5810, n5811, n5813, n5814, n5815, n5816, n5817, n5819, n5820, n5821,
         n5822, n5823, n5825, n5829, n5830, n5831, n5834, n5835, n5836, n5837,
         n5838, n5839, n5841, n5842, n5843, n5844, n5845, n5848, n5849, n5851,
         n5853, n5854, n5855, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5866, n5867, n5869, n5871, n5873, n5874, n5876, n5877, n5878,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5888, n5889, n5890,
         n5891, n5892, n5894, n5895, n5896, n5897, n5899, n5900, n5901, n5902,
         n5905, n5906, n5907, n5908, n5910, n5913, n5914, n5915, n5917, n5918,
         n5919, n5920, n5921, n5923, n5924, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5949, n5951, n5953, n5954,
         n5955, n5956, n5957, n5959, n5960, n5963, n5965, n5966, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5979, n5980,
         n5981, n5982, n5983, n5985, n5986, n5988, n5991, n5992, n5993, n5994,
         n5997, n5998, n5999, n6000, n6001, n6002, n6005, n6007, n6008, n6009,
         n6010, n6012, n6013, n6014, n6015, n6017, n6018, n6019, n6023, n6026,
         n6027, n6029, n6030, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6056, n6057, n6058, n6062, n6064,
         n6065, n6066, n6067, n6068, n6071, n6075, n6077, n6078, n6081, n6083,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6097,
         n6098, n6099, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6112, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6133,
         n6134, n6136, n6137, n6139, n6141, n6142, n6145, n6147, n6148, n6149,
         n6150, n6152, n6153, n6154, n6156, n6158, n6159, n6160, n6161, n6163,
         n6164, n6165, n6169, n6170, n6171, n6172, n6173, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6183, n6184, n6185, n6186, n6187, n6189,
         n6190, n6191, n6192, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6231, n6232, n6233, n6234,
         n6235, n6236, n6241, n6243, n6244, n6245, n6246, n6248, n6252, n6253,
         n6254, n6257, n6261, n6262, n6263, n6264, n6269, n6270, n6271, n6273,
         n6274, n6277, n6281, n6282, n6283, n6285, n6286, n6287, n6289, n6291,
         n6293, n6294, n6295, n6297, n6298, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6327, n6328, n6329, n6331, n6332, n6335, n6336, n6337, n6339, n6340,
         n6341, n6342, n6343, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6355, n6357, n6360, n6361, n6363, n6365, n6366, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6379, n6381,
         n6383, n6384, n6385, n6387, n6388, n6389, n6390, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6405,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6423, n6424, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6435, n6436, n6438, n6440, n6441, n6443,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6453, n6454, n6455,
         n6456, n6457, n6458, n6460, n6461, n6462, n6463, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6477, n6478,
         n6479, n6480, n6481, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6496, n6497, n6498, n6499, n6500, n6501,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6525, n6526, n6527, n6528, n6530, n6531, n6533, n6534, n6535, n6536,
         n6537, n6539, n6540, n6541, n6542, n6543, n6544, n6546, n6548, n6549,
         n6550, n6554, n6555, n6556, n6557, n6559, n6560, n6561, n6562, n6563,
         n6564, n6567, n6569, n6570, n6571, n6572, n6573, n6574, n6576, n6578,
         n6579, n6580, n6581, n6582, n6583, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6595, n6596, n6598, n6599, n6600, n6601,
         n6602, n6604, n6605, n6606, n6608, n6609, n6610, n6611, n6615, n6619,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6652, n6654,
         n6656, n6657, n6658, n6661, n6668, n6669, n6670, n6671, n6672, n6674,
         n6675, n6676, n6677, n6681, n6684, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6696, n6697, n6698, n6703, n6706, n6707,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6717, n6719, n6720,
         n6721, n6722, n6723, n6724, n6727, n6728, n6729, n6731, n6732, n6733,
         n6734, n6739, n6741, n6744, n6746, n6747, n6748, n6749, n6751, n6752,
         n6753, n6756, n6757, n6758, n6759, n6762, n6763, n6764, n6765, n6768,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6788, n6789, n6790, n6791,
         n6795, n6796, n6797, n6799, n6800, n6801, n6802, n6803, n6807, n6808,
         n6809, n6810, n6817, n6818, n6819, n6822, n6825, n6826, n6827, n6830,
         n6831, n6834, n6835, n6836, n6837, n6838, n6839, n6841, n6842, n6843,
         n6844, n6845, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6860, n6862, n6863, n6864, n6865, n6866, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6883, n6885, n6886, n6887, n6891,
         n6892, n6893, n6894, n6895, n6896, n6898, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6916, n6917, n6919, n6920, n6921, n6922, n6923, n6924, n6926, n6927,
         n6930, n6932, n6933, n6934, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6960, n6963, n6965, n6969, n6970, n6972, n6975,
         n6977, n6978, n6980, n6981, n6982, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7017, n7018, n7022, n7023,
         n7024, n7025, n7026, n7028, n7030, n7031, n7032, n7033, n7034, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7044, n7046, n7047, n7048,
         n7049, n7052, n7055, n7056, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7075, n7076,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7088, n7089,
         n7090, n7093, n7096, n7097, n7099, n7100, n7101, n7102, n7104, n7105,
         n7106, n7107, n7108, n7110, n7111, n7112, n7113, n7114, n7115, n7118,
         n7119, n7120, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7140, n7141, n7144,
         n7145, n7146, n7148, n7149, n7150, n7152, n7153, n7154, n7158, n7160,
         n7161, n7162, n7163, n7164, n7166, n7167, n7168, n7170, n7171, n7173,
         n7175, n7176, n7177, n7179, n7180, n7182, n7183, n7185, n7186, n7190,
         n7191, n7193, n7194, n7195, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7206, n7207, n7208, n7209, n7210, n7212, n7216, n7219, n7220,
         n7221, n7223, n7224, n7225, n7227, n7230, n7231, n7232, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7245, n7247,
         n7248, n7250, n7251, n7252, n7253, n7255, n7256, n7257, n7258, n7260,
         n7261, n7263, n7265, n7266, n7267, n7270, n7271, n7273, n7275, n7276,
         n7277, n7278, n7279, n7281, n7282, n7284, n7286, n7287, n7288, n7291,
         n7292, n7293, n7294, n7295, n7296, n7300, n7302, n7303, n7304, n7305,
         n7309, n7310, n7312, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7333, n7335, n7337,
         n7339, n7341, n7342, n7344, n7345, n7346, n7349, n7350, n7352, n7353,
         n7355, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7369, n7370, n7371, n7373, n7374, n7376, n7377, n7379,
         n7380, n7382, n7384, n7387, n7389, n7391, n7392, n7393, n7396, n7397,
         n7399, n7402, n7403, n7404, n7406, n7409, n7414, n7415, n7416, n7418,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7431, n7432, n7434,
         n7435, n7436, n7437, n7439, n7440, n7443, n7445, n7448, n7451, n7454,
         n7457, n7459, n7460, n7462, n7464, n7466, n7467, n7468, n7469, n7471,
         n7472, n7474, n7475, n7478, n7479, n7480, n7481, n7482, n7483, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7502, n7504, n7506, n7507, n7510, n7511,
         n7512, n7513, n7515, n7516, n7517, n7518, n7520, n7523, n7526, n7527,
         n7528, n7529, n7530, n7534, n7535, n7536, n7537, n7539, n7540, n7541,
         n7542, n7543, n7544, n7546, n7547, n7548, n7549, n7551, n7552, n7553,
         n7555, n7558, n7560, n7564, n7565, n7569, n7570, n7571, n7572, n7573,
         n7575, n7577, n7578, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7593, n7595, n7596, n7598, n7600, n7601, n7602,
         n7603, n7606, n7607, n7608, n7610, n7611, n7612, n7613, n7614, n7615,
         n7619, n7620, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7635, n7636, n7637, n7639, n7640, n7643, n7644, n7647,
         n7651, n7654, n7657, n7658, n7659, n7660, n7661, n7663, n7664, n7665,
         n7666, n7667, n7673, n7674, n7676, n7677, n7678, n7680, n7681, n7683,
         n7689, n7690, n7691, n7693, n7694, n7695, n7696, n7698, n7699, n7703,
         n7705, n7706, n7708, n7710, n7712, n7714, n7716, n7717, n7718, n7719,
         n7720, n7722, n7724, n7725, n7726, n7728, n7729, n7730, n7732, n7733,
         n7734, n7737, n7741, n7742, n7744, n7745, n7749, n7751, n7752, n7755,
         n7757, n7759, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7778, n7779, n7780, n7781, n7783, n7785,
         n7786, n7787, n7789, n7790, n7792, n7795, n7796, n7797, n7799, n7800,
         n7801, n7802, n7804, n7805, n7806, n7808, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7825, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7839, n7840, n7843, n7845,
         n7846, n7847, n7848, n7849, n7851, n7852, n7853, n7854, n7855, n7859,
         n7861, n7862, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7874, n7875, n7876, n7877, n7878, n7880, n7882, n7883, n7884,
         n7885, n7886, n7888, n7890, n7892, n7893, n7894, n7895, n7896, n7897,
         n7899, n7900, n7901, n7902, n7904, n7905, n7907, n7908, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7919, n7920, n7921, n7922,
         n7923, n7924, n7926, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7938, n7939, n7941, n7942, n7944, n7945, n7946, n7949, n7950,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7986,
         n7987, n7989, n7990, n7992, n7993, n7998, n7999, n8000, n8002, n8003,
         n8005, n8006, n8008, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8019, n8020, n8021, n8023, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8045, n8046, n8048, n8050, n8052, n8053, n8054, n8056, n8057,
         n8058, n8059, n8060, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8073, n8074, n8075, n8076, n8078, n8080, n8082,
         n8083, n8085, n8087, n8089, n8090, n8092, n8093, n8094, n8096, n8100,
         n8101, n8103, n8105, n8106, n8107, n8108, n8109, n8110, n8112, n8113,
         n8116, n8118, n8119, n8120, n8121, n8122, n8123, n8125, n8127, n8128,
         n8131, n8132, n8133, n8135, n8136, n8137, n8138, n8139, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8151, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8163, n8165, n8166, n8168,
         n8169, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8180, n8181,
         n8182, n8183, n8184, n8186, n8187, n8188, n8189, n8190, n8193, n8194,
         n8196, n8197, n8199, n8200, n8201, n8202, n8204, n8205, n8206, n8207,
         n8208, n8210, n8211, n8212, n8213, n8214, n8216, n8217, n8218, n8219,
         n8221, n8222, n8223, n8228, n8229, n8231, n8232, n8233, n8234, n8235,
         n8236, n8238, n8239, n8240, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8255, n8257, n8260, n8261,
         n8262, n8263, n8264, n8265, n8267, n8268, n8269, n8272, n8275, n8276,
         n8277, n8280, n8281, n8283, n8284, n8285, n8286, n8287, n8289, n8290,
         n8291, n8293, n8294, n8295, n8296, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8307, n8308, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8342, n8343, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8355, n8358, n8359, n8360, n8361, n8362, n8364,
         n8365, n8366, n8368, n8369, n8370, n8371, n8372, n8375, n8376, n8377,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8388, n8389, n8390,
         n8392, n8393, n8395, n8396, n8397, n8399, n8400, n8401, n8402, n8403,
         n8404, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8415,
         n8416, n8419, n8423, n8424, n8425, n8426, n8428, n8430, n8431, n8432,
         n8434, n8436, n8438, n8439, n8440, n8441, n8442, n8443, n8445, n8446,
         n8447, n8449, n8452, n8453, n8454, n8458, n8459, n8460, n8461, n8462,
         n8463, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8485, n8486, n8491, n8493, n8494, n8495, n8496, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8511, n8512,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8537, n8538, n8539, n8540, n8542, n8543, n8544, n8546, n8547,
         n8549, n8552, n8553, n8554, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8574,
         n8575, n8576, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8590, n8591, n8592, n8593, n8594, n8595, n8597, n8598,
         n8599, n8600, n8601, n8602, n8604, n8605, n8606, n8607, n8608, n8618,
         n8621, n8622, n8623, n8625, n8626, n8627, n8628, n8629, n8631, n8632,
         n8634, n8635, n8637, n8640, n8641, n8642, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8656, n8657, n8658,
         n8659, n8660, n8662, n8666, n8668, n8670, n8671, n8673, n8674, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8713, n8714, n8716, n8717, n8719, n8720, n8721,
         n8723, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8769, n8770, n8771, n8773, n8774, n8775, n8776, n8780, n8781, n8782,
         n8784, n8785, n8787, n8788, n8792, n8793, n8794, n8796, n8798, n8799,
         n8800, n8801, n8803, n8804, n8805, n8806, n8809, n8812, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8822, n8824, n8825, n8826, n8830,
         n8833, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8849, n8850, n8852, n8853, n8854, n8856, n8858, n8860, n8863, n8865,
         n8869, n8873, n8874, n8875, n8878, n8879, n8880, n8882, n8883, n8884,
         n8885, n8887, n8888, n8889, n8890, n8891, n8892, n8894, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8913, n8914, n8916, n8917, n8918, n8919, n8920,
         n8922, n8923, n8924, n8925, n8927, n8928, n8929, n8931, n8932, n8933,
         n8934, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8954, n8955, n8957,
         n8958, n8960, n8961, n8963, n8964, n8965, n8966, n8968, n8969, n8970,
         n8971, n8972, n8974, n8975, n8977, n8978, n8979, n8980, n8982, n8983,
         n8985, n8986, n8987, n8988, n8989, n8990, n8993, n8996, n8999, n9000,
         n9001, n9003, n9005, n9007, n9008, n9009, n9010, n9011, n9013, n9014,
         n9015, n9016, n9017, n9018, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9053, n9054, n9056, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9066, n9068, n9071, n9073, n9074, n9075, n9077,
         n9078, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9089,
         n9091, n9092, n9093, n9094, n9095, n9098, n9099, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9129, n9131, n9132, n9133, n9135, n9137, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9151, n9152, n9153, n9154, n9155, n9156, n9159, n9160, n9161, n9162,
         n9164, n9165, n9166, n9168, n9169, n9170, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9187,
         n9188, n9190, n9192, n9193, n9195, n9196, n9197, n9198, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9209, n9211, n9212, n9213,
         n9214, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9230, n9231, n9233, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9255, n9256, n9257, n9261, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9274, n9275,
         n9276, n9277, n9278, n9280, n9286, n9287, n9288, n9290, n9292, n9293,
         n9294, n9295, n9297, n9298, n9299, n9300, n9301, n9303, n9305, n9308,
         n9309, n9310, n9312, n9313, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9346, n9347, n9349, n9350, n9352, n9353, n9355, n9357,
         n9360, n9362, n9363, n9364, n9366, n9367, n9369, n9370, n9371, n9373,
         n9374, n9375, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9398, n9400, n9401, n9404, n9405, n9408, n9409, n9410, n9411, n9412,
         n9413, n9415, n9416, n9417, n9418, n9420, n9422, n9423, n9424, n9425,
         n9427, n9429, n9430, n9431, n9435, n9436, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9448, n9449, n9452, n9454, n9456,
         n9457, n9458, n9459, n9460, n9461, n9466, n9468, n9469, n9470, n9472,
         n9474, n9478, n9479, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9493, n9495, n9496, n9497, n9499, n9500,
         n9501, n9503, n9504, n9506, n9507, n9508, n9509, n9511, n9512, n9513,
         n9514, n9516, n9518, n9519, n9520, n9521, n9523, n9524, n9526, n9528,
         n9529, n9530, n9534, n9535, n9539, n9540, n9541, n9543, n9546, n9547,
         n9548, n9549, n9550, n9552, n9553, n9554, n9555, n9557, n9559, n9563,
         n9564, n9565, n9567, n9568, n9569, n9570, n9572, n9573, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9597, n9598,
         n9599, n9602, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9614, n9616, n9618, n9619, n9621, n9624, n9625, n9626, n9627,
         n9632, n9633, n9634, n9636, n9638, n9639, n9642, n9643, n9646, n9648,
         n9649, n9650, n9651, n9654, n9655, n9656, n9658, n9660, n9663, n9667,
         n9668, n9669, n9670, n9672, n9673, n9674, n9676, n9677, n9680, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9690, n9692, n9694, n9695,
         n9698, n9699, n9700, n9701, n9702, n9703, n9705, n9707, n9708, n9711,
         n9712, n9714, n9715, n9716, n9719, n9721, n9722, n9723, n9725, n9726,
         n9727, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9739, n9740,
         n9743, n9745, n9746, n9748, n9751, n9756, n9757, n9758, n9759, n9762,
         n9763, n9764, n9766, n9768, n9769, n9770, n9772, n9775, n9776, n9777,
         n9780, n9781, n9783, n9786, n9787, n9788, n9790, n9791, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9805, n9806,
         n9807, n9808, n9809, n9811, n9813, n9815, n9816, n9817, n9818, n9821,
         n9822, n9823, n9824, n9825, n9826, n9828, n9829, n9833, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9861, n9862, n9863, n9865, n9868, n9869, n9870, n9872,
         n9873, n9874, n9875, n9876, n9878, n9880, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9891, n9892, n9893, n9894, n9895, n9897,
         n9899, n9900, n9903, n9904, n9907, n9909, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9920, n9921, n9922, n9923, n9924, n9926,
         n9928, n9930, n9931, n9932, n9935, n9937, n9938, n9939, n9941, n9942,
         n9943, n9944, n9945, n9947, n9948, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9975, n9976, n9977, n9979,
         n9980, n9981, n9982, n9983, n9984, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9996, n9997, n9999, n10001, n10002,
         n10003, n10004, n10006, n10008, n10009, n10012, n10013, n10014,
         n10015, n10016, n10018, n10019, n10023, n10024, n10025, n10026,
         n10027, n10029, n10030, n10031, n10032, n10034, n10036, n10037,
         n10038, n10039, n10040, n10041, n10044, n10046, n10047, n10048,
         n10050, n10051, n10052, n10054, n10055, n10056, n10057, n10058,
         n10059, n10061, n10062, n10065, n10066, n10069, n10070, n10071,
         n10073, n10074, n10076, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10087, n10089, n10092, n10096, n10097,
         n10098, n10100, n10101, n10104, n10107, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10120,
         n10122, n10123, n10125, n10126, n10127, n10128, n10129, n10131,
         n10132, n10134, n10136, n10137, n10138, n10139, n10140, n10141,
         n10143, n10144, n10146, n10147, n10148, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10158, n10159, n10160, n10161,
         n10162, n10163, n10166, n10167, n10168, n10169, n10171, n10174,
         n10176, n10177, n10179, n10180, n10181, n10182, n10183, n10185,
         n10186, n10187, n10189, n10190, n10193, n10195, n10196, n10197,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10219, n10220, n10221, n10223, n10224, n10225, n10226,
         n10228, n10230, n10231, n10233, n10234, n10236, n10237, n10239,
         n10240, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10258,
         n10259, n10261, n10263, n10266, n10267, n10268, n10269, n10270,
         n10272, n10273, n10275, n10276, n10278, n10279, n10282, n10284,
         n10287, n10288, n10289, n10290, n10292, n10293, n10294, n10295,
         n10296, n10297, n10299, n10301, n10302, n10303, n10304, n10305,
         n10309, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10321, n10323, n10324, n10325, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10336, n10337, n10338, n10340,
         n10342, n10343, n10345, n10346, n10349, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10361, n10364,
         n10365, n10366, n10369, n10370, n10371, n10373, n10374, n10375,
         n10377, n10378, n10379, n10380, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10393, n10394,
         n10396, n10399, n10400, n10401, n10402, n10403, n10404, n10406,
         n10407, n10408, n10409, n10410, n10412, n10413, n10414, n10417,
         n10418, n10419, n10420, n10421, n10422, n10424, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10447, n10451, n10452, n10455, n10457, n10458, n10461,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10491, n10492, n10493, n10494, n10495, n10498, n10501,
         n10502, n10507, n10508, n10509, n10510, n10511, n10513, n10515,
         n10516, n10518, n10519, n10520, n10521, n10523, n10524, n10525,
         n10526, n10530, n10532, n10534, n10535, n10536, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10546, n10548, n10549,
         n10551, n10552, n10553, n10555, n10556, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10567, n10568, n10569,
         n10570, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10589, n10590, n10592, n10593, n10595, n10596, n10597, n10598,
         n10599, n10605, n10606, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10626, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10638, n10640, n10642, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10662, n10663,
         n10665, n10667, n10668, n10670, n10671, n10673, n10674, n10676,
         n10677, n10678, n10679, n10680, n10681, n10683, n10684, n10685,
         n10686, n10689, n10690, n10691, n10693, n10694, n10695, n10697,
         n10698, n10699, n10702, n10703, n10705, n10706, n10707, n10708,
         n10709, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10729,
         n10731, n10733, n10734, n10735, n10736, n10737, n10739, n10742,
         n10743, n10744, n10746, n10747, n10748, n10751, n10753, n10754,
         n10755, n10756, n10757, n10758, n10762, n10763, n10764, n10765,
         n10766, n10767, n10769, n10770, n10771, n10773, n10774, n10775,
         n10776, n10777, n10779, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10803, n10806, n10807,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10834,
         n10835, n10836, n10837, n10839, n10840, n10841, n10842, n10845,
         n10846, n10847, n10848, n10850, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10862, n10863, n10864, n10866,
         n10867, n10868, n10869, n10870, n10872, n10874, n10875, n10876,
         n10878, n10882, n10883, n10884, n10885, n10887, n10888, n10889,
         n10890, n10891, n10893, n10894, n10896, n10897, n10898, n10899,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10910, n10913, n10914, n10915, n10918, n10920, n10924, n10925,
         n10926, n10928, n10929, n10930, n10931, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10946, n10949,
         n10953, n10955, n10957, n10959, n10961, n10962, n10963, n10965,
         n10966, n10967, n10969, n10970, n10971, n10972, n10973, n10974,
         n10976, n10977, n10978, n10979, n10980, n10982, n10983, n10984,
         n10986, n10987, n10988, n10989, n10992, n10996, n10997, n10998,
         n10999, n11001, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11012, n11013, n11015, n11016, n11017, n11018,
         n11020, n11022, n11024, n11025, n11026, n11028, n11030, n11031,
         n11032, n11033, n11034, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11046, n11047, n11048, n11050,
         n11053, n11054, n11055, n11056, n11057, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11072, n11074,
         n11075, n11076, n11077, n11081, n11082, n11083, n11084, n11087,
         n11088, n11089, n11090, n11091, n11092, n11094, n11095, n11097,
         n11098, n11099, n11102, n11103, n11104, n11105, n11108, n11111,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11136, n11137, n11138, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11180, n11181, n11182, n11183, n11185, n11186, n11187, n11188,
         n11189, n11190, n11192, n11194, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11207, n11208, n11210, n11211, n11213,
         n11214, n11215, n11217, n11218, n11219, n11220, n11222, n11224,
         n11225, n11226, n11227, n11230, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11243, n11245, n11247,
         n11248, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11260, n11261, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11283, n11284, n11286, n11288,
         n11289, n11290, n11291, n11292, n11293, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11321, n11322,
         n11323, n11325, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11339, n11342, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11353, n11354,
         n11355, n11356, n11358, n11361, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11382, n11383, n11384, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11394, n11395, n11397,
         n11398, n11399, n11401, n11402, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11415, n11416,
         n11417, n11418, n11419, n11421, n11423, n11424, n11425, n11428,
         n11429, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11446, n11448,
         n11449, n11451, n11452, n11453, n11455, n11456, n11458, n11459,
         n11461, n11462, n11463, n11464, n11465, n11467, n11468, n11469,
         n11470, n11472, n11473, n11474, n11475, n11476, n11477, n11479,
         n11481, n11482, n11484, n11485, n11486, n11487, n11488, n11490,
         n11491, n11492, n11494, n11495, n11496, n11497, n11498, n11500,
         n11501, n11502, n11503, n11506, n11507, n11508, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11525, n11526, n11528, n11529, n11530,
         n11533, n11534, n11536, n11541, n11542, n11543, n11544, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11562, n11563, n11564,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11581, n11582, n11583, n11584, n11585,
         n11586, n11588, n11589, n11590, n11591, n11594, n11595, n11596,
         n11597, n11598, n11600, n11601, n11602, n11603, n11605, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11620, n11621, n11622, n11623, n11624, n11625, n11627, n11628,
         n11630, n11631, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11641, n11642, n11643, n11644, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11657, n11658, n11659,
         n11661, n11663, n11664, n11665, n11667, n11668, n11669, n11671,
         n11672, n11673, n11674, n11676, n11677, n11678, n11679, n11680,
         n11682, n11683, n11684, n11687, n11688, n11689, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11717, n11718, n11719, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11732,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11742,
         n11743, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11762, n11763, n11764, n11765, n11767, n11768, n11769, n11770,
         n11771, n11773, n11776, n11777, n11778, n11779, n11780, n11782,
         n11783, n11784, n11785, n11787, n11788, n11789, n11790, n11791,
         n11793, n11794, n11795, n11796, n11797, n11800, n11803, n11805,
         n11806, n11807, n11809, n11810, n11814, n11818, n11820, n11822,
         n11823, n11826, n11828, n11830, n11831, n11833, n11834, n11835,
         n11838, n11842, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11858, n11859,
         n11860, n11861, n11864, n11866, n11867, n11868, n11869, n11870,
         n11871, n11873, n11874, n11875, n11876, n11877, n11878, n11880,
         n11881, n11882, n11883, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11893, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11910, n11911, n11912, n11913, n11914, n11916, n11917,
         n11918, n11919, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11935, n11937, n11938, n11939, n11940, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11950, n11951, n11952,
         n11954, n11956, n11957, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11972, n11973,
         n11974, n11975, n11976, n11977, n11980, n11981, n11984, n11985,
         n11986, n11987, n11989, n11994, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12008, n12009, n12011, n12012,
         n12014, n12015, n12016, n12017, n12018, n12020, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12036, n12038, n12039, n12040, n12044, n12045,
         n12046, n12049, n12050, n12053, n12054, n12055, n12056, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12069,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12083, n12084, n12085, n12086, n12090, n12091,
         n12093, n12094, n12096, n12097, n12100, n12101, n12102, n12103,
         n12104, n12105, n12107, n12108, n12109, n12111, n12112, n12113,
         n12114, n12115, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12130, n12131, n12132, n12133, n12138, n12139,
         n12141, n12142, n12144, n12145, n12146, n12148, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12159, n12160,
         n12161, n12162, n12163, n12165, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12183, n12184, n12185, n12187, n12189,
         n12191, n12192, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12212, n12213, n12214, n12215, n12218, n12220, n12221, n12225,
         n12227, n12228, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12242, n12243, n12244,
         n12245, n12246, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12265, n12266, n12267, n12268, n12269, n12272, n12273,
         n12275, n12276, n12277, n12279, n12282, n12283, n12286, n12287,
         n12288, n12289, n12290, n12293, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12306, n12307, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12336, n12337, n12339, n12340, n12341, n12342, n12343, n12345,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12360, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12377, n12378, n12379, n12381, n12382, n12383, n12385,
         n12387, n12388, n12391, n12392, n12393, n12394, n12396, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12420, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12435, n12437, n12438, n12439, n12441, n12442, n12443,
         n12446, n12447, n12448, n12449, n12450, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12460, n12461, n12462, n12463,
         n12464, n12466, n12468, n12469, n12470, n12471, n12472, n12473,
         n12475, n12477, n12478, n12479, n12480, n12481, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12497, n12498, n12499, n12500, n12503, n12504, n12505,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12515,
         n12516, n12517, n12518, n12519, n12520, n12522, n12523, n12524,
         n12525, n12526, n12527, n12529, n12531, n12533, n12534, n12535,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12551, n12552, n12553,
         n12556, n12557, n12558, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12572, n12574,
         n12575, n12576, n12578, n12579, n12580, n12586, n12587, n12588,
         n12590, n12592, n12593, n12594, n12597, n12598, n12599, n12601,
         n12604, n12605, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12616, n12617, n12618, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12638, n12639, n12641, n12642, n12643, n12644,
         n12646, n12649, n12650, n12651, n12653, n12654, n12655, n12657,
         n12659, n12660, n12661, n12663, n12664, n12665, n12667, n12669,
         n12670, n12671, n12672, n12673, n12675, n12676, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12689, n12690, n12691,
         n12692, n12694, n12696, n12697, n12698, n12699, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12717, n12718, n12721, n12722,
         n12723, n12726, n12727, n12728, n12729, n12730, n12732, n12733,
         n12735, n12736, n12737, n12738, n12741, n12744, n12745, n12746,
         n12748, n12749, n12751, n12752, n12754, n12755, n12756, n12758,
         n12759, n12760, n12762, n12763, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12775, n12776, n12778, n12779,
         n12780, n12782, n12784, n12785, n12787, n12788, n12790, n12793,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12824, n12825, n12826, n12828, n12829, n12830,
         n12832, n12833, n12834, n12835, n12836, n12838, n12839, n12840,
         n12842, n12844, n12846, n12847, n12848, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12865, n12866, n12869, n12870, n12871,
         n12876, n12878, n12879, n12880, n12882, n12883, n12884, n12885,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12908, n12909, n12910, n12912, n12914, n12915, n12916, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12930, n12931, n12933, n12934, n12935, n12936, n12939,
         n12940, n12941, n12942, n12943, n12944, n12946, n12947, n12950,
         n12951, n12952, n12953, n12954, n12955, n12960, n12961, n12964,
         n12966, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12978, n12979, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12999, n13000, n13001, n13002, n13004,
         n13005, n13006, n13008, n13009, n13010, n13012, n13013, n13014,
         n13015, n13016, n13018, n13019, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13033, n13034, n13035,
         n13036, n13038, n13039, n13040, n13042, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13052, n13053, n13054, n13055,
         n13056, n13059, n13060, n13061, n13062, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13081, n13082, n13083, n13085, n13087,
         n13088, n13090, n13091, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13118, n13119, n13121, n13123, n13124, n13127, n13128,
         n13129, n13131, n13132, n13133, n13134, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13147, n13149,
         n13150, n13151, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13161, n13163, n13164, n13165, n13166, n13167, n13168,
         n13170, n13171, n13172, n13174, n13176, n13177, n13178, n13179,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13199, n13200, n13201, n13202, n13205, n13206, n13207,
         n13208, n13210, n13211, n13212, n13213, n13214, n13215, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13226,
         n13227, n13228, n13229, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13254, n13255, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13266, n13267, n13268, n13270, n13273, n13274,
         n13275, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13298, n13300, n13301, n13302,
         n13304, n13305, n13306, n13308, n13310, n13311, n13312, n13313,
         n13315, n13316, n13317, n13318, n13320, n13321, n13322, n13323,
         n13324, n13326, n13327, n13329, n13332, n13333, n13334, n13335,
         n13336, n13337, n13339, n13340, n13342, n13345, n13348, n13349,
         n13350, n13351, n13352, n13354, n13356, n13358, n13359, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13378, n13379,
         n13381, n13383, n13384, n13386, n13387, n13388, n13389, n13391,
         n13392, n13393, n13395, n13397, n13398, n13400, n13401, n13403,
         n13404, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13417, n13419, n13420, n13421, n13422,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13448, n13450, n13451, n13453,
         n13454, n13455, n13457, n13458, n13460, n13461, n13462, n13465,
         n13466, n13467, n13468, n13469, n13471, n13472, n13473, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13483, n13484,
         n13485, n13487, n13488, n13489, n13491, n13492, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13508, n13510, n13512, n13513, n13514, n13515, n13516,
         n13518, n13519, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13530, n13531, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13542, n13543, n13544, n13545,
         n13547, n13548, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13563, n13564,
         n13565, n13566, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13591, n13592,
         n13593, n13594, n13595, n13596, n13598, n13599, n13600, n13601,
         n13602, n13603, n13605, n13606, n13607, n13608, n13609, n13610,
         n13614, n13615, n13616, n13617, n13618, n13620, n13621, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13644, n13645, n13646, n13649, n13650,
         n13652, n13653, n13654, n13656, n13657, n13658, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13688, n13689, n13690, n13691,
         n13692, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13716, n13717, n13718,
         n13719, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13738, n13739, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13761, n13762,
         n13763, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13782,
         n13784, n13785, n13786, n13787, n13788, n13789, n13791, n13792,
         n13793, n13794, n13797, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13811, n13814,
         n13815, n13817, n13818, n13820, n13823, n13824, n13825, n13826,
         n13827, n13829, n13830, n13831, n13832, n13833, n13834, n13837,
         n13839, n13840, n13842, n13843, n13844, n13845, n13846, n13847,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13858, n13859, n13860, n13861, n13862, n13869, n13870, n13871,
         n13872, n13873, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13883, n13884, n13885, n13886, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13899, n13900, n13901,
         n13903, n13904, n13905, n13906, n13907, n13909, n13910, n13911,
         n13912, n13913, n13914, n13917, n13918, n13919, n13920, n13922,
         n13926, n13927, n13928, n13931, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13942, n13943, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13954, n13955, n13956,
         n13959, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13969, n13970, n13971, n13973, n13976, n13977, n13978, n13980,
         n13981, n13982, n13983, n13984, n13986, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n14000, n14001, n14002, n14003, n14004, n14006, n14007, n14008,
         n14009, n14011, n14012, n14015, n14016, n14017, n14020, n14022,
         n14023, n14024, n14025, n14027, n14028, n14030, n14031, n14034,
         n14035, n14036, n14037, n14038, n14039, n14041, n14043, n14045,
         n14046, n14049, n14050, n14051, n14052, n14053, n14056, n14057,
         n14058, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14069, n14072, n14073, n14075, n14076, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14088, n14089, n14091,
         n14093, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14109, n14110, n14112, n14113,
         n14115, n14116, n14117, n14118, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14139, n14140, n14143, n14144,
         n14145, n14146, n14147, n14148, n14150, n14151, n14152, n14153,
         n14154, n14156, n14157, n14158, n14160, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14173, n14174,
         n14176, n14178, n14179, n14181, n14183, n14184, n14186, n14187,
         n14188, n14189, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14203, n14205, n14206,
         n14209, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14224, n14226, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14237,
         n14239, n14241, n14244, n14245, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14257, n14258, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14269, n14270,
         n14271, n14272, n14273, n14275, n14276, n14277, n14278, n14280,
         n14281, n14282, n14283, n14285, n14286, n14287, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14297, n14300, n14302,
         n14303, n14304, n14305, n14306, n14307, n14309, n14311, n14312,
         n14316, n14318, n14319, n14322, n14323, n14325, n14326, n14327,
         n14330, n14331, n14332, n14333, n14337, n14338, n14339, n14343,
         n14345, n14346, n14347, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14359, n14361, n14362, n14363, n14364, n14365,
         n14367, n14369, n14371, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14385, n14386,
         n14387, n14388, n14389, n14390, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14417, n14418, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14431,
         n14432, n14433, n14435, n14436, n14437, n14438, n14439, n14440,
         n14442, n14443, n14444, n14448, n14449, n14450, n14451, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14469, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14511, n14512, n14513, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14529, n14530, n14532, n14533, n14534, n14535, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14546, n14548,
         n14549, n14551, n14553, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14568, n14569,
         n14571, n14572, n14573, n14576, n14577, n14578, n14579, n14581,
         n14582, n14583, n14585, n14586, n14587, n14588, n14589, n14590,
         n14592, n14593, n14594, n14596, n14597, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14608, n14609, n14610, n14613,
         n14614, n14615, n14617, n14618, n14619, n14621, n14622, n14623,
         n14625, n14626, n14628, n14630, n14631, n14632, n14634, n14635,
         n14636, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14648, n14649, n14650, n14651, n14652, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14662, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14672, n14673,
         n14675, n14677, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14689, n14691, n14692, n14693, n14694,
         n14695, n14696, n14699, n14701, n14703, n14704, n14705, n14708,
         n14709, n14712, n14713, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14724, n14725, n14729, n14732, n14734,
         n14735, n14736, n14737, n14738, n14739, n14742, n14743, n14744,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14762, n14764,
         n14765, n14766, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14787, n14788, n14789, n14790, n14791, n14793, n14794,
         n14795, n14796, n14797, n14798, n14800, n14801, n14802, n14804,
         n14805, n14807, n14808, n14810, n14811, n14813, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14833, n14834,
         n14835, n14837, n14838, n14839, n14840, n14843, n14844, n14845,
         n14846, n14848, n14850, n14851, n14854, n14855, n14856, n14857,
         n14858, n14859, n14861, n14862, n14866, n14867, n14868, n14869,
         n14872, n14873, n14874, n14875, n14876, n14877, n14879, n14880,
         n14881, n14882, n14887, n14888, n14890, n14891, n14892, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14907, n14908, n14909, n14910, n14911, n14912,
         n14914, n14915, n14916, n14919, n14920, n14921, n14922, n14924,
         n14925, n14926, n14927, n14928, n14929, n14931, n14933, n14934,
         n14935, n14936, n14939, n14940, n14941, n14945, n14946, n14947,
         n14949, n14952, n14953, n14955, n14956, n14957, n14962, n14966,
         n14967, n14968, n14969, n14970, n14971, n14974, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14993, n14994, n14995,
         n14997, n14998, n14999, n15001, n15003, n15004, n15005, n15006,
         n15007, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15056, n15058, n15062, n15063, n15068,
         n15069, n15071, n15072, n15073, n15074, n15075, n15077, n15078,
         n15079, n15080, n15081, n15082, n15084, n15085, n15087, n15089,
         n15090, n15091, n15093, n15094, n15096, n15097, n15099, n15102,
         n15109, n15110, n15112, n15113, n15114, n15115, n15118, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15131, n15132, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15145, n15146, n15148, n15149,
         n15151, n15152, n15153, n15155, n15156, n15157, n15158, n15159,
         n15160, n15162, n15163, n15164, n15165, n15168, n15169, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15180,
         n15181, n15183, n15184, n15186, n15187, n15189, n15193, n15194,
         n15195, n15196, n15197, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15218, n15219, n15220, n15222,
         n15223, n15224, n15226, n15227, n15229, n15230, n15232, n15233,
         n15235, n15237, n15238, n15239, n15240, n15242, n15243, n15245,
         n15246, n15248, n15249, n15250, n15251, n15254, n15256, n15257,
         n15258, n15259, n15261, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15280, n15281, n15282, n15283, n15284, n15286, n15287, n15288,
         n15289, n15290, n15292, n15293, n15294, n15295, n15296, n15298,
         n15299, n15301, n15303, n15304, n15305, n15307, n15308, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15319,
         n15320, n15321, n15323, n15324, n15325, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15336, n15337, n15338,
         n15339, n15340, n15341, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15364, n15365, n15368,
         n15369, n15370, n15371, n15372, n15373, n15375, n15376, n15377,
         n15378, n15380, n15381, n15382, n15384, n15385, n15386, n15388,
         n15389, n15391, n15393, n15394, n15395, n15398, n15400, n15401,
         n15404, n15405, n15406, n15410, n15411, n15412, n15413, n15414,
         n15419, n15420, n15421, n15422, n15423, n15424, n15426, n15427,
         n15429, n15430, n15432, n15433, n15434, n15435, n15436, n15437,
         n15439, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15455, n15456,
         n15457, n15458, n15459, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15471, n15473, n15476, n15477, n15480,
         n15481, n15482, n15483, n15485, n15487, n15488, n15490, n15491,
         n15492, n15493, n15495, n15496, n15497, n15499, n15500, n15502,
         n15503, n15507, n15508, n15509, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15534, n15535, n15540, n15541, n15542, n15543, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15558, n15559, n15560, n15562, n15564, n15565, n15566,
         n15568, n15569, n15570, n15571, n15572, n15573, n15575, n15577,
         n15579, n15580, n15581, n15583, n15584, n15585, n15586, n15588,
         n15589, n15591, n15592, n15594, n15595, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15607, n15608,
         n15609, n15610, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15629, n15630, n15631, n15633, n15634, n15635, n15638,
         n15641, n15642, n15643, n15644, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15656, n15660, n15663, n15664,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15676, n15677, n15678, n15679, n15681, n15682, n15684, n15685,
         n15686, n15688, n15689, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15700, n15701, n15702, n15703, n15704, n15706,
         n15707, n15708, n15709, n15710, n15712, n15713, n15715, n15716,
         n15717, n15718, n15719, n15721, n15722, n15723, n15726, n15727,
         n15728, n15729, n15730, n15733, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15745, n15748, n15750,
         n15751, n15752, n15753, n15754, n15755, n15757, n15758, n15761,
         n15762, n15763, n15765, n15767, n15768, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15779, n15780, n15782,
         n15785, n15787, n15788, n15789, n15790, n15791, n15792, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15808, n15809, n15810, n15811,
         n15812, n15814, n15816, n15817, n15818, n15819, n15821, n15822,
         n15823, n15824, n15825, n15826, n15828, n15829, n15831, n15832,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15844, n15846, n15848, n15849, n15850, n15852, n15853,
         n15854, n15855, n15857, n15858, n15859, n15860, n15861, n15862,
         n15864, n15865, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15888, n15890, n15891, n15892, n15893,
         n15894, n15896, n15897, n15898, n15899, n15903, n15904, n15907,
         n15909, n15910, n15911, n15912, n15913, n15915, n15916, n15917,
         n15918, n15919, n15922, n15924, n15925, n15926, n15928, n15929,
         n15930, n15932, n15933, n15935, n15936, n15937, n15938, n15940,
         n15941, n15943, n15945, n15946, n15947, n15949, n15951, n15952,
         n15953, n15955, n15956, n15957, n15958, n15959, n15960, n15963,
         n15964, n15966, n15967, n15968, n15969, n15971, n15972, n15973,
         n15974, n15975, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15991, n15992,
         n15993, n15994, n15995, n15996, n15998, n15999, n16000, n16004,
         n16006, n16007, n16009, n16010, n16013, n16014, n16015, n16016,
         n16017, n16019, n16021, n16022, n16024, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16038, n16039, n16040, n16041, n16042, n16043, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16091,
         n16093, n16094, n16095, n16096, n16097, n16098, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16113, n16114, n16115, n16116, n16117, n16118, n16121, n16123,
         n16124, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16137, n16138, n16140, n16141, n16144,
         n16146, n16147, n16149, n16150, n16151, n16153, n16154, n16158,
         n16159, n16160, n16161, n16162, n16163, n16165, n16167, n16168,
         n16169, n16170, n16171, n16173, n16174, n16175, n16177, n16179,
         n16180, n16181, n16182, n16183, n16184, n16186, n16187, n16190,
         n16191, n16192, n16193, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16206, n16208, n16209, n16210,
         n16211, n16213, n16216, n16217, n16218, n16220, n16221, n16222,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16252, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16275, n16277, n16278,
         n16281, n16282, n16283, n16284, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16298, n16299,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16315, n16316, n16317,
         n16318, n16320, n16321, n16324, n16325, n16327, n16328, n16332,
         n16333, n16334, n16336, n16337, n16338, n16339, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16350, n16351, n16353,
         n16355, n16356, n16357, n16358, n16359, n16360, n16362, n16363,
         n16364, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16385, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16397, n16398, n16400, n16401, n16402,
         n16403, n16406, n16407, n16410, n16411, n16412, n16416, n16417,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16427,
         n16428, n16430, n16431, n16432, n16435, n16439, n16440, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16452,
         n16453, n16454, n16455, n16456, n16458, n16459, n16460, n16461,
         n16463, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16482, n16484, n16487, n16488, n16489, n16490, n16492, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16502, n16503,
         n16505, n16508, n16510, n16511, n16513, n16514, n16516, n16517,
         n16520, n16522, n16523, n16524, n16525, n16526, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16539, n16540, n16541, n16542, n16543, n16544, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16565,
         n16566, n16567, n16569, n16570, n16573, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16587, n16589, n16590, n16591, n16593, n16595, n16596, n16597,
         n16598, n16599, n16601, n16604, n16605, n16606, n16607, n16610,
         n16612, n16613, n16615, n16617, n16618, n16619, n16621, n16623,
         n16624, n16625, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16647, n16648, n16650, n16651,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16663, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16676, n16677, n16678, n16679, n16682,
         n16683, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16704, n16705, n16706, n16707, n16708, n16709, n16712,
         n16713, n16715, n16716, n16720, n16721, n16722, n16723, n16726,
         n16728, n16729, n16731, n16732, n16733, n16735, n16736, n16737,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16749, n16750, n16751, n16753, n16755, n16757, n16758,
         n16759, n16760, n16762, n16763, n16765, n16766, n16767, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16781, n16782, n16783, n16785, n16786, n16787, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16809,
         n16810, n16813, n16814, n16815, n16816, n16819, n16820, n16825,
         n16828, n16829, n16830, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16845,
         n16847, n16848, n16849, n16851, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16863, n16864, n16867,
         n16868, n16869, n16871, n16873, n16874, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16886, n16887,
         n16888, n16889, n16890, n16892, n16893, n16896, n16897, n16898,
         n16900, n16901, n16902, n16903, n16904, n16905, n16907, n16908,
         n16911, n16912, n16917, n16918, n16919, n16920, n16921, n16922,
         n16924, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16939, n16941, n16942, n16945, n16946, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16960, n16961, n16962, n16963, n16964, n16966, n16967, n16968,
         n16970, n16971, n16972, n16975, n16976, n16977, n16982, n16985,
         n16987, n16988, n16989, n16990, n16992, n16993, n16994, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17006,
         n17007, n17008, n17009, n17013, n17017, n17018, n17020, n17021,
         n17022, n17023, n17024, n17025, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17037, n17038, n17039,
         n17040, n17041, n17043, n17045, n17047, n17048, n17051, n17055,
         n17057, n17058, n17060, n17062, n17063, n17064, n17066, n17067,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17080,
         n17081, n17083, n17084, n17085, n17086, n17087, n17089, n17090,
         n17091, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17110, n17112, n17113, n17114, n17115, n17117, n17118,
         n17119, n17120, n17121, n17122, n17124, n17125, n17126, n17127,
         n17128, n17129, n17131, n17132, n17134, n17136, n17137, n17138,
         n17139, n17140, n17142, n17143, n17144, n17145, n17147, n17148,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17158,
         n17159, n17160, n17161, n17163, n17166, n17167, n17168, n17169,
         n17171, n17172, n17173, n17176, n17177, n17178, n17179, n17180,
         n17182, n17183, n17184, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17197, n17198, n17201, n17202,
         n17205, n17207, n17209, n17210, n17211, n17212, n17213, n17214,
         n17217, n17219, n17220, n17221, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17231, n17232, n17233, n17234, n17236,
         n17237, n17238, n17240, n17242, n17243, n17245, n17246, n17248,
         n17249, n17250, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17301, n17302, n17303,
         n17304, n17305, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17325, n17326, n17328, n17329, n17331, n17332,
         n17333, n17334, n17335, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17346, n17347, n17348, n17349, n17350, n17351,
         n17353, n17354, n17356, n17357, n17358, n17359, n17360, n17361,
         n17363, n17364, n17365, n17366, n17368, n17369, n17371, n17372,
         n17373, n17374, n17377, n17378, n17381, n17382, n17383, n17388,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17415,
         n17416, n17417, n17418, n17420, n17422, n17423, n17424, n17425,
         n17426, n17428, n17429, n17430, n17433, n17435, n17436, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17480, n17482, n17483, n17484,
         n17485, n17486, n17487, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17508, n17509, n17511, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17544, n17546, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17583, n17584, n17586, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17612, n17613,
         n17615, n17616, n17617, n17618, n17621, n17623, n17624, n17627,
         n17628, n17630, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17650, n17651, n17653, n17655, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17668, n17669,
         n17673, n17674, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17691, n17692,
         n17693, n17696, n17697, n17698, n17699, n17700, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17723, n17724, n17725, n17726, n17727, n17730, n17731, n17732,
         n17735, n17737, n17738, n17739, n17740, n17742, n17744, n17745,
         n17747, n17748, n17750, n17751, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17763, n17764, n17765, n17767,
         n17768, n17770, n17771, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17781, n17782, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17797, n17798, n17799, n17800, n17801, n17803, n17804, n17806,
         n17810, n17811, n17812, n17813, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17823, n17824, n17826, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17841, n17842, n17844, n17847, n17848, n17849, n17850,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17871, n17872, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17882, n17884, n17885, n17886, n17887, n17888,
         n17890, n17891, n17893, n17894, n17896, n17897, n17898, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17915, n17916, n17917, n17918,
         n17920, n17921, n17922, n17923, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17951, n17952, n17954, n17955, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18012, n18013, n18014, n18015,
         n18017, n18018, n18019, n18020, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18031, n18032, n18034, n18035, n18036,
         n18037, n18038, n18039, n18041, n18042, n18043, n18044, n18047,
         n18048, n18049, n18050, n18051, n18054, n18055, n18056, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18070, n18071, n18072, n18073, n18074, n18075, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18094, n18095, n18096, n18098,
         n18101, n18103, n18104, n18106, n18107, n18108, n18109, n18110,
         n18112, n18113, n18114, n18115, n18116, n18120, n18121, n18122,
         n18123, n18124, n18125, n18127, n18129, n18131, n18133, n18134,
         n18135, n18137, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18152, n18153, n18155,
         n18156, n18157, n18159, n18160, n18162, n18163, n18164, n18166,
         n18168, n18170, n18171, n18172, n18174, n18175, n18176, n18178,
         n18179, n18180, n18182, n18183, n18184, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18204, n18205, n18207,
         n18208, n18209, n18210, n18211, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18246, n18249, n18250, n18251, n18253,
         n18255, n18256, n18257, n18259, n18261, n18263, n18264, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18276, n18277, n18278, n18279, n18281, n18282, n18283, n18284,
         n18288, n18289, n18290, n18291, n18293, n18294, n18295, n18296,
         n18298, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18319, n18320, n18322, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18335, n18338, n18339,
         n18340, n18341, n18342, n18345, n18346, n18347, n18348, n18349,
         n18350, n18352, n18353, n18354, n18357, n18359, n18360, n18362,
         n18363, n18364, n18365, n18366, n18367, n18369, n18370, n18371,
         n18372, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18386, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18398, n18399, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18410,
         n18412, n18413, n18415, n18416, n18417, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18436, n18438, n18439, n18440,
         n18445, n18446, n18447, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18487, n18488,
         n18489, n18490, n18491, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18515, n18516,
         n18518, n18519, n18520, n18522, n18523, n18524, n18525, n18526,
         n18527, n18529, n18530, n18532, n18534, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18554, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18582, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18597, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18608, n18609,
         n18610, n18611, n18612, n18615, n18616, n18617, n18618, n18619,
         n18620, n18622, n18623, n18624, n18625, n18626, n18628, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18640,
         n18641, n18642, n18643, n18645, n18647, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18665, n18667, n18668, n18669, n18670,
         n18671, n18673, n18674, n18675, n18679, n18680, n18681, n18682,
         n18683, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18694, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18725, n18726, n18728, n18729, n18730,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18755, n18757, n18758, n18759,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18773, n18774, n18776, n18777, n18778, n18780,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18790,
         n18792, n18793, n18794, n18795, n18796, n18797, n18800, n18801,
         n18803, n18804, n18806, n18807, n18808, n18809, n18810, n18811,
         n18813, n18814, n18815, n18816, n18817, n18819, n18822, n18825,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18836, n18837, n18838, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18869, n18870, n18871,
         n18872, n18873, n18875, n18876, n18877, n18879, n18880, n18883,
         n18884, n18886, n18887, n18888, n18889, n18890, n18891, n18893,
         n18894, n18896, n18897, n18898, n18900, n18901, n18902, n18903,
         n18904, n18905, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18917, n18918, n18920, n18921, n18922,
         n18923, n18924, n18926, n18927, n18928, n18929, n18930, n18931,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18950,
         n18951, n18952, n18953, n18954, n18956, n18958, n18959, n18960,
         n18961, n18962, n18966, n18967, n18968, n18969, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18979, n18980, n18981,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19005, n19006, n19007, n19008,
         n19009, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19024, n19025, n19026,
         n19027, n19028, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19041, n19042, n19043, n19045,
         n19047, n19048, n19050, n19051, n19052, n19053, n19054, n19055,
         n19059, n19060, n19061, n19062, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19077, n19078, n19080, n19081, n19082, n19083, n19084, n19085,
         n19088, n19089, n19090, n19091, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19108, n19109, n19111, n19112, n19113, n19115, n19118,
         n19119, n19120, n19121, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19142, n19143, n19145,
         n19146, n19147, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19175,
         n19177, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19191, n19193, n19194, n19195, n19196,
         n19197, n19198, n19200, n19201, n19202, n19203, n19204, n19206,
         n19207, n19209, n19210, n19211, n19213, n19214, n19215, n19216,
         n19217, n19218, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19240, n19241, n19242, n19244,
         n19246, n19249, n19250, n19252, n19253, n19254, n19255, n19257,
         n19258, n19259, n19260, n19261, n19262, n19264, n19266, n19268,
         n19270, n19271, n19272, n19274, n19276, n19277, n19278, n19279,
         n19280, n19281, n19283, n19284, n19285, n19287, n19288, n19289,
         n19290, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19300, n19302, n19303, n19304, n19305, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19316, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19331, n19332, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19358, n19359, n19360, n19361, n19362, n19364, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19379, n19380, n19381, n19382, n19384, n19385,
         n19387, n19388, n19389, n19391, n19392, n19393, n19395, n19396,
         n19397, n19398, n19400, n19401, n19402, n19403, n19404, n19405,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19428, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19438, n19439, n19440, n19442, n19443,
         n19444, n19445, n19446, n19448, n19449, n19450, n19452, n19453,
         n19454, n19455, n19456, n19458, n19459, n19460, n19463, n19464,
         n19465, n19466, n19467, n19469, n19470, n19471, n19472, n19473,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19486, n19488, n19490, n19492, n19493, n19495,
         n19496, n19497, n19498, n19499, n19501, n19503, n19504, n19505,
         n19507, n19508, n19511, n19513, n19514, n19515, n19516, n19517,
         n19518, n19521, n19524, n19525, n19527, n19528, n19529, n19530,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19557, n19559,
         n19560, n19561, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19579, n19580, n19581, n19582, n19583, n19584, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19599, n19600, n19601, n19604, n19605,
         n19606, n19608, n19609, n19610, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19627, n19629, n19630, n19631, n19632, n19633, n19636,
         n19637, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19704, n19706, n19707, n19708,
         n19709, n19712, n19713, n19714, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19754,
         n19755, n19756, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19777, n19778, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19788, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19827, n19828, n19829, n19830, n19831, n19833, n19835, n19836,
         n19837, n19838, n19839, n19840, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19855, n19856,
         n19857, n19859, n19860, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19913, n19914, n19915, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19971,
         n19972, n19973, n19975, n19976, n19978, n19979, n19980, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20002, n20003, n20004, n20006, n20007, n20008,
         n20010, n20013, n20016, n20018, n20019, n20020, n20021, n20022,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20041, n20042, n20043, n20044, n20045, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20056, n20057, n20058, n20059,
         n20061, n20062, n20063, n20064, n20065, n20066, n20068, n20069,
         n20070, n20074, n20076, n20077, n20078, n20080, n20082, n20083,
         n20084, n20085, n20087, n20088, n20089, n20090, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20105, n20107, n20108, n20109, n20111, n20112,
         n20113, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20125, n20126, n20128, n20129, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20139, n20140, n20143, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20164,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20180, n20184, n20185, n20186,
         n20187, n20188, n20190, n20191, n20194, n20196, n20197, n20198,
         n20199, n20200, n20201, n20203, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20216, n20217,
         n20219, n20221, n20222, n20223, n20225, n20226, n20227, n20229,
         n20230, n20232, n20234, n20235, n20236, n20237, n20238, n20239,
         n20241, n20242, n20243, n20244, n20245, n20250, n20251, n20254,
         n20255, n20256, n20257, n20260, n20261, n20262, n20263, n20264,
         n20266, n20267, n20268, n20270, n20274, n20276, n20277, n20278,
         n20279, n20280, n20282, n20284, n20286, n20287, n20288, n20289,
         n20290, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20316, n20317,
         n20319, n20321, n20322, n20323, n20324, n20325, n20326, n20328,
         n20329, n20330, n20331, n20332, n20333, n20335, n20336, n20337,
         n20339, n20340, n20341, n20342, n20343, n20344, n20346, n20347,
         n20348, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20361, n20362, n20363, n20364, n20365,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20381, n20384, n20386, n20387,
         n20388, n20389, n20391, n20392, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20414, n20416,
         n20418, n20419, n20420, n20421, n20423, n20424, n20425, n20426,
         n20427, n20429, n20430, n20431, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20460, n20462,
         n20463, n20464, n20465, n20468, n20469, n20470, n20472, n20473,
         n20474, n20476, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20522, n20524, n20525, n20526, n20528, n20530, n20531,
         n20533, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20544, n20545, n20546, n20547, n20549, n20550, n20551, n20554,
         n20555, n20559, n20560, n20561, n20562, n20564, n20565, n20566,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20600, n20601, n20602, n20604, n20605,
         n20607, n20608, n20609, n20611, n20612, n20613, n20614, n20615,
         n20616, n20618, n20619, n20620, n20621, n20622, n20623, n20625,
         n20626, n20627, n20628, n20629, n20632, n20634, n20635, n20636,
         n20637, n20638, n20639, n20641, n20642, n20643, n20644, n20646,
         n20648, n20649, n20651, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20665, n20666,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20701, n20702,
         n20703, n20704, n20706, n20707, n20708, n20709, n20713, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20723, n20724,
         n20725, n20726, n20727, n20728, n20730, n20731, n20732, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20743,
         n20744, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20756, n20758, n20759, n20761, n20762, n20764,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20787, n20788, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20813, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20835, n20836, n20838, n20839, n20840,
         n20841, n20843, n20844, n20845, n20846, n20849, n20850, n20851,
         n20852, n20855, n20856, n20858, n20859, n20860, n20862, n20863,
         n20864, n20865, n20866, n20867, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20901, n20903, n20907, n20910, n20911, n20912, n20914, n20915,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20936, n20939, n20941,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20951,
         n20952, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20984, n20986, n20987,
         n20988, n20989, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21017, n21018, n21019, n21020, n21021, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21071, n21072, n21073,
         n21074, n21076, n21077, n21079, n21080, n21081, n21084, n21085,
         n21086, n21087, n21090, n21091, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21103, n21104, n21105,
         n21108, n21109, n21110, n21111, n21114, n21116, n21117, n21118,
         n21119, n21120, n21121, n21124, n21125, n21126, n21127, n21128,
         n21130, n21132, n21133, n21134, n21135, n21136, n21137, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21152, n21154, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21174, n21176, n21177,
         n21181, n21182, n21184, n21186, n21187, n21188, n21190, n21191,
         n21192, n21195, n21196, n21197, n21198, n21201, n21202, n21204,
         n21206, n21207, n21208, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21223, n21224, n21225,
         n21226, n21227, n21229, n21231, n21232, n21233, n21234, n21235,
         n21236, n21238, n21239, n21241, n21242, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21274, n21277, n21278, n21279, n21280, n21282, n21283, n21284,
         n21285, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21305, n21306, n21307, n21308, n21309, n21310, n21316, n21317,
         n21318, n21319, n21322, n21323, n21324, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21345,
         n21346, n21347, n21349, n21350, n21351, n21352, n21354, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21397, n21398,
         n21399, n21401, n21402, n21403, n21405, n21406, n21407, n21408,
         n21409, n21410, n21412, n21413, n21414, n21415, n21416, n21417,
         n21419, n21420, n21421, n21422, n21423, n21424, n21426, n21428,
         n21429, n21431, n21432, n21433, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21445, n21446, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21467, n21468, n21469, n21472, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21488, n21489, n21491, n21492, n21493, n21494, n21496,
         n21497, n21498, n21499, n21501, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21524, n21527, n21528, n21529, n21531, n21532, n21533, n21534,
         n21535, n21536, n21539, n21540, n21541, n21542, n21543, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21573, n21574, n21575, n21576, n21577, n21579, n21580,
         n21581, n21582, n21583, n21584, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21596, n21597, n21598,
         n21599, n21601, n21602, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21612, n21614, n21616, n21617, n21618, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21644, n21645,
         n21646, n21647, n21648, n21649, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21678, n21679, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21745, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
         n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
         n21766, n21767, n21768, n21770, n21771, n21772, n21773, n21774,
         n21775, n21776, n21777, n21778, n21779, n21780, n21782, n21783,
         n21784, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21808, n21809, n21810,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21820,
         n21821, n21822, n21823, n21825, n21826, n21827, n21828, n21829,
         n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837,
         n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845,
         n21846, n21847, n21848, n21849, n21850, n21852, n21853, n21854,
         n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
         n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870,
         n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
         n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
         n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
         n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
         n21903, n21904, n21905, n21906, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21919, n21920,
         n21921, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21949, n21950, n21951, n21952, n21953, n21954,
         n21956, n21957, n21958, n21959, n21960, n21961, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21971, n21972, n21973,
         n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21982,
         n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990,
         n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
         n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
         n22007, n22008, n22009, n22010, n22012, n22013, n22014, n22015,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22029, n22030, n22032, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22047, n22048, n22050, n22051, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22110, n22111, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22143, n22144, n22145, n22146, n22147, n22148, n22149,
         n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157,
         n22159, n22160, n22161, n22162, n22163, n22165, n22166, n22167,
         n22168, n22170, n22171, n22172, n22173, n22174, n22176, n22177,
         n22178, n22181, n22182, n22183, n22184, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22203, n22204, n22205,
         n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
         n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221,
         n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229,
         n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22252, n22253, n22254, n22255,
         n22256, n22258, n22259, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22270, n22271, n22272, n22274, n22275,
         n22277, n22278, n22279, n22280, n22281, n22282, n22284, n22285,
         n22286, n22287, n22288, n22289, n22291, n22292, n22293, n22294,
         n22295, n22296, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22332, n22333, n22334, n22335, n22337, n22340,
         n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
         n22349, n22350, n22351, n22352, n22353, n22354, n22356, n22358,
         n22359, n22360, n22361, n22362, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22424, n22425, n22426, n22427,
         n22429, n22430, n22431, n22432, n22433, n22435, n22436, n22438,
         n22439, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22456,
         n22457, n22458, n22459, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22473, n22474, n22475, n22476,
         n22478, n22479, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
         n22497, n22498, n22499, n22500, n22501, n22503, n22505, n22506,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22536, n22537, n22538, n22541, n22542,
         n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550,
         n22551, n22552, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22579, n22580, n22581, n22582, n22583, n22584, n22586,
         n22587, n22588, n22590, n22592, n22594, n22595, n22596, n22597,
         n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605,
         n22606, n22607, n22608, n22609, n22610, n22611, n22613, n22614,
         n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622,
         n22623, n22624, n22625, n22627, n22628, n22629, n22630, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22680, n22681, n22682, n22683,
         n22684, n22686, n22687, n22688, n22689, n22690, n22693, n22694,
         n22695, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22740,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22757,
         n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
         n22766, n22767, n22768, n22769, n22771, n22772, n22773, n22774,
         n22775, n22776, n22778, n22780, n22781, n22782, n22783, n22784,
         n22787, n22789, n22790, n22791, n22792, n22793, n22795, n22796,
         n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804,
         n22805, n22806, n22807, n22809, n22810, n22811, n22812, n22813,
         n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22822,
         n22823, n22824, n22825, n22826, n22828, n22829, n22830, n22831,
         n22833, n22834, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22845, n22846, n22849, n22850, n22851, n22852,
         n22853, n22854, n22856, n22857, n22858, n22859, n22860, n22861,
         n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869,
         n22870, n22871, n22872, n22873, n22875, n22876, n22877, n22878,
         n22879, n22880, n22881, n22882, n22884, n22885, n22886, n22887,
         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
         n22897, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22931, n22932, n22934, n22935, n22937, n22939, n22940, n22942,
         n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950,
         n22951, n22952, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22962, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23003, n23004, n23005,
         n23006, n23007, n23009, n23010, n23011, n23012, n23013, n23015,
         n23016, n23017, n23018, n23019, n23020, n23022, n23023, n23024,
         n23025, n23026, n23027, n23028, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
         n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23093, n23094, n23095, n23096, n23098, n23099, n23100, n23101,
         n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23110,
         n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118,
         n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23127,
         n23128, n23129, n23131, n23132, n23133, n23134, n23135, n23136,
         n23137, n23138, n23140, n23141, n23142, n23143, n23145, n23146,
         n23147, n23148, n23149, n23151, n23152, n23154, n23155, n23156,
         n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164,
         n23165, n23166, n23167, n23169, n23171, n23172, n23173, n23174,
         n23175, n23177, n23178, n23180, n23181, n23182, n23183, n23184,
         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
         n23193, n23194, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23206, n23207, n23209, n23210, n23211, n23212, n23213,
         n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221,
         n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229,
         n23232, n23234, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23255, n23256, n23257, n23259, n23262, n23263,
         n23264, n23265, n23266, n23267, n23270, n23271, n23272, n23274,
         n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
         n23283, n23284, n23286, n23289, n23290, n23291, n23292, n23293,
         n23294, n23295, n23296, n23297, n23298, n23299, n23301, n23302,
         n23303, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23320,
         n23321, n23322, n23324, n23325, n23328, n23329, n23330, n23331,
         n23333, n23334, n23335, n23337, n23338, n23340, n23341, n23342,
         n23343, n23344, n23345, n23346, n23347, n23349, n23350, n23351,
         n23352, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
         n23361, n23362, n23363, n23364, n23365, n23367, n23368, n23369,
         n23370, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
         n23379, n23380, n23381, n23382, n23383, n23385, n23386, n23387,
         n23389, n23390, n23391, n23392, n23393, n23394, n23396, n23397,
         n23399, n23400, n23401, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23412, n23413, n23414, n23416, n23418,
         n23419, n23420, n23421, n23422, n23423, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23439, n23440, n23441, n23442, n23444, n23447, n23450, n23452,
         n23453, n23455, n23456, n23458, n23459, n23460, n23461, n23462,
         n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
         n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
         n23480, n23482, n23483, n23484, n23485, n23487, n23488, n23489,
         n23493, n23494, n23496, n23500, n23502, n23504, n23505, n23506,
         n23508, n23509, n23510, n23511, n23512, n23513, n23515, n23516,
         n23517, n23518, n23520, n23521, n23522, n23523, n23525, n23526,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23537, n23538, n23539, n23540, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23552, n23553, n23554,
         n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562,
         n23563, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23574, n23575, n23576, n23577, n23578, n23579, n23580,
         n23581, n23582, n23583, n23584, n23586, n23587, n23588, n23589,
         n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
         n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
         n23606, n23607, n23608, n23609, n23610, n23611, n23613, n23614,
         n23616, n23617, n23619, n23620, n23621, n23622, n23623, n23624,
         n23625, n23627, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23645, n23648,
         n23649, n23652, n23653, n23654, n23655, n23656, n23658, n23659,
         n23660, n23661, n23662, n23663, n23665, n23666, n23667, n23668,
         n23669, n23670, n23671, n23672, n23674, n23675, n23676, n23677,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23702, n23704, n23705,
         n23707, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23719, n23720, n23722, n23723, n23724, n23725,
         n23727, n23728, n23729, n23730, n23732, n23733, n23734, n23736,
         n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,
         n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23792, n23793, n23794,
         n23795, n23796, n23797, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23812, n23813,
         n23814, n23816, n23817, n23818, n23819, n23820, n23821, n23822,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23838, n23839, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23855, n23857, n23858, n23859,
         n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868,
         n23869, n23870, n23871, n23873, n23874, n23876, n23878, n23879,
         n23880, n23882, n23883, n23884, n23885, n23886, n23887, n23888,
         n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,
         n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904,
         n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,
         n23913, n23914, n23915, n23917, n23918, n23919, n23920, n23921,
         n23922, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
         n23931, n23933, n23934, n23936, n23937, n23938, n23939, n23940,
         n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948,
         n23949, n23950, n23952, n23953, n23954, n23955, n23957, n23958,
         n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966,
         n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974,
         n23975, n23976, n23977, n23979, n23980, n23981, n23982, n23983,
         n23984, n23985, n23987, n23988, n23989, n23990, n23991, n23992,
         n23993, n23994, n23995, n23996, n23997, n24000, n24001, n24002,
         n24005, n24006, n24007, n24009, n24011, n24012, n24013, n24014,
         n24015, n24016, n24017, n24018, n24019, n24020, n24022, n24023,
         n24024, n24025, n24026, n24028, n24029, n24030, n24031, n24032,
         n24033, n24034, n24036, n24037, n24038, n24039, n24040, n24042,
         n24043, n24045, n24047, n24048, n24049, n24050, n24051, n24052,
         n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060,
         n24061, n24062, n24063, n24064, n24065, n24067, n24068, n24069,
         n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
         n24078, n24079, n24081, n24082, n24083, n24084, n24085, n24086,
         n24087, n24088, n24089, n24090, n24091, n24094, n24095, n24096,
         n24098, n24100, n24101, n24102, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24116,
         n24117, n24118, n24119, n24120, n24121, n24123, n24125, n24126,
         n24127, n24128, n24129, n24131, n24132, n24133, n24134, n24135,
         n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143,
         n24145, n24146, n24147, n24148, n24149, n24150, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24161, n24162,
         n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24180,
         n24181, n24182, n24184, n24185, n24187, n24191, n24192, n24193,
         n24194, n24195, n24196, n24198, n24199, n24202, n24203, n24205,
         n24206, n24207, n24208, n24209, n24210, n24214, n24216, n24217,
         n24218, n24219, n24221, n24222, n24223, n24224, n24225, n24226,
         n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234,
         n24235, n24238, n24240, n24241, n24242, n24243, n24244, n24245,
         n24246, n24247, n24250, n24251, n24253, n24254, n24257, n24258,
         n24261, n24263, n24265, n24266, n24267, n24268, n24269, n24270,
         n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
         n24279, n24280, n24282, n24283, n24284, n24285, n24287, n24290,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24300,
         n24301, n24302, n24303, n24304, n24305, n24307, n24308, n24309,
         n24310, n24311, n24312, n24313, n24314, n24316, n24317, n24318,
         n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24331, n24332, n24333, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24345, n24346, n24347, n24348,
         n24349, n24350, n24351, n24353, n24355, n24357, n24359, n24360,
         n24363, n24364, n24365, n24366, n24369, n24370, n24371, n24372,
         n24373, n24374, n24377, n24378, n24380, n24381, n24382, n24383,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24406, n24407, n24408, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24419, n24420,
         n24421, n24424, n24425, n24426, n24427, n24429, n24430, n24431,
         n24432, n24433, n24434, n24436, n24437, n24438, n24439, n24440,
         n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
         n24449, n24451, n24452, n24453, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24463, n24464, n24465, n24466, n24467,
         n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476,
         n24477, n24478, n24479, n24481, n24483, n24484, n24485, n24490,
         n24491, n24492, n24493, n24494, n24495, n24496, n24498, n24499,
         n24500, n24502, n24504, n24506, n24507, n24509, n24510, n24511,
         n24514, n24515, n24516, n24517, n24518, n24524, n24525, n24526,
         n24527, n24528, n24529, n24530, n24531, n24532, n24534, n24535,
         n24536, n24538, n24539, n24540, n24541, n24542, n24543, n24544,
         n24545, n24546, n24547, n24550, n24551, n24552, n24553, n24554,
         n24556, n24557, n24558, n24560, n24561, n24563, n24565, n24566,
         n24568, n24569, n24571, n24572, n24573, n24574, n24575, n24576,
         n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,
         n24585, n24586, n24588, n24589, n24590, n24591, n24592, n24593,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24605, n24606, n24607, n24608, n24609, n24610, n24612,
         n24613, n24614, n24615, n24616, n24618, n24619, n24620, n24621,
         n24622, n24623, n24624, n24625, n24626, n24627, n24629, n24630,
         n24631, n24632, n24633, n24634, n24635, n24637, n24638, n24639,
         n24641, n24643, n24644, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24655, n24656, n24657, n24658, n24659, n24660,
         n24661, n24662, n24663, n24664, n24665, n24666, n24668, n24669,
         n24670, n24671, n24672, n24673, n24674, n24676, n24678, n24679,
         n24680, n24681, n24683, n24685, n24686, n24687, n24689, n24690,
         n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
         n24699, n24700, n24701, n24702, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24715, n24716,
         n24717, n24719, n24720, n24721, n24723, n24724, n24725, n24726,
         n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734,
         n24735, n24736, n24737, n24738, n24740, n24741, n24743, n24744,
         n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752,
         n24753, n24754, n24755, n24757, n24759, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24774, n24775, n24776, n24777, n24778, n24779, n24780,
         n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789,
         n24792, n24793, n24794, n24795, n24798, n24799, n24800, n24801,
         n24802, n24804, n24805, n24806, n24810, n24811, n24812, n24813,
         n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821,
         n24822, n24823, n24824, n24826, n24827, n24828, n24829, n24832,
         n24833, n24834, n24836, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24847, n24849, n24850, n24852, n24853,
         n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861,
         n24862, n24863, n24864, n24866, n24868, n24869, n24871, n24872,
         n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24882,
         n24883, n24884, n24885, n24886, n24887, n24891, n24892, n24894,
         n24895, n24896, n24897, n24898, n24899, n24900, n24902, n24903,
         n24904, n24905, n24906, n24907, n24909, n24910, n24912, n24913,
         n24914, n24915, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24935, n24936, n24937, n24938, n24940,
         n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948,
         n24949, n24950, n24952, n24953, n24954, n24955, n24957, n24958,
         n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966,
         n24967, n24968, n24970, n24971, n24972, n24973, n24974, n24975,
         n24976, n24977, n24978, n24981, n24982, n24984, n24985, n24987,
         n24988, n24989, n24990, n24991, n24992, n24994, n24997, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25014, n25015, n25016,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25051,
         n25052, n25053, n25054, n25055, n25056, n25059, n25060, n25061,
         n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25070,
         n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
         n25079, n25080, n25081, n25083, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25108, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25132, n25133,
         n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
         n25142, n25143, n25144, n25145, n25146, n25148, n25149, n25150,
         n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158,
         n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166,
         n25167, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25200, n25201,
         n25202, n25203, n25204, n25206, n25207, n25208, n25210, n25211,
         n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220,
         n25221, n25222, n25224, n25225, n25226, n25229, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25283,
         n25284, n25285, n25286, n25288, n25289, n25290, n25291, n25292,
         n25293, n25295, n25296, n25298, n25299, n25300, n25301, n25302,
         n25303, n25304, n25305, n25307, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25322, n25323, n25324, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25339,
         n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
         n25349, n25351, n25352, n25353, n25354, n25355, n25358, n25359,
         n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367,
         n25368, n25369, n25370, n25371, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25392, n25393,
         n25394, n25395, n25396, n25397, n25399, n25400, n25401, n25402,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25412,
         n25416, n25418, n25420, n25421, n25422, n25424, n25425, n25427,
         n25428, n25429, n25430, n25431, n25433, n25434, n25435, n25436,
         n25437, n25438, n25439, n25440, n25441, n25443, n25444, n25445,
         n25447, n25448, n25449, n25450, n25451, n25452, n25454, n25455,
         n25456, n25457, n25458, n25459, n25460, n25462, n25464, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25486, n25487, n25488, n25489, n25490, n25491, n25495,
         n25497, n25498, n25499, n25501, n25502, n25503, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25519, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25562, n25563,
         n25564, n25566, n25567, n25568, n25569, n25571, n25572, n25573,
         n25574, n25575, n25576, n25577, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25592, n25593, n25594, n25595, n25596,
         n25597, n25598, n25600, n25601, n25602, n25603, n25604, n25605,
         n25606, n25608, n25609, n25611, n25612, n25613, n25614, n25615,
         n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623,
         n25625, n25627, n25628, n25630, n25631, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25641, n25642, n25643, n25644,
         n25645, n25647, n25649, n25650, n25651, n25655, n25657, n25658,
         n25659, n25660, n25661, n25662, n25665, n25666, n25667, n25669,
         n25670, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25702, n25705, n25706, n25707, n25708, n25712,
         n25713, n25714, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25751, n25753, n25754, n25755, n25756,
         n25758, n25759, n25760, n25761, n25762, n25764, n25766, n25767,
         n25768, n25769, n25770, n25771, n25772, n25774, n25775, n25776,
         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
         n25785, n25787, n25788, n25790, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25803, n25804,
         n25805, n25807, n25808, n25809, n25810, n25812, n25813, n25814,
         n25815, n25817, n25818, n25819, n25820, n25821, n25822, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25833, n25834,
         n25835, n25836, n25837, n25838, n25840, n25841, n25842, n25844,
         n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852,
         n25853, n25854, n25855, n25856, n25857, n25858, n25860, n25861,
         n25862, n25865, n25866, n25867, n25868, n25869, n25870, n25871,
         n25872, n25874, n25875, n25876, n25877, n25878, n25879, n25882,
         n25883, n25886, n25887, n25888, n25889, n25891, n25892, n25894,
         n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903,
         n25904, n25905, n25907, n25910, n25911, n25912, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25930, n25931, n25933,
         n25934, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
         n25943, n25945, n25946, n25947, n25949, n25950, n25951, n25954,
         n25955, n25956, n25957, n25958, n25959, n25961, n25962, n25964,
         n25965, n25966, n25967, n25970, n25971, n25972, n25975, n25977,
         n25978, n25979, n25981, n25982, n25983, n25984, n25985, n25986,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25998, n25999, n26000, n26001, n26003, n26004, n26005,
         n26006, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
         n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022,
         n26023, n26024, n26026, n26027, n26028, n26029, n26030, n26031,
         n26032, n26034, n26035, n26036, n26037, n26038, n26039, n26041,
         n26042, n26045, n26048, n26050, n26051, n26052, n26053, n26054,
         n26055, n26056, n26058, n26059, n26060, n26061, n26063, n26065,
         n26066, n26067, n26068, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26081, n26083, n26084,
         n26085, n26086, n26088, n26089, n26090, n26092, n26093, n26094,
         n26095, n26096, n26097, n26098, n26099, n26101, n26103, n26104,
         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
         n26121, n26122, n26123, n26124, n26125, n26126, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26137, n26138,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26160, n26161, n26162, n26163, n26165,
         n26166, n26167, n26168, n26169, n26171, n26172, n26173, n26176,
         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
         n26185, n26186, n26187, n26188, n26190, n26191, n26192, n26194,
         n26195, n26196, n26197, n26198, n26200, n26201, n26204, n26205,
         n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213,
         n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
         n26222, n26223, n26224, n26225, n26227, n26228, n26229, n26230,
         n26231, n26232, n26233, n26234, n26236, n26237, n26238, n26239,
         n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247,
         n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26268, n26269, n26270, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26299, n26301,
         n26302, n26303, n26304, n26305, n26307, n26308, n26309, n26310,
         n26311, n26312, n26313, n26314, n26316, n26317, n26318, n26319,
         n26320, n26321, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26346,
         n26347, n26348, n26349, n26350, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26363, n26364,
         n26365, n26366, n26368, n26369, n26370, n26371, n26372, n26373,
         n26374, n26375, n26376, n26377, n26379, n26380, n26381, n26382,
         n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390,
         n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
         n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26407,
         n26408, n26409, n26410, n26411, n26412, n26413, n26415, n26417,
         n26418, n26419, n26420, n26421, n26422, n26424, n26425, n26426,
         n26427, n26428, n26429, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460,
         n26461, n26462, n26463, n26464, n26465, n26466, n26468, n26470,
         n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478,
         n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26500, n26502, n26503, n26504,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532,
         n26536, n26537, n26538, n26539, n26541, n26542, n26544, n26545,
         n26547, n26548, n26550, n26551, n26553, n26554, n26555, n26556,
         n26557, n26558, n26559, n26560, n26561, n26562, n26564, n26565,
         n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573,
         n26574, n26575, n26577, n26578, n26579, n26580, n26581, n26582,
         n26584, n26585, n26587, n26588, n26590, n26591, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26605, n26606, n26607, n26608, n26609, n26610, n26612, n26614,
         n26618, n26619, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26630, n26632, n26634, n26635, n26636, n26637,
         n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645,
         n26647, n26648, n26650, n26651, n26652, n26653, n26655, n26657,
         n26659, n26660, n26661, n26662, n26663, n26665, n26666, n26667,
         n26668, n26670, n26671, n26672, n26674, n26675, n26678, n26679,
         n26682, n26684, n26686, n26687, n26688, n26689, n26691, n26692,
         n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
         n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709,
         n26710, n26713, n26717, n26718, n26719, n26720, n26721, n26722,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26737, n26738, n26740, n26741, n26743,
         n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
         n26752, n26754, n26755, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26783, n26784, n26785, n26786, n26787, n26788, n26789,
         n26790, n26791, n26793, n26794, n26795, n26796, n26797, n26798,
         n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
         n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26815,
         n26816, n26817, n26818, n26819, n26822, n26823, n26824, n26825,
         n26826, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26856, n26857, n26858, n26859, n26860,
         n26861, n26862, n26863, n26864, n26865, n26866, n26868, n26869,
         n26870, n26871, n26872, n26876, n26877, n26878, n26879, n26882,
         n26885, n26887, n26888, n26889, n26890, n26892, n26893, n26895,
         n26897, n26898, n26899, n26901, n26902, n26903, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26918, n26919, n26920, n26921, n26922, n26923,
         n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
         n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
         n26942, n26943, n26944, n26945, n26946, n26948, n26950, n26951,
         n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
         n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
         n26970, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26998, n26999, n27000, n27001, n27004, n27006,
         n27007, n27009, n27010, n27011, n27013, n27014, n27015, n27017,
         n27018, n27020, n27021, n27023, n27024, n27026, n27027, n27028,
         n27029, n27030, n27031, n27032, n27033, n27035, n27036, n27037,
         n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045,
         n27046, n27047, n27048, n27049, n27051, n27052, n27053, n27054,
         n27055, n27056, n27057, n27059, n27060, n27061, n27062, n27063,
         n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
         n27072, n27073, n27076, n27078, n27079, n27080, n27081, n27083,
         n27084, n27085, n27087, n27088, n27089, n27090, n27092, n27093,
         n27094, n27095, n27096, n27097, n27098, n27099, n27102, n27103,
         n27106, n27107, n27108, n27109, n27110, n27111, n27113, n27114,
         n27115, n27116, n27118, n27119, n27121, n27122, n27123, n27124,
         n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27133,
         n27135, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
         n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151,
         n27152, n27153, n27154, n27155, n27158, n27159, n27161, n27163,
         n27164, n27165, n27166, n27167, n27169, n27170, n27171, n27172,
         n27174, n27175, n27176, n27178, n27180, n27181, n27182, n27184,
         n27185, n27187, n27189, n27192, n27193, n27194, n27196, n27197,
         n27198, n27199, n27200, n27201, n27203, n27204, n27205, n27206,
         n27207, n27211, n27213, n27214, n27215, n27218, n27220, n27221,
         n27224, n27225, n27226, n27228, n27229, n27230, n27231, n27232,
         n27233, n27234, n27235, n27236, n27237, n27238, n27240, n27242,
         n27244, n27245, n27247, n27248, n27249, n27250, n27251, n27252,
         n27253, n27255, n27256, n27257, n27258, n27259, n27263, n27265,
         n27266, n27267, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27278, n27279, n27282, n27283, n27284, n27285,
         n27286, n27287, n27288, n27289, n27291, n27292, n27295, n27296,
         n27297, n27298, n27299, n27300, n27302, n27304, n27305, n27306,
         n27307, n27310, n27311, n27312, n27314, n27315, n27316, n27317,
         n27318, n27319, n27320, n27321, n27324, n27325, n27326, n27328,
         n27329, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27353, n27354, n27356, n27357,
         n27358, n27360, n27361, n27362, n27363, n27364, n27365, n27366,
         n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375,
         n27376, n27377, n27378, n27379, n27381, n27382, n27383, n27384,
         n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
         n27393, n27395, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27415, n27416, n27417, n27419, n27420,
         n27421, n27422, n27424, n27426, n27428, n27429, n27430, n27431,
         n27433, n27434, n27435, n27436, n27438, n27440, n27441, n27444,
         n27445, n27446, n27447, n27448, n27449, n27451, n27452, n27453,
         n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462,
         n27463, n27464, n27465, n27466, n27467, n27469, n27470, n27471,
         n27472, n27473, n27474, n27475, n27477, n27478, n27479, n27480,
         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,
         n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
         n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,
         n27505, n27506, n27507, n27508, n27509, n27511, n27513, n27514,
         n27515, n27516, n27517, n27518, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27546, n27547, n27548, n27549,
         n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557,
         n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565,
         n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573,
         n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581,
         n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590,
         n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598,
         n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607,
         n27608, n27609, n27611, n27612, n27613, n27614, n27615, n27617,
         n27618, n27619, n27620, n27621, n27622, n27624, n27626, n27627,
         n27628, n27630, n27631, n27632, n27633, n27634, n27635, n27636,
         n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27645,
         n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
         n27654, n27655, n27657, n27658, n27659, n27661, n27662, n27663,
         n27664, n27665, n27666, n27667, n27668, n27669, n27671, n27672,
         n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680,
         n27681, n27683, n27685, n27686, n27687, n27688, n27689, n27690,
         n27692, n27695, n27696, n27697, n27698, n27700, n27701, n27703,
         n27704, n27705, n27706, n27707, n27709, n27710, n27711, n27712,
         n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720,
         n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728,
         n27729, n27730, n27731, n27732, n27733, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27745, n27746,
         n27748, n27749, n27750, n27751, n27753, n27754, n27755, n27756,
         n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
         n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
         n27773, n27774, n27776, n27777, n27778, n27779, n27781, n27782,
         n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
         n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799,
         n27800, n27802, n27803, n27804, n27805, n27806, n27807, n27808,
         n27809, n27810, n27812, n27813, n27815, n27816, n27817, n27818,
         n27819, n27820, n27822, n27823, n27825, n27826, n27827, n27828,
         n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
         n27837, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
         n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854,
         n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862,
         n27863, n27864, n27865, n27866, n27867, n27868, n27870, n27871,
         n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879,
         n27880, n27881, n27882, n27883, n27884, n27885, n27887, n27888,
         n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896,
         n27897, n27898, n27900, n27901, n27902, n27903, n27904, n27906,
         n27907, n27908, n27909, n27910, n27911, n27913, n27914, n27915,
         n27917, n27918, n27919, n27920, n27921, n27925, n27926, n27927,
         n27928, n27929, n27930, n27932, n27934, n27935, n27936, n27938,
         n27940, n27941, n27942, n27943, n27944, n27946, n27948, n27951,
         n27955, n27956, n27957, n27958, n27959, n27962, n27963, n27964,
         n27966, n27967, n27969, n27970, n27972, n27973, n27974, n27976,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n28001, n28002, n28004,
         n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
         n28014, n28015, n28017, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28038, n28039, n28040, n28041, n28042,
         n28043, n28045, n28047, n28048, n28049, n28050, n28051, n28052,
         n28053, n28054, n28056, n28057, n28058, n28059, n28060, n28061,
         n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069,
         n28073, n28074, n28075, n28079, n28080, n28081, n28082, n28083,
         n28085, n28086, n28087, n28089, n28091, n28093, n28095, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28111, n28112, n28113, n28114, n28115,
         n28117, n28118, n28119, n28122, n28123, n28124, n28125, n28126,
         n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134,
         n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144,
         n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152,
         n28153, n28154, n28155, n28156, n28157, n28159, n28161, n28162,
         n28163, n28164, n28165, n28167, n28168, n28170, n28171, n28172,
         n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
         n28181, n28182, n28184, n28185, n28186, n28187, n28188, n28189,
         n28190, n28191, n28192, n28193, n28194, n28195, n28197, n28199,
         n28200, n28202, n28203, n28204, n28205, n28206, n28207, n28209,
         n28210, n28212, n28213, n28214, n28215, n28216, n28217, n28219,
         n28220, n28221, n28222, n28223, n28224, n28226, n28227, n28228,
         n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236,
         n28237, n28238, n28240, n28242, n28243, n28244, n28245, n28246,
         n28247, n28248, n28249, n28250, n28251, n28255, n28256, n28257,
         n28258, n28259, n28260, n28262, n28263, n28264, n28265, n28266,
         n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
         n28276, n28278, n28279, n28281, n28282, n28283, n28284, n28285,
         n28286, n28287, n28288, n28289, n28290, n28291, n28293, n28297,
         n28298, n28299, n28301, n28302, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28322, n28323, n28324,
         n28325, n28326, n28327, n28328, n28330, n28331, n28332, n28333,
         n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342,
         n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350,
         n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358,
         n28359, n28360, n28361, n28362, n28364, n28365, n28366, n28368,
         n28369, n28370, n28372, n28373, n28375, n28376, n28377, n28378,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28389, n28390, n28391, n28392, n28394, n28395, n28396, n28398,
         n28399, n28400, n28401, n28402, n28403, n28406, n28408, n28409,
         n28410, n28411, n28412, n28414, n28415, n28416, n28417, n28418,
         n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
         n28427, n28428, n28429, n28430, n28431, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28442, n28443, n28444,
         n28445, n28448, n28450, n28452, n28453, n28454, n28455, n28456,
         n28457, n28458, n28460, n28463, n28464, n28465, n28466, n28467,
         n28468, n28470, n28471, n28473, n28475, n28477, n28478, n28479,
         n28480, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28507, n28508, n28509, n28510, n28513, n28514, n28515, n28516,
         n28518, n28520, n28521, n28522, n28523, n28524, n28525, n28528,
         n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28553, n28554,
         n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
         n28563, n28564, n28565, n28568, n28569, n28570, n28571, n28573,
         n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28583,
         n28584, n28585, n28586, n28587, n28589, n28590, n28591, n28592,
         n28594, n28595, n28596, n28598, n28601, n28603, n28604, n28605,
         n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28614,
         n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622,
         n28623, n28625, n28626, n28627, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28643, n28644, n28647, n28648, n28649, n28650, n28651, n28652,
         n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
         n28661, n28662, n28664, n28665, n28666, n28669, n28670, n28671,
         n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680,
         n28681, n28682, n28683, n28685, n28686, n28689, n28690, n28691,
         n28692, n28693, n28695, n28696, n28697, n28698, n28699, n28700,
         n28704, n28705, n28707, n28708, n28709, n28710, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28732, n28733, n28735, n28736, n28738, n28739, n28740,
         n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749,
         n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757,
         n28758, n28759, n28761, n28762, n28763, n28764, n28765, n28767,
         n28768, n28769, n28770, n28771, n28772, n28773, n28775, n28776,
         n28777, n28778, n28779, n28780, n28782, n28783, n28785, n28786,
         n28787, n28788, n28789, n28790, n28791, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28811, n28812, n28813,
         n28814, n28815, n28817, n28819, n28820, n28821, n28822, n28823,
         n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28857, n28858, n28859, n28860,
         n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869,
         n28870, n28871, n28873, n28874, n28876, n28878, n28880, n28882,
         n28883, n28885, n28886, n28887, n28888, n28889, n28891, n28892,
         n28893, n28894, n28895, n28896, n28898, n28899, n28900, n28901,
         n28902, n28903, n28904, n28905, n28906, n28907, n28909, n28910,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28923, n28924, n28925, n28927, n28928, n28930, n28931,
         n28933, n28934, n28935, n28940, n28943, n28944, n28945, n28946,
         n28947, n28948, n28949, n28950, n28951, n28953, n28954, n28955,
         n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964,
         n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973,
         n28975, n28976, n28977, n28978, n28979, n28980, n28982, n28983,
         n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991,
         n28992, n28993, n28994, n28996, n28997, n28998, n28999, n29000,
         n29001, n29002, n29003, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29014, n29015, n29016, n29017, n29019,
         n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028,
         n29029, n29030, n29031, n29033, n29034, n29035, n29036, n29037,
         n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045,
         n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29054,
         n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29063,
         n29064, n29065, n29066, n29067, n29068, n29070, n29071, n29072,
         n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
         n29081, n29082, n29083, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29102, n29103, n29104, n29105, n29107,
         n29108, n29109, n29110, n29111, n29113, n29114, n29115, n29119,
         n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127,
         n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135,
         n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144,
         n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
         n29153, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29171, n29173, n29174, n29175, n29176, n29180, n29181, n29182,
         n29183, n29184, n29185, n29187, n29188, n29189, n29190, n29191,
         n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199,
         n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207,
         n29208, n29209, n29210, n29211, n29212, n29214, n29217, n29218,
         n29219, n29220, n29221, n29222, n29223, n29224, n29226, n29228,
         n29229, n29230, n29231, n29232, n29233, n29234, n29236, n29237,
         n29238, n29239, n29241, n29242, n29243, n29244, n29245, n29246,
         n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254,
         n29255, n29257, n29258, n29260, n29262, n29263, n29265, n29266,
         n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274,
         n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
         n29284, n29285, n29286, n29287, n29289, n29290, n29291, n29292,
         n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300,
         n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29309,
         n29310, n29312, n29313, n29314, n29315, n29316, n29317, n29318,
         n29319, n29320, n29321, n29323, n29324, n29325, n29326, n29327,
         n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335,
         n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29344,
         n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29365, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29375, n29377, n29378, n29379, n29380, n29381,
         n29382, n29383, n29384, n29385, n29389, n29390, n29391, n29392,
         n29393, n29394, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
         n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
         n29427, n29430, n29431, n29432, n29433, n29434, n29435, n29436,
         n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444,
         n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452,
         n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29461,
         n29462, n29463, n29464, n29466, n29467, n29468, n29469, n29470,
         n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479,
         n29480, n29481, n29482, n29483, n29485, n29486, n29488, n29489,
         n29490, n29491, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516,
         n29517, n29519, n29520, n29521, n29522, n29523, n29524, n29525,
         n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533,
         n29534, n29535, n29536, n29538, n29539, n29540, n29541, n29542,
         n29543, n29546, n29547, n29548, n29549, n29550, n29551, n29552,
         n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560,
         n29562, n29563, n29565, n29566, n29567, n29568, n29569, n29570,
         n29571, n29572, n29573, n29574, n29575, n29577, n29578, n29579,
         n29580, n29581, n29583, n29586, n29587, n29591, n29592, n29593,
         n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
         n29604, n29605, n29607, n29608, n29610, n29611, n29612, n29613,
         n29614, n29615, n29616, n29617, n29618, n29619, n29621, n29622,
         n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630,
         n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
         n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
         n29648, n29649, n29652, n29654, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29682, n29683, n29684,
         n29685, n29686, n29687, n29688, n29689, n29690, n29692, n29693,
         n29694, n29696, n29697, n29698, n29699, n29700, n29701, n29702,
         n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
         n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718,
         n29719, n29720, n29721, n29722, n29723, n29725, n29726, n29727,
         n29728, n29729, n29730, n29731, n29732, n29733, n29735, n29736,
         n29737, n29739, n29740, n29741, n29747, n29749, n29750, n29751,
         n29752, n29753, n29754, n29755, n29756, n29758, n29759, n29760,
         n29761, n29762, n29763, n29764, n29767, n29768, n29769, n29770,
         n29771, n29774, n29775, n29776, n29777, n29779, n29780, n29781,
         n29782, n29783, n29784, n29785, n29787, n29788, n29789, n29790,
         n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
         n29799, n29800, n29801, n29802, n29803, n29805, n29806, n29807,
         n29808, n29809, n29810, n29811, n29812, n29813, n29815, n29816,
         n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824,
         n29825, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29849, n29851,
         n29852, n29854, n29855, n29856, n29857, n29858, n29859, n29860,
         n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29869,
         n29870, n29871, n29873, n29874, n29875, n29876, n29877, n29879,
         n29880, n29881, n29883, n29884, n29885, n29887, n29888, n29889,
         n29890, n29892, n29895, n29896, n29897, n29898, n29899, n29900,
         n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908,
         n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916,
         n29918, n29919, n29920, n29922, n29923, n29924, n29925, n29927,
         n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
         n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943,
         n29946, n29947, n29948, n29949, n29951, n29952, n29953, n29954,
         n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
         n29963, n29964, n29965, n29966, n29967, n29968, n29970, n29971,
         n29973, n29974, n29975, n29977, n29978, n29979, n29980, n29981,
         n29982, n29983, n29985, n29986, n29987, n29988, n29989, n29990,
         n29991, n29992, n29993, n29994, n29996, n29997, n29998, n30000,
         n30001, n30002, n30003, n30004, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30030, n30031, n30032, n30033, n30034,
         n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042,
         n30043, n30045, n30046, n30047, n30048, n30049, n30051, n30052,
         n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060,
         n30062, n30063, n30065, n30066, n30067, n30068, n30069, n30070,
         n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
         n30079, n30080, n30081, n30083, n30084, n30085, n30086, n30087,
         n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096,
         n30097, n30098, n30099, n30100, n30101, n30102, n30104, n30105,
         n30106, n30107, n30109, n30110, n30111, n30112, n30113, n30114,
         n30115, n30116, n30117, n30118, n30119, n30120, n30122, n30126,
         n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134,
         n30135, n30136, n30138, n30139, n30140, n30141, n30143, n30144,
         n30145, n30146, n30147, n30150, n30152, n30153, n30154, n30155,
         n30156, n30158, n30159, n30160, n30161, n30162, n30163, n30165,
         n30166, n30168, n30169, n30170, n30171, n30172, n30173, n30174,
         n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
         n30183, n30184, n30185, n30186, n30187, n30190, n30191, n30192,
         n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30201,
         n30203, n30204, n30205, n30206, n30207, n30210, n30211, n30212,
         n30213, n30214, n30215, n30216, n30217, n30220, n30221, n30222,
         n30223, n30225, n30228, n30229, n30230, n30231, n30232, n30233,
         n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244,
         n30245, n30246, n30247, n30248, n30249, n30250, n30252, n30253,
         n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
         n30263, n30272, n30274, n30275, n30276, n30279, n30280, n30282,
         n30283, n30284, n30285, n30288, n30290, n30292, n30293, n30295,
         n30299, n30302, n30304, n30306, n30311, n30315, n30317, n30318,
         n30320, n30321, n30322, n30323, n30324, n30326, n30329, n30330,
         n30333, n30334, n30335, n30336, n30338, n30339, n30340, n30342,
         n30345, n30347, n30348, n30350, n30352, n30353, n30354, n30355,
         n30356, n30357, n30358, n30360, n30363, n30364, n30365, n30366,
         n30368, n30369, n30370, n30371, n30372, n30373, n30377, n30378,
         n30379, n30380, n30381, n30384, n30385, n30386, n30388, n30389,
         n30391, n30392, n30393, n30394, n30396, n30397, n30399, n30400,
         n30401, n30402, n30403, n30404, n30405, n30406, n30408, n30409,
         n30410, n30412, n30413, n30414, n30416, n30417, n30419, n30420,
         n30421, n30422, n30423, n30424, n30425, n30427, n30429, n30431,
         n30432, n30433, n30434, n30435, n30436, n30440, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30450, n30451, n30452,
         n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460,
         n30461, n30463, n30464, n30465, n30468, n30469, n30470, n30471,
         n30473, n30475, n30478, n30479, n30480, n30481, n30482, n30483,
         n30484, n30485, n30486, n30487, n30488, n30489, n30494, n30496,
         n30499, n30500, n30502, n30503, n30504, n30506, n30507, n30509,
         n30512, n30519, n30520, n30524, n30526, n30528, n30529, n30530,
         n30534, n30539, n30541, n30542, n30544, n30546, n30547, n30548,
         n30550, n30551, n30554, n30555, n30556, n30558, n30560, n30561,
         n30562, n30565, n30568, n30571, n30572, n30574, n30577, n30578,
         n30580, n30581, n30582, n30584, n30585, n30587, n30588, n30594,
         n30595, n30596, n30597, n30598, n30599, n30602, n30603, n30607,
         n30608, n30609, n30610, n30611, n30612, n30613, n30615, n30616,
         n30617, n30619, n30621, n30623, n30625, n30626, n30629, n30631,
         n30632, n30633, n30635, n30636, n30642, n30643, n30644, n30645,
         n30646, n30647, n30648, n30649, n30651, n30652, n30653, n30655,
         n30656, n30657, n30659, n30661, n30663, n30664, n30665, n30667,
         n30668, n30671, n30674, n30675, n30676, n30677, n30678, n30680,
         n30682, n30684, n30687, n30688, n30689, n30694, n30695, n30696,
         n30698, n30699, n30700, n30701, n30702, n30704, n30705, n30706,
         n30709, n30711, n30712, n30714, n30715, n30716, n30720, n30722,
         n30724, n30725, n30726, n30727, n30728, n30730, n30731, n30732,
         n30733, n30734, n30736, n30738, n30740, n30741, n30745, n30746,
         n30747, n30748, n30756, n30757, n30758, n30761, n30764, n30766,
         n30768, n30771, n30773, n30775, n30776, n30778, n30780, n30781,
         n30785, n30786, n30788, n30789, n30793, n30794, n30795, n30796,
         n30798, n30799, n30800, n30803, n30805, n30806, n30808, n30811,
         n30813, n30815, n30817, n30818, n30819, n30822, n30824, n30825,
         n30826, n30828, n30831, n30833, n30835, n30837, n30838, n30839,
         n30840, n30842, n30843, n30844, n30845, n30846, n30847, n30849,
         n30850, n30851, n30853, n30854, n30856, n30857, n30858, n30859,
         n30862, n30863, n30865, n30871, n30872, n30874, n30877, n30878,
         n30881, n30883, n30886, n30888, n30890, n30891, n30893, n30894,
         n30895, n30897, n30898, n30900, n30905, n30907, n30908, n30910,
         n30913, n30914, n30915, n30917, n30925, n30927, n30928, n30929,
         n30930, n30931, n30933, n30934, n30936, n30937, n30938, n30939,
         n30941, n30942, n30944, n30945, n30946, n30947, n30948, n30949,
         n30950, n30951, n30952, n30953, n30955, n30956, n30957, n30958,
         n30959, n30960, n30962, n30963, n30964, n30965, n30966, n30967,
         n30971, n30972, n30973, n30974, n30976, n30980, n30981, n30982,
         n30983, n30986, n30988, n30989, n30990, n30991, n30993, n30994,
         n30995, n30996, n31000, n31001, n31002, n31003, n31004, n31005,
         n31006, n31010, n31012, n31014, n31015, n31016, n31017, n31018,
         n31019, n31020, n31022, n31023, n31025, n31027, n31028, n31030,
         n31031, n31034, n31035, n31036, n31037, n31038, n31042, n31043,
         n31044, n31045, n31046, n31047, n31048, n31049, n31052, n31055,
         n31059, n31060, n31061, n31062, n31065, n31070, n31073, n31074,
         n31075, n31077, n31078, n31079, n31080, n31081, n31082, n31086,
         n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
         n31095, n31098, n31102, n31103, n31107, n31108, n31110, n31112,
         n31114, n31115, n31116, n31118, n31119, n31120, n31121, n31122,
         n31123, n31124, n31125, n31127, n31129, n31130, n31131, n31132,
         n31133, n31137, n31138, n31139, n31143, n31144, n31146, n31147,
         n31149, n31150, n31151, n31152, n31154, n31156, n31157, n31158,
         n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31168,
         n31170, n31173, n31175, n31177, n31178, n31179, n31180, n31181,
         n31183, n31184, n31185, n31191, n31192, n31194, n31196, n31197,
         n31198, n31199, n31200, n31202, n31204, n31205, n31206, n31207,
         n31211, n31212, n31213, n31214, n31215, n31218, n31220, n31222,
         n31223, n31225, n31226, n31227, n31230, n31231, n31233, n31234,
         n31235, n31236, n31237, n31238, n31240, n31242, n31245, n31247,
         n31248, n31249, n31250, n31252, n31253, n31254, n31257, n31258,
         n31261, n31263, n31264, n31267, n31268, n31269, n31270, n31271,
         n31272, n31273, n31274, n31275, n31277, n31278, n31279, n31280,
         n31281, n31283, n31284, n31287, n31289, n31290, n31292, n31293,
         n31294, n31295, n31296, n31298, n31299, n31300, n31302, n31304,
         n31305, n31307, n31310, n31311, n31312, n31313, n31314, n31318,
         n31319, n31320, n31321, n31322, n31325, n31326, n31327, n31328,
         n31329, n31331, n31332, n31334, n31335, n31339, n31340, n31341,
         n31343, n31345, n31346, n31347, n31348, n31349, n31350, n31351,
         n31352, n31353, n31355, n31356, n31357, n31358, n31359, n31360,
         n31361, n31362, n31364, n31365, n31366, n31367, n31369, n31370,
         n31371, n31374, n31375, n31376, n31377, n31378, n31379, n31381,
         n31383, n31385, n31386, n31388, n31389, n31390, n31393, n31396,
         n31398, n31399, n31400, n31401, n31403, n31404, n31406, n31407,
         n31410, n31412, n31414, n31416, n31418, n31421, n31424, n31425,
         n31426, n31427, n31428, n31430, n31432, n31433, n31437, n31438,
         n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31452,
         n31453, n31455, n31457, n31458, n31459, n31461, n31464, n31465,
         n31466, n31470, n31471, n31473, n31474, n31475, n31476, n31477,
         n31480, n31481, n31483, n31484, n31485, n31486, n31488, n31490,
         n31492, n31494, n31495, n31496, n31498, n31499, n31500, n31502,
         n31504, n31505, n31507, n31508, n31509, n31511, n31512, n31513,
         n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522,
         n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530,
         n31532, n31533, n31534, n31535, n31537, n31538, n31539, n31540,
         n31541, n31542, n31543, n31545, n31546, n31547, n31548, n31549,
         n31550, n31551, n31552, n31554, n31555, n31557, n31558, n31559,
         n31562, n31563, n31564, n31565, n31566, n31568, n31569, n31570,
         n31571, n31573, n31574, n31575, n31576, n31579, n31580, n31581,
         n31582, n31583, n31584, n31585, n31586, n31587, n31591, n31594,
         n31595, n31596, n31597, n31598, n31599, n31601, n31602, n31603,
         n31604, n31605, n31606, n31607, n31608, n31611, n31612, n31615,
         n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31624,
         n31625, n31626, n31627, n31628, n31629, n31630, n31633, n31634,
         n31636, n31637, n31638, n31640, n31643, n31644, n31647, n31648,
         n31649, n31650, n31651, n31652, n31654, n31655, n31656, n31657,
         n31660, n31661, n31662, n31663, n31664, n31665, n31667, n31668,
         n31669, n31670, n31672, n31673, n31678, n31679, n31680, n31682,
         n31683, n31684, n31685, n31688, n31689, n31692, n31693, n31695,
         n31696, n31697, n31698, n31699, n31701, n31702, n31704, n31705,
         n31707, n31708, n31710, n31711, n31712, n31713, n31714, n31716,
         n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
         n31725, n31726, n31727, n31731, n31734, n31735, n31736, n31737,
         n31739, n31743, n31744, n31745, n31748, n31749, n31751, n31752,
         n31755, n31759, n31760, n31762, n31764, n31765, n31766, n31767,
         n31769, n31771, n31772, n31773, n31774, n31775, n31777, n31778,
         n31779, n31780, n31781, n31782, n31784, n31785, n31786, n31787,
         n31788, n31790, n31791, n31794, n31795, n31796, n31797, n31798,
         n31799, n31801, n31805, n31806, n31807, n31808, n31809, n31810,
         n31811, n31812, n31815, n31816, n31820, n31821, n31822, n31823,
         n31824, n31825, n31827, n31829, n31830, n31831, n31832, n31835,
         n31836, n31838, n31840, n31841, n31842, n31843, n31845, n31846,
         n31847, n31848, n31849, n31851, n31852, n31854, n31855, n31857,
         n31859, n31860, n31861, n31862, n31863, n31867, n31869, n31871,
         n31872, n31875, n31876, n31880, n31882, n31883, n31887, n31888,
         n31889, n31891, n31893, n31895, n31897, n31898, n31899, n31900,
         n31904, n31906, n31908, n31909, n31911, n31912, n31913, n31914,
         n31916, n31917, n31918, n31919, n31920, n31921, n31924, n31925,
         n31926, n31927, n31931, n31932, n31933, n31934, n31937, n31939,
         n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947,
         n31948, n31949, n31951, n31953, n31954, n31955, n31958, n31959,
         n31960, n31963, n31964, n31965, n31966, n31967, n31968, n31971,
         n31972, n31975, n31976, n31978, n31980, n31982, n31983, n31984,
         n31985, n31986, n31987, n31994, n31996, n31997, n31999, n32001,
         n32002, n32003, n32004, n32005, n32006, n32009, n32010, n32011,
         n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019,
         n32020, n32021, n32022, n32024, n32025, n32026, n32032, n32033,
         n32035, n32036, n32039, n32040, n32041, n32042, n32043, n32044,
         n32045, n32046, n32049, n32050, n32051, n32052, n32053, n32054,
         n32056, n32057, n32059, n32060, n32061, n32062, n32063, n32064,
         n32068, n32069, n32071, n32072, n32073, n32075, n32076, n32077,
         n32079, n32080, n32081, n32083, n32084, n32085, n32087, n32089,
         n32090, n32091, n32092, n32093, n32095, n32096, n32097, n32099,
         n32101, n32103, n32105, n32106, n32107, n32109, n32110, n32111,
         n32113, n32114, n32118, n32120, n32122, n32123, n32125, n32126,
         n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134,
         n32135, n32136, n32137, n32138, n32141, n32142, n32146, n32149,
         n32150, n32151, n32152, n32153, n32154, n32156, n32157, n32158,
         n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166,
         n32167, n32168, n32169, n32170, n32172, n32174, n32175, n32176,
         n32178, n32181, n32182, n32183, n32184, n32185, n32186, n32188,
         n32189, n32190, n32191, n32192, n32193, n32195, n32196, n32197,
         n32200, n32202, n32203, n32204, n32205, n32206, n32207, n32208,
         n32209, n32210, n32211, n32215, n32216, n32217, n32218, n32219,
         n32221, n32223, n32226, n32227, n32228, n32230, n32232, n32233,
         n32234, n32235, n32236, n32239, n32243, n32245, n32246, n32247,
         n32248, n32250, n32251, n32253, n32255, n32256, n32258, n32259,
         n32260, n32261, n32262, n32263, n32266, n32267, n32268, n32270,
         n32273, n32274, n32275, n32276, n32278, n32279, n32280, n32282,
         n32283, n32284, n32286, n32288, n32290, n32291, n32292, n32293,
         n32294, n32297, n32298, n32301, n32302, n32303, n32304, n32306,
         n32308, n32309, n32310, n32312, n32313, n32314, n32315, n32317,
         n32318, n32319, n32322, n32324, n32325, n32326, n32327, n32331,
         n32332, n32333, n32335, n32337, n32338, n32339, n32340, n32343,
         n32344, n32345, n32346, n32347, n32348, n32349, n32351, n32352,
         n32353, n32354, n32355, n32358, n32359, n32360, n32361, n32362,
         n32363, n32365, n32366, n32367, n32368, n32369, n32370, n32372,
         n32374, n32375, n32376, n32377, n32380, n32382, n32383, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32394, n32396,
         n32397, n32398, n32400, n32401, n32402, n32403, n32404, n32406,
         n32407, n32408, n32410, n32411, n32412, n32413, n32415, n32418,
         n32419, n32420, n32423, n32424, n32425, n32427, n32430, n32431,
         n32432, n32433, n32434, n32436, n32440, n32441, n32442, n32443,
         n32444, n32446, n32447, n32448, n32449, n32450, n32452, n32456,
         n32457, n32460, n32462, n32463, n32464, n32465, n32466, n32467,
         n32468, n32469, n32470, n32471, n32472, n32474, n32477, n32478,
         n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486,
         n32487, n32488, n32490, n32491, n32492, n32494, n32495, n32497,
         n32498, n32499, n32504, n32505, n32506, n32507, n32508, n32510,
         n32512, n32515, n32516, n32518, n32519, n32520, n32524, n32525,
         n32526, n32527, n32528, n32531, n32532, n32534, n32535, n32536,
         n32537, n32539, n32540, n32542, n32543, n32544, n32545, n32546,
         n32548, n32549, n32551, n32552, n32555, n32556, n32557, n32558,
         n32559, n32562, n32563, n32566, n32567, n32570, n32571, n32572,
         n32573, n32574, n32575, n32577, n32579, n32580, n32581, n32583,
         n32584, n32585, n32586, n32588, n32590, n32594, n32595, n32596,
         n32598, n32599, n32601, n32602, n32604, n32607, n32608, n32609,
         n32610, n32613, n32614, n32615, n32616, n32617, n32618, n32619,
         n32620, n32621, n32622, n32623, n32625, n32626, n32628, n32630,
         n32631, n32633, n32634, n32636, n32637, n32638, n32639, n32640,
         n32641, n32643, n32644, n32646, n32647, n32648, n32649, n32650,
         n32651, n32654, n32657, n32658, n32660, n32661, n32662, n32663,
         n32664, n32666, n32667, n32668, n32669, n32670, n32671, n32675,
         n32676, n32677, n32678, n32681, n32682, n32683, n32684, n32685,
         n32686, n32689, n32690, n32691, n32693, n32695, n32696, n32697,
         n32698, n32699, n32702, n32703, n32704, n32705, n32706, n32708,
         n32712, n32714, n32718, n32719, n32720, n32721, n32722, n32725,
         n32727, n32728, n32734, n32740, n32741, n32742, n32743, n32745,
         n32746, n32747, n32748, n32750, n32752, n32753, n32755, n32756,
         n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32765,
         n32766, n32767, n32768, n32769, n32771, n32773, n32775, n32776,
         n32777, n32778, n32779, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32789, n32790, n32791, n32795, n32796, n32797,
         n32798, n32799, n32800, n32802, n32803, n32805, n32806, n32807,
         n32808, n32811, n32813, n32814, n32815, n32817, n32818, n32820,
         n32821, n32822, n32825, n32826, n32827, n32829, n32831, n32832,
         n32833, n32836, n32837, n32838, n32839, n32842, n32843, n32844,
         n32847, n32849, n32850, n32851, n32852, n32853, n32854, n32855,
         n32856, n32857, n32858, n32860, n32861, n32863, n32865, n32866,
         n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32877,
         n32878, n32879, n32881, n32882, n32883, n32884, n32885, n32886,
         n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896,
         n32897, n32898, n32899, n32902, n32903, n32904, n32906, n32909,
         n32910, n32911, n32913, n32915, n32916, n32917, n32918, n32924,
         n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932,
         n32933, n32934, n32937, n32938, n32940, n32941, n32942, n32943,
         n32944, n32945, n32946, n32948, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32958, n32959, n32960, n32961, n32962,
         n32963, n32971, n32972, n32973, n32974, n32976, n32977, n32979,
         n32980, n32981, n32983, n32984, n32985, n32986, n32987, n32989,
         n32993, n32994, n32999, n33001, n33002, n33004, n33005, n33006,
         n33007, n33008, n33010, n33011, n33012, n33013, n33015, n33016,
         n33017, n33020, n33022, n33023, n33025, n33026, n33027, n33028,
         n33029, n33030, n33032, n33034, n33036, n33037, n33038, n33039,
         n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048,
         n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056,
         n33057, n33058, n33059, n33061, n33062, n33063, n33067, n33070,
         n33071, n33072, n33073, n33074, n33075, n33077, n33080, n33081,
         n33082, n33083, n33085, n33086, n33087, n33088, n33091, n33092,
         n33093, n33094, n33097, n33098, n33100, n33101, n33102, n33104,
         n33106, n33107, n33108, n33109, n33111, n33112, n33113, n33114,
         n33115, n33116, n33118, n33120, n33121, n33123, n33125, n33128,
         n33129, n33130, n33131, n33132, n33133, n33135, n33138, n33139,
         n33140, n33141, n33142, n33144, n33145, n33146, n33147, n33148,
         n33151, n33152, n33153, n33154, n33155, n33156, n33158, n33160,
         n33161, n33163, n33165, n33166, n33168, n33170, n33176, n33177,
         n33178, n33179, n33180, n33182, n33183, n33184, n33185, n33186,
         n33187, n33188, n33190, n33192, n33193, n33194, n33195, n33196,
         n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204,
         n33206, n33207, n33208, n33209, n33215, n33216, n33217, n33218,
         n33219, n33220, n33223, n33224, n33226, n33227, n33228, n33229,
         n33230, n33231, n33232, n33233, n33234, n33235, n33237, n33239,
         n33240, n33242, n33243, n33244, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33254, n33255, n33256, n33257, n33258,
         n33261, n33262, n33263, n33264, n33266, n33267, n33268, n33270,
         n33271, n33272, n33273, n33276, n33277, n33278, n33279, n33280,
         n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288,
         n33289, n33291, n33292, n33293, n33295, n33296, n33297, n33299,
         n33300, n33301, n33302, n33303, n33304, n33307, n33308, n33309,
         n33310, n33311, n33313, n33314, n33315, n33316, n33317, n33318,
         n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
         n33327, n33328, n33331, n33333, n33334, n33335, n33336, n33337,
         n33340, n33344, n33346, n33347, n33348, n33349, n33350, n33352,
         n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360,
         n33361, n33362, n33363, n33364, n33365, n33366, n33368, n33369,
         n33370, n33371, n33372, n33373, n33375, n33376, n33379, n33380,
         n33383, n33384, n33385, n33387, n33388, n33389, n33392, n33393,
         n33394, n33395, n33396, n33398, n33399, n33400, n33401, n33402,
         n33403, n33404, n33405, n33407, n33409, n33410, n33412, n33413,
         n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33422,
         n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33431,
         n33433, n33434, n33436, n33437, n33438, n33439, n33440, n33442,
         n33446, n33449, n33450, n33452, n33453, n33455, n33456, n33457,
         n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466,
         n33468, n33470, n33472, n33473, n33474, n33476, n33478, n33479,
         n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487,
         n33488, n33489, n33491, n33493, n33495, n33496, n33498, n33500,
         n33503, n33504, n33505, n33506, n33509, n33510, n33511, n33512,
         n33513, n33514, n33515, n33516, n33517, n33519, n33520, n33521,
         n33522, n33524, n33526, n33527, n33528, n33529, n33530, n33531,
         n33532, n33533, n33534, n33535, n33538, n33539, n33541, n33544,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33557, n33558, n33559, n33561, n33563, n33565,
         n33566, n33567, n33568, n33569, n33571, n33572, n33573, n33574,
         n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33584,
         n33585, n33586, n33587, n33591, n33593, n33594, n33595, n33597,
         n33598, n33599, n33601, n33603, n33604, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33616, n33619, n33620,
         n33621, n33622, n33623, n33625, n33628, n33629, n33630, n33631,
         n33633, n33636, n33638, n33640, n33642, n33643, n33644, n33645,
         n33646, n33647, n33648, n33649, n33650, n33651, n33653, n33655,
         n33656, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33671, n33672, n33674, n33675,
         n33676, n33677, n33678, n33679, n33686, n33687, n33689, n33690,
         n33693, n33694, n33695, n33696, n33697, n33698, n33700, n33701,
         n33702, n33703, n33705, n33706, n33707, n33708, n33709, n33712,
         n33713, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33724, n33725, n33726, n33727, n33730, n33731, n33733,
         n33734, n33735, n33736, n33737, n33738, n33743, n33745, n33746,
         n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754,
         n33755, n33756, n33757, n33758, n33759, n33760, n33763, n33764,
         n33765, n33766, n33767, n33771, n33773, n33775, n33776, n33777,
         n33780, n33781, n33782, n33784, n33785, n33786, n33788, n33789,
         n33792, n33793, n33795, n33799, n33802, n33803, n33804, n33805,
         n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813,
         n33815, n33816, n33817, n33818, n33821, n33824, n33825, n33826,
         n33829, n33831, n33832, n33833, n33834, n33837, n33839, n33840,
         n33841, n33842, n33843, n33844, n33845, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33855, n33856, n33858, n33859,
         n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867,
         n33868, n33869, n33870, n33871, n33876, n33879, n33883, n33885,
         n33886, n33887, n33888, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33899, n33902, n33904, n33905, n33906,
         n33908, n33909, n33910, n33911, n33912, n33913, n33916, n33919,
         n33921, n33924, n33925, n33926, n33928, n33929, n33931, n33933,
         n33934, n33935, n33936, n33937, n33939, n33944, n33945, n33946,
         n33947, n33948, n33949, n33950, n33952, n33954, n33955, n33956,
         n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964,
         n33965, n33966, n33967, n33968, n33969, n33972, n33973, n33976,
         n33978, n33979, n33980, n33981, n33986, n33987, n33990, n33993,
         n33995, n33996, n33997, n33999, n34000, n34001, n34003, n34004,
         n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012,
         n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020,
         n34021, n34022, n34023, n34024, n34025, n34027, n34028, n34030,
         n34031, n34032, n34033, n34034, n34036, n34037, n34038, n34039,
         n34040, n34041, n34042, n34043, n34044, n34046, n34047, n34048,
         n34049, n34050, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34080, n34081, n34082,
         n34083, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
         n34092, n34094, n34096, n34097, n34099, n34103, n34104, n34105,
         n34108, n34111, n34112, n34113, n34114, n34115, n34116, n34117,
         n34120, n34121, n34122, n34123, n34124, n34126, n34128, n34129,
         n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
         n34139, n34141, n34142, n34143, n34144, n34145, n34147, n34148,
         n34149, n34150, n34151, n34152, n34153, n34154, n34156, n34157,
         n34160, n34161, n34162, n34163, n34165, n34166, n34167, n34170,
         n34171, n34172, n34173, n34175, n34176, n34177, n34178, n34179,
         n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34188,
         n34189, n34190, n34192, n34193, n34194, n34195, n34196, n34197,
         n34198, n34199, n34200, n34201, n34202, n34203, n34205, n34206,
         n34208, n34210, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34220, n34221, n34223, n34224, n34225, n34226, n34227,
         n34228, n34231, n34233, n34235, n34237, n34238, n34239, n34244,
         n34245, n34246, n34247, n34249, n34250, n34251, n34252, n34254,
         n34256, n34257, n34259, n34260, n34261, n34262, n34263, n34264,
         n34265, n34266, n34267, n34268, n34269, n34270, n34272, n34274,
         n34275, n34276, n34277, n34279, n34282, n34283, n34284, n34285,
         n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34296,
         n34297, n34298, n34299, n34301, n34303, n34305, n34306, n34307,
         n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34317,
         n34319, n34323, n34324, n34325, n34326, n34329, n34330, n34332,
         n34335, n34336, n34337, n34339, n34340, n34342, n34343, n34344,
         n34345, n34347, n34350, n34351, n34352, n34354, n34357, n34358,
         n34359, n34360, n34365, n34366, n34368, n34370, n34371, n34372,
         n34373, n34374, n34375, n34377, n34378, n34379, n34382, n34383,
         n34384, n34386, n34387, n34389, n34391, n34392, n34393, n34394,
         n34395, n34396, n34397, n34398, n34399, n34401, n34402, n34404,
         n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34413,
         n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421,
         n34422, n34424, n34426, n34427, n34428, n34430, n34433, n34435,
         n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34446,
         n34447, n34448, n34450, n34451, n34452, n34453, n34454, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34472, n34473, n34474,
         n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482,
         n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490,
         n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498,
         n34499, n34501, n34503, n34504, n34506, n34510, n34512, n34513,
         n34514, n34515, n34516, n34518, n34519, n34520, n34521, n34522,
         n34524, n34525, n34526, n34531, n34532, n34533, n34534, n34535,
         n34538, n34539, n34540, n34541, n34544, n34545, n34546, n34547,
         n34549, n34552, n34553, n34554, n34557, n34558, n34559, n34561,
         n34562, n34564, n34565, n34567, n34568, n34569, n34570, n34571,
         n34572, n34573, n34574, n34575, n34576, n34577, n34579, n34580,
         n34581, n34583, n34585, n34586, n34587, n34589, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34601, n34602,
         n34603, n34604, n34606, n34608, n34609, n34610, n34611, n34613,
         n34615, n34616, n34618, n34619, n34620, n34621, n34622, n34627,
         n34630, n34632, n34634, n34635, n34636, n34637, n34638, n34639,
         n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648,
         n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656,
         n34658, n34660, n34662, n34663, n34664, n34666, n34667, n34668,
         n34669, n34670, n34671, n34672, n34673, n34678, n34680, n34681,
         n34682, n34683, n34685, n34686, n34688, n34689, n34690, n34691,
         n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699,
         n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709,
         n34711, n34712, n34713, n34715, n34716, n34717, n34718, n34719,
         n34720, n34722, n34723, n34724, n34726, n34727, n34728, n34733,
         n34737, n34738, n34739, n34740, n34742, n34743, n34745, n34746,
         n34747, n34750, n34751, n34752, n34753, n34755, n34757, n34758,
         n34760, n34761, n34762, n34763, n34764, n34766, n34767, n34768,
         n34769, n34770, n34772, n34773, n34774, n34776, n34777, n34778,
         n34780, n34781, n34783, n34785, n34786, n34787, n34788, n34789,
         n34790, n34793, n34794, n34795, n34796, n34799, n34800, n34801,
         n34802, n34804, n34805, n34806, n34808, n34809, n34811, n34812,
         n34813, n34814, n34815, n34817, n34819, n34820, n34821, n34822,
         n34823, n34825, n34826, n34828, n34829, n34830, n34832, n34836,
         n34837, n34838, n34840, n34841, n34842, n34843, n34844, n34846,
         n34847, n34848, n34849, n34850, n34851, n34853, n34854, n34855,
         n34856, n34857, n34858, n34861, n34863, n34866, n34867, n34868,
         n34869, n34870, n34871, n34876, n34877, n34878, n34881, n34882,
         n34883, n34884, n34885, n34886, n34889, n34890, n34891, n34892,
         n34893, n34894, n34895, n34897, n34898, n34899, n34900, n34901,
         n34902, n34903, n34904, n34905, n34906, n34908, n34909, n34911,
         n34912, n34913, n34914, n34915, n34918, n34920, n34922, n34923,
         n34924, n34925, n34926, n34930, n34931, n34932, n34933, n34934,
         n34935, n34938, n34939, n34940, n34942, n34943, n34944, n34945,
         n34947, n34948, n34949, n34952, n34953, n34955, n34956, n34957,
         n34958, n34959, n34961, n34962, n34963, n34964, n34965, n34966,
         n34967, n34969, n34972, n34973, n34974, n34977, n34979, n34981,
         n34982, n34983, n34984, n34985, n34986, n34987, n34989, n34990,
         n34993, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35003, n35004, n35005, n35006, n35007, n35010, n35012, n35013,
         n35014, n35015, n35016, n35017, n35018, n35019, n35021, n35022,
         n35023, n35025, n35026, n35027, n35028, n35029, n35030, n35031,
         n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039,
         n35040, n35042, n35043, n35045, n35046, n35047, n35048, n35049,
         n35051, n35053, n35054, n35055, n35056, n35057, n35059, n35060,
         n35061, n35062, n35063, n35064, n35065, n35067, n35068, n35070,
         n35071, n35072, n35073, n35075, n35076, n35077, n35078, n35079,
         n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087,
         n35088, n35089, n35092, n35093, n35095, n35096, n35097, n35098,
         n35099, n35102, n35103, n35105, n35107, n35108, n35109, n35112,
         n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120,
         n35121, n35122, n35123, n35124, n35128, n35129, n35130, n35134,
         n35135, n35137, n35138, n35139, n35140, n35141, n35142, n35143,
         n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151,
         n35153, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35168, n35169, n35170, n35171,
         n35172, n35173, n35175, n35176, n35177, n35178, n35179, n35180,
         n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188,
         n35189, n35190, n35191, n35192, n35193, n35194, n35196, n35197,
         n35198, n35199, n35200, n35202, n35203, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35224, n35225, n35227,
         n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235,
         n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244,
         n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252,
         n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260,
         n35262, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
         n35271, n35272, n35273, n35274, n35278, n35279, n35280, n35281,
         n35282, n35285, n35286, n35287, n35288, n35290, n35293, n35294,
         n35295, n35296, n35297, n35299, n35300, n35301, n35302, n35303,
         n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35317,
         n35318, n35320, n35321, n35322, n35323, n35324, n35326, n35327,
         n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336,
         n35339, n35340, n35342, n35343, n35344, n35345, n35347, n35348,
         n35349, n35350, n35351, n35353, n35355, n35357, n35359, n35360,
         n35361, n35362, n35363, n35367, n35368, n35369, n35370, n35371,
         n35373, n35374, n35376, n35377, n35379, n35380, n35381, n35384,
         n35386, n35387, n35389, n35390, n35391, n35392, n35394, n35395,
         n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404,
         n35405, n35407, n35409, n35410, n35414, n35415, n35417, n35419,
         n35420, n35421, n35422, n35423, n35424, n35425, n35427, n35429,
         n35431, n35434, n35435, n35436, n35437, n35438, n35439, n35440,
         n35441, n35442, n35443, n35445, n35446, n35447, n35448, n35449,
         n35450, n35452, n35453, n35454, n35455, n35457, n35462, n35463,
         n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471,
         n35472, n35473, n35474, n35476, n35477, n35478, n35479, n35480,
         n35481, n35483, n35485, n35487, n35489, n35490, n35491, n35492,
         n35494, n35495, n35496, n35498, n35499, n35500, n35501, n35502,
         n35503, n35504, n35505, n35506, n35507, n35508, n35510, n35511,
         n35513, n35514, n35517, n35519, n35520, n35521, n35523, n35525,
         n35526, n35528, n35529, n35532, n35534, n35535, n35536, n35537,
         n35541, n35542, n35543, n35544, n35545, n35547, n35548, n35549,
         n35550, n35551, n35553, n35554, n35556, n35559, n35560, n35561,
         n35563, n35564, n35566, n35567, n35568, n35569, n35570, n35571,
         n35572, n35573, n35574, n35576, n35577, n35578, n35579, n35580,
         n35583, n35584, n35585, n35586, n35588, n35590, n35591, n35594,
         n35595, n35596, n35598, n35599, n35600, n35601, n35603, n35604,
         n35607, n35608, n35610, n35611, n35612, n35613, n35614, n35616,
         n35617, n35618, n35619, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35629, n35630, n35631, n35632, n35633, n35636,
         n35637, n35639, n35640, n35642, n35644, n35645, n35646, n35647,
         n35648, n35649, n35651, n35652, n35653, n35654, n35655, n35656,
         n35657, n35658, n35659, n35660, n35663, n35664, n35665, n35666,
         n35667, n35668, n35670, n35671, n35673, n35675, n35676, n35677,
         n35678, n35679, n35681, n35684, n35685, n35686, n35687, n35688,
         n35689, n35690, n35693, n35694, n35695, n35696, n35697, n35699,
         n35702, n35704, n35705, n35706, n35707, n35708, n35709, n35710,
         n35711, n35712, n35715, n35718, n35720, n35721, n35722, n35723,
         n35724, n35726, n35727, n35728, n35729, n35730, n35731, n35732,
         n35733, n35734, n35735, n35737, n35741, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35752, n35753, n35754,
         n35755, n35756, n35757, n35758, n35760, n35761, n35762, n35763,
         n35764, n35765, n35766, n35767, n35768, n35769, n35771, n35772,
         n35774, n35776, n35777, n35779, n35780, n35781, n35782, n35784,
         n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792,
         n35793, n35794, n35795, n35796, n35801, n35802, n35803, n35804,
         n35805, n35806, n35808, n35809, n35810, n35811, n35812, n35813,
         n35814, n35815, n35816, n35818, n35819, n35820, n35821, n35822,
         n35823, n35824, n35825, n35826, n35827, n35828, n35830, n35832,
         n35833, n35834, n35835, n35836, n35837, n35839, n35840, n35841,
         n35842, n35843, n35844, n35846, n35847, n35848, n35849, n35851,
         n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859,
         n35860, n35862, n35863, n35864, n35867, n35868, n35869, n35870,
         n35871, n35872, n35873, n35874, n35875, n35877, n35878, n35879,
         n35880, n35881, n35882, n35883, n35885, n35886, n35887, n35888,
         n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896,
         n35897, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35908, n35909, n35910, n35911, n35912, n35914, n35915,
         n35916, n35917, n35918, n35919, n35920, n35921, n35923, n35924,
         n35925, n35926, n35928, n35931, n35932, n35935, n35936, n35938,
         n35939, n35941, n35942, n35943, n35944, n35947, n35948, n35950,
         n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959,
         n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967,
         n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975,
         n35976, n35977, n35978, n35979, n35981, n35983, n35984, n35985,
         n35986, n35987, n35988, n35990, n35992, n35993, n35994, n35996,
         n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004,
         n36005, n36006, n36007, n36008, n36011, n36013, n36016, n36017,
         n36019, n36020, n36021, n36022, n36023, n36024, n36026, n36027,
         n36029, n36030, n36031, n36032, n36034, n36035, n36036, n36038,
         n36039, n36040, n36041, n36043, n36044, n36046, n36048, n36050,
         n36051, n36052, n36053, n36055, n36057, n36058, n36059, n36060,
         n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069,
         n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078,
         n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086,
         n36087, n36090, n36091, n36092, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36117,
         n36119, n36120, n36123, n36124, n36125, n36126, n36127, n36128,
         n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136,
         n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144,
         n36145, n36146, n36147, n36150, n36151, n36152, n36154, n36157,
         n36159, n36160, n36162, n36163, n36164, n36165, n36166, n36167,
         n36168, n36170, n36171, n36172, n36173, n36175, n36176, n36177,
         n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187,
         n36188, n36190, n36191, n36193, n36194, n36195, n36196, n36197,
         n36199, n36200, n36201, n36203, n36204, n36205, n36206, n36207,
         n36209, n36210, n36211, n36212, n36214, n36216, n36217, n36218,
         n36219, n36222, n36223, n36224, n36225, n36226, n36227, n36228,
         n36229, n36230, n36231, n36232, n36233, n36234, n36236, n36237,
         n36238, n36239, n36240, n36241, n36243, n36244, n36245, n36246,
         n36247, n36248, n36249, n36250, n36251, n36253, n36254, n36255,
         n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264,
         n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272,
         n36273, n36275, n36277, n36279, n36280, n36281, n36283, n36284,
         n36286, n36287, n36289, n36290, n36291, n36292, n36293, n36295,
         n36296, n36297, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36313, n36314,
         n36317, n36320, n36321, n36322, n36323, n36324, n36325, n36326,
         n36327, n36328, n36329, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36348, n36349, n36351, n36352, n36353, n36354, n36355,
         n36357, n36358, n36360, n36361, n36362, n36363, n36364, n36365,
         n36366, n36368, n36369, n36371, n36372, n36373, n36374, n36375,
         n36376, n36377, n36378, n36379, n36380, n36382, n36383, n36384,
         n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392,
         n36393, n36394, n36395, n36396, n36397, n36400, n36402, n36403,
         n36404, n36406, n36407, n36408, n36410, n36411, n36412, n36413,
         n36414, n36415, n36416, n36418, n36420, n36421, n36422, n36423,
         n36424, n36425, n36426, n36428, n36429, n36430, n36431, n36433,
         n36434, n36435, n36436, n36441, n36442, n36443, n36444, n36445,
         n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453,
         n36454, n36455, n36456, n36457, n36458, n36459, n36460, n36461,
         n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470,
         n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
         n36480, n36481, n36483, n36485, n36486, n36487, n36488, n36490,
         n36491, n36492, n36493, n36494, n36496, n36497, n36498, n36499,
         n36500, n36501, n36502, n36506, n36507, n36508, n36509, n36510,
         n36511, n36513, n36514, n36515, n36516, n36517, n36518, n36519,
         n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527,
         n36528, n36529, n36530, n36532, n36535, n36537, n36538, n36539,
         n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36548,
         n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556,
         n36558, n36559, n36560, n36561, n36563, n36564, n36566, n36567,
         n36568, n36569, n36571, n36572, n36573, n36574, n36575, n36576,
         n36577, n36578, n36579, n36581, n36582, n36583, n36584, n36585,
         n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594,
         n36595, n36596, n36598, n36601, n36602, n36603, n36604, n36605,
         n36606, n36607, n36608, n36609, n36611, n36612, n36613, n36615,
         n36616, n36617, n36618, n36620, n36621, n36622, n36623, n36624,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36637, n36638, n36639, n36640, n36641, n36643,
         n36644, n36645, n36646, n36647, n36649, n36651, n36654, n36655,
         n36656, n36658, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36668, n36669, n36671, n36672, n36673, n36674, n36676,
         n36677, n36678, n36679, n36680, n36682, n36683, n36685, n36686,
         n36687, n36689, n36690, n36691, n36692, n36693, n36694, n36696,
         n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36705,
         n36706, n36707, n36708, n36709, n36711, n36712, n36716, n36717,
         n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725,
         n36726, n36727, n36728, n36729, n36730, n36731, n36734, n36735,
         n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743,
         n36744, n36745, n36746, n36748, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36769, n36772,
         n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780,
         n36781, n36782, n36783, n36785, n36786, n36787, n36788, n36789,
         n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797,
         n36798, n36799, n36800, n36801, n36803, n36804, n36805, n36806,
         n36807, n36808, n36809, n36810, n36812, n36814, n36815, n36816,
         n36817, n36818, n36819, n36821, n36822, n36824, n36827, n36828,
         n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36837,
         n36838, n36839, n36840, n36842, n36843, n36844, n36846, n36847,
         n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36856,
         n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864,
         n36865, n36866, n36867, n36868, n36869, n36871, n36872, n36873,
         n36876, n36877, n36878, n36880, n36882, n36884, n36885, n36886,
         n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894,
         n36895, n36896, n36897, n36899, n36900, n36902, n36903, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36918, n36919, n36920, n36922, n36923,
         n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931,
         n36932, n36935, n36936, n36938, n36939, n36940, n36941, n36942,
         n36944, n36945, n36946, n36947, n36949, n36951, n36952, n36953,
         n36954, n36955, n36957, n36958, n36959, n36960, n36961, n36962,
         n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
         n36972, n36974, n36976, n36977, n36979, n36980, n36981, n36984,
         n36985, n36986, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37001, n37002,
         n37003, n37005, n37006, n37007, n37008, n37010, n37011, n37012,
         n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020,
         n37021, n37023, n37024, n37025, n37026, n37027, n37028, n37030,
         n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038,
         n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37047,
         n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055,
         n37056, n37057, n37059, n37060, n37061, n37062, n37063, n37064,
         n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072,
         n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080,
         n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088,
         n37089, n37092, n37093, n37094, n37095, n37096, n37097, n37098,
         n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106,
         n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114,
         n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122,
         n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130,
         n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138,
         n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146,
         n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154,
         n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
         n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170,
         n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178,
         n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186,
         n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194,
         n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202,
         n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210,
         n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218,
         n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226,
         n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
         n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242,
         n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250,
         n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258,
         n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266,
         n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274,
         n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282,
         n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290,
         n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298,
         n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
         n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314,
         n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322,
         n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331,
         n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339,
         n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347,
         n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355,
         n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363,
         n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371,
         n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379,
         n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387,
         n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395,
         n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403,
         n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411,
         n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419,
         n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427,
         n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435,
         n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443,
         n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451,
         n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459,
         n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467,
         n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475,
         n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483,
         n37484, n37485, n37486, n37487, n37489, n37490, n37491, n37492,
         n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500,
         n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508,
         n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516,
         n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524,
         n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532,
         n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540,
         n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548,
         n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556,
         n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564,
         n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572,
         n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580,
         n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588,
         n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596,
         n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604,
         n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612,
         n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620,
         n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628,
         n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636,
         n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644,
         n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652,
         n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660,
         n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668,
         n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676,
         n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684,
         n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692,
         n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700,
         n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708,
         n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716,
         n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724,
         n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732,
         n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740,
         n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748,
         n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756,
         n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764,
         n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772,
         n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780,
         n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788,
         n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796,
         n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804,
         n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812,
         n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820,
         n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828,
         n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836,
         n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844,
         n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852,
         n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860,
         n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868,
         n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876,
         n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884,
         n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892,
         n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900,
         n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908,
         n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916,
         n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925,
         n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933,
         n37934, n37935, n37936, n37937, n37938, n37939, n37940, n37941,
         n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949,
         n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957,
         n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965,
         n37966, n37967, n37968, n37969, n37970, n37971, n37972, n37973,
         n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981,
         n37982, n37983, n37984, n37985, n37986, n37987, n37988, n37989,
         n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997,
         n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005,
         n38006, n38007, n38008, n38009, n38010, n38011, n38012, n38013,
         n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021,
         n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029,
         n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037,
         n38038, n38039, n38040, n38041, n38042, n38043, n38044, n38045,
         n38046, n38047, n38048, n38049, n38050, n38051, n38052, n38053,
         n38054, n38055, n38056, n38057, n38058, n38059, n38060, n38061,
         n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069,
         n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077,
         n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085,
         n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093,
         n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101,
         n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109,
         n38110, n38111, n38112, n38113, n38114, n38115, n38116, n38117,
         n38118, n38119, n38120, n38121, n38122, n38123, n38124, n38125,
         n38126, n38127, n38128, n38129, n38130, n38131, n38132, n38133,
         n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141,
         n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149,
         n38150, n38151, n38152, n38153, n38154, n38155, n38156, n38157,
         n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165,
         n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173,
         n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181,
         n38182, n38183, n38184, n38185, n38186, n38187, n38188, n38189,
         n38190, n38191, n38192, n38193, n38194, n38195, n38196, n38197,
         n38198, n38199, n38200, n38201, n38202, n38203, n38204, n38205,
         n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213,
         n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221,
         n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229,
         n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237,
         n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245,
         n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253,
         n38254, n38255, n38256, n38257, n38258, n38259, n38260, n38261,
         n38262, n38263, n38264, n38265, n38266, n38267, n38268, n38269,
         n38270, n38271, n38272, n38273, n38274, n38275, n38276, n38277,
         n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285,
         n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293,
         n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301,
         n38302, n38303, n38305, n38306, n38307, n38308, n38309, n38310,
         n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318,
         n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326,
         n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334,
         n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342,
         n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350,
         n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358,
         n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
         n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374,
         n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382,
         n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390,
         n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398,
         n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406,
         n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414,
         n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
         n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430,
         n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
         n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446,
         n38448, n38450, n38451, n38452, n38453, n38454, n38455, n38456,
         n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464,
         n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472,
         n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480,
         n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488,
         n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496,
         n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504,
         n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
         n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520,
         n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528,
         n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536,
         n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544,
         n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552,
         n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560,
         n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568,
         n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576,
         n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
         n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592,
         n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600,
         n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608,
         n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616,
         n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624,
         n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632,
         n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640,
         n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648,
         n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656,
         n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664,
         n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672,
         n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680,
         n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688,
         n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696,
         n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704,
         n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712,
         n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720,
         n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728,
         n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736,
         n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744,
         n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752,
         n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760,
         n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768,
         n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776,
         n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784,
         n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792,
         n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
         n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808,
         n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816,
         n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824,
         n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832,
         n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840,
         n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848,
         n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856,
         n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864,
         n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872,
         n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880,
         n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888,
         n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896,
         n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904,
         n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912,
         n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920,
         n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928,
         n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936,
         n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944,
         n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952,
         n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960,
         n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968,
         n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976,
         n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984,
         n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992,
         n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000,
         n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008,
         n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016,
         n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024,
         n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032,
         n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040,
         n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048,
         n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056,
         n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064,
         n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072,
         n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080,
         n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088,
         n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096,
         n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104,
         n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112,
         n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120,
         n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128,
         n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136,
         n39137, n39138, n39139, n39140, n39141, n39142, n39143, n39144,
         n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152,
         n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160,
         n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168,
         n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176,
         n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184,
         n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192,
         n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200,
         n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208,
         n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216,
         n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224,
         n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232,
         n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240,
         n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248,
         n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256,
         n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264,
         n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272,
         n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280,
         n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288,
         n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296,
         n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304,
         n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312,
         n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320,
         n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328,
         n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336,
         n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344,
         n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352,
         n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360,
         n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368,
         n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376,
         n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384,
         n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392,
         n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400,
         n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408,
         n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416,
         n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424,
         n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432,
         n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440,
         n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448,
         n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456,
         n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464,
         n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472,
         n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480,
         n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488,
         n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496,
         n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504,
         n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512,
         n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520,
         n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528,
         n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
         n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
         n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552,
         n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560,
         n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568,
         n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576,
         n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584,
         n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592,
         n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600,
         n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608,
         n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616,
         n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624,
         n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632,
         n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640,
         n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648,
         n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656,
         n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664,
         n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672,
         n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680,
         n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688,
         n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696,
         n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704,
         n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712,
         n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720,
         n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728,
         n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
         n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744,
         n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752,
         n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760,
         n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768,
         n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776,
         n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784,
         n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
         n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800,
         n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808,
         n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816,
         n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824,
         n39825, n39826, n39827, n39828, n39829, n39830;

  INV_X1 U42 ( .I(n29438), .ZN(n1383) );
  NAND2_X1 U65 ( .A1(n17238), .A2(n30229), .ZN(n18043) );
  NOR2_X1 U73 ( .A1(n29491), .A2(n37099), .ZN(n28649) );
  INV_X1 U108 ( .I(n32304), .ZN(n30187) );
  AND2_X1 U115 ( .A1(n15153), .A2(n9393), .Z(n15605) );
  NOR2_X1 U117 ( .A1(n30232), .A2(n29263), .ZN(n19310) );
  INV_X1 U150 ( .I(n19910), .ZN(n29614) );
  INV_X1 U153 ( .I(n29045), .ZN(n5741) );
  INV_X1 U157 ( .I(n19833), .ZN(n20329) );
  NOR2_X1 U231 ( .A1(n9686), .A2(n14278), .ZN(n450) );
  AOI21_X1 U234 ( .A1(n36814), .A2(n39664), .B(n37460), .ZN(n15110) );
  INV_X2 U268 ( .I(n28689), .ZN(n17771) );
  NAND2_X1 U293 ( .A1(n11283), .A2(n7690), .ZN(n76) );
  INV_X1 U361 ( .I(n27671), .ZN(n14828) );
  INV_X1 U375 ( .I(n30101), .ZN(n1703) );
  INV_X1 U376 ( .I(n19774), .ZN(n29854) );
  INV_X1 U377 ( .I(n19947), .ZN(n17275) );
  INV_X1 U378 ( .I(n29538), .ZN(n1698) );
  INV_X1 U384 ( .I(n29838), .ZN(n1702) );
  INV_X1 U385 ( .I(n19751), .ZN(n21226) );
  INV_X1 U403 ( .I(n19877), .ZN(n27465) );
  NAND2_X1 U419 ( .A1(n27455), .A2(n5101), .ZN(n19030) );
  INV_X1 U449 ( .I(n27108), .ZN(n27230) );
  INV_X1 U459 ( .I(n37075), .ZN(n943) );
  NAND2_X1 U471 ( .A1(n1079), .A2(n995), .ZN(n1797) );
  NOR2_X1 U487 ( .A1(n998), .A2(n27508), .ZN(n27421) );
  INV_X1 U518 ( .I(n26784), .ZN(n3) );
  OAI22_X1 U527 ( .A1(n36873), .A2(n925), .B1(n9147), .B2(n17034), .ZN(n7006)
         );
  NAND3_X1 U533 ( .A1(n2292), .A2(n33858), .A3(n8651), .ZN(n27125) );
  NOR3_X1 U538 ( .A1(n32168), .A2(n13181), .A3(n38483), .ZN(n17573) );
  NAND2_X1 U540 ( .A1(n9654), .A2(n925), .ZN(n81) );
  OAI22_X1 U546 ( .A1(n17823), .A2(n32797), .B1(n26284), .B2(n1229), .ZN(n5221) );
  INV_X1 U552 ( .I(n19615), .ZN(n20021) );
  OR2_X1 U560 ( .A1(n14455), .A2(n26876), .Z(n13184) );
  INV_X1 U629 ( .I(n28968), .ZN(n15046) );
  INV_X1 U633 ( .I(n26587), .ZN(n12383) );
  INV_X1 U641 ( .I(n28910), .ZN(n1730) );
  INV_X1 U642 ( .I(n19952), .ZN(n19799) );
  INV_X1 U643 ( .I(n19887), .ZN(n16498) );
  INV_X1 U644 ( .I(n29671), .ZN(n19432) );
  AOI21_X1 U781 ( .A1(n6300), .A2(n34010), .B(n18837), .ZN(n13533) );
  AOI21_X1 U783 ( .A1(n1535), .A2(n2581), .B(n25466), .ZN(n1933) );
  INV_X1 U794 ( .I(n579), .ZN(n25443) );
  AOI21_X1 U822 ( .A1(n25681), .A2(n7705), .B(n24536), .ZN(n242) );
  NOR3_X1 U827 ( .A1(n18810), .A2(n14436), .A3(n1543), .ZN(n5710) );
  NAND2_X1 U830 ( .A1(n20052), .A2(n31809), .ZN(n25554) );
  NAND2_X1 U852 ( .A1(n36105), .A2(n34427), .ZN(n25519) );
  INV_X1 U892 ( .I(n19729), .ZN(n1733) );
  INV_X1 U893 ( .I(n29319), .ZN(n14969) );
  INV_X1 U900 ( .I(n19851), .ZN(n1719) );
  INV_X1 U903 ( .I(n29707), .ZN(n21280) );
  INV_X1 U904 ( .I(n19885), .ZN(n1735) );
  INV_X1 U905 ( .I(n29801), .ZN(n20781) );
  INV_X1 U906 ( .I(n19913), .ZN(n18993) );
  INV_X1 U912 ( .I(n29298), .ZN(n17646) );
  INV_X1 U913 ( .I(n30207), .ZN(n20804) );
  INV_X1 U922 ( .I(n19649), .ZN(n20748) );
  OR2_X1 U925 ( .A1(n25184), .A2(n7967), .Z(n817) );
  NAND2_X1 U933 ( .A1(n39817), .A2(n18845), .ZN(n24754) );
  NAND2_X1 U938 ( .A1(n35560), .A2(n1580), .ZN(n24490) );
  NAND3_X1 U939 ( .A1(n9921), .A2(n24685), .A3(n24686), .ZN(n7969) );
  INV_X1 U985 ( .I(n24795), .ZN(n7177) );
  NAND2_X1 U1004 ( .A1(n24734), .A2(n5390), .ZN(n5389) );
  INV_X1 U1020 ( .I(n18983), .ZN(n24614) );
  INV_X1 U1041 ( .I(n37227), .ZN(n24275) );
  NOR2_X1 U1052 ( .A1(n14686), .A2(n37994), .ZN(n12) );
  NAND2_X1 U1117 ( .A1(n15892), .A2(n9383), .ZN(n3398) );
  INV_X1 U1143 ( .I(n23846), .ZN(n20594) );
  NAND2_X1 U1168 ( .A1(n1861), .A2(n1632), .ZN(n530) );
  OR2_X1 U1171 ( .A1(n23567), .A2(n1643), .Z(n788) );
  INV_X1 U1181 ( .I(n23484), .ZN(n23364) );
  INV_X1 U1189 ( .I(n38704), .ZN(n98) );
  INV_X1 U1218 ( .I(n7644), .ZN(n16729) );
  NAND2_X1 U1284 ( .A1(n18415), .A2(n22859), .ZN(n5110) );
  INV_X1 U1288 ( .I(n19440), .ZN(n14188) );
  NOR2_X1 U1294 ( .A1(n19698), .A2(n23103), .ZN(n23105) );
  INV_X1 U1304 ( .I(n36453), .ZN(n19769) );
  OAI21_X1 U1309 ( .A1(n22860), .A2(n22861), .B(n22859), .ZN(n4760) );
  NOR2_X1 U1311 ( .A1(n23032), .A2(n22958), .ZN(n22954) );
  INV_X1 U1331 ( .I(n407), .ZN(n8809) );
  INV_X1 U1341 ( .I(n19167), .ZN(n22875) );
  INV_X1 U1351 ( .I(n22879), .ZN(n5892) );
  INV_X1 U1362 ( .I(n11778), .ZN(n22900) );
  BUF_X2 U1369 ( .I(n17628), .Z(n906) );
  NAND2_X1 U1388 ( .A1(n9546), .A2(n64), .ZN(n9521) );
  INV_X1 U1390 ( .I(n6014), .ZN(n1808) );
  NAND2_X1 U1409 ( .A1(n35193), .A2(n4497), .ZN(n367) );
  INV_X2 U1453 ( .I(n16760), .ZN(n22310) );
  AOI21_X1 U1470 ( .A1(n21524), .A2(n21478), .B(n533), .ZN(n532) );
  OR2_X1 U1484 ( .A1(n21688), .A2(n21339), .Z(n5047) );
  NOR2_X1 U1490 ( .A1(n19470), .A2(n13472), .ZN(n3943) );
  INV_X1 U1499 ( .I(n21750), .ZN(n21029) );
  NOR2_X1 U1504 ( .A1(n19545), .A2(n7536), .ZN(n10918) );
  NAND2_X1 U1508 ( .A1(n37200), .A2(n18576), .ZN(n18699) );
  INV_X1 U1529 ( .I(n17964), .ZN(n15338) );
  AND2_X1 U1532 ( .A1(n21722), .A2(n20685), .Z(n12738) );
  INV_X1 U1541 ( .I(n688), .ZN(n1348) );
  INV_X2 U1571 ( .I(n1897), .ZN(n4734) );
  INV_X2 U1572 ( .I(n10004), .ZN(n14635) );
  OAI22_X2 U1587 ( .A1(n6542), .A2(n24576), .B1(n958), .B2(n24723), .ZN(n6541)
         );
  OAI21_X2 U1608 ( .A1(n4636), .A2(n17353), .B(n5355), .ZN(n25567) );
  INV_X2 U1611 ( .I(n28054), .ZN(n6788) );
  INV_X4 U1638 ( .I(n27235), .ZN(n945) );
  AND2_X1 U1640 ( .A1(n27314), .A2(n33417), .Z(n18436) );
  INV_X4 U1646 ( .I(n26839), .ZN(n1092) );
  NAND2_X2 U1682 ( .A1(n10140), .A2(n26107), .ZN(n10139) );
  OAI21_X2 U1722 ( .A1(n5022), .A2(n7431), .B(n27215), .ZN(n28350) );
  INV_X2 U1761 ( .I(n6657), .ZN(n21042) );
  AOI21_X2 U1792 ( .A1(n14541), .A2(n18143), .B(n17866), .ZN(n17865) );
  OAI21_X2 U1827 ( .A1(n22230), .A2(n17156), .B(n36237), .ZN(n17155) );
  INV_X4 U1830 ( .I(n22160), .ZN(n1333) );
  AOI21_X2 U1831 ( .A1(n24599), .A2(n24597), .B(n1563), .ZN(n7443) );
  BUF_X2 U1846 ( .I(n37043), .Z(n4714) );
  INV_X2 U1860 ( .I(n30464), .ZN(n11846) );
  INV_X2 U1871 ( .I(n29574), .ZN(n1393) );
  BUF_X4 U1873 ( .I(n17696), .Z(n603) );
  OAI21_X2 U1876 ( .A1(n26003), .A2(n603), .B(n26005), .ZN(n9667) );
  INV_X4 U1883 ( .I(n17712), .ZN(n1236) );
  NOR2_X2 U1884 ( .A1(n37106), .A2(n259), .ZN(n9217) );
  AOI21_X2 U1912 ( .A1(n15585), .A2(n24695), .B(n38777), .ZN(n12504) );
  NOR2_X1 U1913 ( .A1(n13036), .A2(n17824), .ZN(n207) );
  AOI21_X2 U1922 ( .A1(n21836), .A2(n21837), .B(n14911), .ZN(n14910) );
  INV_X2 U1927 ( .I(n882), .ZN(n1202) );
  AOI21_X2 U1942 ( .A1(n16353), .A2(n20102), .B(n37021), .ZN(n8446) );
  OAI21_X2 U1966 ( .A1(n7972), .A2(n7966), .B(n3655), .ZN(n3654) );
  AOI21_X2 U1967 ( .A1(n25388), .A2(n25389), .B(n25582), .ZN(n4827) );
  INV_X2 U1973 ( .I(n30465), .ZN(n1545) );
  INV_X2 U2044 ( .I(n27253), .ZN(n27115) );
  INV_X2 U2057 ( .I(n20858), .ZN(n17712) );
  OAI21_X2 U2066 ( .A1(n37151), .A2(n26005), .B(n26004), .ZN(n20050) );
  INV_X2 U2079 ( .I(n19223), .ZN(n25677) );
  OAI21_X2 U2093 ( .A1(n39446), .A2(n23095), .B(n8594), .ZN(n14305) );
  OAI21_X2 U2111 ( .A1(n15737), .A2(n35224), .B(n1424), .ZN(n8008) );
  NAND2_X2 U2132 ( .A1(n23391), .A2(n37093), .ZN(n15642) );
  INV_X2 U2152 ( .I(n7364), .ZN(n15385) );
  INV_X4 U2194 ( .I(n13758), .ZN(n1494) );
  NAND2_X1 U2222 ( .A1(n31527), .A2(n17469), .ZN(n4768) );
  NOR2_X1 U2228 ( .A1(n15768), .A2(n37096), .ZN(n29358) );
  NAND2_X2 U2274 ( .A1(n6257), .A2(n17348), .ZN(n17347) );
  NOR3_X1 U2291 ( .A1(n23110), .A2(n20782), .A3(n12392), .ZN(n16132) );
  AND2_X1 U2295 ( .A1(n9725), .A2(n22920), .Z(n22858) );
  INV_X1 U2304 ( .I(n9516), .ZN(n7904) );
  INV_X1 U2307 ( .I(n22571), .ZN(n629) );
  NOR2_X1 U2352 ( .A1(n33966), .A2(n5579), .ZN(n633) );
  INV_X2 U2357 ( .I(n24247), .ZN(n1130) );
  INV_X1 U2393 ( .I(n28940), .ZN(n110) );
  INV_X2 U2403 ( .I(n8519), .ZN(n8518) );
  INV_X1 U2423 ( .I(n28204), .ZN(n1208) );
  NAND2_X1 U2424 ( .A1(n8583), .A2(n29924), .ZN(n8582) );
  OR2_X2 U2426 ( .A1(n13425), .A2(n26177), .Z(n26655) );
  NOR2_X1 U2428 ( .A1(n5089), .A2(n27284), .ZN(n4716) );
  AND2_X2 U2442 ( .A1(n21567), .A2(n3294), .Z(n3821) );
  AOI21_X1 U2455 ( .A1(n11067), .A2(n13981), .B(n37096), .ZN(n13273) );
  OAI21_X2 U2469 ( .A1(n11773), .A2(n14774), .B(n11771), .ZN(n2546) );
  INV_X2 U2483 ( .I(n853), .ZN(n19712) );
  INV_X2 U2504 ( .I(n33966), .ZN(n2347) );
  AND2_X1 U2515 ( .A1(n27910), .A2(n33845), .Z(n15372) );
  XOR2_X1 U2519 ( .A1(n9205), .A2(n22382), .Z(n2781) );
  NAND2_X2 U2522 ( .A1(n2607), .A2(n2610), .ZN(n9701) );
  OAI21_X2 U2544 ( .A1(n37124), .A2(n7590), .B(n21094), .ZN(n10) );
  INV_X2 U2545 ( .I(n11), .ZN(n6163) );
  AOI22_X2 U2559 ( .A1(n22193), .A2(n22194), .B1(n22191), .B2(n22192), .ZN(
        n9982) );
  INV_X2 U2560 ( .I(n25307), .ZN(n18837) );
  NAND3_X1 U2587 ( .A1(n21063), .A2(n21062), .A3(n13352), .ZN(n21061) );
  INV_X2 U2597 ( .I(n22904), .ZN(n4862) );
  OAI21_X2 U2613 ( .A1(n28190), .A2(n28191), .B(n7310), .ZN(n14030) );
  NAND2_X2 U2641 ( .A1(n8053), .A2(n8052), .ZN(n23609) );
  NOR2_X2 U2643 ( .A1(n1821), .A2(n29078), .ZN(n16839) );
  NOR2_X2 U2646 ( .A1(n20112), .A2(n27315), .ZN(n20111) );
  XOR2_X1 U2660 ( .A1(n507), .A2(n30324), .Z(n2446) );
  AOI21_X2 U2688 ( .A1(n37069), .A2(n25512), .B(n36486), .ZN(n46) );
  NAND2_X2 U2727 ( .A1(n13624), .A2(n13636), .ZN(n15332) );
  INV_X2 U2730 ( .I(n63), .ZN(n21285) );
  INV_X1 U2788 ( .I(n9616), .ZN(n19089) );
  OR2_X1 U2802 ( .A1(n24902), .A2(n20158), .Z(n812) );
  INV_X1 U2812 ( .I(n20207), .ZN(n24146) );
  NAND2_X2 U2815 ( .A1(n27967), .A2(n27966), .ZN(n28559) );
  NAND2_X1 U2821 ( .A1(n170), .A2(n4095), .ZN(n29991) );
  NOR3_X2 U2828 ( .A1(n29448), .A2(n19791), .A3(n29447), .ZN(n85) );
  OAI21_X2 U2831 ( .A1(n19579), .A2(n3821), .B(n3295), .ZN(n3327) );
  AOI21_X2 U2869 ( .A1(n5972), .A2(n5973), .B(n5971), .ZN(n5579) );
  XOR2_X1 U2877 ( .A1(n15671), .A2(n2352), .Z(n2351) );
  NAND2_X2 U2893 ( .A1(n12030), .A2(n22161), .ZN(n22162) );
  NAND2_X2 U2897 ( .A1(n2413), .A2(n109), .ZN(n13217) );
  XOR2_X1 U2900 ( .A1(n110), .A2(n5755), .Z(n5889) );
  XOR2_X1 U2918 ( .A1(n22639), .A2(n6329), .Z(n8313) );
  NAND2_X2 U2940 ( .A1(n19963), .A2(n25587), .ZN(n6448) );
  INV_X2 U2941 ( .I(n118), .ZN(n759) );
  XOR2_X1 U2942 ( .A1(n5096), .A2(n12919), .Z(n118) );
  XOR2_X1 U2971 ( .A1(n5031), .A2(n19910), .Z(n11881) );
  XOR2_X1 U2994 ( .A1(n22640), .A2(n22551), .Z(n12102) );
  OAI21_X2 U3023 ( .A1(n6043), .A2(n8800), .B(n1194), .ZN(n137) );
  XOR2_X1 U3044 ( .A1(n15336), .A2(n39073), .Z(n16270) );
  XOR2_X1 U3058 ( .A1(n8015), .A2(n8016), .Z(n16271) );
  XOR2_X1 U3094 ( .A1(n1458), .A2(n27776), .Z(n27675) );
  OR2_X1 U3099 ( .A1(n25772), .A2(n25939), .Z(n155) );
  AOI21_X2 U3105 ( .A1(n2405), .A2(n21924), .B(n8076), .ZN(n2404) );
  INV_X2 U3107 ( .I(n157), .ZN(n8000) );
  XOR2_X1 U3115 ( .A1(n158), .A2(n2592), .Z(n11335) );
  XOR2_X1 U3116 ( .A1(n159), .A2(n31605), .Z(n158) );
  NAND2_X2 U3119 ( .A1(n6263), .A2(n17094), .ZN(n8249) );
  INV_X2 U3140 ( .I(n170), .ZN(n775) );
  XOR2_X1 U3150 ( .A1(n27831), .A2(n20796), .Z(n18663) );
  AOI21_X2 U3152 ( .A1(n20209), .A2(n16074), .B(n14151), .ZN(n14150) );
  NAND2_X2 U3153 ( .A1(n171), .A2(n24498), .ZN(n25266) );
  XOR2_X1 U3163 ( .A1(n22757), .A2(n15753), .Z(n3530) );
  OR2_X1 U3201 ( .A1(n26116), .A2(n30302), .Z(n187) );
  NAND4_X2 U3211 ( .A1(n26426), .A2(n26425), .A3(n26427), .A4(n26674), .ZN(
        n19135) );
  XOR2_X1 U3213 ( .A1(n18512), .A2(n190), .Z(n27671) );
  XOR2_X1 U3214 ( .A1(n18510), .A2(n18511), .Z(n190) );
  XOR2_X1 U3224 ( .A1(n30322), .A2(n12437), .Z(n13235) );
  NOR2_X2 U3225 ( .A1(n11275), .A2(n4619), .ZN(n22465) );
  INV_X2 U3228 ( .I(n37678), .ZN(n21410) );
  NAND3_X2 U3253 ( .A1(n10774), .A2(n17961), .A3(n24757), .ZN(n25197) );
  CLKBUF_X2 U3260 ( .I(Key[63]), .Z(n19953) );
  BUF_X2 U3261 ( .I(Key[74]), .Z(n30150) );
  NAND2_X1 U3266 ( .A1(n16692), .A2(n34073), .ZN(n19013) );
  INV_X2 U3269 ( .I(n25203), .ZN(n3655) );
  AOI21_X1 U3288 ( .A1(n263), .A2(n10152), .B(n1603), .ZN(n7813) );
  AOI21_X2 U3294 ( .A1(n37201), .A2(n20981), .B(n19569), .ZN(n17829) );
  XOR2_X1 U3295 ( .A1(n35463), .A2(n26573), .Z(n5447) );
  NOR2_X2 U3308 ( .A1(n207), .A2(n5221), .ZN(n27385) );
  OR2_X1 U3323 ( .A1(n11375), .A2(n28286), .Z(n6714) );
  NOR2_X2 U3330 ( .A1(n13111), .A2(n13110), .ZN(n26996) );
  INV_X2 U3331 ( .I(n20613), .ZN(n13110) );
  NAND2_X1 U3334 ( .A1(n33703), .A2(n23399), .ZN(n214) );
  NOR2_X1 U3371 ( .A1(n230), .A2(n10050), .ZN(n10190) );
  NOR2_X1 U3372 ( .A1(n3415), .A2(n32209), .ZN(n230) );
  XOR2_X1 U3379 ( .A1(n33736), .A2(n9981), .Z(n13001) );
  INV_X2 U3382 ( .I(n15337), .ZN(n21571) );
  XNOR2_X1 U3390 ( .A1(n23670), .A2(n19890), .ZN(n540) );
  NAND2_X2 U3398 ( .A1(n23826), .A2(n23825), .ZN(n25040) );
  INV_X4 U3399 ( .I(n19718), .ZN(n20376) );
  NAND2_X2 U3401 ( .A1(n2276), .A2(n237), .ZN(n22239) );
  AND2_X1 U3423 ( .A1(n37157), .A2(n19085), .Z(n5825) );
  OAI21_X1 U3425 ( .A1(n18298), .A2(n25681), .B(n242), .ZN(n19503) );
  NOR2_X1 U3443 ( .A1(n251), .A2(n30845), .ZN(n11957) );
  XOR2_X1 U3452 ( .A1(n19472), .A2(n26158), .Z(n254) );
  XOR2_X1 U3457 ( .A1(n15912), .A2(n16498), .Z(n648) );
  XOR2_X1 U3481 ( .A1(n27794), .A2(n1214), .Z(n27497) );
  XOR2_X1 U3498 ( .A1(n266), .A2(n17737), .Z(n29450) );
  OR2_X1 U3503 ( .A1(n13637), .A2(n13638), .Z(n13019) );
  XNOR2_X1 U3514 ( .A1(n16359), .A2(n16358), .ZN(n523) );
  NAND3_X2 U3522 ( .A1(n23818), .A2(n24184), .A3(n39703), .ZN(n13782) );
  XOR2_X1 U3532 ( .A1(n27737), .A2(n20479), .Z(n27483) );
  OAI21_X2 U3545 ( .A1(n27391), .A2(n14881), .B(n37246), .ZN(n26869) );
  OAI22_X1 U3552 ( .A1(n11939), .A2(n15601), .B1(n280), .B2(n3462), .ZN(n5811)
         );
  OAI21_X2 U3555 ( .A1(n24700), .A2(n6791), .B(n6490), .ZN(n8388) );
  XOR2_X1 U3568 ( .A1(n22703), .A2(n4493), .Z(n22571) );
  NAND2_X2 U3570 ( .A1(n15787), .A2(n23560), .ZN(n23340) );
  AOI22_X2 U3574 ( .A1(n11517), .A2(n14377), .B1(n26759), .B2(n6891), .ZN(
        n11516) );
  XOR2_X1 U3581 ( .A1(n17342), .A2(n1162), .Z(n5692) );
  INV_X2 U3590 ( .I(n18829), .ZN(n30109) );
  NAND2_X2 U3606 ( .A1(n6898), .A2(n13252), .ZN(n5218) );
  INV_X1 U3613 ( .I(n26818), .ZN(n26990) );
  BUF_X2 U3648 ( .I(n12961), .Z(n301) );
  XOR2_X1 U3653 ( .A1(n476), .A2(n36065), .Z(n23793) );
  BUF_X2 U3660 ( .I(n28673), .Z(n306) );
  XOR2_X1 U3661 ( .A1(n35654), .A2(n26532), .Z(n6879) );
  NAND2_X1 U3663 ( .A1(n12150), .A2(n12547), .ZN(n307) );
  INV_X2 U3666 ( .I(n26919), .ZN(n3606) );
  INV_X4 U3674 ( .I(n14379), .ZN(n24390) );
  XOR2_X1 U3715 ( .A1(n320), .A2(n9563), .Z(n15159) );
  NAND2_X2 U3747 ( .A1(n24646), .A2(n36321), .ZN(n24599) );
  XOR2_X1 U3758 ( .A1(n23723), .A2(n9153), .Z(n6516) );
  XOR2_X1 U3762 ( .A1(n331), .A2(n9003), .Z(n14290) );
  OR2_X1 U3776 ( .A1(n31518), .A2(n27424), .Z(n336) );
  XOR2_X1 U3807 ( .A1(n7022), .A2(n342), .Z(n19888) );
  AND2_X1 U3813 ( .A1(n21023), .A2(n344), .Z(n8761) );
  NAND2_X2 U3816 ( .A1(n346), .A2(n24485), .ZN(n24874) );
  AOI21_X2 U3826 ( .A1(n37165), .A2(n11243), .B(n11241), .ZN(n26124) );
  NOR2_X2 U3838 ( .A1(n5098), .A2(n4516), .ZN(n4515) );
  XOR2_X1 U3853 ( .A1(n353), .A2(n6223), .Z(n5656) );
  XOR2_X1 U3856 ( .A1(n6033), .A2(n19355), .Z(n27194) );
  OAI21_X2 U3857 ( .A1(n37), .A2(n7872), .B(n28215), .ZN(n3928) );
  NAND2_X2 U3880 ( .A1(n21231), .A2(n24735), .ZN(n24620) );
  XOR2_X1 U3882 ( .A1(n2615), .A2(n6436), .Z(n13207) );
  AOI22_X2 U3884 ( .A1(n9461), .A2(n37837), .B1(n15298), .B2(n36819), .ZN(
        n26163) );
  INV_X2 U3945 ( .I(n27798), .ZN(n379) );
  NAND2_X2 U3958 ( .A1(n1289), .A2(n1596), .ZN(n23983) );
  INV_X2 U3961 ( .I(n29923), .ZN(n29924) );
  INV_X4 U3966 ( .I(n11120), .ZN(n12543) );
  AOI21_X2 U3974 ( .A1(n21362), .A2(n21361), .B(n21360), .ZN(n19718) );
  NOR2_X2 U3981 ( .A1(n21847), .A2(n21672), .ZN(n20469) );
  INV_X2 U3985 ( .I(n23083), .ZN(n23188) );
  XOR2_X1 U3991 ( .A1(n387), .A2(n18416), .Z(n9176) );
  XOR2_X1 U4002 ( .A1(n15656), .A2(n15660), .Z(n391) );
  NAND3_X2 U4010 ( .A1(n25707), .A2(n25706), .A3(n25705), .ZN(n26602) );
  OR2_X1 U4011 ( .A1(n20776), .A2(n32471), .Z(n12642) );
  NAND2_X2 U4012 ( .A1(n24353), .A2(n24477), .ZN(n1898) );
  NAND2_X1 U4023 ( .A1(n36552), .A2(n8193), .ZN(n4761) );
  INV_X2 U4025 ( .I(n9942), .ZN(n21902) );
  BUF_X2 U4029 ( .I(n7757), .Z(n6445) );
  INV_X4 U4033 ( .I(n17307), .ZN(n22265) );
  NAND2_X2 U4039 ( .A1(n13986), .A2(n2792), .ZN(n13606) );
  OAI21_X1 U4041 ( .A1(n20474), .A2(n29704), .B(n29581), .ZN(n20473) );
  OAI21_X1 U4044 ( .A1(n28699), .A2(n16295), .B(n28696), .ZN(n10303) );
  XOR2_X1 U4052 ( .A1(n2317), .A2(n16133), .Z(n10026) );
  BUF_X2 U4054 ( .I(Key[109]), .Z(n19825) );
  XOR2_X1 U4060 ( .A1(n27724), .A2(n27640), .Z(n27798) );
  INV_X2 U4070 ( .I(n22665), .ZN(n1324) );
  NAND2_X2 U4079 ( .A1(n13293), .A2(n13292), .ZN(n13289) );
  NOR2_X2 U4093 ( .A1(n21416), .A2(n21415), .ZN(n21982) );
  XOR2_X1 U4100 ( .A1(n412), .A2(n851), .Z(n3486) );
  XOR2_X1 U4106 ( .A1(n416), .A2(n17642), .Z(n20702) );
  XOR2_X1 U4107 ( .A1(n29148), .A2(n14221), .Z(n416) );
  NAND2_X1 U4123 ( .A1(n16158), .A2(n34783), .ZN(n422) );
  AND2_X1 U4127 ( .A1(n7536), .A2(n21410), .Z(n10915) );
  XOR2_X1 U4138 ( .A1(n2473), .A2(n427), .Z(n3027) );
  XOR2_X1 U4139 ( .A1(n2471), .A2(n22654), .Z(n427) );
  XOR2_X1 U4147 ( .A1(n431), .A2(n33965), .Z(n15854) );
  AOI21_X1 U4156 ( .A1(n29918), .A2(n29919), .B(n434), .ZN(n16992) );
  INV_X1 U4194 ( .I(n10144), .ZN(n440) );
  XOR2_X1 U4197 ( .A1(n29085), .A2(n28826), .Z(n4141) );
  XOR2_X1 U4213 ( .A1(n16523), .A2(n5370), .Z(n3709) );
  INV_X2 U4220 ( .I(n18959), .ZN(n21730) );
  AOI21_X2 U4225 ( .A1(n16578), .A2(n12793), .B(n5147), .ZN(n5146) );
  AOI22_X1 U4230 ( .A1(n9907), .A2(n13108), .B1(n13106), .B2(n29222), .ZN(
        n13105) );
  NAND2_X2 U4235 ( .A1(n3867), .A2(n3864), .ZN(n3863) );
  NAND2_X2 U4239 ( .A1(n22300), .A2(n35431), .ZN(n9941) );
  OAI21_X2 U4254 ( .A1(n9723), .A2(n9722), .B(n1608), .ZN(n13073) );
  XOR2_X1 U4278 ( .A1(n17756), .A2(n29974), .Z(n3478) );
  AOI21_X2 U4280 ( .A1(n30364), .A2(n8757), .B(n462), .ZN(n7150) );
  XOR2_X1 U4289 ( .A1(n14986), .A2(n27533), .Z(n18060) );
  INV_X1 U4294 ( .I(n1740), .ZN(n29163) );
  INV_X2 U4306 ( .I(n26729), .ZN(n8814) );
  NOR2_X1 U4320 ( .A1(n37160), .A2(n25630), .ZN(n17855) );
  INV_X2 U4328 ( .I(n474), .ZN(n12365) );
  NAND2_X2 U4334 ( .A1(n2341), .A2(n17101), .ZN(n15136) );
  NAND3_X2 U4343 ( .A1(n4660), .A2(n15966), .A3(n5552), .ZN(n4875) );
  INV_X4 U4351 ( .I(n19594), .ZN(n1316) );
  XOR2_X1 U4363 ( .A1(n485), .A2(n6802), .Z(n6801) );
  XOR2_X1 U4364 ( .A1(n4796), .A2(n11688), .Z(n485) );
  INV_X2 U4371 ( .I(n8454), .ZN(n12081) );
  NAND3_X2 U4376 ( .A1(n22095), .A2(n22097), .A3(n22096), .ZN(n22648) );
  INV_X4 U4385 ( .I(n22337), .ZN(n22100) );
  INV_X2 U4389 ( .I(n22092), .ZN(n22356) );
  XOR2_X1 U4397 ( .A1(n31127), .A2(n29131), .Z(n489) );
  OR2_X1 U4404 ( .A1(n2257), .A2(n22019), .Z(n2709) );
  NOR2_X2 U4412 ( .A1(n19609), .A2(n19641), .ZN(n21433) );
  XOR2_X1 U4413 ( .A1(n2997), .A2(n27493), .Z(n8425) );
  INV_X4 U4441 ( .I(n18144), .ZN(n1200) );
  INV_X4 U4445 ( .I(n20476), .ZN(n1354) );
  NAND2_X2 U4456 ( .A1(n8971), .A2(n10044), .ZN(n18059) );
  AOI21_X2 U4457 ( .A1(n18059), .A2(n21371), .B(n9253), .ZN(n9251) );
  NAND2_X2 U4477 ( .A1(n16642), .A2(n16643), .ZN(n19847) );
  XOR2_X1 U4482 ( .A1(n10653), .A2(n10622), .Z(n6212) );
  XOR2_X1 U4487 ( .A1(n18597), .A2(n509), .Z(n784) );
  XOR2_X1 U4492 ( .A1(n26482), .A2(n9398), .Z(n3459) );
  INV_X1 U4494 ( .I(n26483), .ZN(n2711) );
  XOR2_X1 U4511 ( .A1(n514), .A2(n22057), .Z(n9420) );
  NAND2_X2 U4519 ( .A1(n25830), .A2(n1512), .ZN(n25919) );
  OAI21_X1 U4521 ( .A1(n11718), .A2(n902), .B(n515), .ZN(n11719) );
  AND2_X1 U4525 ( .A1(n10171), .A2(n2722), .Z(n12213) );
  XOR2_X1 U4528 ( .A1(n11355), .A2(n33936), .Z(n11354) );
  OR3_X1 U4540 ( .A1(n15354), .A2(n114), .A3(n1816), .Z(n1766) );
  INV_X2 U4553 ( .I(n3526), .ZN(n20405) );
  INV_X4 U4558 ( .I(n4553), .ZN(n25978) );
  XOR2_X1 U4570 ( .A1(n28999), .A2(n28998), .Z(n18452) );
  XOR2_X1 U4574 ( .A1(n525), .A2(n30479), .Z(n1455) );
  XOR2_X1 U4575 ( .A1(n16218), .A2(n11996), .Z(n525) );
  INV_X2 U4583 ( .I(n11643), .ZN(n19293) );
  NAND2_X2 U4592 ( .A1(n34404), .A2(n9524), .ZN(n9523) );
  INV_X2 U4609 ( .I(n855), .ZN(n17515) );
  AOI22_X2 U4618 ( .A1(n9705), .A2(n18112), .B1(n9886), .B2(n39650), .ZN(n7759) );
  INV_X2 U4623 ( .I(n19978), .ZN(n25623) );
  AOI21_X2 U4638 ( .A1(n538), .A2(n21764), .B(n15148), .ZN(n15614) );
  AOI21_X2 U4640 ( .A1(n14899), .A2(n33580), .B(n14898), .ZN(n14897) );
  XOR2_X1 U4644 ( .A1(n540), .A2(n23684), .Z(n16893) );
  XOR2_X1 U4653 ( .A1(n10200), .A2(n1867), .Z(n12410) );
  NAND2_X2 U4660 ( .A1(n4597), .A2(n11434), .ZN(n5044) );
  XOR2_X1 U4677 ( .A1(n7944), .A2(n7148), .Z(n19112) );
  NAND2_X2 U4678 ( .A1(n7144), .A2(n7145), .ZN(n7148) );
  AOI22_X2 U4684 ( .A1(n919), .A2(n21833), .B1(n21834), .B2(n19620), .ZN(
        n15951) );
  NOR2_X1 U4686 ( .A1(n19349), .A2(n7905), .ZN(n551) );
  AOI21_X2 U4695 ( .A1(n18104), .A2(n38215), .B(n29956), .ZN(n19093) );
  INV_X2 U4713 ( .I(n39823), .ZN(n11707) );
  NOR2_X2 U4717 ( .A1(n13964), .A2(n13963), .ZN(n13962) );
  XOR2_X1 U4729 ( .A1(n562), .A2(n18301), .Z(n16905) );
  OAI21_X2 U4746 ( .A1(n24147), .A2(n5360), .B(n5359), .ZN(n24794) );
  INV_X2 U4780 ( .I(n21792), .ZN(n21660) );
  INV_X2 U4786 ( .I(n21432), .ZN(n21822) );
  XOR2_X1 U4810 ( .A1(n588), .A2(n29983), .Z(Ciphertext[137]) );
  OAI22_X1 U4811 ( .A1(n29982), .A2(n29981), .B1(n18200), .B2(n5678), .ZN(n588) );
  AND2_X1 U4812 ( .A1(n17867), .A2(n7883), .Z(n2058) );
  AOI21_X2 U4828 ( .A1(n13409), .A2(n10536), .B(n19969), .ZN(n28656) );
  NAND2_X2 U4835 ( .A1(n5479), .A2(n5477), .ZN(n12685) );
  NAND2_X2 U4838 ( .A1(n13669), .A2(n13671), .ZN(n13442) );
  INV_X2 U4850 ( .I(n38210), .ZN(n25472) );
  NOR2_X1 U4859 ( .A1(n35604), .A2(n15245), .ZN(n15243) );
  INV_X2 U4870 ( .I(n9626), .ZN(n22652) );
  NOR2_X2 U4880 ( .A1(n9050), .A2(n23032), .ZN(n22956) );
  XOR2_X1 U4882 ( .A1(n17277), .A2(n18434), .Z(n7327) );
  NAND2_X2 U4883 ( .A1(n28272), .A2(n13609), .ZN(n12644) );
  INV_X2 U4884 ( .I(n12644), .ZN(n20663) );
  XOR2_X1 U4888 ( .A1(n25124), .A2(n25125), .Z(n606) );
  XOR2_X1 U4890 ( .A1(n608), .A2(n16861), .Z(n27538) );
  XOR2_X1 U4916 ( .A1(n6635), .A2(n2979), .Z(n2215) );
  INV_X2 U4930 ( .I(n615), .ZN(n10896) );
  XOR2_X1 U4931 ( .A1(n10899), .A2(n10897), .Z(n615) );
  AOI21_X1 U4934 ( .A1(n29480), .A2(n29466), .B(n616), .ZN(n29467) );
  AOI21_X1 U4938 ( .A1(n619), .A2(n29753), .B(n30555), .ZN(n29725) );
  NAND2_X1 U4939 ( .A1(n38143), .A2(n29740), .ZN(n619) );
  NAND2_X2 U4941 ( .A1(n27386), .A2(n7680), .ZN(n27492) );
  NAND2_X2 U4942 ( .A1(n21057), .A2(n21060), .ZN(n21961) );
  XOR2_X1 U4943 ( .A1(n23882), .A2(n23724), .Z(n5412) );
  NOR2_X1 U4947 ( .A1(n6202), .A2(n1183), .ZN(n6201) );
  NOR2_X1 U4965 ( .A1(n4613), .A2(n20391), .ZN(n15719) );
  BUF_X4 U4973 ( .I(n4381), .Z(n2625) );
  AOI21_X2 U4978 ( .A1(n14118), .A2(n28129), .B(n14117), .ZN(n13690) );
  NAND2_X2 U4980 ( .A1(n4978), .A2(n4977), .ZN(n28207) );
  INV_X4 U4983 ( .I(n38204), .ZN(n11700) );
  XOR2_X1 U4985 ( .A1(n3203), .A2(n629), .Z(n628) );
  INV_X4 U4987 ( .I(n13285), .ZN(n1351) );
  XOR2_X1 U4995 ( .A1(n18305), .A2(n13639), .Z(n632) );
  XOR2_X1 U4999 ( .A1(n2943), .A2(n8940), .Z(n29148) );
  XOR2_X1 U5001 ( .A1(n14977), .A2(n5873), .Z(n635) );
  XOR2_X1 U5003 ( .A1(n636), .A2(n18976), .Z(n18269) );
  INV_X1 U5005 ( .I(n36735), .ZN(n8970) );
  NOR3_X1 U5011 ( .A1(n21693), .A2(n21410), .A3(n36735), .ZN(n9040) );
  NAND2_X1 U5012 ( .A1(n21814), .A2(n21352), .ZN(n21431) );
  AOI21_X1 U5013 ( .A1(n10822), .A2(n36735), .B(n21693), .ZN(n10821) );
  INV_X1 U5017 ( .I(n8026), .ZN(n22590) );
  INV_X1 U5044 ( .I(n19775), .ZN(n26330) );
  INV_X1 U5049 ( .I(n19929), .ZN(n1727) );
  INV_X1 U5056 ( .I(n11562), .ZN(n923) );
  NOR3_X1 U5062 ( .A1(n36344), .A2(n19728), .A3(n38591), .ZN(n27123) );
  INV_X1 U5065 ( .I(n19903), .ZN(n1704) );
  NAND2_X1 U5066 ( .A1(n27421), .A2(n30768), .ZN(n27509) );
  INV_X1 U5067 ( .I(n19845), .ZN(n19020) );
  INV_X1 U5079 ( .I(n29875), .ZN(n28868) );
  INV_X1 U5086 ( .I(n19875), .ZN(n29109) );
  INV_X1 U5088 ( .I(n29432), .ZN(n15181) );
  INV_X1 U5090 ( .I(n29003), .ZN(n1365) );
  INV_X1 U5091 ( .I(n19817), .ZN(n29730) );
  INV_X1 U5092 ( .I(n19905), .ZN(n15273) );
  INV_X1 U5094 ( .I(n19904), .ZN(n15700) );
  INV_X1 U5095 ( .I(n19755), .ZN(n1738) );
  AND2_X1 U5096 ( .A1(n22188), .A2(n39607), .Z(n637) );
  XNOR2_X1 U5097 ( .A1(n23680), .A2(n30006), .ZN(n638) );
  XNOR2_X1 U5098 ( .A1(n22613), .A2(n15762), .ZN(n639) );
  XNOR2_X1 U5105 ( .A1(n29680), .A2(n1010), .ZN(n646) );
  XNOR2_X1 U5108 ( .A1(n4302), .A2(n27739), .ZN(n650) );
  XNOR2_X1 U5111 ( .A1(n35610), .A2(n21280), .ZN(n654) );
  XNOR2_X1 U5112 ( .A1(n18300), .A2(n17428), .ZN(n655) );
  XNOR2_X1 U5113 ( .A1(n17605), .A2(n37110), .ZN(n656) );
  XNOR2_X1 U5114 ( .A1(n25271), .A2(n19937), .ZN(n657) );
  XNOR2_X1 U5115 ( .A1(n22510), .A2(n20206), .ZN(n658) );
  XNOR2_X1 U5118 ( .A1(n24065), .A2(n29671), .ZN(n661) );
  XNOR2_X1 U5119 ( .A1(n16492), .A2(n28831), .ZN(n662) );
  XNOR2_X1 U5120 ( .A1(n30612), .A2(n31771), .ZN(n663) );
  XNOR2_X1 U5121 ( .A1(n25175), .A2(n19950), .ZN(n664) );
  XNOR2_X1 U5122 ( .A1(n35262), .A2(n29229), .ZN(n665) );
  XNOR2_X1 U5124 ( .A1(n23874), .A2(n23591), .ZN(n666) );
  XNOR2_X1 U5126 ( .A1(n36867), .A2(n22763), .ZN(n669) );
  XNOR2_X1 U5129 ( .A1(n24050), .A2(n19758), .ZN(n672) );
  XNOR2_X1 U5130 ( .A1(n27595), .A2(n19676), .ZN(n673) );
  XNOR2_X1 U5131 ( .A1(n34902), .A2(n15046), .ZN(n674) );
  XNOR2_X1 U5132 ( .A1(n23884), .A2(n29964), .ZN(n675) );
  XNOR2_X1 U5134 ( .A1(n27799), .A2(n1161), .ZN(n677) );
  XNOR2_X1 U5135 ( .A1(n23894), .A2(n1367), .ZN(n678) );
  XNOR2_X1 U5137 ( .A1(n29041), .A2(n19913), .ZN(n680) );
  XNOR2_X1 U5138 ( .A1(n29095), .A2(n1377), .ZN(n681) );
  XNOR2_X1 U5139 ( .A1(n27617), .A2(n30114), .ZN(n682) );
  XOR2_X1 U5142 ( .A1(Plaintext[10]), .A2(Key[10]), .Z(n686) );
  INV_X2 U5144 ( .I(n22219), .ZN(n1688) );
  XOR2_X1 U5145 ( .A1(Plaintext[22]), .A2(Key[22]), .Z(n688) );
  XNOR2_X1 U5148 ( .A1(Plaintext[30]), .A2(Key[30]), .ZN(n690) );
  XOR2_X1 U5151 ( .A1(Plaintext[114]), .A2(Key[114]), .Z(n694) );
  INV_X1 U5152 ( .I(n21805), .ZN(n21693) );
  XNOR2_X1 U5153 ( .A1(n22651), .A2(n22430), .ZN(n696) );
  XNOR2_X1 U5154 ( .A1(n22463), .A2(n16648), .ZN(n697) );
  XNOR2_X1 U5155 ( .A1(n4493), .A2(n19648), .ZN(n698) );
  XNOR2_X1 U5156 ( .A1(n22474), .A2(n32993), .ZN(n699) );
  XNOR2_X1 U5157 ( .A1(n32135), .A2(n19885), .ZN(n700) );
  XNOR2_X1 U5158 ( .A1(n10268), .A2(n10267), .ZN(n701) );
  XNOR2_X1 U5160 ( .A1(n20392), .A2(n29363), .ZN(n704) );
  XNOR2_X1 U5161 ( .A1(n22731), .A2(n19254), .ZN(n705) );
  XNOR2_X1 U5162 ( .A1(n22775), .A2(n29689), .ZN(n706) );
  AND2_X1 U5163 ( .A1(n21461), .A2(n21870), .Z(n707) );
  XOR2_X1 U5164 ( .A1(n17285), .A2(n17283), .Z(n708) );
  XNOR2_X1 U5166 ( .A1(n5185), .A2(n29320), .ZN(n710) );
  XNOR2_X1 U5167 ( .A1(n14322), .A2(n9496), .ZN(n711) );
  XNOR2_X1 U5170 ( .A1(n33672), .A2(n30253), .ZN(n713) );
  XNOR2_X1 U5171 ( .A1(n19932), .A2(n37957), .ZN(n714) );
  XNOR2_X1 U5176 ( .A1(n2145), .A2(n23658), .ZN(n718) );
  XNOR2_X1 U5177 ( .A1(n14385), .A2(n19876), .ZN(n719) );
  XNOR2_X1 U5178 ( .A1(n36218), .A2(n29411), .ZN(n720) );
  XNOR2_X1 U5179 ( .A1(n25301), .A2(n16618), .ZN(n721) );
  XNOR2_X1 U5181 ( .A1(n24932), .A2(n25160), .ZN(n723) );
  XNOR2_X1 U5182 ( .A1(n25216), .A2(n25123), .ZN(n724) );
  XNOR2_X1 U5185 ( .A1(n9701), .A2(n25296), .ZN(n727) );
  XNOR2_X1 U5187 ( .A1(n25030), .A2(n28934), .ZN(n729) );
  XNOR2_X1 U5189 ( .A1(n25241), .A2(n29649), .ZN(n731) );
  XNOR2_X1 U5194 ( .A1(n10012), .A2(n1733), .ZN(n736) );
  XNOR2_X1 U5195 ( .A1(n26262), .A2(n19761), .ZN(n737) );
  XNOR2_X1 U5196 ( .A1(n26455), .A2(n19677), .ZN(n738) );
  XNOR2_X1 U5197 ( .A1(n26340), .A2(n26357), .ZN(n739) );
  XNOR2_X1 U5199 ( .A1(n24933), .A2(n25177), .ZN(n741) );
  XNOR2_X1 U5200 ( .A1(n23970), .A2(n23697), .ZN(n742) );
  XNOR2_X1 U5201 ( .A1(n9246), .A2(n965), .ZN(n743) );
  XNOR2_X1 U5203 ( .A1(n5084), .A2(n29223), .ZN(n745) );
  XNOR2_X1 U5205 ( .A1(n26255), .A2(n1050), .ZN(n747) );
  XNOR2_X1 U5206 ( .A1(n6989), .A2(n29514), .ZN(n748) );
  XNOR2_X1 U5207 ( .A1(n6989), .A2(n29831), .ZN(n749) );
  XNOR2_X1 U5208 ( .A1(n26587), .A2(n19805), .ZN(n750) );
  INV_X1 U5211 ( .I(n19226), .ZN(n26895) );
  XNOR2_X1 U5215 ( .A1(n27664), .A2(n19936), .ZN(n756) );
  XNOR2_X1 U5219 ( .A1(n35188), .A2(n30090), .ZN(n760) );
  XNOR2_X1 U5220 ( .A1(n31620), .A2(n35140), .ZN(n761) );
  XNOR2_X1 U5221 ( .A1(n27528), .A2(n19355), .ZN(n763) );
  XNOR2_X1 U5222 ( .A1(n28966), .A2(n30150), .ZN(n764) );
  XNOR2_X1 U5223 ( .A1(n28940), .A2(n1369), .ZN(n765) );
  XNOR2_X1 U5226 ( .A1(n13852), .A2(n19786), .ZN(n769) );
  XNOR2_X1 U5227 ( .A1(n10343), .A2(n29067), .ZN(n770) );
  XNOR2_X1 U5229 ( .A1(n31535), .A2(n19887), .ZN(n772) );
  XNOR2_X1 U5230 ( .A1(n35832), .A2(n1733), .ZN(n774) );
  XNOR2_X1 U5233 ( .A1(n6311), .A2(n22469), .ZN(n778) );
  XOR2_X1 U5238 ( .A1(n6610), .A2(n6608), .Z(n782) );
  XNOR2_X1 U5253 ( .A1(n23623), .A2(n29974), .ZN(n790) );
  XNOR2_X1 U5257 ( .A1(n23927), .A2(n20594), .ZN(n794) );
  XOR2_X1 U5267 ( .A1(n15730), .A2(n15728), .Z(n801) );
  BUF_X2 U5269 ( .I(n24285), .Z(n13970) );
  INV_X2 U5271 ( .I(n24307), .ZN(n14371) );
  NAND2_X2 U5282 ( .A1(n24300), .A2(n39815), .ZN(n14206) );
  AND2_X1 U5283 ( .A1(n24191), .A2(n18466), .Z(n808) );
  XNOR2_X1 U5291 ( .A1(n25241), .A2(n19677), .ZN(n810) );
  XOR2_X1 U5295 ( .A1(n39765), .A2(n30122), .Z(n814) );
  NAND2_X2 U5301 ( .A1(n12914), .A2(n4840), .ZN(n6759) );
  XNOR2_X1 U5305 ( .A1(n824), .A2(n741), .ZN(n823) );
  XOR2_X1 U5307 ( .A1(n4551), .A2(n4550), .Z(n825) );
  XOR2_X1 U5313 ( .A1(n3187), .A2(n3188), .Z(n830) );
  AND2_X2 U5320 ( .A1(n25714), .A2(n25713), .Z(n834) );
  XOR2_X1 U5326 ( .A1(n19384), .A2(n29282), .Z(n837) );
  XNOR2_X1 U5334 ( .A1(n26359), .A2(n30068), .ZN(n838) );
  XNOR2_X1 U5335 ( .A1(n25595), .A2(n25594), .ZN(n839) );
  XNOR2_X1 U5342 ( .A1(n26191), .A2(n26192), .ZN(n845) );
  XNOR2_X1 U5345 ( .A1(n26488), .A2(n8950), .ZN(n848) );
  XNOR2_X1 U5354 ( .A1(n14770), .A2(n14771), .ZN(n856) );
  XNOR2_X1 U5359 ( .A1(n9300), .A2(n9297), .ZN(n859) );
  AND2_X1 U5364 ( .A1(n26934), .A2(n17993), .Z(n863) );
  XOR2_X1 U5371 ( .A1(n26410), .A2(n3858), .Z(n866) );
  INV_X1 U5373 ( .I(n867), .ZN(n9690) );
  XNOR2_X1 U5385 ( .A1(n35189), .A2(n27823), .ZN(n869) );
  XNOR2_X1 U5386 ( .A1(n27491), .A2(n900), .ZN(n870) );
  XNOR2_X1 U5389 ( .A1(n27513), .A2(n27514), .ZN(n873) );
  XNOR2_X1 U5396 ( .A1(n20140), .A2(n19421), .ZN(n877) );
  INV_X1 U5399 ( .I(n20531), .ZN(n28222) );
  XNOR2_X1 U5408 ( .A1(n9139), .A2(n7764), .ZN(n886) );
  BUF_X2 U5421 ( .I(n28883), .Z(n29486) );
  BUF_X2 U5422 ( .I(n30243), .Z(n6443) );
  XNOR2_X1 U5425 ( .A1(n28574), .A2(n28493), .ZN(n893) );
  AOI21_X2 U5430 ( .A1(n16144), .A2(n7612), .B(n14764), .ZN(n3923) );
  OAI21_X2 U5434 ( .A1(n9319), .A2(n9318), .B(n9317), .ZN(n22219) );
  NAND2_X1 U5443 ( .A1(n5402), .A2(n6285), .ZN(n28017) );
  OAI21_X2 U5446 ( .A1(n4375), .A2(n28215), .B(n3928), .ZN(n28326) );
  AOI21_X2 U5456 ( .A1(n1319), .A2(n1654), .B(n5437), .ZN(n22851) );
  NAND2_X1 U5460 ( .A1(n918), .A2(n21478), .ZN(n14527) );
  NAND2_X1 U5461 ( .A1(n20266), .A2(n21478), .ZN(n2278) );
  NAND2_X1 U5462 ( .A1(n21478), .A2(n37200), .ZN(n1814) );
  OAI21_X2 U5469 ( .A1(n22927), .A2(n8141), .B(n37087), .ZN(n23611) );
  INV_X2 U5505 ( .I(n16382), .ZN(n26780) );
  NOR2_X1 U5507 ( .A1(n23057), .A2(n3310), .ZN(n8142) );
  NAND2_X1 U5508 ( .A1(n18450), .A2(n11576), .ZN(n21450) );
  OAI21_X2 U5509 ( .A1(n2237), .A2(n2236), .B(n2233), .ZN(n2082) );
  BUF_X4 U5519 ( .I(n22813), .Z(n23078) );
  AOI22_X2 U5537 ( .A1(n3268), .A2(n22301), .B1(n22039), .B2(n22299), .ZN(
        n3267) );
  OAI22_X2 U5549 ( .A1(n7911), .A2(n9546), .B1(n3181), .B2(n22147), .ZN(n1965)
         );
  NOR2_X1 U5557 ( .A1(n7240), .A2(n1921), .ZN(n8359) );
  OAI21_X1 U5565 ( .A1(n9231), .A2(n30038), .B(n30009), .ZN(n5369) );
  NOR3_X1 U5577 ( .A1(n12081), .A2(n30187), .A3(n30240), .ZN(n6864) );
  BUF_X4 U5600 ( .I(n27908), .Z(n28755) );
  INV_X4 U5609 ( .I(n876), .ZN(n18392) );
  NAND3_X1 U5612 ( .A1(n28054), .A2(n34008), .A3(n1072), .ZN(n13697) );
  INV_X1 U5618 ( .I(n33958), .ZN(n18451) );
  NAND3_X1 U5640 ( .A1(n26976), .A2(n12065), .A3(n10902), .ZN(n26977) );
  INV_X1 U5653 ( .I(n924), .ZN(n13801) );
  INV_X1 U5665 ( .I(n26165), .ZN(n1096) );
  NAND3_X1 U5669 ( .A1(n37683), .A2(n25992), .A3(n1012), .ZN(n8161) );
  INV_X2 U5670 ( .I(n33440), .ZN(n1101) );
  INV_X2 U5672 ( .I(n7901), .ZN(n14375) );
  INV_X4 U5684 ( .I(n11060), .ZN(n17353) );
  NOR2_X1 U5699 ( .A1(n24500), .A2(n933), .ZN(n12207) );
  INV_X2 U5725 ( .I(n10659), .ZN(n19682) );
  OAI21_X2 U5749 ( .A1(n22959), .A2(n22960), .B(n7639), .ZN(n5357) );
  NOR2_X1 U5755 ( .A1(n7960), .A2(n8151), .ZN(n23057) );
  INV_X2 U5766 ( .I(n18433), .ZN(n23053) );
  NOR3_X1 U5779 ( .A1(n22038), .A2(n8899), .A3(n21802), .ZN(n5698) );
  NAND2_X2 U5804 ( .A1(n16014), .A2(n16015), .ZN(n22122) );
  BUF_X2 U5817 ( .I(n33506), .Z(n19470) );
  NOR3_X1 U5839 ( .A1(n971), .A2(n16510), .A3(n21285), .ZN(n9048) );
  NAND3_X1 U5841 ( .A1(n3986), .A2(n4095), .A3(n1058), .ZN(n11217) );
  INV_X1 U5852 ( .I(n9930), .ZN(n12765) );
  NAND2_X2 U5858 ( .A1(n28350), .A2(n28351), .ZN(n28496) );
  NOR2_X1 U5874 ( .A1(n1473), .A2(n35500), .ZN(n4254) );
  INV_X1 U5906 ( .I(n17097), .ZN(n26686) );
  INV_X2 U5910 ( .I(n18390), .ZN(n26688) );
  INV_X2 U5913 ( .I(n14121), .ZN(n924) );
  INV_X1 U5939 ( .I(n252), .ZN(n14460) );
  OAI22_X1 U5950 ( .A1(n24603), .A2(n1270), .B1(n32391), .B2(n5282), .ZN(
        n20807) );
  NAND2_X2 U5961 ( .A1(n10777), .A2(n10784), .ZN(n20039) );
  INV_X4 U5962 ( .I(n13779), .ZN(n933) );
  AND2_X1 U5963 ( .A1(n1597), .A2(n1586), .Z(n10069) );
  NOR2_X1 U5966 ( .A1(n7364), .A2(n5986), .ZN(n24335) );
  INV_X1 U5981 ( .I(n23582), .ZN(n14855) );
  NAND2_X1 U5988 ( .A1(n7584), .A2(n37815), .ZN(n7071) );
  NAND3_X1 U6007 ( .A1(n11091), .A2(n39075), .A3(n5497), .ZN(n5496) );
  NAND2_X1 U6009 ( .A1(n22325), .A2(n12365), .ZN(n17781) );
  NAND3_X1 U6011 ( .A1(n37113), .A2(n18253), .A3(n17976), .ZN(n1864) );
  INV_X1 U6012 ( .I(n9485), .ZN(n9483) );
  NOR2_X1 U6018 ( .A1(n17440), .A2(n22047), .ZN(n22111) );
  INV_X1 U6026 ( .I(n19017), .ZN(n22496) );
  NAND3_X1 U6031 ( .A1(n6420), .A2(n1690), .A3(n21762), .ZN(n6419) );
  NOR2_X1 U6034 ( .A1(n18784), .A2(n21881), .ZN(n9669) );
  OAI21_X1 U6039 ( .A1(n21551), .A2(n21762), .B(n21308), .ZN(n6672) );
  INV_X1 U6040 ( .I(n21765), .ZN(n1690) );
  INV_X2 U6049 ( .I(n16496), .ZN(n21668) );
  INV_X1 U6050 ( .I(n21641), .ZN(n21908) );
  CLKBUF_X2 U6051 ( .I(Key[18]), .Z(n19677) );
  CLKBUF_X2 U6052 ( .I(Key[28]), .Z(n19732) );
  CLKBUF_X2 U6056 ( .I(Key[172]), .Z(n29689) );
  AOI22_X1 U6060 ( .A1(n29340), .A2(n29339), .B1(n12848), .B2(n20481), .ZN(
        n12847) );
  INV_X4 U6071 ( .I(n12726), .ZN(n939) );
  INV_X1 U6095 ( .I(n30243), .ZN(n30192) );
  AOI21_X1 U6130 ( .A1(n984), .A2(n1205), .B(n1072), .ZN(n11147) );
  INV_X2 U6133 ( .I(n28237), .ZN(n982) );
  INV_X1 U6140 ( .I(n11694), .ZN(n27848) );
  NAND2_X1 U6146 ( .A1(n27337), .A2(n1225), .ZN(n11431) );
  AOI21_X1 U6150 ( .A1(n991), .A2(n32046), .B(n4782), .ZN(n16847) );
  INV_X1 U6163 ( .I(n35750), .ZN(n27286) );
  INV_X1 U6164 ( .I(n27446), .ZN(n27447) );
  NAND3_X1 U6203 ( .A1(n26101), .A2(n1021), .A3(n35207), .ZN(n26105) );
  NOR2_X1 U6238 ( .A1(n39599), .A2(n1024), .ZN(n25436) );
  INV_X1 U6247 ( .I(n25694), .ZN(n25630) );
  NAND2_X1 U6260 ( .A1(n24648), .A2(n15850), .ZN(n15848) );
  NAND3_X1 U6263 ( .A1(n16210), .A2(n24660), .A3(n24783), .ZN(n12133) );
  NAND2_X1 U6287 ( .A1(n1586), .A2(n18302), .ZN(n13310) );
  NAND2_X1 U6289 ( .A1(n32297), .A2(n8175), .ZN(n24340) );
  INV_X1 U6298 ( .I(n36552), .ZN(n14699) );
  NOR2_X1 U6301 ( .A1(n7273), .A2(n17709), .ZN(n23797) );
  NOR3_X1 U6303 ( .A1(n14392), .A2(n37045), .A3(n24300), .ZN(n3227) );
  BUF_X4 U6305 ( .I(n23934), .Z(n1129) );
  INV_X1 U6308 ( .I(n8116), .ZN(n20312) );
  OAI22_X1 U6325 ( .A1(n23597), .A2(n23314), .B1(n23055), .B2(n23373), .ZN(
        n23073) );
  OAI21_X1 U6351 ( .A1(n23115), .A2(n9699), .B(n1146), .ZN(n12508) );
  NAND3_X1 U6357 ( .A1(n11658), .A2(n23098), .A3(n21094), .ZN(n12473) );
  NOR2_X1 U6358 ( .A1(n33697), .A2(n35576), .ZN(n22850) );
  NAND2_X1 U6361 ( .A1(n23083), .A2(n23190), .ZN(n2163) );
  INV_X1 U6390 ( .I(n22181), .ZN(n2842) );
  OAI21_X1 U6408 ( .A1(n21906), .A2(n9886), .B(n21908), .ZN(n5305) );
  NAND3_X1 U6416 ( .A1(n21699), .A2(n1353), .A3(n19709), .ZN(n9424) );
  NOR2_X1 U6423 ( .A1(n21550), .A2(n21506), .ZN(n21765) );
  INV_X1 U6429 ( .I(n695), .ZN(n21555) );
  INV_X1 U6432 ( .I(n19516), .ZN(n1367) );
  INV_X1 U6438 ( .I(n19822), .ZN(n21539) );
  INV_X1 U6447 ( .I(n16333), .ZN(n21888) );
  INV_X1 U6449 ( .I(n29657), .ZN(n1724) );
  CLKBUF_X2 U6452 ( .I(Key[133]), .Z(n19816) );
  CLKBUF_X2 U6458 ( .I(Key[37]), .Z(n19905) );
  NOR2_X1 U6478 ( .A1(n35187), .A2(n30107), .ZN(n19033) );
  NOR2_X1 U6479 ( .A1(n4378), .A2(n30079), .ZN(n6687) );
  NOR2_X1 U6483 ( .A1(n29721), .A2(n29719), .ZN(n5779) );
  NAND3_X1 U6531 ( .A1(n9143), .A2(n30052), .A3(n1057), .ZN(n9142) );
  NAND2_X1 U6532 ( .A1(n18816), .A2(n5471), .ZN(n2860) );
  NOR2_X1 U6535 ( .A1(n29862), .A2(n38215), .ZN(n13132) );
  NOR2_X1 U6539 ( .A1(n32906), .A2(n31279), .ZN(n12880) );
  NOR3_X1 U6543 ( .A1(n30154), .A2(n5414), .A3(n892), .ZN(n5415) );
  INV_X1 U6548 ( .I(n30049), .ZN(n8731) );
  NAND2_X1 U6551 ( .A1(n30153), .A2(n30192), .ZN(n30244) );
  OR2_X1 U6569 ( .A1(n14559), .A2(n29174), .Z(n4387) );
  INV_X1 U6576 ( .I(n28983), .ZN(n1413) );
  OAI21_X1 U6586 ( .A1(n28720), .A2(n33646), .B(n4980), .ZN(n16474) );
  INV_X1 U6597 ( .I(n28454), .ZN(n12990) );
  NAND2_X1 U6601 ( .A1(n35182), .A2(n1433), .ZN(n17801) );
  NAND2_X1 U6607 ( .A1(n30304), .A2(n28728), .ZN(n28061) );
  OAI21_X1 U6612 ( .A1(n15792), .A2(n1197), .B(n10369), .ZN(n28658) );
  NAND2_X1 U6669 ( .A1(n27997), .A2(n11461), .ZN(n8523) );
  INV_X1 U6670 ( .I(n27997), .ZN(n27876) );
  INV_X1 U6675 ( .I(n14456), .ZN(n1447) );
  INV_X2 U6693 ( .I(n15410), .ZN(n18689) );
  BUF_X4 U6694 ( .I(n18474), .Z(n988) );
  INV_X2 U6698 ( .I(n15219), .ZN(n16613) );
  AND3_X1 U6706 ( .A1(n27409), .A2(n7706), .A3(n34689), .Z(n27315) );
  NOR2_X1 U6709 ( .A1(n18374), .A2(n18743), .ZN(n15918) );
  NAND2_X1 U6713 ( .A1(n27410), .A2(n32131), .ZN(n4568) );
  INV_X1 U6717 ( .I(n19529), .ZN(n20057) );
  NAND2_X1 U6743 ( .A1(n8000), .A2(n26269), .ZN(n4582) );
  INV_X1 U6746 ( .I(n27043), .ZN(n17227) );
  NAND3_X1 U6747 ( .A1(n26794), .A2(n26793), .A3(n36873), .ZN(n12170) );
  NAND2_X1 U6751 ( .A1(n26708), .A2(n5960), .ZN(n14097) );
  AND2_X1 U6759 ( .A1(n26815), .A2(n1490), .Z(n18956) );
  OAI21_X1 U6780 ( .A1(n13393), .A2(n26763), .B(n26895), .ZN(n12713) );
  INV_X2 U6790 ( .I(n17535), .ZN(n1003) );
  BUF_X2 U6793 ( .I(n26803), .Z(n1091) );
  INV_X1 U6794 ( .I(n11335), .ZN(n26936) );
  INV_X1 U6798 ( .I(n14752), .ZN(n16834) );
  INV_X2 U6804 ( .I(n26689), .ZN(n17252) );
  INV_X2 U6810 ( .I(n26478), .ZN(n1009) );
  AND2_X1 U6812 ( .A1(n6179), .A2(n25875), .Z(n6178) );
  NAND2_X1 U6827 ( .A1(n15020), .A2(n37582), .ZN(n10476) );
  NOR2_X1 U6840 ( .A1(n7110), .A2(n1101), .ZN(n15020) );
  INV_X1 U6858 ( .I(n25900), .ZN(n26122) );
  OAI21_X1 U6881 ( .A1(n25385), .A2(n10158), .B(n7284), .ZN(n25353) );
  NAND2_X1 U6886 ( .A1(n25687), .A2(n14518), .ZN(n20122) );
  NOR3_X1 U6888 ( .A1(n25574), .A2(n18031), .A3(n25614), .ZN(n12097) );
  NAND3_X1 U6895 ( .A1(n7986), .A2(n8070), .A3(n4947), .ZN(n8770) );
  NAND3_X1 U6904 ( .A1(n25036), .A2(n19785), .A3(n17894), .ZN(n8863) );
  INV_X1 U6916 ( .I(n25379), .ZN(n11951) );
  INV_X2 U6921 ( .I(n25543), .ZN(n1539) );
  NAND2_X1 U6955 ( .A1(n7693), .A2(n5388), .ZN(n5387) );
  NOR3_X1 U6960 ( .A1(n10667), .A2(n934), .A3(n17658), .ZN(n17663) );
  NOR2_X1 U6976 ( .A1(n24782), .A2(n1121), .ZN(n4775) );
  NOR3_X1 U6981 ( .A1(n39513), .A2(n16502), .A3(n5768), .ZN(n1996) );
  NAND2_X1 U6997 ( .A1(n23797), .A2(n1586), .ZN(n5740) );
  INV_X2 U7011 ( .I(n30447), .ZN(n1595) );
  AND2_X1 U7026 ( .A1(n24223), .A2(n24088), .Z(n24089) );
  INV_X1 U7031 ( .I(n24327), .ZN(n24229) );
  INV_X1 U7034 ( .I(n205), .ZN(n1280) );
  INV_X1 U7038 ( .I(n12519), .ZN(n17081) );
  INV_X4 U7042 ( .I(n24241), .ZN(n1033) );
  NOR2_X1 U7057 ( .A1(n5044), .A2(n33747), .ZN(n23575) );
  OAI21_X1 U7071 ( .A1(n13830), .A2(n23506), .B(n13833), .ZN(n13829) );
  NAND3_X1 U7075 ( .A1(n35808), .A2(n9823), .A3(n5083), .ZN(n4290) );
  NAND2_X1 U7085 ( .A1(n960), .A2(n14477), .ZN(n23748) );
  OAI21_X1 U7090 ( .A1(n21247), .A2(n11970), .B(n1862), .ZN(n1861) );
  NOR2_X1 U7098 ( .A1(n33840), .A2(n14477), .ZN(n8239) );
  NAND2_X1 U7107 ( .A1(n34506), .A2(n23472), .ZN(n23746) );
  NAND3_X1 U7120 ( .A1(n14234), .A2(n22934), .A3(n9699), .ZN(n8101) );
  NAND3_X1 U7133 ( .A1(n15151), .A2(n23099), .A3(n20570), .ZN(n12472) );
  NOR3_X1 U7139 ( .A1(n1647), .A2(n38524), .A3(n19865), .ZN(n20362) );
  OAI21_X1 U7145 ( .A1(n16419), .A2(n1646), .B(n19469), .ZN(n13093) );
  NAND3_X1 U7147 ( .A1(n11913), .A2(n22937), .A3(n1141), .ZN(n11912) );
  NAND2_X1 U7148 ( .A1(n15330), .A2(n23098), .ZN(n22905) );
  OAI21_X1 U7149 ( .A1(n5581), .A2(n17226), .B(n1313), .ZN(n13640) );
  NAND2_X1 U7166 ( .A1(n22993), .A2(n22866), .ZN(n14749) );
  INV_X1 U7173 ( .I(n12315), .ZN(n1646) );
  INV_X1 U7174 ( .I(n22857), .ZN(n22890) );
  OR2_X2 U7183 ( .A1(n2386), .A2(n2384), .Z(n2383) );
  NOR2_X1 U7191 ( .A1(n39075), .A2(n1149), .ZN(n13570) );
  NAND2_X1 U7192 ( .A1(n21002), .A2(n21001), .ZN(n21000) );
  NAND3_X1 U7193 ( .A1(n11345), .A2(n1812), .A3(n1866), .ZN(n1865) );
  NAND2_X1 U7195 ( .A1(n3840), .A2(n17530), .ZN(n21958) );
  NOR2_X1 U7200 ( .A1(n7916), .A2(n22239), .ZN(n8118) );
  NAND3_X1 U7207 ( .A1(n31940), .A2(n11327), .A3(n1672), .ZN(n22218) );
  INV_X1 U7214 ( .I(n22243), .ZN(n22241) );
  NAND3_X1 U7218 ( .A1(n32107), .A2(n4239), .A3(n2910), .ZN(n8623) );
  INV_X1 U7228 ( .I(n22019), .ZN(n22084) );
  INV_X1 U7231 ( .I(n18303), .ZN(n17086) );
  BUF_X2 U7233 ( .I(n22041), .Z(n2839) );
  BUF_X4 U7237 ( .I(n17440), .Z(n1048) );
  INV_X1 U7239 ( .I(n22113), .ZN(n13191) );
  OAI21_X1 U7243 ( .A1(n21901), .A2(n21902), .B(n35921), .ZN(n5822) );
  NAND2_X1 U7255 ( .A1(n18576), .A2(n20266), .ZN(n2157) );
  AND2_X1 U7257 ( .A1(n21401), .A2(n668), .Z(n9705) );
  NAND2_X1 U7259 ( .A1(n21817), .A2(n32820), .ZN(n21479) );
  INV_X1 U7268 ( .I(n21606), .ZN(n2645) );
  INV_X1 U7277 ( .I(n21550), .ZN(n21763) );
  INV_X1 U7279 ( .I(n21352), .ZN(n4094) );
  INV_X1 U7291 ( .I(n13679), .ZN(n21521) );
  NOR2_X1 U7292 ( .A1(n20778), .A2(n19496), .ZN(n21561) );
  INV_X1 U7294 ( .I(n30104), .ZN(n1163) );
  CLKBUF_X2 U7295 ( .I(n21330), .Z(n21697) );
  INV_X1 U7297 ( .I(n30150), .ZN(n1161) );
  BUF_X2 U7298 ( .I(n21938), .Z(n8700) );
  INV_X1 U7302 ( .I(n29970), .ZN(n1162) );
  INV_X1 U7303 ( .I(n19805), .ZN(n1167) );
  INV_X1 U7307 ( .I(n30126), .ZN(n1165) );
  INV_X1 U7308 ( .I(n29831), .ZN(n1169) );
  CLKBUF_X2 U7309 ( .I(Key[183]), .Z(n30126) );
  CLKBUF_X2 U7312 ( .I(Key[75]), .Z(n30179) );
  CLKBUF_X2 U7320 ( .I(Key[27]), .Z(n29371) );
  NAND3_X1 U7324 ( .A1(n37632), .A2(n939), .A3(n13142), .ZN(n12452) );
  NAND2_X1 U7331 ( .A1(n29874), .A2(n17286), .ZN(n10293) );
  NAND2_X1 U7332 ( .A1(n29881), .A2(n17286), .ZN(n10292) );
  OR2_X1 U7334 ( .A1(n35180), .A2(n16084), .Z(n16083) );
  NAND2_X1 U7340 ( .A1(n37632), .A2(n939), .ZN(n11973) );
  AOI21_X1 U7341 ( .A1(n18039), .A2(n15509), .B(n939), .ZN(n12033) );
  NAND2_X1 U7342 ( .A1(n31160), .A2(n8955), .ZN(n5813) );
  NAND2_X1 U7349 ( .A1(n31569), .A2(n29929), .ZN(n29912) );
  INV_X1 U7351 ( .I(n31569), .ZN(n8561) );
  INV_X1 U7354 ( .I(n29722), .ZN(n5951) );
  NOR2_X1 U7357 ( .A1(n30086), .A2(n30096), .ZN(n2484) );
  AND2_X1 U7376 ( .A1(n2858), .A2(n5579), .Z(n2507) );
  NOR2_X1 U7377 ( .A1(n4377), .A2(n30076), .ZN(n30056) );
  AOI22_X1 U7378 ( .A1(n29708), .A2(n29721), .B1(n29720), .B2(n14337), .ZN(
        n16577) );
  INV_X1 U7383 ( .I(n4449), .ZN(n4447) );
  NOR2_X1 U7384 ( .A1(n3861), .A2(n5579), .ZN(n2073) );
  INV_X1 U7387 ( .I(n13786), .ZN(n11701) );
  NOR2_X1 U7392 ( .A1(n12081), .A2(n19544), .ZN(n6863) );
  NOR2_X1 U7405 ( .A1(n12940), .A2(n33928), .ZN(n15584) );
  NOR2_X1 U7406 ( .A1(n1177), .A2(n1399), .ZN(n2321) );
  NAND3_X1 U7411 ( .A1(n11415), .A2(n30046), .A3(n30162), .ZN(n3819) );
  OAI21_X1 U7416 ( .A1(n9572), .A2(n13132), .B(n18104), .ZN(n9569) );
  NOR2_X1 U7421 ( .A1(n31511), .A2(n37061), .ZN(n28744) );
  AOI21_X1 U7430 ( .A1(n2160), .A2(n8529), .B(n16224), .ZN(n18445) );
  INV_X1 U7433 ( .I(n30232), .ZN(n15062) );
  NAND2_X1 U7436 ( .A1(n19137), .A2(n29892), .ZN(n6803) );
  NOR2_X1 U7450 ( .A1(n19050), .A2(n30220), .ZN(n4807) );
  NOR2_X1 U7455 ( .A1(n21167), .A2(n39828), .ZN(n15301) );
  AND2_X1 U7456 ( .A1(n18816), .A2(n3631), .Z(n4445) );
  NAND2_X1 U7457 ( .A1(n29998), .A2(n30043), .ZN(n4858) );
  AND3_X1 U7464 ( .A1(n19765), .A2(n10590), .A3(n30229), .Z(n9996) );
  NAND2_X1 U7465 ( .A1(n17597), .A2(n19783), .ZN(n29317) );
  NOR2_X1 U7473 ( .A1(n30238), .A2(n31788), .ZN(n11886) );
  INV_X1 U7496 ( .I(n4341), .ZN(n29048) );
  NOR2_X1 U7506 ( .A1(n28360), .A2(n14677), .ZN(n16475) );
  OAI21_X1 U7520 ( .A1(n35172), .A2(n28484), .B(n32543), .ZN(n6694) );
  INV_X2 U7524 ( .I(n5115), .ZN(n1065) );
  OAI22_X1 U7533 ( .A1(n28765), .A2(n35203), .B1(n28812), .B2(n5465), .ZN(
        n12545) );
  NOR2_X1 U7537 ( .A1(n1431), .A2(n28553), .ZN(n8759) );
  NAND3_X1 U7548 ( .A1(n15447), .A2(n39355), .A3(n19827), .ZN(n6071) );
  NAND2_X1 U7551 ( .A1(n976), .A2(n35203), .ZN(n8914) );
  NAND2_X1 U7559 ( .A1(n9329), .A2(n17771), .ZN(n10676) );
  NAND3_X1 U7563 ( .A1(n15112), .A2(n9141), .A3(n5093), .ZN(n16183) );
  INV_X1 U7564 ( .I(n1882), .ZN(n18369) );
  NOR2_X1 U7571 ( .A1(n5383), .A2(n39435), .ZN(n12611) );
  NOR2_X1 U7576 ( .A1(n2790), .A2(n28723), .ZN(n2785) );
  NOR2_X1 U7580 ( .A1(n28323), .A2(n30304), .ZN(n17596) );
  INV_X1 U7600 ( .I(n28569), .ZN(n28614) );
  NAND2_X1 U7608 ( .A1(n10825), .A2(n27980), .ZN(n10824) );
  NAND2_X1 U7618 ( .A1(n8787), .A2(n20445), .ZN(n28612) );
  OAI21_X1 U7637 ( .A1(n28064), .A2(n16513), .B(n981), .ZN(n6980) );
  AOI21_X1 U7638 ( .A1(n27624), .A2(n37056), .B(n16576), .ZN(n7365) );
  AOI21_X1 U7641 ( .A1(n16576), .A2(n8960), .B(n35694), .ZN(n9170) );
  NAND3_X1 U7653 ( .A1(n10836), .A2(n983), .A3(n28050), .ZN(n10443) );
  NAND2_X1 U7660 ( .A1(n27900), .A2(n16461), .ZN(n8525) );
  AND2_X1 U7672 ( .A1(n14397), .A2(n1200), .Z(n4456) );
  NAND2_X1 U7673 ( .A1(n2716), .A2(n5266), .ZN(n5905) );
  NOR2_X1 U7679 ( .A1(n37), .A2(n1448), .ZN(n11838) );
  INV_X1 U7726 ( .I(n27964), .ZN(n28137) );
  BUF_X2 U7736 ( .I(n16339), .Z(n11461) );
  INV_X1 U7747 ( .I(n17378), .ZN(n27997) );
  INV_X1 U7749 ( .I(n39442), .ZN(n7755) );
  INV_X1 U7753 ( .I(n27556), .ZN(n14325) );
  INV_X1 U7755 ( .I(n27574), .ZN(n1215) );
  NAND2_X1 U7765 ( .A1(n30871), .A2(n35115), .ZN(n18050) );
  AOI21_X1 U7768 ( .A1(n26941), .A2(n12156), .B(n18489), .ZN(n26942) );
  AND2_X1 U7787 ( .A1(n4434), .A2(n34689), .Z(n11735) );
  OR2_X1 U7789 ( .A1(n39065), .A2(n1470), .Z(n26967) );
  OAI21_X1 U7791 ( .A1(n33593), .A2(n36496), .B(n16782), .ZN(n4231) );
  NAND2_X1 U7794 ( .A1(n992), .A2(n1227), .ZN(n2259) );
  AND2_X1 U7822 ( .A1(n34562), .A2(n19203), .Z(n4610) );
  NOR3_X1 U7831 ( .A1(n20402), .A2(n17795), .A3(n27123), .ZN(n6415) );
  NOR2_X1 U7837 ( .A1(n33503), .A2(n7975), .ZN(n6975) );
  INV_X2 U7838 ( .I(n7611), .ZN(n12156) );
  OAI21_X1 U7840 ( .A1(n26767), .A2(n9690), .B(n33396), .ZN(n8331) );
  OR2_X1 U7843 ( .A1(n11467), .A2(n14412), .Z(n3809) );
  NOR2_X1 U7849 ( .A1(n26639), .A2(n17515), .ZN(n26767) );
  NOR2_X1 U7854 ( .A1(n26859), .A2(n32256), .ZN(n14469) );
  OAI21_X1 U7864 ( .A1(n19206), .A2(n19207), .B(n38797), .ZN(n9891) );
  OR2_X1 U7865 ( .A1(n13854), .A2(n26988), .Z(n13334) );
  NOR2_X1 U7883 ( .A1(n19448), .A2(n8556), .ZN(n11130) );
  NAND2_X1 U7885 ( .A1(n3350), .A2(n7527), .ZN(n3349) );
  NAND2_X1 U7889 ( .A1(n26962), .A2(n17601), .ZN(n17600) );
  NAND3_X1 U7893 ( .A1(n13605), .A2(n5405), .A3(n35912), .ZN(n26642) );
  AND2_X1 U7900 ( .A1(n26922), .A2(n26895), .Z(n26304) );
  AND2_X1 U7923 ( .A1(n26961), .A2(n20936), .Z(n3224) );
  OAI21_X1 U7929 ( .A1(n14355), .A2(n7752), .B(n3351), .ZN(n3350) );
  INV_X1 U7955 ( .I(n26666), .ZN(n26179) );
  NAND2_X1 U7959 ( .A1(n11105), .A2(n26598), .ZN(n3098) );
  AND2_X1 U7974 ( .A1(n26000), .A2(n13971), .Z(n16239) );
  NAND2_X1 U7981 ( .A1(n16200), .A2(n1017), .ZN(n10138) );
  NOR2_X1 U7987 ( .A1(n2835), .A2(n2833), .ZN(n2832) );
  AND2_X1 U7995 ( .A1(n25847), .A2(n1514), .Z(n11770) );
  OAI21_X1 U8005 ( .A1(n25867), .A2(n37306), .B(n26022), .ZN(n21198) );
  OAI21_X1 U8011 ( .A1(n4190), .A2(n26125), .B(n929), .ZN(n6883) );
  NAND3_X1 U8023 ( .A1(n31192), .A2(n2888), .A3(n4772), .ZN(n12448) );
  NAND2_X1 U8025 ( .A1(n18289), .A2(n26075), .ZN(n26076) );
  AND2_X1 U8048 ( .A1(n1521), .A2(n2534), .Z(n11386) );
  NAND2_X1 U8056 ( .A1(n26029), .A2(n18320), .ZN(n25922) );
  NAND2_X1 U8063 ( .A1(n31133), .A2(n31626), .ZN(n8255) );
  OAI21_X1 U8064 ( .A1(n8883), .A2(n18142), .B(n17791), .ZN(n7732) );
  INV_X2 U8073 ( .I(n18320), .ZN(n1102) );
  BUF_X2 U8074 ( .I(n7136), .Z(n7110) );
  OR2_X1 U8089 ( .A1(n13467), .A2(n954), .Z(n13466) );
  NAND3_X1 U8091 ( .A1(n5860), .A2(n32105), .A3(n25452), .ZN(n5858) );
  NAND2_X1 U8097 ( .A1(n4455), .A2(n13129), .ZN(n4452) );
  NOR2_X1 U8101 ( .A1(n728), .A2(n2799), .ZN(n5455) );
  NAND2_X1 U8113 ( .A1(n1539), .A2(n25482), .ZN(n2250) );
  NAND3_X1 U8115 ( .A1(n1253), .A2(n16677), .A3(n24896), .ZN(n17303) );
  AND2_X1 U8119 ( .A1(n17029), .A2(n36708), .Z(n9429) );
  NOR2_X1 U8121 ( .A1(n5227), .A2(n12500), .ZN(n5010) );
  OAI22_X1 U8135 ( .A1(n14081), .A2(n14082), .B1(n25642), .B2(n25674), .ZN(
        n14056) );
  NAND3_X1 U8143 ( .A1(n1545), .A2(n6747), .A3(n25361), .ZN(n9145) );
  OAI21_X1 U8155 ( .A1(n16933), .A2(n25482), .B(n25548), .ZN(n10786) );
  INV_X1 U8179 ( .I(n20924), .ZN(n25533) );
  OR2_X1 U8180 ( .A1(n15052), .A2(n15051), .Z(n25548) );
  INV_X1 U8186 ( .I(n25722), .ZN(n25721) );
  BUF_X4 U8190 ( .I(n3785), .Z(n25361) );
  INV_X2 U8196 ( .I(n825), .ZN(n1257) );
  INV_X1 U8198 ( .I(n11497), .ZN(n7876) );
  INV_X1 U8201 ( .I(n25176), .ZN(n1554) );
  NAND3_X1 U8203 ( .A1(n25203), .A2(n7968), .A3(n7969), .ZN(n3653) );
  OR2_X1 U8208 ( .A1(n20800), .A2(n4973), .Z(n16747) );
  NAND2_X1 U8215 ( .A1(n7065), .A2(n24608), .ZN(n4908) );
  NOR2_X1 U8244 ( .A1(n7693), .A2(n10116), .ZN(n20689) );
  AND2_X1 U8249 ( .A1(n24887), .A2(n15467), .Z(n16745) );
  NOR2_X1 U8263 ( .A1(n7286), .A2(n19420), .ZN(n8954) );
  INV_X1 U8274 ( .I(n24565), .ZN(n1573) );
  INV_X2 U8277 ( .I(n24673), .ZN(n16547) );
  NOR2_X1 U8284 ( .A1(n1586), .A2(n37227), .ZN(n19027) );
  AOI21_X1 U8290 ( .A1(n4666), .A2(n24153), .B(n16377), .ZN(n24154) );
  OAI21_X1 U8291 ( .A1(n19466), .A2(n24303), .B(n21310), .ZN(n11170) );
  NOR3_X1 U8293 ( .A1(n15240), .A2(n12975), .A3(n1608), .ZN(n20653) );
  INV_X1 U8294 ( .I(n3133), .ZN(n8175) );
  NOR2_X1 U8300 ( .A1(n12366), .A2(n7086), .ZN(n7085) );
  OR2_X1 U8317 ( .A1(n6933), .A2(n33450), .Z(n12974) );
  NAND2_X1 U8322 ( .A1(n33712), .A2(n24245), .ZN(n24582) );
  NOR2_X1 U8323 ( .A1(n24274), .A2(n35954), .ZN(n5358) );
  OAI21_X1 U8327 ( .A1(n12975), .A2(n24087), .B(n1608), .ZN(n7406) );
  INV_X1 U8331 ( .I(n38224), .ZN(n19653) );
  INV_X2 U8341 ( .I(n39816), .ZN(n1596) );
  CLKBUF_X2 U8357 ( .I(n39814), .Z(n7440) );
  AOI22_X1 U8371 ( .A1(n21251), .A2(n21130), .B1(n1633), .B2(n21250), .ZN(
        n12175) );
  NAND2_X1 U8375 ( .A1(n3715), .A2(n31644), .ZN(n2919) );
  NOR3_X1 U8380 ( .A1(n10480), .A2(n9395), .A3(n33496), .ZN(n1918) );
  NOR2_X1 U8385 ( .A1(n1290), .A2(n9862), .ZN(n12851) );
  OAI21_X1 U8388 ( .A1(n20841), .A2(n1308), .B(n33349), .ZN(n17442) );
  NOR2_X1 U8421 ( .A1(n36810), .A2(n33703), .ZN(n23243) );
  NAND2_X1 U8431 ( .A1(n19559), .A2(n13733), .ZN(n1862) );
  INV_X4 U8439 ( .I(n2600), .ZN(n23567) );
  INV_X1 U8443 ( .I(n23516), .ZN(n1623) );
  OAI22_X1 U8466 ( .A1(n20637), .A2(n23209), .B1(n5464), .B2(n23135), .ZN(
        n23136) );
  NAND2_X1 U8469 ( .A1(n35442), .A2(n8812), .ZN(n19181) );
  NOR2_X1 U8470 ( .A1(n1319), .A2(n1654), .ZN(n6500) );
  OAI21_X1 U8473 ( .A1(n1645), .A2(n23124), .B(n22875), .ZN(n13450) );
  NOR2_X1 U8486 ( .A1(n22890), .A2(n22682), .ZN(n15242) );
  NAND2_X1 U8489 ( .A1(n38601), .A2(n23212), .ZN(n3041) );
  OR2_X1 U8494 ( .A1(n18229), .A2(n19697), .Z(n13337) );
  OR2_X1 U8512 ( .A1(n39810), .A2(n2047), .Z(n2049) );
  OAI21_X1 U8517 ( .A1(n19440), .A2(n19134), .B(n23124), .ZN(n14187) );
  INV_X1 U8542 ( .I(n34757), .ZN(n23172) );
  INV_X2 U8545 ( .I(n13572), .ZN(n1145) );
  INV_X1 U8548 ( .I(n23122), .ZN(n11295) );
  BUF_X2 U8552 ( .I(n12315), .Z(n5657) );
  AND2_X2 U8563 ( .A1(n5205), .A2(n5204), .Z(n5203) );
  NAND2_X1 U8564 ( .A1(n37089), .A2(n34808), .ZN(n4851) );
  NAND2_X1 U8568 ( .A1(n22340), .A2(n20238), .ZN(n10630) );
  NOR2_X1 U8569 ( .A1(n30800), .A2(n11329), .ZN(n7896) );
  NAND2_X1 U8570 ( .A1(n22143), .A2(n34808), .ZN(n8753) );
  NAND2_X1 U8574 ( .A1(n19261), .A2(n1329), .ZN(n5877) );
  AND3_X1 U8580 ( .A1(n31940), .A2(n11171), .A3(n22361), .Z(n4800) );
  NAND2_X1 U8584 ( .A1(n32889), .A2(n5929), .ZN(n21969) );
  NOR2_X1 U8585 ( .A1(n11329), .A2(n5302), .ZN(n9484) );
  OR2_X1 U8598 ( .A1(n32889), .A2(n5929), .Z(n11511) );
  NOR2_X1 U8599 ( .A1(n21503), .A2(n30306), .ZN(n19453) );
  NAND2_X1 U8605 ( .A1(n474), .A2(n14349), .ZN(n2211) );
  NOR2_X1 U8610 ( .A1(n6576), .A2(n36397), .ZN(n5617) );
  NOR2_X1 U8612 ( .A1(n32107), .A2(n14423), .ZN(n8622) );
  NAND2_X1 U8614 ( .A1(n17685), .A2(n12077), .ZN(n12930) );
  NAND3_X1 U8615 ( .A1(n18360), .A2(n1344), .A3(n22086), .ZN(n9341) );
  NOR2_X1 U8620 ( .A1(n2839), .A2(n1338), .ZN(n14028) );
  NAND2_X1 U8621 ( .A1(n19958), .A2(n6297), .ZN(n14233) );
  NOR2_X1 U8627 ( .A1(n1338), .A2(n18303), .ZN(n7434) );
  AOI21_X1 U8629 ( .A1(n6347), .A2(n22019), .B(n36006), .ZN(n5462) );
  INV_X2 U8632 ( .I(n4179), .ZN(n12814) );
  NOR2_X1 U8635 ( .A1(n6347), .A2(n2696), .ZN(n21664) );
  BUF_X2 U8636 ( .I(n22497), .Z(n7131) );
  NAND4_X1 U8638 ( .A1(n5304), .A2(n5303), .A3(n5305), .A4(n7608), .ZN(n5302)
         );
  NAND2_X1 U8641 ( .A1(n7357), .A2(n22364), .ZN(n12169) );
  INV_X2 U8649 ( .I(n22354), .ZN(n1152) );
  NAND3_X1 U8650 ( .A1(n2278), .A2(n21817), .A3(n2092), .ZN(n2276) );
  OAI22_X1 U8656 ( .A1(n13701), .A2(n21898), .B1(n21838), .B2(n10120), .ZN(
        n10085) );
  AOI22_X1 U8659 ( .A1(n543), .A2(n6418), .B1(n33771), .B2(n21765), .ZN(n6417)
         );
  AOI22_X1 U8667 ( .A1(n15031), .A2(n275), .B1(n21440), .B2(n18152), .ZN(n5823) );
  OR2_X1 U8668 ( .A1(n2759), .A2(n18219), .Z(n9746) );
  NAND3_X1 U8669 ( .A1(n20898), .A2(n21899), .A3(n21897), .ZN(n3438) );
  NAND2_X1 U8670 ( .A1(n38011), .A2(n5531), .ZN(n5023) );
  NOR2_X1 U8676 ( .A1(n18774), .A2(n14373), .ZN(n19554) );
  NOR2_X1 U8685 ( .A1(n9642), .A2(n20328), .ZN(n15706) );
  NOR2_X1 U8688 ( .A1(n33771), .A2(n21761), .ZN(n6418) );
  NOR2_X1 U8692 ( .A1(n1346), .A2(n5751), .ZN(n9286) );
  NOR2_X1 U8693 ( .A1(n15839), .A2(n3784), .ZN(n15523) );
  NAND2_X1 U8696 ( .A1(n7703), .A2(n7654), .ZN(n10822) );
  INV_X1 U8700 ( .I(n21475), .ZN(n6350) );
  NAND2_X1 U8701 ( .A1(n33154), .A2(n21912), .ZN(n13437) );
  NOR2_X1 U8704 ( .A1(n8799), .A2(n21898), .ZN(n15369) );
  NAND2_X1 U8706 ( .A1(n8293), .A2(n21339), .ZN(n7367) );
  AND2_X1 U8707 ( .A1(n21666), .A2(n690), .Z(n10464) );
  INV_X1 U8709 ( .I(n21905), .ZN(n21462) );
  INV_X1 U8710 ( .I(n21894), .ZN(n21581) );
  INV_X1 U8720 ( .I(n21898), .ZN(n1694) );
  NAND2_X1 U8724 ( .A1(n7304), .A2(n526), .ZN(n16035) );
  INV_X2 U8725 ( .I(n18450), .ZN(n21897) );
  INV_X1 U8726 ( .I(n13997), .ZN(n18496) );
  NOR2_X1 U8727 ( .A1(n19395), .A2(n21875), .ZN(n11916) );
  AOI21_X1 U8728 ( .A1(n21546), .A2(n21696), .B(n21330), .ZN(n11917) );
  INV_X1 U8732 ( .I(n29649), .ZN(n1708) );
  INV_X1 U8733 ( .I(n19804), .ZN(n1371) );
  INV_X1 U8734 ( .I(n29666), .ZN(n1361) );
  INV_X1 U8735 ( .I(n15370), .ZN(n12044) );
  INV_X1 U8737 ( .I(n19683), .ZN(n1356) );
  INV_X1 U8739 ( .I(n19720), .ZN(n1370) );
  INV_X1 U8740 ( .I(n19622), .ZN(n1358) );
  INV_X1 U8741 ( .I(n29506), .ZN(n1357) );
  INV_X1 U8744 ( .I(n30010), .ZN(n1374) );
  BUF_X2 U8746 ( .I(n19871), .Z(n20328) );
  INV_X1 U8750 ( .I(n18270), .ZN(n23591) );
  INV_X1 U8752 ( .I(n19800), .ZN(n1366) );
  INV_X1 U8753 ( .I(n29978), .ZN(n1368) );
  CLKBUF_X2 U8756 ( .I(Key[62]), .Z(n19800) );
  CLKBUF_X2 U8759 ( .I(Key[153]), .Z(n19786) );
  CLKBUF_X2 U8762 ( .I(Key[157]), .Z(n19720) );
  CLKBUF_X2 U8763 ( .I(Key[24]), .Z(n19925) );
  CLKBUF_X2 U8764 ( .I(Key[17]), .Z(n30101) );
  CLKBUF_X2 U8765 ( .I(Key[118]), .Z(n19683) );
  CLKBUF_X2 U8767 ( .I(Key[15]), .Z(n30016) );
  CLKBUF_X2 U8768 ( .I(Key[10]), .Z(n19622) );
  CLKBUF_X2 U8772 ( .I(Key[94]), .Z(n19516) );
  CLKBUF_X2 U8773 ( .I(Key[168]), .Z(n19902) );
  CLKBUF_X2 U8781 ( .I(Key[173]), .Z(n19940) );
  CLKBUF_X2 U8789 ( .I(Key[78]), .Z(n19629) );
  CLKBUF_X2 U8790 ( .I(Key[113]), .Z(n29538) );
  NAND3_X1 U8794 ( .A1(n29369), .A2(n11067), .A3(n15768), .ZN(n4669) );
  OAI21_X1 U8795 ( .A1(n1380), .A2(n6147), .B(n7600), .ZN(n16472) );
  NOR2_X1 U8802 ( .A1(n17369), .A2(n16598), .ZN(n16597) );
  NOR2_X1 U8804 ( .A1(n2489), .A2(n6147), .ZN(n2488) );
  INV_X1 U8806 ( .I(n1385), .ZN(n11448) );
  AOI21_X1 U8808 ( .A1(n969), .A2(n38200), .B(n6341), .ZN(n6340) );
  INV_X1 U8811 ( .I(n29219), .ZN(n1378) );
  OAI21_X1 U8812 ( .A1(n29812), .A2(n29811), .B(n38141), .ZN(n6441) );
  AOI21_X1 U8815 ( .A1(n11898), .A2(n29859), .B(n36764), .ZN(n2506) );
  OAI21_X1 U8816 ( .A1(n15601), .A2(n8955), .B(n968), .ZN(n11972) );
  AOI21_X1 U8818 ( .A1(n8561), .A2(n19097), .B(n18081), .ZN(n8560) );
  AOI21_X1 U8819 ( .A1(n29851), .A2(n11898), .B(n29855), .ZN(n5580) );
  BUF_X2 U8826 ( .I(n33966), .Z(n10003) );
  NAND2_X1 U8828 ( .A1(n29318), .A2(n38156), .ZN(n9627) );
  AOI21_X1 U8829 ( .A1(n6147), .A2(n30096), .B(n13559), .ZN(n6149) );
  NAND2_X1 U8830 ( .A1(n13442), .A2(n29574), .ZN(n14075) );
  NOR2_X1 U8832 ( .A1(n2944), .A2(n5579), .ZN(n29846) );
  OAI21_X1 U8834 ( .A1(n29756), .A2(n29754), .B(n29739), .ZN(n8063) );
  INV_X2 U8838 ( .I(n29980), .ZN(n1170) );
  OAI21_X1 U8849 ( .A1(n30192), .A2(n30153), .B(n30152), .ZN(n5300) );
  NAND2_X1 U8857 ( .A1(n28996), .A2(n1057), .ZN(n7167) );
  NOR3_X1 U8859 ( .A1(n31629), .A2(n6019), .A3(n34179), .ZN(n6372) );
  AOI21_X1 U8860 ( .A1(n6851), .A2(n8918), .B(n32946), .ZN(n12992) );
  NAND2_X1 U8864 ( .A1(n7208), .A2(n4169), .ZN(n21052) );
  NOR2_X1 U8873 ( .A1(n29777), .A2(n17726), .ZN(n15424) );
  NOR2_X1 U8876 ( .A1(n7789), .A2(n29059), .ZN(n7989) );
  NAND2_X1 U8878 ( .A1(n29595), .A2(n1404), .ZN(n6254) );
  NOR2_X1 U8881 ( .A1(n16907), .A2(n7790), .ZN(n7479) );
  NOR2_X1 U8882 ( .A1(n29904), .A2(n6204), .ZN(n6203) );
  NOR2_X1 U8883 ( .A1(n1402), .A2(n29776), .ZN(n7448) );
  NOR2_X1 U8886 ( .A1(n21074), .A2(n30041), .ZN(n9817) );
  NOR2_X1 U8888 ( .A1(n30041), .A2(n21074), .ZN(n20125) );
  NOR2_X1 U8890 ( .A1(n5736), .A2(n3986), .ZN(n3154) );
  BUF_X2 U8893 ( .I(n14438), .Z(n2121) );
  NOR2_X1 U8897 ( .A1(n29992), .A2(n775), .ZN(n3169) );
  NOR2_X1 U8898 ( .A1(n1060), .A2(n29699), .ZN(n9000) );
  NOR2_X1 U8899 ( .A1(n14891), .A2(n18667), .ZN(n11635) );
  INV_X1 U8910 ( .I(n29450), .ZN(n29418) );
  INV_X1 U8917 ( .I(n29907), .ZN(n29955) );
  INV_X2 U8919 ( .I(n29493), .ZN(n1179) );
  INV_X1 U8920 ( .I(n16009), .ZN(n19994) );
  NAND3_X1 U8928 ( .A1(n28632), .A2(n28634), .A3(n14209), .ZN(n28636) );
  NAND2_X1 U8937 ( .A1(n10303), .A2(n32014), .ZN(n10302) );
  NAND3_X1 U8945 ( .A1(n28453), .A2(n13379), .A3(n9668), .ZN(n13378) );
  NOR2_X1 U8948 ( .A1(n28759), .A2(n3014), .ZN(n28408) );
  NAND2_X1 U8955 ( .A1(n17800), .A2(n11164), .ZN(n14239) );
  AOI21_X1 U8964 ( .A1(n8093), .A2(n3845), .B(n28473), .ZN(n8159) );
  NOR2_X1 U8965 ( .A1(n28514), .A2(n28716), .ZN(n5243) );
  INV_X2 U8968 ( .I(n9878), .ZN(n11488) );
  NAND2_X1 U8971 ( .A1(n5343), .A2(n28735), .ZN(n5342) );
  NOR2_X1 U8974 ( .A1(n2639), .A2(n8476), .ZN(n13061) );
  NAND2_X1 U8986 ( .A1(n28570), .A2(n39020), .ZN(n19322) );
  INV_X1 U9004 ( .I(n28715), .ZN(n28509) );
  NAND2_X1 U9005 ( .A1(n3899), .A2(n979), .ZN(n4119) );
  INV_X2 U9013 ( .I(n9597), .ZN(n13508) );
  NOR2_X1 U9022 ( .A1(n39786), .A2(n32080), .ZN(n11743) );
  OAI21_X1 U9031 ( .A1(n28048), .A2(n28258), .B(n11025), .ZN(n11024) );
  NOR2_X1 U9049 ( .A1(n27915), .A2(n1451), .ZN(n19748) );
  NOR2_X1 U9053 ( .A1(n11461), .A2(n28001), .ZN(n8801) );
  OR2_X1 U9054 ( .A1(n1439), .A2(n1441), .Z(n18777) );
  NAND2_X1 U9063 ( .A1(n28206), .A2(n156), .ZN(n4977) );
  NOR2_X1 U9072 ( .A1(n32783), .A2(n15357), .ZN(n10236) );
  NOR2_X1 U9077 ( .A1(n28258), .A2(n34410), .ZN(n27883) );
  NOR2_X1 U9083 ( .A1(n28236), .A2(n2262), .ZN(n4153) );
  NAND3_X1 U9086 ( .A1(n27894), .A2(n17410), .A3(n28273), .ZN(n20639) );
  NAND2_X1 U9090 ( .A1(n36517), .A2(n13366), .ZN(n11407) );
  NOR3_X1 U9094 ( .A1(n13927), .A2(n11461), .A3(n28200), .ZN(n13906) );
  AND2_X1 U9102 ( .A1(n15357), .A2(n1447), .Z(n14615) );
  NAND2_X1 U9103 ( .A1(n28236), .A2(n28237), .ZN(n12623) );
  INV_X1 U9104 ( .I(n38202), .ZN(n3511) );
  NOR2_X1 U9116 ( .A1(n17410), .A2(n14399), .ZN(n12477) );
  NAND2_X1 U9117 ( .A1(n12257), .A2(n28230), .ZN(n27063) );
  INV_X2 U9137 ( .I(n18383), .ZN(n1212) );
  INV_X2 U9142 ( .I(n15287), .ZN(n1214) );
  NAND2_X1 U9151 ( .A1(n9037), .A2(n27395), .ZN(n3851) );
  NOR2_X1 U9156 ( .A1(n38488), .A2(n6191), .ZN(n7499) );
  NAND3_X1 U9159 ( .A1(n13213), .A2(n7975), .A3(n7676), .ZN(n21232) );
  NAND2_X1 U9160 ( .A1(n27084), .A2(n5675), .ZN(n16360) );
  NOR2_X1 U9163 ( .A1(n9488), .A2(n1481), .ZN(n9487) );
  NOR2_X1 U9176 ( .A1(n1473), .A2(n17132), .ZN(n17422) );
  AND2_X1 U9184 ( .A1(n26074), .A2(n1470), .Z(n11485) );
  OAI21_X1 U9185 ( .A1(n10581), .A2(n9633), .B(n38193), .ZN(n10577) );
  NAND2_X1 U9199 ( .A1(n39628), .A2(n15616), .ZN(n7921) );
  NAND2_X1 U9208 ( .A1(n27285), .A2(n33254), .ZN(n10284) );
  NAND2_X1 U9211 ( .A1(n1480), .A2(n33503), .ZN(n27119) );
  OR2_X1 U9213 ( .A1(n19455), .A2(n27197), .Z(n6507) );
  NAND2_X1 U9221 ( .A1(n5089), .A2(n27284), .ZN(n27285) );
  NOR2_X1 U9224 ( .A1(n27357), .A2(n15360), .ZN(n5559) );
  NAND2_X1 U9231 ( .A1(n7975), .A2(n9144), .ZN(n6972) );
  NOR2_X1 U9235 ( .A1(n27127), .A2(n27126), .ZN(n27128) );
  NAND2_X1 U9247 ( .A1(n12373), .A2(n9690), .ZN(n4325) );
  NOR2_X1 U9252 ( .A1(n15594), .A2(n26804), .ZN(n10891) );
  OAI21_X1 U9256 ( .A1(n32168), .A2(n26970), .B(n2226), .ZN(n26250) );
  NOR2_X1 U9263 ( .A1(n2079), .A2(n36801), .ZN(n2078) );
  NAND2_X1 U9269 ( .A1(n18870), .A2(n15485), .ZN(n26750) );
  NOR3_X1 U9275 ( .A1(n20120), .A2(n26802), .A3(n8479), .ZN(n2801) );
  NAND3_X1 U9278 ( .A1(n33333), .A2(n6606), .A3(n26932), .ZN(n14457) );
  NOR2_X1 U9295 ( .A1(n19762), .A2(n36882), .ZN(n18901) );
  AND2_X1 U9296 ( .A1(n26719), .A2(n10111), .Z(n26471) );
  OR2_X1 U9298 ( .A1(n20936), .A2(n33858), .Z(n12505) );
  NAND2_X1 U9304 ( .A1(n34160), .A2(n26968), .ZN(n2079) );
  NAND2_X1 U9306 ( .A1(n17515), .A2(n6454), .ZN(n16402) );
  NOR2_X1 U9312 ( .A1(n26862), .A2(n17712), .ZN(n9731) );
  AOI21_X1 U9313 ( .A1(n26783), .A2(n8814), .B(n8817), .ZN(n26784) );
  INV_X2 U9314 ( .I(n26768), .ZN(n10355) );
  NOR2_X1 U9332 ( .A1(n26734), .A2(n4138), .ZN(n10202) );
  NAND2_X1 U9337 ( .A1(n14382), .A2(n13004), .ZN(n7778) );
  NAND3_X1 U9338 ( .A1(n13777), .A2(n875), .A3(n26937), .ZN(n18024) );
  INV_X1 U9342 ( .I(n3449), .ZN(n26773) );
  NOR2_X1 U9347 ( .A1(n34005), .A2(n26901), .ZN(n5174) );
  INV_X1 U9352 ( .I(n9117), .ZN(n26910) );
  INV_X2 U9354 ( .I(n11188), .ZN(n26961) );
  INV_X2 U9355 ( .I(n20974), .ZN(n26935) );
  BUF_X2 U9356 ( .I(n26713), .Z(n19425) );
  AOI22_X1 U9368 ( .A1(n25846), .A2(n25928), .B1(n25847), .B2(n26116), .ZN(
        n12489) );
  NAND3_X1 U9372 ( .A1(n11552), .A2(n18406), .A3(n318), .ZN(n25896) );
  NOR2_X1 U9376 ( .A1(n25928), .A2(n4154), .ZN(n7544) );
  OAI21_X1 U9377 ( .A1(n25971), .A2(n951), .B(n14215), .ZN(n3916) );
  OAI21_X1 U9381 ( .A1(n31192), .A2(n7961), .B(n26088), .ZN(n20490) );
  OAI21_X1 U9386 ( .A1(n25868), .A2(n31375), .B(n5885), .ZN(n5884) );
  OR2_X1 U9392 ( .A1(n25822), .A2(n1511), .Z(n14660) );
  OAI21_X1 U9399 ( .A1(n26125), .A2(n4190), .B(n4515), .ZN(n26011) );
  NOR2_X1 U9403 ( .A1(n14703), .A2(n6222), .ZN(n12449) );
  NAND3_X1 U9406 ( .A1(n31375), .A2(n26020), .A3(n25867), .ZN(n5885) );
  NAND3_X1 U9423 ( .A1(n38247), .A2(n18801), .A3(n25820), .ZN(n25706) );
  NAND2_X1 U9427 ( .A1(n36546), .A2(n2888), .ZN(n14703) );
  NOR2_X1 U9429 ( .A1(n25829), .A2(n17624), .ZN(n6062) );
  NOR2_X1 U9431 ( .A1(n26055), .A2(n38198), .ZN(n25744) );
  NAND2_X1 U9433 ( .A1(n26185), .A2(n38185), .ZN(n17952) );
  INV_X1 U9438 ( .I(n25936), .ZN(n26130) );
  NOR2_X1 U9441 ( .A1(n19121), .A2(n35138), .ZN(n19120) );
  INV_X1 U9445 ( .I(n4382), .ZN(n4385) );
  NAND2_X1 U9466 ( .A1(n25349), .A2(n25073), .ZN(n25108) );
  OAI21_X1 U9471 ( .A1(n15543), .A2(n15541), .B(n15542), .ZN(n15184) );
  OR2_X1 U9480 ( .A1(n35157), .A2(n15541), .Z(n25593) );
  AOI21_X1 U9481 ( .A1(n4726), .A2(n25575), .B(n25574), .ZN(n16466) );
  NAND2_X1 U9484 ( .A1(n19095), .A2(n19171), .ZN(n20358) );
  NOR3_X1 U9485 ( .A1(n12896), .A2(n6747), .A3(n25361), .ZN(n6748) );
  AOI22_X1 U9486 ( .A1(n8879), .A2(n31780), .B1(n953), .B2(n1548), .ZN(n12062)
         );
  OAI22_X1 U9490 ( .A1(n1117), .A2(n25380), .B1(n19863), .B2(n1109), .ZN(n7173) );
  INV_X1 U9492 ( .I(n33950), .ZN(n18894) );
  NAND2_X1 U9493 ( .A1(n25571), .A2(n19235), .ZN(n19234) );
  NAND2_X1 U9494 ( .A1(n25480), .A2(n10786), .ZN(n10785) );
  NAND3_X1 U9496 ( .A1(n18298), .A2(n25649), .A3(n32291), .ZN(n25650) );
  NAND2_X1 U9513 ( .A1(n13218), .A2(n19235), .ZN(n20876) );
  NAND2_X1 U9519 ( .A1(n25481), .A2(n25543), .ZN(n12625) );
  NAND2_X1 U9521 ( .A1(n1535), .A2(n10938), .ZN(n6762) );
  NOR2_X1 U9522 ( .A1(n6696), .A2(n7583), .ZN(n6763) );
  NAND2_X1 U9524 ( .A1(n25601), .A2(n33947), .ZN(n3058) );
  NAND2_X1 U9526 ( .A1(n34576), .A2(n17594), .ZN(n2721) );
  NOR2_X1 U9533 ( .A1(n220), .A2(n2366), .ZN(n3005) );
  NOR2_X1 U9542 ( .A1(n37050), .A2(n1552), .ZN(n8738) );
  OAI21_X1 U9543 ( .A1(n19581), .A2(n12825), .B(n20052), .ZN(n10082) );
  NOR2_X1 U9552 ( .A1(n5541), .A2(n31509), .ZN(n5483) );
  NOR2_X1 U9558 ( .A1(n14436), .A2(n835), .ZN(n6573) );
  INV_X1 U9576 ( .I(n25552), .ZN(n12828) );
  INV_X1 U9582 ( .I(n21031), .ZN(n17183) );
  NAND2_X1 U9586 ( .A1(n1560), .A2(n11601), .ZN(n7263) );
  INV_X1 U9589 ( .I(n25218), .ZN(n24873) );
  INV_X2 U9590 ( .I(n33132), .ZN(n1258) );
  INV_X1 U9598 ( .I(n19670), .ZN(n6598) );
  NOR2_X1 U9602 ( .A1(n16745), .A2(n17270), .ZN(n20000) );
  INV_X2 U9606 ( .I(n19691), .ZN(n1261) );
  INV_X2 U9610 ( .I(n25140), .ZN(n1262) );
  NOR2_X1 U9616 ( .A1(n13583), .A2(n24806), .ZN(n13582) );
  NAND2_X1 U9620 ( .A1(n1567), .A2(n7831), .ZN(n24491) );
  NAND2_X1 U9622 ( .A1(n7248), .A2(n38073), .ZN(n7245) );
  NAND2_X1 U9631 ( .A1(n6273), .A2(n24529), .ZN(n1784) );
  NAND2_X1 U9633 ( .A1(n1583), .A2(n7177), .ZN(n7176) );
  NAND2_X1 U9635 ( .A1(n19484), .A2(n24680), .ZN(n6335) );
  AOI21_X1 U9642 ( .A1(n24692), .A2(n30764), .B(n24717), .ZN(n6539) );
  AOI21_X1 U9643 ( .A1(n35250), .A2(n37395), .B(n14211), .ZN(n20505) );
  NAND2_X1 U9647 ( .A1(n24785), .A2(n32045), .ZN(n13817) );
  INV_X1 U9658 ( .I(n24613), .ZN(n1567) );
  NOR2_X1 U9659 ( .A1(n1583), .A2(n16238), .ZN(n8803) );
  AOI21_X1 U9663 ( .A1(n19431), .A2(n34458), .B(n37341), .ZN(n13553) );
  OAI21_X1 U9664 ( .A1(n20155), .A2(n24712), .B(n19279), .ZN(n20154) );
  NOR2_X1 U9670 ( .A1(n38749), .A2(n24515), .ZN(n24776) );
  NOR2_X1 U9673 ( .A1(n1030), .A2(n3697), .ZN(n4176) );
  NAND2_X1 U9677 ( .A1(n24707), .A2(n34526), .ZN(n6274) );
  INV_X1 U9678 ( .I(n24866), .ZN(n19339) );
  INV_X2 U9683 ( .I(n20728), .ZN(n14999) );
  NAND2_X1 U9684 ( .A1(n24148), .A2(n24274), .ZN(n5360) );
  NAND2_X1 U9687 ( .A1(n8846), .A2(n1598), .ZN(n8845) );
  AOI21_X1 U9712 ( .A1(n6998), .A2(n13692), .B(n1595), .ZN(n6997) );
  OAI21_X1 U9719 ( .A1(n24272), .A2(n1604), .B(n24273), .ZN(n10713) );
  AOI21_X1 U9721 ( .A1(n38224), .A2(n8690), .B(n12692), .ZN(n9362) );
  NAND2_X1 U9731 ( .A1(n24231), .A2(n1127), .ZN(n18256) );
  NOR2_X1 U9737 ( .A1(n13808), .A2(n1598), .ZN(n9634) );
  OAI21_X1 U9751 ( .A1(n24406), .A2(n37934), .B(n24410), .ZN(n18615) );
  OAI22_X1 U9762 ( .A1(n16884), .A2(n1596), .B1(n250), .B2(n24442), .ZN(n10783) );
  NAND2_X1 U9763 ( .A1(n39467), .A2(n19880), .ZN(n9584) );
  NAND2_X1 U9765 ( .A1(n19402), .A2(n6515), .ZN(n9822) );
  NAND2_X1 U9776 ( .A1(n4243), .A2(n36500), .ZN(n3453) );
  NOR2_X1 U9784 ( .A1(n18304), .A2(n7210), .ZN(n24123) );
  NOR2_X1 U9795 ( .A1(n24146), .A2(n232), .ZN(n12692) );
  OR2_X1 U9797 ( .A1(n13144), .A2(n30280), .Z(n23855) );
  INV_X1 U9799 ( .I(n24445), .ZN(n24448) );
  INV_X2 U9807 ( .I(n15865), .ZN(n24469) );
  NAND2_X1 U9813 ( .A1(n24294), .A2(n33939), .ZN(n24297) );
  BUF_X2 U9826 ( .I(n24431), .Z(n12975) );
  INV_X1 U9832 ( .I(n23794), .ZN(n23670) );
  NAND2_X1 U9839 ( .A1(n23751), .A2(n11452), .ZN(n23987) );
  NOR2_X1 U9846 ( .A1(n12638), .A2(n23399), .ZN(n11723) );
  NAND2_X1 U9857 ( .A1(n2961), .A2(n23588), .ZN(n2960) );
  NOR2_X1 U9865 ( .A1(n1918), .A2(n23622), .ZN(n1917) );
  NOR2_X1 U9866 ( .A1(n23251), .A2(n23592), .ZN(n17888) );
  NOR2_X1 U9868 ( .A1(n4207), .A2(n14235), .ZN(n10840) );
  NAND2_X1 U9880 ( .A1(n52), .A2(n33496), .ZN(n15842) );
  NAND2_X1 U9881 ( .A1(n23243), .A2(n38981), .ZN(n12641) );
  INV_X1 U9885 ( .I(n11669), .ZN(n4637) );
  NOR2_X1 U9887 ( .A1(n32424), .A2(n1635), .ZN(n6993) );
  OAI21_X1 U9889 ( .A1(n32377), .A2(n23578), .B(n1138), .ZN(n10612) );
  INV_X1 U9899 ( .I(n23637), .ZN(n23641) );
  NOR2_X1 U9915 ( .A1(n16443), .A2(n35506), .ZN(n9621) );
  NAND3_X1 U9916 ( .A1(n37622), .A2(n38042), .A3(n23515), .ZN(n11842) );
  NAND2_X1 U9922 ( .A1(n4207), .A2(n14235), .ZN(n10711) );
  NOR2_X1 U9924 ( .A1(n23458), .A2(n23238), .ZN(n4707) );
  NAND3_X1 U9929 ( .A1(n6303), .A2(n6176), .A3(n23484), .ZN(n23362) );
  NOR2_X1 U9935 ( .A1(n20835), .A2(n16013), .ZN(n13602) );
  INV_X1 U9937 ( .I(n38724), .ZN(n19665) );
  OAI21_X1 U9945 ( .A1(n36829), .A2(n30574), .B(n37014), .ZN(n9796) );
  INV_X1 U9949 ( .I(n23517), .ZN(n6373) );
  NAND2_X1 U9953 ( .A1(n7335), .A2(n23624), .ZN(n3498) );
  NAND2_X1 U9966 ( .A1(n6827), .A2(n6826), .ZN(n11245) );
  OAI22_X1 U9967 ( .A1(n2049), .A2(n1989), .B1(n20439), .B2(n23146), .ZN(
        n23147) );
  INV_X1 U9970 ( .I(n3713), .ZN(n3717) );
  NAND2_X1 U9972 ( .A1(n6916), .A2(n20373), .ZN(n4959) );
  AOI21_X1 U9978 ( .A1(n6581), .A2(n4472), .B(n15388), .ZN(n6826) );
  NOR2_X1 U9979 ( .A1(n19469), .A2(n8462), .ZN(n8461) );
  NAND3_X1 U9991 ( .A1(n17131), .A2(n22368), .A3(n1143), .ZN(n6916) );
  AOI21_X1 U10002 ( .A1(n11307), .A2(n23111), .B(n12392), .ZN(n13262) );
  OR3_X1 U10004 ( .A1(n8809), .A2(n32677), .A3(n31300), .Z(n22805) );
  AND2_X1 U10005 ( .A1(n38524), .A2(n1647), .Z(n2927) );
  AND3_X1 U10011 ( .A1(n37791), .A2(n22368), .A3(n2047), .Z(n5942) );
  NOR2_X1 U10013 ( .A1(n1650), .A2(n6499), .ZN(n6498) );
  NAND2_X1 U10014 ( .A1(n1645), .A2(n14187), .ZN(n14186) );
  NAND2_X1 U10022 ( .A1(n23214), .A2(n4472), .ZN(n3040) );
  NAND2_X1 U10025 ( .A1(n22682), .A2(n22921), .ZN(n13515) );
  NAND2_X1 U10033 ( .A1(n272), .A2(n1655), .ZN(n21062) );
  NOR2_X1 U10034 ( .A1(n17080), .A2(n22920), .ZN(n22922) );
  NAND2_X1 U10038 ( .A1(n22890), .A2(n17080), .ZN(n22924) );
  NOR2_X1 U10046 ( .A1(n5657), .A2(n19645), .ZN(n8458) );
  AND3_X1 U10050 ( .A1(n33934), .A2(n19586), .A3(n33745), .Z(n23187) );
  AND2_X1 U10051 ( .A1(n18750), .A2(n3273), .Z(n3543) );
  INV_X1 U10058 ( .I(n12925), .ZN(n22901) );
  NOR2_X1 U10060 ( .A1(n9472), .A2(n10074), .ZN(n22860) );
  INV_X1 U10062 ( .I(n23088), .ZN(n23090) );
  NAND2_X1 U10066 ( .A1(n12392), .A2(n23108), .ZN(n13339) );
  NOR2_X1 U10068 ( .A1(n23111), .A2(n23110), .ZN(n23112) );
  NOR2_X1 U10069 ( .A1(n8197), .A2(n12630), .ZN(n22908) );
  NOR2_X1 U10076 ( .A1(n22709), .A2(n550), .ZN(n5214) );
  NOR2_X1 U10077 ( .A1(n18708), .A2(n1654), .ZN(n4162) );
  NOR2_X1 U10079 ( .A1(n3906), .A2(n23142), .ZN(n2116) );
  NAND2_X1 U10083 ( .A1(n1648), .A2(n16104), .ZN(n20175) );
  CLKBUF_X2 U10090 ( .I(n22897), .Z(n10074) );
  INV_X1 U10107 ( .I(n22862), .ZN(n18708) );
  INV_X1 U10114 ( .I(n22610), .ZN(n2838) );
  OAI21_X1 U10115 ( .A1(n13565), .A2(n13566), .B(n22348), .ZN(n3024) );
  INV_X1 U10117 ( .I(n22622), .ZN(n1657) );
  INV_X1 U10118 ( .I(n22657), .ZN(n1660) );
  NAND2_X1 U10129 ( .A1(n19515), .A2(n12023), .ZN(n8343) );
  NAND2_X1 U10131 ( .A1(n22055), .A2(n8089), .ZN(n13765) );
  OAI21_X1 U10137 ( .A1(n22143), .A2(n8754), .B(n8753), .ZN(n8752) );
  NAND2_X1 U10153 ( .A1(n5053), .A2(n22286), .ZN(n3954) );
  NOR2_X1 U10154 ( .A1(n11542), .A2(n22388), .ZN(n5204) );
  OAI21_X1 U10156 ( .A1(n21958), .A2(n17531), .B(n16989), .ZN(n2386) );
  NAND2_X1 U10160 ( .A1(n1672), .A2(n5617), .ZN(n5616) );
  NAND2_X1 U10161 ( .A1(n35822), .A2(n12793), .ZN(n12812) );
  OAI22_X1 U10165 ( .A1(n31092), .A2(n22324), .B1(n1812), .B2(n22323), .ZN(
        n21830) );
  NAND2_X1 U10171 ( .A1(n21090), .A2(n22326), .ZN(n8342) );
  NAND2_X1 U10179 ( .A1(n22181), .A2(n2840), .ZN(n9843) );
  AOI21_X1 U10181 ( .A1(n4239), .A2(n19873), .B(n14423), .ZN(n5207) );
  AND2_X1 U10183 ( .A1(n11149), .A2(n19773), .Z(n12023) );
  NAND2_X1 U10188 ( .A1(n7955), .A2(n12230), .ZN(n7818) );
  NOR2_X1 U10193 ( .A1(n37217), .A2(n22132), .ZN(n14311) );
  NAND2_X1 U10194 ( .A1(n6128), .A2(n22295), .ZN(n5497) );
  AND2_X1 U10198 ( .A1(n22265), .A2(n19515), .Z(n13900) );
  NAND2_X1 U10210 ( .A1(n9387), .A2(n1688), .ZN(n11013) );
  NAND2_X1 U10211 ( .A1(n1686), .A2(n36371), .ZN(n14020) );
  NAND2_X1 U10212 ( .A1(n8520), .A2(n8518), .ZN(n5053) );
  AOI21_X1 U10218 ( .A1(n33168), .A2(n9422), .B(n20376), .ZN(n21363) );
  AND2_X1 U10219 ( .A1(n1680), .A2(n6128), .Z(n13627) );
  AND2_X1 U10222 ( .A1(n22143), .A2(n37089), .Z(n8687) );
  AOI21_X1 U10238 ( .A1(n33860), .A2(n22177), .B(n6451), .ZN(n5878) );
  AND2_X1 U10241 ( .A1(n35526), .A2(n22264), .Z(n19211) );
  NAND2_X1 U10256 ( .A1(n22226), .A2(n22225), .ZN(n20123) );
  AND2_X1 U10261 ( .A1(n19373), .A2(n9165), .Z(n22249) );
  OAI21_X1 U10264 ( .A1(n33168), .A2(n5821), .B(n31649), .ZN(n21364) );
  NAND2_X1 U10272 ( .A1(n3325), .A2(n21583), .ZN(n3323) );
  NAND2_X1 U10278 ( .A1(n3676), .A2(n32817), .ZN(n3680) );
  NOR2_X1 U10280 ( .A1(n33168), .A2(n19017), .ZN(n20374) );
  OAI22_X1 U10289 ( .A1(n3692), .A2(n938), .B1(n1155), .B2(n5132), .ZN(n3691)
         );
  AOI21_X1 U10296 ( .A1(n8438), .A2(n21838), .B(n1159), .ZN(n8442) );
  NOR2_X1 U10297 ( .A1(n10875), .A2(n37678), .ZN(n10125) );
  INV_X2 U10302 ( .I(n8040), .ZN(n1342) );
  NOR3_X1 U10303 ( .A1(n38546), .A2(n21712), .A3(n17266), .ZN(n17265) );
  AOI21_X1 U10305 ( .A1(n21551), .A2(n19871), .B(n21550), .ZN(n11238) );
  AND2_X1 U10306 ( .A1(n21654), .A2(n6732), .Z(n12546) );
  AOI22_X1 U10312 ( .A1(n8598), .A2(n19543), .B1(n17792), .B2(n8600), .ZN(
        n15382) );
  AOI22_X1 U10318 ( .A1(n8466), .A2(n19323), .B1(n8468), .B2(n670), .ZN(n5417)
         );
  OAI21_X1 U10319 ( .A1(n21911), .A2(n21910), .B(n21909), .ZN(n7608) );
  AOI21_X1 U10322 ( .A1(n21665), .A2(n919), .B(n21833), .ZN(n9319) );
  NAND2_X1 U10324 ( .A1(n21723), .A2(n1689), .ZN(n4924) );
  AOI22_X1 U10328 ( .A1(n1156), .A2(n21691), .B1(n21690), .B2(n21339), .ZN(
        n7998) );
  NAND2_X1 U10330 ( .A1(n13996), .A2(n13998), .ZN(n12513) );
  NOR2_X1 U10334 ( .A1(n21410), .A2(n21804), .ZN(n21371) );
  INV_X1 U10339 ( .I(n21885), .ZN(n2045) );
  OAI21_X1 U10340 ( .A1(n18542), .A2(n17792), .B(n21561), .ZN(n21562) );
  INV_X1 U10342 ( .I(n20328), .ZN(n21764) );
  AND2_X1 U10344 ( .A1(n1159), .A2(n21897), .Z(n11008) );
  AOI21_X1 U10346 ( .A1(n17848), .A2(n21450), .B(n17242), .ZN(n17544) );
  NAND2_X1 U10347 ( .A1(n21784), .A2(n37111), .ZN(n18339) );
  NOR2_X1 U10349 ( .A1(n19620), .A2(n8936), .ZN(n8434) );
  OAI22_X1 U10351 ( .A1(n293), .A2(n670), .B1(n18412), .B2(n34867), .ZN(n13098) );
  OAI21_X1 U10352 ( .A1(n7935), .A2(n21923), .B(n4116), .ZN(n5187) );
  AND2_X1 U10354 ( .A1(n21565), .A2(n17534), .Z(n3912) );
  NAND2_X1 U10357 ( .A1(n1816), .A2(n15839), .ZN(n13859) );
  NAND2_X1 U10358 ( .A1(n1816), .A2(n15338), .ZN(n13861) );
  NOR3_X1 U10360 ( .A1(n917), .A2(n21928), .A3(n19372), .ZN(n7640) );
  NAND2_X1 U10362 ( .A1(n33771), .A2(n21762), .ZN(n17886) );
  NAND2_X1 U10364 ( .A1(n21640), .A2(n21923), .ZN(n4925) );
  OAI21_X1 U10367 ( .A1(n275), .A2(n21440), .B(n16035), .ZN(n21442) );
  NOR2_X1 U10368 ( .A1(n21887), .A2(n19850), .ZN(n5980) );
  NOR2_X1 U10369 ( .A1(n21450), .A2(n1694), .ZN(n16901) );
  AND2_X1 U10373 ( .A1(n1694), .A2(n452), .Z(n12439) );
  NAND2_X1 U10375 ( .A1(n21899), .A2(n10120), .ZN(n11007) );
  INV_X1 U10379 ( .I(n37200), .ZN(n2277) );
  INV_X1 U10390 ( .I(n1697), .ZN(n8951) );
  INV_X1 U10392 ( .I(n21688), .ZN(n1693) );
  NAND2_X1 U10395 ( .A1(n21893), .A2(n3294), .ZN(n3295) );
  NOR2_X1 U10396 ( .A1(n37200), .A2(n20266), .ZN(n2187) );
  NAND2_X1 U10397 ( .A1(n21730), .A2(n10211), .ZN(n21554) );
  BUF_X2 U10400 ( .I(n21577), .Z(n19238) );
  NOR2_X1 U10401 ( .A1(n2533), .A2(n2532), .ZN(n2531) );
  BUF_X2 U10403 ( .I(n21750), .Z(n21889) );
  INV_X1 U10404 ( .I(n19733), .ZN(n1734) );
  INV_X1 U10405 ( .I(n19874), .ZN(n1695) );
  INV_X1 U10408 ( .I(n19616), .ZN(n1710) );
  INV_X1 U10410 ( .I(n29785), .ZN(n1711) );
  INV_X1 U10415 ( .I(n28831), .ZN(n1723) );
  INV_X1 U10421 ( .I(n19527), .ZN(n1707) );
  INV_X1 U10422 ( .I(n19722), .ZN(n1714) );
  INV_X1 U10424 ( .I(n21428), .ZN(n21682) );
  CLKBUF_X2 U10425 ( .I(n10212), .Z(n9863) );
  INV_X1 U10430 ( .I(n19770), .ZN(n1700) );
  INV_X1 U10432 ( .I(n29509), .ZN(n1699) );
  INV_X1 U10433 ( .I(n29647), .ZN(n1725) );
  INV_X1 U10436 ( .I(n29357), .ZN(n1717) );
  CLKBUF_X2 U10438 ( .I(Key[174]), .Z(n29785) );
  CLKBUF_X2 U10440 ( .I(Key[188]), .Z(n29221) );
  CLKBUF_X2 U10443 ( .I(Key[38]), .Z(n29808) );
  CLKBUF_X2 U10444 ( .I(Key[90]), .Z(n29711) );
  CLKBUF_X2 U10446 ( .I(Key[104]), .Z(n30253) );
  CLKBUF_X2 U10449 ( .I(Key[26]), .Z(n29334) );
  CLKBUF_X2 U10453 ( .I(Key[191]), .Z(n29357) );
  CLKBUF_X2 U10455 ( .I(Key[182]), .Z(n30114) );
  CLKBUF_X2 U10459 ( .I(Key[144]), .Z(n19616) );
  CLKBUF_X2 U10460 ( .I(Key[116]), .Z(n29657) );
  CLKBUF_X2 U10461 ( .I(Key[158]), .Z(n19831) );
  CLKBUF_X2 U10463 ( .I(Key[125]), .Z(n30063) );
  CLKBUF_X2 U10466 ( .I(Key[135]), .Z(n29285) );
  CLKBUF_X2 U10469 ( .I(Key[55]), .Z(n19929) );
  CLKBUF_X2 U10470 ( .I(Key[48]), .Z(n30207) );
  CLKBUF_X2 U10471 ( .I(Key[149]), .Z(n29875) );
  CLKBUF_X2 U10472 ( .I(Key[179]), .Z(n30006) );
  CLKBUF_X2 U10474 ( .I(Key[117]), .Z(n29680) );
  CLKBUF_X2 U10477 ( .I(Key[23]), .Z(n19770) );
  CLKBUF_X2 U10478 ( .I(Key[68]), .Z(n29920) );
  CLKBUF_X2 U10479 ( .I(Key[185]), .Z(n30203) );
  CLKBUF_X2 U10481 ( .I(Key[119]), .Z(n28831) );
  CLKBUF_X2 U10484 ( .I(Key[136]), .Z(n19733) );
  CLKBUF_X2 U10485 ( .I(Key[122]), .Z(n28910) );
  CLKBUF_X2 U10486 ( .I(Key[56]), .Z(n29141) );
  CLKBUF_X2 U10487 ( .I(Key[2]), .Z(n29474) );
  CLKBUF_X2 U10488 ( .I(Key[77]), .Z(n19875) );
  CLKBUF_X2 U10490 ( .I(Key[29]), .Z(n29463) );
  CLKBUF_X2 U10492 ( .I(Key[105]), .Z(n29206) );
  NOR2_X1 U10493 ( .A1(n5369), .A2(n30010), .ZN(n5194) );
  NAND2_X1 U10497 ( .A1(n12942), .A2(n29369), .ZN(n29362) );
  NAND2_X1 U10510 ( .A1(n6440), .A2(n29802), .ZN(n6438) );
  AOI21_X1 U10513 ( .A1(n14073), .A2(n29572), .B(n14072), .ZN(n29573) );
  AOI21_X1 U10515 ( .A1(n12033), .A2(n5813), .B(n5811), .ZN(n15600) );
  AOI21_X1 U10516 ( .A1(n29543), .A2(n29560), .B(n21177), .ZN(n29019) );
  OR2_X1 U10519 ( .A1(n9591), .A2(n29932), .Z(n16187) );
  NAND2_X1 U10522 ( .A1(n9837), .A2(n19380), .ZN(n29552) );
  NAND2_X1 U10526 ( .A1(n7015), .A2(n5970), .ZN(n6440) );
  AOI21_X1 U10532 ( .A1(n3287), .A2(n29318), .B(n3285), .ZN(n3284) );
  AOI21_X1 U10540 ( .A1(n29372), .A2(n29373), .B(n29355), .ZN(n15957) );
  NAND2_X1 U10542 ( .A1(n18041), .A2(n31538), .ZN(n3118) );
  NOR2_X1 U10543 ( .A1(n6342), .A2(n29468), .ZN(n6341) );
  OAI21_X1 U10544 ( .A1(n19097), .A2(n29922), .B(n8560), .ZN(n18085) );
  AOI21_X1 U10546 ( .A1(n29932), .A2(n29922), .B(n1174), .ZN(n29919) );
  OAI22_X1 U10550 ( .A1(n30099), .A2(n30098), .B1(n30097), .B2(n6149), .ZN(
        n6148) );
  OAI21_X1 U10554 ( .A1(n14007), .A2(n4910), .B(n29807), .ZN(n29809) );
  NAND2_X1 U10561 ( .A1(n6843), .A2(n16233), .ZN(n11394) );
  NAND2_X1 U10562 ( .A1(n29207), .A2(n920), .ZN(n13143) );
  OAI22_X1 U10565 ( .A1(n5580), .A2(n29860), .B1(n1171), .B2(n8727), .ZN(n5065) );
  NAND2_X1 U10567 ( .A1(n29923), .A2(n39709), .ZN(n21283) );
  NOR2_X1 U10571 ( .A1(n14009), .A2(n14008), .ZN(n4910) );
  NAND2_X1 U10574 ( .A1(n29540), .A2(n29541), .ZN(n7435) );
  NAND2_X1 U10575 ( .A1(n29846), .A2(n29851), .ZN(n5108) );
  NOR2_X1 U10579 ( .A1(n21146), .A2(n29739), .ZN(n8064) );
  NAND2_X1 U10580 ( .A1(n29275), .A2(n3378), .ZN(n6842) );
  NAND2_X1 U10581 ( .A1(n29795), .A2(n32050), .ZN(n5467) );
  AOI21_X1 U10582 ( .A1(n19090), .A2(n16233), .B(n29277), .ZN(n16232) );
  NAND2_X1 U10589 ( .A1(n14414), .A2(n15841), .ZN(n12340) );
  OAI21_X1 U10590 ( .A1(n29437), .A2(n29441), .B(n29433), .ZN(n12339) );
  NAND2_X1 U10591 ( .A1(n13363), .A2(n30257), .ZN(n30247) );
  NOR3_X1 U10592 ( .A1(n29677), .A2(n20672), .A3(n1173), .ZN(n9610) );
  NAND2_X1 U10597 ( .A1(n29670), .A2(n5067), .ZN(n2110) );
  NAND2_X1 U10598 ( .A1(n29979), .A2(n29980), .ZN(n5018) );
  NOR2_X1 U10600 ( .A1(n969), .A2(n29477), .ZN(n9103) );
  INV_X1 U10603 ( .I(n15259), .ZN(n11940) );
  NAND2_X1 U10605 ( .A1(n12301), .A2(n30183), .ZN(n10513) );
  AOI21_X1 U10606 ( .A1(n2113), .A2(n29675), .B(n2112), .ZN(n2111) );
  INV_X2 U10609 ( .I(n7303), .ZN(n13433) );
  AOI21_X1 U10611 ( .A1(n19663), .A2(n1172), .B(n11700), .ZN(n13991) );
  NAND2_X1 U10612 ( .A1(n8955), .A2(n13142), .ZN(n13014) );
  NOR2_X1 U10615 ( .A1(n2944), .A2(n2858), .ZN(n2205) );
  AND2_X1 U10616 ( .A1(n6720), .A2(n16803), .Z(n11182) );
  INV_X1 U10619 ( .I(n3614), .ZN(n3611) );
  AND2_X1 U10621 ( .A1(n29806), .A2(n38141), .Z(n14007) );
  NAND2_X1 U10622 ( .A1(n29858), .A2(n3725), .ZN(n2945) );
  OAI21_X1 U10626 ( .A1(n29439), .A2(n15841), .B(n18502), .ZN(n15131) );
  NAND2_X1 U10630 ( .A1(n17192), .A2(n17469), .ZN(n9264) );
  OR2_X1 U10631 ( .A1(n8287), .A2(n20274), .Z(n10289) );
  INV_X1 U10632 ( .I(n8063), .ZN(n8062) );
  INV_X1 U10633 ( .I(n36096), .ZN(n29791) );
  INV_X1 U10635 ( .I(n30033), .ZN(n18780) );
  AND4_X1 U10636 ( .A1(n29273), .A2(n29272), .A3(n29270), .A4(n29271), .Z(
        n29274) );
  OR2_X1 U10641 ( .A1(n29407), .A2(n9790), .Z(n20131) );
  NAND2_X1 U10642 ( .A1(n16683), .A2(n9839), .ZN(n7376) );
  AOI21_X1 U10643 ( .A1(n31539), .A2(n29683), .B(n18042), .ZN(n29674) );
  AND4_X1 U10648 ( .A1(n30174), .A2(n10101), .A3(n30173), .A4(n30172), .Z(
        n30175) );
  OR2_X1 U10654 ( .A1(n17262), .A2(n29574), .Z(n29572) );
  CLKBUF_X2 U10667 ( .I(n29687), .Z(n5067) );
  INV_X1 U10670 ( .I(n29687), .ZN(n29676) );
  NAND2_X1 U10684 ( .A1(n9573), .A2(n29957), .ZN(n9570) );
  NAND2_X1 U10690 ( .A1(n20436), .A2(n20435), .ZN(n20434) );
  OAI22_X1 U10698 ( .A1(n29499), .A2(n36275), .B1(n29498), .B2(n29497), .ZN(
        n29503) );
  NAND2_X1 U10700 ( .A1(n5300), .A2(n33784), .ZN(n5299) );
  INV_X1 U10706 ( .I(n9885), .ZN(n9884) );
  INV_X1 U10707 ( .I(n4220), .ZN(n9818) );
  OAI21_X1 U10712 ( .A1(n16116), .A2(n1179), .B(n4655), .ZN(n29496) );
  NAND2_X1 U10722 ( .A1(n37544), .A2(n15584), .ZN(n15583) );
  NAND2_X1 U10728 ( .A1(n18658), .A2(n19994), .ZN(n6257) );
  INV_X1 U10731 ( .I(n14281), .ZN(n12657) );
  AOI21_X1 U10733 ( .A1(n39830), .A2(n21023), .B(n344), .ZN(n20435) );
  NOR2_X1 U10736 ( .A1(n15267), .A2(n7194), .ZN(n7191) );
  NOR2_X1 U10741 ( .A1(n30152), .A2(n33784), .ZN(n10976) );
  NAND2_X1 U10743 ( .A1(n29702), .A2(n9000), .ZN(n8999) );
  OAI21_X1 U10746 ( .A1(n7790), .A2(n30240), .B(n31603), .ZN(n8338) );
  INV_X1 U10748 ( .I(n13069), .ZN(n11218) );
  NOR2_X1 U10752 ( .A1(n2001), .A2(n19878), .ZN(n9572) );
  OAI21_X1 U10755 ( .A1(n2001), .A2(n29960), .B(n29955), .ZN(n9573) );
  INV_X1 U10762 ( .I(n7166), .ZN(n7163) );
  NAND2_X1 U10765 ( .A1(n34086), .A2(n7167), .ZN(n7164) );
  NAND2_X1 U10769 ( .A1(n13657), .A2(n12992), .ZN(n12991) );
  NAND2_X1 U10770 ( .A1(n13942), .A2(n16116), .ZN(n7614) );
  NAND2_X1 U10774 ( .A1(n8477), .A2(n29997), .ZN(n8419) );
  NAND2_X1 U10775 ( .A1(n7448), .A2(n29779), .ZN(n21038) );
  NOR2_X1 U10780 ( .A1(n30153), .A2(n1059), .ZN(n8716) );
  NOR2_X1 U10784 ( .A1(n21168), .A2(n21167), .ZN(n21166) );
  OR2_X1 U10788 ( .A1(n6851), .A2(n8918), .Z(n10452) );
  NOR2_X1 U10792 ( .A1(n8529), .A2(n30049), .ZN(n29864) );
  OR2_X1 U10794 ( .A1(n29643), .A2(n19734), .Z(n29485) );
  NAND2_X1 U10796 ( .A1(n14151), .A2(n29494), .ZN(n28902) );
  OAI21_X1 U10800 ( .A1(n34006), .A2(n20979), .B(n19962), .ZN(n28885) );
  NAND2_X1 U10806 ( .A1(n1059), .A2(n30192), .ZN(n8031) );
  OAI21_X1 U10807 ( .A1(n29006), .A2(n1058), .B(n29992), .ZN(n13069) );
  NOR2_X1 U10809 ( .A1(n3700), .A2(n5471), .ZN(n3246) );
  AND2_X1 U10813 ( .A1(n19508), .A2(n3700), .Z(n29703) );
  CLKBUF_X2 U10816 ( .I(n37083), .Z(n10101) );
  NAND2_X1 U10826 ( .A1(n9872), .A2(n10590), .ZN(n7193) );
  AND2_X1 U10829 ( .A1(n29701), .A2(n5977), .Z(n14511) );
  NOR2_X1 U10833 ( .A1(n16490), .A2(n29940), .ZN(n7363) );
  INV_X1 U10834 ( .I(n11677), .ZN(n9836) );
  NOR2_X1 U10836 ( .A1(n10702), .A2(n7789), .ZN(n8892) );
  INV_X1 U10845 ( .I(n9649), .ZN(n2001) );
  OR2_X1 U10846 ( .A1(n29450), .A2(n28899), .Z(n29380) );
  INV_X1 U10847 ( .I(n29904), .ZN(n29902) );
  AND2_X1 U10849 ( .A1(n10569), .A2(n6938), .Z(n28788) );
  AND2_X1 U10852 ( .A1(n16224), .A2(n16060), .Z(n15521) );
  NOR3_X1 U10853 ( .A1(n14449), .A2(n29310), .A3(n1406), .ZN(n29078) );
  INV_X1 U10863 ( .I(n15293), .ZN(n18461) );
  INV_X1 U10865 ( .I(n35551), .ZN(n11826) );
  NOR2_X1 U10866 ( .A1(n15293), .A2(n20018), .ZN(n12056) );
  INV_X2 U10867 ( .I(n34175), .ZN(n29635) );
  INV_X1 U10868 ( .I(n14438), .ZN(n7295) );
  NAND2_X1 U10870 ( .A1(n20931), .A2(n3986), .ZN(n3951) );
  INV_X1 U10872 ( .I(n30058), .ZN(n3671) );
  INV_X1 U10873 ( .I(n20508), .ZN(n13349) );
  AND2_X1 U10874 ( .A1(n30042), .A2(n30041), .Z(n29150) );
  AND2_X1 U10875 ( .A1(n2216), .A2(n29957), .Z(n11830) );
  OR2_X1 U10876 ( .A1(n39828), .A2(n20102), .Z(n29173) );
  NOR2_X1 U10877 ( .A1(n28882), .A2(n21023), .ZN(n17681) );
  NOR2_X1 U10878 ( .A1(n971), .A2(n39745), .ZN(n9049) );
  OR2_X1 U10882 ( .A1(n30047), .A2(n16217), .Z(n14664) );
  INV_X1 U10883 ( .I(n29347), .ZN(n14178) );
  AND2_X1 U10884 ( .A1(n15651), .A2(n5414), .Z(n18962) );
  CLKBUF_X2 U10886 ( .I(n29907), .Z(n19878) );
  INV_X4 U10887 ( .I(n29185), .ZN(n1400) );
  NOR2_X1 U10894 ( .A1(n21187), .A2(n29862), .ZN(n2216) );
  INV_X2 U10897 ( .I(n19599), .ZN(n29760) );
  CLKBUF_X2 U10902 ( .I(n14405), .Z(n12353) );
  INV_X1 U10915 ( .I(n29049), .ZN(n12574) );
  INV_X1 U10917 ( .I(n29153), .ZN(n5041) );
  INV_X1 U10918 ( .I(n29114), .ZN(n9436) );
  NAND2_X1 U10921 ( .A1(n15006), .A2(n15005), .ZN(n3551) );
  INV_X1 U10922 ( .I(n29026), .ZN(n2914) );
  INV_X1 U10924 ( .I(n38147), .ZN(n6854) );
  INV_X1 U10925 ( .I(n29162), .ZN(n2995) );
  NAND2_X1 U10927 ( .A1(n7384), .A2(n28747), .ZN(n28751) );
  NAND2_X1 U10928 ( .A1(n19957), .A2(n7296), .ZN(n13484) );
  INV_X1 U10936 ( .I(n15271), .ZN(n11347) );
  INV_X1 U10944 ( .I(n28852), .ZN(n28707) );
  INV_X1 U10946 ( .I(n28529), .ZN(n28343) );
  NAND2_X1 U10955 ( .A1(n28522), .A2(n28747), .ZN(n12608) );
  NAND2_X1 U10961 ( .A1(n18473), .A2(n18470), .ZN(n28953) );
  AOI21_X1 U10968 ( .A1(n20314), .A2(n28331), .B(n29474), .ZN(n15007) );
  NAND2_X1 U10972 ( .A1(n28480), .A2(n32575), .ZN(n4665) );
  AND2_X1 U10976 ( .A1(n6405), .A2(n3927), .Z(n8323) );
  INV_X1 U10980 ( .I(n1815), .ZN(n4371) );
  OR2_X1 U11003 ( .A1(n28095), .A2(n19827), .Z(n14049) );
  INV_X1 U11006 ( .I(n28747), .ZN(n4025) );
  NAND2_X1 U11026 ( .A1(n20952), .A2(n28748), .ZN(n20951) );
  AND2_X1 U11032 ( .A1(n6287), .A2(n37204), .Z(n12882) );
  NOR2_X1 U11033 ( .A1(n28289), .A2(n1187), .ZN(n13963) );
  INV_X1 U11035 ( .I(n28455), .ZN(n12883) );
  OR3_X1 U11041 ( .A1(n28720), .A2(n28722), .A3(n38145), .Z(n13593) );
  INV_X1 U11044 ( .I(n28431), .ZN(n16307) );
  AND2_X1 U11057 ( .A1(n28612), .A2(n7454), .Z(n2060) );
  AND2_X1 U11060 ( .A1(n6892), .A2(n12237), .Z(n12238) );
  AND2_X1 U11065 ( .A1(n9878), .A2(n32146), .Z(n28528) );
  NOR2_X1 U11067 ( .A1(n10544), .A2(n10543), .ZN(n13563) );
  INV_X1 U11069 ( .I(n28576), .ZN(n2703) );
  NOR2_X1 U11077 ( .A1(n39355), .A2(n28464), .ZN(n28302) );
  INV_X1 U11081 ( .I(n28535), .ZN(n7869) );
  INV_X1 U11082 ( .I(n15752), .ZN(n5399) );
  NOR2_X1 U11092 ( .A1(n1190), .A2(n30894), .ZN(n17542) );
  NAND2_X1 U11095 ( .A1(n13508), .A2(n28408), .ZN(n20878) );
  AND2_X1 U11099 ( .A1(n28551), .A2(n28659), .Z(n14652) );
  AND2_X1 U11100 ( .A1(n10907), .A2(n18871), .Z(n10857) );
  NAND2_X1 U11102 ( .A1(n3903), .A2(n28569), .ZN(n28571) );
  OR2_X1 U11105 ( .A1(n28606), .A2(n8349), .Z(n12045) );
  NOR2_X1 U11106 ( .A1(n28391), .A2(n28486), .ZN(n12343) );
  NAND2_X1 U11107 ( .A1(n28313), .A2(n19844), .ZN(n28209) );
  AND2_X1 U11110 ( .A1(n28532), .A2(n36796), .Z(n13894) );
  AND2_X1 U11113 ( .A1(n28759), .A2(n2022), .Z(n13237) );
  NOR2_X1 U11114 ( .A1(n7251), .A2(n31554), .ZN(n5343) );
  INV_X1 U11118 ( .I(n28515), .ZN(n9638) );
  INV_X1 U11120 ( .I(n1193), .ZN(n5152) );
  AND2_X1 U11124 ( .A1(n28433), .A2(n28434), .Z(n8322) );
  AND2_X1 U11126 ( .A1(n28681), .A2(n15473), .Z(n14677) );
  INV_X1 U11128 ( .I(n13601), .ZN(n6017) );
  OAI21_X1 U11129 ( .A1(n38998), .A2(n36623), .B(n5028), .ZN(n3191) );
  NOR2_X1 U11130 ( .A1(n28606), .A2(n2639), .ZN(n10757) );
  NOR2_X1 U11134 ( .A1(n20199), .A2(n20198), .ZN(n20197) );
  NAND2_X1 U11136 ( .A1(n13133), .A2(n496), .ZN(n8714) );
  OR2_X1 U11140 ( .A1(n8349), .A2(n36827), .Z(n14339) );
  AND2_X1 U11141 ( .A1(n18369), .A2(n28717), .Z(n4428) );
  AND2_X1 U11144 ( .A1(n28772), .A2(n17771), .Z(n28773) );
  NOR2_X1 U11147 ( .A1(n31597), .A2(n14760), .ZN(n28635) );
  INV_X1 U11151 ( .I(n28444), .ZN(n14003) );
  INV_X1 U11153 ( .I(n1192), .ZN(n11128) );
  NAND3_X1 U11156 ( .A1(n28424), .A2(n17818), .A3(n28423), .ZN(n9405) );
  OAI21_X1 U11165 ( .A1(n1206), .A2(n3231), .B(n3230), .ZN(n4028) );
  NOR2_X1 U11178 ( .A1(n18020), .A2(n17447), .ZN(n17057) );
  NAND2_X1 U11195 ( .A1(n11743), .A2(n37623), .ZN(n11742) );
  AND4_X1 U11200 ( .A1(n28347), .A2(n28346), .A3(n28345), .A4(n28344), .Z(
        n28348) );
  AND3_X1 U11204 ( .A1(n20019), .A2(n20020), .A3(n28104), .Z(n14596) );
  INV_X1 U11205 ( .I(n11717), .ZN(n12061) );
  INV_X1 U11208 ( .I(n10167), .ZN(n3534) );
  NAND2_X1 U11216 ( .A1(n1198), .A2(n27892), .ZN(n13755) );
  NAND2_X1 U11223 ( .A1(n28053), .A2(n18392), .ZN(n13847) );
  NAND2_X1 U11235 ( .A1(n8290), .A2(n1073), .ZN(n8289) );
  NAND2_X1 U11243 ( .A1(n1445), .A2(n981), .ZN(n17856) );
  INV_X1 U11245 ( .I(n8819), .ZN(n28243) );
  NAND2_X1 U11252 ( .A1(n28022), .A2(n27951), .ZN(n11705) );
  NAND2_X1 U11257 ( .A1(n27948), .A2(n28022), .ZN(n19039) );
  NAND2_X1 U11259 ( .A1(n11024), .A2(n28260), .ZN(n10150) );
  OAI21_X1 U11260 ( .A1(n7719), .A2(n984), .B(n7718), .ZN(n28058) );
  OAI21_X1 U11262 ( .A1(n4767), .A2(n14389), .B(n4766), .ZN(n28185) );
  NAND2_X1 U11268 ( .A1(n18530), .A2(n19743), .ZN(n18529) );
  NOR2_X1 U11272 ( .A1(n27963), .A2(n14404), .ZN(n21318) );
  NAND2_X1 U11276 ( .A1(n28259), .A2(n28258), .ZN(n9990) );
  NOR2_X1 U11277 ( .A1(n16115), .A2(n580), .ZN(n6693) );
  NAND2_X1 U11278 ( .A1(n5939), .A2(n28045), .ZN(n4889) );
  INV_X1 U11293 ( .I(n13984), .ZN(n10536) );
  AND2_X1 U11296 ( .A1(n1202), .A2(n16115), .Z(n6245) );
  OAI21_X1 U11299 ( .A1(n8801), .A2(n18061), .B(n27998), .ZN(n4788) );
  INV_X1 U11307 ( .I(n6777), .ZN(n3198) );
  INV_X1 U11311 ( .I(n28223), .ZN(n28227) );
  INV_X1 U11312 ( .I(n15695), .ZN(n15693) );
  NAND2_X1 U11313 ( .A1(n8291), .A2(n17032), .ZN(n8290) );
  AOI21_X1 U11314 ( .A1(n33980), .A2(n13457), .B(n36844), .ZN(n3067) );
  OAI21_X1 U11316 ( .A1(n16461), .A2(n878), .B(n4507), .ZN(n4506) );
  NOR2_X1 U11319 ( .A1(n33957), .A2(n28283), .ZN(n13993) );
  INV_X1 U11330 ( .I(n28235), .ZN(n3832) );
  INV_X1 U11335 ( .I(n28285), .ZN(n6374) );
  OR2_X1 U11341 ( .A1(n1211), .A2(n28089), .Z(n6118) );
  NAND2_X1 U11351 ( .A1(n2302), .A2(n17314), .ZN(n27888) );
  OR2_X1 U11353 ( .A1(n1209), .A2(n882), .Z(n27911) );
  INV_X1 U11354 ( .I(n11408), .ZN(n8351) );
  AND3_X1 U11359 ( .A1(n33656), .A2(n37783), .A3(n288), .Z(n6115) );
  OAI21_X1 U11361 ( .A1(n27772), .A2(n36877), .B(n30846), .ZN(n10825) );
  NOR2_X1 U11363 ( .A1(n5940), .A2(n6990), .ZN(n5939) );
  OR2_X1 U11369 ( .A1(n18841), .A2(n16065), .Z(n4825) );
  NAND2_X1 U11371 ( .A1(n28257), .A2(n3989), .ZN(n3164) );
  NAND2_X1 U11375 ( .A1(n12623), .A2(n28238), .ZN(n2983) );
  AND2_X1 U11386 ( .A1(n759), .A2(n28205), .Z(n14791) );
  INV_X1 U11391 ( .I(n27901), .ZN(n4507) );
  INV_X1 U11394 ( .I(n28282), .ZN(n12807) );
  INV_X1 U11396 ( .I(n10009), .ZN(n14829) );
  INV_X2 U11400 ( .I(n12298), .ZN(n27910) );
  OR2_X1 U11405 ( .A1(n27995), .A2(n16461), .Z(n4502) );
  OR2_X1 U11406 ( .A1(n5266), .A2(n20053), .Z(n20993) );
  AND2_X1 U11409 ( .A1(n19667), .A2(n28137), .Z(n16987) );
  NOR2_X1 U11411 ( .A1(n36854), .A2(n11283), .ZN(n2613) );
  INV_X1 U11412 ( .I(n12663), .ZN(n19525) );
  BUF_X2 U11413 ( .I(n19855), .Z(n6643) );
  NAND2_X1 U11414 ( .A1(n39488), .A2(n28237), .ZN(n2982) );
  NOR2_X1 U11417 ( .A1(n16115), .A2(n39571), .ZN(n15048) );
  INV_X2 U11418 ( .I(n17177), .ZN(n1445) );
  INV_X1 U11419 ( .I(n28127), .ZN(n28124) );
  INV_X2 U11424 ( .I(n9791), .ZN(n15925) );
  CLKBUF_X2 U11425 ( .I(n28132), .Z(n19946) );
  BUF_X2 U11428 ( .I(n28127), .Z(n11891) );
  INV_X4 U11429 ( .I(n28236), .ZN(n1453) );
  INV_X1 U11430 ( .I(n27675), .ZN(n6471) );
  INV_X1 U11432 ( .I(n14977), .ZN(n3499) );
  INV_X1 U11433 ( .I(n27732), .ZN(n27733) );
  OAI21_X1 U11441 ( .A1(n13291), .A2(n13290), .B(n27523), .ZN(n12240) );
  INV_X1 U11451 ( .I(n13293), .ZN(n13290) );
  NAND2_X2 U11453 ( .A1(n12415), .A2(n26967), .ZN(n12556) );
  NAND2_X1 U11455 ( .A1(n27466), .A2(n19877), .ZN(n17686) );
  AND2_X1 U11459 ( .A1(n27346), .A2(n27345), .Z(n6689) );
  NOR2_X1 U11463 ( .A1(n10576), .A2(n10575), .ZN(n10573) );
  OAI21_X1 U11471 ( .A1(n17524), .A2(n21110), .B(n17523), .ZN(n4419) );
  INV_X1 U11476 ( .I(n26942), .ZN(n10575) );
  INV_X1 U11477 ( .I(n13245), .ZN(n27597) );
  INV_X1 U11481 ( .I(n27178), .ZN(n27860) );
  INV_X1 U11482 ( .I(n10580), .ZN(n10576) );
  INV_X1 U11487 ( .I(n27549), .ZN(n27863) );
  NAND2_X1 U11489 ( .A1(n27199), .A2(n35919), .ZN(n9202) );
  AND3_X1 U11493 ( .A1(n27563), .A2(n27562), .A3(n27561), .Z(n18927) );
  INV_X1 U11497 ( .I(n27501), .ZN(n7910) );
  INV_X1 U11499 ( .I(n27632), .ZN(n12970) );
  INV_X1 U11501 ( .I(n27509), .ZN(n15245) );
  INV_X2 U11502 ( .I(n27541), .ZN(n1466) );
  INV_X2 U11505 ( .I(n27755), .ZN(n1467) );
  NAND2_X1 U11508 ( .A1(n30981), .A2(n27368), .ZN(n13462) );
  NAND2_X1 U11514 ( .A1(n27351), .A2(n11682), .ZN(n8168) );
  INV_X1 U11516 ( .I(n10177), .ZN(n10176) );
  NAND2_X1 U11517 ( .A1(n27559), .A2(n8252), .ZN(n27563) );
  NAND3_X1 U11531 ( .A1(n20143), .A2(n20145), .A3(n27288), .ZN(n12446) );
  NAND2_X1 U11534 ( .A1(n8931), .A2(n36159), .ZN(n7312) );
  NAND2_X1 U11536 ( .A1(n27351), .A2(n8988), .ZN(n27051) );
  AND3_X1 U11540 ( .A1(n27428), .A2(n4964), .A3(n10461), .Z(n9452) );
  NAND2_X1 U11557 ( .A1(n27366), .A2(n9310), .ZN(n5774) );
  OR3_X1 U11563 ( .A1(n39711), .A2(n35904), .A3(n1084), .Z(n14116) );
  NOR2_X1 U11566 ( .A1(n5101), .A2(n6534), .ZN(n7894) );
  NOR2_X1 U11578 ( .A1(n2259), .A2(n5559), .ZN(n2258) );
  OAI21_X1 U11579 ( .A1(n38305), .A2(n27197), .B(n19455), .ZN(n16127) );
  NAND3_X1 U11580 ( .A1(n27412), .A2(n36200), .A3(n997), .ZN(n20203) );
  OR2_X1 U11588 ( .A1(n18562), .A2(n12018), .Z(n12017) );
  NAND2_X1 U11597 ( .A1(n27430), .A2(n10051), .ZN(n10755) );
  NAND2_X1 U11616 ( .A1(n9512), .A2(n27009), .ZN(n10574) );
  NAND2_X1 U11621 ( .A1(n27220), .A2(n39546), .ZN(n6192) );
  OR2_X1 U11627 ( .A1(n27289), .A2(n1223), .Z(n14682) );
  NAND2_X1 U11628 ( .A1(n27020), .A2(n11140), .ZN(n16919) );
  NAND2_X1 U11633 ( .A1(n1080), .A2(n17662), .ZN(n17465) );
  NOR2_X1 U11636 ( .A1(n27248), .A2(n6972), .ZN(n11853) );
  NAND2_X1 U11637 ( .A1(n991), .A2(n3531), .ZN(n8932) );
  NAND2_X1 U11643 ( .A1(n26428), .A2(n35299), .ZN(n9680) );
  NAND2_X1 U11652 ( .A1(n994), .A2(n35258), .ZN(n1798) );
  AND2_X1 U11654 ( .A1(n27484), .A2(n1218), .Z(n11042) );
  NAND2_X1 U11658 ( .A1(n18549), .A2(n34562), .ZN(n12018) );
  NAND2_X1 U11664 ( .A1(n11039), .A2(n39296), .ZN(n7227) );
  AND2_X1 U11665 ( .A1(n27387), .A2(n6908), .Z(n20870) );
  NAND2_X1 U11669 ( .A1(n18669), .A2(n14881), .ZN(n18668) );
  AND2_X1 U11674 ( .A1(n27385), .A2(n34562), .Z(n5219) );
  AND2_X1 U11682 ( .A1(n39671), .A2(n20740), .Z(n14482) );
  NAND2_X1 U11693 ( .A1(n27298), .A2(n8137), .ZN(n4038) );
  INV_X1 U11696 ( .I(n5630), .ZN(n2006) );
  INV_X1 U11700 ( .I(n27128), .ZN(n6416) );
  NOR2_X1 U11702 ( .A1(n31672), .A2(n27269), .ZN(n3466) );
  NAND2_X1 U11706 ( .A1(n27383), .A2(n27064), .ZN(n12022) );
  NOR2_X1 U11720 ( .A1(n12685), .A2(n27417), .ZN(n7175) );
  INV_X1 U11722 ( .I(n20871), .ZN(n2846) );
  AOI21_X1 U11723 ( .A1(n31672), .A2(n27267), .B(n27372), .ZN(n15748) );
  NAND2_X1 U11739 ( .A1(n26612), .A2(n14496), .ZN(n17467) );
  NAND2_X1 U11740 ( .A1(n26037), .A2(n10890), .ZN(n12510) );
  NAND2_X1 U11742 ( .A1(n20797), .A2(n10187), .ZN(n7912) );
  INV_X2 U11743 ( .I(n9144), .ZN(n26870) );
  NAND2_X1 U11762 ( .A1(n38120), .A2(n26515), .ZN(n4489) );
  NAND2_X1 U11780 ( .A1(n20462), .A2(n21202), .ZN(n10203) );
  INV_X1 U11784 ( .I(n8311), .ZN(n26684) );
  NAND2_X1 U11792 ( .A1(n26731), .A2(n17712), .ZN(n9075) );
  NAND2_X1 U11817 ( .A1(n26697), .A2(n26269), .ZN(n4937) );
  OR2_X1 U11824 ( .A1(n7742), .A2(n4218), .Z(n20912) );
  NOR2_X1 U11825 ( .A1(n14825), .A2(n17047), .ZN(n13159) );
  NOR2_X1 U11833 ( .A1(n3368), .A2(n1229), .ZN(n20549) );
  OR2_X1 U11836 ( .A1(n16773), .A2(n3388), .Z(n26138) );
  NAND2_X1 U11838 ( .A1(n4486), .A2(n11334), .ZN(n4485) );
  NAND2_X1 U11840 ( .A1(n26926), .A2(n26470), .ZN(n6503) );
  NAND2_X1 U11843 ( .A1(n26283), .A2(n19353), .ZN(n13252) );
  NAND2_X1 U11846 ( .A1(n14382), .A2(n860), .ZN(n8746) );
  NOR2_X1 U11848 ( .A1(n26299), .A2(n26763), .ZN(n7320) );
  NAND2_X1 U11856 ( .A1(n17655), .A2(n13110), .ZN(n17823) );
  NAND2_X1 U11857 ( .A1(n17466), .A2(n36392), .ZN(n11388) );
  NOR2_X1 U11859 ( .A1(n15124), .A2(n13181), .ZN(n4173) );
  NAND2_X1 U11864 ( .A1(n19206), .A2(n19425), .ZN(n26717) );
  INV_X2 U11866 ( .I(n19762), .ZN(n26826) );
  OAI21_X1 U11868 ( .A1(n26842), .A2(n34004), .B(n9650), .ZN(n21181) );
  OR2_X1 U11871 ( .A1(n26671), .A2(n26672), .Z(n14583) );
  NAND2_X1 U11879 ( .A1(n26734), .A2(n9188), .ZN(n9763) );
  NAND2_X1 U11880 ( .A1(n10913), .A2(n26978), .ZN(n5438) );
  INV_X1 U11883 ( .I(n18792), .ZN(n4887) );
  AND2_X1 U11886 ( .A1(n26686), .A2(n26979), .Z(n17098) );
  NOR2_X1 U11894 ( .A1(n26819), .A2(n37104), .ZN(n13948) );
  NOR2_X1 U11898 ( .A1(n13110), .A2(n26993), .ZN(n4656) );
  NOR2_X1 U11899 ( .A1(n38491), .A2(n19332), .ZN(n18706) );
  OR2_X1 U11914 ( .A1(n33726), .A2(n3328), .Z(n26813) );
  NAND2_X1 U11915 ( .A1(n5869), .A2(n26932), .ZN(n16633) );
  AND2_X1 U11923 ( .A1(n13758), .A2(n3134), .Z(n3135) );
  NOR2_X1 U11924 ( .A1(n3574), .A2(n1008), .ZN(n3573) );
  OAI22_X1 U11925 ( .A1(n26979), .A2(n26978), .B1(n17097), .B2(n17252), .ZN(
        n26981) );
  OR3_X1 U11929 ( .A1(n26901), .A2(n10231), .A3(n19821), .Z(n26902) );
  NOR2_X1 U11931 ( .A1(n26930), .A2(n19222), .ZN(n7523) );
  INV_X1 U11932 ( .I(n14347), .ZN(n16970) );
  INV_X1 U11935 ( .I(n26926), .ZN(n26928) );
  NOR2_X1 U11938 ( .A1(n1232), .A2(n19371), .ZN(n8989) );
  NOR2_X1 U11939 ( .A1(n2966), .A2(n19338), .ZN(n2965) );
  INV_X1 U11940 ( .I(n13777), .ZN(n4486) );
  INV_X1 U11941 ( .I(n33561), .ZN(n19045) );
  OR2_X1 U11944 ( .A1(n26724), .A2(n14355), .Z(n26725) );
  AND2_X1 U11956 ( .A1(n6190), .A2(n10440), .Z(n8010) );
  NOR2_X1 U11960 ( .A1(n26708), .A2(n17034), .ZN(n4946) );
  INV_X1 U11974 ( .I(n13131), .ZN(n26346) );
  INV_X1 U11975 ( .I(n26309), .ZN(n13928) );
  INV_X1 U11977 ( .I(n34009), .ZN(n19882) );
  INV_X1 U11979 ( .I(n26348), .ZN(n7474) );
  INV_X1 U11986 ( .I(n26154), .ZN(n7571) );
  INV_X1 U11987 ( .I(n26201), .ZN(n3802) );
  INV_X1 U11991 ( .I(n9001), .ZN(n6413) );
  INV_X1 U11993 ( .I(n26434), .ZN(n3639) );
  INV_X1 U12000 ( .I(n3219), .ZN(n3218) );
  INV_X1 U12002 ( .I(n17757), .ZN(n26291) );
  NAND2_X1 U12007 ( .A1(n14546), .A2(n26333), .ZN(n12859) );
  INV_X1 U12010 ( .I(n7481), .ZN(n2178) );
  INV_X1 U12013 ( .I(n5241), .ZN(n5691) );
  INV_X1 U12017 ( .I(n36522), .ZN(n26550) );
  INV_X1 U12019 ( .I(n26514), .ZN(n12915) );
  OR2_X1 U12033 ( .A1(n10724), .A2(n25989), .Z(n20336) );
  NAND2_X1 U12039 ( .A1(n4293), .A2(n37502), .ZN(n4292) );
  NOR2_X1 U12041 ( .A1(n33440), .A2(n26001), .ZN(n9375) );
  OAI21_X1 U12048 ( .A1(n424), .A2(n927), .B(n5162), .ZN(n5161) );
  NAND2_X1 U12052 ( .A1(n18958), .A2(n7544), .ZN(n12490) );
  NAND2_X1 U12060 ( .A1(n8710), .A2(n26027), .ZN(n8709) );
  NOR2_X1 U12061 ( .A1(n26214), .A2(n5908), .ZN(n17125) );
  NAND2_X1 U12062 ( .A1(n25958), .A2(n25959), .ZN(n2125) );
  INV_X1 U12070 ( .I(n14157), .ZN(n26238) );
  AND2_X1 U12071 ( .A1(n26187), .A2(n14375), .Z(n16878) );
  INV_X1 U12073 ( .I(n26190), .ZN(n3333) );
  NAND2_X1 U12077 ( .A1(n17035), .A2(n25970), .ZN(n9811) );
  AND2_X1 U12078 ( .A1(n25770), .A2(n25941), .Z(n14685) );
  NAND2_X1 U12084 ( .A1(n8898), .A2(n26045), .ZN(n20965) );
  NAND2_X1 U12091 ( .A1(n6883), .A2(n11904), .ZN(n1850) );
  NAND2_X1 U12092 ( .A1(n1239), .A2(n25744), .ZN(n7415) );
  OAI21_X1 U12094 ( .A1(n4163), .A2(n3517), .B(n5356), .ZN(n3516) );
  NAND2_X1 U12097 ( .A1(n37306), .A2(n5886), .ZN(n5883) );
  AND3_X1 U12101 ( .A1(n19259), .A2(n2830), .A3(n1021), .Z(n4794) );
  AND2_X1 U12105 ( .A1(n26010), .A2(n26012), .Z(n3555) );
  INV_X1 U12107 ( .I(n26131), .ZN(n14146) );
  AND2_X1 U12108 ( .A1(n14133), .A2(n14131), .Z(n25938) );
  OAI22_X1 U12111 ( .A1(n7369), .A2(n31205), .B1(n1014), .B2(n26024), .ZN(
        n6400) );
  INV_X1 U12113 ( .I(n6180), .ZN(n25875) );
  NAND2_X1 U12118 ( .A1(n18037), .A2(n25961), .ZN(n13164) );
  NAND2_X1 U12124 ( .A1(n17439), .A2(n840), .ZN(n5683) );
  OAI21_X1 U12127 ( .A1(n25982), .A2(n25981), .B(n39375), .ZN(n25983) );
  OAI21_X1 U12133 ( .A1(n4190), .A2(n5098), .B(n10834), .ZN(n11904) );
  AOI21_X1 U12135 ( .A1(n26111), .A2(n14228), .B(n951), .ZN(n6589) );
  AOI21_X1 U12139 ( .A1(n926), .A2(n26018), .B(n1020), .ZN(n11763) );
  NAND2_X1 U12142 ( .A1(n950), .A2(n4699), .ZN(n12522) );
  NAND2_X1 U12146 ( .A1(n11762), .A2(n34898), .ZN(n13586) );
  AND3_X1 U12147 ( .A1(n32690), .A2(n34961), .A3(n38835), .Z(n4884) );
  NAND2_X1 U12153 ( .A1(n25915), .A2(n25978), .ZN(n16977) );
  NOR2_X1 U12156 ( .A1(n25852), .A2(n13391), .ZN(n13067) );
  NAND2_X1 U12160 ( .A1(n25927), .A2(n5356), .ZN(n18958) );
  NAND2_X1 U12165 ( .A1(n7370), .A2(n26024), .ZN(n7369) );
  INV_X1 U12167 ( .I(n17008), .ZN(n20530) );
  AOI21_X1 U12170 ( .A1(n26109), .A2(n14228), .B(n1019), .ZN(n17035) );
  NAND2_X1 U12171 ( .A1(n33293), .A2(n36922), .ZN(n4832) );
  OR2_X1 U12176 ( .A1(n25852), .A2(n31523), .Z(n2946) );
  INV_X1 U12181 ( .I(n26110), .ZN(n11945) );
  AND3_X1 U12183 ( .A1(n1240), .A2(n26330), .A3(n931), .Z(n14407) );
  CLKBUF_X2 U12191 ( .I(n26328), .Z(n19574) );
  NAND2_X1 U12198 ( .A1(n26130), .A2(n9916), .ZN(n7370) );
  INV_X1 U12203 ( .I(n26113), .ZN(n8393) );
  AND2_X1 U12207 ( .A1(n18162), .A2(n17180), .Z(n25783) );
  INV_X1 U12208 ( .I(n26024), .ZN(n20769) );
  NAND2_X1 U12215 ( .A1(n15575), .A2(n17624), .ZN(n10234) );
  NOR3_X1 U12216 ( .A1(n26108), .A2(n1017), .A3(n38760), .ZN(n10137) );
  NOR2_X1 U12218 ( .A1(n31205), .A2(n25813), .ZN(n7699) );
  NOR2_X1 U12220 ( .A1(n4385), .A2(n2625), .ZN(n8376) );
  NAND2_X1 U12224 ( .A1(n5753), .A2(n33440), .ZN(n7134) );
  INV_X1 U12235 ( .I(n36546), .ZN(n6221) );
  AND2_X1 U12246 ( .A1(n25836), .A2(n33997), .Z(n14694) );
  NAND2_X1 U12250 ( .A1(n25567), .A2(n19438), .ZN(n16569) );
  NOR2_X1 U12257 ( .A1(n4048), .A2(n8906), .ZN(n8905) );
  NAND2_X1 U12269 ( .A1(n13195), .A2(n19367), .ZN(n13194) );
  INV_X1 U12274 ( .I(n17305), .ZN(n4433) );
  NOR2_X1 U12275 ( .A1(n7853), .A2(n5519), .ZN(n5711) );
  NAND2_X1 U12286 ( .A1(n20876), .A2(n19237), .ZN(n20875) );
  NAND2_X1 U12296 ( .A1(n6762), .A2(n6763), .ZN(n1932) );
  INV_X1 U12298 ( .I(n38825), .ZN(n25904) );
  CLKBUF_X2 U12300 ( .I(n26124), .Z(n9682) );
  INV_X1 U12307 ( .I(n25479), .ZN(n8978) );
  AND3_X1 U12308 ( .A1(n25719), .A2(n18519), .A3(n18831), .Z(n8689) );
  NOR2_X1 U12310 ( .A1(n7235), .A2(n25721), .ZN(n7234) );
  AND2_X1 U12313 ( .A1(n39289), .A2(n953), .Z(n8878) );
  OAI21_X1 U12318 ( .A1(n25437), .A2(n39389), .B(n39599), .ZN(n25438) );
  OAI21_X1 U12323 ( .A1(n25427), .A2(n19302), .B(n34150), .ZN(n25714) );
  OAI21_X1 U12337 ( .A1(n12478), .A2(n33950), .B(n20648), .ZN(n11333) );
  OAI21_X1 U12340 ( .A1(n25698), .A2(n17774), .B(n11641), .ZN(n16229) );
  AND2_X1 U12343 ( .A1(n17303), .A2(n25389), .Z(n4988) );
  NAND2_X1 U12344 ( .A1(n1022), .A2(n36019), .ZN(n18694) );
  NAND2_X1 U12345 ( .A1(n38178), .A2(n8033), .ZN(n8032) );
  AND2_X1 U12349 ( .A1(n25719), .A2(n25557), .Z(n17282) );
  NAND2_X1 U12350 ( .A1(n14056), .A2(n34464), .ZN(n14192) );
  NAND2_X1 U12352 ( .A1(n17450), .A2(n18831), .ZN(n13195) );
  NOR2_X1 U12356 ( .A1(n24894), .A2(n25449), .ZN(n8122) );
  NOR2_X1 U12365 ( .A1(n32101), .A2(n7802), .ZN(n18988) );
  AND2_X1 U12368 ( .A1(n38359), .A2(n3736), .Z(n3735) );
  NAND2_X1 U12371 ( .A1(n14947), .A2(n11874), .ZN(n5901) );
  NAND2_X1 U12373 ( .A1(n25577), .A2(n25660), .ZN(n11806) );
  OR2_X1 U12374 ( .A1(n1109), .A2(n25660), .Z(n13826) );
  NAND2_X1 U12376 ( .A1(n25012), .A2(n25337), .ZN(n6939) );
  NOR2_X1 U12378 ( .A1(n32419), .A2(n4048), .ZN(n4047) );
  NAND2_X1 U12380 ( .A1(n33826), .A2(n25425), .ZN(n4791) );
  NAND2_X1 U12386 ( .A1(n4755), .A2(n5798), .ZN(n4754) );
  OAI21_X1 U12389 ( .A1(n25448), .A2(n38782), .B(n17304), .ZN(n4989) );
  NAND2_X1 U12390 ( .A1(n18734), .A2(n1256), .ZN(n7878) );
  INV_X1 U12397 ( .I(n25548), .ZN(n12417) );
  OR2_X1 U12398 ( .A1(n18909), .A2(n21254), .Z(n4976) );
  AND3_X1 U12409 ( .A1(n25689), .A2(n19548), .A3(n31557), .Z(n25506) );
  NAND3_X1 U12410 ( .A1(n25681), .A2(n25680), .A3(n25679), .ZN(n13589) );
  INV_X1 U12413 ( .I(n9441), .ZN(n9241) );
  AND3_X1 U12414 ( .A1(n25540), .A2(n5042), .A3(n25513), .Z(n14613) );
  AND2_X1 U12425 ( .A1(n12500), .A2(n7866), .Z(n12768) );
  AND2_X1 U12432 ( .A1(n541), .A2(n319), .Z(n14666) );
  OR2_X1 U12433 ( .A1(n20052), .A2(n25477), .Z(n11924) );
  OR2_X1 U12434 ( .A1(n33130), .A2(n14460), .Z(n14490) );
  AND2_X1 U12444 ( .A1(n25355), .A2(n24896), .Z(n4674) );
  NOR2_X1 U12445 ( .A1(n14472), .A2(n24963), .ZN(n10973) );
  OAI21_X1 U12446 ( .A1(n14475), .A2(n15180), .B(n25401), .ZN(n20859) );
  NAND2_X1 U12449 ( .A1(n17281), .A2(n18519), .ZN(n7238) );
  OR2_X1 U12452 ( .A1(n19701), .A2(n16933), .Z(n25333) );
  NAND2_X1 U12455 ( .A1(n17183), .A2(n14602), .ZN(n11063) );
  INV_X1 U12458 ( .I(n19636), .ZN(n25385) );
  OR2_X1 U12460 ( .A1(n25670), .A2(n18164), .Z(n11647) );
  NAND2_X1 U12461 ( .A1(n25408), .A2(n25606), .ZN(n4647) );
  INV_X1 U12465 ( .I(n25725), .ZN(n25633) );
  AND2_X1 U12472 ( .A1(n25412), .A2(n25307), .Z(n16911) );
  AND2_X1 U12476 ( .A1(n8304), .A2(n37926), .Z(n14475) );
  NAND3_X1 U12486 ( .A1(n8764), .A2(n5501), .A3(n7990), .ZN(n5500) );
  INV_X1 U12492 ( .I(n25022), .ZN(n8764) );
  OAI21_X1 U12496 ( .A1(n9183), .A2(n9182), .B(n7967), .ZN(n9181) );
  INV_X1 U12500 ( .I(n9177), .ZN(n5501) );
  INV_X1 U12505 ( .I(n39541), .ZN(n9564) );
  INV_X1 U12506 ( .I(n16819), .ZN(n16420) );
  INV_X1 U12508 ( .I(n6759), .ZN(n8447) );
  INV_X1 U12509 ( .I(n7968), .ZN(n7966) );
  INV_X1 U12511 ( .I(n17904), .ZN(n9182) );
  INV_X1 U12518 ( .I(n25127), .ZN(n17445) );
  INV_X1 U12519 ( .I(n18211), .ZN(n6896) );
  INV_X2 U12521 ( .I(n18395), .ZN(n1553) );
  INV_X1 U12523 ( .I(n16581), .ZN(n9438) );
  NAND2_X1 U12526 ( .A1(n1118), .A2(n2747), .ZN(n16820) );
  INV_X1 U12527 ( .I(n16751), .ZN(n8608) );
  NOR2_X1 U12531 ( .A1(n10988), .A2(n10648), .ZN(n2847) );
  INV_X1 U12533 ( .I(n15945), .ZN(n8607) );
  INV_X1 U12534 ( .I(n4063), .ZN(n4062) );
  INV_X1 U12546 ( .I(n9528), .ZN(n17100) );
  NAND2_X1 U12548 ( .A1(n13582), .A2(n13581), .ZN(n14534) );
  INV_X1 U12549 ( .I(n24813), .ZN(n9183) );
  NAND2_X1 U12564 ( .A1(n36955), .A2(n3750), .ZN(n3749) );
  NAND2_X1 U12567 ( .A1(n1907), .A2(n19279), .ZN(n1906) );
  NOR2_X1 U12569 ( .A1(n15527), .A2(n5933), .ZN(n15526) );
  OAI21_X1 U12570 ( .A1(n10114), .A2(n9849), .B(n24735), .ZN(n4688) );
  INV_X1 U12571 ( .I(n7969), .ZN(n7972) );
  INV_X1 U12572 ( .I(n24540), .ZN(n16750) );
  NAND2_X1 U12587 ( .A1(n24755), .A2(n19339), .ZN(n17962) );
  NAND2_X1 U12592 ( .A1(n7242), .A2(n24691), .ZN(n7241) );
  NAND2_X1 U12594 ( .A1(n24733), .A2(n16815), .ZN(n3630) );
  NAND2_X1 U12598 ( .A1(n13553), .A2(n13554), .ZN(n12363) );
  NAND2_X1 U12604 ( .A1(n8428), .A2(n8426), .ZN(n11610) );
  NOR2_X1 U12609 ( .A1(n2634), .A2(n1029), .ZN(n20926) );
  NOR2_X1 U12612 ( .A1(n6038), .A2(n36186), .ZN(n6037) );
  NAND2_X1 U12613 ( .A1(n14167), .A2(n24820), .ZN(n4349) );
  INV_X1 U12615 ( .I(n24704), .ZN(n2697) );
  INV_X1 U12616 ( .I(n24494), .ZN(n13214) );
  NOR2_X1 U12623 ( .A1(n31722), .A2(n18508), .ZN(n13628) );
  NAND2_X1 U12632 ( .A1(n35250), .A2(n14211), .ZN(n24842) );
  INV_X1 U12639 ( .I(n24581), .ZN(n16871) );
  NAND2_X1 U12651 ( .A1(n4008), .A2(n24764), .ZN(n10353) );
  INV_X1 U12652 ( .I(n24602), .ZN(n3374) );
  INV_X1 U12672 ( .I(n24591), .ZN(n6838) );
  NAND2_X1 U12674 ( .A1(n5934), .A2(n16547), .ZN(n5933) );
  INV_X1 U12677 ( .I(n5934), .ZN(n2537) );
  INV_X1 U12681 ( .I(n32831), .ZN(n13518) );
  NAND2_X1 U12686 ( .A1(n24788), .A2(n24787), .ZN(n7065) );
  NAND2_X1 U12697 ( .A1(n17618), .A2(n14276), .ZN(n14275) );
  INV_X1 U12705 ( .I(n24847), .ZN(n11714) );
  NAND2_X1 U12707 ( .A1(n24614), .A2(n24812), .ZN(n12160) );
  NOR2_X1 U12708 ( .A1(n39523), .A2(n38317), .ZN(n2698) );
  NAND2_X1 U12712 ( .A1(n24818), .A2(n17618), .ZN(n4350) );
  NOR2_X1 U12714 ( .A1(n1029), .A2(n19422), .ZN(n20013) );
  INV_X1 U12715 ( .I(n24779), .ZN(n7515) );
  NAND3_X1 U12722 ( .A1(n8842), .A2(n8843), .A3(n8839), .ZN(n18508) );
  NOR2_X1 U12733 ( .A1(n8841), .A2(n8840), .ZN(n8839) );
  OR2_X1 U12734 ( .A1(n19422), .A2(n17101), .Z(n18771) );
  NOR2_X1 U12736 ( .A1(n24811), .A2(n24810), .ZN(n3626) );
  NAND2_X1 U12738 ( .A1(n16238), .A2(n35981), .ZN(n9149) );
  NAND2_X1 U12740 ( .A1(n24874), .A2(n31519), .ZN(n5607) );
  INV_X2 U12744 ( .I(n24878), .ZN(n1570) );
  NAND2_X1 U12756 ( .A1(n20654), .A2(n24222), .ZN(n5712) );
  INV_X1 U12760 ( .I(n15365), .ZN(n8841) );
  INV_X1 U12761 ( .I(n7813), .ZN(n7812) );
  AOI21_X1 U12771 ( .A1(n2400), .A2(n16106), .B(n24330), .ZN(n15497) );
  NOR2_X1 U12779 ( .A1(n11316), .A2(n23797), .ZN(n7624) );
  NAND2_X1 U12795 ( .A1(n24441), .A2(n24440), .ZN(n10784) );
  NAND3_X1 U12799 ( .A1(n16313), .A2(n24086), .A3(n13513), .ZN(n16312) );
  NAND2_X1 U12809 ( .A1(n24297), .A2(n8847), .ZN(n8846) );
  NAND2_X1 U12813 ( .A1(n1031), .A2(n19895), .ZN(n2977) );
  NAND2_X1 U12818 ( .A1(n12665), .A2(n38431), .ZN(n20172) );
  OAI21_X1 U12824 ( .A1(n39818), .A2(n7210), .B(n24121), .ZN(n24125) );
  OAI21_X1 U12827 ( .A1(n35712), .A2(n19653), .B(n4687), .ZN(n5140) );
  INV_X1 U12830 ( .I(n21114), .ZN(n8842) );
  NAND2_X1 U12839 ( .A1(n7773), .A2(n7772), .ZN(n24096) );
  NAND2_X1 U12848 ( .A1(n24355), .A2(n1128), .ZN(n8361) );
  NAND2_X1 U12850 ( .A1(n24141), .A2(n24359), .ZN(n13227) );
  NAND2_X1 U12855 ( .A1(n11134), .A2(n1285), .ZN(n6954) );
  NAND2_X1 U12872 ( .A1(n11261), .A2(n1035), .ZN(n11260) );
  INV_X1 U12880 ( .I(n10421), .ZN(n24627) );
  NAND2_X1 U12882 ( .A1(n8501), .A2(n8500), .ZN(n8499) );
  NAND2_X1 U12890 ( .A1(n3142), .A2(n37047), .ZN(n24377) );
  NAND2_X1 U12898 ( .A1(n12248), .A2(n20839), .ZN(n13808) );
  AND2_X1 U12900 ( .A1(n24303), .A2(n1126), .Z(n24304) );
  INV_X1 U12902 ( .I(n23855), .ZN(n6175) );
  NAND2_X1 U12904 ( .A1(n24400), .A2(n1284), .ZN(n23817) );
  OR2_X1 U12905 ( .A1(n24275), .A2(n24180), .Z(n14654) );
  NAND2_X1 U12907 ( .A1(n12759), .A2(n1276), .ZN(n13692) );
  NOR2_X1 U12909 ( .A1(n20312), .A2(n15320), .ZN(n2268) );
  NAND2_X1 U12912 ( .A1(n24198), .A2(n32891), .ZN(n24199) );
  AND2_X1 U12914 ( .A1(n18466), .A2(n24373), .Z(n24374) );
  NOR2_X1 U12915 ( .A1(n3453), .A2(n30454), .ZN(n14898) );
  NOR2_X1 U12919 ( .A1(n24223), .A2(n24432), .ZN(n5714) );
  NOR2_X1 U12921 ( .A1(n24360), .A2(n39814), .ZN(n15256) );
  NAND2_X1 U12924 ( .A1(n24426), .A2(n38972), .ZN(n18532) );
  NOR2_X1 U12927 ( .A1(n1276), .A2(n5985), .ZN(n12277) );
  OR2_X1 U12929 ( .A1(n24238), .A2(n20313), .Z(n13636) );
  NOR2_X1 U12931 ( .A1(n23855), .A2(n12771), .ZN(n10691) );
  AND2_X1 U12934 ( .A1(n37229), .A2(n21125), .Z(n21124) );
  NAND2_X1 U12935 ( .A1(n19990), .A2(n24461), .ZN(n24460) );
  AOI21_X1 U12939 ( .A1(n1274), .A2(n19653), .B(n13970), .ZN(n9360) );
  AND2_X1 U12946 ( .A1(n14255), .A2(n24119), .Z(n7950) );
  NAND3_X1 U12950 ( .A1(n14718), .A2(n14717), .A3(n24309), .ZN(n13548) );
  OR2_X1 U12952 ( .A1(n24152), .A2(n14491), .Z(n5432) );
  NAND2_X1 U12953 ( .A1(n14699), .A2(n20537), .ZN(n12120) );
  AND2_X1 U12955 ( .A1(n24446), .A2(n24445), .Z(n24447) );
  AND2_X1 U12958 ( .A1(n24296), .A2(n8825), .Z(n9084) );
  AND2_X1 U12961 ( .A1(n23819), .A2(n24116), .Z(n8500) );
  AND2_X1 U12967 ( .A1(n24309), .A2(n24446), .Z(n18141) );
  NAND2_X1 U12969 ( .A1(n24232), .A2(n545), .ZN(n4361) );
  INV_X2 U12976 ( .I(n39467), .ZN(n1587) );
  NAND2_X1 U12978 ( .A1(n24446), .A2(n24445), .ZN(n14717) );
  INV_X1 U12980 ( .I(n5985), .ZN(n18295) );
  OR2_X1 U12984 ( .A1(n24267), .A2(n24445), .Z(n13513) );
  INV_X1 U12985 ( .I(n24207), .ZN(n24218) );
  NOR3_X1 U12989 ( .A1(n94), .A2(n3869), .A3(n370), .ZN(n15205) );
  NAND2_X1 U12997 ( .A1(n1282), .A2(n1288), .ZN(n13040) );
  INV_X2 U12999 ( .I(n13444), .ZN(n19007) );
  NAND2_X1 U13001 ( .A1(n24372), .A2(n24225), .ZN(n16644) );
  NOR2_X1 U13002 ( .A1(n5985), .A2(n19915), .ZN(n20068) );
  NAND2_X1 U13003 ( .A1(n36380), .A2(n1131), .ZN(n16141) );
  OR2_X1 U13007 ( .A1(n800), .A2(n33937), .Z(n14686) );
  NOR2_X1 U13008 ( .A1(n17871), .A2(n14491), .ZN(n7880) );
  NOR2_X1 U13012 ( .A1(n37230), .A2(n20404), .ZN(n7835) );
  INV_X2 U13023 ( .I(n11795), .ZN(n18697) );
  INV_X1 U13026 ( .I(n24245), .ZN(n9519) );
  OR2_X1 U13039 ( .A1(n24445), .A2(n24266), .Z(n14718) );
  NOR2_X1 U13040 ( .A1(n39815), .A2(n24110), .ZN(n10800) );
  INV_X1 U13044 ( .I(n14471), .ZN(n11004) );
  INV_X2 U13051 ( .I(n13540), .ZN(n1609) );
  INV_X1 U13055 ( .I(n23920), .ZN(n5441) );
  INV_X1 U13057 ( .I(n23802), .ZN(n7673) );
  NAND2_X1 U13058 ( .A1(n12820), .A2(n12819), .ZN(n15971) );
  INV_X1 U13061 ( .I(n12798), .ZN(n5005) );
  INV_X1 U13066 ( .I(n24062), .ZN(n20715) );
  INV_X1 U13077 ( .I(n12821), .ZN(n12820) );
  INV_X1 U13080 ( .I(n33322), .ZN(n23805) );
  INV_X1 U13081 ( .I(n38175), .ZN(n23919) );
  NOR2_X1 U13083 ( .A1(n22806), .A2(n10174), .ZN(n10614) );
  INV_X1 U13084 ( .I(n23710), .ZN(n23769) );
  INV_X1 U13085 ( .I(n5841), .ZN(n11116) );
  INV_X1 U13090 ( .I(n15800), .ZN(n5914) );
  INV_X1 U13097 ( .I(n24047), .ZN(n6626) );
  NOR2_X1 U13098 ( .A1(n10205), .A2(n10204), .ZN(n10110) );
  INV_X1 U13100 ( .I(n24053), .ZN(n12842) );
  INV_X1 U13105 ( .I(n23685), .ZN(n23851) );
  NAND2_X1 U13116 ( .A1(n9795), .A2(n9794), .ZN(n18889) );
  INV_X1 U13119 ( .I(n10207), .ZN(n10204) );
  INV_X1 U13120 ( .I(n10208), .ZN(n10205) );
  INV_X2 U13129 ( .I(n14219), .ZN(n1618) );
  NAND2_X1 U13132 ( .A1(n17888), .A2(n23315), .ZN(n16370) );
  NAND2_X1 U13140 ( .A1(n11723), .A2(n23400), .ZN(n18918) );
  INV_X1 U13141 ( .I(n17423), .ZN(n8986) );
  INV_X1 U13152 ( .I(n6561), .ZN(n21046) );
  INV_X1 U13166 ( .I(n23217), .ZN(n2599) );
  NAND2_X1 U13173 ( .A1(n6637), .A2(n6993), .ZN(n6992) );
  NOR2_X1 U13177 ( .A1(n23512), .A2(n23513), .ZN(n7333) );
  AOI21_X1 U13185 ( .A1(n23247), .A2(n14011), .B(n7008), .ZN(n20118) );
  NAND2_X1 U13192 ( .A1(n23471), .A2(n23636), .ZN(n20504) );
  NOR2_X1 U13201 ( .A1(n21051), .A2(n8965), .ZN(n8964) );
  NAND2_X1 U13205 ( .A1(n37209), .A2(n37757), .ZN(n22824) );
  NAND2_X1 U13208 ( .A1(n21156), .A2(n23641), .ZN(n3274) );
  NAND2_X1 U13209 ( .A1(n23575), .A2(n20955), .ZN(n3743) );
  INV_X1 U13210 ( .I(n9796), .ZN(n9795) );
  NAND3_X1 U13214 ( .A1(n8432), .A2(n11186), .A3(n15176), .ZN(n11185) );
  NAND2_X1 U13219 ( .A1(n6217), .A2(n6216), .ZN(n14623) );
  INV_X1 U13221 ( .I(n20100), .ZN(n3383) );
  INV_X1 U13231 ( .I(n17875), .ZN(n7146) );
  OR2_X1 U13232 ( .A1(n23194), .A2(n33349), .Z(n20629) );
  NAND2_X1 U13241 ( .A1(n36829), .A2(n1039), .ZN(n9794) );
  NAND2_X1 U13242 ( .A1(n1295), .A2(n34506), .ZN(n17768) );
  NAND2_X1 U13243 ( .A1(n38248), .A2(n14477), .ZN(n19068) );
  INV_X1 U13251 ( .I(n11186), .ZN(n11187) );
  OAI21_X1 U13253 ( .A1(n17511), .A2(n1139), .B(n20343), .ZN(n12011) );
  NAND2_X1 U13263 ( .A1(n38244), .A2(n1306), .ZN(n2961) );
  NAND2_X1 U13269 ( .A1(n23747), .A2(n39805), .ZN(n23752) );
  AOI21_X1 U13274 ( .A1(n39300), .A2(n10216), .B(n32366), .ZN(n4534) );
  AOI21_X1 U13276 ( .A1(n22987), .A2(n22986), .B(n18762), .ZN(n16033) );
  NOR2_X1 U13283 ( .A1(n31908), .A2(n13414), .ZN(n23555) );
  INV_X1 U13289 ( .I(n23543), .ZN(n2921) );
  INV_X1 U13292 ( .I(n8249), .ZN(n2812) );
  NAND2_X1 U13294 ( .A1(n3716), .A2(n4618), .ZN(n2928) );
  AND2_X1 U13301 ( .A1(n32377), .A2(n13150), .Z(n13560) );
  NAND2_X1 U13303 ( .A1(n9321), .A2(n14477), .ZN(n2683) );
  INV_X1 U13305 ( .I(n23576), .ZN(n6301) );
  OR2_X1 U13312 ( .A1(n35331), .A2(n14235), .Z(n10122) );
  AND2_X1 U13313 ( .A1(n52), .A2(n37431), .Z(n19379) );
  NAND2_X1 U13314 ( .A1(n34012), .A2(n8249), .ZN(n1894) );
  AND2_X1 U13320 ( .A1(n33894), .A2(n7335), .Z(n16575) );
  AND2_X1 U13325 ( .A1(n23580), .A2(n10174), .Z(n23257) );
  AND2_X1 U13327 ( .A1(n34959), .A2(n18866), .Z(n9192) );
  NAND2_X1 U13336 ( .A1(n13095), .A2(n11588), .ZN(n13094) );
  NAND2_X1 U13337 ( .A1(n3717), .A2(n23566), .ZN(n3716) );
  NAND2_X1 U13339 ( .A1(n9340), .A2(n23158), .ZN(n6346) );
  NAND2_X1 U13355 ( .A1(n22369), .A2(n3289), .ZN(n6917) );
  NAND2_X1 U13360 ( .A1(n22858), .A2(n13515), .ZN(n16301) );
  AND2_X1 U13365 ( .A1(n5657), .A2(n38282), .Z(n8459) );
  NAND2_X1 U13366 ( .A1(n16053), .A2(n22894), .ZN(n22896) );
  NOR2_X1 U13375 ( .A1(n15947), .A2(n23120), .ZN(n13095) );
  NAND2_X1 U13381 ( .A1(n9472), .A2(n36453), .ZN(n15345) );
  NAND2_X1 U13383 ( .A1(n11197), .A2(n14725), .ZN(n18856) );
  AND2_X1 U13390 ( .A1(n23042), .A2(n1144), .Z(n9322) );
  NOR2_X1 U13392 ( .A1(n22791), .A2(n23172), .ZN(n20076) );
  AND3_X1 U13397 ( .A1(n11584), .A2(n11582), .A3(n34184), .Z(n11583) );
  AOI21_X1 U13398 ( .A1(n20175), .A2(n20174), .B(n20173), .ZN(n22885) );
  NOR2_X1 U13400 ( .A1(n23046), .A2(n11582), .ZN(n4963) );
  NOR2_X1 U13402 ( .A1(n19082), .A2(n1143), .ZN(n5806) );
  NAND2_X1 U13403 ( .A1(n16957), .A2(n16956), .ZN(n12253) );
  INV_X1 U13408 ( .I(n23044), .ZN(n2726) );
  OR2_X1 U13413 ( .A1(n23005), .A2(n19823), .Z(n5895) );
  NAND2_X1 U13416 ( .A1(n22909), .A2(n22908), .ZN(n21229) );
  NAND2_X1 U13419 ( .A1(n22792), .A2(n22804), .ZN(n8806) );
  NOR2_X1 U13433 ( .A1(n15741), .A2(n32032), .ZN(n15740) );
  NOR2_X1 U13437 ( .A1(n22947), .A2(n23175), .ZN(n15742) );
  INV_X1 U13438 ( .I(n23072), .ZN(n16617) );
  INV_X1 U13440 ( .I(n22947), .ZN(n22960) );
  INV_X1 U13441 ( .I(n22924), .ZN(n5747) );
  INV_X1 U13472 ( .I(n13373), .ZN(n18462) );
  OR2_X2 U13487 ( .A1(n34073), .A2(n16692), .Z(n7130) );
  NAND2_X1 U13498 ( .A1(n22916), .A2(n19870), .ZN(n8143) );
  AOI21_X1 U13505 ( .A1(n33082), .A2(n11658), .B(n34184), .ZN(n16957) );
  AND2_X1 U13507 ( .A1(n38282), .A2(n23198), .Z(n10552) );
  NAND2_X1 U13512 ( .A1(n22850), .A2(n37335), .ZN(n14658) );
  AND2_X1 U13513 ( .A1(n5515), .A2(n14442), .Z(n5786) );
  NOR2_X1 U13516 ( .A1(n640), .A2(n39527), .ZN(n6902) );
  INV_X1 U13517 ( .I(n11704), .ZN(n9660) );
  INV_X1 U13527 ( .I(n23030), .ZN(n5621) );
  NAND2_X1 U13528 ( .A1(n11295), .A2(n23124), .ZN(n22769) );
  INV_X1 U13532 ( .I(n19319), .ZN(n23068) );
  AND2_X1 U13538 ( .A1(n22915), .A2(n23163), .Z(n22916) );
  NOR2_X1 U13540 ( .A1(n36724), .A2(n19535), .ZN(n19246) );
  CLKBUF_X2 U13543 ( .I(n10071), .Z(n9725) );
  INV_X1 U13544 ( .I(n12032), .ZN(n22807) );
  NAND2_X1 U13550 ( .A1(n10634), .A2(n19859), .ZN(n7013) );
  AND2_X1 U13556 ( .A1(n39155), .A2(n18415), .Z(n6385) );
  CLKBUF_X2 U13557 ( .I(n22857), .Z(n7537) );
  INV_X2 U13570 ( .I(n9176), .ZN(n18415) );
  NAND2_X1 U13582 ( .A1(n9334), .A2(n4413), .ZN(n10729) );
  INV_X1 U13583 ( .I(n9334), .ZN(n22587) );
  NAND2_X1 U13584 ( .A1(n10556), .A2(n10555), .ZN(n11255) );
  INV_X1 U13587 ( .I(n15413), .ZN(n12194) );
  INV_X1 U13589 ( .I(n22654), .ZN(n13354) );
  INV_X1 U13590 ( .I(n3969), .ZN(n2236) );
  INV_X1 U13592 ( .I(n22531), .ZN(n22291) );
  INV_X1 U13596 ( .I(n22500), .ZN(n3623) );
  INV_X1 U13599 ( .I(n14309), .ZN(n7593) );
  NAND2_X1 U13603 ( .A1(n38099), .A2(n9483), .ZN(n8549) );
  INV_X2 U13610 ( .I(n22348), .ZN(n1658) );
  INV_X1 U13615 ( .I(n22488), .ZN(n10862) );
  CLKBUF_X2 U13616 ( .I(n19328), .Z(n4819) );
  INV_X1 U13619 ( .I(n9116), .ZN(n9115) );
  INV_X1 U13620 ( .I(n8552), .ZN(n22666) );
  INV_X1 U13621 ( .I(n22485), .ZN(n2986) );
  INV_X2 U13622 ( .I(n16667), .ZN(n1661) );
  INV_X1 U13624 ( .I(n19221), .ZN(n22675) );
  AOI21_X1 U13626 ( .A1(n12567), .A2(n22162), .B(n19890), .ZN(n6773) );
  INV_X1 U13627 ( .I(n12324), .ZN(n6121) );
  NOR2_X1 U13628 ( .A1(n12325), .A2(n19801), .ZN(n6120) );
  OAI21_X1 U13629 ( .A1(n12324), .A2(n12325), .B(n19801), .ZN(n6125) );
  INV_X1 U13630 ( .I(n31504), .ZN(n14322) );
  NAND3_X1 U13631 ( .A1(n12661), .A2(n29334), .A3(n12660), .ZN(n10555) );
  NAND2_X1 U13635 ( .A1(n22381), .A2(n22380), .ZN(n22637) );
  INV_X2 U13636 ( .I(n36886), .ZN(n1663) );
  INV_X1 U13642 ( .I(n22298), .ZN(n6015) );
  NAND2_X1 U13645 ( .A1(n19976), .A2(n17096), .ZN(n3236) );
  OAI21_X1 U13647 ( .A1(n8749), .A2(n37089), .B(n4851), .ZN(n7058) );
  NAND2_X1 U13648 ( .A1(n18950), .A2(n18953), .ZN(n17041) );
  NAND2_X1 U13649 ( .A1(n13570), .A2(n11091), .ZN(n4662) );
  INV_X1 U13654 ( .I(n3967), .ZN(n2237) );
  NAND2_X1 U13657 ( .A1(n22242), .A2(n8749), .ZN(n2590) );
  NAND2_X1 U13661 ( .A1(n13279), .A2(n17147), .ZN(n7490) );
  OAI21_X1 U13665 ( .A1(n39075), .A2(n1149), .B(n10092), .ZN(n19284) );
  AND2_X1 U13675 ( .A1(n21801), .A2(n33886), .Z(n19292) );
  NAND2_X1 U13677 ( .A1(n22123), .A2(n11149), .ZN(n12345) );
  NAND2_X1 U13692 ( .A1(n22134), .A2(n1327), .ZN(n11047) );
  NAND2_X1 U13693 ( .A1(n7818), .A2(n7817), .ZN(n7816) );
  NAND2_X1 U13696 ( .A1(n22271), .A2(n12814), .ZN(n5149) );
  AND2_X1 U13700 ( .A1(n22325), .A2(n31092), .Z(n14535) );
  NOR2_X1 U13705 ( .A1(n21363), .A2(n31649), .ZN(n6557) );
  NOR2_X1 U13711 ( .A1(n22089), .A2(n18656), .ZN(n13279) );
  OAI21_X1 U13714 ( .A1(n37089), .A2(n34808), .B(n13055), .ZN(n22403) );
  OAI22_X1 U13718 ( .A1(n6722), .A2(n10261), .B1(n5819), .B2(n22189), .ZN(
        n6721) );
  NAND2_X1 U13719 ( .A1(n1149), .A2(n6129), .ZN(n4661) );
  INV_X1 U13720 ( .I(n10631), .ZN(n7771) );
  NOR2_X1 U13729 ( .A1(n22349), .A2(n916), .ZN(n5577) );
  OAI21_X1 U13730 ( .A1(n14423), .A2(n1332), .B(n19873), .ZN(n5576) );
  NOR3_X1 U13733 ( .A1(n3003), .A2(n3001), .A3(n17359), .ZN(n3002) );
  INV_X1 U13738 ( .I(n5302), .ZN(n20759) );
  INV_X1 U13742 ( .I(n4283), .ZN(n18675) );
  NOR2_X1 U13743 ( .A1(n22147), .A2(n22239), .ZN(n13633) );
  NOR2_X1 U13746 ( .A1(n22267), .A2(n33782), .ZN(n21262) );
  NAND2_X1 U13747 ( .A1(n10434), .A2(n32889), .ZN(n10433) );
  NAND2_X1 U13748 ( .A1(n19486), .A2(n22282), .ZN(n13980) );
  OR2_X1 U13749 ( .A1(n22360), .A2(n31939), .Z(n14683) );
  AOI21_X1 U13750 ( .A1(n22289), .A2(n22041), .B(n2840), .ZN(n13420) );
  NOR2_X1 U13751 ( .A1(n22367), .A2(n22365), .ZN(n13296) );
  NAND2_X1 U13753 ( .A1(n1331), .A2(n36237), .ZN(n4629) );
  NAND2_X1 U13755 ( .A1(n22151), .A2(n33678), .ZN(n17973) );
  INV_X1 U13764 ( .I(n16511), .ZN(n16772) );
  NOR2_X1 U13766 ( .A1(n20869), .A2(n2910), .ZN(n11542) );
  NAND2_X1 U13769 ( .A1(n17639), .A2(n22184), .ZN(n17638) );
  NOR2_X1 U13770 ( .A1(n10681), .A2(n34488), .ZN(n4110) );
  INV_X1 U13771 ( .I(n22111), .ZN(n4932) );
  NAND2_X1 U13772 ( .A1(n36151), .A2(n15493), .ZN(n7294) );
  NAND2_X1 U13776 ( .A1(n9224), .A2(n9223), .ZN(n9222) );
  OR2_X1 U13784 ( .A1(n22030), .A2(n5075), .Z(n9126) );
  OR2_X1 U13785 ( .A1(n34813), .A2(n19873), .Z(n5206) );
  AND4_X1 U13788 ( .A1(n10650), .A2(n685), .A3(n10649), .A4(n10652), .Z(n10651) );
  NOR2_X1 U13794 ( .A1(n17307), .A2(n19773), .ZN(n21261) );
  NOR3_X1 U13796 ( .A1(n22263), .A2(n22262), .A3(n22264), .ZN(n4336) );
  AND2_X1 U13797 ( .A1(n21961), .A2(n22130), .Z(n12255) );
  AND2_X1 U13799 ( .A1(n21961), .A2(n12892), .Z(n6722) );
  INV_X2 U13807 ( .I(n21973), .ZN(n22184) );
  OR2_X1 U13813 ( .A1(n22086), .A2(n36006), .Z(n13837) );
  CLKBUF_X2 U13817 ( .I(n22215), .Z(n9938) );
  INV_X1 U13818 ( .I(n18656), .ZN(n9129) );
  INV_X1 U13823 ( .I(n37089), .ZN(n8439) );
  NAND2_X1 U13824 ( .A1(n1342), .A2(n20679), .ZN(n3678) );
  NAND2_X1 U13826 ( .A1(n21891), .A2(n18758), .ZN(n10417) );
  NAND2_X1 U13834 ( .A1(n5451), .A2(n5391), .ZN(n5448) );
  NOR2_X1 U13835 ( .A1(n12513), .A2(n21733), .ZN(n12512) );
  AOI21_X1 U13842 ( .A1(n21708), .A2(n19271), .B(n21886), .ZN(n21709) );
  INV_X1 U13843 ( .I(n21695), .ZN(n10325) );
  NAND2_X1 U13845 ( .A1(n21710), .A2(n20535), .ZN(n10323) );
  NOR2_X1 U13849 ( .A1(n2458), .A2(n29411), .ZN(n17940) );
  NAND2_X1 U13852 ( .A1(n20037), .A2(n21910), .ZN(n13240) );
  INV_X1 U13854 ( .I(n9102), .ZN(n7183) );
  NAND2_X1 U13856 ( .A1(n7414), .A2(n9863), .ZN(n4241) );
  NAND2_X1 U13857 ( .A1(n13098), .A2(n21557), .ZN(n6799) );
  OAI21_X1 U13867 ( .A1(n12737), .A2(n4116), .B(n5187), .ZN(n12358) );
  OR2_X1 U13869 ( .A1(n21843), .A2(n15031), .Z(n14572) );
  AOI21_X1 U13872 ( .A1(n19822), .A2(n14493), .B(n19708), .ZN(n19707) );
  INV_X1 U13873 ( .I(n21867), .ZN(n10657) );
  NAND2_X1 U13875 ( .A1(n21550), .A2(n20328), .ZN(n6420) );
  AND2_X1 U13877 ( .A1(n16951), .A2(n21789), .Z(n21796) );
  NAND2_X1 U13888 ( .A1(n21443), .A2(n15031), .ZN(n2479) );
  NAND2_X1 U13889 ( .A1(n21442), .A2(n33285), .ZN(n2478) );
  NAND2_X1 U13892 ( .A1(n2045), .A2(n11274), .ZN(n21708) );
  NAND2_X1 U13893 ( .A1(n2990), .A2(n18205), .ZN(n17965) );
  NAND2_X1 U13896 ( .A1(n17886), .A2(n21653), .ZN(n7601) );
  AOI21_X1 U13897 ( .A1(n21373), .A2(n21372), .B(n35973), .ZN(n21374) );
  NAND2_X1 U13898 ( .A1(n8969), .A2(n21410), .ZN(n21127) );
  NAND2_X1 U13899 ( .A1(n14909), .A2(n21833), .ZN(n14908) );
  AND2_X1 U13901 ( .A1(n21901), .A2(n21900), .Z(n14526) );
  OR2_X1 U13904 ( .A1(n33771), .A2(n11851), .Z(n11850) );
  INV_X2 U13907 ( .I(n19091), .ZN(n18710) );
  AND2_X1 U13909 ( .A1(n13959), .A2(n13997), .Z(n13685) );
  NOR2_X1 U13911 ( .A1(n21569), .A2(n3326), .ZN(n3325) );
  NAND2_X1 U13912 ( .A1(n15381), .A2(n6504), .ZN(n15380) );
  AND2_X1 U13913 ( .A1(n21750), .A2(n2532), .Z(n16163) );
  NAND2_X1 U13914 ( .A1(n17233), .A2(n32370), .ZN(n13348) );
  NAND2_X1 U13915 ( .A1(n19169), .A2(n18496), .ZN(n10263) );
  NAND2_X1 U13917 ( .A1(n21545), .A2(n19650), .ZN(n13522) );
  AOI21_X1 U13921 ( .A1(n21923), .A2(n21640), .B(n12738), .ZN(n12737) );
  INV_X1 U13926 ( .I(n10875), .ZN(n9253) );
  NAND2_X1 U13929 ( .A1(n19768), .A2(n4094), .ZN(n21372) );
  INV_X1 U13933 ( .I(n11851), .ZN(n11239) );
  NOR2_X1 U13935 ( .A1(n21718), .A2(n1352), .ZN(n5503) );
  INV_X1 U13939 ( .I(n1814), .ZN(n1813) );
  INV_X1 U13940 ( .I(n21450), .ZN(n16873) );
  NOR2_X1 U13941 ( .A1(n21749), .A2(n21748), .ZN(n18274) );
  INV_X1 U13942 ( .I(n17848), .ZN(n12109) );
  OR3_X1 U13944 ( .A1(n4759), .A2(n21029), .A3(n19850), .Z(n21891) );
  NAND2_X1 U13945 ( .A1(n20587), .A2(n21509), .ZN(n17820) );
  NAND2_X1 U13946 ( .A1(n13997), .A2(n10211), .ZN(n13158) );
  AND2_X1 U13951 ( .A1(n10212), .A2(n695), .Z(n21397) );
  CLKBUF_X2 U13952 ( .I(n21688), .Z(n21853) );
  NOR2_X1 U13956 ( .A1(n21465), .A2(n34922), .ZN(n20752) );
  NOR2_X1 U13960 ( .A1(n19699), .A2(n21894), .ZN(n3326) );
  AND2_X1 U13962 ( .A1(n21699), .A2(n18266), .Z(n19037) );
  INV_X2 U13966 ( .I(n8799), .ZN(n7278) );
  AND2_X1 U13972 ( .A1(n19542), .A2(n21748), .Z(n14542) );
  CLKBUF_X2 U13976 ( .I(n21506), .Z(n9642) );
  CLKBUF_X2 U13980 ( .I(n21846), .Z(n19392) );
  INV_X1 U13986 ( .I(n29689), .ZN(n29690) );
  INV_X1 U13987 ( .I(n30179), .ZN(n3711) );
  INV_X1 U13993 ( .I(n29661), .ZN(n16641) );
  INV_X1 U13994 ( .I(n29849), .ZN(n18691) );
  INV_X1 U13995 ( .I(n30006), .ZN(n30007) );
  CLKBUF_X2 U13998 ( .I(n21849), .Z(n18219) );
  INV_X1 U14001 ( .I(n30114), .ZN(n30115) );
  INV_X1 U14003 ( .I(n19950), .ZN(n6462) );
  INV_X1 U14004 ( .I(n19801), .ZN(n6429) );
  INV_X1 U14005 ( .I(n29857), .ZN(n20420) );
  INV_X1 U14009 ( .I(n19758), .ZN(n17316) );
  INV_X1 U14010 ( .I(n29808), .ZN(n22285) );
  INV_X1 U14011 ( .I(n29320), .ZN(n29321) );
  CLKBUF_X2 U14013 ( .I(n21776), .Z(n19350) );
  INV_X1 U14014 ( .I(n29238), .ZN(n29239) );
  INV_X1 U14015 ( .I(n19732), .ZN(n21048) );
  INV_X2 U14017 ( .I(n8653), .ZN(n8799) );
  INV_X1 U14019 ( .I(n19761), .ZN(n15599) );
  INV_X1 U14020 ( .I(n19583), .ZN(n15888) );
  INV_X1 U14023 ( .I(n15009), .ZN(n21782) );
  CLKBUF_X2 U14024 ( .I(Key[134]), .Z(n19913) );
  INV_X1 U14025 ( .I(Key[178]), .ZN(n11200) );
  CLKBUF_X2 U14030 ( .I(Key[87]), .Z(n28934) );
  CLKBUF_X2 U14035 ( .I(Key[131]), .Z(n30248) );
  CLKBUF_X2 U14037 ( .I(Key[83]), .Z(n29432) );
  CLKBUF_X2 U14038 ( .I(Key[152]), .Z(n19883) );
  CLKBUF_X2 U14039 ( .I(Key[53]), .Z(n29319) );
  INV_X1 U14042 ( .I(n29295), .ZN(n1706) );
  CLKBUF_X2 U14045 ( .I(Key[111]), .Z(n19814) );
  CLKBUF_X2 U14046 ( .I(Key[89]), .Z(n29671) );
  CLKBUF_X2 U14048 ( .I(Key[71]), .Z(n10027) );
  CLKBUF_X2 U14050 ( .I(Key[32]), .Z(n28968) );
  CLKBUF_X2 U14051 ( .I(Key[57]), .Z(n29476) );
  CLKBUF_X2 U14056 ( .I(Key[101]), .Z(n29298) );
  CLKBUF_X2 U14057 ( .I(Key[186]), .Z(n19936) );
  INV_X1 U14058 ( .I(n19825), .ZN(n1726) );
  CLKBUF_X2 U14059 ( .I(Key[35]), .Z(n29707) );
  CLKBUF_X2 U14060 ( .I(Key[161]), .Z(n29229) );
  CLKBUF_X2 U14064 ( .I(Key[128]), .Z(n19649) );
  CLKBUF_X2 U14066 ( .I(Key[171]), .Z(n29661) );
  INV_X1 U14067 ( .I(n30063), .ZN(n1737) );
  CLKBUF_X2 U14069 ( .I(Key[59]), .Z(n29562) );
  CLKBUF_X2 U14070 ( .I(Key[178]), .Z(n19749) );
  XOR2_X1 U14071 ( .A1(n1740), .A2(n4041), .Z(n1769) );
  NOR3_X1 U14082 ( .A1(n14791), .A2(n9514), .A3(n1753), .ZN(n1752) );
  XOR2_X1 U14086 ( .A1(n36895), .A2(n23609), .Z(n23771) );
  XOR2_X1 U14087 ( .A1(n17478), .A2(n36895), .Z(n10885) );
  NOR2_X1 U14088 ( .A1(n20873), .A2(n906), .ZN(n18851) );
  XOR2_X1 U14089 ( .A1(n1758), .A2(n22385), .Z(n17628) );
  NAND2_X1 U14092 ( .A1(n1759), .A2(n15038), .ZN(n19327) );
  NAND2_X2 U14095 ( .A1(n3380), .A2(n1760), .ZN(n26553) );
  XOR2_X1 U14099 ( .A1(n10026), .A2(n16134), .Z(n18966) );
  XOR2_X1 U14105 ( .A1(n22416), .A2(n22417), .Z(n1765) );
  NAND2_X2 U14107 ( .A1(n3226), .A2(n1284), .ZN(n23818) );
  NAND2_X1 U14113 ( .A1(n1771), .A2(n13113), .ZN(n13047) );
  NAND2_X1 U14114 ( .A1(n1771), .A2(n13112), .ZN(n13048) );
  XOR2_X1 U14115 ( .A1(n29029), .A2(n9952), .Z(n2217) );
  XOR2_X1 U14120 ( .A1(n1775), .A2(n28783), .Z(n28945) );
  XOR2_X1 U14122 ( .A1(n1775), .A2(n19816), .Z(n8774) );
  XOR2_X1 U14123 ( .A1(n1775), .A2(n29831), .Z(n29834) );
  NAND3_X1 U14125 ( .A1(n35287), .A2(n4434), .A3(n38079), .ZN(n27317) );
  NAND2_X1 U14130 ( .A1(n27298), .A2(n1788), .ZN(n5082) );
  XOR2_X1 U14136 ( .A1(n13395), .A2(n19733), .Z(n1790) );
  XOR2_X1 U14137 ( .A1(n23712), .A2(n18006), .Z(n24062) );
  NOR2_X2 U14138 ( .A1(n16033), .A2(n16032), .ZN(n18006) );
  XOR2_X1 U14145 ( .A1(n29073), .A2(n1793), .Z(n1792) );
  XOR2_X1 U14146 ( .A1(n20452), .A2(n29509), .Z(n1793) );
  XOR2_X1 U14150 ( .A1(n13289), .A2(n19875), .Z(n18182) );
  AOI21_X2 U14151 ( .A1(n34036), .A2(n35258), .B(n1796), .ZN(n13293) );
  OAI21_X1 U14152 ( .A1(n29862), .A2(n29960), .B(n29955), .ZN(n15140) );
  NOR2_X2 U14154 ( .A1(n24863), .A2(n13966), .ZN(n24862) );
  NAND2_X2 U14155 ( .A1(n4178), .A2(n4177), .ZN(n24863) );
  INV_X1 U14158 ( .I(n29844), .ZN(n5972) );
  NAND2_X1 U14159 ( .A1(n1063), .A2(n20284), .ZN(n29844) );
  XOR2_X1 U14163 ( .A1(n16898), .A2(n1808), .Z(n1807) );
  XOR2_X1 U14164 ( .A1(n17908), .A2(n22568), .Z(n1809) );
  NAND2_X1 U14168 ( .A1(n11344), .A2(n1812), .ZN(n21989) );
  INV_X2 U14170 ( .I(n1816), .ZN(n21886) );
  INV_X2 U14177 ( .I(n10962), .ZN(n13042) );
  INV_X1 U14178 ( .I(n23080), .ZN(n23104) );
  XOR2_X1 U14179 ( .A1(n10963), .A2(n7708), .Z(n10962) );
  NOR2_X1 U14185 ( .A1(n425), .A2(n1827), .ZN(n20850) );
  NAND2_X1 U14187 ( .A1(n25738), .A2(n34485), .ZN(n5236) );
  XOR2_X1 U14188 ( .A1(n35215), .A2(n16296), .Z(n16338) );
  MUX2_X1 U14191 ( .I0(n1836), .I1(n1835), .S(n34520), .Z(n1834) );
  NAND2_X1 U14192 ( .A1(n30358), .A2(n27390), .ZN(n1836) );
  OAI22_X2 U14198 ( .A1(n8316), .A2(n38369), .B1(n8315), .B2(n1844), .ZN(
        n24985) );
  XOR2_X1 U14206 ( .A1(n23833), .A2(n23801), .Z(n21268) );
  XOR2_X1 U14207 ( .A1(n23695), .A2(n23707), .Z(n23833) );
  XOR2_X1 U14220 ( .A1(n22758), .A2(n1868), .Z(n1867) );
  XOR2_X1 U14228 ( .A1(n1878), .A2(n19627), .Z(n4853) );
  XNOR2_X1 U14229 ( .A1(n10965), .A2(n26554), .ZN(n19627) );
  XOR2_X1 U14231 ( .A1(n1880), .A2(n1879), .Z(n1878) );
  XOR2_X1 U14237 ( .A1(n16864), .A2(n19843), .Z(n1884) );
  XOR2_X1 U14239 ( .A1(n24857), .A2(n25132), .Z(n1885) );
  XOR2_X1 U14241 ( .A1(n25016), .A2(n25266), .Z(n19797) );
  MUX2_X1 U14245 ( .I0(n30134), .I1(n37117), .S(n35234), .Z(n3898) );
  XOR2_X1 U14256 ( .A1(n1897), .A2(n10617), .Z(n1896) );
  XOR2_X1 U14259 ( .A1(n39637), .A2(n29357), .Z(n1902) );
  INV_X2 U14260 ( .I(n5966), .ZN(n2716) );
  XOR2_X1 U14268 ( .A1(n1913), .A2(n1912), .Z(n1911) );
  XOR2_X1 U14269 ( .A1(n5652), .A2(n39082), .Z(n1912) );
  XOR2_X1 U14271 ( .A1(n28948), .A2(n38195), .Z(n1913) );
  NAND2_X2 U14276 ( .A1(n15321), .A2(n15323), .ZN(n29147) );
  NAND2_X1 U14288 ( .A1(n5570), .A2(n2121), .ZN(n2856) );
  NAND3_X1 U14292 ( .A1(n25480), .A2(n36083), .A3(n1539), .ZN(n25332) );
  XOR2_X1 U14301 ( .A1(n1930), .A2(n25015), .Z(n2623) );
  NAND2_X1 U14307 ( .A1(n10015), .A2(n26215), .ZN(n1934) );
  OAI21_X2 U14311 ( .A1(n10336), .A2(n10337), .B(n9493), .ZN(n19606) );
  XOR2_X1 U14322 ( .A1(n1945), .A2(n1947), .Z(n17564) );
  XOR2_X1 U14323 ( .A1(n22723), .A2(n1946), .Z(n1945) );
  XOR2_X1 U14324 ( .A1(n22444), .A2(n30803), .Z(n1946) );
  NAND3_X1 U14334 ( .A1(n26101), .A2(n11148), .A3(n35207), .ZN(n1954) );
  INV_X2 U14340 ( .I(n1961), .ZN(n20673) );
  OR2_X1 U14346 ( .A1(n22145), .A2(n19180), .Z(n1966) );
  NAND2_X2 U14350 ( .A1(n1003), .A2(n865), .ZN(n26743) );
  XOR2_X1 U14351 ( .A1(n7543), .A2(n857), .Z(n9618) );
  XOR2_X1 U14362 ( .A1(n38180), .A2(n1366), .Z(n1980) );
  XOR2_X1 U14364 ( .A1(n26165), .A2(n26180), .Z(n26229) );
  INV_X2 U14372 ( .I(n13994), .ZN(n2047) );
  AND2_X1 U14376 ( .A1(n25528), .A2(n36083), .Z(n1991) );
  OAI21_X2 U14380 ( .A1(n2698), .A2(n19836), .B(n1995), .ZN(n19725) );
  XOR2_X1 U14388 ( .A1(n2004), .A2(n2003), .Z(n2002) );
  XOR2_X1 U14389 ( .A1(n29247), .A2(n19681), .Z(n2003) );
  XOR2_X1 U14393 ( .A1(n36596), .A2(n35559), .Z(n10201) );
  NAND2_X1 U14396 ( .A1(n21925), .A2(n2008), .ZN(n3437) );
  OAI21_X2 U14399 ( .A1(n2017), .A2(n2016), .B(n2013), .ZN(n29672) );
  INV_X1 U14404 ( .I(n24404), .ZN(n13443) );
  NAND2_X2 U14409 ( .A1(n20200), .A2(n20201), .ZN(n9597) );
  XOR2_X1 U14414 ( .A1(n25183), .A2(n24936), .Z(n2025) );
  NOR2_X1 U14419 ( .A1(n2423), .A2(n2029), .ZN(n17371) );
  NOR2_X1 U14420 ( .A1(n30302), .A2(n2029), .ZN(n25847) );
  NOR2_X1 U14421 ( .A1(n5356), .A2(n2029), .ZN(n4154) );
  XOR2_X1 U14427 ( .A1(n2032), .A2(n28871), .Z(n2031) );
  XOR2_X1 U14429 ( .A1(n29289), .A2(n28790), .Z(n28871) );
  NOR2_X2 U14433 ( .A1(n16968), .A2(n3093), .ZN(n3092) );
  XOR2_X1 U14438 ( .A1(n35241), .A2(n11755), .Z(n2041) );
  XOR2_X1 U14449 ( .A1(n15202), .A2(n2044), .Z(n23739) );
  NAND2_X1 U14452 ( .A1(n7210), .A2(n24383), .ZN(n6570) );
  XOR2_X1 U14460 ( .A1(n14260), .A2(n29647), .Z(n20513) );
  NOR2_X2 U14461 ( .A1(n21110), .A2(n21109), .ZN(n14260) );
  XOR2_X1 U14469 ( .A1(n37312), .A2(n1559), .Z(n2064) );
  XOR2_X1 U14471 ( .A1(n9939), .A2(n657), .Z(n2065) );
  XOR2_X1 U14477 ( .A1(n31062), .A2(n35238), .Z(n2067) );
  AOI21_X2 U14482 ( .A1(n25924), .A2(n25961), .B(n25805), .ZN(n26554) );
  XOR2_X1 U14484 ( .A1(n2070), .A2(n1367), .Z(Ciphertext[119]) );
  XOR2_X1 U14486 ( .A1(n34564), .A2(n19730), .Z(n16555) );
  NAND2_X1 U14489 ( .A1(n1573), .A2(n24812), .ZN(n2075) );
  NAND2_X1 U14490 ( .A1(n24615), .A2(n18983), .ZN(n2076) );
  OAI21_X2 U14492 ( .A1(n31214), .A2(n2233), .B(n2082), .ZN(n2234) );
  AOI21_X2 U14493 ( .A1(n3972), .A2(n22204), .B(n3971), .ZN(n2233) );
  INV_X2 U14497 ( .I(n3021), .ZN(n18576) );
  NAND2_X1 U14498 ( .A1(n21820), .A2(n18722), .ZN(n2092) );
  INV_X2 U14499 ( .I(n2094), .ZN(n18815) );
  XOR2_X1 U14502 ( .A1(n28835), .A2(n2097), .Z(n2096) );
  XOR2_X1 U14503 ( .A1(n14039), .A2(n19947), .Z(n2097) );
  XOR2_X1 U14506 ( .A1(n542), .A2(n9035), .Z(n28834) );
  AOI21_X2 U14513 ( .A1(n24780), .A2(n24783), .B(n17936), .ZN(n25298) );
  INV_X2 U14517 ( .I(n21277), .ZN(n26959) );
  XOR2_X1 U14518 ( .A1(n27690), .A2(n2281), .Z(n27756) );
  XOR2_X1 U14523 ( .A1(n2106), .A2(n2105), .Z(n2104) );
  XOR2_X1 U14524 ( .A1(n23728), .A2(n29522), .Z(n2105) );
  NOR3_X1 U14528 ( .A1(n29683), .A2(n31538), .A3(n38206), .ZN(n2112) );
  XOR2_X1 U14540 ( .A1(n2122), .A2(n28841), .Z(n14438) );
  XOR2_X1 U14551 ( .A1(n32298), .A2(n29221), .Z(n2135) );
  XOR2_X1 U14552 ( .A1(n33470), .A2(n27862), .Z(n2136) );
  NAND2_X2 U14553 ( .A1(n27375), .A2(n27376), .ZN(n27862) );
  XOR2_X1 U14557 ( .A1(n38144), .A2(n27178), .Z(n2138) );
  NAND2_X1 U14568 ( .A1(n2147), .A2(n28745), .ZN(n4024) );
  XOR2_X1 U14584 ( .A1(n29840), .A2(n4268), .Z(n2162) );
  XOR2_X1 U14585 ( .A1(n29070), .A2(n28948), .Z(n29840) );
  OAI21_X2 U14592 ( .A1(n25430), .A2(n30633), .B(n2167), .ZN(n17180) );
  XOR2_X1 U14597 ( .A1(n24043), .A2(n24042), .Z(n2170) );
  XOR2_X1 U14606 ( .A1(n2177), .A2(n39579), .Z(n2176) );
  XOR2_X1 U14607 ( .A1(n18051), .A2(n2178), .Z(n2177) );
  XOR2_X1 U14617 ( .A1(n25263), .A2(n19359), .Z(n2185) );
  NOR2_X1 U14620 ( .A1(n2187), .A2(n18576), .ZN(n2189) );
  NAND2_X1 U14623 ( .A1(n16237), .A2(n8537), .ZN(n16243) );
  OAI21_X1 U14627 ( .A1(n31875), .A2(n16237), .B(n8538), .ZN(n8534) );
  XOR2_X1 U14631 ( .A1(n36758), .A2(n18180), .Z(n2195) );
  XOR2_X1 U14636 ( .A1(n2199), .A2(n14609), .Z(n2198) );
  XOR2_X1 U14637 ( .A1(n1659), .A2(n4139), .Z(n2199) );
  AOI21_X2 U14641 ( .A1(n22849), .A2(n12925), .B(n6018), .ZN(n23200) );
  NOR2_X1 U14643 ( .A1(n22849), .A2(n36369), .ZN(n2202) );
  XOR2_X1 U14644 ( .A1(n2203), .A2(n19874), .Z(Ciphertext[118]) );
  NAND2_X1 U14645 ( .A1(n21018), .A2(n524), .ZN(n21017) );
  XOR2_X1 U14647 ( .A1(n4135), .A2(n2209), .Z(n4137) );
  XOR2_X1 U14652 ( .A1(n2215), .A2(n2214), .Z(n20687) );
  XOR2_X1 U14653 ( .A1(n2978), .A2(n11151), .Z(n2214) );
  XOR2_X1 U14659 ( .A1(n2221), .A2(n32973), .Z(n2220) );
  XOR2_X1 U14663 ( .A1(n24031), .A2(n24032), .Z(n2222) );
  NOR2_X2 U14664 ( .A1(n10109), .A2(n2223), .ZN(n24031) );
  AOI21_X1 U14670 ( .A1(n3697), .A2(n1030), .B(n20728), .ZN(n2231) );
  XOR2_X1 U14671 ( .A1(n8083), .A2(n34553), .Z(n2235) );
  NAND2_X2 U14672 ( .A1(n2707), .A2(n2705), .ZN(n8083) );
  XOR2_X1 U14674 ( .A1(n2234), .A2(n2235), .Z(n3999) );
  INV_X2 U14675 ( .I(n8083), .ZN(n7287) );
  NAND2_X2 U14682 ( .A1(n35059), .A2(n26039), .ZN(n26214) );
  XOR2_X1 U14689 ( .A1(n828), .A2(n2263), .Z(n15050) );
  XOR2_X1 U14691 ( .A1(n449), .A2(n29602), .Z(n2263) );
  INV_X2 U14692 ( .I(n2264), .ZN(n28163) );
  MUX2_X1 U14694 ( .I0(n4945), .I1(n16363), .S(n28163), .Z(n28164) );
  NAND2_X2 U14698 ( .A1(n2270), .A2(n28308), .ZN(n29122) );
  NAND3_X1 U14703 ( .A1(n23521), .A2(n30835), .A3(n2273), .ZN(n23406) );
  AOI22_X1 U14706 ( .A1(n21821), .A2(n38246), .B1(n22240), .B2(n22239), .ZN(
        n19012) );
  NOR2_X1 U14707 ( .A1(n1349), .A2(n2277), .ZN(n2279) );
  AND2_X1 U14708 ( .A1(n918), .A2(n19388), .Z(n2280) );
  XOR2_X1 U14714 ( .A1(n29066), .A2(n2285), .Z(n2284) );
  XOR2_X1 U14715 ( .A1(n1413), .A2(n19571), .Z(n2285) );
  XOR2_X1 U14731 ( .A1(n2301), .A2(Plaintext[65]), .Z(n3021) );
  INV_X1 U14732 ( .I(Key[65]), .ZN(n2301) );
  INV_X2 U14736 ( .I(n2309), .ZN(n19966) );
  XOR2_X1 U14742 ( .A1(n35062), .A2(n23846), .Z(n7127) );
  XOR2_X1 U14743 ( .A1(n24061), .A2(n35062), .Z(n23711) );
  XOR2_X1 U14745 ( .A1(n35062), .A2(n36895), .Z(n16004) );
  AOI21_X1 U14754 ( .A1(n26039), .A2(n31340), .B(n20813), .ZN(n2326) );
  NAND2_X2 U14757 ( .A1(n2328), .A2(n2327), .ZN(n28850) );
  OR2_X1 U14758 ( .A1(n18875), .A2(n31663), .Z(n2330) );
  MUX2_X1 U14759 ( .I0(n28735), .I1(n32682), .S(n31554), .Z(n2331) );
  AOI21_X2 U14760 ( .A1(n28058), .A2(n28057), .B(n28056), .ZN(n28735) );
  INV_X1 U14766 ( .I(n11390), .ZN(n2335) );
  NOR2_X1 U14773 ( .A1(n35187), .A2(n10118), .ZN(n16275) );
  OR2_X1 U14776 ( .A1(n10734), .A2(n16792), .Z(n15701) );
  XOR2_X1 U14777 ( .A1(n12200), .A2(n15987), .Z(n10734) );
  XOR2_X1 U14784 ( .A1(n3475), .A2(n37974), .Z(n2354) );
  NAND2_X1 U14794 ( .A1(n38364), .A2(n38013), .ZN(n14444) );
  NOR2_X1 U14797 ( .A1(n10938), .A2(n2366), .ZN(n10444) );
  XOR2_X1 U14799 ( .A1(n23807), .A2(n2367), .Z(n3376) );
  XOR2_X1 U14800 ( .A1(n23910), .A2(n1369), .Z(n2367) );
  OAI21_X2 U14803 ( .A1(n2369), .A2(n17454), .B(n2368), .ZN(n5841) );
  XOR2_X1 U14810 ( .A1(n12430), .A2(n39359), .Z(n2371) );
  NOR2_X2 U14819 ( .A1(n19918), .A2(n7974), .ZN(n27027) );
  NAND2_X2 U14820 ( .A1(n27249), .A2(n7974), .ZN(n27250) );
  NAND2_X1 U14821 ( .A1(n29441), .A2(n29437), .ZN(n29423) );
  XOR2_X1 U14822 ( .A1(n2382), .A2(n2379), .Z(n20032) );
  XOR2_X1 U14823 ( .A1(n35266), .A2(n1698), .Z(n2379) );
  XOR2_X1 U14826 ( .A1(n27850), .A2(n27672), .Z(n2382) );
  XOR2_X1 U14830 ( .A1(n17398), .A2(n2389), .Z(n2387) );
  XOR2_X1 U14831 ( .A1(n19194), .A2(n9271), .Z(n2388) );
  XOR2_X1 U14832 ( .A1(n2390), .A2(n12972), .Z(n19194) );
  XOR2_X1 U14833 ( .A1(n16138), .A2(n19845), .Z(n2389) );
  INV_X2 U14836 ( .I(n2391), .ZN(n28033) );
  XOR2_X1 U14855 ( .A1(n23677), .A2(n23891), .Z(n2402) );
  NOR2_X2 U14858 ( .A1(n21557), .A2(n21917), .ZN(n21622) );
  INV_X2 U14864 ( .I(n10665), .ZN(n25365) );
  INV_X1 U14870 ( .I(n2424), .ZN(n26068) );
  NAND2_X1 U14872 ( .A1(n38914), .A2(n26070), .ZN(n25371) );
  XOR2_X1 U14886 ( .A1(n38219), .A2(n29838), .Z(n14772) );
  XOR2_X1 U14888 ( .A1(n13496), .A2(n38218), .Z(n26374) );
  XOR2_X1 U14893 ( .A1(n24970), .A2(n2446), .Z(n2445) );
  XNOR2_X1 U14894 ( .A1(n20707), .A2(n25163), .ZN(n24970) );
  NAND2_X1 U14897 ( .A1(n9103), .A2(n13433), .ZN(n2450) );
  INV_X2 U14900 ( .I(n25636), .ZN(n25637) );
  NOR2_X1 U14911 ( .A1(n2467), .A2(n28128), .ZN(n14117) );
  XOR2_X1 U14915 ( .A1(n20335), .A2(n22790), .Z(n22654) );
  NOR2_X2 U14918 ( .A1(n22024), .A2(n22023), .ZN(n22491) );
  XOR2_X1 U14920 ( .A1(n2476), .A2(n2475), .Z(n2474) );
  XOR2_X1 U14921 ( .A1(n23776), .A2(n1711), .Z(n2475) );
  NAND2_X2 U14929 ( .A1(n2479), .A2(n2478), .ZN(n8431) );
  NAND2_X2 U14930 ( .A1(n2482), .A2(n2481), .ZN(n4424) );
  OAI21_X1 U14931 ( .A1(n16873), .A2(n12109), .B(n5733), .ZN(n2482) );
  XOR2_X1 U14933 ( .A1(n2485), .A2(n1713), .Z(Ciphertext[152]) );
  XOR2_X1 U14935 ( .A1(n35404), .A2(n32765), .Z(n9695) );
  XOR2_X1 U14937 ( .A1(n25214), .A2(n32765), .Z(n3427) );
  XOR2_X1 U14938 ( .A1(n32765), .A2(n17395), .Z(n10617) );
  XOR2_X1 U14955 ( .A1(n23865), .A2(n7129), .Z(n2510) );
  XOR2_X1 U14956 ( .A1(n23712), .A2(n3601), .Z(n23865) );
  XOR2_X1 U14959 ( .A1(n20509), .A2(n2656), .Z(n7129) );
  NOR2_X2 U14961 ( .A1(n6911), .A2(n6910), .ZN(n2656) );
  XOR2_X1 U14970 ( .A1(n31537), .A2(n14069), .Z(n2515) );
  XOR2_X1 U14972 ( .A1(n2526), .A2(n2525), .Z(n2524) );
  XOR2_X1 U14973 ( .A1(n24049), .A2(n1370), .Z(n2525) );
  XOR2_X1 U14977 ( .A1(n3609), .A2(n17462), .Z(n2529) );
  XOR2_X1 U14980 ( .A1(n38581), .A2(n31543), .Z(n24892) );
  XOR2_X1 U14982 ( .A1(n35707), .A2(n31543), .Z(n13918) );
  XNOR2_X1 U14986 ( .A1(Plaintext[106]), .A2(Key[106]), .ZN(n2533) );
  NAND2_X1 U14988 ( .A1(n11033), .A2(n2534), .ZN(n2679) );
  NAND2_X2 U14997 ( .A1(n16820), .A2(n2537), .ZN(n16819) );
  XOR2_X1 U14999 ( .A1(Plaintext[128]), .A2(Key[128]), .Z(n11702) );
  XOR2_X1 U15001 ( .A1(n35208), .A2(n37110), .Z(n2543) );
  XOR2_X1 U15003 ( .A1(n871), .A2(n2544), .Z(n14174) );
  XOR2_X1 U15004 ( .A1(n27749), .A2(n19815), .Z(n2544) );
  NAND3_X1 U15009 ( .A1(n30699), .A2(n37983), .A3(n32882), .ZN(n24748) );
  NAND2_X2 U15020 ( .A1(n939), .A2(n3462), .ZN(n11939) );
  INV_X2 U15021 ( .I(n2572), .ZN(n20309) );
  NAND2_X2 U15023 ( .A1(n2667), .A2(n2666), .ZN(n6287) );
  XOR2_X1 U15039 ( .A1(n26491), .A2(n26493), .Z(n2592) );
  XOR2_X1 U15043 ( .A1(n2596), .A2(n18179), .Z(n19142) );
  OAI21_X1 U15048 ( .A1(n2599), .A2(n2601), .B(n2598), .ZN(n23219) );
  XOR2_X1 U15055 ( .A1(n13090), .A2(n5090), .Z(n20406) );
  NAND2_X1 U15058 ( .A1(n24581), .A2(n24904), .ZN(n2610) );
  INV_X2 U15065 ( .I(n13207), .ZN(n17105) );
  NAND2_X1 U15067 ( .A1(n17351), .A2(n2616), .ZN(n24800) );
  XOR2_X1 U15072 ( .A1(n25148), .A2(n724), .Z(n2622) );
  XOR2_X1 U15075 ( .A1(n282), .A2(n2627), .Z(n6351) );
  XOR2_X1 U15076 ( .A1(n2627), .A2(n27540), .Z(n12495) );
  XOR2_X1 U15077 ( .A1(n2627), .A2(n19952), .Z(n12855) );
  XOR2_X1 U15079 ( .A1(n2627), .A2(n27802), .Z(n27630) );
  INV_X1 U15081 ( .I(n33703), .ZN(n23263) );
  NOR2_X2 U15089 ( .A1(n6636), .A2(n2340), .ZN(n10988) );
  NAND2_X1 U15090 ( .A1(n2634), .A2(n9825), .ZN(n24662) );
  OR2_X1 U15093 ( .A1(n18573), .A2(n1029), .Z(n2635) );
  XOR2_X1 U15095 ( .A1(n28836), .A2(n770), .Z(n2637) );
  XOR2_X1 U15100 ( .A1(n2646), .A2(n2648), .Z(n11224) );
  XOR2_X1 U15101 ( .A1(n26241), .A2(n2647), .Z(n2646) );
  XOR2_X1 U15102 ( .A1(n26439), .A2(n36958), .Z(n2647) );
  XOR2_X1 U15103 ( .A1(n15010), .A2(n2649), .Z(n2648) );
  XOR2_X1 U15104 ( .A1(n9989), .A2(n3413), .Z(n2649) );
  OAI21_X2 U15105 ( .A1(n18273), .A2(n34148), .B(n7862), .ZN(n15010) );
  XOR2_X1 U15106 ( .A1(n2650), .A2(n711), .Z(n22897) );
  XOR2_X1 U15108 ( .A1(n9497), .A2(n2838), .Z(n2651) );
  XOR2_X1 U15110 ( .A1(n2653), .A2(n25290), .Z(n25291) );
  NAND2_X1 U15113 ( .A1(n21982), .A2(n2654), .ZN(n3137) );
  XOR2_X1 U15117 ( .A1(n2656), .A2(n29838), .Z(n10402) );
  XOR2_X1 U15118 ( .A1(n2656), .A2(n19683), .Z(n17006) );
  NOR2_X1 U15128 ( .A1(n7355), .A2(n32434), .ZN(n2671) );
  OAI21_X2 U15130 ( .A1(n2677), .A2(n2674), .B(n2675), .ZN(n16502) );
  AND2_X1 U15131 ( .A1(n24162), .A2(n1603), .Z(n2677) );
  NAND2_X2 U15136 ( .A1(n26447), .A2(n14682), .ZN(n27556) );
  NAND3_X1 U15151 ( .A1(n1337), .A2(n36006), .A3(n32434), .ZN(n22021) );
  OAI21_X1 U15152 ( .A1(n22019), .A2(n2816), .B(n32434), .ZN(n2705) );
  XOR2_X1 U15159 ( .A1(n2714), .A2(n2713), .Z(n2712) );
  XOR2_X1 U15160 ( .A1(n26531), .A2(n19592), .Z(n2713) );
  NOR2_X1 U15165 ( .A1(n27305), .A2(n34853), .ZN(n12427) );
  XOR2_X1 U15171 ( .A1(n3126), .A2(n2728), .Z(n2727) );
  XOR2_X1 U15173 ( .A1(n37059), .A2(n18430), .Z(n2728) );
  AOI21_X2 U15180 ( .A1(n9580), .A2(n9581), .B(n9579), .ZN(n24674) );
  XOR2_X1 U15181 ( .A1(n22552), .A2(n22743), .Z(n18943) );
  XOR2_X1 U15184 ( .A1(n23894), .A2(n3601), .Z(n23663) );
  XOR2_X1 U15191 ( .A1(n9979), .A2(n23695), .Z(n2738) );
  XOR2_X1 U15196 ( .A1(n15165), .A2(n3110), .Z(n11603) );
  INV_X2 U15203 ( .I(n2742), .ZN(n8245) );
  XOR2_X1 U15205 ( .A1(n22438), .A2(n5247), .Z(n2743) );
  XOR2_X1 U15212 ( .A1(n20212), .A2(n14569), .Z(n2753) );
  NOR2_X1 U15218 ( .A1(n4105), .A2(n36840), .ZN(n9489) );
  NAND2_X1 U15220 ( .A1(n9756), .A2(n36840), .ZN(n27113) );
  XOR2_X1 U15224 ( .A1(n27565), .A2(n674), .Z(n2757) );
  XOR2_X1 U15225 ( .A1(n27829), .A2(n27766), .Z(n27565) );
  NOR2_X1 U15233 ( .A1(n34808), .A2(n2765), .ZN(n22242) );
  INV_X2 U15248 ( .I(n2778), .ZN(n7705) );
  XOR2_X1 U15253 ( .A1(n2781), .A2(n2780), .Z(n22813) );
  XOR2_X1 U15254 ( .A1(n9206), .A2(n9207), .Z(n2780) );
  NOR2_X2 U15258 ( .A1(n10052), .A2(n17254), .ZN(n28722) );
  XOR2_X1 U15269 ( .A1(n10582), .A2(n25245), .Z(n2800) );
  XOR2_X1 U15270 ( .A1(n27831), .A2(n15736), .Z(n2815) );
  NAND2_X1 U15273 ( .A1(n25484), .A2(n2803), .ZN(n25375) );
  NAND2_X1 U15274 ( .A1(n32904), .A2(n2803), .ZN(n25462) );
  XOR2_X1 U15277 ( .A1(n2806), .A2(n2808), .Z(n2805) );
  XOR2_X1 U15279 ( .A1(n24038), .A2(n23886), .Z(n2808) );
  OAI21_X2 U15282 ( .A1(n2814), .A2(n34245), .B(n2813), .ZN(n23894) );
  INV_X2 U15283 ( .I(n2819), .ZN(n26863) );
  XOR2_X1 U15290 ( .A1(n39798), .A2(n39482), .Z(n2825) );
  INV_X2 U15294 ( .I(n9133), .ZN(n24366) );
  XOR2_X1 U15312 ( .A1(n26275), .A2(n17428), .Z(n2864) );
  INV_X1 U15314 ( .I(n2867), .ZN(n5900) );
  XOR2_X1 U15316 ( .A1(n29964), .A2(n2867), .Z(n9270) );
  XOR2_X1 U15317 ( .A1(n2867), .A2(n27776), .Z(n16551) );
  NAND2_X2 U15318 ( .A1(n3468), .A2(n3467), .ZN(n2867) );
  INV_X2 U15319 ( .I(n19888), .ZN(n28224) );
  NAND3_X2 U15325 ( .A1(n2873), .A2(n2874), .A3(n2872), .ZN(n3538) );
  INV_X2 U15331 ( .I(n2881), .ZN(n4472) );
  XOR2_X1 U15333 ( .A1(n3999), .A2(n4000), .Z(n2881) );
  INV_X2 U15335 ( .I(n2895), .ZN(n24536) );
  XOR2_X1 U15340 ( .A1(n467), .A2(n29131), .Z(n29047) );
  INV_X2 U15351 ( .I(n16704), .ZN(n30238) );
  NAND2_X2 U15361 ( .A1(n2920), .A2(n2919), .ZN(n23774) );
  OAI21_X2 U15362 ( .A1(n19281), .A2(n13262), .B(n23086), .ZN(n17017) );
  XOR2_X1 U15369 ( .A1(n27466), .A2(n29238), .Z(n8397) );
  NAND2_X2 U15373 ( .A1(n14351), .A2(n14352), .ZN(n4618) );
  XOR2_X1 U15374 ( .A1(n25263), .A2(n31568), .Z(n13711) );
  XOR2_X1 U15375 ( .A1(n25182), .A2(n31568), .Z(n20805) );
  XOR2_X1 U15377 ( .A1(n13076), .A2(n2931), .Z(n15451) );
  XOR2_X1 U15379 ( .A1(n23996), .A2(n38880), .Z(n9271) );
  XOR2_X1 U15384 ( .A1(n22648), .A2(n19950), .Z(n2935) );
  NOR2_X2 U15388 ( .A1(n20226), .A2(n20225), .ZN(n9878) );
  AOI21_X1 U15390 ( .A1(n15360), .A2(n32020), .B(n27357), .ZN(n21169) );
  MUX2_X1 U15391 ( .I0(n27066), .I1(n27067), .S(n1000), .Z(n27068) );
  XOR2_X1 U15399 ( .A1(n2943), .A2(n5652), .Z(n16587) );
  XOR2_X1 U15400 ( .A1(n2943), .A2(n28886), .Z(n28794) );
  AOI21_X1 U15405 ( .A1(n2947), .A2(n495), .B(n27406), .ZN(n2949) );
  XNOR2_X1 U15406 ( .A1(n23419), .A2(n23965), .ZN(n24026) );
  AND2_X1 U15410 ( .A1(n13468), .A2(n6894), .Z(n2957) );
  XOR2_X1 U15422 ( .A1(n29142), .A2(n19035), .Z(n2978) );
  XOR2_X1 U15424 ( .A1(n38222), .A2(n31548), .Z(n2979) );
  XOR2_X1 U15426 ( .A1(n3649), .A2(n8447), .Z(n3651) );
  NAND2_X2 U15428 ( .A1(n18571), .A2(n20410), .ZN(n3014) );
  XOR2_X1 U15430 ( .A1(n22699), .A2(n39136), .Z(n18834) );
  XOR2_X1 U15432 ( .A1(n2988), .A2(n2985), .Z(n20874) );
  XOR2_X1 U15433 ( .A1(n2986), .A2(n3953), .Z(n2985) );
  NAND2_X2 U15434 ( .A1(n2987), .A2(n3954), .ZN(n3953) );
  AND2_X1 U15435 ( .A1(n22198), .A2(n22199), .Z(n2987) );
  NAND2_X2 U15439 ( .A1(n5006), .A2(n2991), .ZN(n7497) );
  XOR2_X1 U15444 ( .A1(n28889), .A2(n5862), .Z(n29162) );
  XOR2_X1 U15445 ( .A1(n29164), .A2(n29163), .Z(n2996) );
  XOR2_X1 U15450 ( .A1(n12114), .A2(n12111), .Z(n7742) );
  NAND2_X2 U15451 ( .A1(n15801), .A2(n15804), .ZN(n3003) );
  NOR2_X1 U15465 ( .A1(n22022), .A2(n39010), .ZN(n22023) );
  XOR2_X1 U15466 ( .A1(n22661), .A2(n18888), .Z(n3022) );
  XOR2_X1 U15469 ( .A1(n15311), .A2(n11908), .Z(n3023) );
  OAI21_X2 U15474 ( .A1(n3464), .A2(n29059), .B(n3463), .ZN(n3462) );
  INV_X2 U15476 ( .I(n3027), .ZN(n22895) );
  NAND2_X1 U15477 ( .A1(n16104), .A2(n20174), .ZN(n22884) );
  XNOR2_X1 U15479 ( .A1(n35220), .A2(n38201), .ZN(n14563) );
  XOR2_X1 U15489 ( .A1(n3036), .A2(n3037), .Z(n3035) );
  XOR2_X1 U15490 ( .A1(n38844), .A2(n1704), .Z(n3036) );
  XOR2_X1 U15491 ( .A1(n26594), .A2(n10221), .Z(n3037) );
  NAND2_X1 U15497 ( .A1(n3045), .A2(n39828), .ZN(n3599) );
  XOR2_X1 U15506 ( .A1(n3060), .A2(n38189), .Z(n29169) );
  XOR2_X1 U15507 ( .A1(n3082), .A2(n29300), .Z(n3060) );
  OAI21_X2 U15514 ( .A1(n3072), .A2(n1000), .B(n3071), .ZN(n27663) );
  AOI21_X1 U15516 ( .A1(n34952), .A2(n3313), .B(n32557), .ZN(n3072) );
  XOR2_X1 U15525 ( .A1(n10638), .A2(n10635), .Z(n12480) );
  OAI21_X2 U15532 ( .A1(n17531), .A2(n22182), .B(n3085), .ZN(n16487) );
  XOR2_X1 U15537 ( .A1(n27785), .A2(n29785), .Z(n3090) );
  NOR2_X1 U15542 ( .A1(n18257), .A2(n3096), .ZN(n20963) );
  XOR2_X1 U15551 ( .A1(n26194), .A2(n26360), .Z(n4022) );
  XOR2_X1 U15554 ( .A1(n12282), .A2(n3105), .Z(n7708) );
  XOR2_X1 U15555 ( .A1(n22476), .A2(n19866), .Z(n3105) );
  OAI22_X2 U15557 ( .A1(n8549), .A2(n3107), .B1(n8552), .B2(n3106), .ZN(n12282) );
  AOI21_X1 U15564 ( .A1(n37093), .A2(n31944), .B(n38173), .ZN(n20809) );
  NOR2_X1 U15565 ( .A1(n1642), .A2(n37093), .ZN(n15519) );
  NOR2_X1 U15566 ( .A1(n1633), .A2(n37093), .ZN(n21251) );
  AOI22_X1 U15572 ( .A1(n28708), .A2(n16108), .B1(n18369), .B2(n28716), .ZN(
        n3128) );
  OAI21_X2 U15573 ( .A1(n27458), .A2(n36609), .B(n3129), .ZN(n28943) );
  INV_X2 U15575 ( .I(n5410), .ZN(n20313) );
  INV_X2 U15576 ( .I(n3134), .ZN(n26837) );
  INV_X2 U15581 ( .I(n16102), .ZN(n18261) );
  XOR2_X1 U15587 ( .A1(n791), .A2(n3141), .Z(n24427) );
  XOR2_X1 U15592 ( .A1(n38584), .A2(n33515), .Z(n3150) );
  XOR2_X1 U15594 ( .A1(n26595), .A2(n18004), .Z(n3152) );
  AND2_X1 U15599 ( .A1(n5736), .A2(n29182), .Z(n3155) );
  OR2_X1 U15600 ( .A1(n775), .A2(n4095), .Z(n3156) );
  NAND2_X2 U15615 ( .A1(n25441), .A2(n25440), .ZN(n18051) );
  NAND3_X2 U15621 ( .A1(n28173), .A2(n18192), .A3(n3164), .ZN(n28673) );
  XOR2_X1 U15626 ( .A1(n16523), .A2(n19991), .Z(n3166) );
  XOR2_X1 U15629 ( .A1(n22729), .A2(n29671), .Z(n3172) );
  XOR2_X1 U15639 ( .A1(n27664), .A2(n27663), .Z(n27835) );
  OAI22_X1 U15642 ( .A1(n21826), .A2(n34407), .B1(n21827), .B2(n3181), .ZN(
        n21828) );
  INV_X2 U15644 ( .I(n21187), .ZN(n18104) );
  XOR2_X1 U15647 ( .A1(n14639), .A2(n25035), .Z(n3186) );
  XOR2_X1 U15649 ( .A1(n15531), .A2(n20069), .Z(n3188) );
  XOR2_X1 U15661 ( .A1(n6560), .A2(n35196), .Z(n5915) );
  XOR2_X1 U15662 ( .A1(n6560), .A2(n23902), .Z(n14230) );
  MUX2_X1 U15664 ( .I0(n1069), .I1(n989), .S(n28023), .Z(n3199) );
  OAI21_X1 U15666 ( .A1(n1042), .A2(n33817), .B(n3200), .ZN(n17202) );
  XOR2_X1 U15671 ( .A1(n13035), .A2(n27839), .Z(n3206) );
  XOR2_X1 U15675 ( .A1(n27581), .A2(n27580), .Z(n27837) );
  XOR2_X1 U15677 ( .A1(n39093), .A2(n35200), .Z(n18106) );
  XOR2_X1 U15678 ( .A1(n39093), .A2(n12838), .Z(n10920) );
  NAND3_X2 U15680 ( .A1(n24964), .A2(n3214), .A3(n16785), .ZN(n25274) );
  OAI22_X1 U15681 ( .A1(n3215), .A2(n2277), .B1(n21479), .B2(n18576), .ZN(
        n21481) );
  AOI21_X1 U15682 ( .A1(n1349), .A2(n3215), .B(n21820), .ZN(n21480) );
  NAND3_X1 U15683 ( .A1(n6844), .A2(n6845), .A3(n1377), .ZN(n3217) );
  XOR2_X1 U15685 ( .A1(n35654), .A2(n29983), .Z(n17363) );
  XOR2_X1 U15688 ( .A1(n35867), .A2(n29269), .Z(n3223) );
  XOR2_X1 U15692 ( .A1(n3229), .A2(n4235), .Z(n25636) );
  NAND2_X2 U15694 ( .A1(n8096), .A2(n25358), .ZN(n9743) );
  NOR2_X2 U15696 ( .A1(n5592), .A2(n23313), .ZN(n6561) );
  NAND2_X1 U15699 ( .A1(n13539), .A2(n3235), .ZN(n28146) );
  OAI21_X2 U15702 ( .A1(n1663), .A2(n4139), .B(n3237), .ZN(n22663) );
  XOR2_X1 U15707 ( .A1(n22663), .A2(n8136), .Z(n3240) );
  XOR2_X1 U15708 ( .A1(n3242), .A2(n10718), .Z(n3241) );
  XOR2_X1 U15709 ( .A1(n33690), .A2(n31620), .Z(n3242) );
  AOI21_X2 U15710 ( .A1(n12375), .A2(n16041), .B(n12374), .ZN(n10621) );
  NOR2_X2 U15715 ( .A1(n23468), .A2(n3256), .ZN(n23635) );
  XOR2_X1 U15723 ( .A1(n3262), .A2(n27819), .Z(n3261) );
  NOR2_X2 U15724 ( .A1(n27489), .A2(n27488), .ZN(n27819) );
  XOR2_X1 U15725 ( .A1(n19642), .A2(n1160), .Z(n3262) );
  NAND3_X1 U15727 ( .A1(n29236), .A2(n3263), .A3(n8728), .ZN(n29234) );
  OAI22_X1 U15729 ( .A1(n14198), .A2(n3263), .B1(n14199), .B2(n29231), .ZN(
        n14197) );
  NAND2_X1 U15730 ( .A1(n29230), .A2(n3263), .ZN(n15026) );
  OAI22_X2 U15735 ( .A1(n3271), .A2(n21810), .B1(n3270), .B2(n19470), .ZN(
        n21214) );
  XOR2_X1 U15739 ( .A1(n28852), .A2(n3280), .Z(n29023) );
  XOR2_X1 U15741 ( .A1(n3280), .A2(n1374), .Z(n29250) );
  XOR2_X1 U15742 ( .A1(n3280), .A2(n13639), .Z(n5648) );
  INV_X2 U15747 ( .I(n14060), .ZN(n19914) );
  XOR2_X1 U15751 ( .A1(n3284), .A2(n14969), .Z(Ciphertext[24]) );
  NAND2_X1 U15754 ( .A1(n3288), .A2(n29333), .ZN(n3287) );
  XOR2_X1 U15757 ( .A1(n26393), .A2(n11057), .Z(n3290) );
  XOR2_X1 U15758 ( .A1(n26421), .A2(n26436), .Z(n11057) );
  XOR2_X1 U15774 ( .A1(n7287), .A2(n38920), .Z(n3301) );
  XOR2_X1 U15775 ( .A1(n12437), .A2(n22775), .Z(n3303) );
  XOR2_X1 U15776 ( .A1(n3305), .A2(n16131), .Z(n3304) );
  XOR2_X1 U15777 ( .A1(n15513), .A2(n4139), .Z(n3305) );
  AOI22_X1 U15783 ( .A1(n3312), .A2(n13754), .B1(n27282), .B2(n3313), .ZN(
        n17697) );
  NOR2_X1 U15784 ( .A1(n1227), .A2(n3313), .ZN(n3312) );
  NAND2_X2 U15786 ( .A1(n16147), .A2(n9008), .ZN(n20333) );
  XOR2_X1 U15789 ( .A1(n5820), .A2(n23964), .Z(n3316) );
  XOR2_X1 U15797 ( .A1(n26311), .A2(n26232), .Z(n3331) );
  OAI21_X1 U15798 ( .A1(n21574), .A2(n3337), .B(n21571), .ZN(n20581) );
  INV_X1 U15800 ( .I(n29023), .ZN(n3342) );
  INV_X2 U15801 ( .I(n14834), .ZN(n13153) );
  XOR2_X1 U15808 ( .A1(n11739), .A2(n19879), .Z(n3346) );
  INV_X1 U15810 ( .I(n8705), .ZN(n3352) );
  OAI21_X2 U15822 ( .A1(n23318), .A2(n23589), .B(n3364), .ZN(n23883) );
  OAI21_X1 U15829 ( .A1(n34177), .A2(n30141), .B(n18588), .ZN(n3373) );
  XOR2_X1 U15831 ( .A1(n23835), .A2(n16781), .Z(n3375) );
  NAND2_X1 U15834 ( .A1(n6843), .A2(n29278), .ZN(n6841) );
  NOR3_X1 U15842 ( .A1(n34813), .A2(n19873), .A3(n22349), .ZN(n22388) );
  XOR2_X1 U15846 ( .A1(n57), .A2(n1163), .Z(n3387) );
  NAND2_X1 U15847 ( .A1(n26666), .A2(n3388), .ZN(n9646) );
  NAND2_X1 U15848 ( .A1(n11523), .A2(n3388), .ZN(n11522) );
  XOR2_X1 U15849 ( .A1(n3604), .A2(n8874), .Z(n8741) );
  AOI21_X2 U15873 ( .A1(n3412), .A2(n36662), .B(n3409), .ZN(n13733) );
  MUX2_X1 U15875 ( .I0(n19698), .I1(n4846), .S(n13042), .Z(n3412) );
  AOI21_X2 U15878 ( .A1(n25955), .A2(n365), .B(n9589), .ZN(n4828) );
  XOR2_X1 U15880 ( .A1(n32190), .A2(n18279), .Z(n13025) );
  XOR2_X1 U15881 ( .A1(n23832), .A2(n32190), .Z(n13102) );
  XOR2_X1 U15886 ( .A1(n29098), .A2(n3127), .Z(n29100) );
  XOR2_X1 U15892 ( .A1(Plaintext[187]), .A2(Key[187]), .Z(n3443) );
  XOR2_X1 U15896 ( .A1(n8885), .A2(n26247), .Z(n3422) );
  INV_X2 U15897 ( .I(n14122), .ZN(n17709) );
  XOR2_X1 U15902 ( .A1(n3424), .A2(n7329), .Z(n15051) );
  NAND2_X2 U15911 ( .A1(n6214), .A2(n14654), .ZN(n17658) );
  INV_X2 U15916 ( .I(n3445), .ZN(n5988) );
  XNOR2_X1 U15917 ( .A1(n3446), .A2(n3603), .ZN(n3445) );
  XOR2_X1 U15919 ( .A1(n27749), .A2(n9981), .Z(n3447) );
  NAND2_X2 U15922 ( .A1(n12269), .A2(n12268), .ZN(n3448) );
  INV_X1 U15924 ( .I(Plaintext[191]), .ZN(n3450) );
  XOR2_X1 U15925 ( .A1(n3450), .A2(Key[191]), .Z(n3507) );
  NAND2_X1 U15926 ( .A1(n3452), .A2(n17464), .ZN(n23003) );
  XOR2_X1 U15933 ( .A1(n3458), .A2(n3457), .Z(n3456) );
  XOR2_X1 U15934 ( .A1(n34768), .A2(n3413), .Z(n3457) );
  XOR2_X1 U15935 ( .A1(n1009), .A2(n26480), .Z(n3458) );
  XOR2_X1 U15940 ( .A1(n3473), .A2(n3472), .Z(n3471) );
  XOR2_X1 U15941 ( .A1(n27796), .A2(n37112), .Z(n3472) );
  XOR2_X1 U15942 ( .A1(n27633), .A2(n8059), .Z(n3473) );
  MUX2_X1 U15953 ( .I0(n19322), .I1(n28571), .S(n31513), .Z(n28573) );
  AOI21_X1 U15954 ( .A1(n37938), .A2(n18854), .B(n35290), .ZN(n18952) );
  INV_X2 U15958 ( .I(n3486), .ZN(n17993) );
  NAND2_X1 U15961 ( .A1(n3760), .A2(n30464), .ZN(n5401) );
  XOR2_X1 U15964 ( .A1(n17399), .A2(n3488), .Z(n3489) );
  XOR2_X1 U15965 ( .A1(n29047), .A2(n29046), .Z(n3490) );
  XOR2_X1 U15970 ( .A1(n25240), .A2(n19947), .Z(n3493) );
  NAND2_X2 U15979 ( .A1(n23433), .A2(n23431), .ZN(n23624) );
  NAND2_X2 U15981 ( .A1(n23434), .A2(n23432), .ZN(n7335) );
  INV_X2 U15982 ( .I(n3507), .ZN(n4116) );
  NAND2_X1 U15986 ( .A1(n24909), .A2(n3510), .ZN(n24729) );
  NAND3_X2 U15992 ( .A1(n26579), .A2(n26580), .A3(n26581), .ZN(n5831) );
  AND2_X1 U15995 ( .A1(n26116), .A2(n30302), .Z(n3517) );
  XOR2_X1 U15996 ( .A1(n3521), .A2(n19897), .Z(n6781) );
  XOR2_X1 U15998 ( .A1(n3521), .A2(n19902), .Z(n23995) );
  XOR2_X1 U15999 ( .A1(n3521), .A2(n19887), .Z(n15862) );
  XOR2_X1 U16003 ( .A1(n3523), .A2(n25003), .Z(n3522) );
  XOR2_X1 U16004 ( .A1(n33038), .A2(n31891), .Z(n3523) );
  XNOR2_X1 U16005 ( .A1(n38581), .A2(n25115), .ZN(n25003) );
  XOR2_X1 U16006 ( .A1(n24970), .A2(n4015), .Z(n3525) );
  OAI21_X2 U16009 ( .A1(n33861), .A2(n30196), .B(n37083), .ZN(n3527) );
  INV_X4 U16011 ( .I(n20405), .ZN(n30196) );
  NOR2_X1 U16015 ( .A1(n34014), .A2(n3273), .ZN(n3546) );
  INV_X1 U16016 ( .I(n13688), .ZN(n3547) );
  XOR2_X1 U16017 ( .A1(n6635), .A2(n3549), .Z(n3548) );
  XOR2_X1 U16018 ( .A1(n29165), .A2(n35249), .Z(n3549) );
  XOR2_X1 U16020 ( .A1(n3552), .A2(n3551), .Z(n3550) );
  XOR2_X1 U16023 ( .A1(n26363), .A2(n3554), .Z(n3553) );
  XOR2_X1 U16024 ( .A1(n18012), .A2(n39082), .Z(n3554) );
  XOR2_X1 U16025 ( .A1(n26587), .A2(n26387), .Z(n26363) );
  NAND2_X2 U16026 ( .A1(n3555), .A2(n26011), .ZN(n26387) );
  NOR2_X2 U16027 ( .A1(n7517), .A2(n26017), .ZN(n26587) );
  XOR2_X1 U16041 ( .A1(Plaintext[99]), .A2(Key[99]), .Z(n3839) );
  XOR2_X1 U16042 ( .A1(Key[101]), .A2(Plaintext[101]), .Z(n7696) );
  INV_X2 U16043 ( .I(n10629), .ZN(n21870) );
  NOR2_X1 U16059 ( .A1(n6390), .A2(n3575), .ZN(n6179) );
  OAI21_X2 U16065 ( .A1(n24209), .A2(n326), .B(n23816), .ZN(n8646) );
  AOI21_X1 U16069 ( .A1(n17618), .A2(n8646), .B(n7529), .ZN(n23824) );
  XOR2_X1 U16072 ( .A1(n25269), .A2(n449), .Z(n3576) );
  XOR2_X1 U16073 ( .A1(n6778), .A2(n3578), .Z(n3577) );
  XOR2_X1 U16074 ( .A1(n25115), .A2(n24944), .Z(n3578) );
  XOR2_X1 U16077 ( .A1(n3585), .A2(n3584), .Z(n8765) );
  XOR2_X1 U16078 ( .A1(n4301), .A2(n698), .Z(n3584) );
  NAND2_X1 U16087 ( .A1(n23529), .A2(n31685), .ZN(n6611) );
  NOR2_X1 U16089 ( .A1(n18883), .A2(n28578), .ZN(n14516) );
  XOR2_X1 U16096 ( .A1(n3601), .A2(n19534), .Z(n23984) );
  XOR2_X1 U16097 ( .A1(n39014), .A2(n19674), .Z(n23809) );
  XOR2_X1 U16098 ( .A1(n39014), .A2(n19903), .Z(n23842) );
  XOR2_X1 U16104 ( .A1(n3604), .A2(n27750), .Z(n3603) );
  NAND2_X1 U16107 ( .A1(n35427), .A2(n11820), .ZN(n18488) );
  NOR2_X1 U16110 ( .A1(n3606), .A2(n13393), .ZN(n17024) );
  NAND2_X1 U16111 ( .A1(n26897), .A2(n3606), .ZN(n9203) );
  XOR2_X1 U16114 ( .A1(n3609), .A2(n19816), .Z(n13023) );
  XOR2_X1 U16115 ( .A1(n3609), .A2(n19843), .Z(n23759) );
  XOR2_X1 U16116 ( .A1(n16858), .A2(n34844), .Z(n24015) );
  XOR2_X1 U16117 ( .A1(n2585), .A2(n29017), .Z(n22690) );
  XOR2_X1 U16120 ( .A1(n23931), .A2(n23609), .Z(n3616) );
  XOR2_X1 U16126 ( .A1(n3621), .A2(n13845), .Z(n8694) );
  XOR2_X1 U16128 ( .A1(n22634), .A2(n3623), .Z(n3622) );
  OAI21_X2 U16134 ( .A1(n3627), .A2(n3626), .B(n33821), .ZN(n17904) );
  XOR2_X1 U16135 ( .A1(n17907), .A2(n17909), .Z(n3952) );
  INV_X2 U16136 ( .I(n20482), .ZN(n22795) );
  XOR2_X1 U16139 ( .A1(n28836), .A2(n665), .Z(n3632) );
  INV_X2 U16141 ( .I(n11784), .ZN(n8527) );
  XOR2_X1 U16143 ( .A1(n3639), .A2(n13154), .Z(n3638) );
  XOR2_X1 U16145 ( .A1(n26437), .A2(n1506), .Z(n3641) );
  NAND2_X1 U16147 ( .A1(n8393), .A2(n3642), .ZN(n8392) );
  XNOR2_X1 U16152 ( .A1(n19156), .A2(n25030), .ZN(n25201) );
  XOR2_X1 U16158 ( .A1(n3657), .A2(n3651), .Z(n3650) );
  XOR2_X1 U16159 ( .A1(n3656), .A2(n25043), .Z(n3652) );
  XOR2_X1 U16160 ( .A1(n39541), .A2(n19874), .Z(n3656) );
  XOR2_X1 U16162 ( .A1(n26403), .A2(n18432), .Z(n15717) );
  NAND2_X1 U16172 ( .A1(n28654), .A2(n3664), .ZN(n28443) );
  XOR2_X1 U16174 ( .A1(n39798), .A2(n29165), .Z(n3666) );
  XOR2_X1 U16184 ( .A1(n38816), .A2(n29514), .Z(n16606) );
  INV_X2 U16186 ( .I(n3675), .ZN(n4947) );
  XOR2_X1 U16187 ( .A1(n1664), .A2(n22604), .Z(n4270) );
  NAND2_X2 U16188 ( .A1(n3679), .A2(n3677), .ZN(n10488) );
  XOR2_X1 U16189 ( .A1(n7848), .A2(n28610), .Z(n28959) );
  OAI21_X1 U16197 ( .A1(n13900), .A2(n11684), .B(n3687), .ZN(n11683) );
  NOR2_X1 U16200 ( .A1(n15996), .A2(n3694), .ZN(n20882) );
  XNOR2_X1 U16203 ( .A1(n22635), .A2(n22619), .ZN(n3695) );
  XOR2_X1 U16204 ( .A1(n19819), .A2(n13564), .Z(n22619) );
  XOR2_X1 U16206 ( .A1(n22760), .A2(n8890), .Z(n3696) );
  NAND2_X1 U16211 ( .A1(n4449), .A2(n3700), .ZN(n4448) );
  XOR2_X1 U16213 ( .A1(n10382), .A2(n14648), .Z(n3701) );
  NOR2_X2 U16222 ( .A1(n18364), .A2(n28518), .ZN(n29042) );
  XOR2_X1 U16225 ( .A1(n9776), .A2(n3711), .Z(n3710) );
  XOR2_X1 U16228 ( .A1(n13155), .A2(n38979), .Z(n3712) );
  INV_X1 U16232 ( .I(n30076), .ZN(n30081) );
  NOR2_X1 U16233 ( .A1(n20078), .A2(n30076), .ZN(n30060) );
  NOR2_X2 U16235 ( .A1(n23567), .A2(n23566), .ZN(n3715) );
  NOR2_X1 U16238 ( .A1(n29856), .A2(n3725), .ZN(n14160) );
  XOR2_X1 U16241 ( .A1(n27497), .A2(n3727), .Z(n3726) );
  XOR2_X1 U16242 ( .A1(n27672), .A2(n28831), .Z(n3727) );
  XOR2_X1 U16244 ( .A1(n34829), .A2(n27556), .Z(n27673) );
  XOR2_X1 U16248 ( .A1(n26487), .A2(n39129), .Z(n3731) );
  NOR2_X1 U16256 ( .A1(n19863), .A2(n25498), .ZN(n3736) );
  XOR2_X1 U16259 ( .A1(n25163), .A2(n25096), .Z(n24987) );
  XOR2_X1 U16260 ( .A1(n25163), .A2(n1369), .Z(n14687) );
  XOR2_X1 U16263 ( .A1(n23938), .A2(n9518), .Z(n23387) );
  XOR2_X1 U16267 ( .A1(n12101), .A2(n12282), .Z(n3747) );
  XOR2_X1 U16269 ( .A1(n17651), .A2(n22782), .Z(n3748) );
  OAI21_X2 U16270 ( .A1(n3751), .A2(n24731), .B(n3749), .ZN(n15186) );
  XOR2_X1 U16279 ( .A1(n26522), .A2(n3769), .Z(n4412) );
  XOR2_X1 U16280 ( .A1(n291), .A2(n1723), .Z(n3769) );
  INV_X2 U16285 ( .I(n3770), .ZN(n16363) );
  INV_X2 U16286 ( .I(n3771), .ZN(n4945) );
  INV_X2 U16293 ( .I(n31775), .ZN(n3917) );
  XOR2_X1 U16297 ( .A1(n35320), .A2(n14307), .Z(n3776) );
  XOR2_X1 U16298 ( .A1(n8585), .A2(n30324), .Z(n3777) );
  XOR2_X1 U16299 ( .A1(n38495), .A2(n35251), .Z(n3778) );
  NAND2_X1 U16301 ( .A1(n2302), .A2(n3779), .ZN(n12486) );
  XOR2_X1 U16302 ( .A1(n3780), .A2(n3782), .Z(n19436) );
  NAND2_X2 U16304 ( .A1(n25795), .A2(n25794), .ZN(n26396) );
  NAND2_X2 U16306 ( .A1(n14145), .A2(n25938), .ZN(n12649) );
  XOR2_X1 U16307 ( .A1(n26497), .A2(n30471), .Z(n3782) );
  XOR2_X1 U16315 ( .A1(n33310), .A2(n19925), .Z(n3787) );
  XOR2_X1 U16319 ( .A1(n33584), .A2(n1215), .Z(n3790) );
  XOR2_X1 U16320 ( .A1(n27845), .A2(n31551), .Z(n3791) );
  NOR2_X1 U16325 ( .A1(n28622), .A2(n9917), .ZN(n3799) );
  XOR2_X1 U16326 ( .A1(n3800), .A2(n3801), .Z(n12770) );
  XOR2_X1 U16328 ( .A1(n22689), .A2(n22410), .Z(n3801) );
  NAND2_X2 U16330 ( .A1(n17155), .A2(n17154), .ZN(n22775) );
  INV_X2 U16331 ( .I(n26265), .ZN(n10440) );
  XOR2_X1 U16337 ( .A1(n5086), .A2(n3804), .Z(n6331) );
  INV_X1 U16349 ( .I(n10029), .ZN(n3826) );
  XOR2_X1 U16352 ( .A1(n15581), .A2(n14969), .Z(n11882) );
  OAI21_X1 U16353 ( .A1(n22299), .A2(n22073), .B(n22038), .ZN(n3833) );
  NAND2_X2 U16354 ( .A1(n33886), .A2(n4388), .ZN(n22304) );
  NAND2_X1 U16359 ( .A1(n39098), .A2(n24764), .ZN(n6038) );
  AOI21_X1 U16362 ( .A1(n36186), .A2(n39098), .B(n5896), .ZN(n8579) );
  OAI21_X1 U16364 ( .A1(n1269), .A2(n39098), .B(n4008), .ZN(n7242) );
  INV_X2 U16371 ( .I(n3852), .ZN(n8805) );
  NOR2_X2 U16373 ( .A1(n9016), .A2(n10712), .ZN(n11923) );
  XOR2_X1 U16377 ( .A1(n39698), .A2(n38160), .Z(n3855) );
  OR2_X1 U16380 ( .A1(n3951), .A2(n29182), .Z(n3857) );
  XOR2_X1 U16381 ( .A1(n26408), .A2(n26409), .Z(n3858) );
  NOR2_X1 U16383 ( .A1(n3860), .A2(n31570), .ZN(n18083) );
  NAND2_X1 U16384 ( .A1(n3860), .A2(n39709), .ZN(n29913) );
  OAI21_X1 U16387 ( .A1(n12439), .A2(n7278), .B(n3868), .ZN(n3867) );
  XOR2_X1 U16391 ( .A1(n3929), .A2(n7783), .Z(n3872) );
  AND2_X1 U16396 ( .A1(n19005), .A2(n23381), .Z(n3884) );
  XOR2_X1 U16406 ( .A1(n31620), .A2(n38154), .Z(n3891) );
  XOR2_X1 U16409 ( .A1(n3895), .A2(n3894), .Z(n3893) );
  XOR2_X1 U16410 ( .A1(n9325), .A2(n9324), .Z(n3894) );
  XOR2_X1 U16411 ( .A1(n15186), .A2(n37357), .Z(n3895) );
  NAND2_X2 U16413 ( .A1(n28014), .A2(n28013), .ZN(n28570) );
  XOR2_X1 U16418 ( .A1(n23780), .A2(n3917), .Z(n6628) );
  NAND2_X1 U16432 ( .A1(n9711), .A2(n39489), .ZN(n3930) );
  MUX2_X1 U16433 ( .I0(n6361), .I1(n22069), .S(n22327), .Z(n20090) );
  AOI21_X2 U16446 ( .A1(n14971), .A2(n17190), .B(n28754), .ZN(n28852) );
  XOR2_X1 U16447 ( .A1(n28943), .A2(n19845), .Z(n3941) );
  NOR2_X2 U16449 ( .A1(n34016), .A2(n6241), .ZN(n10961) );
  XNOR2_X1 U16454 ( .A1(n25179), .A2(n20707), .ZN(n14644) );
  XOR2_X1 U16457 ( .A1(n20212), .A2(n11057), .Z(n3956) );
  XOR2_X1 U16461 ( .A1(n2711), .A2(n4258), .Z(n4257) );
  XOR2_X1 U16462 ( .A1(n10653), .A2(n21121), .Z(n18893) );
  XOR2_X1 U16464 ( .A1(n27535), .A2(n10653), .Z(n9732) );
  INV_X2 U16470 ( .I(n3973), .ZN(n19615) );
  XOR2_X1 U16473 ( .A1(n11399), .A2(n14293), .Z(n3975) );
  XOR2_X1 U16479 ( .A1(n4273), .A2(n816), .Z(n16203) );
  INV_X2 U16485 ( .I(n28174), .ZN(n28258) );
  XOR2_X1 U16494 ( .A1(n8785), .A2(n22505), .Z(n4000) );
  NOR2_X2 U16495 ( .A1(n7041), .A2(n7042), .ZN(n4117) );
  XOR2_X1 U16498 ( .A1(n654), .A2(n27628), .Z(n4009) );
  OR2_X1 U16500 ( .A1(n9334), .A2(n4413), .Z(n4010) );
  NAND3_X2 U16502 ( .A1(n11921), .A2(n22217), .A3(n22218), .ZN(n22615) );
  XOR2_X1 U16506 ( .A1(n25301), .A2(n29432), .Z(n4015) );
  INV_X2 U16507 ( .I(n4016), .ZN(n22920) );
  XOR2_X1 U16508 ( .A1(n14106), .A2(n7593), .Z(n15331) );
  XOR2_X1 U16514 ( .A1(n33308), .A2(n2150), .Z(n4021) );
  XOR2_X1 U16518 ( .A1(n5848), .A2(n39652), .Z(n4039) );
  XOR2_X1 U16520 ( .A1(n29303), .A2(n29934), .Z(n4041) );
  INV_X2 U16528 ( .I(n17084), .ZN(n24360) );
  XOR2_X1 U16538 ( .A1(n25330), .A2(n18898), .Z(n4061) );
  XOR2_X1 U16542 ( .A1(n4066), .A2(n4065), .Z(n4064) );
  XOR2_X1 U16543 ( .A1(n27525), .A2(n30207), .Z(n4065) );
  XOR2_X1 U16544 ( .A1(n33584), .A2(n27663), .Z(n4066) );
  XOR2_X1 U16554 ( .A1(n792), .A2(n23940), .Z(n4070) );
  OAI21_X2 U16559 ( .A1(n4429), .A2(n4428), .B(n4076), .ZN(n18362) );
  XOR2_X1 U16562 ( .A1(n39637), .A2(n1357), .Z(n4079) );
  XOR2_X1 U16563 ( .A1(n26571), .A2(n8585), .Z(n4080) );
  XOR2_X1 U16569 ( .A1(n22625), .A2(n22650), .Z(n4085) );
  NOR2_X2 U16573 ( .A1(n10025), .A2(n20042), .ZN(n19221) );
  XOR2_X1 U16580 ( .A1(n32349), .A2(n4092), .Z(n4091) );
  XOR2_X1 U16582 ( .A1(n5026), .A2(n24923), .Z(n4090) );
  XOR2_X1 U16585 ( .A1(n7352), .A2(n15186), .Z(n4092) );
  NOR2_X2 U16586 ( .A1(n23148), .A2(n23147), .ZN(n23560) );
  AOI22_X1 U16588 ( .A1(n19262), .A2(n4093), .B1(n21812), .B2(n4094), .ZN(
        n18825) );
  NOR2_X1 U16589 ( .A1(n19768), .A2(n4094), .ZN(n4093) );
  OR2_X1 U16591 ( .A1(n22871), .A2(n19293), .Z(n4100) );
  NOR2_X1 U16594 ( .A1(n38193), .A2(n27253), .ZN(n4104) );
  NAND2_X2 U16598 ( .A1(n4111), .A2(n4109), .ZN(n19152) );
  INV_X1 U16600 ( .I(n4108), .ZN(n4114) );
  XOR2_X1 U16603 ( .A1(n20586), .A2(n5185), .Z(n23565) );
  NOR2_X2 U16608 ( .A1(n21374), .A2(n21375), .ZN(n22131) );
  XOR2_X1 U16611 ( .A1(n8875), .A2(n38174), .Z(n27750) );
  XOR2_X1 U16619 ( .A1(n25202), .A2(n24918), .Z(n4129) );
  XOR2_X1 U16622 ( .A1(n5293), .A2(n718), .Z(n4131) );
  XOR2_X1 U16626 ( .A1(n35972), .A2(n19862), .Z(n4136) );
  INV_X2 U16627 ( .I(n4137), .ZN(n10414) );
  XOR2_X1 U16628 ( .A1(n4139), .A2(n1356), .Z(n4436) );
  XOR2_X1 U16629 ( .A1(n4441), .A2(n4139), .Z(n19956) );
  XOR2_X1 U16630 ( .A1(n28969), .A2(n29840), .Z(n4140) );
  XOR2_X1 U16632 ( .A1(n11997), .A2(n4142), .Z(n11996) );
  INV_X1 U16633 ( .I(n27828), .ZN(n4142) );
  NOR2_X1 U16654 ( .A1(n954), .A2(n728), .ZN(n5453) );
  NAND2_X2 U16659 ( .A1(n17142), .A2(n35500), .ZN(n27328) );
  MUX2_X1 U16662 ( .I0(n24378), .I1(n24377), .S(n8041), .Z(n4177) );
  NOR2_X1 U16671 ( .A1(n17217), .A2(n38377), .ZN(n4194) );
  XOR2_X1 U16677 ( .A1(n4201), .A2(n9027), .Z(n9026) );
  XOR2_X1 U16678 ( .A1(n4201), .A2(n11392), .Z(n6906) );
  XOR2_X1 U16683 ( .A1(n334), .A2(n10027), .Z(n4204) );
  XOR2_X1 U16685 ( .A1(n4205), .A2(n26477), .Z(n20536) );
  NOR2_X1 U16689 ( .A1(n35915), .A2(n31931), .ZN(n5723) );
  NAND3_X1 U16693 ( .A1(n1231), .A2(n33858), .A3(n4211), .ZN(n26964) );
  NAND2_X1 U16696 ( .A1(n25584), .A2(n25449), .ZN(n4214) );
  XOR2_X1 U16700 ( .A1(n38221), .A2(n4222), .Z(n4221) );
  XOR2_X1 U16701 ( .A1(n7710), .A2(n29325), .Z(n4222) );
  NAND2_X2 U16709 ( .A1(n13073), .A2(n13072), .ZN(n13966) );
  XOR2_X1 U16711 ( .A1(Plaintext[11]), .A2(Key[11]), .Z(n5131) );
  OAI21_X1 U16714 ( .A1(n18453), .A2(n4232), .B(n10544), .ZN(n18398) );
  NAND3_X1 U16715 ( .A1(n10544), .A2(n18453), .A3(n4232), .ZN(n17045) );
  XOR2_X1 U16720 ( .A1(n4237), .A2(n25276), .Z(n4235) );
  XOR2_X1 U16721 ( .A1(n18600), .A2(n25275), .Z(n4237) );
  XOR2_X1 U16731 ( .A1(n4256), .A2(n4257), .Z(n20995) );
  XOR2_X1 U16733 ( .A1(n19450), .A2(n19583), .Z(n4258) );
  XOR2_X1 U16741 ( .A1(n16096), .A2(n23591), .Z(n4268) );
  XOR2_X1 U16744 ( .A1(n20668), .A2(n4270), .Z(n4269) );
  XOR2_X1 U16745 ( .A1(n10525), .A2(n22525), .Z(n4271) );
  NAND2_X2 U16746 ( .A1(n22856), .A2(n17080), .ZN(n22923) );
  XOR2_X1 U16756 ( .A1(n22615), .A2(n29920), .Z(n4277) );
  XOR2_X1 U16757 ( .A1(n10558), .A2(n4493), .Z(n4278) );
  XOR2_X1 U16765 ( .A1(n14023), .A2(n9272), .Z(n4282) );
  NAND2_X1 U16768 ( .A1(n14927), .A2(n4283), .ZN(n14926) );
  NAND2_X2 U16769 ( .A1(n22315), .A2(n9616), .ZN(n4283) );
  NOR2_X1 U16771 ( .A1(n35911), .A2(n1414), .ZN(n17115) );
  MUX2_X1 U16772 ( .I0(n28113), .I1(n28112), .S(n1414), .Z(n28122) );
  NAND2_X1 U16773 ( .A1(n32796), .A2(n9677), .ZN(n22840) );
  NAND2_X1 U16775 ( .A1(n31601), .A2(n30096), .ZN(n18134) );
  NOR2_X1 U16777 ( .A1(n9543), .A2(n4294), .ZN(n13408) );
  NAND2_X1 U16778 ( .A1(n33431), .A2(n10334), .ZN(n4294) );
  INV_X2 U16779 ( .I(n4300), .ZN(n11496) );
  XOR2_X1 U16797 ( .A1(n29824), .A2(n29785), .Z(n4313) );
  XOR2_X1 U16798 ( .A1(n4314), .A2(n15157), .Z(n29129) );
  OR2_X1 U16806 ( .A1(n16999), .A2(n37067), .Z(n4321) );
  XOR2_X1 U16814 ( .A1(n4327), .A2(n12174), .Z(n4326) );
  NAND2_X2 U16815 ( .A1(n5946), .A2(n4328), .ZN(n4644) );
  OAI21_X1 U16816 ( .A1(n15230), .A2(n22833), .B(n11914), .ZN(n4329) );
  XOR2_X1 U16817 ( .A1(n21098), .A2(n18322), .Z(n4330) );
  XOR2_X1 U16819 ( .A1(n4332), .A2(n4334), .Z(n5050) );
  XOR2_X1 U16820 ( .A1(n24610), .A2(n4333), .Z(n4332) );
  XOR2_X1 U16821 ( .A1(n6066), .A2(n965), .Z(n4333) );
  XOR2_X1 U16823 ( .A1(n25254), .A2(n4335), .Z(n4334) );
  XOR2_X1 U16824 ( .A1(n38665), .A2(n32195), .Z(n4335) );
  NAND2_X1 U16826 ( .A1(n4340), .A2(n1648), .ZN(n20971) );
  INV_X2 U16830 ( .I(n4342), .ZN(n22335) );
  XOR2_X1 U16831 ( .A1(n32239), .A2(n19774), .Z(n23782) );
  XOR2_X1 U16836 ( .A1(n22624), .A2(n34239), .Z(n4346) );
  XOR2_X1 U16839 ( .A1(n5566), .A2(n5565), .Z(n5402) );
  INV_X2 U16840 ( .I(n4352), .ZN(n25601) );
  NAND2_X2 U16842 ( .A1(n19495), .A2(n25601), .ZN(n17613) );
  NAND3_X1 U16845 ( .A1(n27199), .A2(n13471), .A3(n4353), .ZN(n26915) );
  XOR2_X1 U16848 ( .A1(n29060), .A2(n4357), .Z(n4355) );
  INV_X2 U16850 ( .I(n4356), .ZN(n14559) );
  XOR2_X1 U16851 ( .A1(n15960), .A2(n30682), .Z(n4357) );
  NAND2_X2 U16860 ( .A1(n8169), .A2(n8168), .ZN(n9013) );
  OAI21_X1 U16862 ( .A1(n30181), .A2(n12198), .B(n4368), .ZN(n30182) );
  INV_X2 U16867 ( .I(n4386), .ZN(n30161) );
  NOR2_X1 U16875 ( .A1(n28458), .A2(n39423), .ZN(n28098) );
  XOR2_X1 U16877 ( .A1(n4399), .A2(n4398), .Z(n4397) );
  XOR2_X1 U16878 ( .A1(n19561), .A2(n17428), .Z(n4398) );
  XOR2_X1 U16879 ( .A1(n282), .A2(n27504), .Z(n4399) );
  INV_X2 U16885 ( .I(n4409), .ZN(n13605) );
  MUX2_X1 U16891 ( .I0(n4417), .I1(n788), .S(n1298), .Z(n4416) );
  NAND2_X2 U16895 ( .A1(n15982), .A2(n15985), .ZN(n27754) );
  AOI21_X1 U16898 ( .A1(n6938), .A2(n1399), .B(n19050), .ZN(n4423) );
  INV_X1 U16899 ( .I(n4424), .ZN(n15663) );
  NAND2_X1 U16901 ( .A1(n22063), .A2(n4424), .ZN(n16499) );
  XNOR2_X1 U16913 ( .A1(n26514), .A2(n26245), .ZN(n26287) );
  NAND2_X1 U16925 ( .A1(n13982), .A2(n4439), .ZN(n23513) );
  XOR2_X1 U16926 ( .A1(n4440), .A2(n4443), .Z(n4442) );
  XOR2_X1 U16927 ( .A1(n37699), .A2(n1707), .Z(n4443) );
  MUX2_X1 U16931 ( .I0(n28181), .I1(n36573), .S(n14397), .Z(n27742) );
  MUX2_X1 U16932 ( .I0(n1200), .I1(n1074), .S(n14397), .Z(n27904) );
  NOR2_X1 U16933 ( .A1(n4458), .A2(n2752), .ZN(n9014) );
  XOR2_X1 U16937 ( .A1(n38212), .A2(n1362), .Z(n15785) );
  INV_X1 U16939 ( .I(n4469), .ZN(n25645) );
  INV_X1 U16944 ( .I(n9155), .ZN(n8339) );
  INV_X2 U16945 ( .I(n12900), .ZN(n14561) );
  XOR2_X1 U16948 ( .A1(n4477), .A2(n1464), .Z(n4476) );
  XOR2_X1 U16949 ( .A1(n7106), .A2(n19825), .Z(n4477) );
  OAI21_X1 U16959 ( .A1(n30041), .A2(n30042), .B(n4498), .ZN(n8477) );
  XOR2_X1 U16961 ( .A1(n4499), .A2(n4501), .Z(n25722) );
  XOR2_X1 U16962 ( .A1(n25206), .A2(n4500), .Z(n4499) );
  XOR2_X1 U16963 ( .A1(n449), .A2(n30063), .Z(n4500) );
  XOR2_X1 U16964 ( .A1(n25301), .A2(n24984), .Z(n25206) );
  AOI21_X1 U16975 ( .A1(n9559), .A2(n1391), .B(n4518), .ZN(n18137) );
  OAI21_X1 U16976 ( .A1(n29318), .A2(n29333), .B(n4519), .ZN(n4518) );
  XOR2_X1 U16988 ( .A1(n36516), .A2(n12972), .Z(n23922) );
  NAND2_X1 U16989 ( .A1(n8416), .A2(n23414), .ZN(n4536) );
  XOR2_X1 U16991 ( .A1(n360), .A2(n9246), .Z(n4540) );
  XOR2_X1 U16994 ( .A1(n25046), .A2(n4549), .Z(n4551) );
  XOR2_X1 U16995 ( .A1(n16897), .A2(n31771), .Z(n4549) );
  XOR2_X1 U16997 ( .A1(n19967), .A2(n4552), .Z(n4550) );
  XOR2_X1 U16999 ( .A1(n1555), .A2(n3110), .Z(n4552) );
  NAND2_X2 U17002 ( .A1(n19258), .A2(n19257), .ZN(n4553) );
  XOR2_X1 U17008 ( .A1(n38850), .A2(n19534), .Z(n4558) );
  XOR2_X1 U17010 ( .A1(n22637), .A2(n31214), .Z(n4559) );
  XOR2_X1 U17014 ( .A1(n39310), .A2(n30104), .Z(n4561) );
  NAND2_X2 U17018 ( .A1(n5186), .A2(n16393), .ZN(n5185) );
  XOR2_X1 U17020 ( .A1(n4572), .A2(n10230), .Z(n9235) );
  NAND3_X2 U17023 ( .A1(n26104), .A2(n10234), .A3(n26105), .ZN(n26436) );
  XNOR2_X1 U17030 ( .A1(n778), .A2(n6308), .ZN(n4574) );
  XOR2_X1 U17037 ( .A1(n4591), .A2(n739), .Z(n4587) );
  XOR2_X1 U17038 ( .A1(n11667), .A2(n19516), .Z(n4589) );
  XOR2_X1 U17042 ( .A1(n4592), .A2(n23783), .Z(n15160) );
  XOR2_X1 U17052 ( .A1(n12838), .A2(n8585), .Z(n6526) );
  AOI21_X2 U17077 ( .A1(n4611), .A2(n20971), .B(n14544), .ZN(n23307) );
  NOR2_X2 U17084 ( .A1(n15915), .A2(n27111), .ZN(n27478) );
  INV_X1 U17095 ( .I(n19366), .ZN(n28147) );
  OR2_X1 U17099 ( .A1(n29687), .A2(n29678), .Z(n29673) );
  NAND2_X1 U17101 ( .A1(n5357), .A2(n23251), .ZN(n19358) );
  CLKBUF_X2 U17102 ( .I(Key[177]), .Z(n29887) );
  INV_X2 U17106 ( .I(n11782), .ZN(n20522) );
  OAI21_X1 U17111 ( .A1(n15246), .A2(n27506), .B(n15243), .ZN(n16861) );
  INV_X1 U17114 ( .I(n20546), .ZN(n7468) );
  NAND2_X1 U17119 ( .A1(n7303), .A2(n38200), .ZN(n4621) );
  NAND2_X2 U17124 ( .A1(n11141), .A2(n11143), .ZN(n12015) );
  OAI21_X2 U17128 ( .A1(n22224), .A2(n22166), .B(n13008), .ZN(n22485) );
  AND2_X1 U17129 ( .A1(n16261), .A2(n1208), .Z(n9850) );
  XOR2_X1 U17130 ( .A1(n29122), .A2(n29072), .Z(n28917) );
  NAND2_X1 U17133 ( .A1(n19060), .A2(n11067), .ZN(n4631) );
  OR2_X1 U17134 ( .A1(n27150), .A2(n27149), .Z(n27151) );
  INV_X2 U17139 ( .I(n4632), .ZN(n29643) );
  XOR2_X1 U17140 ( .A1(n27944), .A2(n4834), .Z(n4632) );
  INV_X1 U17141 ( .I(n22647), .ZN(n7056) );
  INV_X2 U17142 ( .I(n4633), .ZN(n20638) );
  XOR2_X1 U17143 ( .A1(n24935), .A2(n11698), .Z(n12181) );
  XNOR2_X1 U17149 ( .A1(n18765), .A2(n18764), .ZN(n5517) );
  OAI22_X1 U17150 ( .A1(n24720), .A2(n24719), .B1(n30764), .B2(n24723), .ZN(
        n24726) );
  XOR2_X1 U17151 ( .A1(n30179), .A2(n16017), .Z(n7548) );
  NAND3_X1 U17162 ( .A1(n20314), .A2(n28331), .A3(n29474), .ZN(n15005) );
  NAND2_X2 U17163 ( .A1(n10798), .A2(n10799), .ZN(n10667) );
  XOR2_X1 U17166 ( .A1(n5794), .A2(n23378), .Z(n5793) );
  XOR2_X1 U17171 ( .A1(n17552), .A2(n17553), .Z(n9748) );
  XOR2_X1 U17174 ( .A1(n27460), .A2(n1461), .Z(n4646) );
  INV_X1 U17179 ( .I(n19088), .ZN(n6862) );
  XOR2_X1 U17183 ( .A1(n5649), .A2(n5651), .Z(n28186) );
  XOR2_X1 U17184 ( .A1(n29085), .A2(n17832), .Z(n6855) );
  OAI21_X2 U17185 ( .A1(n6866), .A2(n17821), .B(n6865), .ZN(n16233) );
  XOR2_X1 U17197 ( .A1(n5889), .A2(n19186), .Z(n4658) );
  AND2_X1 U17199 ( .A1(n18077), .A2(n10004), .Z(n17332) );
  NOR2_X2 U17217 ( .A1(n4670), .A2(n10751), .ZN(n24492) );
  NOR2_X1 U17221 ( .A1(n26847), .A2(n26945), .ZN(n15669) );
  XOR2_X1 U17228 ( .A1(n9776), .A2(n26588), .Z(n4673) );
  NAND2_X1 U17238 ( .A1(n29946), .A2(n105), .ZN(n10146) );
  XNOR2_X1 U17239 ( .A1(n17937), .A2(n30114), .ZN(n14053) );
  XOR2_X1 U17246 ( .A1(n13235), .A2(n5861), .Z(n17461) );
  XNOR2_X1 U17262 ( .A1(n24525), .A2(n24524), .ZN(n7957) );
  OAI21_X1 U17268 ( .A1(n38173), .A2(n15519), .B(n23450), .ZN(n22913) );
  XOR2_X1 U17269 ( .A1(n23954), .A2(n23953), .Z(n11575) );
  NOR2_X2 U17277 ( .A1(n4704), .A2(n22885), .ZN(n23296) );
  XOR2_X1 U17278 ( .A1(n39739), .A2(n29857), .Z(n10040) );
  NAND2_X1 U17282 ( .A1(n22910), .A2(n10828), .ZN(n12697) );
  OR2_X1 U17292 ( .A1(n15320), .A2(n14471), .Z(n10937) );
  AOI21_X2 U17293 ( .A1(n1249), .A2(n20924), .B(n4715), .ZN(n25491) );
  OR2_X1 U17302 ( .A1(n15267), .A2(n9872), .Z(n20994) );
  OAI21_X1 U17316 ( .A1(n19686), .A2(n37757), .B(n9856), .ZN(n22823) );
  XOR2_X1 U17319 ( .A1(n9626), .A2(n29229), .Z(n4720) );
  INV_X1 U17325 ( .I(n5762), .ZN(n21324) );
  OR2_X1 U17327 ( .A1(n18815), .A2(n7295), .Z(n29187) );
  OR2_X1 U17334 ( .A1(n26634), .A2(n26905), .Z(n26579) );
  XOR2_X1 U17336 ( .A1(n8703), .A2(n10364), .Z(n5583) );
  AOI21_X1 U17337 ( .A1(n29527), .A2(n29526), .B(n4730), .ZN(n29529) );
  OR2_X1 U17340 ( .A1(n9177), .A2(n25022), .Z(n4736) );
  XOR2_X1 U17343 ( .A1(n19973), .A2(n26314), .Z(n9577) );
  XOR2_X1 U17346 ( .A1(n4738), .A2(n13680), .Z(n17918) );
  XOR2_X1 U17350 ( .A1(n36750), .A2(n19681), .Z(n15765) );
  INV_X2 U17356 ( .I(n21074), .ZN(n30042) );
  XOR2_X1 U17358 ( .A1(n4739), .A2(n1730), .Z(Ciphertext[123]) );
  NOR2_X1 U17371 ( .A1(n27904), .A2(n18832), .ZN(n13976) );
  NAND3_X1 U17377 ( .A1(n16630), .A2(n16628), .A3(n20499), .ZN(n7589) );
  XOR2_X1 U17380 ( .A1(n25072), .A2(n6410), .Z(n25270) );
  NAND2_X1 U17384 ( .A1(n13097), .A2(n26956), .ZN(n13096) );
  OR2_X1 U17402 ( .A1(n18168), .A2(n24768), .Z(n9418) );
  XOR2_X1 U17404 ( .A1(n4752), .A2(n27803), .Z(n15995) );
  NAND2_X1 U17421 ( .A1(n2910), .A2(n32107), .ZN(n7817) );
  NAND2_X2 U17422 ( .A1(n8578), .A2(n7971), .ZN(n25203) );
  XOR2_X1 U17433 ( .A1(n17138), .A2(n17139), .Z(n28179) );
  INV_X1 U17440 ( .I(n13018), .ZN(n20648) );
  AND2_X1 U17441 ( .A1(n25692), .A2(n12500), .Z(n5011) );
  NAND3_X2 U17450 ( .A1(n22972), .A2(n22970), .A3(n22971), .ZN(n17478) );
  XOR2_X1 U17468 ( .A1(n4780), .A2(n33515), .Z(Ciphertext[179]) );
  XOR2_X1 U17470 ( .A1(n9137), .A2(n779), .Z(n4899) );
  INV_X2 U17476 ( .I(n17064), .ZN(n20010) );
  OR2_X1 U17480 ( .A1(n16671), .A2(n24737), .Z(n14681) );
  INV_X2 U17481 ( .I(n4786), .ZN(n14417) );
  XOR2_X1 U17483 ( .A1(n13177), .A2(n16310), .Z(n13176) );
  NAND2_X2 U17489 ( .A1(n4897), .A2(n13905), .ZN(n15224) );
  XOR2_X1 U17493 ( .A1(n22454), .A2(n35590), .Z(n21134) );
  NAND2_X2 U17494 ( .A1(n8135), .A2(n16070), .ZN(n8585) );
  AND2_X1 U17499 ( .A1(n30162), .A2(n1400), .Z(n17842) );
  XOR2_X1 U17511 ( .A1(n6642), .A2(n9887), .Z(n6641) );
  NAND2_X2 U17512 ( .A1(n9053), .A2(n11605), .ZN(n14425) );
  NOR2_X1 U17513 ( .A1(n14618), .A2(n6643), .ZN(n13620) );
  AND2_X1 U17517 ( .A1(n3977), .A2(n3092), .Z(n11088) );
  INV_X1 U17530 ( .I(n29174), .ZN(n30046) );
  INV_X1 U17532 ( .I(n22346), .ZN(n13565) );
  NAND3_X1 U17537 ( .A1(n5110), .A2(n18708), .A3(n10074), .ZN(n16202) );
  OR2_X1 U17538 ( .A1(n25825), .A2(n18162), .Z(n25784) );
  XOR2_X1 U17542 ( .A1(n11779), .A2(n697), .Z(n11778) );
  NAND3_X2 U17551 ( .A1(n10056), .A2(n24598), .A3(n24599), .ZN(n24991) );
  XNOR2_X1 U17566 ( .A1(n1065), .A2(n29067), .ZN(n9054) );
  XNOR2_X1 U17569 ( .A1(n27942), .A2(n27943), .ZN(n4834) );
  AND2_X1 U17579 ( .A1(n25539), .A2(n30317), .Z(n12908) );
  NAND2_X1 U17584 ( .A1(n1120), .A2(n24764), .ZN(n9417) );
  INV_X2 U17590 ( .I(n4850), .ZN(n17424) );
  NAND3_X1 U17597 ( .A1(n28717), .A2(n28716), .A3(n16108), .ZN(n16505) );
  OR2_X1 U17598 ( .A1(n5044), .A2(n23542), .Z(n6235) );
  NAND3_X1 U17606 ( .A1(n13586), .A2(n26077), .A3(n9883), .ZN(n13585) );
  XOR2_X1 U17615 ( .A1(n35376), .A2(n23846), .Z(n10888) );
  NAND2_X2 U17616 ( .A1(n23279), .A2(n15562), .ZN(n23846) );
  AND2_X1 U17618 ( .A1(n906), .A2(n4862), .Z(n10018) );
  INV_X2 U17627 ( .I(n4866), .ZN(n17412) );
  XOR2_X1 U17628 ( .A1(n4869), .A2(n11960), .Z(n13827) );
  XOR2_X1 U17636 ( .A1(n4876), .A2(n16641), .Z(Ciphertext[82]) );
  NOR3_X1 U17637 ( .A1(n20443), .A2(n21032), .A3(n20444), .ZN(n4876) );
  XOR2_X1 U17649 ( .A1(n18843), .A2(n22694), .Z(n4883) );
  XOR2_X1 U17658 ( .A1(n17403), .A2(n17402), .Z(n14367) );
  AND2_X1 U17668 ( .A1(n21310), .A2(n19864), .Z(n14617) );
  NOR2_X1 U17673 ( .A1(n5669), .A2(n16704), .ZN(n4893) );
  OAI21_X1 U17674 ( .A1(n13123), .A2(n13771), .B(n10190), .ZN(n10189) );
  AND2_X1 U17677 ( .A1(n19750), .A2(n10836), .Z(n10518) );
  XOR2_X1 U17681 ( .A1(n4894), .A2(n12330), .Z(n5080) );
  OAI21_X1 U17682 ( .A1(n4713), .A2(n12952), .B(n4895), .ZN(n16006) );
  NAND2_X1 U17690 ( .A1(n17202), .A2(n935), .ZN(n17201) );
  OR2_X1 U17691 ( .A1(n28203), .A2(n28001), .Z(n4897) );
  INV_X2 U17693 ( .I(n4899), .ZN(n20408) );
  XOR2_X1 U17695 ( .A1(n29027), .A2(n681), .Z(n4900) );
  NAND2_X2 U17702 ( .A1(n4901), .A2(n18108), .ZN(n26109) );
  OR2_X1 U17704 ( .A1(n21989), .A2(n12365), .Z(n15652) );
  XOR2_X1 U17706 ( .A1(n11319), .A2(n16460), .Z(n11318) );
  XNOR2_X1 U17707 ( .A1(n3528), .A2(n17727), .ZN(n8785) );
  XOR2_X1 U17711 ( .A1(n17554), .A2(n9748), .Z(n20194) );
  NAND2_X2 U17716 ( .A1(n28467), .A2(n16840), .ZN(n29247) );
  NAND2_X1 U17728 ( .A1(n6488), .A2(n6489), .ZN(n6487) );
  OR2_X1 U17730 ( .A1(n22783), .A2(n38725), .Z(n15375) );
  OR2_X1 U17731 ( .A1(n20407), .A2(n20408), .Z(n13373) );
  XOR2_X1 U17735 ( .A1(n29837), .A2(n28840), .Z(n6536) );
  NAND2_X1 U17742 ( .A1(n18670), .A2(n29341), .ZN(n4919) );
  AND2_X1 U17745 ( .A1(n12964), .A2(n36006), .Z(n5461) );
  NOR2_X2 U17751 ( .A1(n12537), .A2(n32535), .ZN(n11438) );
  XOR2_X1 U17755 ( .A1(n14955), .A2(n21279), .Z(n4929) );
  XOR2_X1 U17772 ( .A1(n13012), .A2(n13013), .Z(n13286) );
  NAND2_X2 U17776 ( .A1(n4936), .A2(n20302), .ZN(n13038) );
  XOR2_X1 U17777 ( .A1(n26181), .A2(n26182), .Z(n17922) );
  XNOR2_X1 U17779 ( .A1(n22670), .A2(n2383), .ZN(n12806) );
  NOR2_X2 U17790 ( .A1(n11443), .A2(n27010), .ZN(n19642) );
  OR2_X1 U17795 ( .A1(n25327), .A2(n5080), .Z(n25535) );
  NAND3_X2 U17798 ( .A1(n10577), .A2(n10578), .A3(n27106), .ZN(n20976) );
  NAND2_X1 U17800 ( .A1(n30845), .A2(n7529), .ZN(n14276) );
  INV_X2 U17802 ( .I(n21846), .ZN(n21672) );
  OAI21_X1 U17807 ( .A1(n14551), .A2(n18755), .B(n21751), .ZN(n10419) );
  XOR2_X1 U17812 ( .A1(n22699), .A2(n13768), .Z(n10382) );
  NAND2_X2 U17813 ( .A1(n8649), .A2(n22106), .ZN(n22699) );
  AOI21_X1 U17816 ( .A1(n29806), .A2(n29811), .B(n39018), .ZN(n5144) );
  XOR2_X1 U17817 ( .A1(n25029), .A2(n24588), .Z(n6109) );
  XOR2_X1 U17823 ( .A1(n5291), .A2(n4958), .Z(n19995) );
  INV_X1 U17824 ( .I(n27538), .ZN(n4958) );
  NOR2_X1 U17825 ( .A1(n11300), .A2(n22856), .ZN(n11299) );
  NOR2_X2 U17826 ( .A1(n24717), .A2(n6944), .ZN(n24591) );
  NOR2_X2 U17827 ( .A1(n6917), .A2(n4959), .ZN(n18425) );
  NAND2_X2 U17831 ( .A1(n13075), .A2(n7884), .ZN(n23832) );
  NAND2_X1 U17834 ( .A1(n11202), .A2(n22008), .ZN(n5618) );
  XOR2_X1 U17841 ( .A1(n21087), .A2(n5742), .Z(n4967) );
  NAND2_X1 U17842 ( .A1(n35506), .A2(n1308), .ZN(n4968) );
  INV_X1 U17843 ( .I(n10419), .ZN(n10418) );
  INV_X1 U17846 ( .I(n27690), .ZN(n15547) );
  INV_X1 U17849 ( .I(n13420), .ZN(n13419) );
  XOR2_X1 U17853 ( .A1(n35303), .A2(n27672), .Z(n6026) );
  NAND2_X2 U17856 ( .A1(n11822), .A2(n4972), .ZN(n12028) );
  XNOR2_X1 U17860 ( .A1(n17567), .A2(n29818), .ZN(n5636) );
  XOR2_X1 U17862 ( .A1(n27692), .A2(n756), .Z(n6927) );
  NOR2_X1 U17871 ( .A1(n6322), .A2(n6321), .ZN(n6320) );
  NAND2_X1 U17881 ( .A1(n9725), .A2(n7537), .ZN(n11300) );
  XOR2_X1 U17883 ( .A1(n26375), .A2(n16046), .Z(n26377) );
  XOR2_X1 U17885 ( .A1(n25180), .A2(n4987), .Z(n15517) );
  XOR2_X1 U17886 ( .A1(n24926), .A2(n19904), .Z(n4987) );
  AND2_X1 U17887 ( .A1(n16250), .A2(n35003), .Z(n13885) );
  XOR2_X1 U17890 ( .A1(n5443), .A2(n23919), .Z(n5442) );
  AOI22_X1 U17892 ( .A1(n13143), .A2(n11981), .B1(n13141), .B2(n19303), .ZN(
        n13140) );
  XOR2_X1 U17897 ( .A1(n29096), .A2(n29253), .Z(n28767) );
  XOR2_X1 U17901 ( .A1(n13729), .A2(n16245), .Z(n20384) );
  NAND2_X1 U17905 ( .A1(n19994), .A2(n17644), .ZN(n17684) );
  XOR2_X1 U17909 ( .A1(n29074), .A2(n5648), .Z(n4999) );
  XOR2_X1 U17916 ( .A1(n34009), .A2(n15717), .Z(n5003) );
  NOR2_X2 U17923 ( .A1(n6999), .A2(n6997), .ZN(n24829) );
  AOI21_X2 U17928 ( .A1(n23605), .A2(n23604), .B(n23603), .ZN(n23654) );
  NAND2_X1 U17929 ( .A1(n24232), .A2(n5985), .ZN(n6998) );
  INV_X2 U17938 ( .I(n5012), .ZN(n11795) );
  NOR2_X1 U17944 ( .A1(n30059), .A2(n36166), .ZN(n21168) );
  OR2_X1 U17946 ( .A1(n6623), .A2(n29980), .Z(n5019) );
  XOR2_X1 U17956 ( .A1(n29304), .A2(n29305), .Z(n14872) );
  XOR2_X1 U17957 ( .A1(n29113), .A2(n29254), .Z(n29305) );
  NAND2_X2 U17963 ( .A1(n6110), .A2(n27122), .ZN(n27786) );
  XOR2_X1 U17966 ( .A1(n5033), .A2(n24915), .Z(n19572) );
  NAND2_X1 U17968 ( .A1(n32450), .A2(n7467), .ZN(n7466) );
  OAI22_X1 U17969 ( .A1(n9954), .A2(n14390), .B1(n34073), .B2(n23071), .ZN(
        n16693) );
  XOR2_X1 U17973 ( .A1(n18094), .A2(n5037), .Z(n5525) );
  XOR2_X1 U17974 ( .A1(n27628), .A2(n27627), .Z(n5037) );
  INV_X1 U17977 ( .I(n23686), .ZN(n6227) );
  AND2_X1 U17980 ( .A1(n25851), .A2(n11858), .Z(n6399) );
  XOR2_X1 U17984 ( .A1(n21235), .A2(n5048), .Z(n21234) );
  XOR2_X1 U17985 ( .A1(n18526), .A2(n31515), .Z(n5048) );
  XOR2_X1 U17996 ( .A1(n17195), .A2(n1050), .Z(n12598) );
  OR2_X1 U18003 ( .A1(n8245), .A2(n12631), .Z(n7626) );
  NAND2_X2 U18005 ( .A1(n5054), .A2(n18589), .ZN(n20307) );
  XOR2_X1 U18009 ( .A1(n28946), .A2(n28945), .Z(n5587) );
  XOR2_X1 U18013 ( .A1(n3953), .A2(n17189), .Z(n5055) );
  NAND2_X1 U18015 ( .A1(n9616), .A2(n22155), .ZN(n15435) );
  XOR2_X1 U18019 ( .A1(n8401), .A2(n15197), .Z(n5651) );
  NAND2_X2 U18020 ( .A1(n5623), .A2(n5622), .ZN(n8401) );
  XOR2_X1 U18021 ( .A1(n25253), .A2(n19022), .Z(n5058) );
  AOI21_X2 U18028 ( .A1(n11869), .A2(n19055), .B(n11868), .ZN(n11867) );
  XOR2_X1 U18031 ( .A1(n5065), .A2(n14820), .Z(Ciphertext[115]) );
  XOR2_X1 U18033 ( .A1(n15758), .A2(n25178), .Z(n17108) );
  XOR2_X1 U18034 ( .A1(n23965), .A2(n5071), .Z(n23966) );
  XOR2_X1 U18035 ( .A1(n5073), .A2(n19950), .Z(Ciphertext[106]) );
  NOR2_X1 U18041 ( .A1(n29719), .A2(n5921), .ZN(n16629) );
  NAND2_X2 U18049 ( .A1(n8961), .A2(n12974), .ZN(n13779) );
  OR2_X1 U18051 ( .A1(n17496), .A2(n16841), .Z(n17495) );
  NAND2_X1 U18061 ( .A1(n5773), .A2(n5772), .ZN(n5771) );
  XOR2_X1 U18065 ( .A1(n5088), .A2(n19845), .Z(Ciphertext[19]) );
  XOR2_X1 U18070 ( .A1(n29086), .A2(n13497), .Z(n5090) );
  NAND2_X1 U18071 ( .A1(n8231), .A2(n39083), .ZN(n8229) );
  XOR2_X1 U18072 ( .A1(n7031), .A2(n5091), .Z(n28961) );
  XOR2_X1 U18073 ( .A1(n29026), .A2(n28849), .Z(n5091) );
  XOR2_X1 U18077 ( .A1(n5094), .A2(n23910), .Z(n5293) );
  XOR2_X1 U18086 ( .A1(n16218), .A2(n677), .Z(n5096) );
  OR2_X1 U18091 ( .A1(n31564), .A2(n17790), .Z(n23958) );
  NAND3_X2 U18097 ( .A1(n6521), .A2(n6520), .A3(n9988), .ZN(n6527) );
  XOR2_X1 U18107 ( .A1(n25164), .A2(n10431), .Z(n5114) );
  XOR2_X1 U18112 ( .A1(n5119), .A2(n5120), .Z(n5118) );
  XOR2_X1 U18113 ( .A1(n26531), .A2(n26305), .Z(n5120) );
  NAND2_X1 U18118 ( .A1(n5126), .A2(n26128), .ZN(n25892) );
  NAND2_X1 U18119 ( .A1(n26126), .A2(n5126), .ZN(n5687) );
  XOR2_X1 U18128 ( .A1(n16781), .A2(n5142), .Z(n14258) );
  XOR2_X1 U18129 ( .A1(n14219), .A2(n23658), .Z(n5142) );
  XOR2_X1 U18130 ( .A1(n5143), .A2(n20781), .Z(Ciphertext[108]) );
  XOR2_X1 U18132 ( .A1(n5153), .A2(n28889), .Z(n29036) );
  NOR2_X2 U18133 ( .A1(n5151), .A2(n5150), .ZN(n28889) );
  OAI21_X1 U18140 ( .A1(n27385), .A2(n27064), .B(n34562), .ZN(n5167) );
  XOR2_X1 U18141 ( .A1(n5171), .A2(n13564), .Z(n6310) );
  XOR2_X1 U18142 ( .A1(n5171), .A2(n22598), .Z(n13844) );
  XOR2_X1 U18143 ( .A1(n5171), .A2(n4624), .Z(n22686) );
  XOR2_X1 U18152 ( .A1(n5185), .A2(n14820), .Z(n14819) );
  NAND2_X1 U18154 ( .A1(n5192), .A2(n5188), .ZN(Ciphertext[139]) );
  NAND2_X1 U18155 ( .A1(n5189), .A2(n5369), .ZN(n5188) );
  NOR2_X1 U18156 ( .A1(n5191), .A2(n5190), .ZN(n5189) );
  NAND2_X1 U18157 ( .A1(n5270), .A2(n30010), .ZN(n5190) );
  NOR2_X1 U18158 ( .A1(n30032), .A2(n39407), .ZN(n5191) );
  NOR3_X1 U18159 ( .A1(n5195), .A2(n5194), .A3(n5193), .ZN(n5192) );
  NOR2_X1 U18160 ( .A1(n5270), .A2(n30010), .ZN(n5193) );
  NOR3_X1 U18161 ( .A1(n30032), .A2(n39407), .A3(n30010), .ZN(n5195) );
  INV_X2 U18164 ( .I(n11727), .ZN(n25727) );
  OAI22_X2 U18166 ( .A1(n25491), .A2(n14947), .B1(n25142), .B2(n30470), .ZN(
        n9833) );
  INV_X2 U18171 ( .I(n18707), .ZN(n22709) );
  XOR2_X1 U18173 ( .A1(n28500), .A2(n1160), .Z(n28793) );
  XOR2_X1 U18176 ( .A1(n13853), .A2(n26162), .Z(n5226) );
  XOR2_X1 U18177 ( .A1(n25063), .A2(n5271), .Z(n5228) );
  XNOR2_X1 U18178 ( .A1(n25266), .A2(n25290), .ZN(n5271) );
  XOR2_X1 U18180 ( .A1(n25159), .A2(n813), .Z(n5229) );
  XOR2_X1 U18186 ( .A1(n20353), .A2(n29432), .Z(n5235) );
  XOR2_X1 U18188 ( .A1(n7148), .A2(n30065), .Z(n5238) );
  XOR2_X1 U18190 ( .A1(n5241), .A2(n26325), .Z(n8189) );
  XOR2_X1 U18193 ( .A1(n5242), .A2(n4413), .Z(n11967) );
  XOR2_X1 U18194 ( .A1(n5242), .A2(n29282), .Z(n22057) );
  XOR2_X1 U18199 ( .A1(n19094), .A2(n21048), .Z(n5247) );
  AND2_X1 U18201 ( .A1(n25618), .A2(n19264), .Z(n5249) );
  INV_X1 U18203 ( .I(n31767), .ZN(n5251) );
  NAND2_X2 U18215 ( .A1(n9231), .A2(n15643), .ZN(n5270) );
  XOR2_X1 U18226 ( .A1(n19781), .A2(n5285), .Z(n19692) );
  XOR2_X1 U18227 ( .A1(n5286), .A2(n22487), .Z(n5285) );
  XOR2_X1 U18228 ( .A1(n22644), .A2(n5284), .Z(n5286) );
  XOR2_X1 U18232 ( .A1(n6559), .A2(n5290), .Z(n18622) );
  XOR2_X1 U18235 ( .A1(n32464), .A2(n18004), .Z(n8780) );
  NAND3_X1 U18238 ( .A1(n36989), .A2(n6445), .A3(n8137), .ZN(n5295) );
  INV_X2 U18242 ( .I(n19224), .ZN(n30153) );
  XOR2_X1 U18254 ( .A1(n10424), .A2(n9309), .Z(n5316) );
  XOR2_X1 U18257 ( .A1(n5320), .A2(n17859), .Z(n5318) );
  XNOR2_X1 U18265 ( .A1(n5338), .A2(n5339), .ZN(n5337) );
  XOR2_X1 U18269 ( .A1(n5340), .A2(n14530), .Z(n5339) );
  INV_X1 U18283 ( .I(n12916), .ZN(n5367) );
  XOR2_X1 U18285 ( .A1(n14333), .A2(Key[71]), .Z(n21518) );
  MUX2_X1 U18286 ( .I0(n21039), .I1(n36404), .S(n25975), .Z(n16201) );
  NOR2_X1 U18288 ( .A1(n14838), .A2(n3487), .ZN(n10089) );
  XOR2_X1 U18289 ( .A1(n16524), .A2(n23814), .Z(n23676) );
  XOR2_X1 U18291 ( .A1(n5323), .A2(n29514), .Z(n5370) );
  XOR2_X1 U18294 ( .A1(n27566), .A2(n27767), .Z(n27721) );
  OR2_X1 U18296 ( .A1(n27220), .A2(n37077), .Z(n5377) );
  NOR2_X1 U18297 ( .A1(n3273), .A2(n5380), .ZN(n15885) );
  NAND2_X1 U18298 ( .A1(n5929), .A2(n8882), .ZN(n10434) );
  NAND2_X2 U18301 ( .A1(n23994), .A2(n23993), .ZN(n24814) );
  XOR2_X1 U18306 ( .A1(n5625), .A2(n11755), .Z(n5394) );
  XOR2_X1 U18308 ( .A1(n27716), .A2(n7801), .Z(n5395) );
  XOR2_X1 U18316 ( .A1(n8163), .A2(n1361), .Z(n5407) );
  INV_X2 U18321 ( .I(n11543), .ZN(n30154) );
  NAND3_X1 U18325 ( .A1(n30177), .A2(n35899), .A3(n30184), .ZN(n5422) );
  INV_X1 U18326 ( .I(Plaintext[9]), .ZN(n5423) );
  XOR2_X1 U18327 ( .A1(n5423), .A2(Key[9]), .Z(n13397) );
  AOI21_X1 U18331 ( .A1(n30069), .A2(n30071), .B(n30078), .ZN(n20948) );
  XOR2_X1 U18332 ( .A1(n35215), .A2(n17850), .Z(n23920) );
  XOR2_X1 U18333 ( .A1(n39038), .A2(n19833), .Z(n5443) );
  XOR2_X1 U18334 ( .A1(n20540), .A2(n1096), .Z(n26373) );
  XOR2_X1 U18336 ( .A1(n5447), .A2(n5445), .Z(n5444) );
  XOR2_X1 U18337 ( .A1(n5446), .A2(n26244), .Z(n5445) );
  XOR2_X1 U18338 ( .A1(n26252), .A2(n19866), .Z(n5446) );
  OAI21_X1 U18341 ( .A1(n29338), .A2(n16889), .B(n31532), .ZN(n12848) );
  NOR2_X1 U18350 ( .A1(n28812), .A2(n5465), .ZN(n18471) );
  NAND2_X1 U18351 ( .A1(n28811), .A2(n5465), .ZN(n18473) );
  XOR2_X1 U18354 ( .A1(n39600), .A2(n25074), .Z(n5472) );
  XOR2_X1 U18356 ( .A1(n6352), .A2(n12438), .Z(n5473) );
  XOR2_X1 U18365 ( .A1(n27745), .A2(n29661), .Z(n5486) );
  OAI21_X2 U18366 ( .A1(n21140), .A2(n38305), .B(n21139), .ZN(n27745) );
  INV_X4 U18367 ( .I(n23634), .ZN(n23468) );
  OAI21_X2 U18368 ( .A1(n23635), .A2(n5491), .B(n5488), .ZN(n24050) );
  NAND2_X1 U18371 ( .A1(n5798), .A2(n1530), .ZN(n15882) );
  XOR2_X1 U18375 ( .A1(n5510), .A2(n5511), .Z(n24104) );
  XOR2_X1 U18379 ( .A1(n13977), .A2(n23674), .Z(n5511) );
  INV_X1 U18386 ( .I(n5709), .ZN(n18810) );
  XOR2_X1 U18392 ( .A1(n35270), .A2(n5524), .Z(n5522) );
  NAND2_X1 U18394 ( .A1(n28286), .A2(n11375), .ZN(n6375) );
  XOR2_X1 U18395 ( .A1(n9030), .A2(n26396), .Z(n25853) );
  XOR2_X1 U18396 ( .A1(n9030), .A2(n19885), .Z(n14102) );
  INV_X1 U18397 ( .I(n5527), .ZN(n20147) );
  NOR2_X1 U18401 ( .A1(n5530), .A2(n29284), .ZN(n29276) );
  NOR2_X1 U18402 ( .A1(n37157), .A2(n5530), .ZN(n9445) );
  OAI21_X1 U18403 ( .A1(n18611), .A2(n18610), .B(n36676), .ZN(n29280) );
  XOR2_X1 U18406 ( .A1(n7464), .A2(n8475), .Z(n12400) );
  XOR2_X1 U18409 ( .A1(n5540), .A2(n5538), .Z(n13572) );
  XOR2_X1 U18410 ( .A1(n17413), .A2(n5539), .Z(n5538) );
  XOR2_X1 U18411 ( .A1(n13564), .A2(n29514), .Z(n5539) );
  NAND2_X1 U18424 ( .A1(n36763), .A2(n936), .ZN(n23141) );
  AOI21_X2 U18432 ( .A1(n20504), .A2(n20503), .B(n15564), .ZN(n23710) );
  XOR2_X1 U18433 ( .A1(n5561), .A2(n5562), .Z(n5986) );
  XOR2_X1 U18434 ( .A1(n23756), .A2(n7017), .Z(n5561) );
  XOR2_X1 U18435 ( .A1(n5563), .A2(n23653), .Z(n5562) );
  XOR2_X1 U18436 ( .A1(n8045), .A2(n5564), .Z(n5563) );
  XOR2_X1 U18438 ( .A1(n27713), .A2(n761), .Z(n5565) );
  XOR2_X1 U18446 ( .A1(n22567), .A2(n2383), .Z(n17528) );
  XOR2_X1 U18450 ( .A1(n12464), .A2(n5583), .Z(n8943) );
  XOR2_X1 U18452 ( .A1(n5639), .A2(n18609), .Z(n5584) );
  XOR2_X1 U18453 ( .A1(n10079), .A2(n29050), .Z(n5586) );
  NOR2_X1 U18459 ( .A1(n20924), .A2(n16114), .ZN(n5596) );
  NAND2_X1 U18461 ( .A1(n19587), .A2(n686), .ZN(n5598) );
  XOR2_X1 U18462 ( .A1(n743), .A2(n17680), .Z(n5600) );
  AOI21_X2 U18488 ( .A1(n15651), .A2(n30239), .B(n5632), .ZN(n30262) );
  XOR2_X1 U18492 ( .A1(n5637), .A2(n5636), .Z(n5635) );
  NAND2_X1 U18495 ( .A1(n10836), .A2(n11890), .ZN(n27915) );
  NAND2_X2 U18499 ( .A1(n5930), .A2(n5931), .ZN(n5929) );
  XOR2_X1 U18505 ( .A1(n31550), .A2(n6854), .Z(n6853) );
  XOR2_X1 U18506 ( .A1(n29024), .A2(n5647), .Z(n5646) );
  XOR2_X1 U18507 ( .A1(n29122), .A2(n19897), .Z(n5647) );
  XOR2_X1 U18513 ( .A1(n27781), .A2(n27637), .Z(n5650) );
  XOR2_X1 U18516 ( .A1(n5652), .A2(n29071), .Z(n10258) );
  XOR2_X1 U18517 ( .A1(n5652), .A2(n1165), .Z(n17832) );
  XOR2_X1 U18518 ( .A1(n27823), .A2(n35229), .Z(n5655) );
  INV_X2 U18519 ( .I(n5656), .ZN(n19469) );
  XOR2_X1 U18526 ( .A1(n9719), .A2(n1167), .Z(n11189) );
  INV_X1 U18528 ( .I(n11166), .ZN(n5670) );
  NAND2_X1 U18529 ( .A1(n28159), .A2(n6548), .ZN(n11166) );
  NAND2_X1 U18532 ( .A1(n1104), .A2(n26055), .ZN(n5674) );
  AOI21_X1 U18536 ( .A1(n29977), .A2(n5678), .B(n13705), .ZN(n5677) );
  OAI21_X1 U18537 ( .A1(n26126), .A2(n15677), .B(n5687), .ZN(n5686) );
  XOR2_X1 U18541 ( .A1(n5692), .A2(n5691), .Z(n5690) );
  XOR2_X1 U18544 ( .A1(n12865), .A2(n18487), .Z(n5694) );
  XOR2_X1 U18546 ( .A1(n1460), .A2(n27676), .Z(n5697) );
  XOR2_X1 U18547 ( .A1(n10370), .A2(n18981), .Z(n18980) );
  XOR2_X1 U18549 ( .A1(n23924), .A2(n5699), .Z(n17874) );
  MUX2_X1 U18554 ( .I0(n27866), .I1(n27928), .S(n28193), .Z(n5707) );
  INV_X2 U18558 ( .I(n5717), .ZN(n18342) );
  XOR2_X1 U18561 ( .A1(n6951), .A2(n6952), .Z(n5719) );
  XOR2_X1 U18564 ( .A1(n9567), .A2(n16093), .Z(n5722) );
  XOR2_X1 U18568 ( .A1(n5726), .A2(n5725), .Z(n5724) );
  XOR2_X1 U18569 ( .A1(n29819), .A2(n29818), .Z(n5725) );
  AOI21_X2 U18570 ( .A1(n20951), .A2(n28750), .B(n13656), .ZN(n29818) );
  XOR2_X1 U18571 ( .A1(n38160), .A2(n15617), .Z(n5726) );
  XOR2_X1 U18575 ( .A1(n25247), .A2(n30126), .Z(n5730) );
  XOR2_X1 U18577 ( .A1(n25245), .A2(n11905), .Z(n5731) );
  INV_X1 U18579 ( .I(n31528), .ZN(n24071) );
  XOR2_X1 U18580 ( .A1(n15916), .A2(n31528), .Z(n7017) );
  XOR2_X1 U18582 ( .A1(n31528), .A2(n19646), .Z(n20045) );
  XOR2_X1 U18584 ( .A1(n5737), .A2(n12412), .Z(n14121) );
  XOR2_X1 U18590 ( .A1(n29045), .A2(n1163), .Z(n14195) );
  XOR2_X1 U18591 ( .A1(n5741), .A2(n28707), .Z(n7665) );
  XOR2_X1 U18592 ( .A1(n35266), .A2(n29298), .Z(n5742) );
  XOR2_X1 U18596 ( .A1(n15368), .A2(n1214), .Z(n5744) );
  AOI21_X2 U18597 ( .A1(n5748), .A2(n5837), .B(n5747), .ZN(n23610) );
  XOR2_X1 U18599 ( .A1(n5750), .A2(n29506), .Z(n18487) );
  XOR2_X1 U18604 ( .A1(n37044), .A2(n661), .Z(n5760) );
  XOR2_X1 U18605 ( .A1(n24031), .A2(n11267), .Z(n5761) );
  OAI22_X1 U18607 ( .A1(n29869), .A2(n5762), .B1(n20793), .B2(n4879), .ZN(
        n5971) );
  XOR2_X1 U18609 ( .A1(n5766), .A2(n5763), .Z(n18210) );
  XOR2_X1 U18610 ( .A1(n5765), .A2(n5764), .Z(n5763) );
  XOR2_X1 U18611 ( .A1(n26402), .A2(n37109), .Z(n5764) );
  XOR2_X1 U18614 ( .A1(n12429), .A2(n26242), .Z(n5766) );
  OAI21_X1 U18616 ( .A1(n1581), .A2(n5768), .B(n36395), .ZN(n19836) );
  OR2_X1 U18618 ( .A1(n27270), .A2(n5772), .Z(n5775) );
  XOR2_X1 U18620 ( .A1(n5778), .A2(n29718), .Z(Ciphertext[93]) );
  XOR2_X1 U18621 ( .A1(n28958), .A2(n28959), .Z(n5781) );
  XOR2_X1 U18627 ( .A1(n25257), .A2(n24960), .Z(n5789) );
  AOI21_X2 U18628 ( .A1(n11769), .A2(n11768), .B(n17663), .ZN(n6066) );
  XOR2_X1 U18629 ( .A1(n18427), .A2(n5793), .Z(n24202) );
  INV_X1 U18630 ( .I(n23945), .ZN(n5794) );
  XOR2_X1 U18631 ( .A1(n23929), .A2(n24040), .Z(n23945) );
  XOR2_X1 U18636 ( .A1(n17623), .A2(n24962), .Z(n5801) );
  XOR2_X1 U18638 ( .A1(n15288), .A2(n25865), .Z(n5803) );
  XOR2_X1 U18640 ( .A1(n26492), .A2(n26210), .Z(n5804) );
  NAND2_X2 U18643 ( .A1(n5807), .A2(n5805), .ZN(n18866) );
  XOR2_X1 U18644 ( .A1(n5814), .A2(n6112), .Z(n5815) );
  XOR2_X1 U18645 ( .A1(n15186), .A2(n25079), .Z(n5814) );
  AND2_X1 U18653 ( .A1(n22282), .A2(n5819), .Z(n6485) );
  XOR2_X1 U18656 ( .A1(n23873), .A2(n29711), .Z(n5820) );
  OAI21_X2 U18657 ( .A1(n5823), .A2(n526), .B(n5822), .ZN(n8071) );
  XOR2_X1 U18663 ( .A1(n5830), .A2(n1554), .Z(n5829) );
  XOR2_X1 U18664 ( .A1(n6759), .A2(n29661), .Z(n5830) );
  NAND2_X2 U18672 ( .A1(n8358), .A2(n8361), .ZN(n24764) );
  XOR2_X1 U18674 ( .A1(n5841), .A2(n15203), .Z(n5842) );
  XOR2_X1 U18675 ( .A1(n23714), .A2(n23883), .Z(n24068) );
  XOR2_X1 U18678 ( .A1(n15531), .A2(n5844), .Z(n5843) );
  XOR2_X1 U18679 ( .A1(n25216), .A2(n19516), .Z(n5844) );
  AOI22_X2 U18680 ( .A1(n21028), .A2(n24749), .B1(n20944), .B2(n18858), .ZN(
        n25216) );
  NAND2_X2 U18682 ( .A1(n24965), .A2(n16819), .ZN(n24942) );
  XOR2_X1 U18691 ( .A1(n9719), .A2(n7056), .Z(n22516) );
  XOR2_X1 U18692 ( .A1(n37660), .A2(n1361), .Z(n5861) );
  XOR2_X1 U18693 ( .A1(n5862), .A2(n29034), .Z(n28888) );
  XOR2_X1 U18694 ( .A1(n28982), .A2(n5862), .Z(n12561) );
  AOI21_X2 U18697 ( .A1(n14339), .A2(n11680), .B(n7647), .ZN(n5862) );
  XOR2_X1 U18701 ( .A1(n23686), .A2(n29562), .Z(n5866) );
  XOR2_X1 U18704 ( .A1(n10253), .A2(n10252), .Z(n5867) );
  NAND2_X1 U18708 ( .A1(n5871), .A2(n31679), .ZN(n24539) );
  XOR2_X1 U18710 ( .A1(n27736), .A2(n19874), .Z(n5873) );
  NOR3_X1 U18716 ( .A1(n4674), .A2(n17091), .A3(n36792), .ZN(n25450) );
  NAND3_X1 U18725 ( .A1(n24709), .A2(n5897), .A3(n34526), .ZN(n7595) );
  OAI21_X1 U18726 ( .A1(n24708), .A2(n24529), .B(n5897), .ZN(n6083) );
  INV_X2 U18736 ( .I(n18186), .ZN(n27866) );
  XOR2_X1 U18741 ( .A1(n360), .A2(n5914), .Z(n5913) );
  XOR2_X1 U18744 ( .A1(n10424), .A2(n723), .Z(n5917) );
  XOR2_X1 U18745 ( .A1(n6896), .A2(n25271), .Z(n10424) );
  XOR2_X1 U18747 ( .A1(n23868), .A2(n5919), .Z(n5918) );
  XOR2_X1 U18748 ( .A1(n23774), .A2(n23686), .Z(n5919) );
  NAND2_X2 U18749 ( .A1(n10208), .A2(n10207), .ZN(n19656) );
  XOR2_X1 U18750 ( .A1(n23740), .A2(n23687), .Z(n5920) );
  NAND2_X1 U18756 ( .A1(n21377), .A2(n21565), .ZN(n5931) );
  XOR2_X1 U18760 ( .A1(n23848), .A2(n16258), .Z(n5936) );
  XOR2_X1 U18761 ( .A1(n24031), .A2(n16257), .Z(n5937) );
  AND2_X1 U18762 ( .A1(n34279), .A2(n31433), .Z(n5941) );
  AOI21_X1 U18764 ( .A1(n17731), .A2(n29719), .B(n5921), .ZN(n5949) );
  OAI21_X1 U18768 ( .A1(n7835), .A2(n1288), .B(n5953), .ZN(n24485) );
  XOR2_X1 U18770 ( .A1(n5956), .A2(n13681), .Z(n8812) );
  XOR2_X1 U18771 ( .A1(n17569), .A2(n22321), .Z(n5956) );
  XOR2_X1 U18778 ( .A1(n10635), .A2(n34848), .Z(n5959) );
  NAND2_X2 U18786 ( .A1(n5969), .A2(n5968), .ZN(n20460) );
  INV_X2 U18788 ( .I(n5975), .ZN(n19823) );
  XOR2_X1 U18792 ( .A1(n12863), .A2(n12861), .Z(n5974) );
  NAND3_X2 U18801 ( .A1(n17393), .A2(n17391), .A3(n14457), .ZN(n7611) );
  INV_X2 U18802 ( .I(n5986), .ZN(n19915) );
  XOR2_X1 U18807 ( .A1(n5993), .A2(n5992), .Z(n5991) );
  OAI22_X1 U18810 ( .A1(n33864), .A2(n30299), .B1(n23381), .B2(n31594), .ZN(
        n5999) );
  NOR2_X1 U18812 ( .A1(n29220), .A2(n35264), .ZN(n13123) );
  AOI21_X1 U18814 ( .A1(n31772), .A2(n18240), .B(n6002), .ZN(n13108) );
  NOR2_X1 U18815 ( .A1(n10685), .A2(n6002), .ZN(n10050) );
  NAND2_X1 U18817 ( .A1(n13761), .A2(n6002), .ZN(n6001) );
  XOR2_X1 U18819 ( .A1(n26358), .A2(n6008), .Z(n6007) );
  XOR2_X1 U18820 ( .A1(n26596), .A2(n19751), .Z(n6008) );
  NOR3_X1 U18821 ( .A1(n5314), .A2(n10882), .A3(n953), .ZN(n11944) );
  XOR2_X1 U18827 ( .A1(n5284), .A2(n22743), .Z(n7277) );
  OAI21_X2 U18828 ( .A1(n22305), .A2(n6015), .B(n22304), .ZN(n22743) );
  INV_X2 U18830 ( .I(n8694), .ZN(n12925) );
  OR2_X2 U18831 ( .A1(n20649), .A2(n6449), .Z(n16468) );
  NAND2_X1 U18832 ( .A1(n30053), .A2(n6019), .ZN(n29180) );
  XOR2_X1 U18834 ( .A1(n12053), .A2(n6029), .Z(n7462) );
  XOR2_X1 U18835 ( .A1(n7854), .A2(n6030), .Z(n6029) );
  XOR2_X1 U18836 ( .A1(n35240), .A2(n33811), .Z(n6030) );
  XOR2_X1 U18842 ( .A1(n6035), .A2(n22563), .Z(n6034) );
  XOR2_X1 U18843 ( .A1(n22485), .A2(n33661), .Z(n6035) );
  NOR2_X1 U18845 ( .A1(n19089), .A2(n6036), .ZN(n13910) );
  OAI21_X1 U18847 ( .A1(n22156), .A2(n6036), .B(n16935), .ZN(n13912) );
  INV_X4 U18850 ( .I(n19604), .ZN(n6036) );
  OAI21_X2 U18851 ( .A1(n15955), .A2(n24094), .B(n9909), .ZN(n24878) );
  INV_X1 U18856 ( .I(n4441), .ZN(n9074) );
  XOR2_X1 U18857 ( .A1(n4441), .A2(n4123), .Z(n6047) );
  NAND2_X1 U18868 ( .A1(n23583), .A2(n1626), .ZN(n6053) );
  XOR2_X1 U18871 ( .A1(n6412), .A2(n26206), .Z(n6057) );
  XOR2_X1 U18874 ( .A1(n6066), .A2(n25184), .Z(n25042) );
  INV_X2 U18886 ( .I(n7140), .ZN(n20931) );
  XOR2_X1 U18887 ( .A1(n6092), .A2(n6090), .Z(n17660) );
  XOR2_X1 U18890 ( .A1(n19608), .A2(n29554), .Z(n6091) );
  OAI21_X2 U18892 ( .A1(n28531), .A2(n6095), .B(n6094), .ZN(n29082) );
  XOR2_X1 U18896 ( .A1(n12251), .A2(n6108), .Z(n6107) );
  XOR2_X1 U18897 ( .A1(n13917), .A2(n39765), .Z(n6108) );
  XNOR2_X1 U18899 ( .A1(n27786), .A2(n27632), .ZN(n16066) );
  XOR2_X1 U18904 ( .A1(n33921), .A2(n19749), .Z(n6112) );
  NAND2_X1 U18905 ( .A1(n6121), .A2(n6120), .ZN(n6126) );
  NAND2_X1 U18909 ( .A1(n6126), .A2(n6125), .ZN(n6124) );
  NAND3_X1 U18911 ( .A1(n5061), .A2(n6128), .A3(n22248), .ZN(n21739) );
  XOR2_X1 U18914 ( .A1(n9085), .A2(n6131), .Z(n6133) );
  NOR2_X1 U18921 ( .A1(n35990), .A2(n27267), .ZN(n27055) );
  AOI21_X1 U18923 ( .A1(n27129), .A2(n27128), .B(n36177), .ZN(n9727) );
  NOR2_X1 U18924 ( .A1(n19662), .A2(n35990), .ZN(n27130) );
  XOR2_X1 U18925 ( .A1(n6148), .A2(n19903), .Z(Ciphertext[155]) );
  XOR2_X1 U18929 ( .A1(n13961), .A2(n17117), .Z(n17060) );
  NAND2_X2 U18933 ( .A1(n18748), .A2(n19177), .ZN(n6159) );
  XOR2_X1 U18934 ( .A1(Key[131]), .A2(Plaintext[131]), .Z(n6161) );
  INV_X2 U18935 ( .I(n6161), .ZN(n21308) );
  NAND2_X1 U18938 ( .A1(n19941), .A2(n25449), .ZN(n6172) );
  XOR2_X1 U18940 ( .A1(n11165), .A2(n11266), .Z(n13144) );
  XOR2_X1 U18941 ( .A1(n6177), .A2(n29298), .Z(n20232) );
  NOR2_X1 U18948 ( .A1(n11126), .A2(n39268), .ZN(n6189) );
  NOR2_X1 U18950 ( .A1(n19951), .A2(n6190), .ZN(n10442) );
  NAND2_X1 U18957 ( .A1(n6198), .A2(n21667), .ZN(n6197) );
  AOI21_X1 U18959 ( .A1(n13574), .A2(n1407), .B(n14158), .ZN(n6207) );
  XOR2_X1 U18962 ( .A1(n6677), .A2(n6212), .Z(n6211) );
  NAND2_X1 U18964 ( .A1(n23528), .A2(n6218), .ZN(n23221) );
  INV_X1 U18965 ( .I(n6218), .ZN(n6216) );
  NAND2_X1 U18966 ( .A1(n18086), .A2(n6218), .ZN(n20978) );
  NOR2_X2 U18967 ( .A1(n15588), .A2(n15589), .ZN(n6218) );
  XOR2_X1 U18968 ( .A1(n6224), .A2(n6225), .Z(n6223) );
  XOR2_X1 U18970 ( .A1(n12243), .A2(n19860), .Z(n6225) );
  XOR2_X1 U18974 ( .A1(n6233), .A2(n6231), .Z(n25322) );
  XOR2_X1 U18976 ( .A1(n31579), .A2(n1167), .Z(n6232) );
  NAND2_X1 U18983 ( .A1(n6241), .A2(n261), .ZN(n14124) );
  NAND2_X2 U18984 ( .A1(n17534), .A2(n6241), .ZN(n9102) );
  NOR2_X1 U18988 ( .A1(n39140), .A2(n38198), .ZN(n6783) );
  XOR2_X1 U18990 ( .A1(n6527), .A2(n23776), .Z(n23804) );
  XOR2_X1 U18992 ( .A1(n39231), .A2(n6429), .Z(n6428) );
  XOR2_X1 U18993 ( .A1(n38207), .A2(n1938), .Z(n8896) );
  INV_X2 U18999 ( .I(n11084), .ZN(n16828) );
  XOR2_X1 U19006 ( .A1(n22656), .A2(n17428), .Z(n12125) );
  XOR2_X1 U19007 ( .A1(n22656), .A2(n13564), .Z(n11289) );
  INV_X2 U19017 ( .I(n21214), .ZN(n22146) );
  XOR2_X1 U19023 ( .A1(n19960), .A2(n6281), .Z(n19959) );
  XOR2_X1 U19024 ( .A1(n23709), .A2(n8929), .Z(n6281) );
  XOR2_X1 U19025 ( .A1(n8447), .A2(n24927), .Z(n6283) );
  OAI22_X2 U19027 ( .A1(n6286), .A2(n39812), .B1(n23553), .B2(n18747), .ZN(
        n14219) );
  OAI21_X1 U19028 ( .A1(n6287), .A2(n1420), .B(n38155), .ZN(n15964) );
  XOR2_X1 U19031 ( .A1(n7944), .A2(n29649), .Z(n6289) );
  XOR2_X1 U19032 ( .A1(n26400), .A2(n1509), .Z(n26555) );
  XOR2_X1 U19033 ( .A1(n35239), .A2(n26359), .Z(n26400) );
  XOR2_X1 U19035 ( .A1(n6294), .A2(n20136), .Z(n20135) );
  INV_X1 U19036 ( .I(n17493), .ZN(n6294) );
  NAND2_X1 U19042 ( .A1(n26060), .A2(n6302), .ZN(n7677) );
  MUX2_X1 U19044 ( .I0(n18176), .I1(n26063), .S(n25943), .Z(n26065) );
  XOR2_X1 U19047 ( .A1(n6305), .A2(n6306), .Z(n6304) );
  XOR2_X1 U19048 ( .A1(n5021), .A2(n1727), .Z(n6305) );
  XOR2_X1 U19050 ( .A1(n25272), .A2(n19797), .Z(n6307) );
  XOR2_X1 U19051 ( .A1(n6310), .A2(n6309), .Z(n6308) );
  XOR2_X1 U19052 ( .A1(n22620), .A2(n22488), .Z(n6309) );
  INV_X2 U19056 ( .I(n18574), .ZN(n26893) );
  XOR2_X1 U19063 ( .A1(n28909), .A2(n6319), .Z(n6318) );
  XOR2_X1 U19064 ( .A1(n10343), .A2(n29849), .Z(n6319) );
  XOR2_X1 U19067 ( .A1(n6320), .A2(n33811), .Z(Ciphertext[53]) );
  NAND2_X1 U19068 ( .A1(n9913), .A2(n38200), .ZN(n6323) );
  XOR2_X1 U19070 ( .A1(n6325), .A2(n20047), .Z(n6324) );
  XOR2_X1 U19074 ( .A1(n6329), .A2(n14979), .Z(n6328) );
  INV_X2 U19076 ( .I(n6331), .ZN(n7834) );
  NOR2_X1 U19082 ( .A1(n32091), .A2(n6756), .ZN(n6706) );
  NOR2_X1 U19085 ( .A1(n9105), .A2(n9913), .ZN(n6339) );
  NAND2_X2 U19087 ( .A1(n29472), .A2(n29469), .ZN(n29477) );
  NAND2_X1 U19088 ( .A1(n38629), .A2(n34695), .ZN(n28112) );
  XOR2_X1 U19092 ( .A1(n6351), .A2(n16606), .Z(n16605) );
  OAI21_X1 U19093 ( .A1(n39495), .A2(n10211), .B(n33148), .ZN(n19169) );
  XOR2_X1 U19094 ( .A1(n6352), .A2(n24325), .Z(n15989) );
  NOR2_X1 U19095 ( .A1(n6355), .A2(n34969), .ZN(n8538) );
  NAND2_X1 U19096 ( .A1(n6355), .A2(n34969), .ZN(n8642) );
  XOR2_X1 U19105 ( .A1(n23885), .A2(n39161), .Z(n6360) );
  XOR2_X1 U19115 ( .A1(n22542), .A2(n19952), .Z(n6368) );
  XNOR2_X1 U19116 ( .A1(n22488), .A2(n19254), .ZN(n22372) );
  XOR2_X1 U19118 ( .A1(n13564), .A2(n7659), .Z(n18153) );
  AOI21_X2 U19127 ( .A1(n26749), .A2(n11682), .B(n6383), .ZN(n13569) );
  XOR2_X1 U19130 ( .A1(n28850), .A2(n6384), .Z(n29031) );
  XOR2_X1 U19131 ( .A1(n31599), .A2(n19808), .Z(n6387) );
  XOR2_X1 U19132 ( .A1(n6389), .A2(n6467), .Z(n20801) );
  XOR2_X1 U19135 ( .A1(n6395), .A2(n6392), .Z(n7281) );
  XOR2_X1 U19136 ( .A1(n6394), .A2(n6393), .Z(n6392) );
  XOR2_X1 U19137 ( .A1(n27710), .A2(n1707), .Z(n6393) );
  XOR2_X1 U19138 ( .A1(n5625), .A2(n21093), .Z(n6394) );
  NAND3_X2 U19142 ( .A1(n17312), .A2(n6397), .A3(n6396), .ZN(n26519) );
  OAI21_X2 U19143 ( .A1(n6399), .A2(n17311), .B(n6398), .ZN(n26259) );
  NAND3_X1 U19148 ( .A1(n30078), .A2(n20078), .A3(n3815), .ZN(n30074) );
  XOR2_X1 U19155 ( .A1(n6413), .A2(n26476), .Z(n6412) );
  AOI21_X2 U19164 ( .A1(n15457), .A2(n19892), .B(n33318), .ZN(n10712) );
  XOR2_X1 U19167 ( .A1(n21108), .A2(n6428), .Z(n6427) );
  XOR2_X1 U19169 ( .A1(n34091), .A2(n29138), .Z(n6430) );
  XOR2_X1 U19170 ( .A1(n6431), .A2(n6432), .Z(n6991) );
  XOR2_X1 U19171 ( .A1(n34829), .A2(n30006), .Z(n6431) );
  XOR2_X1 U19172 ( .A1(n15368), .A2(n13289), .Z(n6432) );
  XOR2_X1 U19173 ( .A1(n6433), .A2(n19761), .Z(n29248) );
  XOR2_X1 U19174 ( .A1(n6433), .A2(n19839), .Z(n28785) );
  XOR2_X1 U19176 ( .A1(n18886), .A2(n769), .Z(n6436) );
  INV_X2 U19179 ( .I(n13258), .ZN(n7062) );
  INV_X1 U19185 ( .I(Key[134]), .ZN(n6447) );
  XOR2_X1 U19193 ( .A1(n26335), .A2(n9554), .Z(n6455) );
  XOR2_X1 U19195 ( .A1(n6458), .A2(n6457), .Z(n6456) );
  XOR2_X1 U19199 ( .A1(n25274), .A2(n6461), .Z(n6460) );
  XOR2_X1 U19201 ( .A1(n23707), .A2(n6462), .Z(n6881) );
  INV_X2 U19207 ( .I(n20801), .ZN(n24244) );
  XOR2_X1 U19208 ( .A1(n6468), .A2(n23906), .Z(n6467) );
  XOR2_X1 U19212 ( .A1(n27626), .A2(n6471), .Z(n6470) );
  AOI21_X1 U19215 ( .A1(n6481), .A2(n6480), .B(n6479), .ZN(n16249) );
  NOR3_X1 U19216 ( .A1(n31534), .A2(n29237), .A3(n14933), .ZN(n6479) );
  OAI21_X1 U19217 ( .A1(n29237), .A2(n1387), .B(n1388), .ZN(n6480) );
  NAND3_X1 U19218 ( .A1(n29228), .A2(n8728), .A3(n38945), .ZN(n6481) );
  INV_X2 U19219 ( .I(n6484), .ZN(n19543) );
  XNOR2_X1 U19220 ( .A1(Plaintext[74]), .A2(Key[74]), .ZN(n6484) );
  NAND2_X2 U19221 ( .A1(n9328), .A2(n9327), .ZN(n28768) );
  NAND2_X1 U19223 ( .A1(n30067), .A2(n31120), .ZN(n6486) );
  NAND2_X2 U19226 ( .A1(n23818), .A2(n13881), .ZN(n23796) );
  INV_X2 U19229 ( .I(n6493), .ZN(n14562) );
  NAND2_X2 U19232 ( .A1(n15343), .A2(n6497), .ZN(n18762) );
  INV_X1 U19235 ( .I(n19455), .ZN(n27276) );
  NAND2_X1 U19236 ( .A1(n20027), .A2(n37480), .ZN(n6509) );
  XOR2_X1 U19239 ( .A1(n22597), .A2(n6512), .Z(n6511) );
  XOR2_X1 U19240 ( .A1(n12243), .A2(n19905), .Z(n6512) );
  XOR2_X1 U19241 ( .A1(n22658), .A2(n18634), .Z(n6513) );
  XOR2_X1 U19242 ( .A1(n11541), .A2(n5203), .Z(n22658) );
  XOR2_X1 U19246 ( .A1(n12839), .A2(n18296), .Z(n6525) );
  XOR2_X1 U19248 ( .A1(n6530), .A2(n6528), .Z(n19576) );
  XOR2_X1 U19250 ( .A1(n23794), .A2(n1699), .Z(n6531) );
  XOR2_X1 U19252 ( .A1(n6536), .A2(n28820), .Z(n6535) );
  NAND2_X2 U19256 ( .A1(n24717), .A2(n6944), .ZN(n24724) );
  NOR2_X2 U19257 ( .A1(n6543), .A2(n19580), .ZN(n25862) );
  XOR2_X1 U19259 ( .A1(n10705), .A2(n22448), .Z(n6544) );
  XOR2_X1 U19260 ( .A1(n57), .A2(n22784), .Z(n22448) );
  XOR2_X1 U19267 ( .A1(n27413), .A2(n11365), .Z(n6549) );
  XOR2_X1 U19274 ( .A1(n6562), .A2(n6563), .Z(n18602) );
  XOR2_X1 U19275 ( .A1(n31581), .A2(n23785), .Z(n6562) );
  XOR2_X1 U19276 ( .A1(n23316), .A2(n6564), .Z(n6563) );
  XOR2_X1 U19285 ( .A1(n6817), .A2(n6580), .Z(n6581) );
  XOR2_X1 U19286 ( .A1(n6633), .A2(n6632), .Z(n6580) );
  XOR2_X1 U19287 ( .A1(n6630), .A2(n17513), .Z(n6817) );
  OAI21_X2 U19292 ( .A1(n14665), .A2(n15702), .B(n14012), .ZN(n10635) );
  NAND2_X2 U19294 ( .A1(n6587), .A2(n6586), .ZN(n28807) );
  NAND2_X1 U19295 ( .A1(n28288), .A2(n11375), .ZN(n6586) );
  NAND2_X1 U19296 ( .A1(n6590), .A2(n13712), .ZN(n25970) );
  XOR2_X1 U19304 ( .A1(n13919), .A2(n13918), .Z(n6595) );
  OAI21_X1 U19310 ( .A1(n6600), .A2(n11861), .B(n16510), .ZN(n6599) );
  XOR2_X1 U19316 ( .A1(n22442), .A2(n6609), .Z(n6608) );
  XOR2_X1 U19317 ( .A1(n11201), .A2(n1661), .Z(n6609) );
  XOR2_X1 U19321 ( .A1(n22484), .A2(n22459), .Z(n22441) );
  INV_X1 U19326 ( .I(n26088), .ZN(n20545) );
  AOI21_X1 U19328 ( .A1(n29979), .A2(n29980), .B(n6623), .ZN(n18200) );
  NAND2_X1 U19331 ( .A1(n6623), .A2(n29979), .ZN(n6622) );
  NAND2_X2 U19332 ( .A1(n17983), .A2(n29961), .ZN(n6623) );
  XOR2_X1 U19333 ( .A1(n6624), .A2(n6627), .Z(n7364) );
  XOR2_X1 U19334 ( .A1(n24013), .A2(n6625), .Z(n6624) );
  XOR2_X1 U19335 ( .A1(n24079), .A2(n6626), .Z(n6625) );
  XOR2_X1 U19337 ( .A1(n6628), .A2(n19623), .Z(n6627) );
  OR2_X1 U19338 ( .A1(n6629), .A2(n8082), .Z(n6697) );
  XOR2_X1 U19343 ( .A1(n17189), .A2(n22508), .Z(n6632) );
  NAND2_X1 U19345 ( .A1(n6772), .A2(n6771), .ZN(n6634) );
  NOR2_X2 U19347 ( .A1(n10648), .A2(n10988), .ZN(n10987) );
  XOR2_X1 U19349 ( .A1(n6644), .A2(n16886), .Z(n19855) );
  OAI21_X1 U19355 ( .A1(n10096), .A2(n29870), .B(n20793), .ZN(n20895) );
  MUX2_X1 U19360 ( .I0(n841), .I1(n6656), .S(n25669), .Z(n19971) );
  NOR3_X1 U19365 ( .A1(n38529), .A2(n28695), .A3(n28696), .ZN(n10680) );
  NAND2_X2 U19367 ( .A1(n10304), .A2(n10302), .ZN(n29054) );
  OR2_X1 U19373 ( .A1(n1486), .A2(n34001), .Z(n6668) );
  XOR2_X1 U19382 ( .A1(n12101), .A2(n6676), .Z(n9595) );
  XOR2_X1 U19383 ( .A1(n22703), .A2(n19676), .Z(n6676) );
  XOR2_X1 U19385 ( .A1(n2281), .A2(n27736), .Z(n6677) );
  INV_X2 U19395 ( .I(n4378), .ZN(n30071) );
  XOR2_X1 U19397 ( .A1(n10653), .A2(n1738), .Z(n6688) );
  XOR2_X1 U19401 ( .A1(n12763), .A2(n10059), .Z(n16217) );
  INV_X2 U19402 ( .I(n8532), .ZN(n16639) );
  INV_X1 U19404 ( .I(n8082), .ZN(n6698) );
  XOR2_X1 U19409 ( .A1(n22634), .A2(n5203), .Z(n6711) );
  NAND2_X2 U19411 ( .A1(n1275), .A2(n39699), .ZN(n6715) );
  XOR2_X1 U19412 ( .A1(n8402), .A2(n11755), .Z(n6717) );
  XOR2_X1 U19417 ( .A1(n38161), .A2(n29394), .Z(n28372) );
  XOR2_X1 U19418 ( .A1(n30856), .A2(n38161), .Z(n29138) );
  XOR2_X1 U19424 ( .A1(n26370), .A2(n26323), .Z(n12228) );
  AOI21_X2 U19429 ( .A1(n27297), .A2(n35473), .B(n27296), .ZN(n27525) );
  XOR2_X1 U19431 ( .A1(n25153), .A2(n20803), .Z(n6728) );
  XOR2_X1 U19433 ( .A1(n25152), .A2(n20805), .Z(n6729) );
  OAI21_X1 U19437 ( .A1(n21654), .A2(n33771), .B(n6732), .ZN(n11849) );
  XOR2_X1 U19447 ( .A1(n26510), .A2(n36579), .Z(n26172) );
  XOR2_X1 U19449 ( .A1(n26233), .A2(n25930), .Z(n6739) );
  XOR2_X1 U19450 ( .A1(n26157), .A2(n26389), .Z(n26233) );
  XOR2_X1 U19452 ( .A1(n16254), .A2(n22693), .Z(n6741) );
  XOR2_X1 U19460 ( .A1(n16066), .A2(n6752), .Z(n6751) );
  XOR2_X1 U19461 ( .A1(n27729), .A2(n37101), .Z(n6752) );
  XOR2_X1 U19462 ( .A1(n27515), .A2(n10766), .Z(n6753) );
  XOR2_X1 U19463 ( .A1(n5284), .A2(n19904), .Z(n18843) );
  XOR2_X1 U19464 ( .A1(n6014), .A2(n29649), .Z(n18941) );
  XOR2_X1 U19465 ( .A1(n5284), .A2(n19677), .Z(n22427) );
  NAND3_X1 U19466 ( .A1(n36376), .A2(n36920), .A3(n38884), .ZN(n8109) );
  XOR2_X1 U19468 ( .A1(n6757), .A2(n19877), .Z(n25865) );
  XOR2_X1 U19470 ( .A1(n38584), .A2(n6757), .Z(n13814) );
  XOR2_X1 U19472 ( .A1(n38195), .A2(n19874), .Z(n28306) );
  XOR2_X1 U19474 ( .A1(n19725), .A2(n61), .Z(n25075) );
  XOR2_X1 U19479 ( .A1(n6765), .A2(n34815), .Z(n6764) );
  XOR2_X1 U19480 ( .A1(n1613), .A2(n23900), .Z(n6765) );
  NAND3_X1 U19490 ( .A1(n12567), .A2(n22162), .A3(n19890), .ZN(n6771) );
  INV_X1 U19491 ( .I(n6773), .ZN(n6772) );
  INV_X2 U19493 ( .I(n29943), .ZN(n16353) );
  NOR2_X1 U19495 ( .A1(n6776), .A2(n9727), .ZN(n6775) );
  XOR2_X1 U19501 ( .A1(n35379), .A2(n19875), .Z(n6778) );
  XOR2_X1 U19502 ( .A1(n6782), .A2(n6781), .Z(n6780) );
  XOR2_X1 U19503 ( .A1(n6527), .A2(n23829), .Z(n6782) );
  XOR2_X1 U19507 ( .A1(n22689), .A2(n2234), .Z(n7346) );
  INV_X2 U19509 ( .I(n6801), .ZN(n12162) );
  XOR2_X1 U19510 ( .A1(n24946), .A2(n11689), .Z(n6802) );
  XOR2_X1 U19516 ( .A1(n7352), .A2(n25123), .Z(n25011) );
  NOR2_X1 U19518 ( .A1(n23502), .A2(n32366), .ZN(n23048) );
  OAI21_X2 U19521 ( .A1(n19104), .A2(n21622), .B(n18900), .ZN(n22364) );
  XOR2_X1 U19527 ( .A1(Plaintext[21]), .A2(Key[21]), .Z(n8267) );
  XOR2_X1 U19531 ( .A1(n12442), .A2(n15158), .Z(n6825) );
  XOR2_X1 U19538 ( .A1(n6835), .A2(n6834), .Z(n6836) );
  INV_X2 U19540 ( .I(n6836), .ZN(n30055) );
  INV_X1 U19542 ( .I(n9310), .ZN(n27271) );
  XOR2_X1 U19545 ( .A1(n12730), .A2(n31562), .Z(n11908) );
  XOR2_X1 U19546 ( .A1(n31562), .A2(n1718), .Z(n16753) );
  XOR2_X1 U19547 ( .A1(n31562), .A2(n19761), .Z(n13846) );
  NAND2_X1 U19552 ( .A1(n6851), .A2(n20018), .ZN(n12994) );
  OAI21_X1 U19554 ( .A1(n18461), .A2(n13153), .B(n6851), .ZN(n16121) );
  XOR2_X1 U19556 ( .A1(n29031), .A2(n6853), .Z(n6852) );
  INV_X1 U19568 ( .I(n34001), .ZN(n27196) );
  NAND2_X1 U19570 ( .A1(n27368), .A2(n5772), .ZN(n6874) );
  XOR2_X1 U19571 ( .A1(n6879), .A2(n6878), .Z(n6877) );
  XOR2_X1 U19572 ( .A1(n26234), .A2(n1362), .Z(n6878) );
  XOR2_X1 U19573 ( .A1(n208), .A2(n6881), .Z(n6880) );
  NAND2_X1 U19577 ( .A1(n31533), .A2(n16803), .ZN(n10294) );
  NAND2_X1 U19578 ( .A1(n31533), .A2(n967), .ZN(n17885) );
  XOR2_X1 U19580 ( .A1(n6886), .A2(n12076), .Z(n8069) );
  XOR2_X1 U19581 ( .A1(n25126), .A2(n6887), .Z(n6886) );
  XOR2_X1 U19582 ( .A1(n25080), .A2(n19733), .Z(n6887) );
  XOR2_X1 U19583 ( .A1(n25259), .A2(n25216), .Z(n25126) );
  NAND2_X2 U19585 ( .A1(n10826), .A2(n10824), .ZN(n6892) );
  XOR2_X1 U19588 ( .A1(n35112), .A2(n22615), .Z(n22479) );
  XOR2_X1 U19591 ( .A1(n10424), .A2(n6895), .Z(n9808) );
  XOR2_X1 U19592 ( .A1(n35053), .A2(n1697), .Z(n6895) );
  XOR2_X1 U19598 ( .A1(n7416), .A2(n11391), .Z(n6905) );
  NAND2_X1 U19602 ( .A1(n6908), .A2(n27389), .ZN(n26428) );
  XOR2_X1 U19611 ( .A1(n6923), .A2(n25262), .Z(n6922) );
  XOR2_X1 U19613 ( .A1(n15779), .A2(n13711), .Z(n6924) );
  XOR2_X1 U19619 ( .A1(n6930), .A2(n30006), .Z(n29068) );
  XOR2_X1 U19620 ( .A1(n6930), .A2(n29671), .Z(n29028) );
  XOR2_X1 U19622 ( .A1(n38703), .A2(n29538), .Z(n20136) );
  NAND3_X2 U19625 ( .A1(n10476), .A2(n10475), .A3(n25378), .ZN(n7133) );
  XOR2_X1 U19627 ( .A1(n19384), .A2(n26244), .Z(n9490) );
  XOR2_X1 U19631 ( .A1(n6942), .A2(n6941), .Z(n6940) );
  XOR2_X1 U19632 ( .A1(n23658), .A2(n29357), .Z(n6941) );
  XOR2_X1 U19633 ( .A1(n33322), .A2(n24002), .Z(n6942) );
  OAI21_X1 U19636 ( .A1(n24590), .A2(n5056), .B(n6944), .ZN(n16077) );
  NOR2_X2 U19640 ( .A1(n8496), .A2(n9165), .ZN(n21995) );
  NOR2_X1 U19641 ( .A1(n36303), .A2(n39489), .ZN(n6948) );
  INV_X1 U19642 ( .I(n17478), .ZN(n10560) );
  XOR2_X1 U19643 ( .A1(n23888), .A2(n18006), .Z(n6951) );
  XOR2_X1 U19644 ( .A1(n23988), .A2(n23609), .Z(n6952) );
  XNOR2_X1 U19645 ( .A1(n17478), .A2(n23762), .ZN(n23745) );
  AOI21_X2 U19648 ( .A1(n6956), .A2(n23828), .B(n6955), .ZN(n24696) );
  NAND2_X1 U19649 ( .A1(n39196), .A2(n24805), .ZN(n6957) );
  OAI22_X1 U19666 ( .A1(n6981), .A2(n22157), .B1(n22225), .B2(n6982), .ZN(
        n22087) );
  NAND2_X1 U19667 ( .A1(n6982), .A2(n7357), .ZN(n6981) );
  NAND2_X1 U19669 ( .A1(n8275), .A2(n22364), .ZN(n6982) );
  NAND2_X2 U19670 ( .A1(n21625), .A2(n15468), .ZN(n8275) );
  XOR2_X1 U19674 ( .A1(n6987), .A2(n6986), .Z(n6985) );
  XOR2_X1 U19675 ( .A1(n23903), .A2(n29476), .Z(n6986) );
  NAND3_X2 U19677 ( .A1(n6994), .A2(n11842), .A3(n6992), .ZN(n23755) );
  XOR2_X1 U19680 ( .A1(n24982), .A2(n29223), .Z(n6996) );
  NAND3_X1 U19685 ( .A1(n1595), .A2(n1127), .A3(n15385), .ZN(n7000) );
  OAI21_X2 U19690 ( .A1(n7007), .A2(n7006), .B(n7005), .ZN(n9144) );
  NAND2_X2 U19694 ( .A1(n21213), .A2(n7009), .ZN(n23331) );
  AOI21_X1 U19703 ( .A1(n24804), .A2(n24829), .B(n15664), .ZN(n10521) );
  INV_X2 U19705 ( .I(n14367), .ZN(n23042) );
  NAND2_X2 U19707 ( .A1(n28565), .A2(n28564), .ZN(n28983) );
  XOR2_X1 U19711 ( .A1(n19571), .A2(n29303), .Z(n7032) );
  XOR2_X1 U19716 ( .A1(n7039), .A2(n7038), .Z(n7037) );
  XOR2_X1 U19720 ( .A1(n37023), .A2(n22167), .Z(n7040) );
  NAND2_X1 U19726 ( .A1(n7046), .A2(n33713), .ZN(n18951) );
  INV_X1 U19727 ( .I(n21795), .ZN(n7047) );
  XOR2_X1 U19731 ( .A1(n27672), .A2(n29229), .Z(n7060) );
  NAND3_X1 U19738 ( .A1(n10906), .A2(n28686), .A3(n36663), .ZN(n28587) );
  OAI21_X1 U19741 ( .A1(n24789), .A2(n31161), .B(n20039), .ZN(n7066) );
  XOR2_X1 U19747 ( .A1(n19606), .A2(n29411), .Z(n7069) );
  XOR2_X1 U19748 ( .A1(n29824), .A2(n19722), .Z(n7070) );
  XOR2_X1 U19755 ( .A1(n10794), .A2(n1370), .Z(n7089) );
  NAND2_X1 U19770 ( .A1(n9875), .A2(n27197), .ZN(n12031) );
  XOR2_X1 U19775 ( .A1(n12838), .A2(n29849), .Z(n7101) );
  AOI21_X1 U19780 ( .A1(n20376), .A2(n19017), .B(n1154), .ZN(n7104) );
  XOR2_X1 U19785 ( .A1(n23970), .A2(n39482), .Z(n7113) );
  XOR2_X1 U19790 ( .A1(n1658), .A2(n19127), .Z(n7119) );
  INV_X2 U19792 ( .I(n18732), .ZN(n28205) );
  XOR2_X1 U19793 ( .A1(n7120), .A2(n7123), .Z(n22864) );
  XOR2_X1 U19796 ( .A1(n7510), .A2(n17153), .Z(n7123) );
  INV_X2 U19797 ( .I(n7124), .ZN(n7304) );
  XNOR2_X1 U19798 ( .A1(Plaintext[20]), .A2(Key[20]), .ZN(n7124) );
  XOR2_X1 U19799 ( .A1(n24925), .A2(n15912), .Z(n18584) );
  XOR2_X1 U19800 ( .A1(n15912), .A2(n30065), .Z(n25035) );
  XOR2_X1 U19803 ( .A1(n7127), .A2(n7126), .Z(n7125) );
  XOR2_X1 U19804 ( .A1(n24040), .A2(n1362), .Z(n7126) );
  XOR2_X1 U19809 ( .A1(n26244), .A2(n1096), .Z(n10317) );
  NOR2_X1 U19811 ( .A1(n15121), .A2(n7134), .ZN(n15021) );
  NAND2_X2 U19814 ( .A1(n22211), .A2(n22210), .ZN(n22665) );
  NAND2_X1 U19817 ( .A1(n7146), .A2(n23229), .ZN(n7145) );
  XOR2_X1 U19820 ( .A1(n25254), .A2(n25001), .Z(n7152) );
  XOR2_X1 U19821 ( .A1(n20333), .A2(n38148), .Z(n25001) );
  XOR2_X1 U19822 ( .A1(n25002), .A2(n10905), .Z(n7153) );
  XOR2_X1 U19824 ( .A1(n25118), .A2(n24982), .Z(n25002) );
  XOR2_X1 U19833 ( .A1(n57), .A2(n7162), .Z(n7161) );
  AOI21_X2 U19834 ( .A1(n34086), .A2(n7167), .B(n7166), .ZN(n17469) );
  XOR2_X1 U19839 ( .A1(n15216), .A2(n18905), .Z(n7180) );
  XOR2_X1 U19844 ( .A1(n39631), .A2(n1413), .Z(n7182) );
  NOR2_X1 U19853 ( .A1(n13088), .A2(n7195), .ZN(n13951) );
  XOR2_X1 U19860 ( .A1(n1662), .A2(n17195), .Z(n7200) );
  XOR2_X1 U19862 ( .A1(n19071), .A2(n7202), .Z(n9894) );
  XOR2_X1 U19863 ( .A1(n19656), .A2(n29229), .Z(n7202) );
  XOR2_X1 U19864 ( .A1(n7203), .A2(n7206), .Z(n17764) );
  XOR2_X1 U19865 ( .A1(n25313), .A2(n7204), .Z(n7203) );
  XOR2_X1 U19866 ( .A1(n39295), .A2(n24926), .Z(n7204) );
  XOR2_X1 U19867 ( .A1(n35237), .A2(n20828), .Z(n7206) );
  NAND2_X1 U19869 ( .A1(n29952), .A2(n7208), .ZN(n29953) );
  XOR2_X1 U19873 ( .A1(n3082), .A2(n15617), .Z(n8285) );
  XOR2_X1 U19874 ( .A1(n35320), .A2(n3082), .Z(n20137) );
  AND2_X1 U19875 ( .A1(n19017), .A2(n1154), .Z(n22149) );
  OAI21_X2 U19878 ( .A1(n7232), .A2(n7230), .B(n26998), .ZN(n27503) );
  NAND2_X2 U19879 ( .A1(n37393), .A2(n33263), .ZN(n25940) );
  INV_X2 U19882 ( .I(n25719), .ZN(n19237) );
  XNOR2_X1 U19883 ( .A1(n27854), .A2(n38158), .ZN(n27628) );
  XOR2_X1 U19884 ( .A1(n10782), .A2(n7257), .Z(n7256) );
  XOR2_X1 U19886 ( .A1(n27674), .A2(n1467), .Z(n7257) );
  NAND2_X1 U19888 ( .A1(n37160), .A2(n32722), .ZN(n14840) );
  NAND2_X1 U19890 ( .A1(n1147), .A2(n7266), .ZN(n23191) );
  NAND3_X1 U19892 ( .A1(n7267), .A2(n24799), .A3(n17350), .ZN(n16570) );
  AOI21_X1 U19893 ( .A1(n7267), .A2(n19679), .B(n33409), .ZN(n8575) );
  NAND2_X2 U19896 ( .A1(n17980), .A2(n17982), .ZN(n29980) );
  XOR2_X1 U19898 ( .A1(n16667), .A2(n17310), .Z(n7275) );
  XOR2_X1 U19899 ( .A1(n37023), .A2(n7277), .Z(n7276) );
  INV_X2 U19901 ( .I(n12951), .ZN(n19857) );
  NAND2_X1 U19903 ( .A1(n21383), .A2(n21384), .ZN(n19911) );
  NAND2_X1 U19912 ( .A1(n23639), .A2(n35232), .ZN(n23470) );
  AND2_X1 U19914 ( .A1(n17648), .A2(n23617), .Z(n12426) );
  NAND2_X1 U19923 ( .A1(n27278), .A2(n7291), .ZN(n7300) );
  INV_X1 U19928 ( .I(n10413), .ZN(n7737) );
  XNOR2_X1 U19932 ( .A1(n39063), .A2(n19851), .ZN(n17921) );
  XOR2_X1 U19937 ( .A1(n7316), .A2(n7667), .Z(n28841) );
  XOR2_X1 U19938 ( .A1(n29145), .A2(n14956), .Z(n7316) );
  OAI21_X1 U19947 ( .A1(n20538), .A2(n20342), .B(n7318), .ZN(n10409) );
  NAND2_X2 U19950 ( .A1(n18641), .A2(n18640), .ZN(n27830) );
  NOR2_X1 U19952 ( .A1(n9276), .A2(n17087), .ZN(n9849) );
  AND2_X1 U19955 ( .A1(n18406), .A2(n9413), .Z(n11835) );
  XOR2_X1 U19957 ( .A1(n17455), .A2(n19919), .Z(n17396) );
  XOR2_X1 U19958 ( .A1(n23912), .A2(n29857), .Z(n10312) );
  XOR2_X1 U19966 ( .A1(n11318), .A2(n24988), .Z(n7329) );
  NOR2_X2 U19967 ( .A1(n13922), .A2(n20356), .ZN(n9626) );
  NAND2_X1 U19969 ( .A1(n34004), .A2(n35269), .ZN(n9650) );
  XOR2_X1 U19975 ( .A1(n18267), .A2(n26368), .Z(n26832) );
  NAND2_X1 U19976 ( .A1(n8000), .A2(n17934), .ZN(n12844) );
  AND2_X1 U19983 ( .A1(n24335), .A2(n545), .Z(n14581) );
  XOR2_X1 U19987 ( .A1(n22755), .A2(n704), .Z(n7341) );
  OAI21_X2 U19988 ( .A1(n27661), .A2(n27557), .B(n10801), .ZN(n27648) );
  NOR2_X2 U19991 ( .A1(n26853), .A2(n7349), .ZN(n27320) );
  NOR3_X1 U19992 ( .A1(n26944), .A2(n19425), .A3(n15670), .ZN(n7349) );
  XOR2_X1 U19999 ( .A1(n27606), .A2(n18817), .Z(n7353) );
  XOR2_X1 U20000 ( .A1(n22712), .A2(n22617), .Z(n13840) );
  INV_X1 U20001 ( .I(n14991), .ZN(n14990) );
  XOR2_X1 U20006 ( .A1(n24060), .A2(n7360), .Z(n7359) );
  NAND3_X1 U20019 ( .A1(n8568), .A2(n15173), .A3(n36708), .ZN(n7362) );
  INV_X2 U20022 ( .I(n25782), .ZN(n26108) );
  XOR2_X1 U20030 ( .A1(n334), .A2(n30169), .Z(n7698) );
  OR2_X1 U20037 ( .A1(n29794), .A2(n18257), .Z(n29787) );
  XOR2_X1 U20045 ( .A1(n25000), .A2(n810), .Z(n7380) );
  XOR2_X1 U20047 ( .A1(n28985), .A2(n765), .Z(n7382) );
  MUX2_X1 U20052 ( .I0(n27363), .I1(n34001), .S(n21101), .Z(n27056) );
  INV_X1 U20056 ( .I(n13004), .ZN(n7393) );
  NOR2_X1 U20058 ( .A1(n18377), .A2(n22991), .ZN(n8011) );
  OAI21_X1 U20060 ( .A1(n9460), .A2(n9459), .B(n10220), .ZN(n10219) );
  OR2_X1 U20072 ( .A1(n10634), .A2(n18072), .Z(n21120) );
  XNOR2_X1 U20074 ( .A1(n26246), .A2(n35212), .ZN(n26166) );
  AND2_X1 U20079 ( .A1(n20734), .A2(n31452), .Z(n8927) );
  INV_X1 U20082 ( .I(n20243), .ZN(n15058) );
  XOR2_X1 U20100 ( .A1(n27825), .A2(n27540), .Z(n27667) );
  XOR2_X1 U20104 ( .A1(n8199), .A2(n11475), .Z(n10970) );
  XOR2_X1 U20106 ( .A1(n8401), .A2(n27577), .Z(n8403) );
  AOI21_X1 U20109 ( .A1(n7303), .A2(n38200), .B(n969), .ZN(n29466) );
  AND2_X1 U20113 ( .A1(n29662), .A2(n19297), .Z(n29654) );
  XOR2_X1 U20115 ( .A1(n23680), .A2(n7917), .Z(n10279) );
  NOR2_X1 U20118 ( .A1(n26133), .A2(n13678), .ZN(n13677) );
  NAND2_X1 U20119 ( .A1(n20807), .A2(n20696), .ZN(n11963) );
  XOR2_X1 U20122 ( .A1(n22435), .A2(n12598), .Z(n7498) );
  NOR2_X2 U20123 ( .A1(n7443), .A2(n9148), .ZN(n17184) );
  XOR2_X1 U20124 ( .A1(n1667), .A2(n22766), .Z(n22606) );
  OAI21_X2 U20125 ( .A1(n17409), .A2(n17408), .B(n17407), .ZN(n22766) );
  XOR2_X1 U20127 ( .A1(n29070), .A2(n1409), .Z(n20675) );
  INV_X1 U20128 ( .I(n25897), .ZN(n16444) );
  OR2_X1 U20129 ( .A1(n29218), .A2(n29219), .Z(n13104) );
  XOR2_X1 U20138 ( .A1(n7451), .A2(n15432), .Z(Ciphertext[72]) );
  AOI22_X1 U20139 ( .A1(n20126), .A2(n29618), .B1(n29601), .B2(n29616), .ZN(
        n7451) );
  OR3_X1 U20146 ( .A1(n34906), .A2(n24733), .A3(n24839), .Z(n11367) );
  AND2_X1 U20149 ( .A1(n22900), .A2(n2350), .Z(n14483) );
  XOR2_X1 U20152 ( .A1(n26497), .A2(n26496), .Z(n26502) );
  INV_X2 U20154 ( .I(n7459), .ZN(n8818) );
  INV_X2 U20157 ( .I(n7462), .ZN(n14459) );
  OAI21_X1 U20163 ( .A1(n17262), .A2(n29567), .B(n1053), .ZN(n13926) );
  OR2_X1 U20165 ( .A1(n27233), .A2(n12306), .Z(n7472) );
  NAND2_X1 U20172 ( .A1(n17939), .A2(n16534), .ZN(n16533) );
  AOI21_X1 U20173 ( .A1(n14582), .A2(n30323), .B(n16533), .ZN(n16532) );
  INV_X1 U20174 ( .I(n16179), .ZN(n24294) );
  NAND2_X1 U20175 ( .A1(n25937), .A2(n1105), .ZN(n14133) );
  XOR2_X1 U20176 ( .A1(n13035), .A2(n18800), .Z(n8564) );
  XOR2_X1 U20177 ( .A1(n26396), .A2(n12649), .Z(n19051) );
  NAND3_X2 U20178 ( .A1(n25478), .A2(n11063), .A3(n25460), .ZN(n11064) );
  AOI22_X1 U20180 ( .A1(n17318), .A2(n1389), .B1(n17317), .B2(n29437), .ZN(
        n7572) );
  XOR2_X1 U20184 ( .A1(n27728), .A2(n17721), .Z(n8975) );
  INV_X2 U20190 ( .I(n7492), .ZN(n25540) );
  INV_X1 U20191 ( .I(n1283), .ZN(n13185) );
  AND2_X1 U20193 ( .A1(n36162), .A2(n3985), .Z(n25373) );
  AOI21_X1 U20199 ( .A1(n7502), .A2(n29633), .B(n29700), .ZN(n29198) );
  AND3_X1 U20206 ( .A1(n13770), .A2(n26811), .A3(n26810), .Z(n7628) );
  XNOR2_X1 U20208 ( .A1(n31823), .A2(n18273), .ZN(n10546) );
  XOR2_X1 U20210 ( .A1(n32298), .A2(n27830), .Z(n27657) );
  XOR2_X1 U20213 ( .A1(n7507), .A2(n29964), .Z(Ciphertext[132]) );
  OAI22_X1 U20214 ( .A1(n29963), .A2(n29977), .B1(n29962), .B2(n1170), .ZN(
        n7507) );
  NOR2_X2 U20224 ( .A1(n31569), .A2(n29927), .ZN(n29923) );
  NAND2_X1 U20234 ( .A1(n32865), .A2(n11700), .ZN(n19164) );
  AND2_X1 U20237 ( .A1(n30158), .A2(n20541), .Z(n14539) );
  OAI22_X2 U20238 ( .A1(n21553), .A2(n21908), .B1(n7526), .B2(n21645), .ZN(
        n19604) );
  OR2_X1 U20246 ( .A1(n22324), .A2(n22322), .Z(n11345) );
  NOR2_X1 U20252 ( .A1(n12168), .A2(n11330), .ZN(n7539) );
  XOR2_X1 U20254 ( .A1(n10668), .A2(n16591), .Z(n7543) );
  XOR2_X1 U20256 ( .A1(n29159), .A2(n7546), .Z(n28805) );
  XOR2_X1 U20257 ( .A1(n973), .A2(n29828), .Z(n7546) );
  XOR2_X1 U20258 ( .A1(n10156), .A2(n7547), .Z(n10155) );
  XOR2_X1 U20259 ( .A1(n28914), .A2(n7548), .Z(n7547) );
  NAND2_X2 U20260 ( .A1(n9382), .A2(n9381), .ZN(n9385) );
  NAND3_X1 U20261 ( .A1(n26635), .A2(n26634), .A3(n4748), .ZN(n26638) );
  INV_X4 U20263 ( .I(n10632), .ZN(n22342) );
  OR2_X1 U20270 ( .A1(n26976), .A2(n36262), .Z(n10853) );
  NAND2_X1 U20271 ( .A1(n9737), .A2(n13997), .ZN(n11124) );
  XOR2_X1 U20272 ( .A1(n26537), .A2(n26538), .Z(n8020) );
  NAND2_X1 U20280 ( .A1(n12526), .A2(n12525), .ZN(n12524) );
  XOR2_X1 U20287 ( .A1(n25072), .A2(n7569), .Z(n7762) );
  XOR2_X1 U20288 ( .A1(n25179), .A2(n35707), .Z(n7569) );
  XOR2_X1 U20289 ( .A1(n7570), .A2(n846), .Z(n7959) );
  XOR2_X1 U20290 ( .A1(n11374), .A2(n7571), .Z(n7570) );
  XOR2_X1 U20291 ( .A1(n7572), .A2(n17316), .Z(Ciphertext[44]) );
  XOR2_X1 U20293 ( .A1(n26276), .A2(n11902), .Z(n7573) );
  OAI21_X1 U20302 ( .A1(n19570), .A2(n19569), .B(n27286), .ZN(n11487) );
  XNOR2_X1 U20309 ( .A1(n29026), .A2(n14689), .ZN(n11405) );
  NAND3_X1 U20310 ( .A1(n5921), .A2(n29721), .A3(n20498), .ZN(n29713) );
  XOR2_X1 U20314 ( .A1(n7589), .A2(n19953), .Z(Ciphertext[94]) );
  XNOR2_X1 U20327 ( .A1(n27825), .A2(n35229), .ZN(n11031) );
  XOR2_X1 U20329 ( .A1(n20811), .A2(n28829), .Z(n16380) );
  XOR2_X1 U20330 ( .A1(n28991), .A2(n29247), .Z(n28829) );
  AND2_X1 U20344 ( .A1(n23550), .A2(n35191), .Z(n18617) );
  INV_X1 U20350 ( .I(n28523), .ZN(n12609) );
  XOR2_X1 U20352 ( .A1(n13247), .A2(n23995), .Z(n13246) );
  XOR2_X1 U20354 ( .A1(n23889), .A2(n32230), .Z(n23724) );
  XOR2_X1 U20356 ( .A1(n20101), .A2(n839), .Z(n14440) );
  OR2_X1 U20358 ( .A1(n13415), .A2(n34666), .Z(n18264) );
  XOR2_X1 U20363 ( .A1(n9120), .A2(n738), .Z(n7623) );
  AOI21_X1 U20373 ( .A1(n16722), .A2(n30109), .B(n1052), .ZN(n16721) );
  XOR2_X1 U20377 ( .A1(n19112), .A2(n23672), .Z(n7981) );
  XOR2_X1 U20379 ( .A1(n25161), .A2(n17457), .Z(n11161) );
  OAI22_X1 U20385 ( .A1(n11939), .A2(n15509), .B1(n8955), .B2(n15535), .ZN(
        n7637) );
  XOR2_X1 U20389 ( .A1(n18133), .A2(n28982), .Z(n28913) );
  OR2_X1 U20392 ( .A1(n1630), .A2(n23325), .Z(n19666) );
  XOR2_X1 U20399 ( .A1(n8563), .A2(n8564), .Z(n16327) );
  NAND3_X1 U20401 ( .A1(n1172), .A2(n13786), .A3(n38204), .ZN(n18231) );
  XOR2_X1 U20407 ( .A1(n7661), .A2(n26455), .Z(n26309) );
  XOR2_X1 U20412 ( .A1(n7663), .A2(n9270), .Z(n18923) );
  XOR2_X1 U20413 ( .A1(n18924), .A2(n27672), .Z(n7663) );
  XOR2_X1 U20417 ( .A1(n28710), .A2(n7665), .Z(n7664) );
  INV_X2 U20418 ( .I(n7666), .ZN(n10422) );
  NOR3_X1 U20422 ( .A1(n3989), .A2(n19467), .A3(n28255), .ZN(n9880) );
  NAND2_X1 U20433 ( .A1(n25769), .A2(n25943), .ZN(n7678) );
  XOR2_X1 U20434 ( .A1(n7681), .A2(n1362), .Z(Ciphertext[191]) );
  XNOR2_X1 U20438 ( .A1(n13243), .A2(n13242), .ZN(n7720) );
  XOR2_X1 U20444 ( .A1(n27539), .A2(n12495), .Z(n12494) );
  XOR2_X1 U20453 ( .A1(n9980), .A2(n12283), .Z(n22862) );
  XOR2_X1 U20459 ( .A1(n7698), .A2(n8585), .Z(n8586) );
  XOR2_X1 U20473 ( .A1(n25204), .A2(n1735), .Z(n24962) );
  AOI21_X2 U20474 ( .A1(n13893), .A2(n13894), .B(n8733), .ZN(n7710) );
  AND3_X1 U20484 ( .A1(n27048), .A2(n27047), .A3(n27046), .Z(n7716) );
  XNOR2_X1 U20493 ( .A1(n29253), .A2(n19730), .ZN(n10087) );
  NAND2_X1 U20494 ( .A1(n14132), .A2(n25813), .ZN(n7724) );
  OR3_X1 U20496 ( .A1(n1276), .A2(n1127), .A3(n24232), .Z(n18759) );
  NOR2_X1 U20497 ( .A1(n16924), .A2(n9178), .ZN(n20462) );
  OR2_X1 U20498 ( .A1(n11805), .A2(n35919), .Z(n26913) );
  NAND3_X2 U20507 ( .A1(n16312), .A2(n24268), .A3(n16311), .ZN(n24912) );
  XOR2_X1 U20509 ( .A1(n31627), .A2(n26287), .Z(n10967) );
  XOR2_X1 U20512 ( .A1(n31339), .A2(n35596), .Z(n22321) );
  XNOR2_X1 U20524 ( .A1(n38152), .A2(n19592), .ZN(n7801) );
  XOR2_X1 U20538 ( .A1(n14219), .A2(n16055), .Z(n23715) );
  XOR2_X1 U20549 ( .A1(n35505), .A2(n7287), .Z(n9093) );
  XOR2_X1 U20554 ( .A1(n7763), .A2(n18371), .Z(n8002) );
  XOR2_X1 U20557 ( .A1(n27813), .A2(n673), .Z(n7764) );
  OR2_X2 U20561 ( .A1(n29198), .A2(n7765), .Z(n29732) );
  OAI21_X1 U20562 ( .A1(n29197), .A2(n29702), .B(n34180), .ZN(n7765) );
  XOR2_X1 U20563 ( .A1(n12265), .A2(n12266), .Z(n12759) );
  OAI21_X1 U20565 ( .A1(n29611), .A2(n29618), .B(n9045), .ZN(n9044) );
  XOR2_X1 U20568 ( .A1(n7779), .A2(n7780), .Z(n26768) );
  XOR2_X1 U20569 ( .A1(n26442), .A2(n15750), .Z(n7779) );
  XOR2_X1 U20573 ( .A1(n18849), .A2(n1368), .Z(n7783) );
  XOR2_X1 U20576 ( .A1(n26324), .A2(n1237), .Z(n7785) );
  XOR2_X1 U20577 ( .A1(n20425), .A2(n7787), .Z(n7786) );
  XNOR2_X1 U20578 ( .A1(n26223), .A2(n26598), .ZN(n20425) );
  NOR2_X1 U20579 ( .A1(n5077), .A2(n22215), .ZN(n11202) );
  NAND2_X1 U20580 ( .A1(n9938), .A2(n5077), .ZN(n22009) );
  NAND2_X1 U20581 ( .A1(n15488), .A2(n5077), .ZN(n15487) );
  AOI21_X1 U20586 ( .A1(n30214), .A2(n14387), .B(n30217), .ZN(n7795) );
  NAND2_X1 U20587 ( .A1(n7892), .A2(n30210), .ZN(n7796) );
  XOR2_X1 U20600 ( .A1(n23700), .A2(n7832), .Z(n13369) );
  XOR2_X1 U20601 ( .A1(n7833), .A2(n23973), .Z(n7832) );
  NOR2_X2 U20606 ( .A1(n15072), .A2(n14526), .ZN(n7843) );
  XOR2_X1 U20608 ( .A1(n23980), .A2(n21046), .Z(n21045) );
  XOR2_X1 U20609 ( .A1(n7848), .A2(n29021), .Z(n28333) );
  NAND3_X1 U20610 ( .A1(n1438), .A2(n39235), .A3(n9514), .ZN(n14790) );
  NAND2_X2 U20622 ( .A1(n7868), .A2(n7867), .ZN(n20352) );
  XOR2_X1 U20623 ( .A1(n7870), .A2(n10794), .Z(n19308) );
  XOR2_X1 U20624 ( .A1(n9108), .A2(n19929), .Z(n7870) );
  INV_X2 U20625 ( .I(n12686), .ZN(n19420) );
  OR2_X1 U20629 ( .A1(n19731), .A2(n21132), .Z(n22947) );
  XOR2_X1 U20630 ( .A1(n21133), .A2(n22415), .Z(n19731) );
  XOR2_X1 U20635 ( .A1(n8473), .A2(n8939), .Z(n12357) );
  INV_X1 U20644 ( .I(n7914), .ZN(n14713) );
  NAND2_X1 U20646 ( .A1(n7914), .A2(n28625), .ZN(n21004) );
  XOR2_X1 U20648 ( .A1(n11938), .A2(n23696), .Z(n7920) );
  XOR2_X1 U20651 ( .A1(n1618), .A2(n1357), .Z(n7919) );
  XOR2_X1 U20656 ( .A1(n8729), .A2(n35262), .Z(n28987) );
  XOR2_X1 U20658 ( .A1(n29820), .A2(n1050), .Z(n7929) );
  XOR2_X1 U20659 ( .A1(n7931), .A2(n7932), .Z(n13635) );
  XOR2_X1 U20662 ( .A1(n18595), .A2(n22411), .Z(n22447) );
  NAND3_X1 U20664 ( .A1(n34179), .A2(n9918), .A3(n31629), .ZN(n7933) );
  NOR2_X2 U20665 ( .A1(n7591), .A2(n20053), .ZN(n8498) );
  AOI22_X2 U20672 ( .A1(n20037), .A2(n21645), .B1(n21462), .B2(n21910), .ZN(
        n21553) );
  NOR2_X2 U20673 ( .A1(n20037), .A2(n39650), .ZN(n21719) );
  XOR2_X1 U20677 ( .A1(n7980), .A2(n7979), .Z(n26704) );
  NAND2_X2 U20680 ( .A1(n7969), .A2(n7968), .ZN(n25278) );
  XOR2_X1 U20683 ( .A1(n25853), .A2(n747), .Z(n7979) );
  OAI22_X2 U20690 ( .A1(n21439), .A2(n21853), .B1(n21438), .B2(n21687), .ZN(
        n8040) );
  OAI22_X2 U20693 ( .A1(n33978), .A2(n9312), .B1(n9320), .B2(n18801), .ZN(
        n26180) );
  NAND3_X1 U20696 ( .A1(n36183), .A2(n1225), .A3(n27337), .ZN(n18268) );
  NOR2_X2 U20706 ( .A1(n8012), .A2(n8011), .ZN(n23607) );
  XOR2_X1 U20710 ( .A1(n16270), .A2(n14053), .Z(n8015) );
  NAND4_X1 U20715 ( .A1(n8213), .A2(n8211), .A3(n18381), .A4(n18382), .ZN(
        n8023) );
  NOR2_X2 U20718 ( .A1(n21855), .A2(n21856), .ZN(n22243) );
  NAND2_X1 U20720 ( .A1(n6443), .A2(n30153), .ZN(n8030) );
  XOR2_X1 U20722 ( .A1(n22629), .A2(n29602), .Z(n8037) );
  XOR2_X1 U20723 ( .A1(n12267), .A2(n39548), .Z(n8038) );
  NOR2_X1 U20725 ( .A1(n30022), .A2(n8039), .ZN(n30009) );
  INV_X1 U20731 ( .I(n11956), .ZN(n28548) );
  INV_X1 U20732 ( .I(n28735), .ZN(n16206) );
  XOR2_X1 U20739 ( .A1(n19910), .A2(n8059), .Z(n19183) );
  XOR2_X1 U20741 ( .A1(n8060), .A2(n1169), .Z(Ciphertext[98]) );
  XOR2_X1 U20743 ( .A1(n8067), .A2(n8066), .Z(n8065) );
  XOR2_X1 U20744 ( .A1(n36750), .A2(n29051), .Z(n8066) );
  XOR2_X1 U20745 ( .A1(n22620), .A2(n12243), .Z(n8067) );
  OAI21_X2 U20747 ( .A1(n17358), .A2(n20798), .B(n17356), .ZN(n22371) );
  XOR2_X1 U20749 ( .A1(n8075), .A2(n26600), .Z(n8074) );
  NOR2_X1 U20751 ( .A1(n14837), .A2(n33899), .ZN(n8076) );
  NOR2_X1 U20753 ( .A1(n20632), .A2(n8078), .ZN(n10806) );
  XNOR2_X1 U20756 ( .A1(n17276), .A2(n17273), .ZN(n8078) );
  NOR2_X1 U20758 ( .A1(n28486), .A2(n8082), .ZN(n28031) );
  NAND2_X1 U20759 ( .A1(n1066), .A2(n8082), .ZN(n28392) );
  NOR2_X1 U20760 ( .A1(n28483), .A2(n8082), .ZN(n19610) );
  NOR2_X1 U20761 ( .A1(n16559), .A2(n8082), .ZN(n8658) );
  NAND2_X1 U20762 ( .A1(n12343), .A2(n8082), .ZN(n12342) );
  NAND2_X1 U20763 ( .A1(n36573), .A2(n18144), .ZN(n8085) );
  XOR2_X1 U20768 ( .A1(n27712), .A2(n16759), .Z(n8100) );
  AND2_X1 U20771 ( .A1(n24681), .A2(n8109), .Z(n8108) );
  NOR2_X1 U20775 ( .A1(n124), .A2(n20313), .ZN(n11757) );
  XOR2_X1 U20777 ( .A1(n6522), .A2(n21003), .Z(n8119) );
  NOR2_X1 U20778 ( .A1(n24895), .A2(n25583), .ZN(n8123) );
  OAI21_X2 U20782 ( .A1(n8127), .A2(n24877), .B(n8125), .ZN(n21028) );
  INV_X2 U20783 ( .I(n8128), .ZN(n16080) );
  XOR2_X1 U20789 ( .A1(n26476), .A2(n8585), .Z(n8132) );
  XOR2_X1 U20790 ( .A1(n38951), .A2(n19717), .Z(n8136) );
  NAND2_X2 U20795 ( .A1(n13748), .A2(n13747), .ZN(n8139) );
  INV_X2 U20798 ( .I(n8151), .ZN(n22915) );
  XOR2_X1 U20804 ( .A1(n8163), .A2(n19624), .Z(n25260) );
  XOR2_X1 U20805 ( .A1(n8163), .A2(n29238), .Z(n24952) );
  XOR2_X1 U20811 ( .A1(n8171), .A2(n17060), .Z(n23152) );
  XOR2_X1 U20812 ( .A1(n8172), .A2(n13295), .Z(n8171) );
  XOR2_X1 U20813 ( .A1(n8176), .A2(n8180), .Z(n26746) );
  XOR2_X1 U20815 ( .A1(n12839), .A2(n35984), .Z(n8177) );
  XOR2_X1 U20817 ( .A1(n8502), .A2(n9018), .Z(n8180) );
  INV_X2 U20823 ( .I(n8186), .ZN(n14383) );
  XNOR2_X1 U20824 ( .A1(n8187), .A2(n8188), .ZN(n8186) );
  XOR2_X1 U20826 ( .A1(n8189), .A2(n26429), .Z(n8188) );
  NAND2_X1 U20829 ( .A1(n8201), .A2(n8193), .ZN(n8200) );
  OAI21_X2 U20831 ( .A1(n8338), .A2(n8892), .B(n8202), .ZN(n13786) );
  NAND2_X2 U20833 ( .A1(n9251), .A2(n21127), .ZN(n8882) );
  INV_X2 U20834 ( .I(n8205), .ZN(n14478) );
  NOR2_X2 U20835 ( .A1(n8205), .A2(n16081), .ZN(n10815) );
  NAND2_X1 U20836 ( .A1(n7424), .A2(n14949), .ZN(n27035) );
  NOR2_X2 U20839 ( .A1(n27036), .A2(n19034), .ZN(n27570) );
  XOR2_X1 U20840 ( .A1(n31214), .A2(n19877), .Z(n18969) );
  XOR2_X1 U20848 ( .A1(n32448), .A2(n21280), .Z(n14476) );
  XOR2_X1 U20849 ( .A1(n32448), .A2(n33320), .Z(n28857) );
  MUX2_X1 U20851 ( .I0(n8236), .I1(n26077), .S(n11807), .Z(n8235) );
  XOR2_X1 U20854 ( .A1(n8244), .A2(n8242), .Z(n11497) );
  XOR2_X1 U20855 ( .A1(n25081), .A2(n8243), .Z(n8242) );
  XOR2_X1 U20856 ( .A1(n16627), .A2(n1358), .Z(n8243) );
  XOR2_X1 U20857 ( .A1(n25032), .A2(n25314), .Z(n8244) );
  XOR2_X1 U20859 ( .A1(n8247), .A2(n8246), .Z(n12634) );
  XOR2_X1 U20860 ( .A1(n26560), .A2(n30473), .Z(n8246) );
  XOR2_X1 U20861 ( .A1(n26594), .A2(n26305), .Z(n26560) );
  NAND2_X1 U20864 ( .A1(n27560), .A2(n8253), .ZN(n27561) );
  NOR2_X1 U20867 ( .A1(n27456), .A2(n27455), .ZN(n8257) );
  NAND2_X2 U20869 ( .A1(n26638), .A2(n26637), .ZN(n27240) );
  XOR2_X1 U20878 ( .A1(n25080), .A2(n1260), .Z(n8276) );
  XOR2_X1 U20883 ( .A1(n27464), .A2(n27503), .Z(n27650) );
  XOR2_X1 U20884 ( .A1(n27848), .A2(n35189), .Z(n8280) );
  XOR2_X1 U20888 ( .A1(n38190), .A2(n30324), .Z(n8283) );
  NAND2_X1 U20892 ( .A1(n8287), .A2(n20274), .ZN(n20510) );
  INV_X2 U20895 ( .I(n12001), .ZN(n9751) );
  XOR2_X1 U20901 ( .A1(n8299), .A2(n15160), .Z(n8298) );
  XOR2_X1 U20903 ( .A1(n25303), .A2(n25252), .Z(n17804) );
  XOR2_X1 U20906 ( .A1(n8303), .A2(n29978), .Z(n12003) );
  XOR2_X1 U20907 ( .A1(n16096), .A2(n8303), .Z(n17643) );
  XOR2_X1 U20908 ( .A1(n8303), .A2(n30016), .Z(n28607) );
  NOR2_X1 U20909 ( .A1(n8304), .A2(n16080), .ZN(n14515) );
  OAI21_X1 U20910 ( .A1(n34150), .A2(n8305), .B(n15180), .ZN(n25712) );
  XOR2_X1 U20922 ( .A1(n8335), .A2(n8334), .Z(n8333) );
  XOR2_X1 U20923 ( .A1(n27778), .A2(n1704), .Z(n8334) );
  XOR2_X1 U20928 ( .A1(n26495), .A2(n29229), .Z(n8340) );
  NOR2_X1 U20935 ( .A1(n10940), .A2(n15873), .ZN(n24410) );
  NAND2_X1 U20937 ( .A1(n21929), .A2(n917), .ZN(n21060) );
  NAND2_X2 U20938 ( .A1(n20525), .A2(n20522), .ZN(n30245) );
  AOI21_X1 U20950 ( .A1(n5675), .A2(n32191), .B(n33662), .ZN(n8384) );
  AOI21_X1 U20952 ( .A1(n23049), .A2(n8491), .B(n8386), .ZN(n23051) );
  XOR2_X1 U20957 ( .A1(n18633), .A2(n8397), .Z(n8396) );
  XOR2_X1 U20964 ( .A1(n26448), .A2(n7602), .Z(n8409) );
  XOR2_X1 U20965 ( .A1(n26449), .A2(n9152), .Z(n8410) );
  NAND2_X1 U20967 ( .A1(n8412), .A2(n27211), .ZN(n27096) );
  OAI21_X1 U20970 ( .A1(n27438), .A2(n4771), .B(n8412), .ZN(n12916) );
  XOR2_X1 U20975 ( .A1(n31293), .A2(n26519), .Z(n26176) );
  XOR2_X1 U20978 ( .A1(n8425), .A2(n27494), .Z(n8424) );
  NAND2_X1 U20985 ( .A1(n18148), .A2(n8430), .ZN(n11609) );
  NAND3_X1 U20987 ( .A1(n32817), .A2(n20679), .A3(n3676), .ZN(n14904) );
  AOI21_X1 U20988 ( .A1(n1341), .A2(n32817), .B(n3676), .ZN(n9223) );
  NAND2_X1 U20990 ( .A1(n8799), .A2(n31381), .ZN(n8438) );
  NAND3_X1 U20994 ( .A1(n7278), .A2(n17242), .A3(n21898), .ZN(n8441) );
  INV_X2 U20995 ( .I(n8443), .ZN(n30057) );
  NAND2_X1 U21002 ( .A1(n8463), .A2(n24294), .ZN(n24208) );
  AOI21_X2 U21004 ( .A1(n20680), .A2(n20682), .B(n15490), .ZN(n20679) );
  OAI21_X1 U21008 ( .A1(n293), .A2(n8468), .B(n19323), .ZN(n21734) );
  NOR2_X1 U21009 ( .A1(n18926), .A2(n8468), .ZN(n8466) );
  XOR2_X1 U21012 ( .A1(n8474), .A2(n8470), .Z(n8469) );
  XOR2_X1 U21013 ( .A1(n29147), .A2(n19498), .Z(n8470) );
  XOR2_X1 U21014 ( .A1(n8472), .A2(n29148), .Z(n8471) );
  NAND2_X2 U21015 ( .A1(n27914), .A2(n27913), .ZN(n8476) );
  NOR2_X2 U21019 ( .A1(n1245), .A2(n834), .ZN(n18884) );
  XOR2_X1 U21021 ( .A1(n25295), .A2(n8483), .Z(n8482) );
  XOR2_X1 U21022 ( .A1(n19359), .A2(n29509), .Z(n8483) );
  XOR2_X1 U21023 ( .A1(n2145), .A2(n23805), .Z(n8632) );
  XOR2_X1 U21026 ( .A1(n22574), .A2(n22576), .Z(n13550) );
  NAND2_X1 U21031 ( .A1(n19604), .A2(n396), .ZN(n16936) );
  NOR2_X1 U21032 ( .A1(n22313), .A2(n396), .ZN(n15294) );
  NAND2_X1 U21033 ( .A1(n13912), .A2(n396), .ZN(n13911) );
  NOR2_X1 U21036 ( .A1(n21929), .A2(n8495), .ZN(n21059) );
  OAI22_X2 U21037 ( .A1(n14813), .A2(n21928), .B1(n14811), .B2(n8495), .ZN(
        n22337) );
  INV_X1 U21038 ( .I(n21927), .ZN(n8495) );
  XOR2_X1 U21044 ( .A1(n8671), .A2(n13215), .Z(n8505) );
  XOR2_X1 U21050 ( .A1(n8512), .A2(n8511), .Z(n13904) );
  XOR2_X1 U21051 ( .A1(n23918), .A2(n12553), .Z(n8511) );
  XOR2_X1 U21054 ( .A1(n13483), .A2(n8515), .Z(n8514) );
  XOR2_X1 U21055 ( .A1(n18785), .A2(n19835), .Z(n8515) );
  XNOR2_X1 U21058 ( .A1(Plaintext[12]), .A2(Key[12]), .ZN(n8517) );
  XOR2_X1 U21062 ( .A1(n12690), .A2(n8528), .Z(n11870) );
  XOR2_X1 U21063 ( .A1(n19355), .A2(n1702), .Z(n8528) );
  XOR2_X1 U21066 ( .A1(n29823), .A2(n8531), .Z(n8530) );
  XOR2_X1 U21067 ( .A1(n31524), .A2(n30964), .Z(n29823) );
  XOR2_X1 U21070 ( .A1(n29824), .A2(n8532), .Z(n8531) );
  XOR2_X1 U21071 ( .A1(n29822), .A2(n29827), .Z(n8533) );
  XOR2_X1 U21072 ( .A1(n8852), .A2(n28943), .Z(n29822) );
  NAND2_X1 U21073 ( .A1(n8517), .A2(n21898), .ZN(n20898) );
  INV_X2 U21074 ( .I(n14217), .ZN(n14426) );
  XOR2_X1 U21075 ( .A1(n27619), .A2(n27618), .Z(n8540) );
  XOR2_X1 U21077 ( .A1(n30761), .A2(n32218), .Z(n16843) );
  XOR2_X1 U21078 ( .A1(n25149), .A2(n30761), .Z(n24953) );
  XOR2_X1 U21080 ( .A1(n30761), .A2(n25014), .Z(n24631) );
  NOR2_X1 U21081 ( .A1(n29951), .A2(n29997), .ZN(n19197) );
  XOR2_X1 U21087 ( .A1(n10579), .A2(n27467), .Z(n8553) );
  XOR2_X1 U21091 ( .A1(n1503), .A2(n16735), .Z(n8559) );
  INV_X1 U21092 ( .I(Plaintext[116]), .ZN(n8562) );
  XOR2_X1 U21093 ( .A1(n8562), .A2(Key[116]), .Z(n9308) );
  XOR2_X1 U21095 ( .A1(n8566), .A2(n18482), .Z(n8565) );
  XOR2_X1 U21096 ( .A1(n10526), .A2(n23931), .Z(n18482) );
  XOR2_X1 U21097 ( .A1(n24043), .A2(n23763), .Z(n8567) );
  OR2_X1 U21098 ( .A1(n21969), .A2(n34015), .Z(n8570) );
  AOI21_X1 U21104 ( .A1(n16187), .A2(n8584), .B(n8582), .ZN(n19138) );
  AOI21_X1 U21105 ( .A1(n31570), .A2(n9591), .B(n1174), .ZN(n8584) );
  NAND3_X1 U21110 ( .A1(n8731), .A2(n33256), .A3(n16224), .ZN(n8590) );
  NAND2_X1 U21111 ( .A1(n30049), .A2(n29936), .ZN(n8593) );
  XOR2_X1 U21120 ( .A1(n26432), .A2(n26517), .Z(n8625) );
  XOR2_X1 U21122 ( .A1(n26431), .A2(n14148), .Z(n8626) );
  XOR2_X1 U21127 ( .A1(n8632), .A2(n23806), .Z(n8631) );
  INV_X2 U21128 ( .I(n8824), .ZN(n13453) );
  XNOR2_X1 U21132 ( .A1(Plaintext[15]), .A2(Key[15]), .ZN(n8653) );
  NAND2_X1 U21136 ( .A1(n29901), .A2(n13607), .ZN(n8666) );
  OR2_X1 U21146 ( .A1(n23078), .A2(n20873), .Z(n8674) );
  OAI21_X2 U21149 ( .A1(n21143), .A2(n23076), .B(n23078), .ZN(n14804) );
  XOR2_X1 U21150 ( .A1(n8678), .A2(n15808), .Z(n14403) );
  NAND2_X1 U21154 ( .A1(n22243), .A2(n37089), .ZN(n8754) );
  NOR2_X1 U21155 ( .A1(n37089), .A2(n21864), .ZN(n8688) );
  XOR2_X1 U21162 ( .A1(Plaintext[164]), .A2(Key[164]), .Z(n21938) );
  NOR3_X1 U21163 ( .A1(n22349), .A2(n14423), .A3(n7955), .ZN(n8701) );
  INV_X2 U21165 ( .I(n10733), .ZN(n13584) );
  NAND3_X1 U21174 ( .A1(n1477), .A2(n27412), .A3(n34969), .ZN(n27159) );
  XOR2_X1 U21180 ( .A1(n13374), .A2(n38962), .Z(n8723) );
  NAND2_X1 U21186 ( .A1(n14933), .A2(n8728), .ZN(n14199) );
  AOI21_X1 U21187 ( .A1(n16837), .A2(n16839), .B(n8728), .ZN(n16838) );
  XOR2_X1 U21191 ( .A1(n29829), .A2(n29832), .Z(n8732) );
  INV_X2 U21192 ( .I(n8736), .ZN(n21436) );
  XNOR2_X1 U21193 ( .A1(Plaintext[33]), .A2(Key[33]), .ZN(n8736) );
  NAND2_X1 U21195 ( .A1(n955), .A2(n8738), .ZN(n8737) );
  XOR2_X1 U21205 ( .A1(n27502), .A2(n8748), .Z(n8747) );
  XOR2_X1 U21206 ( .A1(n29292), .A2(n29291), .Z(n8755) );
  XOR2_X1 U21211 ( .A1(n38154), .A2(n1938), .Z(n11153) );
  NAND2_X1 U21213 ( .A1(n8762), .A2(n29704), .ZN(n20436) );
  NAND2_X1 U21214 ( .A1(n28843), .A2(n29635), .ZN(n20474) );
  XOR2_X1 U21216 ( .A1(n28838), .A2(n8774), .Z(n8773) );
  XOR2_X1 U21217 ( .A1(n28920), .A2(n8776), .Z(n8775) );
  XOR2_X1 U21219 ( .A1(n28977), .A2(n10079), .Z(n8776) );
  XOR2_X1 U21224 ( .A1(n27662), .A2(n19953), .Z(n8782) );
  OAI21_X1 U21226 ( .A1(n22165), .A2(n8792), .B(n22221), .ZN(n18804) );
  XOR2_X1 U21227 ( .A1(n37899), .A2(n35215), .Z(n23975) );
  XOR2_X1 U21229 ( .A1(n27665), .A2(n8794), .Z(n8793) );
  XOR2_X1 U21230 ( .A1(n13569), .A2(n1699), .Z(n8794) );
  XOR2_X1 U21232 ( .A1(n25215), .A2(n19800), .Z(n8796) );
  NAND2_X1 U21236 ( .A1(n8799), .A2(n21898), .ZN(n17847) );
  XNOR2_X1 U21237 ( .A1(n27540), .A2(n9013), .ZN(n14986) );
  NOR2_X2 U21238 ( .A1(n11463), .A2(n11462), .ZN(n27540) );
  INV_X2 U21242 ( .I(n8812), .ZN(n22368) );
  INV_X2 U21249 ( .I(n12634), .ZN(n12755) );
  XOR2_X1 U21251 ( .A1(n23802), .A2(n23803), .Z(n8826) );
  NAND3_X1 U21261 ( .A1(n15121), .A2(n9380), .A3(n34577), .ZN(n25378) );
  NAND2_X1 U21276 ( .A1(n8882), .A2(n22131), .ZN(n21968) );
  AOI21_X1 U21277 ( .A1(n36457), .A2(n31573), .B(n35780), .ZN(n14323) );
  XOR2_X1 U21278 ( .A1(n38041), .A2(n29051), .Z(n8885) );
  XOR2_X1 U21281 ( .A1(n29260), .A2(n31591), .Z(n8887) );
  INV_X2 U21283 ( .I(n8889), .ZN(n10436) );
  XOR2_X1 U21284 ( .A1(n4819), .A2(n1713), .Z(n8890) );
  INV_X1 U21285 ( .I(Plaintext[97]), .ZN(n8891) );
  XOR2_X1 U21286 ( .A1(n8891), .A2(Key[97]), .Z(n9552) );
  XOR2_X1 U21296 ( .A1(n8902), .A2(n8901), .Z(n8900) );
  XOR2_X1 U21297 ( .A1(n35239), .A2(n1370), .Z(n8901) );
  NAND2_X1 U21300 ( .A1(n32419), .A2(n833), .ZN(n8906) );
  INV_X2 U21306 ( .I(n14170), .ZN(n14415) );
  AND2_X1 U21314 ( .A1(n5282), .A2(n1270), .Z(n24516) );
  XOR2_X1 U21316 ( .A1(n23590), .A2(n29223), .Z(n8929) );
  XOR2_X1 U21319 ( .A1(n8939), .A2(n29206), .Z(n28887) );
  AND2_X1 U21320 ( .A1(n9745), .A2(n28508), .Z(n8934) );
  NOR2_X1 U21322 ( .A1(n1158), .A2(n8936), .ZN(n20681) );
  XNOR2_X1 U21323 ( .A1(Plaintext[31]), .A2(Key[31]), .ZN(n8936) );
  XOR2_X1 U21324 ( .A1(n19991), .A2(n8938), .Z(n8937) );
  XOR2_X1 U21327 ( .A1(n23831), .A2(n19729), .Z(n8938) );
  XOR2_X1 U21330 ( .A1(n8940), .A2(n1167), .Z(n13497) );
  AOI21_X1 U21332 ( .A1(n22221), .A2(n22219), .B(n9387), .ZN(n8949) );
  XOR2_X1 U21335 ( .A1(n26489), .A2(n8951), .Z(n8950) );
  XOR2_X1 U21336 ( .A1(n10621), .A2(n19835), .Z(n8952) );
  XOR2_X1 U21339 ( .A1(n37129), .A2(n28868), .Z(n8957) );
  INV_X2 U21341 ( .I(n16907), .ZN(n29059) );
  XOR2_X1 U21344 ( .A1(Plaintext[79]), .A2(Key[79]), .Z(n17209) );
  NOR2_X1 U21345 ( .A1(n8970), .A2(n7536), .ZN(n8969) );
  XOR2_X1 U21348 ( .A1(n33083), .A2(n1010), .Z(n26468) );
  XOR2_X1 U21352 ( .A1(n27729), .A2(n17884), .Z(n8974) );
  XOR2_X1 U21357 ( .A1(n38208), .A2(n19801), .Z(n8982) );
  INV_X2 U21359 ( .I(n8983), .ZN(n25696) );
  XOR2_X1 U21360 ( .A1(n15361), .A2(n17255), .Z(n8983) );
  XOR2_X1 U21362 ( .A1(n24071), .A2(n8985), .Z(n12912) );
  XOR2_X1 U21363 ( .A1(n15916), .A2(n8986), .Z(n8985) );
  NAND3_X1 U21364 ( .A1(n34379), .A2(n7916), .A3(n38246), .ZN(n22032) );
  XOR2_X1 U21368 ( .A1(n23852), .A2(n23853), .Z(n9003) );
  XOR2_X1 U21373 ( .A1(n25280), .A2(n1371), .Z(n9005) );
  XOR2_X1 U21376 ( .A1(n9010), .A2(n9009), .Z(n19840) );
  XOR2_X1 U21377 ( .A1(n22650), .A2(n22649), .Z(n9009) );
  XOR2_X1 U21378 ( .A1(n10384), .A2(n14194), .Z(n9010) );
  XOR2_X1 U21381 ( .A1(n26396), .A2(n26460), .Z(n9018) );
  AOI22_X2 U21383 ( .A1(n15554), .A2(n9021), .B1(n18744), .B2(n15553), .ZN(
        n25160) );
  NAND2_X2 U21384 ( .A1(n16999), .A2(n37067), .ZN(n9021) );
  XOR2_X1 U21385 ( .A1(n9023), .A2(n9022), .Z(n14709) );
  NOR2_X2 U21391 ( .A1(n16230), .A2(n16229), .ZN(n18142) );
  XOR2_X1 U21393 ( .A1(n9013), .A2(n1733), .Z(n9027) );
  XOR2_X1 U21394 ( .A1(n15653), .A2(n22441), .Z(n9028) );
  XOR2_X1 U21397 ( .A1(n9030), .A2(n35251), .Z(n26293) );
  OR2_X1 U21398 ( .A1(n24607), .A2(n29285), .Z(n9032) );
  XOR2_X1 U21399 ( .A1(n24610), .A2(n9033), .Z(n13938) );
  AOI21_X1 U21402 ( .A1(n29613), .A2(n29612), .B(n9044), .ZN(n29615) );
  OAI21_X2 U21403 ( .A1(n9049), .A2(n21289), .B(n9047), .ZN(n29859) );
  XOR2_X1 U21404 ( .A1(n9054), .A2(n11347), .Z(n11349) );
  NOR2_X1 U21406 ( .A1(n9062), .A2(n15411), .ZN(n9058) );
  AOI21_X1 U21407 ( .A1(n9061), .A2(n9060), .B(n11226), .ZN(n9059) );
  INV_X2 U21414 ( .I(n16160), .ZN(n26619) );
  XOR2_X1 U21417 ( .A1(n17519), .A2(n17516), .Z(n16179) );
  XOR2_X1 U21421 ( .A1(n9246), .A2(n15916), .Z(n9247) );
  XOR2_X1 U21422 ( .A1(n9093), .A2(n9092), .Z(n9091) );
  XOR2_X1 U21423 ( .A1(n22483), .A2(n29238), .Z(n9092) );
  XOR2_X1 U21424 ( .A1(n13596), .A2(n9095), .Z(n9094) );
  XOR2_X1 U21425 ( .A1(n25243), .A2(n19592), .Z(n9095) );
  XOR2_X1 U21431 ( .A1(n9114), .A2(n1713), .Z(n10485) );
  XOR2_X1 U21432 ( .A1(n9114), .A2(n17428), .Z(n19824) );
  XOR2_X1 U21433 ( .A1(n25093), .A2(n9113), .Z(n25095) );
  XOR2_X1 U21434 ( .A1(n9114), .A2(n25192), .Z(n17555) );
  XOR2_X1 U21435 ( .A1(n26454), .A2(n26453), .Z(n9119) );
  XOR2_X1 U21436 ( .A1(n26259), .A2(n26402), .Z(n26453) );
  XOR2_X1 U21438 ( .A1(n26456), .A2(n32528), .Z(n9120) );
  XOR2_X1 U21446 ( .A1(n17140), .A2(n655), .Z(n9123) );
  NAND2_X1 U21449 ( .A1(n1331), .A2(n18656), .ZN(n14590) );
  NOR2_X1 U21450 ( .A1(n22229), .A2(n9129), .ZN(n22088) );
  AOI21_X2 U21454 ( .A1(n1024), .A2(n25637), .B(n14410), .ZN(n12866) );
  XOR2_X1 U21459 ( .A1(n27657), .A2(n27463), .Z(n9139) );
  AOI21_X1 U21462 ( .A1(n24795), .A2(n9149), .B(n24646), .ZN(n9148) );
  NOR2_X1 U21464 ( .A1(n3944), .A2(n14448), .ZN(n28468) );
  XOR2_X1 U21468 ( .A1(n26532), .A2(n19407), .Z(n9152) );
  XOR2_X1 U21469 ( .A1(n39163), .A2(n19738), .Z(n9153) );
  AND2_X1 U21470 ( .A1(n26927), .A2(n735), .Z(n9156) );
  XOR2_X1 U21472 ( .A1(n9160), .A2(n16161), .Z(n9159) );
  NAND2_X2 U21477 ( .A1(n18769), .A2(n18767), .ZN(n27730) );
  XOR2_X1 U21484 ( .A1(n7475), .A2(n28821), .Z(n9244) );
  INV_X1 U21486 ( .I(Plaintext[39]), .ZN(n9180) );
  XOR2_X1 U21487 ( .A1(n9180), .A2(Key[39]), .Z(n20361) );
  NOR2_X1 U21488 ( .A1(n15663), .A2(n1342), .ZN(n21451) );
  AOI21_X1 U21489 ( .A1(n1341), .A2(n1342), .B(n32817), .ZN(n13411) );
  INV_X2 U21495 ( .I(n14440), .ZN(n9188) );
  XOR2_X1 U21499 ( .A1(n33587), .A2(n30203), .Z(n9195) );
  XOR2_X1 U21502 ( .A1(n22637), .A2(n32218), .Z(n9206) );
  XOR2_X1 U21503 ( .A1(n12015), .A2(n16226), .Z(n9207) );
  AOI21_X2 U21508 ( .A1(n23909), .A2(n9909), .B(n23908), .ZN(n9218) );
  XOR2_X1 U21512 ( .A1(n23920), .A2(n9220), .Z(n9219) );
  XOR2_X1 U21513 ( .A1(n23890), .A2(n1162), .Z(n9220) );
  NAND2_X1 U21515 ( .A1(n18567), .A2(n14833), .ZN(n9224) );
  XOR2_X1 U21517 ( .A1(n38165), .A2(n17428), .Z(n9230) );
  INV_X2 U21519 ( .I(n9235), .ZN(n19821) );
  XOR2_X1 U21524 ( .A1(n9247), .A2(n9244), .Z(n9243) );
  XOR2_X1 U21534 ( .A1(n33197), .A2(n29657), .Z(n9272) );
  XOR2_X1 U21535 ( .A1(n22429), .A2(n22762), .Z(n19342) );
  XOR2_X1 U21536 ( .A1(n21149), .A2(n9275), .Z(n9274) );
  XOR2_X1 U21537 ( .A1(n27549), .A2(n1724), .Z(n9275) );
  NAND2_X1 U21538 ( .A1(n10589), .A2(n34786), .ZN(n9278) );
  AND2_X1 U21546 ( .A1(n31669), .A2(n25696), .Z(n9292) );
  AOI21_X1 U21547 ( .A1(n11734), .A2(n36666), .B(n1103), .ZN(n9294) );
  XOR2_X1 U21548 ( .A1(n29021), .A2(n12707), .Z(n11077) );
  XOR2_X1 U21549 ( .A1(n12707), .A2(n31515), .Z(n28406) );
  XOR2_X1 U21550 ( .A1(n9299), .A2(n9298), .Z(n9297) );
  XOR2_X1 U21551 ( .A1(n26519), .A2(n1714), .Z(n9298) );
  XOR2_X1 U21552 ( .A1(n26516), .A2(n26518), .Z(n9299) );
  INV_X2 U21559 ( .I(n9308), .ZN(n14493) );
  XOR2_X1 U21560 ( .A1(n25193), .A2(n29805), .Z(n9309) );
  AOI21_X1 U21562 ( .A1(n1511), .A2(n31133), .B(n37378), .ZN(n9312) );
  NAND2_X2 U21565 ( .A1(n10580), .A2(n26942), .ZN(n9315) );
  NOR2_X2 U21567 ( .A1(n12122), .A2(n12121), .ZN(n9920) );
  NAND2_X1 U21570 ( .A1(n9326), .A2(n4602), .ZN(n25891) );
  OAI21_X2 U21574 ( .A1(n25644), .A2(n25361), .B(n9337), .ZN(n11589) );
  INV_X2 U21575 ( .I(n10686), .ZN(n25644) );
  INV_X2 U21576 ( .I(n9338), .ZN(n25699) );
  INV_X1 U21577 ( .I(n9698), .ZN(n9340) );
  NAND3_X1 U21582 ( .A1(n33987), .A2(n24709), .A3(n6273), .ZN(n9357) );
  NAND2_X1 U21586 ( .A1(n32891), .A2(n9371), .ZN(n23799) );
  AOI21_X1 U21587 ( .A1(n39605), .A2(n31452), .B(n9371), .ZN(n9821) );
  INV_X2 U21588 ( .I(n24280), .ZN(n9371) );
  INV_X2 U21590 ( .I(n9373), .ZN(n14389) );
  INV_X2 U21591 ( .I(n9374), .ZN(n18144) );
  XOR2_X1 U21594 ( .A1(n38149), .A2(n26567), .Z(n20139) );
  XOR2_X1 U21599 ( .A1(n9390), .A2(n24929), .Z(n19742) );
  NAND2_X1 U21600 ( .A1(n5669), .A2(n21299), .ZN(n16171) );
  NAND3_X1 U21601 ( .A1(n5414), .A2(n30238), .A3(n5669), .ZN(n12232) );
  XOR2_X1 U21603 ( .A1(n26481), .A2(n29221), .Z(n9398) );
  XOR2_X1 U21609 ( .A1(n26386), .A2(n26474), .Z(n9408) );
  XOR2_X1 U21612 ( .A1(n9411), .A2(n9410), .Z(n9409) );
  XOR2_X1 U21613 ( .A1(n26390), .A2(n29978), .Z(n9410) );
  XOR2_X1 U21614 ( .A1(n9776), .A2(n37024), .Z(n9411) );
  XOR2_X1 U21615 ( .A1(n25201), .A2(n11899), .Z(n9550) );
  NOR2_X2 U21617 ( .A1(n19740), .A2(n9413), .ZN(n25996) );
  MUX2_X1 U21618 ( .I0(n24763), .I1(n9417), .S(n24691), .Z(n9416) );
  XOR2_X1 U21623 ( .A1(n18857), .A2(n9431), .Z(n9430) );
  XOR2_X1 U21624 ( .A1(n23885), .A2(n34672), .Z(n9431) );
  XOR2_X1 U21630 ( .A1(n22755), .A2(n19145), .Z(n9448) );
  NAND3_X1 U21631 ( .A1(n32050), .A2(n29794), .A3(n15867), .ZN(n9457) );
  NOR2_X1 U21635 ( .A1(n16663), .A2(n26932), .ZN(n17394) );
  NOR2_X1 U21636 ( .A1(n26933), .A2(n26932), .ZN(n17392) );
  XOR2_X1 U21637 ( .A1(n14902), .A2(n15171), .Z(n9469) );
  XOR2_X1 U21638 ( .A1(n22669), .A2(n22556), .Z(n9468) );
  XOR2_X1 U21643 ( .A1(n22503), .A2(n7432), .Z(n9496) );
  XOR2_X1 U21644 ( .A1(n22744), .A2(n35211), .Z(n22616) );
  OAI21_X1 U21648 ( .A1(n1654), .A2(n18708), .B(n9507), .ZN(n9506) );
  INV_X2 U21649 ( .I(n9509), .ZN(n22802) );
  NAND2_X2 U21652 ( .A1(n9513), .A2(n27121), .ZN(n27776) );
  INV_X2 U21655 ( .I(n14306), .ZN(n9520) );
  INV_X1 U21657 ( .I(n9529), .ZN(n12624) );
  NAND2_X1 U21668 ( .A1(n9546), .A2(n7916), .ZN(n21816) );
  NAND3_X1 U21669 ( .A1(n16888), .A2(n13632), .A3(n9546), .ZN(n21815) );
  XOR2_X1 U21671 ( .A1(n23922), .A2(n23901), .Z(n9549) );
  XOR2_X1 U21672 ( .A1(n9550), .A2(n17878), .Z(n20614) );
  INV_X2 U21673 ( .I(n9552), .ZN(n21869) );
  XOR2_X1 U21675 ( .A1(n3413), .A2(n15046), .Z(n9554) );
  NOR2_X2 U21682 ( .A1(n12371), .A2(n12372), .ZN(n16889) );
  OAI21_X1 U21685 ( .A1(n9321), .A2(n14477), .B(n33840), .ZN(n17875) );
  XOR2_X1 U21686 ( .A1(n9565), .A2(n9564), .Z(n9563) );
  XOR2_X1 U21687 ( .A1(n12233), .A2(n39559), .Z(n9565) );
  OAI22_X2 U21691 ( .A1(n20180), .A2(n14827), .B1(n24729), .B2(n1273), .ZN(
        n24922) );
  NAND2_X1 U21695 ( .A1(n28380), .A2(n7555), .ZN(n28099) );
  XOR2_X1 U21699 ( .A1(n19973), .A2(n26282), .Z(n12735) );
  OR2_X1 U21703 ( .A1(n12471), .A2(n39811), .Z(n15151) );
  NOR2_X1 U21705 ( .A1(n26813), .A2(n11138), .ZN(n15352) );
  NAND3_X1 U21706 ( .A1(n17308), .A2(n33782), .A3(n21458), .ZN(n11672) );
  NAND2_X1 U21713 ( .A1(n30156), .A2(n16786), .ZN(n10210) );
  AND2_X1 U21715 ( .A1(n26724), .A2(n14318), .Z(n18225) );
  NOR2_X1 U21716 ( .A1(n33230), .A2(n24759), .ZN(n13903) );
  OR2_X1 U21719 ( .A1(n33368), .A2(n14428), .Z(n13723) );
  AND2_X1 U21724 ( .A1(n19609), .A2(n455), .Z(n21343) );
  INV_X2 U21726 ( .I(n9604), .ZN(n13285) );
  XOR2_X1 U21727 ( .A1(Plaintext[143]), .A2(Key[143]), .Z(n9604) );
  NAND2_X1 U21730 ( .A1(n39140), .A2(n38198), .ZN(n9605) );
  AOI21_X1 U21732 ( .A1(n12978), .A2(n29218), .B(n1378), .ZN(n9607) );
  INV_X4 U21733 ( .I(n11304), .ZN(n12077) );
  XNOR2_X1 U21734 ( .A1(n28970), .A2(n20137), .ZN(n9853) );
  NAND2_X1 U21735 ( .A1(n22684), .A2(n37589), .ZN(n9608) );
  NAND2_X2 U21736 ( .A1(n21061), .A2(n21064), .ZN(n23639) );
  NAND2_X1 U21741 ( .A1(n14497), .A2(n28468), .ZN(n28471) );
  XOR2_X1 U21743 ( .A1(n25268), .A2(n814), .Z(n9624) );
  OAI21_X1 U21750 ( .A1(n32697), .A2(n9633), .B(n9632), .ZN(n27116) );
  NOR2_X2 U21752 ( .A1(n27045), .A2(n27044), .ZN(n27253) );
  OR2_X1 U21753 ( .A1(n13300), .A2(n24683), .Z(n14657) );
  INV_X1 U21754 ( .I(n29531), .ZN(n29516) );
  XOR2_X1 U21756 ( .A1(n18612), .A2(n35561), .Z(n9643) );
  AND2_X1 U21758 ( .A1(n19085), .A2(n38142), .Z(n18611) );
  NAND2_X1 U21763 ( .A1(n9917), .A2(n28622), .ZN(n20952) );
  AND2_X1 U21774 ( .A1(n28576), .A2(n35199), .Z(n28177) );
  XOR2_X1 U21783 ( .A1(n25196), .A2(n19670), .Z(n24958) );
  NOR2_X1 U21789 ( .A1(n15256), .A2(n24359), .ZN(n10439) );
  AND3_X1 U21790 ( .A1(n16154), .A2(n28141), .A3(n281), .Z(n15975) );
  XOR2_X1 U21791 ( .A1(n22713), .A2(n22195), .Z(n22203) );
  XOR2_X1 U21800 ( .A1(n39636), .A2(n23841), .Z(n16697) );
  NAND2_X2 U21803 ( .A1(n10349), .A2(n11705), .ZN(n28313) );
  XOR2_X1 U21809 ( .A1(n11810), .A2(n11809), .Z(n9687) );
  XOR2_X1 U21810 ( .A1(n26597), .A2(n19627), .Z(n19772) );
  INV_X1 U21831 ( .I(n6523), .ZN(n10904) );
  XOR2_X1 U21837 ( .A1(n12157), .A2(n28100), .Z(n9712) );
  NOR2_X2 U21839 ( .A1(n10174), .A2(n23582), .ZN(n23508) );
  XOR2_X1 U21845 ( .A1(n10113), .A2(n20279), .Z(n20891) );
  NAND2_X1 U21846 ( .A1(n16854), .A2(n16855), .ZN(n12385) );
  XOR2_X1 U21848 ( .A1(n20454), .A2(n29887), .Z(n19766) );
  NAND2_X2 U21849 ( .A1(n948), .A2(n26660), .ZN(n27141) );
  AND2_X1 U21852 ( .A1(n12032), .A2(n7575), .Z(n13157) );
  XOR2_X1 U21857 ( .A1(n9732), .A2(n27536), .Z(n12104) );
  INV_X2 U21862 ( .I(n9737), .ZN(n13998) );
  XOR2_X1 U21863 ( .A1(Plaintext[179]), .A2(Key[179]), .Z(n9737) );
  OR2_X1 U21865 ( .A1(n32105), .A2(n25349), .Z(n12923) );
  INV_X1 U21873 ( .I(n10012), .ZN(n24678) );
  INV_X1 U21875 ( .I(n10847), .ZN(n10846) );
  XOR2_X1 U21887 ( .A1(n36039), .A2(n721), .Z(n12000) );
  XOR2_X1 U21903 ( .A1(n9766), .A2(n25226), .Z(n13575) );
  XOR2_X1 U21904 ( .A1(n25323), .A2(n25006), .Z(n9766) );
  NOR2_X1 U21909 ( .A1(n15420), .A2(n14869), .ZN(n15419) );
  INV_X1 U21910 ( .I(n13219), .ZN(n10754) );
  INV_X2 U21917 ( .I(n9780), .ZN(n16836) );
  NOR2_X1 U21923 ( .A1(n21071), .A2(n21069), .ZN(n29539) );
  INV_X2 U21932 ( .I(n19313), .ZN(n20476) );
  NAND2_X1 U21934 ( .A1(n15003), .A2(n26092), .ZN(n25883) );
  INV_X2 U21938 ( .I(n9813), .ZN(n10334) );
  XOR2_X1 U21939 ( .A1(n22233), .A2(n22232), .Z(n9813) );
  XOR2_X1 U21941 ( .A1(n17987), .A2(n12806), .Z(n12805) );
  XOR2_X1 U21942 ( .A1(n13155), .A2(n29337), .Z(n13154) );
  XOR2_X1 U21951 ( .A1(Plaintext[4]), .A2(Key[4]), .Z(n12225) );
  OAI22_X1 U21954 ( .A1(n7876), .A2(n7284), .B1(n19637), .B2(n1256), .ZN(
        n25352) );
  XOR2_X1 U21957 ( .A1(n9829), .A2(n10027), .Z(Ciphertext[150]) );
  OAI22_X1 U21958 ( .A1(n30084), .A2(n30093), .B1(n30086), .B2(n30083), .ZN(
        n9829) );
  AND2_X1 U21962 ( .A1(n1548), .A2(n10882), .Z(n14625) );
  NOR2_X2 U21964 ( .A1(n16078), .A2(n16076), .ZN(n24925) );
  XOR2_X1 U21969 ( .A1(n18447), .A2(n18449), .Z(n9845) );
  NOR2_X1 U21973 ( .A1(n13646), .A2(n29359), .ZN(n9857) );
  OAI21_X2 U21975 ( .A1(n22634), .A2(n12243), .B(n12242), .ZN(n18751) );
  AND3_X1 U21977 ( .A1(n914), .A2(n14558), .A3(n20313), .Z(n11758) );
  XOR2_X1 U21979 ( .A1(n9852), .A2(n14867), .Z(n14866) );
  XOR2_X1 U21980 ( .A1(n37024), .A2(n36171), .Z(n9852) );
  XNOR2_X1 U21984 ( .A1(n22717), .A2(n37094), .ZN(n14109) );
  INV_X2 U21988 ( .I(n15621), .ZN(n29452) );
  XOR2_X1 U21989 ( .A1(n20135), .A2(n9853), .Z(n15621) );
  XOR2_X1 U21990 ( .A1(n12300), .A2(n26400), .Z(n20098) );
  XOR2_X1 U21992 ( .A1(n15011), .A2(n25100), .Z(n14859) );
  XOR2_X1 U21996 ( .A1(n9857), .A2(n29360), .Z(Ciphertext[31]) );
  OAI22_X1 U22001 ( .A1(n9865), .A2(n14417), .B1(n29596), .B2(n31667), .ZN(
        n28585) );
  NOR2_X2 U22004 ( .A1(n13000), .A2(n9869), .ZN(n12726) );
  NOR2_X2 U22008 ( .A1(n21401), .A2(n21645), .ZN(n9886) );
  NAND2_X2 U22012 ( .A1(n3293), .A2(n21895), .ZN(n21582) );
  XOR2_X1 U22018 ( .A1(n14986), .A2(n754), .Z(n27827) );
  XOR2_X1 U22020 ( .A1(n29002), .A2(n20324), .Z(n20323) );
  XOR2_X1 U22024 ( .A1(n35227), .A2(n16613), .Z(n9887) );
  XOR2_X1 U22026 ( .A1(n26259), .A2(n29711), .Z(n16427) );
  NAND2_X2 U22027 ( .A1(n9891), .A2(n10535), .ZN(n27407) );
  INV_X2 U22028 ( .I(n9895), .ZN(n14636) );
  XOR2_X1 U22029 ( .A1(n16425), .A2(n16423), .Z(n9895) );
  XOR2_X1 U22031 ( .A1(Plaintext[73]), .A2(Key[73]), .Z(n20778) );
  XNOR2_X1 U22037 ( .A1(n22450), .A2(n22451), .ZN(n13667) );
  XOR2_X1 U22039 ( .A1(n10225), .A2(n1356), .Z(n11902) );
  NAND2_X1 U22041 ( .A1(n13107), .A2(n10803), .ZN(n9907) );
  NOR2_X1 U22044 ( .A1(n19310), .A2(n29262), .ZN(n19475) );
  XOR2_X1 U22045 ( .A1(n11437), .A2(n22522), .Z(n9911) );
  AND2_X1 U22048 ( .A1(n18451), .A2(n14451), .Z(n14484) );
  AND2_X1 U22049 ( .A1(n27150), .A2(n20740), .Z(n26966) );
  XOR2_X1 U22059 ( .A1(n25245), .A2(n25187), .Z(n10928) );
  XOR2_X1 U22065 ( .A1(n35532), .A2(n37094), .Z(n9937) );
  NAND2_X1 U22067 ( .A1(n20997), .A2(n31586), .ZN(n9988) );
  AND2_X1 U22068 ( .A1(n13370), .A2(n32377), .Z(n23583) );
  XNOR2_X1 U22069 ( .A1(Key[18]), .A2(Plaintext[18]), .ZN(n9942) );
  NAND2_X1 U22071 ( .A1(n17965), .A2(n13257), .ZN(n15803) );
  XOR2_X1 U22072 ( .A1(n1412), .A2(n38150), .Z(n18493) );
  OAI22_X1 U22074 ( .A1(n21507), .A2(n21509), .B1(n21484), .B2(n21593), .ZN(
        n21485) );
  XOR2_X1 U22080 ( .A1(n736), .A2(n11989), .Z(n9948) );
  XOR2_X1 U22088 ( .A1(n15581), .A2(n15181), .Z(n9952) );
  XOR2_X1 U22089 ( .A1(n9953), .A2(n29887), .Z(Ciphertext[124]) );
  NOR2_X1 U22093 ( .A1(n34049), .A2(n21626), .ZN(n21627) );
  NAND3_X1 U22095 ( .A1(n29621), .A2(n29622), .A3(n29627), .ZN(n9957) );
  NOR2_X2 U22100 ( .A1(n10041), .A2(n11544), .ZN(n9959) );
  XOR2_X1 U22102 ( .A1(n9960), .A2(n20824), .Z(n11856) );
  XOR2_X1 U22108 ( .A1(n9967), .A2(n29109), .Z(Ciphertext[0]) );
  OAI21_X1 U22109 ( .A1(n10681), .A2(n1681), .B(n6361), .ZN(n10979) );
  XOR2_X1 U22110 ( .A1(n14638), .A2(n29245), .Z(n14136) );
  XOR2_X1 U22113 ( .A1(Plaintext[14]), .A2(Key[14]), .Z(n10925) );
  INV_X2 U22115 ( .I(n9973), .ZN(n14422) );
  XOR2_X1 U22116 ( .A1(n19443), .A2(n750), .Z(n18973) );
  XOR2_X1 U22121 ( .A1(n37044), .A2(n14651), .Z(n9976) );
  XOR2_X1 U22124 ( .A1(n1555), .A2(n15625), .Z(n9977) );
  XOR2_X1 U22125 ( .A1(n12282), .A2(n22501), .Z(n9980) );
  XOR2_X1 U22133 ( .A1(n9986), .A2(n823), .Z(n11046) );
  NAND2_X1 U22136 ( .A1(n9991), .A2(n9990), .ZN(n28264) );
  INV_X1 U22137 ( .I(n9992), .ZN(n9991) );
  AOI21_X1 U22138 ( .A1(n28048), .A2(n28255), .B(n28258), .ZN(n9992) );
  BUF_X2 U22140 ( .I(n29493), .Z(n9993) );
  XOR2_X1 U22141 ( .A1(n33322), .A2(n7917), .Z(n23848) );
  XNOR2_X1 U22143 ( .A1(n35245), .A2(n25274), .ZN(n10644) );
  XOR2_X1 U22145 ( .A1(n1259), .A2(n10791), .Z(n24914) );
  NAND3_X2 U22149 ( .A1(n14903), .A2(n5795), .A3(n14904), .ZN(n16798) );
  XOR2_X1 U22154 ( .A1(n19002), .A2(n10001), .Z(n19001) );
  XOR2_X1 U22155 ( .A1(n18751), .A2(n658), .Z(n10001) );
  XNOR2_X1 U22158 ( .A1(n26343), .A2(n19099), .ZN(n10230) );
  AND2_X1 U22167 ( .A1(n19941), .A2(n36794), .Z(n17304) );
  XOR2_X1 U22170 ( .A1(n10583), .A2(n10585), .Z(n10584) );
  XOR2_X1 U22171 ( .A1(n23688), .A2(n23849), .Z(n10014) );
  NAND2_X1 U22172 ( .A1(n16567), .A2(n13851), .ZN(n13600) );
  XOR2_X1 U22174 ( .A1(n11620), .A2(n11621), .Z(n19423) );
  XOR2_X1 U22175 ( .A1(n22506), .A2(n11230), .Z(n15218) );
  XOR2_X1 U22183 ( .A1(n22622), .A2(n33990), .Z(n15610) );
  AOI22_X1 U22186 ( .A1(n10031), .A2(n30139), .B1(n19098), .B2(n30138), .ZN(
        n30140) );
  OR2_X1 U22188 ( .A1(n13786), .A2(n11700), .Z(n11022) );
  XOR2_X1 U22189 ( .A1(n13229), .A2(n1469), .Z(n10036) );
  XOR2_X1 U22193 ( .A1(n14388), .A2(n21097), .Z(n21096) );
  XOR2_X1 U22196 ( .A1(n28662), .A2(n10040), .Z(n13234) );
  XNOR2_X1 U22197 ( .A1(n15270), .A2(n29067), .ZN(n11127) );
  NOR2_X1 U22202 ( .A1(n27152), .A2(n19750), .ZN(n10393) );
  XOR2_X1 U22204 ( .A1(n29128), .A2(n29107), .Z(n11946) );
  INV_X1 U22217 ( .I(n27252), .ZN(n18717) );
  AND2_X1 U22220 ( .A1(n34561), .A2(n12612), .Z(n16779) );
  OAI21_X1 U22221 ( .A1(n34007), .A2(n32146), .B(n10058), .ZN(n28342) );
  NAND2_X1 U22223 ( .A1(n28068), .A2(n28067), .ZN(n13512) );
  XOR2_X1 U22224 ( .A1(n29836), .A2(n29839), .Z(n10059) );
  AOI21_X1 U22226 ( .A1(n28634), .A2(n28635), .B(n28633), .ZN(n10061) );
  XOR2_X1 U22231 ( .A1(n25257), .A2(n642), .Z(n10070) );
  XOR2_X1 U22233 ( .A1(n12356), .A2(n12354), .Z(n14405) );
  NAND3_X2 U22239 ( .A1(n18125), .A2(n21004), .A3(n28627), .ZN(n10080) );
  XOR2_X1 U22241 ( .A1(n29037), .A2(n10087), .Z(n11747) );
  NAND2_X1 U22242 ( .A1(n27138), .A2(n18074), .ZN(n18073) );
  XOR2_X1 U22245 ( .A1(n19289), .A2(n33866), .Z(n14569) );
  XOR2_X1 U22246 ( .A1(n29140), .A2(n19078), .Z(n10391) );
  NAND3_X1 U22248 ( .A1(n1202), .A2(n15704), .A3(n11676), .ZN(n15446) );
  NAND2_X1 U22253 ( .A1(n20965), .A2(n37306), .ZN(n26052) );
  NOR2_X1 U22265 ( .A1(n24814), .A2(n21231), .ZN(n10114) );
  XOR2_X1 U22267 ( .A1(Plaintext[17]), .A2(Key[17]), .Z(n11576) );
  XOR2_X1 U22269 ( .A1(n33178), .A2(n1165), .Z(n10131) );
  XOR2_X1 U22270 ( .A1(n10136), .A2(n10134), .Z(n10679) );
  XOR2_X1 U22276 ( .A1(n11724), .A2(n11725), .Z(n14471) );
  INV_X2 U22278 ( .I(n10155), .ZN(n19424) );
  AOI21_X1 U22285 ( .A1(n21322), .A2(n28119), .B(n28139), .ZN(n10167) );
  XOR2_X1 U22289 ( .A1(n27496), .A2(n12351), .Z(n10169) );
  INV_X2 U22291 ( .I(n12950), .ZN(n24274) );
  XOR2_X1 U22292 ( .A1(n10182), .A2(n10181), .Z(n12950) );
  XOR2_X1 U22294 ( .A1(n21227), .A2(n18683), .Z(n10182) );
  XOR2_X1 U22298 ( .A1(n10189), .A2(n29223), .Z(Ciphertext[10]) );
  XOR2_X1 U22302 ( .A1(n10197), .A2(n10196), .Z(n10195) );
  XOR2_X1 U22303 ( .A1(n35953), .A2(n19833), .Z(n10196) );
  XOR2_X1 U22304 ( .A1(n37312), .A2(n25226), .Z(n10197) );
  XOR2_X1 U22305 ( .A1(n10201), .A2(n16458), .Z(n10200) );
  XOR2_X1 U22307 ( .A1(Plaintext[177]), .A2(Key[177]), .Z(n10212) );
  NOR2_X1 U22308 ( .A1(n21730), .A2(n9863), .ZN(n21731) );
  XOR2_X1 U22310 ( .A1(n7287), .A2(n19516), .Z(n10214) );
  XOR2_X1 U22314 ( .A1(n27539), .A2(n27826), .Z(n10226) );
  XOR2_X1 U22327 ( .A1(n10240), .A2(n27761), .Z(n10673) );
  XOR2_X1 U22328 ( .A1(n27664), .A2(n19616), .Z(n10240) );
  AOI21_X1 U22331 ( .A1(n17411), .A2(n22252), .B(n10242), .ZN(n17408) );
  XOR2_X1 U22332 ( .A1(n10243), .A2(n10245), .Z(n26666) );
  XOR2_X1 U22333 ( .A1(n21034), .A2(n10244), .Z(n10243) );
  XOR2_X1 U22335 ( .A1(n19760), .A2(n33194), .Z(n10244) );
  XOR2_X1 U22336 ( .A1(n10246), .A2(n26085), .Z(n10245) );
  XOR2_X1 U22337 ( .A1(n12934), .A2(n26518), .Z(n10246) );
  INV_X2 U22338 ( .I(n10247), .ZN(n20077) );
  NAND2_X1 U22339 ( .A1(n38725), .A2(n20077), .ZN(n19054) );
  XOR2_X1 U22340 ( .A1(n17706), .A2(n10250), .Z(n10248) );
  XOR2_X1 U22341 ( .A1(n25149), .A2(n19670), .Z(n10250) );
  INV_X2 U22342 ( .I(n10251), .ZN(n24271) );
  XOR2_X1 U22343 ( .A1(n24064), .A2(n23073), .Z(n10252) );
  XOR2_X1 U22349 ( .A1(n10258), .A2(n12357), .Z(n12356) );
  XOR2_X1 U22355 ( .A1(n22749), .A2(n29647), .Z(n10267) );
  XOR2_X1 U22356 ( .A1(n18595), .A2(n22580), .Z(n10268) );
  XOR2_X1 U22358 ( .A1(n24033), .A2(n10276), .Z(n10275) );
  XOR2_X1 U22359 ( .A1(n19656), .A2(n30248), .Z(n10276) );
  XOR2_X1 U22361 ( .A1(n24022), .A2(n10279), .Z(n10278) );
  XOR2_X1 U22362 ( .A1(n23933), .A2(n15202), .Z(n24022) );
  NAND2_X1 U22363 ( .A1(n1084), .A2(n35750), .ZN(n17900) );
  INV_X2 U22364 ( .I(n10282), .ZN(n12953) );
  XOR2_X1 U22369 ( .A1(n17937), .A2(n23968), .Z(n12799) );
  NAND2_X2 U22370 ( .A1(n15073), .A2(n23228), .ZN(n23968) );
  XOR2_X1 U22375 ( .A1(n32931), .A2(n35318), .Z(n13750) );
  XOR2_X1 U22387 ( .A1(n10319), .A2(n10318), .Z(n10315) );
  XOR2_X1 U22389 ( .A1(n26584), .A2(n29474), .Z(n10318) );
  INV_X1 U22392 ( .I(n22209), .ZN(n22207) );
  OAI21_X2 U22394 ( .A1(n10325), .A2(n21759), .B(n10324), .ZN(n22354) );
  NAND2_X2 U22395 ( .A1(n19650), .A2(n21697), .ZN(n21759) );
  XOR2_X1 U22397 ( .A1(n35222), .A2(n1730), .Z(n10328) );
  XOR2_X1 U22398 ( .A1(n10333), .A2(n10330), .Z(n20595) );
  XOR2_X1 U22399 ( .A1(n10332), .A2(n10331), .Z(n10330) );
  XOR2_X1 U22400 ( .A1(n25182), .A2(n34848), .Z(n10331) );
  XOR2_X1 U22401 ( .A1(n6727), .A2(n25181), .Z(n10332) );
  XOR2_X1 U22405 ( .A1(n30856), .A2(n10343), .Z(n28854) );
  INV_X2 U22407 ( .I(n20883), .ZN(n21270) );
  XOR2_X1 U22412 ( .A1(n39548), .A2(n30063), .Z(n10364) );
  XOR2_X1 U22415 ( .A1(n10371), .A2(n16029), .Z(n10636) );
  XOR2_X1 U22421 ( .A1(n10387), .A2(n10386), .Z(n23992) );
  XOR2_X1 U22422 ( .A1(n15777), .A2(n10389), .Z(n10386) );
  XOR2_X1 U22423 ( .A1(n23981), .A2(n10388), .Z(n10387) );
  XOR2_X1 U22424 ( .A1(n36143), .A2(n35181), .Z(n10388) );
  XOR2_X1 U22425 ( .A1(n23982), .A2(n19498), .Z(n10389) );
  AOI21_X2 U22427 ( .A1(n10394), .A2(n27063), .B(n27062), .ZN(n28537) );
  XOR2_X1 U22432 ( .A1(n10400), .A2(n11464), .Z(n10534) );
  XOR2_X1 U22434 ( .A1(n10402), .A2(n24005), .Z(n10401) );
  XOR2_X1 U22436 ( .A1(n25161), .A2(n14687), .Z(n10406) );
  NAND2_X1 U22438 ( .A1(n30171), .A2(n30177), .ZN(n10410) );
  XOR2_X1 U22439 ( .A1(n10412), .A2(n18927), .Z(n27784) );
  XOR2_X1 U22444 ( .A1(n37094), .A2(n22621), .Z(n15608) );
  XOR2_X1 U22446 ( .A1(n18857), .A2(n663), .Z(n10426) );
  OAI21_X1 U22450 ( .A1(n29220), .A2(n29222), .B(n9914), .ZN(n10428) );
  XOR2_X1 U22451 ( .A1(n10430), .A2(n20560), .Z(n10658) );
  XOR2_X1 U22452 ( .A1(n12534), .A2(n19933), .Z(n10431) );
  XOR2_X1 U22458 ( .A1(n12251), .A2(n19131), .Z(n10447) );
  NAND3_X1 U22462 ( .A1(n21599), .A2(n16305), .A3(n21870), .ZN(n10649) );
  INV_X2 U22467 ( .I(n10455), .ZN(n23198) );
  OAI21_X1 U22469 ( .A1(n10051), .A2(n10461), .B(n20133), .ZN(n16966) );
  NOR2_X1 U22470 ( .A1(n10461), .A2(n27428), .ZN(n26941) );
  XOR2_X1 U22475 ( .A1(n10884), .A2(n10885), .Z(n10478) );
  XOR2_X1 U22477 ( .A1(n17284), .A2(n708), .Z(n10482) );
  XOR2_X1 U22480 ( .A1(n20304), .A2(n25291), .Z(n10486) );
  XOR2_X1 U22482 ( .A1(n26258), .A2(n38502), .Z(n26385) );
  XOR2_X1 U22483 ( .A1(n14386), .A2(n10493), .Z(n11661) );
  XOR2_X1 U22484 ( .A1(n11098), .A2(n29337), .Z(n10493) );
  XOR2_X1 U22487 ( .A1(n16743), .A2(n27785), .Z(n27494) );
  XOR2_X1 U22489 ( .A1(n22541), .A2(n669), .Z(n10502) );
  INV_X1 U22494 ( .I(n24829), .ZN(n18654) );
  XOR2_X1 U22495 ( .A1(n17935), .A2(n845), .Z(n10523) );
  INV_X2 U22498 ( .I(n10534), .ZN(n13444) );
  XOR2_X1 U22500 ( .A1(n32931), .A2(n19950), .Z(n10538) );
  XOR2_X1 U22506 ( .A1(n10541), .A2(n15071), .Z(n29495) );
  OAI21_X1 U22507 ( .A1(n37804), .A2(n36827), .B(n10542), .ZN(n14362) );
  NOR2_X1 U22508 ( .A1(n28690), .A2(n36827), .ZN(n28691) );
  XOR2_X1 U22510 ( .A1(n23898), .A2(n23779), .Z(n10548) );
  XOR2_X1 U22512 ( .A1(n23781), .A2(n12107), .Z(n10549) );
  XOR2_X1 U22518 ( .A1(n13083), .A2(n10561), .Z(n13082) );
  XOR2_X1 U22519 ( .A1(n10562), .A2(n27638), .Z(n10561) );
  XOR2_X1 U22520 ( .A1(n34345), .A2(n29875), .Z(n20047) );
  XOR2_X1 U22521 ( .A1(n37466), .A2(n1717), .Z(n15214) );
  XOR2_X1 U22522 ( .A1(n2383), .A2(n34345), .Z(n22432) );
  XOR2_X1 U22531 ( .A1(n10586), .A2(n664), .Z(n10585) );
  XOR2_X1 U22532 ( .A1(n1554), .A2(n24927), .Z(n10586) );
  XOR2_X1 U22537 ( .A1(n33216), .A2(n26334), .Z(n10593) );
  XOR2_X1 U22539 ( .A1(n29093), .A2(n29146), .Z(n29065) );
  NAND2_X2 U22540 ( .A1(n10596), .A2(n20430), .ZN(n29146) );
  INV_X2 U22543 ( .I(n14061), .ZN(n14408) );
  XOR2_X1 U22544 ( .A1(n10599), .A2(n10597), .Z(n14061) );
  XOR2_X1 U22545 ( .A1(n26204), .A2(n10598), .Z(n10597) );
  XOR2_X1 U22547 ( .A1(n26150), .A2(n16998), .Z(n10599) );
  XOR2_X1 U22552 ( .A1(n10616), .A2(n25027), .Z(n10615) );
  INV_X1 U22554 ( .I(n25959), .ZN(n25334) );
  XOR2_X1 U22556 ( .A1(n10620), .A2(n10619), .Z(n24307) );
  XOR2_X1 U22557 ( .A1(n24045), .A2(n24048), .Z(n10619) );
  XOR2_X1 U22558 ( .A1(n33690), .A2(n27736), .Z(n10706) );
  NAND2_X2 U22561 ( .A1(n21884), .A2(n13856), .ZN(n22042) );
  XNOR2_X1 U22566 ( .A1(Plaintext[96]), .A2(Key[96]), .ZN(n10629) );
  XNOR2_X1 U22580 ( .A1(Plaintext[100]), .A2(Key[100]), .ZN(n10656) );
  MUX2_X1 U22582 ( .I0(n11034), .I1(n2678), .S(n910), .Z(n11036) );
  XOR2_X1 U22583 ( .A1(n19956), .A2(n10663), .Z(n10662) );
  XOR2_X1 U22584 ( .A1(n30322), .A2(n19717), .Z(n10663) );
  NOR2_X1 U22585 ( .A1(n15282), .A2(n10667), .ZN(n12409) );
  XOR2_X1 U22589 ( .A1(n17937), .A2(n1366), .Z(n10684) );
  XOR2_X1 U22593 ( .A1(n13245), .A2(n27534), .Z(n10707) );
  XOR2_X1 U22594 ( .A1(n35268), .A2(n19910), .Z(n11401) );
  XOR2_X1 U22595 ( .A1(n1614), .A2(n35181), .Z(n22957) );
  XOR2_X1 U22596 ( .A1(n10717), .A2(n10714), .Z(n21031) );
  XOR2_X1 U22597 ( .A1(n10715), .A2(n10716), .Z(n10714) );
  XOR2_X1 U22598 ( .A1(n35268), .A2(n20748), .Z(n10715) );
  XOR2_X1 U22599 ( .A1(n7250), .A2(n19096), .Z(n10716) );
  INV_X1 U22600 ( .I(n33178), .ZN(n10718) );
  XOR2_X1 U22601 ( .A1(n36596), .A2(n19674), .Z(n22518) );
  OAI21_X1 U22606 ( .A1(n31564), .A2(n38839), .B(n20864), .ZN(n23962) );
  XOR2_X1 U22609 ( .A1(n10737), .A2(n14101), .Z(n14170) );
  AOI21_X1 U22611 ( .A1(n22045), .A2(n38448), .B(n10743), .ZN(n10742) );
  XOR2_X1 U22614 ( .A1(n14023), .A2(n18992), .Z(n10748) );
  XOR2_X1 U22618 ( .A1(n8402), .A2(n1051), .Z(n10766) );
  OR2_X1 U22626 ( .A1(n24872), .A2(n31161), .Z(n10773) );
  NAND2_X1 U22629 ( .A1(n21256), .A2(n9178), .ZN(n21255) );
  XOR2_X1 U22632 ( .A1(n39320), .A2(n25086), .Z(n15126) );
  XOR2_X1 U22636 ( .A1(n38950), .A2(n10791), .Z(n25000) );
  XOR2_X1 U22637 ( .A1(n10791), .A2(n19808), .Z(n19986) );
  XOR2_X1 U22638 ( .A1(n10797), .A2(n16783), .Z(n11503) );
  OAI21_X1 U22641 ( .A1(n13107), .A2(n10803), .B(n29224), .ZN(n29226) );
  INV_X2 U22646 ( .I(n10810), .ZN(n12235) );
  INV_X2 U22647 ( .I(n16931), .ZN(n18164) );
  INV_X2 U22649 ( .I(n10816), .ZN(n14158) );
  XOR2_X1 U22650 ( .A1(n27757), .A2(n12769), .Z(n10819) );
  XOR2_X1 U22652 ( .A1(n26441), .A2(n29857), .Z(n10823) );
  XOR2_X1 U22653 ( .A1(n26438), .A2(n6131), .Z(n26523) );
  XOR2_X1 U22654 ( .A1(n28928), .A2(n10830), .Z(n10829) );
  XOR2_X1 U22655 ( .A1(n28927), .A2(n10794), .Z(n10830) );
  AOI21_X1 U22656 ( .A1(n10831), .A2(n17750), .B(n17748), .ZN(n17747) );
  NOR2_X1 U22657 ( .A1(n39454), .A2(n32979), .ZN(n25749) );
  INV_X2 U22658 ( .I(n10835), .ZN(n11150) );
  XOR2_X1 U22662 ( .A1(n26450), .A2(n17858), .Z(n10855) );
  XOR2_X1 U22663 ( .A1(n22688), .A2(n10859), .Z(n10858) );
  XOR2_X1 U22664 ( .A1(n5203), .A2(n19843), .Z(n10859) );
  XOR2_X1 U22668 ( .A1(n27606), .A2(n10864), .Z(n10863) );
  XOR2_X1 U22669 ( .A1(n27776), .A2(n29849), .Z(n10864) );
  XOR2_X1 U22673 ( .A1(n3649), .A2(n35169), .Z(n25044) );
  XOR2_X1 U22674 ( .A1(n32195), .A2(n3649), .Z(n17879) );
  XOR2_X1 U22675 ( .A1(n10872), .A2(n10874), .Z(n13248) );
  XOR2_X1 U22679 ( .A1(n9344), .A2(n23996), .Z(n10874) );
  XOR2_X1 U22686 ( .A1(n21093), .A2(n1367), .Z(n27808) );
  XOR2_X1 U22687 ( .A1(n27858), .A2(n21093), .Z(n15068) );
  XOR2_X1 U22688 ( .A1(n21093), .A2(n27781), .Z(n27615) );
  XOR2_X1 U22689 ( .A1(n39636), .A2(n1375), .Z(n10884) );
  XOR2_X1 U22691 ( .A1(n20509), .A2(n33452), .Z(n10887) );
  XOR2_X1 U22696 ( .A1(n10898), .A2(n764), .Z(n10897) );
  XOR2_X1 U22697 ( .A1(n33961), .A2(n35249), .Z(n10898) );
  XOR2_X1 U22699 ( .A1(n25247), .A2(n29554), .Z(n10905) );
  INV_X2 U22706 ( .I(n10925), .ZN(n18450) );
  INV_X1 U22711 ( .I(Plaintext[59]), .ZN(n10929) );
  NOR2_X1 U22713 ( .A1(n1416), .A2(n2022), .ZN(n18701) );
  AOI22_X1 U22714 ( .A1(n33100), .A2(n9597), .B1(n18571), .B2(n20197), .ZN(
        n28409) );
  XOR2_X1 U22728 ( .A1(n17999), .A2(n656), .Z(n10955) );
  XOR2_X1 U22730 ( .A1(n23774), .A2(n23680), .Z(n10957) );
  XOR2_X1 U22735 ( .A1(n10967), .A2(n10966), .Z(n18933) );
  XOR2_X1 U22736 ( .A1(n26222), .A2(n18934), .Z(n10966) );
  XOR2_X1 U22737 ( .A1(n10965), .A2(n26359), .Z(n26222) );
  OR2_X1 U22740 ( .A1(n19159), .A2(n10979), .Z(n19158) );
  XOR2_X1 U22743 ( .A1(n13374), .A2(n11755), .Z(n10983) );
  XOR2_X1 U22744 ( .A1(n27807), .A2(n27808), .Z(n10984) );
  XOR2_X1 U22746 ( .A1(n10987), .A2(n29474), .Z(n24929) );
  XOR2_X1 U22747 ( .A1(n10987), .A2(n16460), .Z(n17836) );
  XOR2_X1 U22750 ( .A1(n18180), .A2(n30114), .Z(n13064) );
  XOR2_X1 U22760 ( .A1(n15617), .A2(n29300), .Z(n11016) );
  NOR2_X1 U22765 ( .A1(n25533), .A2(n9594), .ZN(n11018) );
  NOR2_X1 U22768 ( .A1(n11020), .A2(n15135), .ZN(n27589) );
  XOR2_X1 U22773 ( .A1(n27697), .A2(n27503), .Z(n27826) );
  NOR2_X1 U22775 ( .A1(n30758), .A2(n17095), .ZN(n11043) );
  INV_X2 U22776 ( .I(n11046), .ZN(n19696) );
  NAND2_X2 U22781 ( .A1(n21242), .A2(n21241), .ZN(n17986) );
  AOI21_X1 U22787 ( .A1(n15958), .A2(n12943), .B(n11067), .ZN(n15956) );
  XOR2_X1 U22789 ( .A1(n12393), .A2(n29857), .Z(n14505) );
  XOR2_X1 U22792 ( .A1(Plaintext[153]), .A2(Key[153]), .Z(n15009) );
  XOR2_X1 U22794 ( .A1(n29090), .A2(n11075), .Z(n11074) );
  XOR2_X1 U22795 ( .A1(n296), .A2(n29808), .Z(n11075) );
  XOR2_X1 U22796 ( .A1(n29022), .A2(n11077), .Z(n11076) );
  INV_X1 U22798 ( .I(n24152), .ZN(n21148) );
  XOR2_X1 U22799 ( .A1(n11372), .A2(n24011), .Z(n23915) );
  XOR2_X1 U22800 ( .A1(n11372), .A2(n19947), .Z(n17725) );
  XNOR2_X1 U22804 ( .A1(n16742), .A2(n16740), .ZN(n11084) );
  OAI21_X2 U22806 ( .A1(n27902), .A2(n21020), .B(n16994), .ZN(n28689) );
  XOR2_X1 U22807 ( .A1(n11098), .A2(n29411), .Z(n23316) );
  XOR2_X1 U22808 ( .A1(n23695), .A2(n11098), .Z(n15974) );
  XOR2_X1 U22810 ( .A1(n11102), .A2(n25075), .Z(n11103) );
  XOR2_X1 U22814 ( .A1(n11115), .A2(n23977), .Z(n11114) );
  NOR2_X1 U22819 ( .A1(n11120), .A2(n16619), .ZN(n18971) );
  NAND2_X1 U22821 ( .A1(n25998), .A2(n39165), .ZN(n25842) );
  NAND2_X1 U22831 ( .A1(n20328), .A2(n11146), .ZN(n17219) );
  XOR2_X1 U22832 ( .A1(n16254), .A2(n649), .Z(n22412) );
  NAND3_X2 U22834 ( .A1(n16028), .A2(n21998), .A3(n18401), .ZN(n22644) );
  OAI22_X2 U22836 ( .A1(n12546), .A2(n11239), .B1(n11238), .B2(n543), .ZN(
        n11149) );
  NOR2_X1 U22837 ( .A1(n11149), .A2(n19515), .ZN(n13899) );
  XOR2_X1 U22838 ( .A1(n28966), .A2(n28968), .Z(n11151) );
  XOR2_X1 U22840 ( .A1(n679), .A2(n11153), .Z(n11152) );
  XOR2_X1 U22841 ( .A1(n10129), .A2(n11155), .Z(n11154) );
  XOR2_X1 U22845 ( .A1(n11267), .A2(n722), .Z(n11165) );
  OAI21_X2 U22852 ( .A1(n14189), .A2(n14188), .B(n14186), .ZN(n17511) );
  XOR2_X1 U22858 ( .A1(n11200), .A2(Plaintext[178]), .Z(n13996) );
  XOR2_X1 U22860 ( .A1(n11201), .A2(n3953), .Z(n22694) );
  XOR2_X1 U22866 ( .A1(n27865), .A2(n11211), .Z(n11210) );
  XOR2_X1 U22867 ( .A1(n20454), .A2(n27738), .Z(n11211) );
  INV_X1 U22871 ( .I(n11214), .ZN(n18746) );
  NAND2_X2 U22872 ( .A1(n11218), .A2(n11217), .ZN(n17192) );
  XOR2_X1 U22877 ( .A1(n11233), .A2(n22291), .Z(n22506) );
  XOR2_X1 U22879 ( .A1(n11236), .A2(n27479), .Z(n11235) );
  NAND2_X1 U22882 ( .A1(n15299), .A2(n7577), .ZN(n23249) );
  XOR2_X1 U22883 ( .A1(n11255), .A2(n11254), .Z(n11253) );
  OAI21_X2 U22885 ( .A1(n26940), .A2(n26939), .B(n26938), .ZN(n27184) );
  OAI21_X1 U22886 ( .A1(n13971), .A2(n7317), .B(n11257), .ZN(n25955) );
  XOR2_X1 U22887 ( .A1(n518), .A2(n1051), .Z(n20592) );
  XOR2_X1 U22888 ( .A1(n1558), .A2(n13531), .Z(n13530) );
  NOR2_X1 U22889 ( .A1(n15049), .A2(n1275), .ZN(n11261) );
  NAND2_X1 U22891 ( .A1(n14492), .A2(n11274), .ZN(n16165) );
  XOR2_X1 U22892 ( .A1(Plaintext[95]), .A2(Key[95]), .Z(n15354) );
  XOR2_X1 U22898 ( .A1(n22688), .A2(n11289), .Z(n11288) );
  XOR2_X1 U22899 ( .A1(n22544), .A2(n22409), .Z(n11290) );
  INV_X1 U22901 ( .I(Plaintext[160]), .ZN(n11291) );
  XOR2_X1 U22902 ( .A1(n11291), .A2(Key[160]), .Z(n12036) );
  XOR2_X1 U22905 ( .A1(n22524), .A2(n22523), .Z(n22857) );
  AOI21_X2 U22907 ( .A1(n21636), .A2(n11303), .B(n11302), .ZN(n11304) );
  XOR2_X1 U22909 ( .A1(n11311), .A2(n11310), .Z(n11309) );
  XOR2_X1 U22910 ( .A1(n22621), .A2(n19953), .Z(n11310) );
  XOR2_X1 U22912 ( .A1(n11314), .A2(n11313), .Z(n11312) );
  XOR2_X1 U22913 ( .A1(n9116), .A2(n19221), .Z(n11313) );
  XOR2_X1 U22915 ( .A1(n14304), .A2(n1745), .Z(n21201) );
  INV_X2 U22916 ( .I(n15051), .ZN(n25543) );
  XOR2_X1 U22918 ( .A1(n11321), .A2(n25218), .Z(n25219) );
  OAI22_X2 U22924 ( .A1(n24689), .A2(n24690), .B1(n10019), .B2(n13002), .ZN(
        n25237) );
  NAND2_X1 U22926 ( .A1(n1314), .A2(n33745), .ZN(n15081) );
  XOR2_X1 U22929 ( .A1(n24994), .A2(n25127), .Z(n25171) );
  XOR2_X1 U22933 ( .A1(n15270), .A2(n5755), .Z(n11346) );
  XOR2_X1 U22936 ( .A1(n22606), .A2(n11356), .Z(n11355) );
  XOR2_X1 U22937 ( .A1(n22699), .A2(n11308), .Z(n11356) );
  XOR2_X1 U22941 ( .A1(n33027), .A2(n26554), .Z(n26307) );
  XOR2_X1 U22942 ( .A1(n33027), .A2(n19464), .Z(n20539) );
  XOR2_X1 U22943 ( .A1(n38937), .A2(n1374), .Z(n11365) );
  XOR2_X1 U22950 ( .A1(n11377), .A2(n11376), .Z(n23122) );
  XOR2_X1 U22951 ( .A1(n16278), .A2(n22646), .Z(n11376) );
  XOR2_X1 U22952 ( .A1(n22643), .A2(n22644), .Z(n16278) );
  XOR2_X1 U22958 ( .A1(n20294), .A2(n22636), .Z(n11382) );
  XOR2_X1 U22960 ( .A1(n11384), .A2(n28814), .Z(n11783) );
  INV_X1 U22961 ( .I(n37295), .ZN(n28769) );
  XOR2_X1 U22964 ( .A1(n27773), .A2(n31295), .Z(n11391) );
  XOR2_X1 U22965 ( .A1(n27774), .A2(n36384), .Z(n11392) );
  NAND2_X1 U22969 ( .A1(n19090), .A2(n19085), .ZN(n11397) );
  XOR2_X1 U22974 ( .A1(n14843), .A2(n11405), .Z(n11406) );
  NAND2_X1 U22975 ( .A1(n11406), .A2(n12049), .ZN(n15293) );
  XOR2_X1 U22978 ( .A1(n11419), .A2(n11417), .Z(n11416) );
  XOR2_X1 U22979 ( .A1(n30964), .A2(n11418), .Z(n11417) );
  INV_X1 U22980 ( .I(n28851), .ZN(n11418) );
  XOR2_X1 U22981 ( .A1(n13639), .A2(n15745), .Z(n11419) );
  XOR2_X1 U22987 ( .A1(n11425), .A2(n29974), .Z(n17760) );
  XOR2_X1 U22988 ( .A1(n4622), .A2(n11425), .Z(n12587) );
  XOR2_X1 U22989 ( .A1(n35065), .A2(n23880), .Z(n23737) );
  XOR2_X1 U22990 ( .A1(n22416), .A2(n1657), .Z(n12205) );
  NAND2_X2 U22995 ( .A1(n30128), .A2(n20274), .ZN(n30127) );
  XOR2_X1 U23001 ( .A1(n27539), .A2(n27029), .Z(n11458) );
  INV_X2 U23002 ( .I(n11459), .ZN(n12257) );
  INV_X1 U23005 ( .I(n23926), .ZN(n11464) );
  NAND2_X1 U23006 ( .A1(n26829), .A2(n11467), .ZN(n21182) );
  NAND3_X2 U23007 ( .A1(n11473), .A2(n23180), .A3(n11472), .ZN(n23631) );
  XOR2_X1 U23010 ( .A1(n25194), .A2(n1706), .Z(n11475) );
  NAND2_X2 U23011 ( .A1(n18393), .A2(n18394), .ZN(n25194) );
  NAND2_X1 U23012 ( .A1(n11476), .A2(n22722), .ZN(n22730) );
  NAND2_X1 U23013 ( .A1(n37954), .A2(n24328), .ZN(n11477) );
  INV_X2 U23018 ( .I(n11482), .ZN(n17240) );
  NOR2_X1 U23020 ( .A1(n24206), .A2(n37264), .ZN(n11494) );
  INV_X2 U23025 ( .I(n18502), .ZN(n11506) );
  XOR2_X1 U23030 ( .A1(n11519), .A2(n11520), .Z(n13018) );
  XOR2_X1 U23032 ( .A1(n25162), .A2(n24945), .Z(n11520) );
  NOR2_X1 U23034 ( .A1(n26666), .A2(n924), .ZN(n11523) );
  NAND3_X1 U23041 ( .A1(n31523), .A2(n39729), .A3(n33237), .ZN(n26094) );
  NAND2_X1 U23042 ( .A1(n17008), .A2(n11533), .ZN(n20833) );
  XOR2_X1 U23052 ( .A1(n1258), .A2(n11554), .Z(n11553) );
  NAND2_X1 U23053 ( .A1(n11556), .A2(n11555), .ZN(n11554) );
  OAI21_X1 U23054 ( .A1(n24495), .A2(n24496), .B(n19128), .ZN(n11555) );
  NAND2_X1 U23055 ( .A1(n11558), .A2(n11557), .ZN(n11556) );
  NOR2_X1 U23056 ( .A1(n24496), .A2(n19128), .ZN(n11557) );
  INV_X1 U23057 ( .I(n24495), .ZN(n11558) );
  XOR2_X1 U23058 ( .A1(n38213), .A2(n13054), .Z(n11559) );
  INV_X1 U23061 ( .I(n20840), .ZN(n23175) );
  XOR2_X1 U23063 ( .A1(n19072), .A2(n11572), .Z(n11571) );
  XOR2_X1 U23064 ( .A1(n25242), .A2(n25241), .Z(n11572) );
  XOR2_X1 U23067 ( .A1(n13439), .A2(n17423), .Z(n23953) );
  XOR2_X1 U23068 ( .A1(n27607), .A2(n27707), .Z(n27608) );
  NAND2_X1 U23070 ( .A1(n5892), .A2(n35994), .ZN(n23036) );
  INV_X2 U23071 ( .I(n11586), .ZN(n14379) );
  AND2_X1 U23073 ( .A1(n29237), .A2(n12141), .Z(n14529) );
  XOR2_X1 U23076 ( .A1(n14425), .A2(n11603), .Z(n11602) );
  XOR2_X1 U23079 ( .A1(n11612), .A2(n11611), .Z(n12103) );
  XOR2_X1 U23080 ( .A1(n2281), .A2(n27534), .Z(n11611) );
  XOR2_X1 U23082 ( .A1(n19608), .A2(n39559), .Z(n11615) );
  XOR2_X1 U23084 ( .A1(n12824), .A2(n26350), .Z(n11621) );
  INV_X2 U23086 ( .I(n11622), .ZN(n14436) );
  INV_X2 U23090 ( .I(n11627), .ZN(n15163) );
  INV_X4 U23091 ( .I(n13609), .ZN(n11628) );
  INV_X2 U23092 ( .I(n13787), .ZN(n13609) );
  NAND2_X1 U23097 ( .A1(n20092), .A2(n27438), .ZN(n11637) );
  XOR2_X1 U23099 ( .A1(n10213), .A2(n11644), .Z(n22662) );
  XOR2_X1 U23100 ( .A1(n11644), .A2(n1375), .Z(n14609) );
  XOR2_X1 U23101 ( .A1(n15448), .A2(n11644), .Z(n20350) );
  INV_X2 U23105 ( .I(n11663), .ZN(n15320) );
  NAND2_X1 U23108 ( .A1(n5657), .A2(n22889), .ZN(n23509) );
  XOR2_X1 U23114 ( .A1(n30068), .A2(n24932), .Z(n11688) );
  XOR2_X1 U23115 ( .A1(n25133), .A2(n37296), .Z(n11689) );
  XOR2_X1 U23120 ( .A1(n11694), .A2(n29269), .Z(n27477) );
  XOR2_X1 U23121 ( .A1(n27669), .A2(n282), .Z(n18548) );
  XOR2_X1 U23123 ( .A1(n3703), .A2(n3665), .Z(n28662) );
  XOR2_X1 U23124 ( .A1(n11698), .A2(n30170), .Z(n17134) );
  XOR2_X1 U23125 ( .A1(n12534), .A2(n11698), .Z(n25295) );
  XOR2_X1 U23126 ( .A1(n24978), .A2(n11698), .Z(n19073) );
  INV_X2 U23127 ( .I(n11699), .ZN(n20517) );
  NOR2_X1 U23129 ( .A1(n22901), .A2(n11704), .ZN(n22468) );
  AND2_X1 U23133 ( .A1(n15540), .A2(n31418), .Z(n11718) );
  XOR2_X1 U23136 ( .A1(n23663), .A2(n15094), .Z(n11725) );
  OAI21_X1 U23137 ( .A1(n26954), .A2(n26957), .B(n11726), .ZN(n13097) );
  NAND3_X1 U23142 ( .A1(n30621), .A2(n425), .A3(n11734), .ZN(n25404) );
  INV_X1 U23143 ( .I(n26521), .ZN(n26347) );
  OAI21_X2 U23147 ( .A1(n14503), .A2(n17125), .B(n26218), .ZN(n26407) );
  XOR2_X1 U23149 ( .A1(n29036), .A2(n29035), .Z(n11746) );
  XOR2_X1 U23150 ( .A1(n11750), .A2(n11748), .Z(n16593) );
  XOR2_X1 U23151 ( .A1(n5463), .A2(n11749), .Z(n11748) );
  XOR2_X1 U23152 ( .A1(n22531), .A2(n11974), .Z(n11749) );
  XOR2_X1 U23154 ( .A1(n37951), .A2(n31591), .Z(n16695) );
  XOR2_X1 U23156 ( .A1(n11756), .A2(n25278), .Z(n25279) );
  XOR2_X1 U23157 ( .A1(n39541), .A2(n11756), .Z(n11905) );
  NAND2_X2 U23161 ( .A1(n25573), .A2(n25572), .ZN(n26116) );
  XOR2_X1 U23164 ( .A1(n22533), .A2(n22462), .Z(n11779) );
  NOR2_X2 U23166 ( .A1(n21103), .A2(n21104), .ZN(n22582) );
  OAI21_X2 U23167 ( .A1(n22010), .A2(n21105), .B(n14683), .ZN(n18778) );
  INV_X2 U23168 ( .I(n11780), .ZN(n12931) );
  OR2_X1 U23170 ( .A1(n11783), .A2(n20522), .Z(n29010) );
  XOR2_X1 U23172 ( .A1(n11790), .A2(n11788), .Z(n21187) );
  XOR2_X1 U23173 ( .A1(n28979), .A2(n11789), .Z(n11788) );
  XOR2_X1 U23174 ( .A1(n36905), .A2(n19932), .Z(n11789) );
  XOR2_X1 U23175 ( .A1(n28984), .A2(n19600), .Z(n11790) );
  XOR2_X1 U23177 ( .A1(n22717), .A2(n22514), .Z(n11791) );
  XOR2_X1 U23180 ( .A1(n22515), .A2(n1371), .Z(n11793) );
  NOR2_X1 U23185 ( .A1(n18029), .A2(n25614), .ZN(n12096) );
  INV_X4 U23186 ( .I(n39827), .ZN(n29185) );
  AND2_X1 U23188 ( .A1(n7693), .A2(n19868), .Z(n20690) );
  NAND3_X1 U23192 ( .A1(n22212), .A2(n22213), .A3(n22361), .ZN(n11921) );
  XOR2_X1 U23195 ( .A1(n963), .A2(n29983), .Z(n16061) );
  XOR2_X1 U23196 ( .A1(n963), .A2(n19730), .Z(n22720) );
  XOR2_X1 U23198 ( .A1(n24023), .A2(n29875), .Z(n23806) );
  XOR2_X1 U23202 ( .A1(n22595), .A2(n37042), .Z(n11809) );
  XOR2_X1 U23206 ( .A1(n31181), .A2(n29785), .Z(n12180) );
  XOR2_X1 U23207 ( .A1(n31181), .A2(n30010), .Z(n19074) );
  XOR2_X1 U23208 ( .A1(n35972), .A2(n19845), .Z(n24950) );
  XOR2_X1 U23211 ( .A1(n507), .A2(n14969), .Z(n24588) );
  XOR2_X1 U23216 ( .A1(n6559), .A2(n13617), .Z(n19984) );
  XOR2_X1 U23217 ( .A1(n16639), .A2(n32836), .Z(n14487) );
  NAND2_X2 U23219 ( .A1(n13913), .A2(n14658), .ZN(n23515) );
  AOI21_X2 U23224 ( .A1(n21653), .A2(n11850), .B(n11849), .ZN(n19737) );
  INV_X2 U23230 ( .I(n13499), .ZN(n28141) );
  XOR2_X1 U23232 ( .A1(n27474), .A2(n15068), .Z(n11871) );
  XOR2_X1 U23238 ( .A1(n1410), .A2(n15780), .Z(n11883) );
  OAI21_X1 U23242 ( .A1(n11890), .A2(n28123), .B(n11891), .ZN(n11895) );
  INV_X1 U23245 ( .I(Plaintext[169]), .ZN(n11901) );
  NAND2_X1 U23251 ( .A1(n13512), .A2(n36877), .ZN(n14766) );
  XOR2_X1 U23254 ( .A1(n16566), .A2(n11926), .Z(n11925) );
  XOR2_X1 U23255 ( .A1(n35202), .A2(n19874), .Z(n11926) );
  XOR2_X1 U23258 ( .A1(n18051), .A2(n35200), .Z(n14285) );
  XOR2_X1 U23262 ( .A1(n11962), .A2(n11961), .Z(n11960) );
  XOR2_X1 U23263 ( .A1(n33038), .A2(n19770), .Z(n11961) );
  XOR2_X1 U23264 ( .A1(n25071), .A2(n10273), .Z(n11962) );
  NAND2_X2 U23265 ( .A1(n20697), .A2(n11963), .ZN(n25071) );
  XOR2_X1 U23266 ( .A1(n14258), .A2(n11965), .Z(n12612) );
  XOR2_X1 U23267 ( .A1(n11966), .A2(n23795), .Z(n11965) );
  XOR2_X1 U23268 ( .A1(n36842), .A2(n29394), .Z(n11966) );
  INV_X2 U23271 ( .I(n11975), .ZN(n13770) );
  XOR2_X1 U23273 ( .A1(n27788), .A2(n11977), .Z(n11976) );
  XOR2_X1 U23274 ( .A1(n17884), .A2(n21226), .Z(n11977) );
  XOR2_X1 U23281 ( .A1(n22677), .A2(n22715), .Z(n11984) );
  XOR2_X1 U23282 ( .A1(n20980), .A2(n22675), .Z(n11985) );
  NAND2_X1 U23283 ( .A1(n11987), .A2(n11986), .ZN(n14140) );
  NAND3_X1 U23284 ( .A1(n36701), .A2(n36011), .A3(n1695), .ZN(n11986) );
  XOR2_X1 U23287 ( .A1(n38641), .A2(n25090), .Z(n11989) );
  XOR2_X1 U23291 ( .A1(n27564), .A2(n27640), .Z(n11994) );
  XOR2_X1 U23292 ( .A1(n26221), .A2(n26143), .Z(n11998) );
  XOR2_X1 U23293 ( .A1(n26454), .A2(n26413), .Z(n11999) );
  XOR2_X1 U23294 ( .A1(n12000), .A2(n18869), .Z(n12001) );
  NAND2_X1 U23295 ( .A1(n2771), .A2(n37984), .ZN(n22826) );
  NAND2_X2 U23302 ( .A1(n12025), .A2(n12024), .ZN(n19773) );
  XOR2_X1 U23306 ( .A1(n13430), .A2(n639), .Z(n23196) );
  AOI22_X2 U23307 ( .A1(n25819), .A2(n25940), .B1(n25817), .B2(n25818), .ZN(
        n20600) );
  INV_X2 U23310 ( .I(n12036), .ZN(n21770) );
  XOR2_X1 U23313 ( .A1(n18924), .A2(n35178), .Z(n15222) );
  NAND2_X2 U23318 ( .A1(n8127), .A2(n24668), .ZN(n18858) );
  XOR2_X1 U23321 ( .A1(n26160), .A2(n31605), .Z(n12053) );
  XOR2_X1 U23330 ( .A1(n25170), .A2(n24958), .Z(n12076) );
  INV_X1 U23331 ( .I(n21213), .ZN(n23638) );
  NAND2_X2 U23333 ( .A1(n1424), .A2(n496), .ZN(n28544) );
  INV_X1 U23336 ( .I(n24162), .ZN(n24173) );
  XOR2_X1 U23337 ( .A1(n12086), .A2(n12085), .Z(n12084) );
  XOR2_X1 U23338 ( .A1(n33323), .A2(n19845), .Z(n12085) );
  XOR2_X1 U23339 ( .A1(n22668), .A2(n7432), .Z(n12086) );
  XOR2_X1 U23344 ( .A1(n23778), .A2(n19910), .Z(n12107) );
  XOR2_X1 U23345 ( .A1(Plaintext[82]), .A2(Key[82]), .Z(n12670) );
  NAND2_X1 U23346 ( .A1(n9916), .A2(n25813), .ZN(n13678) );
  XOR2_X1 U23349 ( .A1(n12113), .A2(n12112), .Z(n12111) );
  XOR2_X1 U23350 ( .A1(n26455), .A2(n31771), .Z(n12112) );
  NAND3_X2 U23351 ( .A1(n26095), .A2(n26096), .A3(n26094), .ZN(n26455) );
  XOR2_X1 U23352 ( .A1(n26403), .A2(n26541), .Z(n12113) );
  NAND2_X2 U23353 ( .A1(n12490), .A2(n12489), .ZN(n26541) );
  NOR2_X1 U23356 ( .A1(n26185), .A2(n38185), .ZN(n12115) );
  OAI21_X1 U23359 ( .A1(n15456), .A2(n18152), .B(n21840), .ZN(n12118) );
  NAND2_X1 U23360 ( .A1(n23111), .A2(n20783), .ZN(n12123) );
  XOR2_X1 U23362 ( .A1(n10329), .A2(n731), .Z(n12132) );
  NAND2_X1 U23363 ( .A1(n9913), .A2(n7303), .ZN(n12547) );
  OAI22_X1 U23364 ( .A1(n29462), .A2(n7303), .B1(n29464), .B2(n969), .ZN(
        n13431) );
  XOR2_X1 U23369 ( .A1(n7148), .A2(n19722), .Z(n12139) );
  NAND3_X1 U23370 ( .A1(n1388), .A2(n35185), .A3(n29236), .ZN(n29233) );
  NOR2_X1 U23371 ( .A1(n1388), .A2(n35185), .ZN(n15028) );
  NAND3_X2 U23373 ( .A1(n25950), .A2(n25949), .A3(n12151), .ZN(n26438) );
  OAI22_X2 U23375 ( .A1(n20996), .A2(n133), .B1(n22047), .B2(n21973), .ZN(
        n22188) );
  XOR2_X1 U23382 ( .A1(n557), .A2(n19890), .Z(n12165) );
  XOR2_X1 U23385 ( .A1(n35065), .A2(n1165), .Z(n23674) );
  XOR2_X1 U23390 ( .A1(n23745), .A2(n12184), .Z(n12183) );
  XOR2_X1 U23391 ( .A1(n23789), .A2(n35235), .Z(n12184) );
  XOR2_X1 U23392 ( .A1(n12185), .A2(n20093), .Z(n28250) );
  XOR2_X1 U23393 ( .A1(n379), .A2(n37242), .Z(n12185) );
  XOR2_X1 U23400 ( .A1(n22750), .A2(n12197), .Z(n12196) );
  XOR2_X1 U23401 ( .A1(n35824), .A2(n29506), .Z(n12197) );
  NAND2_X1 U23402 ( .A1(n30106), .A2(n18829), .ZN(n12204) );
  INV_X2 U23405 ( .I(n18188), .ZN(n19435) );
  INV_X2 U23406 ( .I(n15774), .ZN(n19667) );
  INV_X2 U23412 ( .I(n12225), .ZN(n18412) );
  XOR2_X1 U23413 ( .A1(n22695), .A2(n36362), .Z(n20048) );
  XOR2_X1 U23415 ( .A1(n30865), .A2(n12233), .Z(n24525) );
  XOR2_X1 U23417 ( .A1(Plaintext[176]), .A2(Key[176]), .Z(n12535) );
  XOR2_X1 U23418 ( .A1(n15286), .A2(n27843), .Z(n12432) );
  XOR2_X1 U23420 ( .A1(n12243), .A2(n19876), .Z(n22545) );
  XOR2_X1 U23422 ( .A1(n19516), .A2(n39536), .Z(n28493) );
  XOR2_X1 U23429 ( .A1(n24043), .A2(n23892), .Z(n12265) );
  XOR2_X1 U23430 ( .A1(n21316), .A2(n23656), .Z(n12266) );
  INV_X2 U23431 ( .I(n12759), .ZN(n24232) );
  XOR2_X1 U23432 ( .A1(n12267), .A2(n30122), .Z(n21225) );
  XOR2_X1 U23433 ( .A1(n21227), .A2(n12973), .Z(n18582) );
  NOR2_X1 U23434 ( .A1(n16224), .A2(n29935), .ZN(n12273) );
  NOR2_X1 U23441 ( .A1(n23226), .A2(n12289), .ZN(n16394) );
  NAND2_X1 U23442 ( .A1(n23226), .A2(n12289), .ZN(n15075) );
  NOR2_X1 U23444 ( .A1(n31331), .A2(n12289), .ZN(n23278) );
  XOR2_X1 U23452 ( .A1(n17884), .A2(n29442), .Z(n15726) );
  XOR2_X1 U23453 ( .A1(n12970), .A2(n17884), .Z(n12969) );
  INV_X2 U23454 ( .I(n12302), .ZN(n20739) );
  NOR2_X1 U23457 ( .A1(n12306), .A2(n27233), .ZN(n27234) );
  XOR2_X1 U23460 ( .A1(n25089), .A2(n25088), .Z(n12310) );
  XOR2_X1 U23464 ( .A1(n12316), .A2(n1377), .Z(Ciphertext[47]) );
  AOI21_X1 U23465 ( .A1(n15841), .A2(n12318), .B(n11506), .ZN(n12317) );
  NAND2_X1 U23466 ( .A1(n29439), .A2(n29438), .ZN(n12318) );
  INV_X2 U23472 ( .I(n12334), .ZN(n14399) );
  XOR2_X1 U23475 ( .A1(n6522), .A2(n12337), .Z(n12834) );
  XOR2_X1 U23476 ( .A1(n9576), .A2(n33184), .Z(n12337) );
  INV_X1 U23480 ( .I(n17777), .ZN(n20632) );
  XOR2_X1 U23482 ( .A1(n35218), .A2(n4709), .Z(n12351) );
  INV_X2 U23483 ( .I(n14405), .ZN(n15651) );
  XOR2_X1 U23484 ( .A1(n28969), .A2(n12355), .Z(n12354) );
  XOR2_X1 U23485 ( .A1(n28850), .A2(n19950), .Z(n12355) );
  NAND2_X1 U23489 ( .A1(n24403), .A2(n20517), .ZN(n12367) );
  INV_X2 U23492 ( .I(n17198), .ZN(n19147) );
  XOR2_X1 U23496 ( .A1(n27792), .A2(n27511), .Z(n27569) );
  INV_X2 U23502 ( .I(n12403), .ZN(n21898) );
  XNOR2_X1 U23503 ( .A1(Plaintext[13]), .A2(Key[13]), .ZN(n12403) );
  NOR2_X1 U23504 ( .A1(n13142), .A2(n3462), .ZN(n13141) );
  INV_X2 U23506 ( .I(n12414), .ZN(n29241) );
  XOR2_X1 U23507 ( .A1(n12556), .A2(n1169), .Z(n27000) );
  XOR2_X1 U23509 ( .A1(n29260), .A2(n19804), .Z(n13287) );
  XOR2_X1 U23511 ( .A1(n25263), .A2(n19897), .Z(n12438) );
  XOR2_X1 U23515 ( .A1(n35188), .A2(n29522), .Z(n27618) );
  NAND3_X1 U23518 ( .A1(n14433), .A2(n20901), .A3(n12450), .ZN(n14850) );
  XOR2_X1 U23520 ( .A1(n12454), .A2(n28549), .Z(n12453) );
  XOR2_X1 U23521 ( .A1(n35262), .A2(n38160), .Z(n12454) );
  XOR2_X1 U23526 ( .A1(n12470), .A2(n12468), .Z(n14076) );
  XOR2_X1 U23527 ( .A1(n28589), .A2(n12469), .Z(n12468) );
  XOR2_X1 U23528 ( .A1(n19513), .A2(n28889), .Z(n28589) );
  XOR2_X1 U23530 ( .A1(n29092), .A2(n19751), .Z(n12469) );
  XOR2_X1 U23531 ( .A1(n14388), .A2(n29114), .Z(n12470) );
  XOR2_X1 U23532 ( .A1(n28865), .A2(n31396), .Z(n29114) );
  NAND2_X2 U23533 ( .A1(n19482), .A2(n28488), .ZN(n29115) );
  XOR2_X1 U23542 ( .A1(n12493), .A2(n12492), .Z(n12491) );
  XOR2_X1 U23543 ( .A1(n27631), .A2(n19681), .Z(n12492) );
  XOR2_X1 U23544 ( .A1(n27541), .A2(n20976), .Z(n12493) );
  NOR2_X1 U23545 ( .A1(n28271), .A2(n11628), .ZN(n12498) );
  NAND3_X1 U23546 ( .A1(n19290), .A2(n28271), .A3(n28272), .ZN(n12499) );
  NOR2_X1 U23551 ( .A1(n24603), .A2(n36058), .ZN(n18055) );
  XOR2_X1 U23552 ( .A1(n27302), .A2(n12507), .Z(n18847) );
  XOR2_X1 U23553 ( .A1(n23695), .A2(n14289), .Z(n23786) );
  XOR2_X1 U23557 ( .A1(n12516), .A2(n14309), .Z(n12515) );
  INV_X2 U23558 ( .I(n18933), .ZN(n19332) );
  NAND2_X1 U23563 ( .A1(n25957), .A2(n18406), .ZN(n12525) );
  INV_X2 U23564 ( .I(n12535), .ZN(n13997) );
  XOR2_X1 U23565 ( .A1(n29252), .A2(n29253), .Z(n14171) );
  XOR2_X1 U23568 ( .A1(n37101), .A2(n19894), .Z(n27193) );
  XOR2_X1 U23570 ( .A1(n18160), .A2(n29528), .Z(n12553) );
  NOR2_X1 U23574 ( .A1(n32580), .A2(n5519), .ZN(n12558) );
  XOR2_X1 U23579 ( .A1(n12562), .A2(n12561), .Z(n12560) );
  XOR2_X1 U23580 ( .A1(n28866), .A2(n16685), .Z(n12563) );
  XOR2_X1 U23584 ( .A1(n29292), .A2(n12576), .Z(n12575) );
  XOR2_X1 U23585 ( .A1(n16356), .A2(n19741), .Z(n29049) );
  XOR2_X1 U23586 ( .A1(n4341), .A2(n29832), .Z(n12576) );
  XOR2_X1 U23588 ( .A1(n26286), .A2(n12587), .Z(n12586) );
  XOR2_X1 U23589 ( .A1(n11298), .A2(n18180), .Z(n12588) );
  XOR2_X1 U23593 ( .A1(n12593), .A2(n25034), .Z(n12592) );
  XOR2_X1 U23594 ( .A1(n37943), .A2(n25160), .Z(n12593) );
  XOR2_X1 U23596 ( .A1(n14214), .A2(n25033), .Z(n12594) );
  NAND2_X1 U23597 ( .A1(n37105), .A2(n24912), .ZN(n13610) );
  NAND2_X1 U23598 ( .A1(n36634), .A2(n32825), .ZN(n12654) );
  XOR2_X1 U23601 ( .A1(n18568), .A2(n22511), .Z(n22435) );
  XOR2_X1 U23605 ( .A1(n12622), .A2(n16381), .Z(n16382) );
  INV_X2 U23606 ( .I(n17313), .ZN(n28236) );
  INV_X2 U23607 ( .I(n20945), .ZN(n29815) );
  NAND2_X1 U23608 ( .A1(n21397), .A2(n19483), .ZN(n13682) );
  NAND2_X1 U23609 ( .A1(n19327), .A2(n12644), .ZN(n28011) );
  XOR2_X1 U23611 ( .A1(n26197), .A2(n12655), .Z(n20501) );
  XOR2_X1 U23612 ( .A1(n29562), .A2(n12839), .Z(n12655) );
  XOR2_X1 U23613 ( .A1(n5848), .A2(n29875), .Z(n26314) );
  XOR2_X1 U23614 ( .A1(n14307), .A2(n29298), .Z(n29299) );
  XOR2_X1 U23615 ( .A1(n33452), .A2(n19894), .Z(n12664) );
  XOR2_X1 U23617 ( .A1(n6131), .A2(n19649), .Z(n26228) );
  XOR2_X1 U23618 ( .A1(n6131), .A2(n36544), .Z(n12728) );
  XOR2_X1 U23622 ( .A1(n33041), .A2(n30085), .Z(n28928) );
  XOR2_X1 U23625 ( .A1(n16376), .A2(n26594), .Z(n12683) );
  XOR2_X1 U23626 ( .A1(Plaintext[159]), .A2(Key[159]), .Z(n12722) );
  OR2_X1 U23629 ( .A1(n20852), .A2(n20851), .Z(n12689) );
  XOR2_X1 U23630 ( .A1(n12570), .A2(n16697), .Z(n16696) );
  NOR2_X1 U23631 ( .A1(n13849), .A2(n34010), .ZN(n12703) );
  AOI21_X2 U23633 ( .A1(n34459), .A2(n975), .B(n12715), .ZN(n28799) );
  XOR2_X1 U23634 ( .A1(n18601), .A2(n1718), .Z(n29324) );
  INV_X2 U23635 ( .I(n12722), .ZN(n12754) );
  OAI21_X1 U23636 ( .A1(n19601), .A2(n27882), .B(n19467), .ZN(n12723) );
  XOR2_X1 U23639 ( .A1(n12728), .A2(n12727), .Z(n13183) );
  XOR2_X1 U23640 ( .A1(n5031), .A2(n1730), .Z(n12727) );
  XOR2_X1 U23642 ( .A1(n12730), .A2(n1697), .Z(n12862) );
  XOR2_X1 U23643 ( .A1(n12730), .A2(n22762), .Z(n16690) );
  INV_X2 U23644 ( .I(n12732), .ZN(n29591) );
  XOR2_X1 U23645 ( .A1(n12903), .A2(n26281), .Z(n12736) );
  XOR2_X1 U23646 ( .A1(n12741), .A2(n1738), .Z(n28826) );
  XOR2_X1 U23657 ( .A1(n22757), .A2(n16061), .Z(n12762) );
  NAND2_X1 U23660 ( .A1(n15332), .A2(n3120), .ZN(n15333) );
  OAI21_X1 U23661 ( .A1(n33344), .A2(n24847), .B(n3120), .ZN(n24540) );
  XOR2_X1 U23663 ( .A1(n27758), .A2(n30179), .Z(n12769) );
  INV_X2 U23664 ( .I(n12770), .ZN(n21132) );
  XOR2_X1 U23672 ( .A1(n39025), .A2(n29649), .Z(n12796) );
  OAI21_X2 U23673 ( .A1(n39467), .A2(n19880), .B(n24395), .ZN(n12804) );
  AOI21_X2 U23677 ( .A1(n25834), .A2(n39291), .B(n25833), .ZN(n26253) );
  MUX2_X1 U23679 ( .I0(n19581), .I1(n31580), .S(n12828), .Z(n12826) );
  XOR2_X1 U23682 ( .A1(n25003), .A2(n25004), .Z(n12833) );
  XOR2_X1 U23683 ( .A1(n12835), .A2(n12834), .Z(n12836) );
  XOR2_X1 U23684 ( .A1(n7055), .A2(n32174), .Z(n22697) );
  XOR2_X1 U23687 ( .A1(n12847), .A2(n1734), .Z(Ciphertext[29]) );
  NAND2_X1 U23688 ( .A1(n20566), .A2(n29241), .ZN(n29287) );
  XOR2_X1 U23689 ( .A1(n20976), .A2(n900), .Z(n12854) );
  XOR2_X1 U23691 ( .A1(n14230), .A2(n666), .Z(n12858) );
  XOR2_X1 U23693 ( .A1(n18446), .A2(n12862), .Z(n12861) );
  XOR2_X1 U23695 ( .A1(n25285), .A2(n16843), .Z(n12871) );
  NAND3_X1 U23701 ( .A1(n12885), .A2(n28352), .A3(n28351), .ZN(n28353) );
  NAND2_X1 U23702 ( .A1(n28535), .A2(n28495), .ZN(n12888) );
  XOR2_X1 U23705 ( .A1(n20412), .A2(n12897), .Z(n12899) );
  XOR2_X1 U23706 ( .A1(n17195), .A2(n22580), .Z(n12897) );
  XOR2_X1 U23707 ( .A1(n12898), .A2(n12899), .Z(n12900) );
  XOR2_X1 U23711 ( .A1(n22511), .A2(n18296), .Z(n12901) );
  XOR2_X1 U23712 ( .A1(n12902), .A2(Plaintext[23]), .Z(n21441) );
  INV_X1 U23713 ( .I(Key[23]), .ZN(n12902) );
  XOR2_X1 U23717 ( .A1(n39172), .A2(n12915), .Z(n17946) );
  XOR2_X1 U23718 ( .A1(n2782), .A2(n12939), .Z(n12918) );
  XOR2_X1 U23719 ( .A1(n14756), .A2(n17817), .Z(n12919) );
  XOR2_X1 U23720 ( .A1(n12922), .A2(n790), .Z(n12920) );
  XOR2_X1 U23722 ( .A1(n23912), .A2(n23667), .Z(n12922) );
  XOR2_X1 U23724 ( .A1(n24944), .A2(n24984), .Z(n25029) );
  NAND2_X1 U23725 ( .A1(n12926), .A2(n370), .ZN(n24481) );
  NOR2_X1 U23733 ( .A1(n9839), .A2(n29367), .ZN(n19059) );
  NOR2_X1 U23736 ( .A1(n35023), .A2(n28695), .ZN(n17320) );
  NAND2_X1 U23738 ( .A1(n12950), .A2(n12951), .ZN(n24273) );
  OAI21_X2 U23742 ( .A1(n17724), .A2(n16660), .B(n16659), .ZN(n17685) );
  XOR2_X1 U23746 ( .A1(n23812), .A2(n23220), .Z(n12976) );
  NAND2_X1 U23750 ( .A1(n38953), .A2(n16250), .ZN(n12984) );
  XOR2_X1 U23751 ( .A1(n29045), .A2(n29730), .Z(n12985) );
  XOR2_X1 U23752 ( .A1(n29289), .A2(n12989), .Z(n29290) );
  XOR2_X1 U23754 ( .A1(n24932), .A2(n25006), .Z(n25234) );
  OAI22_X2 U23755 ( .A1(n24726), .A2(n24725), .B1(n24724), .B2(n9656), .ZN(
        n25006) );
  NAND2_X2 U23756 ( .A1(n24415), .A2(n24414), .ZN(n24932) );
  NAND2_X1 U23759 ( .A1(n30171), .A2(n17997), .ZN(n13006) );
  XOR2_X1 U23760 ( .A1(n22485), .A2(n19925), .Z(n13255) );
  NOR2_X1 U23761 ( .A1(n13300), .A2(n24515), .ZN(n24292) );
  XNOR2_X1 U23764 ( .A1(n25303), .A2(n18991), .ZN(n25329) );
  XOR2_X1 U23765 ( .A1(n25330), .A2(n25331), .Z(n13013) );
  NAND2_X1 U23766 ( .A1(n21892), .A2(n12670), .ZN(n19376) );
  XOR2_X1 U23767 ( .A1(n13024), .A2(n13022), .Z(n14122) );
  XOR2_X1 U23768 ( .A1(n23741), .A2(n13023), .Z(n13022) );
  XOR2_X1 U23769 ( .A1(n23972), .A2(n13025), .Z(n13024) );
  INV_X1 U23774 ( .I(n20342), .ZN(n30181) );
  NOR2_X1 U23777 ( .A1(n35506), .A2(n13038), .ZN(n19924) );
  XOR2_X1 U23782 ( .A1(n13054), .A2(n30094), .Z(n16161) );
  XOR2_X1 U23784 ( .A1(n39063), .A2(n26365), .Z(n26398) );
  INV_X2 U23793 ( .I(n13082), .ZN(n17410) );
  XOR2_X1 U23794 ( .A1(n27636), .A2(n27639), .Z(n13083) );
  XOR2_X1 U23806 ( .A1(n23831), .A2(n1726), .Z(n13101) );
  AND2_X1 U23807 ( .A1(n25826), .A2(n25825), .Z(n13103) );
  INV_X2 U23813 ( .I(n13124), .ZN(n15290) );
  INV_X2 U23815 ( .I(n13127), .ZN(n14962) );
  NAND3_X1 U23816 ( .A1(n25630), .A2(n13129), .A3(n911), .ZN(n25369) );
  INV_X1 U23820 ( .I(n13132), .ZN(n29906) );
  XOR2_X1 U23821 ( .A1(n37943), .A2(n14374), .Z(n25231) );
  XOR2_X1 U23822 ( .A1(n35953), .A2(n14374), .Z(n25091) );
  XOR2_X1 U23824 ( .A1(n25193), .A2(n14374), .Z(n17553) );
  XOR2_X1 U23826 ( .A1(n18543), .A2(n18546), .Z(n13138) );
  XOR2_X1 U23827 ( .A1(n5021), .A2(n19720), .Z(n16093) );
  XOR2_X1 U23828 ( .A1(n29024), .A2(n13139), .Z(n14835) );
  XOR2_X1 U23829 ( .A1(n19887), .A2(n29824), .Z(n13139) );
  XOR2_X1 U23830 ( .A1(n13140), .A2(n16498), .Z(Ciphertext[1]) );
  NAND2_X1 U23835 ( .A1(n13153), .A2(n37060), .ZN(n13657) );
  NAND2_X1 U23836 ( .A1(n13158), .A2(n13998), .ZN(n13557) );
  NAND2_X1 U23837 ( .A1(n13170), .A2(n31542), .ZN(n14222) );
  XOR2_X1 U23839 ( .A1(n22661), .A2(n22660), .Z(n13172) );
  XOR2_X1 U23841 ( .A1(n13716), .A2(n13183), .Z(n26968) );
  XOR2_X1 U23842 ( .A1(n13188), .A2(n15835), .Z(n13187) );
  XOR2_X1 U23843 ( .A1(n29040), .A2(n30964), .Z(n13188) );
  XOR2_X1 U23846 ( .A1(n24417), .A2(n25133), .Z(n13190) );
  XOR2_X1 U23848 ( .A1(n22710), .A2(n36513), .Z(n13199) );
  NAND2_X1 U23852 ( .A1(n29763), .A2(n13208), .ZN(n28963) );
  AND2_X1 U23853 ( .A1(n13207), .A2(n28961), .Z(n13208) );
  NOR2_X1 U23855 ( .A1(n7676), .A2(n7973), .ZN(n13212) );
  XOR2_X1 U23857 ( .A1(n18279), .A2(n30068), .Z(n13215) );
  NOR2_X1 U23862 ( .A1(n22368), .A2(n13995), .ZN(n13226) );
  XOR2_X1 U23864 ( .A1(n26274), .A2(n39172), .Z(n13232) );
  XOR2_X1 U23866 ( .A1(n29024), .A2(n29823), .Z(n21079) );
  XOR2_X1 U23869 ( .A1(n26389), .A2(n19755), .Z(n13242) );
  XOR2_X1 U23870 ( .A1(n26437), .A2(n26567), .Z(n13243) );
  XOR2_X1 U23871 ( .A1(n31599), .A2(n7944), .Z(n13247) );
  OR2_X1 U23872 ( .A1(n29673), .A2(n18042), .Z(n18795) );
  INV_X2 U23873 ( .I(n19948), .ZN(n29764) );
  XOR2_X1 U23875 ( .A1(n13255), .A2(n7432), .Z(n13254) );
  NAND2_X2 U23878 ( .A1(n19268), .A2(n21967), .ZN(n22621) );
  XOR2_X1 U23881 ( .A1(Plaintext[77]), .A2(Key[77]), .Z(n17833) );
  NAND2_X2 U23882 ( .A1(n29403), .A2(n29400), .ZN(n29410) );
  XOR2_X1 U23884 ( .A1(n33509), .A2(n29522), .Z(n17243) );
  INV_X1 U23887 ( .I(n13278), .ZN(n20708) );
  XOR2_X1 U23888 ( .A1(n13283), .A2(n27658), .Z(n27659) );
  INV_X2 U23892 ( .I(n13286), .ZN(n13545) );
  INV_X1 U23895 ( .I(n13292), .ZN(n13291) );
  XOR2_X1 U23896 ( .A1(n22595), .A2(n28934), .Z(n13295) );
  OR2_X1 U23897 ( .A1(n29493), .A2(n15621), .Z(n13302) );
  NOR2_X1 U23898 ( .A1(n13959), .A2(n13997), .ZN(n13556) );
  AOI21_X2 U23903 ( .A1(n24278), .A2(n13310), .B(n24277), .ZN(n24515) );
  XOR2_X1 U23904 ( .A1(n13315), .A2(n13312), .Z(n13317) );
  XOR2_X1 U23906 ( .A1(n9035), .A2(n19800), .Z(n13313) );
  INV_X2 U23908 ( .I(n13317), .ZN(n29493) );
  NOR3_X1 U23909 ( .A1(n21397), .A2(n13318), .A3(n13997), .ZN(n13684) );
  NOR2_X1 U23910 ( .A1(n695), .A2(n18959), .ZN(n13318) );
  XOR2_X1 U23913 ( .A1(n25247), .A2(n20479), .Z(n13326) );
  XOR2_X1 U23917 ( .A1(n8894), .A2(n27735), .Z(n27547) );
  XOR2_X1 U23918 ( .A1(n13329), .A2(n19929), .Z(Ciphertext[38]) );
  INV_X2 U23921 ( .I(n13332), .ZN(n28283) );
  XOR2_X1 U23922 ( .A1(n31579), .A2(n19786), .Z(n15405) );
  MUX2_X1 U23924 ( .I0(n19737), .I1(n18656), .S(n22228), .Z(n22027) );
  XOR2_X1 U23932 ( .A1(n22651), .A2(n22652), .Z(n13356) );
  XOR2_X1 U23934 ( .A1(n29123), .A2(n14244), .Z(n13358) );
  XNOR2_X1 U23937 ( .A1(Plaintext[54]), .A2(Key[54]), .ZN(n13359) );
  INV_X2 U23939 ( .I(n22837), .ZN(n23101) );
  XOR2_X1 U23940 ( .A1(n13362), .A2(n13361), .Z(n22837) );
  XOR2_X1 U23941 ( .A1(n17988), .A2(n14894), .Z(n13361) );
  XOR2_X1 U23942 ( .A1(n22774), .A2(n22662), .Z(n13362) );
  XOR2_X1 U23943 ( .A1(n23971), .A2(n13368), .Z(n13367) );
  XOR2_X1 U23944 ( .A1(n24049), .A2(n19937), .Z(n13368) );
  XOR2_X1 U23945 ( .A1(n26573), .A2(n29334), .Z(n26575) );
  AND2_X1 U23946 ( .A1(n28466), .A2(n13372), .Z(n16840) );
  XOR2_X1 U23953 ( .A1(n13544), .A2(n26294), .Z(n13543) );
  INV_X2 U23954 ( .I(n13397), .ZN(n21912) );
  XOR2_X1 U23957 ( .A1(n16651), .A2(n33990), .Z(n16650) );
  OAI21_X1 U23959 ( .A1(n19007), .A2(n13412), .B(n1032), .ZN(n17301) );
  INV_X2 U23960 ( .I(n13413), .ZN(n18909) );
  NAND2_X1 U23961 ( .A1(n13415), .A2(n1121), .ZN(n24413) );
  MUX2_X1 U23964 ( .I0(n16853), .I1(n35224), .S(n14193), .Z(n13424) );
  INV_X1 U23965 ( .I(n26177), .ZN(n26703) );
  INV_X2 U23966 ( .I(n13425), .ZN(n19951) );
  INV_X2 U23968 ( .I(n13429), .ZN(n17693) );
  XOR2_X1 U23969 ( .A1(n14303), .A2(n22611), .Z(n13430) );
  AOI21_X1 U23970 ( .A1(n20964), .A2(n34534), .B(n13433), .ZN(n13432) );
  INV_X1 U23971 ( .I(n17594), .ZN(n25575) );
  XOR2_X1 U23972 ( .A1(n13439), .A2(n23880), .Z(n23660) );
  XOR2_X1 U23975 ( .A1(n27864), .A2(n29476), .Z(n13448) );
  AND2_X1 U23976 ( .A1(n1645), .A2(n19351), .Z(n13451) );
  INV_X2 U23977 ( .I(n14332), .ZN(n25539) );
  XOR2_X1 U23978 ( .A1(Plaintext[69]), .A2(Key[69]), .Z(n13473) );
  XOR2_X1 U23979 ( .A1(n13477), .A2(n13475), .Z(n21291) );
  XOR2_X1 U23980 ( .A1(n13476), .A2(n22565), .Z(n13475) );
  XOR2_X1 U23981 ( .A1(n19254), .A2(n22732), .Z(n13476) );
  XOR2_X1 U23983 ( .A1(n13479), .A2(n11541), .Z(n13478) );
  XOR2_X1 U23984 ( .A1(n17605), .A2(n19720), .Z(n13479) );
  XOR2_X1 U23991 ( .A1(n31504), .A2(n29320), .Z(n22200) );
  INV_X2 U23997 ( .I(n13503), .ZN(n24445) );
  XOR2_X1 U24000 ( .A1(n27782), .A2(n13510), .Z(n13969) );
  XOR2_X1 U24001 ( .A1(n27781), .A2(n19749), .Z(n13510) );
  NAND2_X2 U24003 ( .A1(n13523), .A2(n13525), .ZN(n17757) );
  NAND3_X1 U24008 ( .A1(n1340), .A2(n4200), .A3(n13519), .ZN(n21334) );
  NOR2_X1 U24013 ( .A1(n8304), .A2(n1551), .ZN(n19302) );
  XOR2_X1 U24014 ( .A1(n29104), .A2(n29306), .Z(n28869) );
  AND2_X1 U24022 ( .A1(n25717), .A2(n25716), .Z(n13538) );
  MUX2_X1 U24023 ( .I0(n28141), .I1(n20184), .S(n281), .Z(n13539) );
  XOR2_X1 U24025 ( .A1(n23996), .A2(n38813), .Z(n23684) );
  XOR2_X1 U24031 ( .A1(n28574), .A2(n13552), .Z(n13551) );
  XOR2_X1 U24032 ( .A1(n29837), .A2(n19613), .Z(n13552) );
  OAI21_X1 U24036 ( .A1(n16472), .A2(n13559), .B(n13558), .ZN(n16469) );
  AOI22_X1 U24037 ( .A1(n16471), .A2(n30093), .B1(n16470), .B2(n13559), .ZN(
        n13558) );
  INV_X2 U24039 ( .I(n13561), .ZN(n23020) );
  XOR2_X1 U24042 ( .A1(n22659), .A2(n15909), .Z(n20865) );
  INV_X1 U24043 ( .I(n22347), .ZN(n13566) );
  XOR2_X1 U24044 ( .A1(n13569), .A2(n19817), .Z(n27513) );
  XOR2_X1 U24053 ( .A1(n15216), .A2(n28912), .Z(n17905) );
  XOR2_X1 U24057 ( .A1(n13592), .A2(n22559), .Z(n13591) );
  XOR2_X1 U24058 ( .A1(n22773), .A2(n29661), .Z(n13592) );
  INV_X2 U24063 ( .I(n13595), .ZN(n28036) );
  XOR2_X1 U24065 ( .A1(n23830), .A2(n18828), .Z(n17581) );
  NAND2_X1 U24076 ( .A1(n16065), .A2(n19855), .ZN(n13623) );
  XOR2_X1 U24080 ( .A1(n13634), .A2(n29399), .Z(n24936) );
  XOR2_X1 U24085 ( .A1(n23688), .A2(n23465), .Z(n13649) );
  XOR2_X1 U24087 ( .A1(n21332), .A2(Key[102]), .Z(n19387) );
  XOR2_X1 U24089 ( .A1(n35824), .A2(n2383), .Z(n22520) );
  XOR2_X1 U24093 ( .A1(n13658), .A2(n19492), .Z(n18135) );
  XOR2_X1 U24095 ( .A1(n17565), .A2(n13667), .Z(n13668) );
  INV_X2 U24096 ( .I(n13668), .ZN(n14442) );
  NOR2_X1 U24097 ( .A1(n19704), .A2(n33368), .ZN(n13672) );
  XOR2_X1 U24098 ( .A1(n17757), .A2(n12649), .Z(n13674) );
  XOR2_X1 U24100 ( .A1(Plaintext[72]), .A2(Key[72]), .Z(n13679) );
  XOR2_X1 U24101 ( .A1(n705), .A2(n5203), .Z(n13680) );
  XOR2_X1 U24102 ( .A1(n22700), .A2(n14022), .Z(n13681) );
  NAND2_X2 U24103 ( .A1(n13683), .A2(n13682), .ZN(n22315) );
  XOR2_X1 U24104 ( .A1(n25137), .A2(n13689), .Z(n25138) );
  XOR2_X1 U24105 ( .A1(n1258), .A2(n16864), .Z(n13689) );
  NAND2_X1 U24112 ( .A1(n26856), .A2(n11334), .ZN(n13698) );
  NAND2_X1 U24115 ( .A1(n1641), .A2(n35689), .ZN(n23617) );
  XOR2_X1 U24116 ( .A1(n386), .A2(n1718), .Z(n16709) );
  XOR2_X1 U24118 ( .A1(n35505), .A2(n16226), .Z(n22664) );
  NOR2_X1 U24121 ( .A1(n24309), .A2(n807), .ZN(n13710) );
  XOR2_X1 U24126 ( .A1(n26364), .A2(n26482), .Z(n13716) );
  INV_X2 U24128 ( .I(n13725), .ZN(n15153) );
  XOR2_X1 U24129 ( .A1(n23756), .A2(n16244), .Z(n13729) );
  INV_X2 U24131 ( .I(n16993), .ZN(n21484) );
  XOR2_X1 U24132 ( .A1(Plaintext[86]), .A2(Key[86]), .Z(n16993) );
  INV_X2 U24134 ( .I(n13745), .ZN(n23107) );
  XOR2_X1 U24135 ( .A1(n13750), .A2(n27521), .Z(n13749) );
  NAND2_X1 U24136 ( .A1(n13786), .A2(n30262), .ZN(n13990) );
  NOR2_X1 U24137 ( .A1(n13753), .A2(n35114), .ZN(n27331) );
  NOR2_X1 U24139 ( .A1(n11039), .A2(n13753), .ZN(n27332) );
  INV_X2 U24141 ( .I(n13759), .ZN(n26839) );
  NAND2_X2 U24148 ( .A1(n13789), .A2(n13788), .ZN(n19515) );
  XOR2_X1 U24151 ( .A1(n29245), .A2(n29244), .Z(n13797) );
  NOR2_X1 U24153 ( .A1(n26137), .A2(n13801), .ZN(n15684) );
  XOR2_X1 U24154 ( .A1(n13802), .A2(n19879), .Z(n27087) );
  XOR2_X1 U24155 ( .A1(n27679), .A2(n13802), .Z(n27042) );
  INV_X2 U24156 ( .I(n13827), .ZN(n19863) );
  AND2_X1 U24162 ( .A1(n13834), .A2(n13833), .Z(n13832) );
  XOR2_X1 U24165 ( .A1(n22608), .A2(n13846), .Z(n13845) );
  INV_X2 U24167 ( .I(n13862), .ZN(n14404) );
  XOR2_X1 U24175 ( .A1(n900), .A2(n19761), .Z(n13878) );
  OAI21_X1 U24176 ( .A1(n16778), .A2(n33843), .B(n13879), .ZN(n14931) );
  OR2_X1 U24179 ( .A1(n37157), .A2(n19085), .Z(n13886) );
  NOR2_X1 U24182 ( .A1(n11413), .A2(n8944), .ZN(n13892) );
  MUX2_X1 U24185 ( .I0(n27876), .I1(n28200), .S(n18061), .Z(n13907) );
  XOR2_X1 U24189 ( .A1(n20352), .A2(n9626), .Z(n22533) );
  XOR2_X1 U24197 ( .A1(n34178), .A2(n29300), .Z(n13933) );
  XOR2_X1 U24199 ( .A1(n21108), .A2(n29110), .Z(n13934) );
  XOR2_X1 U24200 ( .A1(n14639), .A2(n16417), .Z(n13937) );
  XOR2_X1 U24201 ( .A1(n25277), .A2(n33661), .Z(n13939) );
  OAI21_X1 U24203 ( .A1(n14409), .A2(n33925), .B(n13945), .ZN(n23206) );
  XOR2_X1 U24209 ( .A1(n39765), .A2(n17646), .Z(n13967) );
  NOR2_X1 U24212 ( .A1(n28231), .A2(n18451), .ZN(n13983) );
  INV_X2 U24216 ( .I(n14000), .ZN(n19762) );
  NAND3_X1 U24218 ( .A1(n14006), .A2(n22817), .A3(n6646), .ZN(n22819) );
  OAI21_X1 U24219 ( .A1(n29810), .A2(n966), .B(n15189), .ZN(n14008) );
  INV_X2 U24221 ( .I(n14016), .ZN(n19395) );
  XNOR2_X1 U24222 ( .A1(Plaintext[108]), .A2(Key[108]), .ZN(n14016) );
  XOR2_X1 U24225 ( .A1(n22515), .A2(n30120), .Z(n14022) );
  XOR2_X1 U24228 ( .A1(n20723), .A2(n18539), .Z(n14031) );
  XOR2_X1 U24230 ( .A1(n12839), .A2(n26476), .Z(n14143) );
  NOR3_X1 U24231 ( .A1(n2839), .A2(n14027), .A3(n36428), .ZN(n14034) );
  NOR2_X1 U24232 ( .A1(n17664), .A2(n2839), .ZN(n14035) );
  XOR2_X1 U24233 ( .A1(n25264), .A2(n719), .Z(n14043) );
  XOR2_X1 U24234 ( .A1(n17837), .A2(n24966), .Z(n14046) );
  NAND2_X1 U24237 ( .A1(n34074), .A2(n37377), .ZN(n14050) );
  XOR2_X1 U24241 ( .A1(n7942), .A2(n14063), .Z(n14062) );
  XOR2_X1 U24242 ( .A1(n22741), .A2(n31863), .Z(n14063) );
  XOR2_X1 U24244 ( .A1(n26590), .A2(n29689), .Z(n14069) );
  XOR2_X1 U24250 ( .A1(n14128), .A2(n31547), .Z(n14099) );
  XOR2_X1 U24252 ( .A1(n23676), .A2(n14105), .Z(n14104) );
  XOR2_X1 U24253 ( .A1(n23890), .A2(n19681), .Z(n14105) );
  INV_X1 U24256 ( .I(n22603), .ZN(n19118) );
  XOR2_X1 U24258 ( .A1(n35824), .A2(n28831), .Z(n14112) );
  XOR2_X1 U24259 ( .A1(n22787), .A2(n22447), .Z(n14113) );
  XOR2_X1 U24270 ( .A1(n27567), .A2(n27568), .Z(n14147) );
  XOR2_X1 U24271 ( .A1(n33252), .A2(n30065), .Z(n14148) );
  AOI21_X2 U24273 ( .A1(n29496), .A2(n14151), .B(n14150), .ZN(n20208) );
  OR2_X1 U24275 ( .A1(n37227), .A2(n17693), .Z(n14154) );
  XOR2_X1 U24279 ( .A1(n5208), .A2(n31543), .Z(n24542) );
  XOR2_X1 U24281 ( .A1(Plaintext[88]), .A2(Key[88]), .Z(n21882) );
  XOR2_X1 U24284 ( .A1(n22668), .A2(n22563), .Z(n21994) );
  NAND2_X2 U24286 ( .A1(n23800), .A2(n14169), .ZN(n24821) );
  XOR2_X1 U24287 ( .A1(n31566), .A2(n19851), .Z(n14173) );
  INV_X1 U24288 ( .I(n28290), .ZN(n28155) );
  XOR2_X1 U24291 ( .A1(n9116), .A2(n33990), .Z(n22698) );
  XOR2_X1 U24296 ( .A1(n22647), .A2(n22772), .Z(n14194) );
  NAND2_X2 U24297 ( .A1(n20487), .A2(n27572), .ZN(n15745) );
  AOI21_X1 U24298 ( .A1(n17973), .A2(n17972), .B(n14196), .ZN(n20670) );
  XOR2_X1 U24302 ( .A1(n37499), .A2(n38212), .Z(n18579) );
  NAND2_X1 U24303 ( .A1(n25971), .A2(n35151), .ZN(n14215) );
  XOR2_X1 U24305 ( .A1(n36218), .A2(n19755), .Z(n24524) );
  XOR2_X1 U24306 ( .A1(n36218), .A2(n24982), .Z(n24861) );
  NAND2_X2 U24307 ( .A1(n15038), .A2(n14426), .ZN(n14232) );
  XOR2_X1 U24310 ( .A1(n31522), .A2(n20658), .Z(n14244) );
  XNOR2_X1 U24312 ( .A1(Plaintext[49]), .A2(Key[49]), .ZN(n14245) );
  OAI21_X2 U24316 ( .A1(n14252), .A2(n14251), .B(n14248), .ZN(n22594) );
  XNOR2_X1 U24321 ( .A1(n24065), .A2(n23905), .ZN(n16781) );
  NOR2_X1 U24326 ( .A1(n19193), .A2(n17238), .ZN(n14282) );
  XOR2_X1 U24328 ( .A1(Key[127]), .A2(Plaintext[127]), .Z(n19871) );
  INV_X2 U24329 ( .I(n14287), .ZN(n19594) );
  XOR2_X1 U24331 ( .A1(n33252), .A2(n19904), .Z(n14293) );
  XOR2_X1 U24332 ( .A1(n22771), .A2(n14295), .Z(n14294) );
  XOR2_X1 U24333 ( .A1(n22528), .A2(n11308), .Z(n14295) );
  XOR2_X1 U24336 ( .A1(n26457), .A2(n837), .Z(n14302) );
  XOR2_X1 U24337 ( .A1(n14304), .A2(n14309), .Z(n14303) );
  XOR2_X1 U24339 ( .A1(n14307), .A2(n15203), .Z(n16583) );
  XOR2_X1 U24343 ( .A1(n33038), .A2(n29849), .Z(n19131) );
  XOR2_X1 U24350 ( .A1(n1458), .A2(n27556), .Z(n27573) );
  XOR2_X1 U24351 ( .A1(n27461), .A2(n14325), .Z(n27462) );
  INV_X1 U24354 ( .I(Plaintext[71]), .ZN(n14333) );
  MUX2_X1 U24357 ( .I0(n28006), .I1(n28007), .S(n941), .Z(n28010) );
  OAI22_X2 U24358 ( .A1(n22878), .A2(n14343), .B1(n22877), .B2(n23121), .ZN(
        n23461) );
  XOR2_X1 U24365 ( .A1(n39637), .A2(n29647), .Z(n26344) );
  XOR2_X1 U24369 ( .A1(n18300), .A2(n23675), .Z(n23741) );
  OAI21_X2 U24370 ( .A1(n14363), .A2(n19292), .B(n21803), .ZN(n22773) );
  XOR2_X1 U24371 ( .A1(n6435), .A2(n32174), .Z(n14364) );
  NOR2_X1 U24373 ( .A1(n25048), .A2(n24912), .ZN(n15633) );
  AOI21_X1 U24375 ( .A1(n23311), .A2(n39626), .B(n19869), .ZN(n23015) );
  NOR2_X1 U24386 ( .A1(n28675), .A2(n28676), .ZN(n15631) );
  NOR2_X1 U24390 ( .A1(n14450), .A2(n1354), .ZN(n17724) );
  NAND2_X1 U24393 ( .A1(n19594), .A2(n20590), .ZN(n19361) );
  INV_X1 U24394 ( .I(n27862), .ZN(n20310) );
  NAND2_X1 U24395 ( .A1(n17942), .A2(n17551), .ZN(n16534) );
  NOR2_X1 U24397 ( .A1(n11307), .A2(n20782), .ZN(n23113) );
  NAND2_X1 U24406 ( .A1(n16159), .A2(n10477), .ZN(n16158) );
  NOR2_X1 U24408 ( .A1(n24854), .A2(n24853), .ZN(n18537) );
  NAND2_X1 U24414 ( .A1(n36954), .A2(n20010), .ZN(n19996) );
  NAND2_X1 U24415 ( .A1(n5020), .A2(n28282), .ZN(n28068) );
  NAND3_X1 U24418 ( .A1(n31604), .A2(n21672), .A3(n21667), .ZN(n14912) );
  NAND2_X1 U24419 ( .A1(n18266), .A2(n694), .ZN(n16763) );
  OAI21_X1 U24423 ( .A1(n21551), .A2(n11851), .B(n1690), .ZN(n20330) );
  NAND2_X1 U24430 ( .A1(n1678), .A2(n9685), .ZN(n16455) );
  INV_X1 U24433 ( .I(n20518), .ZN(n23063) );
  NAND2_X1 U24436 ( .A1(n22928), .A2(n22990), .ZN(n18377) );
  NOR2_X1 U24444 ( .A1(n17076), .A2(n24461), .ZN(n20002) );
  NAND3_X1 U24447 ( .A1(n1634), .A2(n23552), .A3(n14845), .ZN(n18915) );
  NAND2_X1 U24448 ( .A1(n6849), .A2(n24469), .ZN(n19053) );
  INV_X1 U24451 ( .I(n20394), .ZN(n24156) );
  NAND2_X1 U24459 ( .A1(n16999), .A2(n39317), .ZN(n19643) );
  INV_X1 U24460 ( .I(n37943), .ZN(n16350) );
  INV_X1 U24462 ( .I(n20627), .ZN(n25390) );
  INV_X1 U24463 ( .I(n25724), .ZN(n16317) );
  NAND2_X1 U24464 ( .A1(n15180), .A2(n37926), .ZN(n25399) );
  INV_X1 U24469 ( .I(n26163), .ZN(n19464) );
  NAND2_X1 U24474 ( .A1(n27321), .A2(n14881), .ZN(n18251) );
  INV_X1 U24477 ( .I(n16169), .ZN(n17051) );
  INV_X1 U24478 ( .I(n27606), .ZN(n27609) );
  NAND2_X1 U24479 ( .A1(n17686), .A2(n17699), .ZN(n15162) );
  NAND3_X1 U24480 ( .A1(n27449), .A2(n33893), .A3(n16043), .ZN(n15277) );
  INV_X1 U24481 ( .I(n27507), .ZN(n15246) );
  INV_X1 U24482 ( .I(n17349), .ZN(n20721) );
  NAND2_X1 U24484 ( .A1(n27989), .A2(n38996), .ZN(n18687) );
  NAND2_X1 U24489 ( .A1(n20053), .A2(n7591), .ZN(n19324) );
  NAND2_X1 U24490 ( .A1(n38874), .A2(n18948), .ZN(n19325) );
  NAND2_X1 U24493 ( .A1(n27984), .A2(n37204), .ZN(n19957) );
  NAND2_X1 U24494 ( .A1(n16777), .A2(n17542), .ZN(n17541) );
  INV_X1 U24495 ( .I(n7667), .ZN(n28931) );
  NAND2_X1 U24498 ( .A1(n21550), .A2(n21506), .ZN(n15149) );
  INV_X1 U24500 ( .I(n21753), .ZN(n21698) );
  NOR3_X1 U24502 ( .A1(n20535), .A2(n3562), .A3(n21870), .ZN(n15155) );
  NOR2_X1 U24506 ( .A1(n21862), .A2(n21823), .ZN(n15097) );
  OR2_X1 U24507 ( .A1(n19016), .A2(n21858), .Z(n15099) );
  INV_X1 U24508 ( .I(n21841), .ZN(n21903) );
  OAI21_X1 U24517 ( .A1(n37200), .A2(n1349), .B(n1990), .ZN(n19320) );
  NAND2_X1 U24520 ( .A1(n39680), .A2(n21488), .ZN(n19377) );
  NAND2_X1 U24521 ( .A1(n39680), .A2(n21568), .ZN(n14919) );
  NOR2_X1 U24522 ( .A1(n20799), .A2(n1333), .ZN(n18728) );
  NAND2_X1 U24523 ( .A1(n9942), .A2(n18152), .ZN(n21843) );
  NAND2_X1 U24524 ( .A1(n21890), .A2(n15910), .ZN(n18758) );
  NOR2_X1 U24525 ( .A1(n21784), .A2(n20241), .ZN(n21505) );
  NOR2_X1 U24527 ( .A1(n19850), .A2(n16333), .ZN(n21694) );
  NOR2_X1 U24529 ( .A1(n34282), .A2(n17989), .ZN(n20280) );
  NAND2_X1 U24530 ( .A1(n21593), .A2(n21484), .ZN(n21590) );
  OAI21_X1 U24534 ( .A1(n32525), .A2(n18028), .B(n1354), .ZN(n21935) );
  AOI21_X1 U24535 ( .A1(n20003), .A2(n20476), .B(n16537), .ZN(n16536) );
  OAI21_X1 U24539 ( .A1(n18412), .A2(n21917), .B(n19105), .ZN(n19104) );
  NAND2_X1 U24541 ( .A1(n21917), .A2(n34867), .ZN(n19105) );
  NOR2_X1 U24544 ( .A1(n9543), .A2(n23042), .ZN(n14851) );
  NOR2_X1 U24553 ( .A1(n22865), .A2(n12331), .ZN(n15239) );
  NOR2_X1 U24554 ( .A1(n18071), .A2(n18072), .ZN(n18506) );
  NAND2_X1 U24555 ( .A1(n33933), .A2(n23076), .ZN(n15039) );
  INV_X1 U24558 ( .I(n22934), .ZN(n22083) );
  NAND2_X1 U24559 ( .A1(n18850), .A2(n23308), .ZN(n23309) );
  INV_X1 U24568 ( .I(n23420), .ZN(n17224) );
  NAND2_X1 U24572 ( .A1(n22992), .A2(n22993), .ZN(n20024) );
  NAND2_X1 U24573 ( .A1(n16292), .A2(n16291), .ZN(n16150) );
  OAI21_X1 U24574 ( .A1(n23346), .A2(n1634), .B(n23550), .ZN(n18618) );
  INV_X1 U24575 ( .I(n24077), .ZN(n15477) );
  NAND2_X1 U24578 ( .A1(n24311), .A2(n19584), .ZN(n16918) );
  NAND3_X1 U24579 ( .A1(n9078), .A2(n20972), .A3(n4542), .ZN(n15534) );
  NAND2_X1 U24582 ( .A1(n32069), .A2(n39074), .ZN(n24153) );
  NAND2_X1 U24583 ( .A1(n24795), .A2(n16238), .ZN(n17453) );
  NOR2_X1 U24585 ( .A1(n24419), .A2(n30494), .ZN(n24090) );
  NAND2_X1 U24592 ( .A1(n24660), .A2(n18110), .ZN(n18263) );
  INV_X1 U24593 ( .I(n24784), .ZN(n24785) );
  OAI21_X1 U24596 ( .A1(n596), .A2(n26061), .B(n9530), .ZN(n25740) );
  NOR2_X1 U24601 ( .A1(n26185), .A2(n25934), .ZN(n26187) );
  INV_X1 U24603 ( .I(n26338), .ZN(n26418) );
  NAND2_X1 U24606 ( .A1(n9859), .A2(n25849), .ZN(n14839) );
  NOR2_X1 U24609 ( .A1(n25754), .A2(n25699), .ZN(n21233) );
  NOR2_X1 U24610 ( .A1(n24896), .A2(n25390), .ZN(n17091) );
  INV_X1 U24611 ( .I(n25418), .ZN(n25600) );
  NOR2_X1 U24614 ( .A1(n36249), .A2(n19637), .ZN(n16810) );
  NAND2_X1 U24620 ( .A1(n26923), .A2(n13393), .ZN(n17025) );
  INV_X1 U24626 ( .I(n18146), .ZN(n18145) );
  NAND2_X1 U24630 ( .A1(n26803), .A2(n26802), .ZN(n20797) );
  NAND2_X1 U24631 ( .A1(n20669), .A2(n26961), .ZN(n17601) );
  OAI21_X1 U24636 ( .A1(n26937), .A2(n875), .B(n17993), .ZN(n26856) );
  NOR2_X1 U24638 ( .A1(n26734), .A2(n9188), .ZN(n16924) );
  NAND2_X1 U24639 ( .A1(n13758), .A2(n13757), .ZN(n14861) );
  NAND2_X1 U24641 ( .A1(n27347), .A2(n993), .ZN(n18651) );
  INV_X1 U24642 ( .I(n18652), .ZN(n27138) );
  NOR3_X1 U24658 ( .A1(n26672), .A2(n17158), .A3(n36480), .ZN(n14989) );
  NOR2_X1 U24659 ( .A1(n1207), .A2(n34166), .ZN(n20305) );
  NAND2_X1 U24661 ( .A1(n3158), .A2(n13457), .ZN(n21224) );
  NAND2_X1 U24664 ( .A1(n27875), .A2(n17378), .ZN(n27901) );
  NOR3_X1 U24671 ( .A1(n17253), .A2(n1212), .A3(n15357), .ZN(n17254) );
  NAND3_X1 U24675 ( .A1(n17410), .A2(n988), .A3(n13081), .ZN(n28075) );
  INV_X1 U24677 ( .I(n29223), .ZN(n15395) );
  NAND2_X1 U24680 ( .A1(n16343), .A2(n28598), .ZN(n16272) );
  INV_X1 U24682 ( .I(n29034), .ZN(n18523) );
  NAND2_X1 U24683 ( .A1(n28577), .A2(n28674), .ZN(n28307) );
  NAND2_X1 U24684 ( .A1(n17644), .A2(n39830), .ZN(n20288) );
  INV_X1 U24686 ( .I(n29768), .ZN(n29692) );
  NOR2_X1 U24687 ( .A1(n19424), .A2(n29900), .ZN(n17779) );
  INV_X1 U24688 ( .I(n30233), .ZN(n14891) );
  NAND2_X1 U24691 ( .A1(n14428), .A2(n21269), .ZN(n28880) );
  NOR2_X1 U24693 ( .A1(n31444), .A2(n29774), .ZN(n18221) );
  NOR2_X1 U24695 ( .A1(n21285), .A2(n32571), .ZN(n17632) );
  INV_X2 U24696 ( .I(n20080), .ZN(n30043) );
  INV_X1 U24698 ( .I(n19050), .ZN(n20251) );
  NAND2_X1 U24699 ( .A1(n29438), .A2(n29439), .ZN(n16960) );
  AOI21_X1 U24701 ( .A1(n29543), .A2(n21072), .B(n29559), .ZN(n21071) );
  NAND2_X1 U24702 ( .A1(n19272), .A2(n29548), .ZN(n21072) );
  AOI21_X1 U24703 ( .A1(n29546), .A2(n29548), .B(n29558), .ZN(n29542) );
  INV_X1 U24704 ( .I(n29558), .ZN(n29550) );
  NAND2_X1 U24706 ( .A1(n29567), .A2(n29574), .ZN(n15308) );
  NAND2_X1 U24707 ( .A1(n29797), .A2(n18257), .ZN(n21012) );
  NAND2_X1 U24710 ( .A1(n15466), .A2(n20277), .ZN(n21058) );
  OAI21_X1 U24712 ( .A1(n21666), .A2(n21833), .B(n21436), .ZN(n21361) );
  NOR2_X1 U24716 ( .A1(n22019), .A2(n36006), .ZN(n19958) );
  OAI22_X1 U24717 ( .A1(n21431), .A2(n21682), .B1(n21681), .B2(n21683), .ZN(
        n21356) );
  NAND2_X1 U24718 ( .A1(n35973), .A2(n21681), .ZN(n21354) );
  NAND3_X1 U24721 ( .A1(n33771), .A2(n21762), .A3(n11851), .ZN(n15613) );
  NAND2_X1 U24723 ( .A1(n21964), .A2(n10261), .ZN(n20043) );
  NAND2_X1 U24727 ( .A1(n19850), .A2(n17102), .ZN(n16231) );
  NAND2_X1 U24730 ( .A1(n9970), .A2(n22234), .ZN(n18064) );
  NOR2_X1 U24731 ( .A1(n9970), .A2(n1329), .ZN(n16228) );
  NAND2_X1 U24735 ( .A1(n21863), .A2(n19609), .ZN(n14995) );
  NOR2_X1 U24739 ( .A1(n22236), .A2(n22235), .ZN(n18129) );
  INV_X1 U24743 ( .I(n15268), .ZN(n18272) );
  NAND2_X1 U24748 ( .A1(n13855), .A2(n21885), .ZN(n15816) );
  AOI21_X1 U24750 ( .A1(n19416), .A2(n18266), .B(n1353), .ZN(n16762) );
  NOR2_X1 U24753 ( .A1(n21656), .A2(n17938), .ZN(n17433) );
  INV_X1 U24757 ( .I(n16347), .ZN(n16345) );
  NOR2_X1 U24758 ( .A1(n39594), .A2(n21478), .ZN(n14945) );
  NOR2_X1 U24761 ( .A1(n17869), .A2(n1676), .ZN(n17334) );
  AOI21_X1 U24763 ( .A1(n18657), .A2(n21924), .B(n21923), .ZN(n20844) );
  NOR2_X1 U24765 ( .A1(n20681), .A2(n21837), .ZN(n20680) );
  OAI21_X1 U24767 ( .A1(n1372), .A2(n19709), .B(n21703), .ZN(n21704) );
  OAI21_X1 U24768 ( .A1(n16302), .A2(n21887), .B(n21889), .ZN(n15929) );
  NOR2_X1 U24770 ( .A1(n18542), .A2(n19543), .ZN(n18561) );
  AOI21_X1 U24772 ( .A1(n21591), .A2(n21590), .B(n19434), .ZN(n21598) );
  NAND2_X1 U24773 ( .A1(n33086), .A2(n22262), .ZN(n16625) );
  NAND2_X1 U24774 ( .A1(n18926), .A2(n21920), .ZN(n21736) );
  NOR2_X1 U24776 ( .A1(n18205), .A2(n21528), .ZN(n17967) );
  NAND2_X1 U24777 ( .A1(n32525), .A2(n15560), .ZN(n21657) );
  NOR2_X1 U24779 ( .A1(n1354), .A2(n18028), .ZN(n15560) );
  AND2_X1 U24780 ( .A1(n22915), .A2(n23164), .Z(n14628) );
  NOR2_X1 U24781 ( .A1(n36095), .A2(n19293), .ZN(n16604) );
  NAND2_X1 U24782 ( .A1(n39418), .A2(n23171), .ZN(n19177) );
  INV_X1 U24784 ( .I(n12392), .ZN(n21292) );
  NAND2_X1 U24793 ( .A1(n1310), .A2(n23637), .ZN(n23471) );
  AOI21_X1 U24794 ( .A1(n38604), .A2(n9699), .B(n19229), .ZN(n19228) );
  NOR2_X1 U24796 ( .A1(n36839), .A2(n23213), .ZN(n16198) );
  NAND2_X1 U24798 ( .A1(n22918), .A2(n18679), .ZN(n14738) );
  NAND2_X1 U24801 ( .A1(n31234), .A2(n39070), .ZN(n23194) );
  NAND2_X1 U24805 ( .A1(n1300), .A2(n18236), .ZN(n18235) );
  NOR2_X1 U24807 ( .A1(n23548), .A2(n9321), .ZN(n17674) );
  OAI21_X1 U24814 ( .A1(n23184), .A2(n19538), .B(n1314), .ZN(n22965) );
  NAND2_X1 U24815 ( .A1(n21094), .A2(n23098), .ZN(n16956) );
  NOR2_X1 U24816 ( .A1(n23060), .A2(n14560), .ZN(n23062) );
  NAND2_X1 U24817 ( .A1(n17127), .A2(n39810), .ZN(n19083) );
  NOR2_X1 U24818 ( .A1(n19823), .A2(n3452), .ZN(n16615) );
  INV_X1 U24819 ( .I(n22870), .ZN(n22998) );
  NAND3_X1 U24820 ( .A1(n32815), .A2(n19293), .A3(n22996), .ZN(n20214) );
  NOR2_X1 U24821 ( .A1(n1648), .A2(n16104), .ZN(n22894) );
  INV_X1 U24822 ( .I(n24065), .ZN(n19102) );
  NOR2_X1 U24823 ( .A1(n38282), .A2(n12029), .ZN(n16419) );
  NAND2_X1 U24825 ( .A1(n23087), .A2(n531), .ZN(n23093) );
  AOI21_X1 U24830 ( .A1(n31049), .A2(n19469), .B(n1044), .ZN(n15588) );
  NOR3_X1 U24831 ( .A1(n20408), .A2(n23211), .A3(n20407), .ZN(n21119) );
  INV_X1 U24832 ( .I(n20788), .ZN(n23614) );
  NAND2_X1 U24840 ( .A1(n15320), .A2(n11004), .ZN(n24238) );
  INV_X1 U24844 ( .I(n24223), .ZN(n20655) );
  NAND3_X1 U24845 ( .A1(n14265), .A2(n24761), .A3(n33230), .ZN(n20787) );
  NAND2_X1 U24849 ( .A1(n24327), .A2(n1589), .ZN(n16106) );
  NAND2_X1 U24850 ( .A1(n19745), .A2(n24267), .ZN(n16313) );
  NAND2_X1 U24854 ( .A1(n24348), .A2(n24347), .ZN(n24349) );
  OAI21_X1 U24857 ( .A1(n20058), .A2(n37227), .B(n24143), .ZN(n24145) );
  NAND3_X1 U24860 ( .A1(n24157), .A2(n24465), .A3(n17546), .ZN(n24159) );
  NAND2_X1 U24862 ( .A1(n23962), .A2(n6849), .ZN(n21241) );
  NAND2_X1 U24863 ( .A1(n24510), .A2(n24608), .ZN(n15208) );
  NAND2_X1 U24866 ( .A1(n24258), .A2(n38972), .ZN(n19069) );
  NOR2_X1 U24867 ( .A1(n34547), .A2(n20839), .ZN(n18937) );
  AOI21_X1 U24873 ( .A1(n24118), .A2(n24373), .B(n24191), .ZN(n18456) );
  NAND2_X1 U24875 ( .A1(n17246), .A2(n955), .ZN(n17451) );
  NAND2_X1 U24879 ( .A1(n25106), .A2(n24896), .ZN(n24895) );
  NOR2_X1 U24884 ( .A1(n911), .A2(n19767), .ZN(n20216) );
  OAI21_X1 U24886 ( .A1(n17645), .A2(n9682), .B(n26125), .ZN(n14983) );
  NAND3_X1 U24888 ( .A1(n25741), .A2(n25742), .A3(n596), .ZN(n16137) );
  INV_X1 U24899 ( .I(n18031), .ZN(n19514) );
  NOR2_X1 U24902 ( .A1(n25431), .A2(n25649), .ZN(n17182) );
  NAND2_X1 U24908 ( .A1(n1102), .A2(n25965), .ZN(n18038) );
  NOR2_X1 U24909 ( .A1(n33644), .A2(n37502), .ZN(n20235) );
  NAND2_X1 U24914 ( .A1(n834), .A2(n17212), .ZN(n15178) );
  NOR2_X1 U24915 ( .A1(n25721), .A2(n18519), .ZN(n25723) );
  NOR2_X1 U24916 ( .A1(n2752), .A2(n35580), .ZN(n26037) );
  NOR2_X1 U24917 ( .A1(n20699), .A2(n32986), .ZN(n20103) );
  NAND2_X1 U24921 ( .A1(n26934), .A2(n17993), .ZN(n19939) );
  NAND3_X1 U24924 ( .A1(n12290), .A2(n26688), .A3(n26979), .ZN(n26659) );
  NAND3_X1 U24927 ( .A1(n12162), .A2(n25721), .A3(n33826), .ZN(n25572) );
  OAI22_X1 U24928 ( .A1(n26101), .A2(n35207), .B1(n25779), .B2(n25780), .ZN(
        n20738) );
  NOR2_X1 U24929 ( .A1(n25866), .A2(n2830), .ZN(n25774) );
  NAND2_X1 U24930 ( .A1(n1021), .A2(n35207), .ZN(n16181) );
  NAND2_X1 U24933 ( .A1(n34279), .A2(n39417), .ZN(n17662) );
  NOR2_X1 U24934 ( .A1(n17575), .A2(n33279), .ZN(n17574) );
  NAND2_X1 U24937 ( .A1(n32191), .A2(n38211), .ZN(n20244) );
  NAND2_X1 U24938 ( .A1(n26776), .A2(n38120), .ZN(n21021) );
  NAND2_X1 U24939 ( .A1(n19222), .A2(n26905), .ZN(n15897) );
  INV_X1 U24940 ( .I(n27436), .ZN(n16173) );
  NOR2_X1 U24945 ( .A1(n33050), .A2(n27364), .ZN(n18232) );
  NOR2_X1 U24946 ( .A1(n1484), .A2(n34001), .ZN(n19619) );
  NAND2_X1 U24959 ( .A1(n31254), .A2(n26734), .ZN(n21202) );
  INV_X1 U24960 ( .I(n7974), .ZN(n27248) );
  NAND2_X1 U24966 ( .A1(n4411), .A2(n17392), .ZN(n17391) );
  OAI21_X1 U24968 ( .A1(n14862), .A2(n20211), .B(n14861), .ZN(n20546) );
  INV_X1 U24969 ( .I(n26982), .ZN(n26983) );
  NOR2_X1 U24971 ( .A1(n26996), .A2(n13111), .ZN(n17824) );
  INV_X1 U24974 ( .I(n19855), .ZN(n28221) );
  AOI21_X1 U24975 ( .A1(n26671), .A2(n33726), .B(n11138), .ZN(n14991) );
  INV_X1 U24978 ( .I(n20200), .ZN(n20198) );
  NAND2_X1 U24979 ( .A1(n20201), .A2(n20410), .ZN(n20199) );
  NAND2_X1 U24983 ( .A1(n28324), .A2(n33331), .ZN(n27867) );
  NAND2_X1 U24985 ( .A1(n17322), .A2(n28698), .ZN(n19591) );
  NAND2_X1 U24987 ( .A1(n3899), .A2(n37018), .ZN(n19321) );
  NAND3_X1 U24991 ( .A1(n28532), .A2(n38159), .A3(n11413), .ZN(n28508) );
  NAND3_X1 U24999 ( .A1(n28652), .A2(n28653), .A3(n28386), .ZN(n28387) );
  NAND2_X1 U25000 ( .A1(n18341), .A2(n19039), .ZN(n28327) );
  NOR2_X1 U25001 ( .A1(n28283), .A2(n28282), .ZN(n20398) );
  AOI21_X1 U25002 ( .A1(n1426), .A2(n3014), .B(n1415), .ZN(n19795) );
  AND2_X1 U25003 ( .A1(n18036), .A2(n28656), .Z(n14621) );
  NAND2_X1 U25005 ( .A1(n28310), .A2(n28723), .ZN(n14816) );
  NOR2_X1 U25006 ( .A1(n28724), .A2(n28722), .ZN(n28310) );
  NOR2_X1 U25011 ( .A1(n1397), .A2(n10702), .ZN(n16988) );
  NAND2_X1 U25013 ( .A1(n20830), .A2(n29455), .ZN(n29457) );
  NAND2_X1 U25015 ( .A1(n29764), .A2(n29696), .ZN(n29636) );
  NOR2_X1 U25018 ( .A1(n29698), .A2(n1060), .ZN(n16392) );
  OAI21_X1 U25019 ( .A1(n29761), .A2(n31516), .B(n19567), .ZN(n29697) );
  AOI21_X1 U25020 ( .A1(n31516), .A2(n19568), .B(n19599), .ZN(n19567) );
  INV_X1 U25021 ( .I(n29940), .ZN(n29989) );
  OAI21_X1 U25025 ( .A1(n1387), .A2(n1388), .B(n29236), .ZN(n15482) );
  NOR2_X1 U25026 ( .A1(n907), .A2(n19088), .ZN(n17821) );
  NAND2_X1 U25027 ( .A1(n29351), .A2(n12876), .ZN(n29309) );
  AOI21_X1 U25028 ( .A1(n1055), .A2(n29314), .B(n29313), .ZN(n19130) );
  NAND2_X1 U25029 ( .A1(n29315), .A2(n357), .ZN(n19129) );
  NOR2_X1 U25030 ( .A1(n16123), .A2(n29317), .ZN(n14787) );
  NAND2_X1 U25031 ( .A1(n12943), .A2(n29367), .ZN(n29373) );
  NAND2_X1 U25034 ( .A1(n38200), .A2(n29478), .ZN(n29462) );
  NAND2_X1 U25038 ( .A1(n28619), .A2(n505), .ZN(n18726) );
  NAND2_X1 U25040 ( .A1(n1390), .A2(n29664), .ZN(n16596) );
  NAND2_X1 U25041 ( .A1(n29641), .A2(n29660), .ZN(n21033) );
  NAND2_X1 U25045 ( .A1(n17684), .A2(n33358), .ZN(n17683) );
  AOI22_X1 U25046 ( .A1(n17681), .A2(n4849), .B1(n39830), .B2(n21023), .ZN(
        n16996) );
  OAI21_X1 U25048 ( .A1(n29761), .A2(n29760), .B(n16962), .ZN(n29767) );
  NOR2_X1 U25049 ( .A1(n29763), .A2(n17105), .ZN(n16962) );
  NAND2_X1 U25051 ( .A1(n1063), .A2(n29870), .ZN(n19393) );
  NAND2_X1 U25052 ( .A1(n19093), .A2(n18104), .ZN(n15138) );
  INV_X1 U25053 ( .I(n28980), .ZN(n15141) );
  NAND2_X1 U25056 ( .A1(n29949), .A2(n35809), .ZN(n29951) );
  NAND2_X1 U25057 ( .A1(n21166), .A2(n30058), .ZN(n17982) );
  NOR2_X1 U25058 ( .A1(n11861), .A2(n29996), .ZN(n17633) );
  NAND2_X1 U25060 ( .A1(n16180), .A2(n35187), .ZN(n16722) );
  INV_X1 U25063 ( .I(n32415), .ZN(n29183) );
  NOR2_X1 U25064 ( .A1(n30177), .A2(n20342), .ZN(n14998) );
  NOR2_X1 U25066 ( .A1(n37659), .A2(n33280), .ZN(n18755) );
  OAI21_X1 U25070 ( .A1(n16016), .A2(n2532), .B(n21889), .ZN(n16014) );
  INV_X1 U25075 ( .I(n1048), .ZN(n17639) );
  NOR2_X1 U25079 ( .A1(n36237), .A2(n20799), .ZN(n20798) );
  NAND2_X1 U25080 ( .A1(n17940), .A2(n15175), .ZN(n17939) );
  NAND2_X1 U25081 ( .A1(n9970), .A2(n20943), .ZN(n22061) );
  NAND2_X1 U25082 ( .A1(n16262), .A2(n21288), .ZN(n16453) );
  NOR2_X1 U25084 ( .A1(n1152), .A2(n16265), .ZN(n16452) );
  INV_X1 U25085 ( .I(n2233), .ZN(n22445) );
  INV_X1 U25086 ( .I(n22495), .ZN(n18189) );
  NAND3_X1 U25087 ( .A1(n22209), .A2(n30315), .A3(n22208), .ZN(n22210) );
  NAND2_X1 U25090 ( .A1(n22345), .A2(n22341), .ZN(n21967) );
  INV_X1 U25098 ( .I(n16348), .ZN(n16346) );
  INV_X1 U25099 ( .I(n22645), .ZN(n20718) );
  NAND2_X1 U25100 ( .A1(n22190), .A2(n9987), .ZN(n22191) );
  OAI21_X1 U25101 ( .A1(n19486), .A2(n22189), .B(n9987), .ZN(n22193) );
  INV_X1 U25102 ( .I(n22743), .ZN(n17513) );
  NAND2_X1 U25103 ( .A1(n17341), .A2(n30323), .ZN(n17339) );
  NAND3_X1 U25105 ( .A1(n30315), .A2(n22204), .A3(n21288), .ZN(n22096) );
  INV_X1 U25110 ( .I(n22043), .ZN(n17668) );
  INV_X1 U25111 ( .I(n22044), .ZN(n17669) );
  NAND2_X1 U25112 ( .A1(n22944), .A2(n23166), .ZN(n16955) );
  NAND3_X1 U25127 ( .A1(n4147), .A2(n17887), .A3(n23493), .ZN(n22970) );
  INV_X1 U25128 ( .I(n32226), .ZN(n20503) );
  AOI21_X1 U25130 ( .A1(n15579), .A2(n23461), .B(n23238), .ZN(n20322) );
  AOI21_X1 U25132 ( .A1(n22988), .A2(n1135), .B(n36829), .ZN(n16032) );
  NOR2_X1 U25135 ( .A1(n19481), .A2(n19686), .ZN(n21118) );
  NAND2_X1 U25137 ( .A1(n20817), .A2(n39001), .ZN(n18389) );
  NAND2_X1 U25141 ( .A1(n23547), .A2(n1295), .ZN(n17677) );
  AND2_X1 U25143 ( .A1(n1038), .A2(n23515), .Z(n14665) );
  NAND2_X1 U25148 ( .A1(n23264), .A2(n38724), .ZN(n16058) );
  OAI21_X1 U25151 ( .A1(n16443), .A2(n34307), .B(n35068), .ZN(n23557) );
  AOI22_X1 U25155 ( .A1(n20661), .A2(n20343), .B1(n17511), .B2(n23477), .ZN(
        n23466) );
  INV_X1 U25156 ( .I(n23969), .ZN(n23698) );
  NAND2_X1 U25159 ( .A1(n23630), .A2(n39070), .ZN(n19922) );
  NOR2_X1 U25161 ( .A1(n23351), .A2(n17090), .ZN(n14720) );
  NAND2_X1 U25162 ( .A1(n20100), .A2(n31331), .ZN(n23118) );
  INV_X1 U25163 ( .I(n23762), .ZN(n18172) );
  OAI21_X1 U25165 ( .A1(n23039), .A2(n20620), .B(n15797), .ZN(n15800) );
  NOR2_X1 U25166 ( .A1(n15949), .A2(n15798), .ZN(n15797) );
  NOR2_X1 U25167 ( .A1(n17995), .A2(n20620), .ZN(n15798) );
  OAI21_X1 U25169 ( .A1(n20002), .A2(n15210), .B(n39067), .ZN(n18552) );
  NOR2_X1 U25170 ( .A1(n19466), .A2(n21310), .ZN(n18551) );
  INV_X1 U25171 ( .I(n24669), .ZN(n24670) );
  NOR2_X1 U25172 ( .A1(n24668), .A2(n3076), .ZN(n24671) );
  AND2_X1 U25174 ( .A1(n20787), .A2(n24762), .Z(n14548) );
  INV_X1 U25181 ( .I(n24965), .ZN(n16421) );
  AND2_X1 U25185 ( .A1(n37229), .A2(n24433), .Z(n14538) );
  NAND2_X1 U25186 ( .A1(n20027), .A2(n24271), .ZN(n19690) );
  AOI21_X1 U25187 ( .A1(n24738), .A2(n24737), .B(n37389), .ZN(n16670) );
  NAND2_X1 U25191 ( .A1(n24117), .A2(n16547), .ZN(n16785) );
  INV_X1 U25193 ( .I(n16900), .ZN(n15158) );
  NAND3_X1 U25194 ( .A1(n9892), .A2(n1240), .A3(n931), .ZN(n26326) );
  AOI22_X1 U25195 ( .A1(n1515), .A2(n26330), .B1(n14407), .B2(n9892), .ZN(
        n15194) );
  INV_X1 U25197 ( .I(n17891), .ZN(n24606) );
  INV_X1 U25200 ( .I(n16542), .ZN(n16540) );
  INV_X1 U25201 ( .I(n17613), .ZN(n25347) );
  OAI21_X1 U25216 ( .A1(n31557), .A2(n25689), .B(n25690), .ZN(n18146) );
  NAND2_X1 U25218 ( .A1(n25803), .A2(n25965), .ZN(n25585) );
  NOR2_X1 U25220 ( .A1(n4699), .A2(n26098), .ZN(n25785) );
  NAND2_X1 U25221 ( .A1(n1528), .A2(n11848), .ZN(n25817) );
  INV_X1 U25222 ( .I(n17372), .ZN(n17261) );
  NAND2_X1 U25223 ( .A1(n951), .A2(n26109), .ZN(n14810) );
  INV_X1 U25224 ( .I(n35209), .ZN(n18371) );
  NOR2_X1 U25225 ( .A1(n25812), .A2(n26131), .ZN(n21305) );
  NAND2_X1 U25226 ( .A1(n1097), .A2(n4604), .ZN(n18282) );
  INV_X1 U25232 ( .I(n26006), .ZN(n20051) );
  INV_X1 U25241 ( .I(n25841), .ZN(n16424) );
  NOR2_X1 U25243 ( .A1(n27054), .A2(n27341), .ZN(n20915) );
  NOR2_X1 U25244 ( .A1(n25803), .A2(n25965), .ZN(n18037) );
  NAND2_X1 U25245 ( .A1(n19980), .A2(n12162), .ZN(n25559) );
  NOR2_X1 U25246 ( .A1(n25558), .A2(n25557), .ZN(n19980) );
  OAI21_X1 U25250 ( .A1(n27230), .A2(n27415), .B(n27109), .ZN(n15915) );
  NAND2_X1 U25252 ( .A1(n39065), .A2(n27069), .ZN(n20145) );
  NAND2_X1 U25261 ( .A1(n20738), .A2(n32193), .ZN(n15869) );
  NAND2_X1 U25265 ( .A1(n8696), .A2(n27586), .ZN(n27041) );
  INV_X1 U25266 ( .I(n19352), .ZN(n27175) );
  OAI21_X1 U25270 ( .A1(n15433), .A2(n15434), .B(n15432), .ZN(n15430) );
  INV_X1 U25273 ( .I(n27076), .ZN(n18170) );
  INV_X1 U25274 ( .I(n27441), .ZN(n27444) );
  OAI21_X1 U25275 ( .A1(n27306), .A2(n27583), .B(n27585), .ZN(n27307) );
  NAND2_X1 U25278 ( .A1(n38571), .A2(n7291), .ZN(n27146) );
  NAND2_X1 U25279 ( .A1(n27145), .A2(n7291), .ZN(n17058) );
  NAND3_X1 U25283 ( .A1(n27429), .A2(n27428), .A3(n12156), .ZN(n27431) );
  OR2_X1 U25284 ( .A1(n27167), .A2(n27166), .Z(n14586) );
  INV_X1 U25291 ( .I(n16848), .ZN(n19669) );
  INV_X1 U25295 ( .I(n28650), .ZN(n18961) );
  NAND2_X1 U25296 ( .A1(n32543), .A2(n28484), .ZN(n28483) );
  NAND3_X1 U25297 ( .A1(n28756), .A2(n28755), .A3(n16691), .ZN(n28757) );
  NAND2_X1 U25298 ( .A1(n28666), .A2(n28665), .ZN(n21212) );
  NAND2_X1 U25303 ( .A1(n37956), .A2(n14968), .ZN(n14967) );
  INV_X1 U25305 ( .I(n29142), .ZN(n21056) );
  INV_X1 U25309 ( .I(n15015), .ZN(n28670) );
  NAND2_X1 U25312 ( .A1(n28061), .A2(n28060), .ZN(n28062) );
  NOR2_X1 U25315 ( .A1(n18472), .A2(n18471), .ZN(n18470) );
  NOR2_X1 U25316 ( .A1(n28758), .A2(n978), .ZN(n19055) );
  NAND2_X1 U25322 ( .A1(n28323), .A2(n30304), .ZN(n19754) );
  INV_X1 U25325 ( .I(n28943), .ZN(n16640) );
  OAI21_X1 U25328 ( .A1(n20931), .A2(n8805), .B(n37013), .ZN(n29006) );
  NAND2_X1 U25332 ( .A1(n28715), .A2(n19844), .ZN(n28210) );
  NOR2_X1 U25335 ( .A1(n29777), .A2(n29781), .ZN(n21037) );
  INV_X1 U25337 ( .I(n35272), .ZN(n29390) );
  NAND2_X1 U25340 ( .A1(n29525), .A2(n29535), .ZN(n16084) );
  NAND2_X1 U25341 ( .A1(n29546), .A2(n29558), .ZN(n19380) );
  NAND2_X1 U25342 ( .A1(n29721), .A2(n29720), .ZN(n17731) );
  NAND2_X1 U25343 ( .A1(n30022), .A2(n9231), .ZN(n18782) );
  NOR2_X1 U25345 ( .A1(n30109), .A2(n35186), .ZN(n19032) );
  OAI21_X1 U25348 ( .A1(n18611), .A2(n29274), .B(n19090), .ZN(n17955) );
  NOR2_X1 U25353 ( .A1(n29409), .A2(n17849), .ZN(n29405) );
  AOI21_X1 U25354 ( .A1(n29423), .A2(n29440), .B(n1383), .ZN(n19618) );
  NAND2_X1 U25355 ( .A1(n1389), .A2(n29438), .ZN(n15127) );
  NOR2_X1 U25356 ( .A1(n29440), .A2(n17293), .ZN(n15128) );
  NAND2_X1 U25357 ( .A1(n29540), .A2(n29550), .ZN(n28906) );
  OAI21_X1 U25359 ( .A1(n29570), .A2(n29571), .B(n1393), .ZN(n20701) );
  NAND3_X1 U25360 ( .A1(n29570), .A2(n31899), .A3(n29571), .ZN(n15310) );
  NOR2_X1 U25362 ( .A1(n30295), .A2(n19318), .ZN(n29656) );
  NOR3_X1 U25363 ( .A1(n6181), .A2(n19297), .A3(n39689), .ZN(n21032) );
  NOR2_X1 U25364 ( .A1(n21033), .A2(n19318), .ZN(n20444) );
  INV_X1 U25366 ( .I(n18042), .ZN(n29686) );
  NAND3_X1 U25368 ( .A1(n20498), .A2(n5921), .A3(n29722), .ZN(n20499) );
  AOI21_X1 U25369 ( .A1(n21013), .A2(n29788), .B(n21010), .ZN(n21009) );
  NAND2_X1 U25371 ( .A1(n18085), .A2(n18082), .ZN(n29915) );
  INV_X1 U25373 ( .I(n30078), .ZN(n19550) );
  AOI21_X1 U25374 ( .A1(n16723), .A2(n30111), .B(n16721), .ZN(n16720) );
  AOI21_X1 U25377 ( .A1(n10289), .A2(n31527), .B(n17192), .ZN(n21006) );
  AOI21_X1 U25378 ( .A1(n13384), .A2(n10813), .B(n17193), .ZN(n21005) );
  NAND2_X1 U25379 ( .A1(n20538), .A2(n14998), .ZN(n14997) );
  NAND2_X1 U25380 ( .A1(n30176), .A2(n17997), .ZN(n17168) );
  OR2_X1 U25386 ( .A1(n16052), .A2(n21606), .Z(n14420) );
  OR2_X1 U25389 ( .A1(n25387), .A2(n25386), .Z(n14431) );
  NAND2_X1 U25390 ( .A1(n1177), .A2(n10569), .ZN(n14435) );
  NOR2_X1 U25399 ( .A1(n21885), .A2(n15839), .ZN(n14492) );
  XOR2_X1 U25400 ( .A1(n22781), .A2(n22780), .Z(n14494) );
  XNOR2_X1 U25404 ( .A1(n24861), .A2(n24860), .ZN(n14507) );
  OR2_X1 U25407 ( .A1(n1076), .A2(n28150), .Z(n14513) );
  OR2_X1 U25408 ( .A1(n25690), .A2(n25689), .Z(n14518) );
  OR2_X1 U25410 ( .A1(n29675), .A2(n29683), .Z(n14522) );
  XNOR2_X1 U25412 ( .A1(n10027), .A2(n22749), .ZN(n14530) );
  XNOR2_X1 U25414 ( .A1(n9576), .A2(n19875), .ZN(n14533) );
  INV_X1 U25416 ( .I(n19819), .ZN(n22565) );
  INV_X1 U25418 ( .I(n37229), .ZN(n24434) );
  AND2_X1 U25419 ( .A1(n35357), .A2(n28812), .Z(n14543) );
  AND2_X1 U25421 ( .A1(n15194), .A2(n26332), .Z(n14546) );
  INV_X1 U25422 ( .I(n22674), .ZN(n23135) );
  NOR2_X1 U25424 ( .A1(n8700), .A2(n19350), .ZN(n14549) );
  AND2_X1 U25425 ( .A1(n19850), .A2(n21887), .Z(n14551) );
  XNOR2_X1 U25428 ( .A1(n38184), .A2(n35267), .ZN(n14565) );
  INV_X1 U25430 ( .I(n29696), .ZN(n19568) );
  XNOR2_X1 U25431 ( .A1(n14264), .A2(n20706), .ZN(n14566) );
  XNOR2_X1 U25433 ( .A1(n33194), .A2(n30207), .ZN(n14568) );
  XNOR2_X1 U25434 ( .A1(n23357), .A2(n1621), .ZN(n14571) );
  AND2_X1 U25436 ( .A1(n18884), .A2(n11848), .Z(n14579) );
  BUF_X2 U25437 ( .I(n21655), .Z(n17938) );
  AND2_X1 U25438 ( .A1(n17943), .A2(n29411), .Z(n14582) );
  INV_X1 U25442 ( .I(n22204), .ZN(n22351) );
  OR2_X1 U25443 ( .A1(n24687), .A2(n14857), .Z(n14593) );
  AND2_X1 U25444 ( .A1(n23107), .A2(n22005), .Z(n14594) );
  NAND2_X1 U25445 ( .A1(n22101), .A2(n20234), .ZN(n14597) );
  XNOR2_X1 U25449 ( .A1(n16017), .A2(n19775), .ZN(n14603) );
  AND2_X1 U25458 ( .A1(n27163), .A2(n20981), .Z(n14626) );
  AND2_X1 U25459 ( .A1(n20919), .A2(n28053), .Z(n14632) );
  INV_X1 U25463 ( .I(n314), .ZN(n21073) );
  XNOR2_X1 U25467 ( .A1(n25094), .A2(n25095), .ZN(n14646) );
  XNOR2_X1 U25469 ( .A1(n19221), .A2(n20479), .ZN(n14648) );
  XNOR2_X1 U25470 ( .A1(n24002), .A2(n1723), .ZN(n14651) );
  XNOR2_X1 U25473 ( .A1(n39063), .A2(n19913), .ZN(n14670) );
  XNOR2_X1 U25476 ( .A1(n22790), .A2(n29707), .ZN(n14673) );
  INV_X1 U25478 ( .I(n21880), .ZN(n21509) );
  XNOR2_X1 U25479 ( .A1(n26394), .A2(n28934), .ZN(n14675) );
  INV_X1 U25482 ( .I(n25502), .ZN(n15647) );
  INV_X1 U25484 ( .I(n22773), .ZN(n16531) );
  XNOR2_X1 U25487 ( .A1(n29252), .A2(n1734), .ZN(n14689) );
  XNOR2_X1 U25488 ( .A1(n20311), .A2(n20310), .ZN(n14691) );
  XNOR2_X1 U25491 ( .A1(n27746), .A2(n35702), .ZN(n14693) );
  NOR2_X1 U25492 ( .A1(n438), .A2(n759), .ZN(n14696) );
  INV_X1 U25499 ( .I(n27129), .ZN(n20402) );
  INV_X1 U25501 ( .I(n19879), .ZN(n17078) );
  INV_X1 U25502 ( .I(n19760), .ZN(n18981) );
  INV_X1 U25503 ( .I(n19937), .ZN(n20206) );
  INV_X1 U25504 ( .I(n19876), .ZN(n16320) );
  INV_X1 U25505 ( .I(n29554), .ZN(n21121) );
  INV_X1 U25506 ( .I(n30090), .ZN(n18109) );
  INV_X1 U25507 ( .I(n19866), .ZN(n17603) );
  INV_X1 U25509 ( .I(n19808), .ZN(n20658) );
  INV_X1 U25510 ( .I(n9981), .ZN(n18432) );
  INV_X1 U25511 ( .I(n10027), .ZN(n16618) );
  INV_X1 U25512 ( .I(n29411), .ZN(n17551) );
  INV_X1 U25513 ( .I(n30169), .ZN(n15203) );
  INV_X1 U25517 ( .I(n19936), .ZN(n16562) );
  INV_X1 U25518 ( .I(n19613), .ZN(n16332) );
  INV_X1 U25520 ( .I(n29221), .ZN(n17257) );
  INV_X1 U25521 ( .I(n19860), .ZN(n17463) );
  INV_X1 U25522 ( .I(n29269), .ZN(n19128) );
  INV_X1 U25524 ( .I(n30068), .ZN(n21294) );
  INV_X1 U25525 ( .I(n30248), .ZN(n18296) );
  INV_X1 U25526 ( .I(n29602), .ZN(n15432) );
  BUF_X2 U25527 ( .I(Key[65]), .Z(n29801) );
  XOR2_X1 U25532 ( .A1(n19862), .A2(n29320), .Z(n18015) );
  XOR2_X1 U25536 ( .A1(n25246), .A2(n14716), .Z(n14715) );
  XOR2_X1 U25537 ( .A1(n19156), .A2(n25280), .Z(n14716) );
  XOR2_X1 U25538 ( .A1(n16318), .A2(n16321), .Z(n24308) );
  NOR2_X1 U25540 ( .A1(n8597), .A2(n21587), .ZN(n21589) );
  AOI21_X2 U25541 ( .A1(n15491), .A2(n14721), .B(n14720), .ZN(n23667) );
  NOR2_X1 U25543 ( .A1(n22964), .A2(n14725), .ZN(n15084) );
  XOR2_X1 U25550 ( .A1(n27594), .A2(n15776), .Z(n14756) );
  INV_X2 U25551 ( .I(n14758), .ZN(n22682) );
  NOR2_X1 U25552 ( .A1(n23533), .A2(n14759), .ZN(n16395) );
  XOR2_X1 U25553 ( .A1(n18273), .A2(n39183), .Z(n19493) );
  NAND2_X1 U25555 ( .A1(n25946), .A2(n39729), .ZN(n14762) );
  XOR2_X1 U25556 ( .A1(n15288), .A2(n14772), .Z(n14771) );
  XOR2_X1 U25561 ( .A1(n15165), .A2(n24999), .Z(n25087) );
  XOR2_X1 U25563 ( .A1(Plaintext[171]), .A2(Key[171]), .Z(n15370) );
  OR2_X1 U25564 ( .A1(n20021), .A2(n14488), .Z(n14798) );
  NAND2_X1 U25569 ( .A1(n1126), .A2(n19864), .ZN(n24069) );
  XOR2_X1 U25575 ( .A1(n14808), .A2(n27834), .Z(n27472) );
  XOR2_X1 U25577 ( .A1(n14818), .A2(n14821), .Z(n19806) );
  XOR2_X1 U25578 ( .A1(n24058), .A2(n14819), .Z(n14818) );
  XOR2_X1 U25582 ( .A1(Plaintext[173]), .A2(Key[173]), .Z(n15152) );
  MUX2_X1 U25585 ( .I0(n28647), .I1(n15296), .S(n30805), .Z(n15295) );
  XOR2_X1 U25586 ( .A1(n29027), .A2(n14844), .Z(n14843) );
  XOR2_X1 U25587 ( .A1(n19513), .A2(n14956), .Z(n14844) );
  XOR2_X1 U25591 ( .A1(n25101), .A2(n14859), .Z(n18121) );
  XOR2_X1 U25592 ( .A1(n7728), .A2(n16492), .Z(n25100) );
  XOR2_X1 U25595 ( .A1(n26511), .A2(n26510), .Z(n14867) );
  XOR2_X1 U25600 ( .A1(n14425), .A2(n24919), .Z(n24920) );
  NAND2_X1 U25602 ( .A1(n23595), .A2(n23596), .ZN(n23314) );
  XOR2_X1 U25605 ( .A1(n35231), .A2(n1734), .Z(n14887) );
  XOR2_X1 U25606 ( .A1(n22465), .A2(n22600), .Z(n14888) );
  NAND2_X1 U25609 ( .A1(n39322), .A2(n14891), .ZN(n29203) );
  XOR2_X1 U25612 ( .A1(n2233), .A2(n19735), .Z(n14894) );
  NOR2_X1 U25615 ( .A1(n28559), .A2(n1197), .ZN(n14900) );
  XOR2_X1 U25618 ( .A1(n27855), .A2(n19885), .Z(n14907) );
  NOR2_X1 U25620 ( .A1(n1158), .A2(n21837), .ZN(n14911) );
  XOR2_X1 U25623 ( .A1(n18974), .A2(n18973), .Z(n26668) );
  XOR2_X1 U25630 ( .A1(n24018), .A2(n35196), .Z(n23981) );
  NAND2_X2 U25632 ( .A1(n25516), .A2(n19209), .ZN(n25798) );
  XOR2_X1 U25638 ( .A1(n28953), .A2(n14956), .Z(n28813) );
  XOR2_X1 U25640 ( .A1(n25071), .A2(n14970), .Z(n17457) );
  XOR2_X1 U25643 ( .A1(n26348), .A2(n1096), .Z(n14978) );
  INV_X1 U25644 ( .I(n23992), .ZN(n24311) );
  XOR2_X1 U25645 ( .A1(n22703), .A2(n4413), .Z(n14979) );
  NOR2_X2 U25646 ( .A1(n21976), .A2(n17027), .ZN(n19931) );
  INV_X2 U25647 ( .I(n19685), .ZN(n23028) );
  XNOR2_X1 U25648 ( .A1(n14981), .A2(n14982), .ZN(n14980) );
  XOR2_X1 U25650 ( .A1(n18127), .A2(n29097), .Z(n14982) );
  OAI22_X1 U25651 ( .A1(n3826), .A2(n17158), .B1(n11226), .B2(n38377), .ZN(
        n26829) );
  OAI21_X1 U25654 ( .A1(n15269), .A2(n14500), .B(n33516), .ZN(n28013) );
  NAND3_X2 U25655 ( .A1(n17221), .A2(n27093), .A3(n27094), .ZN(n17220) );
  INV_X1 U25656 ( .I(n15007), .ZN(n15006) );
  XOR2_X1 U25658 ( .A1(n15012), .A2(n21278), .Z(n22674) );
  XOR2_X1 U25660 ( .A1(n38850), .A2(n19592), .Z(n15013) );
  OAI22_X1 U25661 ( .A1(n28800), .A2(n28799), .B1(n19905), .B2(n15015), .ZN(
        n28801) );
  NAND2_X1 U25662 ( .A1(n15015), .A2(n19905), .ZN(n28800) );
  OAI21_X1 U25664 ( .A1(n21950), .A2(n32664), .B(n15019), .ZN(n21952) );
  XOR2_X1 U25666 ( .A1(n27516), .A2(n35188), .Z(n27169) );
  INV_X2 U25669 ( .I(n15036), .ZN(n25660) );
  INV_X2 U25672 ( .I(n15052), .ZN(n25481) );
  AOI21_X2 U25674 ( .A1(n18340), .A2(n15053), .B(n18338), .ZN(n22058) );
  XOR2_X1 U25677 ( .A1(n38158), .A2(n35266), .Z(n15056) );
  NOR2_X2 U25678 ( .A1(n32791), .A2(n28753), .ZN(n28754) );
  XOR2_X1 U25679 ( .A1(n17423), .A2(n18849), .Z(n15972) );
  XOR2_X1 U25680 ( .A1(n25163), .A2(n33184), .Z(n18643) );
  XOR2_X1 U25681 ( .A1(n38951), .A2(n15888), .Z(n15753) );
  OAI21_X1 U25682 ( .A1(n29497), .A2(n15063), .B(n29498), .ZN(n20720) );
  NOR2_X1 U25683 ( .A1(n38051), .A2(n17424), .ZN(n15063) );
  XOR2_X1 U25685 ( .A1(n28603), .A2(n28607), .Z(n15071) );
  NAND2_X1 U25686 ( .A1(n19871), .A2(n20703), .ZN(n21654) );
  OAI22_X1 U25687 ( .A1(n21904), .A2(n21903), .B1(n21900), .B2(n21902), .ZN(
        n15072) );
  NOR2_X1 U25689 ( .A1(n36530), .A2(n15075), .ZN(n15074) );
  MUX2_X1 U25692 ( .I0(n27484), .I1(n1218), .S(n3977), .Z(n27485) );
  XOR2_X1 U25696 ( .A1(n29297), .A2(n4816), .Z(n15090) );
  XOR2_X1 U25699 ( .A1(n37874), .A2(n29295), .Z(n15093) );
  XOR2_X1 U25700 ( .A1(n23931), .A2(n19732), .Z(n15094) );
  AOI21_X1 U25703 ( .A1(n28717), .A2(n28716), .B(n5093), .ZN(n27941) );
  XOR2_X1 U25710 ( .A1(n15126), .A2(n18584), .Z(n15516) );
  OAI21_X1 U25712 ( .A1(n29435), .A2(n29437), .B(n11506), .ZN(n15132) );
  AOI21_X1 U25714 ( .A1(n29960), .A2(n29957), .B(n15140), .ZN(n15139) );
  INV_X2 U25719 ( .I(n15152), .ZN(n18293) );
  XOR2_X1 U25720 ( .A1(n15156), .A2(n19629), .Z(n28710) );
  XOR2_X1 U25721 ( .A1(n15156), .A2(n20804), .Z(n29155) );
  OR2_X1 U25723 ( .A1(n22976), .A2(n15163), .Z(n21245) );
  XOR2_X1 U25725 ( .A1(n22749), .A2(n1700), .Z(n15171) );
  XOR2_X1 U25730 ( .A1(Plaintext[144]), .A2(Key[144]), .Z(n15619) );
  XOR2_X1 U25733 ( .A1(n15186), .A2(n1377), .Z(n15226) );
  INV_X2 U25737 ( .I(n27985), .ZN(n28054) );
  INV_X2 U25738 ( .I(n15195), .ZN(n21254) );
  XOR2_X1 U25740 ( .A1(n27858), .A2(n19932), .Z(n15197) );
  OAI21_X1 U25744 ( .A1(n15209), .A2(n17262), .B(n29574), .ZN(n29575) );
  NOR2_X1 U25748 ( .A1(n1126), .A2(n21310), .ZN(n15210) );
  NOR2_X2 U25749 ( .A1(n16467), .A2(n27921), .ZN(n19844) );
  XOR2_X1 U25750 ( .A1(n15213), .A2(n15212), .Z(n18308) );
  XOR2_X1 U25751 ( .A1(n22557), .A2(n22556), .Z(n15212) );
  XOR2_X1 U25752 ( .A1(n18778), .A2(n22629), .Z(n22556) );
  XOR2_X1 U25753 ( .A1(n22411), .A2(n36290), .Z(n22557) );
  XOR2_X1 U25754 ( .A1(n17987), .A2(n15214), .Z(n15213) );
  XOR2_X1 U25756 ( .A1(n28860), .A2(n28946), .Z(n21271) );
  XOR2_X1 U25757 ( .A1(n28827), .A2(n19741), .Z(n28860) );
  XOR2_X1 U25758 ( .A1(n15216), .A2(n28777), .Z(n16554) );
  XOR2_X1 U25759 ( .A1(n15220), .A2(n19986), .Z(n15938) );
  XOR2_X1 U25762 ( .A1(n21380), .A2(Key[130]), .Z(n21761) );
  XOR2_X1 U25765 ( .A1(n17606), .A2(n25217), .Z(n15227) );
  NAND2_X2 U25767 ( .A1(n19999), .A2(n20000), .ZN(n25127) );
  NAND2_X1 U25770 ( .A1(n15233), .A2(n19362), .ZN(n15232) );
  INV_X2 U25774 ( .I(n18308), .ZN(n22929) );
  NAND2_X1 U25776 ( .A1(n24193), .A2(n15240), .ZN(n16882) );
  XOR2_X1 U25781 ( .A1(n14454), .A2(n23280), .Z(n15250) );
  NAND3_X1 U25783 ( .A1(n24359), .A2(n24360), .A3(n38431), .ZN(n15257) );
  XOR2_X1 U25790 ( .A1(n27842), .A2(n31438), .Z(n15286) );
  XOR2_X1 U25791 ( .A1(Plaintext[172]), .A2(Key[172]), .Z(n18968) );
  XOR2_X1 U25795 ( .A1(n28925), .A2(n3633), .Z(n15303) );
  XOR2_X1 U25797 ( .A1(n14638), .A2(n14476), .Z(n15305) );
  NAND2_X1 U25798 ( .A1(n29571), .A2(n29570), .ZN(n29563) );
  XOR2_X1 U25801 ( .A1(n15316), .A2(n15315), .Z(n18544) );
  XOR2_X1 U25802 ( .A1(n25093), .A2(n24931), .Z(n15315) );
  MUX2_X1 U25807 ( .I0(n15172), .I1(n9751), .S(n15443), .Z(n15444) );
  XOR2_X1 U25811 ( .A1(n15340), .A2(n22621), .Z(n15339) );
  XOR2_X1 U25812 ( .A1(n22647), .A2(n19755), .Z(n15340) );
  XOR2_X1 U25815 ( .A1(n871), .A2(n15349), .Z(n15348) );
  XOR2_X1 U25816 ( .A1(n27730), .A2(n19763), .Z(n15349) );
  OAI22_X1 U25818 ( .A1(n18558), .A2(n15350), .B1(n9876), .B2(n22341), .ZN(
        n19270) );
  NOR2_X1 U25820 ( .A1(n36754), .A2(n11274), .ZN(n21573) );
  XOR2_X1 U25823 ( .A1(n10647), .A2(n14565), .Z(n15361) );
  NOR2_X1 U25825 ( .A1(n14783), .A2(n19372), .ZN(n21629) );
  NAND2_X1 U25826 ( .A1(n18968), .A2(n14783), .ZN(n21726) );
  NOR2_X1 U25830 ( .A1(n17792), .A2(n19397), .ZN(n15381) );
  NAND2_X1 U25831 ( .A1(n29687), .A2(n38206), .ZN(n29667) );
  INV_X2 U25832 ( .I(n19741), .ZN(n29829) );
  XOR2_X1 U25834 ( .A1(n19308), .A2(n28860), .Z(n15384) );
  INV_X2 U25835 ( .I(n15386), .ZN(n17217) );
  INV_X1 U25836 ( .I(n8585), .ZN(n26477) );
  XOR2_X1 U25837 ( .A1(Plaintext[76]), .A2(Key[76]), .Z(n18542) );
  INV_X2 U25838 ( .I(n25544), .ZN(n16933) );
  XOR2_X1 U25841 ( .A1(n28914), .A2(n15394), .Z(n15393) );
  XOR2_X1 U25842 ( .A1(n13852), .A2(n15395), .Z(n15394) );
  XOR2_X1 U25845 ( .A1(n27683), .A2(n1356), .Z(n15398) );
  XOR2_X1 U25851 ( .A1(n39116), .A2(n19929), .Z(n18604) );
  XOR2_X1 U25852 ( .A1(n36750), .A2(n19729), .Z(n22278) );
  INV_X2 U25853 ( .I(n15412), .ZN(n22935) );
  INV_X1 U25862 ( .I(n18880), .ZN(n19171) );
  NAND2_X1 U25867 ( .A1(n22277), .A2(n9616), .ZN(n15436) );
  XOR2_X1 U25869 ( .A1(n38896), .A2(n37024), .Z(n15442) );
  XOR2_X1 U25873 ( .A1(n15450), .A2(n15451), .Z(n16062) );
  INV_X2 U25878 ( .I(n15463), .ZN(n23163) );
  NOR2_X1 U25880 ( .A1(n24602), .A2(n34011), .ZN(n17270) );
  XOR2_X1 U25885 ( .A1(n5841), .A2(n15679), .Z(n20486) );
  XOR2_X1 U25887 ( .A1(n15476), .A2(n24078), .Z(n20270) );
  XOR2_X1 U25888 ( .A1(n24079), .A2(n15477), .Z(n15476) );
  XOR2_X1 U25891 ( .A1(n35222), .A2(n1724), .Z(n15481) );
  XOR2_X1 U25892 ( .A1(n26548), .A2(n29003), .Z(n25985) );
  XOR2_X1 U25893 ( .A1(n26548), .A2(n19081), .Z(n18808) );
  XOR2_X1 U25894 ( .A1(n20956), .A2(n26548), .Z(n15529) );
  XOR2_X1 U25898 ( .A1(n9757), .A2(n19732), .Z(n15500) );
  NOR2_X1 U25899 ( .A1(n37200), .A2(n918), .ZN(n21524) );
  INV_X2 U25900 ( .I(n20591), .ZN(n20590) );
  XOR2_X1 U25902 ( .A1(n23843), .A2(n15507), .Z(n24106) );
  XOR2_X1 U25903 ( .A1(n14454), .A2(n23839), .Z(n15507) );
  XOR2_X1 U25904 ( .A1(n26489), .A2(n1727), .Z(n15508) );
  INV_X2 U25906 ( .I(n19928), .ZN(n15515) );
  NAND2_X2 U25908 ( .A1(n19701), .A2(n15515), .ZN(n25528) );
  OAI21_X1 U25910 ( .A1(n15357), .A2(n31832), .B(n15518), .ZN(n28008) );
  MUX2_X1 U25911 ( .I0(n36850), .I1(n29864), .S(n29938), .Z(n29866) );
  INV_X1 U25912 ( .I(n18115), .ZN(n25019) );
  XOR2_X1 U25916 ( .A1(n22495), .A2(n16199), .Z(n18416) );
  XOR2_X1 U25918 ( .A1(n20452), .A2(n29025), .Z(n28780) );
  XOR2_X1 U25919 ( .A1(n38844), .A2(n19624), .Z(n26059) );
  XOR2_X1 U25920 ( .A1(n38844), .A2(n1361), .Z(n18322) );
  XOR2_X1 U25921 ( .A1(n11667), .A2(n38844), .Z(n26557) );
  XOR2_X1 U25922 ( .A1(n27688), .A2(n15546), .Z(n15545) );
  XOR2_X1 U25923 ( .A1(n15547), .A2(n27689), .Z(n15546) );
  XOR2_X1 U25927 ( .A1(n25236), .A2(n25235), .Z(n19644) );
  XOR2_X1 U25928 ( .A1(n25323), .A2(n25160), .Z(n25232) );
  XOR2_X1 U25932 ( .A1(n39739), .A2(n38181), .Z(n15565) );
  NAND2_X1 U25934 ( .A1(n39112), .A2(n28228), .ZN(n15572) );
  XOR2_X1 U25936 ( .A1(n33511), .A2(n21294), .Z(n20811) );
  XOR2_X1 U25937 ( .A1(n33511), .A2(n19738), .Z(n28870) );
  XOR2_X1 U25939 ( .A1(n22542), .A2(n19738), .Z(n18888) );
  XOR2_X1 U25940 ( .A1(n15591), .A2(n7602), .Z(n26073) );
  INV_X2 U25943 ( .I(n15598), .ZN(n20896) );
  XOR2_X1 U25944 ( .A1(n15600), .A2(n15599), .Z(Ciphertext[2]) );
  XOR2_X1 U25946 ( .A1(n22624), .A2(n30179), .Z(n15607) );
  NOR2_X1 U25949 ( .A1(n30184), .A2(n30178), .ZN(n15615) );
  NOR2_X2 U25950 ( .A1(n15684), .A2(n15685), .ZN(n15616) );
  XOR2_X1 U25956 ( .A1(n23779), .A2(n37842), .Z(n23691) );
  NAND2_X1 U25961 ( .A1(n9394), .A2(n15651), .ZN(n29201) );
  XOR2_X1 U25966 ( .A1(n22743), .A2(n15654), .Z(n15653) );
  XOR2_X1 U25967 ( .A1(n33323), .A2(n19760), .Z(n15654) );
  XOR2_X1 U25969 ( .A1(n26587), .A2(n33735), .Z(n15656) );
  XOR2_X1 U25971 ( .A1(n34469), .A2(n30094), .Z(n15660) );
  NAND3_X1 U25973 ( .A1(n24804), .A2(n15664), .A3(n14064), .ZN(n15689) );
  MUX2_X1 U25974 ( .I0(n34354), .I1(n15664), .S(n36471), .Z(n24573) );
  AOI21_X1 U25976 ( .A1(n28323), .A2(n13601), .B(n3845), .ZN(n28060) );
  XOR2_X1 U25977 ( .A1(n15674), .A2(n15672), .Z(n20063) );
  XOR2_X1 U25979 ( .A1(n26595), .A2(n26594), .Z(n15673) );
  XOR2_X1 U25982 ( .A1(n24030), .A2(n15679), .Z(n23681) );
  XOR2_X1 U25983 ( .A1(n35936), .A2(n15679), .Z(n23562) );
  NAND2_X2 U25984 ( .A1(n23557), .A2(n23558), .ZN(n15679) );
  AOI21_X2 U25986 ( .A1(n23363), .A2(n23364), .B(n15681), .ZN(n24040) );
  OAI22_X2 U25989 ( .A1(n18025), .A2(n17923), .B1(n21607), .B2(n18026), .ZN(
        n15697) );
  XOR2_X1 U25991 ( .A1(Plaintext[147]), .A2(Key[147]), .Z(n21933) );
  AOI21_X2 U25994 ( .A1(n28083), .A2(n986), .B(n28082), .ZN(n28638) );
  XOR2_X1 U26001 ( .A1(n27794), .A2(n16618), .Z(n15721) );
  XOR2_X1 U26002 ( .A1(n35303), .A2(n27754), .Z(n15722) );
  XOR2_X1 U26004 ( .A1(n27498), .A2(n27850), .Z(n27795) );
  XOR2_X1 U26009 ( .A1(n23662), .A2(n15729), .Z(n15728) );
  XOR2_X1 U26010 ( .A1(n23888), .A2(n19624), .Z(n15729) );
  XOR2_X1 U26011 ( .A1(n12570), .A2(n24028), .Z(n15730) );
  XOR2_X1 U26012 ( .A1(n22588), .A2(n17078), .Z(n22525) );
  INV_X2 U26014 ( .I(n15839), .ZN(n21579) );
  NOR3_X1 U26015 ( .A1(n31530), .A2(n35137), .A3(n9197), .ZN(n15735) );
  NOR2_X1 U26017 ( .A1(n23174), .A2(n14130), .ZN(n15739) );
  XOR2_X1 U26020 ( .A1(n18242), .A2(n15745), .Z(n29251) );
  NAND3_X1 U26022 ( .A1(n1139), .A2(n17511), .A3(n34558), .ZN(n16098) );
  NOR2_X1 U26023 ( .A1(n16094), .A2(n34558), .ZN(n20661) );
  XOR2_X1 U26024 ( .A1(n38816), .A2(n19561), .Z(n27550) );
  XOR2_X1 U26026 ( .A1(n10221), .A2(n29934), .Z(n15750) );
  XOR2_X1 U26028 ( .A1(n27707), .A2(n36894), .Z(n27816) );
  XOR2_X1 U26029 ( .A1(n27524), .A2(n27522), .Z(n15757) );
  XOR2_X1 U26030 ( .A1(n15758), .A2(n30435), .Z(n19198) );
  XOR2_X1 U26033 ( .A1(n22763), .A2(n35211), .Z(n15762) );
  NOR2_X1 U26036 ( .A1(n26135), .A2(n36798), .ZN(n15767) );
  INV_X1 U26037 ( .I(n15768), .ZN(n29355) );
  INV_X2 U26040 ( .I(n16339), .ZN(n16461) );
  NAND2_X1 U26041 ( .A1(n7975), .A2(n7974), .ZN(n19276) );
  NAND2_X1 U26042 ( .A1(n7973), .A2(n7975), .ZN(n27028) );
  NOR2_X1 U26043 ( .A1(n26870), .A2(n7975), .ZN(n26871) );
  XOR2_X1 U26044 ( .A1(n26435), .A2(n38279), .Z(n18975) );
  NAND2_X1 U26046 ( .A1(n15773), .A2(n29883), .ZN(n29876) );
  XOR2_X1 U26047 ( .A1(n27799), .A2(n15776), .Z(n27800) );
  XOR2_X1 U26048 ( .A1(n15776), .A2(n19851), .Z(n18539) );
  XOR2_X1 U26054 ( .A1(n29159), .A2(n21172), .Z(n15782) );
  AOI21_X1 U26059 ( .A1(n28654), .A2(n28617), .B(n15792), .ZN(n28562) );
  NAND2_X1 U26062 ( .A1(n17967), .A2(n39627), .ZN(n15804) );
  NAND2_X2 U26063 ( .A1(n15806), .A2(n15805), .ZN(n22160) );
  NAND2_X1 U26064 ( .A1(n21663), .A2(n21662), .ZN(n15806) );
  XOR2_X1 U26065 ( .A1(n15810), .A2(n15809), .Z(n15808) );
  XOR2_X1 U26066 ( .A1(n29050), .A2(n19820), .Z(n15809) );
  XOR2_X1 U26068 ( .A1(n21142), .A2(n15819), .Z(n15818) );
  XOR2_X1 U26075 ( .A1(n9719), .A2(n33990), .Z(n15824) );
  XOR2_X1 U26079 ( .A1(n18242), .A2(n19677), .Z(n15835) );
  XOR2_X1 U26086 ( .A1(n29253), .A2(n29238), .Z(n29161) );
  NAND2_X1 U26088 ( .A1(n22354), .A2(n22353), .ZN(n16266) );
  INV_X1 U26090 ( .I(n16658), .ZN(n16656) );
  NOR3_X1 U26091 ( .A1(n31542), .A2(n35203), .A3(n1187), .ZN(n18472) );
  OAI21_X1 U26092 ( .A1(n17942), .A2(n1670), .B(n22676), .ZN(n17340) );
  NAND2_X1 U26097 ( .A1(n12537), .A2(n28340), .ZN(n28341) );
  OAI21_X1 U26098 ( .A1(n19657), .A2(n27866), .B(n16476), .ZN(n28195) );
  NOR2_X1 U26101 ( .A1(n29704), .A2(n29635), .ZN(n20433) );
  NAND2_X1 U26108 ( .A1(n19404), .A2(n9993), .ZN(n18494) );
  OAI21_X1 U26111 ( .A1(n18408), .A2(n22274), .B(n35771), .ZN(n16351) );
  NAND2_X1 U26114 ( .A1(n7265), .A2(n39160), .ZN(n25368) );
  NAND2_X1 U26115 ( .A1(n7644), .A2(n32024), .ZN(n16726) );
  NOR2_X1 U26123 ( .A1(n26089), .A2(n9743), .ZN(n17439) );
  NAND2_X1 U26125 ( .A1(n20348), .A2(n1351), .ZN(n17483) );
  AOI21_X1 U26129 ( .A1(n1679), .A2(n22316), .B(n9824), .ZN(n22320) );
  OAI21_X1 U26130 ( .A1(n14422), .A2(n14400), .B(n29446), .ZN(n17089) );
  NOR2_X1 U26140 ( .A1(n37089), .A2(n22243), .ZN(n22244) );
  NOR2_X1 U26141 ( .A1(n19084), .A2(n16128), .ZN(n16130) );
  INV_X1 U26151 ( .I(n10747), .ZN(n18479) );
  INV_X1 U26153 ( .I(n18806), .ZN(n19508) );
  INV_X1 U26156 ( .I(n8473), .ZN(n18623) );
  NAND2_X1 U26163 ( .A1(n28193), .A2(n27866), .ZN(n16476) );
  INV_X1 U26166 ( .I(Key[94]), .ZN(n15838) );
  XOR2_X1 U26170 ( .A1(n38147), .A2(n34239), .Z(n21157) );
  XOR2_X1 U26171 ( .A1(n38147), .A2(n29554), .Z(n28502) );
  NAND2_X1 U26172 ( .A1(n15841), .A2(n29439), .ZN(n15840) );
  OAI22_X1 U26173 ( .A1(n18495), .A2(n15841), .B1(n29435), .B2(n29434), .ZN(
        n19689) );
  XOR2_X1 U26180 ( .A1(n25174), .A2(n15858), .Z(n15857) );
  XOR2_X1 U26181 ( .A1(n25155), .A2(n19952), .Z(n15858) );
  XOR2_X1 U26182 ( .A1(n15862), .A2(n15861), .Z(n15859) );
  XOR2_X1 U26183 ( .A1(n23671), .A2(n12972), .Z(n15861) );
  INV_X1 U26186 ( .I(n15867), .ZN(n21011) );
  NOR2_X1 U26187 ( .A1(n15867), .A2(n29792), .ZN(n29783) );
  MUX2_X1 U26188 ( .I0(n15867), .I1(n18257), .S(n29792), .Z(n29790) );
  OAI21_X1 U26189 ( .A1(n29782), .A2(n15867), .B(n29789), .ZN(n21013) );
  NAND2_X1 U26193 ( .A1(n31412), .A2(n15868), .ZN(n17972) );
  NAND2_X2 U26194 ( .A1(n23859), .A2(n23858), .ZN(n25269) );
  MUX2_X1 U26200 ( .I0(n24490), .I1(n15878), .S(n9212), .Z(n15877) );
  NAND2_X1 U26204 ( .A1(n16302), .A2(n33280), .ZN(n15891) );
  XNOR2_X1 U26206 ( .A1(n20550), .A2(n15893), .ZN(n15892) );
  XOR2_X1 U26207 ( .A1(n20777), .A2(n15894), .Z(n15893) );
  XOR2_X1 U26208 ( .A1(n3917), .A2(n36065), .Z(n15894) );
  INV_X2 U26210 ( .I(n15903), .ZN(n24296) );
  AOI22_X2 U26211 ( .A1(n34547), .A2(n24296), .B1(n13453), .B2(n33939), .ZN(
        n24209) );
  XOR2_X1 U26214 ( .A1(n24038), .A2(n23893), .Z(n24006) );
  INV_X2 U26217 ( .I(n15913), .ZN(n26802) );
  XOR2_X1 U26222 ( .A1(n15916), .A2(n19775), .Z(n16244) );
  XOR2_X1 U26223 ( .A1(n35245), .A2(n29334), .Z(n20678) );
  NAND3_X1 U26232 ( .A1(n37040), .A2(n27416), .A3(n33773), .ZN(n18640) );
  XOR2_X1 U26233 ( .A1(n1468), .A2(n27802), .Z(n15932) );
  XOR2_X1 U26240 ( .A1(n32354), .A2(n34017), .Z(n17721) );
  XOR2_X1 U26242 ( .A1(n20082), .A2(n26392), .Z(n16440) );
  XOR2_X1 U26249 ( .A1(n18482), .A2(n23847), .Z(n15987) );
  XOR2_X1 U26250 ( .A1(n15989), .A2(n16775), .Z(n25392) );
  OAI21_X2 U26257 ( .A1(n17683), .A2(n17682), .B(n16996), .ZN(n29719) );
  MUX2_X1 U26259 ( .I0(n23036), .I1(n23037), .S(n1145), .Z(n16007) );
  XOR2_X1 U26261 ( .A1(n29037), .A2(n28589), .Z(n16010) );
  XOR2_X1 U26266 ( .A1(n23967), .A2(n39073), .Z(n23790) );
  XOR2_X1 U26268 ( .A1(n16022), .A2(n5116), .Z(n16021) );
  XOR2_X1 U26269 ( .A1(n23623), .A2(n1724), .Z(n16022) );
  XOR2_X1 U26271 ( .A1(n30612), .A2(n18432), .Z(n16029) );
  XOR2_X1 U26272 ( .A1(n23892), .A2(n16030), .Z(n23773) );
  XOR2_X1 U26274 ( .A1(n18006), .A2(n23655), .Z(n23892) );
  NAND2_X1 U26275 ( .A1(n16034), .A2(n14596), .ZN(n28113) );
  XOR2_X1 U26281 ( .A1(n38753), .A2(n20206), .Z(n16046) );
  XOR2_X1 U26283 ( .A1(n16054), .A2(n15960), .Z(n28579) );
  NAND2_X2 U26289 ( .A1(n16075), .A2(n30002), .ZN(n30022) );
  NAND2_X1 U26292 ( .A1(n25641), .A2(n38963), .ZN(n16095) );
  OR2_X1 U26293 ( .A1(n19713), .A2(n24874), .Z(n16097) );
  XOR2_X1 U26295 ( .A1(n18362), .A2(n29363), .Z(n18363) );
  NOR2_X1 U26296 ( .A1(n27030), .A2(n2522), .ZN(n27033) );
  XOR2_X1 U26297 ( .A1(n27692), .A2(n772), .Z(n16103) );
  XOR2_X1 U26302 ( .A1(n22758), .A2(n22419), .Z(n22420) );
  XOR2_X1 U26303 ( .A1(n29093), .A2(n29092), .Z(n18127) );
  XOR2_X1 U26309 ( .A1(n33916), .A2(n16332), .Z(n16131) );
  XOR2_X1 U26310 ( .A1(n16135), .A2(n25023), .Z(n16134) );
  XOR2_X1 U26311 ( .A1(n31112), .A2(n25165), .Z(n16135) );
  XOR2_X1 U26317 ( .A1(n16151), .A2(n16150), .Z(n16149) );
  XOR2_X1 U26318 ( .A1(n38880), .A2(n1622), .Z(n16151) );
  XOR2_X1 U26322 ( .A1(n16864), .A2(n1718), .Z(n24575) );
  XOR2_X1 U26325 ( .A1(n39575), .A2(n19883), .Z(n16175) );
  INV_X1 U26328 ( .I(n16182), .ZN(n23361) );
  NOR2_X1 U26329 ( .A1(n16182), .A2(n23482), .ZN(n22513) );
  XOR2_X1 U26330 ( .A1(n35266), .A2(n29357), .Z(n27555) );
  XOR2_X1 U26336 ( .A1(n39756), .A2(n25193), .Z(n16192) );
  XOR2_X1 U26337 ( .A1(n16193), .A2(n16694), .Z(n19838) );
  OAI21_X2 U26340 ( .A1(n22851), .A2(n22861), .B(n16202), .ZN(n23352) );
  NAND2_X1 U26341 ( .A1(n24072), .A2(n21310), .ZN(n24083) );
  NOR2_X1 U26343 ( .A1(n16209), .A2(n4849), .ZN(n28375) );
  NOR2_X1 U26344 ( .A1(n19994), .A2(n16209), .ZN(n17682) );
  AND2_X1 U26347 ( .A1(n13393), .A2(n26763), .Z(n16221) );
  XOR2_X1 U26349 ( .A1(n28913), .A2(n16705), .Z(n16225) );
  XOR2_X1 U26350 ( .A1(n26602), .A2(n30010), .Z(n20261) );
  XOR2_X1 U26351 ( .A1(n26602), .A2(n29320), .Z(n26143) );
  XOR2_X1 U26352 ( .A1(n26602), .A2(n19020), .Z(n19019) );
  XOR2_X1 U26353 ( .A1(n17798), .A2(n26602), .Z(n17797) );
  INV_X1 U26354 ( .I(n16233), .ZN(n17975) );
  NAND2_X1 U26355 ( .A1(n29276), .A2(n16233), .ZN(n29281) );
  XOR2_X1 U26356 ( .A1(n35190), .A2(n19908), .Z(n16269) );
  XOR2_X1 U26357 ( .A1(n35189), .A2(n1697), .Z(n20263) );
  XOR2_X1 U26360 ( .A1(n26157), .A2(n20213), .Z(n26434) );
  XOR2_X1 U26361 ( .A1(n16249), .A2(n17705), .Z(Ciphertext[12]) );
  XOR2_X1 U26362 ( .A1(n23764), .A2(n30063), .Z(n16257) );
  XOR2_X1 U26363 ( .A1(n31247), .A2(n32973), .Z(n16258) );
  OAI21_X1 U26365 ( .A1(n35272), .A2(n16260), .B(n9790), .ZN(n29406) );
  OAI21_X1 U26366 ( .A1(n20724), .A2(n16260), .B(n35272), .ZN(n29392) );
  XOR2_X1 U26368 ( .A1(n27630), .A2(n16269), .Z(n16268) );
  XOR2_X1 U26369 ( .A1(Plaintext[105]), .A2(Key[105]), .Z(n18757) );
  INV_X2 U26370 ( .I(n16356), .ZN(n29828) );
  NAND3_X1 U26375 ( .A1(n21067), .A2(n21066), .A3(n19933), .ZN(n16291) );
  INV_X1 U26376 ( .I(n16293), .ZN(n16292) );
  AOI21_X1 U26377 ( .A1(n21067), .A2(n21066), .B(n19933), .ZN(n16293) );
  INV_X1 U26378 ( .I(n23885), .ZN(n23964) );
  INV_X2 U26379 ( .I(n18741), .ZN(n18870) );
  XOR2_X1 U26380 ( .A1(n25275), .A2(n29141), .Z(n24921) );
  XOR2_X1 U26382 ( .A1(n16342), .A2(n34945), .Z(n23465) );
  NOR2_X1 U26383 ( .A1(n28754), .A2(n16303), .ZN(n17007) );
  NAND3_X1 U26386 ( .A1(n39656), .A2(n19549), .A3(n16305), .ZN(n22116) );
  NAND2_X1 U26392 ( .A1(n1405), .A2(n16328), .ZN(n16874) );
  AOI21_X1 U26393 ( .A1(n1405), .A2(n30043), .B(n16328), .ZN(n29952) );
  XOR2_X1 U26394 ( .A1(n29072), .A2(n28972), .Z(n28319) );
  XOR2_X1 U26398 ( .A1(Key[103]), .A2(Plaintext[103]), .Z(n16333) );
  XOR2_X1 U26401 ( .A1(n23758), .A2(n16338), .Z(n16337) );
  NAND2_X1 U26403 ( .A1(n26090), .A2(n19889), .ZN(n18003) );
  XOR2_X1 U26406 ( .A1(n973), .A2(n16357), .Z(n17452) );
  XOR2_X1 U26407 ( .A1(n25326), .A2(n16350), .Z(n20151) );
  XOR2_X1 U26408 ( .A1(n25093), .A2(n24922), .Z(n25326) );
  XOR2_X1 U26409 ( .A1(n29082), .A2(n20329), .Z(n16358) );
  XOR2_X1 U26411 ( .A1(n27690), .A2(n27736), .Z(n16362) );
  XOR2_X1 U26414 ( .A1(n32863), .A2(n19629), .Z(n22745) );
  XOR2_X1 U26415 ( .A1(n22643), .A2(n32863), .Z(n22387) );
  XOR2_X1 U26420 ( .A1(n16379), .A2(n28945), .Z(n16378) );
  XOR2_X1 U26421 ( .A1(n28927), .A2(n29081), .Z(n16379) );
  XOR2_X1 U26422 ( .A1(n26395), .A2(n14675), .Z(n16381) );
  NAND2_X2 U26423 ( .A1(n16390), .A2(n16389), .ZN(n29720) );
  NOR2_X1 U26424 ( .A1(n29700), .A2(n29699), .ZN(n16391) );
  XOR2_X1 U26426 ( .A1(n33916), .A2(n29838), .Z(n16679) );
  NAND2_X1 U26429 ( .A1(n28153), .A2(n28151), .ZN(n16412) );
  XOR2_X1 U26430 ( .A1(n1262), .A2(n19722), .Z(n16417) );
  INV_X1 U26431 ( .I(n25149), .ZN(n16422) );
  XOR2_X1 U26432 ( .A1(n16424), .A2(n17051), .Z(n16423) );
  XOR2_X1 U26433 ( .A1(n26487), .A2(n26407), .Z(n25841) );
  XOR2_X1 U26436 ( .A1(n17349), .A2(n19897), .Z(n16439) );
  AOI21_X1 U26439 ( .A1(n16455), .A2(n22205), .B(n21288), .ZN(n16454) );
  XOR2_X1 U26442 ( .A1(n16460), .A2(n19676), .Z(n25331) );
  XOR2_X1 U26443 ( .A1(n16460), .A2(n25194), .Z(n17258) );
  XOR2_X1 U26445 ( .A1(n16469), .A2(n30094), .Z(Ciphertext[154]) );
  NOR2_X1 U26446 ( .A1(n30097), .A2(n30096), .ZN(n16470) );
  OR2_X1 U26450 ( .A1(n35903), .A2(n26031), .Z(n16478) );
  INV_X1 U26451 ( .I(n25615), .ZN(n25617) );
  XOR2_X1 U26454 ( .A1(n16492), .A2(n25298), .Z(n25300) );
  XNOR2_X1 U26456 ( .A1(Plaintext[28]), .A2(Key[28]), .ZN(n16496) );
  XOR2_X1 U26457 ( .A1(n26404), .A2(n16498), .Z(n16497) );
  INV_X1 U26458 ( .I(n17716), .ZN(n26028) );
  NOR2_X1 U26464 ( .A1(n14453), .A2(n26945), .ZN(n16522) );
  XOR2_X1 U26465 ( .A1(n29104), .A2(n29661), .Z(n16529) );
  INV_X1 U26469 ( .I(n32637), .ZN(n24810) );
  XOR2_X1 U26471 ( .A1(n1460), .A2(n35178), .Z(n16549) );
  XOR2_X1 U26472 ( .A1(n27850), .A2(n29671), .Z(n16550) );
  XOR2_X1 U26474 ( .A1(n26225), .A2(n16557), .Z(n16556) );
  XOR2_X1 U26475 ( .A1(n12838), .A2(n10904), .Z(n16557) );
  XOR2_X1 U26477 ( .A1(n22508), .A2(n22645), .Z(n22486) );
  XOR2_X1 U26481 ( .A1(n22713), .A2(n16561), .Z(n16560) );
  XOR2_X1 U26482 ( .A1(n1323), .A2(n16562), .Z(n16561) );
  XOR2_X1 U26483 ( .A1(n22712), .A2(n21201), .Z(n16563) );
  XOR2_X1 U26485 ( .A1(n16743), .A2(n19722), .Z(n16565) );
  XOR2_X1 U26486 ( .A1(n22503), .A2(n16667), .Z(n22569) );
  NAND2_X1 U26488 ( .A1(n24394), .A2(n16449), .ZN(n17947) );
  XOR2_X1 U26490 ( .A1(n16584), .A2(n16582), .Z(n28436) );
  XOR2_X1 U26491 ( .A1(n28545), .A2(n16583), .Z(n16582) );
  XOR2_X1 U26495 ( .A1(n26404), .A2(n19763), .Z(n16591) );
  NOR2_X1 U26500 ( .A1(n1390), .A2(n19297), .ZN(n16598) );
  XOR2_X1 U26509 ( .A1(n38208), .A2(n30101), .Z(n24067) );
  NAND2_X1 U26510 ( .A1(n29708), .A2(n16629), .ZN(n16628) );
  NAND2_X1 U26511 ( .A1(n35771), .A2(n16635), .ZN(n16634) );
  XOR2_X1 U26512 ( .A1(n16639), .A2(n16640), .Z(n16976) );
  NAND2_X1 U26514 ( .A1(n35761), .A2(n33580), .ZN(n16645) );
  XOR2_X1 U26515 ( .A1(n22511), .A2(n1369), .Z(n16648) );
  INV_X2 U26516 ( .I(n38901), .ZN(n26972) );
  XOR2_X1 U26518 ( .A1(n22594), .A2(n19775), .Z(n16651) );
  NOR2_X1 U26520 ( .A1(n35151), .A2(n39015), .ZN(n20884) );
  XOR2_X1 U26522 ( .A1(n26525), .A2(n1503), .Z(n16665) );
  AOI21_X1 U26523 ( .A1(n21012), .A2(n16682), .B(n21011), .ZN(n21010) );
  XOR2_X1 U26526 ( .A1(n29254), .A2(n19736), .Z(n16685) );
  XOR2_X1 U26527 ( .A1(n22760), .A2(n16688), .Z(n16687) );
  XOR2_X1 U26528 ( .A1(n22761), .A2(n30068), .Z(n16688) );
  XOR2_X1 U26529 ( .A1(n22759), .A2(n16690), .Z(n16689) );
  XOR2_X1 U26531 ( .A1(n16695), .A2(n28887), .Z(n16694) );
  XOR2_X1 U26532 ( .A1(n23787), .A2(n17150), .Z(n16698) );
  XOR2_X1 U26534 ( .A1(n29093), .A2(n19674), .Z(n16705) );
  NAND2_X1 U26537 ( .A1(n19837), .A2(n16265), .ZN(n18163) );
  NAND3_X1 U26538 ( .A1(n22351), .A2(n19837), .A3(n35060), .ZN(n22012) );
  XOR2_X1 U26541 ( .A1(n16720), .A2(n1703), .Z(Ciphertext[156]) );
  OAI21_X1 U26542 ( .A1(n30100), .A2(n10118), .B(n30112), .ZN(n16723) );
  XOR2_X1 U26547 ( .A1(n4828), .A2(n29363), .Z(n16735) );
  XOR2_X1 U26549 ( .A1(n29064), .A2(n16741), .Z(n16740) );
  XOR2_X1 U26550 ( .A1(n19571), .A2(n29666), .Z(n16741) );
  XOR2_X1 U26551 ( .A1(n29066), .A2(n29065), .Z(n16742) );
  XOR2_X1 U26552 ( .A1(n16743), .A2(n19933), .Z(n27695) );
  XOR2_X1 U26559 ( .A1(n27534), .A2(n19814), .Z(n16759) );
  XOR2_X1 U26562 ( .A1(n12221), .A2(n26460), .Z(n17487) );
  XOR2_X1 U26564 ( .A1(n23869), .A2(n23699), .Z(n16766) );
  XOR2_X1 U26568 ( .A1(n39575), .A2(n28968), .Z(n23665) );
  XOR2_X1 U26571 ( .A1(n16771), .A2(n20748), .Z(n20560) );
  XOR2_X1 U26572 ( .A1(n16771), .A2(n18700), .Z(n29143) );
  XOR2_X1 U26573 ( .A1(n16771), .A2(n36513), .Z(n19445) );
  NOR2_X1 U26574 ( .A1(n9066), .A2(n33939), .ZN(n24149) );
  OAI21_X1 U26575 ( .A1(n19914), .A2(n14458), .B(n16773), .ZN(n26137) );
  XOR2_X1 U26576 ( .A1(n1505), .A2(n26476), .Z(n16998) );
  XOR2_X1 U26577 ( .A1(n38171), .A2(n19359), .Z(n16776) );
  XOR2_X1 U26578 ( .A1(n11974), .A2(n29718), .Z(n16783) );
  XOR2_X1 U26582 ( .A1(n32776), .A2(n19943), .Z(n23683) );
  NAND3_X1 U26584 ( .A1(n10618), .A2(n35777), .A3(n17771), .ZN(n16791) );
  XNOR2_X1 U26585 ( .A1(n16795), .A2(n16793), .ZN(n16792) );
  XOR2_X1 U26586 ( .A1(n16794), .A2(n16796), .Z(n16793) );
  XOR2_X1 U26587 ( .A1(n1618), .A2(n23910), .Z(n16794) );
  XOR2_X1 U26589 ( .A1(n23905), .A2(n29298), .Z(n16796) );
  XOR2_X1 U26590 ( .A1(n38208), .A2(n23686), .Z(n16797) );
  NAND2_X1 U26591 ( .A1(n22818), .A2(n1315), .ZN(n20177) );
  XOR2_X1 U26592 ( .A1(n16802), .A2(n16799), .Z(n19685) );
  XOR2_X1 U26593 ( .A1(n16801), .A2(n16800), .Z(n16799) );
  XOR2_X1 U26594 ( .A1(n22790), .A2(n29394), .Z(n16800) );
  XOR2_X1 U26595 ( .A1(n22789), .A2(n36290), .Z(n16801) );
  NAND2_X2 U26597 ( .A1(n17287), .A2(n17302), .ZN(n16803) );
  XOR2_X1 U26598 ( .A1(n900), .A2(n19839), .Z(n16806) );
  NAND2_X2 U26603 ( .A1(n25018), .A2(n18115), .ZN(n24965) );
  NOR2_X1 U26605 ( .A1(n38193), .A2(n39583), .ZN(n18716) );
  NAND2_X1 U26610 ( .A1(n496), .A2(n16853), .ZN(n19391) );
  NAND2_X1 U26611 ( .A1(n28733), .A2(n16853), .ZN(n27553) );
  NAND2_X1 U26612 ( .A1(n24782), .A2(n24779), .ZN(n16855) );
  NOR2_X1 U26619 ( .A1(n26186), .A2(n16878), .ZN(n26188) );
  OR2_X1 U26624 ( .A1(n34171), .A2(n2937), .Z(n28297) );
  NAND2_X1 U26625 ( .A1(n18671), .A2(n32790), .ZN(n16985) );
  XOR2_X1 U26629 ( .A1(n31320), .A2(n27704), .Z(n16886) );
  NOR2_X1 U26630 ( .A1(n1492), .A2(n19712), .ZN(n26148) );
  NOR2_X1 U26637 ( .A1(n25892), .A2(n15677), .ZN(n16904) );
  NAND3_X1 U26641 ( .A1(n24783), .A2(n1121), .A3(n38658), .ZN(n24414) );
  XOR2_X1 U26644 ( .A1(n18291), .A2(n22666), .Z(n16912) );
  NAND2_X2 U26647 ( .A1(n16929), .A2(n23427), .ZN(n23955) );
  AOI21_X1 U26649 ( .A1(n29431), .A2(n29435), .B(n19618), .ZN(n19617) );
  AND2_X1 U26655 ( .A1(n19692), .A2(n22895), .Z(n20344) );
  NAND3_X1 U26659 ( .A1(n38210), .A2(n10004), .A3(n25609), .ZN(n19257) );
  XOR2_X1 U26660 ( .A1(n21408), .A2(Key[163]), .Z(n18739) );
  XOR2_X1 U26662 ( .A1(n22663), .A2(n22662), .Z(n21278) );
  OAI21_X1 U26664 ( .A1(n29440), .A2(n29438), .B(n16960), .ZN(n17317) );
  NAND2_X2 U26668 ( .A1(n25775), .A2(n25777), .ZN(n18827) );
  XOR2_X1 U26671 ( .A1(n28944), .A2(n16976), .Z(n16975) );
  NAND2_X1 U26676 ( .A1(n18908), .A2(n29682), .ZN(n29688) );
  NOR2_X1 U26677 ( .A1(n25468), .A2(n25606), .ZN(n17480) );
  NAND2_X1 U26678 ( .A1(n19796), .A2(n19795), .ZN(n19794) );
  XOR2_X1 U26679 ( .A1(n16992), .A2(n38265), .Z(Ciphertext[129]) );
  OAI21_X1 U26684 ( .A1(n12290), .A2(n26686), .B(n852), .ZN(n17099) );
  INV_X1 U26686 ( .I(n27875), .ZN(n27998) );
  XOR2_X1 U26687 ( .A1(n25211), .A2(n24886), .Z(n25178) );
  INV_X1 U26688 ( .I(n23394), .ZN(n22912) );
  XOR2_X1 U26690 ( .A1(n25299), .A2(n25300), .Z(n18869) );
  XNOR2_X1 U26691 ( .A1(n26599), .A2(n19876), .ZN(n17858) );
  NAND2_X1 U26699 ( .A1(n29551), .A2(n29558), .ZN(n28907) );
  NAND2_X2 U26701 ( .A1(n25731), .A2(n25732), .ZN(n17915) );
  XOR2_X1 U26702 ( .A1(n17028), .A2(n14646), .Z(n25613) );
  XOR2_X1 U26703 ( .A1(n25091), .A2(n25092), .Z(n17028) );
  XOR2_X1 U26704 ( .A1(n17030), .A2(n29978), .Z(Ciphertext[136]) );
  NOR2_X1 U26705 ( .A1(n22904), .A2(n22813), .ZN(n22903) );
  XOR2_X1 U26709 ( .A1(n27856), .A2(n17033), .Z(n27857) );
  XOR2_X1 U26710 ( .A1(n27854), .A2(n27855), .Z(n17033) );
  NOR2_X1 U26719 ( .A1(n21604), .A2(n21783), .ZN(n18340) );
  XOR2_X1 U26725 ( .A1(n29553), .A2(n29554), .Z(Ciphertext[64]) );
  NAND3_X1 U26726 ( .A1(n17152), .A2(n39305), .A3(n27263), .ZN(n17151) );
  NAND2_X1 U26729 ( .A1(n36191), .A2(n23450), .ZN(n17470) );
  XOR2_X1 U26731 ( .A1(n17063), .A2(n25736), .Z(n26796) );
  XOR2_X1 U26734 ( .A1(n29115), .A2(n29252), .Z(n28574) );
  NAND2_X1 U26738 ( .A1(n1268), .A2(n24900), .ZN(n17377) );
  XOR2_X1 U26739 ( .A1(n29165), .A2(n29614), .Z(n28824) );
  OR2_X1 U26740 ( .A1(n21958), .A2(n17086), .Z(n21959) );
  NAND2_X1 U26741 ( .A1(n19134), .A2(n19840), .ZN(n21065) );
  OR2_X1 U26743 ( .A1(n22340), .A2(n22341), .Z(n21988) );
  XOR2_X1 U26745 ( .A1(n25197), .A2(n25283), .Z(n25060) );
  OAI21_X1 U26751 ( .A1(n17382), .A2(n29662), .B(n1390), .ZN(n17381) );
  XOR2_X1 U26752 ( .A1(n17113), .A2(n1702), .Z(Ciphertext[71]) );
  NAND2_X1 U26761 ( .A1(n21997), .A2(n22265), .ZN(n18401) );
  INV_X2 U26762 ( .I(n17119), .ZN(n17127) );
  XOR2_X1 U26765 ( .A1(n25039), .A2(n25041), .Z(n17129) );
  XOR2_X1 U26766 ( .A1(n7432), .A2(n30207), .Z(n19201) );
  XOR2_X1 U26767 ( .A1(n38330), .A2(n7432), .Z(n20719) );
  NAND3_X1 U26770 ( .A1(n25374), .A2(n25375), .A3(n35508), .ZN(n25376) );
  XOR2_X1 U26772 ( .A1(n26458), .A2(n38177), .Z(n17136) );
  XOR2_X1 U26774 ( .A1(n26572), .A2(n26277), .Z(n17137) );
  XOR2_X1 U26776 ( .A1(n10579), .A2(n20263), .Z(n17139) );
  XOR2_X1 U26777 ( .A1(n35707), .A2(n17705), .Z(n17704) );
  INV_X1 U26778 ( .I(n27325), .ZN(n27400) );
  NAND2_X1 U26782 ( .A1(n1333), .A2(n22228), .ZN(n17147) );
  XOR2_X1 U26784 ( .A1(n23886), .A2(n19919), .Z(n17150) );
  XOR2_X1 U26785 ( .A1(n37094), .A2(n29371), .Z(n17153) );
  XOR2_X1 U26786 ( .A1(n22453), .A2(n11308), .Z(n22550) );
  NAND2_X2 U26787 ( .A1(n21658), .A2(n21657), .ZN(n19655) );
  NAND2_X1 U26791 ( .A1(n14418), .A2(n21779), .ZN(n17160) );
  XOR2_X1 U26793 ( .A1(n39129), .A2(n30104), .Z(n25734) );
  XOR2_X1 U26794 ( .A1(n39129), .A2(n19817), .Z(n26323) );
  XOR2_X1 U26795 ( .A1(n17171), .A2(n17172), .Z(n20389) );
  XOR2_X1 U26797 ( .A1(n26154), .A2(n26156), .Z(n17172) );
  XOR2_X1 U26801 ( .A1(n27731), .A2(n31551), .Z(n18511) );
  XOR2_X1 U26802 ( .A1(n19231), .A2(n14691), .Z(n17177) );
  NOR2_X2 U26803 ( .A1(n20369), .A2(n29631), .ZN(n29662) );
  XOR2_X1 U26805 ( .A1(n17189), .A2(n30010), .Z(n22001) );
  XOR2_X1 U26806 ( .A1(n17189), .A2(n29785), .Z(n22568) );
  XOR2_X1 U26809 ( .A1(Plaintext[126]), .A2(Key[126]), .Z(n20703) );
  INV_X2 U26810 ( .I(n31596), .ZN(n20979) );
  INV_X2 U26812 ( .I(n17210), .ZN(n20267) );
  OAI21_X1 U26813 ( .A1(n17212), .A2(n1245), .B(n17211), .ZN(n17213) );
  NAND3_X1 U26814 ( .A1(n28143), .A2(n28142), .A3(n17114), .ZN(n28145) );
  INV_X2 U26815 ( .I(n19806), .ZN(n24461) );
  NOR2_X1 U26817 ( .A1(n29347), .A2(n29120), .ZN(n20508) );
  NOR3_X1 U26819 ( .A1(n17233), .A2(n1351), .A3(n19202), .ZN(n17678) );
  XOR2_X1 U26821 ( .A1(n7667), .A2(n35702), .Z(n17245) );
  XOR2_X1 U26823 ( .A1(n25097), .A2(n24924), .Z(n18765) );
  NAND2_X1 U26825 ( .A1(n17249), .A2(n6604), .ZN(n21552) );
  NOR2_X1 U26828 ( .A1(n18603), .A2(n34120), .ZN(n17253) );
  XOR2_X1 U26829 ( .A1(n17256), .A2(n17258), .Z(n17255) );
  XOR2_X1 U26830 ( .A1(n25250), .A2(n17257), .Z(n17256) );
  NOR2_X1 U26833 ( .A1(n30731), .A2(n19542), .ZN(n17264) );
  XOR2_X1 U26835 ( .A1(n35241), .A2(n27858), .Z(n17272) );
  XOR2_X1 U26836 ( .A1(n27362), .A2(n17274), .Z(n17273) );
  XOR2_X1 U26837 ( .A1(n27564), .A2(n17275), .Z(n17274) );
  XOR2_X1 U26838 ( .A1(n27724), .A2(n27516), .Z(n27362) );
  NOR2_X1 U26841 ( .A1(n20223), .A2(n26619), .ZN(n17278) );
  NAND2_X1 U26843 ( .A1(n19367), .A2(n17281), .ZN(n25571) );
  XOR2_X1 U26844 ( .A1(n22728), .A2(n36290), .Z(n17283) );
  XOR2_X1 U26845 ( .A1(n22729), .A2(n30006), .Z(n17285) );
  XOR2_X1 U26847 ( .A1(n17292), .A2(n24859), .Z(n25106) );
  AOI21_X1 U26848 ( .A1(n29435), .A2(n18502), .B(n17293), .ZN(n17318) );
  NOR2_X1 U26850 ( .A1(n25454), .A2(n31375), .ZN(n17297) );
  INV_X1 U26855 ( .I(n28696), .ZN(n17322) );
  XOR2_X1 U26857 ( .A1(n29303), .A2(n28889), .Z(n17325) );
  XOR2_X1 U26859 ( .A1(n31112), .A2(n30090), .Z(n17328) );
  NAND2_X2 U26863 ( .A1(n22312), .A2(n22311), .ZN(n22453) );
  NAND2_X1 U26865 ( .A1(n14590), .A2(n17357), .ZN(n17356) );
  AOI21_X1 U26866 ( .A1(n1675), .A2(n22228), .B(n1333), .ZN(n17357) );
  OR2_X1 U26867 ( .A1(n22089), .A2(n17359), .Z(n17358) );
  XOR2_X1 U26869 ( .A1(n26484), .A2(n21100), .Z(n17361) );
  XOR2_X1 U26870 ( .A1(n17366), .A2(n34945), .Z(Ciphertext[68]) );
  OR2_X1 U26872 ( .A1(n26114), .A2(n31624), .Z(n17373) );
  AOI21_X1 U26873 ( .A1(n29658), .A2(n17382), .B(n17381), .ZN(n20443) );
  XOR2_X1 U26876 ( .A1(Plaintext[148]), .A2(Key[148]), .Z(n18027) );
  XOR2_X1 U26877 ( .A1(n7402), .A2(n19905), .Z(n20730) );
  OAI21_X1 U26879 ( .A1(n28679), .A2(n33646), .B(n28719), .ZN(n19304) );
  XOR2_X1 U26881 ( .A1(n17850), .A2(n1713), .Z(n17404) );
  XOR2_X1 U26882 ( .A1(n27471), .A2(n27472), .Z(n17406) );
  XOR2_X1 U26883 ( .A1(n27728), .A2(n14693), .Z(n20693) );
  XOR2_X1 U26885 ( .A1(n22776), .A2(n39787), .Z(n17429) );
  NAND3_X1 U26889 ( .A1(n32616), .A2(n31234), .A3(n34307), .ZN(n23632) );
  NOR2_X1 U26892 ( .A1(n20364), .A2(n5515), .ZN(n20363) );
  NAND2_X1 U26899 ( .A1(n20274), .A2(n17469), .ZN(n29008) );
  NOR2_X1 U26901 ( .A1(n24713), .A2(n24899), .ZN(n17473) );
  XOR2_X1 U26906 ( .A1(n17492), .A2(n17489), .Z(n19949) );
  XOR2_X1 U26907 ( .A1(n17491), .A2(n17490), .Z(n17489) );
  XOR2_X1 U26908 ( .A1(n23686), .A2(n29849), .Z(n17490) );
  XOR2_X1 U26909 ( .A1(n23952), .A2(n35942), .Z(n17491) );
  XOR2_X1 U26911 ( .A1(n28867), .A2(n20033), .Z(n17494) );
  XOR2_X1 U26914 ( .A1(n38370), .A2(n19905), .Z(n23940) );
  XOR2_X1 U26915 ( .A1(n39038), .A2(n29051), .Z(n23960) );
  XOR2_X1 U26916 ( .A1(n17518), .A2(n17517), .Z(n17516) );
  XOR2_X1 U26917 ( .A1(n17462), .A2(n19929), .Z(n17517) );
  XOR2_X1 U26918 ( .A1(n23961), .A2(n17520), .Z(n17519) );
  XOR2_X1 U26919 ( .A1(n24050), .A2(n23814), .Z(n17520) );
  OAI21_X1 U26920 ( .A1(n21110), .A2(n21109), .B(n30169), .ZN(n17523) );
  OR2_X1 U26921 ( .A1(n21109), .A2(n30169), .Z(n17524) );
  XOR2_X1 U26922 ( .A1(n22750), .A2(n17528), .Z(n20836) );
  XOR2_X1 U26923 ( .A1(n21378), .A2(Key[67]), .Z(n19370) );
  NAND2_X2 U26926 ( .A1(n21513), .A2(n21512), .ZN(n22322) );
  XOR2_X1 U26933 ( .A1(n10012), .A2(n19905), .Z(n17552) );
  XOR2_X1 U26934 ( .A1(n25234), .A2(n17555), .Z(n17554) );
  INV_X1 U26935 ( .I(n35529), .ZN(n20025) );
  XOR2_X1 U26936 ( .A1(n35255), .A2(n29131), .Z(n29133) );
  INV_X1 U26940 ( .I(n22448), .ZN(n17566) );
  NAND2_X2 U26941 ( .A1(n29193), .A2(n29192), .ZN(n29740) );
  NAND2_X1 U26943 ( .A1(n17989), .A2(n17499), .ZN(n22050) );
  XOR2_X1 U26944 ( .A1(n17580), .A2(n38880), .Z(n17579) );
  XOR2_X1 U26949 ( .A1(n39797), .A2(n30006), .Z(n17595) );
  XOR2_X1 U26950 ( .A1(n31163), .A2(n17603), .Z(n20311) );
  INV_X2 U26951 ( .I(n17604), .ZN(n25557) );
  XOR2_X1 U26952 ( .A1(n35238), .A2(n39172), .Z(n26167) );
  XOR2_X1 U26959 ( .A1(n27466), .A2(n35241), .Z(n17621) );
  NAND2_X2 U26962 ( .A1(n28063), .A2(n28062), .ZN(n29254) );
  XOR2_X1 U26963 ( .A1(n28983), .A2(n19527), .Z(n17627) );
  NAND2_X1 U26965 ( .A1(n906), .A2(n20873), .ZN(n17630) );
  NAND2_X1 U26966 ( .A1(n17636), .A2(n1048), .ZN(n17635) );
  XOR2_X1 U26967 ( .A1(n28306), .A2(n17643), .Z(n17642) );
  INV_X2 U26971 ( .I(n17660), .ZN(n24287) );
  NOR2_X1 U26973 ( .A1(n21780), .A2(n12144), .ZN(n17679) );
  NAND3_X1 U26978 ( .A1(n17687), .A2(n18986), .A3(n27465), .ZN(n17699) );
  XOR2_X1 U26981 ( .A1(Plaintext[129]), .A2(Key[129]), .Z(n20300) );
  XOR2_X1 U26982 ( .A1(n24801), .A2(n17704), .Z(n18556) );
  XOR2_X1 U26983 ( .A1(n16627), .A2(n1557), .Z(n17706) );
  XOR2_X1 U26984 ( .A1(n24991), .A2(n19534), .Z(n17707) );
  INV_X1 U26985 ( .I(Plaintext[146]), .ZN(n17717) );
  XOR2_X1 U26986 ( .A1(n17717), .A2(Key[146]), .Z(n17799) );
  INV_X2 U26988 ( .I(n17726), .ZN(n29781) );
  XOR2_X1 U26990 ( .A1(n467), .A2(n17738), .Z(n17737) );
  XOR2_X1 U26991 ( .A1(n29040), .A2(n13639), .Z(n17738) );
  AND2_X1 U26992 ( .A1(n23550), .A2(n17094), .Z(n17744) );
  XOR2_X1 U26994 ( .A1(n17747), .A2(n29879), .Z(Ciphertext[122]) );
  NAND2_X1 U26996 ( .A1(n39019), .A2(n17286), .ZN(n17750) );
  INV_X2 U27001 ( .I(n17764), .ZN(n25558) );
  INV_X2 U27002 ( .I(n25558), .ZN(n25719) );
  INV_X2 U27003 ( .I(n17767), .ZN(n18841) );
  XOR2_X1 U27007 ( .A1(n8833), .A2(n29801), .Z(n21003) );
  XOR2_X1 U27008 ( .A1(n17776), .A2(n19714), .Z(n20526) );
  AOI21_X1 U27015 ( .A1(n25799), .A2(n31263), .B(n38168), .ZN(n19048) );
  MUX2_X1 U27019 ( .I0(n23221), .I1(n23222), .S(n18236), .Z(n23223) );
  XOR2_X1 U27020 ( .A1(n27830), .A2(n27862), .Z(n17817) );
  XOR2_X1 U27022 ( .A1(n23707), .A2(n19755), .Z(n19344) );
  INV_X2 U27024 ( .I(n17830), .ZN(n23108) );
  OR2_X1 U27025 ( .A1(n20493), .A2(n20492), .Z(n17831) );
  XOR2_X1 U27028 ( .A1(n17836), .A2(n17835), .Z(n17839) );
  XOR2_X1 U27029 ( .A1(n1261), .A2(n25104), .Z(n17835) );
  XOR2_X1 U27035 ( .A1(n17854), .A2(n17853), .Z(n17852) );
  XOR2_X1 U27036 ( .A1(n39682), .A2(n18700), .Z(n17853) );
  XOR2_X1 U27038 ( .A1(n29071), .A2(n20479), .Z(n17859) );
  NOR2_X1 U27039 ( .A1(n17864), .A2(n22240), .ZN(n19180) );
  OAI21_X1 U27040 ( .A1(n24449), .A2(n24453), .B(n17867), .ZN(n24246) );
  XOR2_X1 U27045 ( .A1(n23922), .A2(n37521), .Z(n17872) );
  OAI21_X1 U27046 ( .A1(n18720), .A2(n29494), .B(n29451), .ZN(n28619) );
  XOR2_X1 U27048 ( .A1(n38137), .A2(n19738), .Z(n26339) );
  XOR2_X1 U27051 ( .A1(n17910), .A2(n22764), .Z(n17909) );
  INV_X2 U27052 ( .I(n19959), .ZN(n17911) );
  NOR2_X1 U27053 ( .A1(n24195), .A2(n17911), .ZN(n20734) );
  XOR2_X1 U27056 ( .A1(n17921), .A2(n26183), .Z(n17920) );
  XOR2_X1 U27058 ( .A1(n17937), .A2(n23898), .Z(n23669) );
  XOR2_X1 U27059 ( .A1(n17945), .A2(n17944), .Z(n20573) );
  XOR2_X1 U27060 ( .A1(n844), .A2(n838), .Z(n17944) );
  XOR2_X1 U27061 ( .A1(n26263), .A2(n17946), .Z(n17945) );
  XNOR2_X1 U27062 ( .A1(Plaintext[91]), .A2(Key[91]), .ZN(n17964) );
  XOR2_X1 U27063 ( .A1(n17974), .A2(n19592), .Z(Ciphertext[23]) );
  NAND2_X1 U27066 ( .A1(n29958), .A2(n29959), .ZN(n17983) );
  XOR2_X1 U27067 ( .A1(n1667), .A2(n39136), .Z(n18912) );
  XOR2_X1 U27070 ( .A1(n22509), .A2(n39787), .Z(n17999) );
  AOI21_X1 U27071 ( .A1(n993), .A2(n27137), .B(n19477), .ZN(n18074) );
  NOR2_X1 U27072 ( .A1(n7304), .A2(n1348), .ZN(n18005) );
  XOR2_X1 U27073 ( .A1(n18006), .A2(n39636), .Z(n18410) );
  XOR2_X1 U27074 ( .A1(n18012), .A2(n30016), .Z(n18367) );
  XOR2_X1 U27075 ( .A1(n18012), .A2(n29285), .Z(n26295) );
  XOR2_X1 U27076 ( .A1(n25152), .A2(n18015), .Z(n18014) );
  NAND3_X1 U27081 ( .A1(n20672), .A2(n1173), .A3(n18042), .ZN(n20862) );
  INV_X1 U27082 ( .I(n14387), .ZN(n30215) );
  XOR2_X1 U27085 ( .A1(n18931), .A2(n12707), .Z(n18317) );
  NAND2_X1 U27086 ( .A1(n28717), .A2(n32759), .ZN(n28497) );
  OAI21_X1 U27088 ( .A1(n26122), .A2(n31719), .B(n25903), .ZN(n25905) );
  XOR2_X1 U27089 ( .A1(n27862), .A2(n29295), .Z(n27680) );
  XOR2_X1 U27090 ( .A1(n20602), .A2(n18078), .Z(n20601) );
  XOR2_X1 U27091 ( .A1(n18080), .A2(n18079), .Z(n18078) );
  XOR2_X1 U27092 ( .A1(n23707), .A2(n29661), .Z(n18079) );
  OAI21_X1 U27095 ( .A1(n18084), .A2(n18083), .B(n39709), .ZN(n18082) );
  AND2_X1 U27096 ( .A1(n31570), .A2(n29927), .Z(n18084) );
  NAND2_X1 U27098 ( .A1(n18089), .A2(n18088), .ZN(n28770) );
  AND2_X1 U27105 ( .A1(n37674), .A2(n23155), .Z(n23157) );
  XOR2_X1 U27107 ( .A1(n24012), .A2(n18109), .Z(n19623) );
  XOR2_X1 U27113 ( .A1(n23955), .A2(n24012), .Z(n23717) );
  XOR2_X1 U27115 ( .A1(n1466), .A2(n1468), .Z(n18122) );
  NOR3_X1 U27117 ( .A1(n15338), .A2(n15839), .A3(n21571), .ZN(n20580) );
  XOR2_X1 U27125 ( .A1(n18137), .A2(n39482), .Z(Ciphertext[27]) );
  INV_X2 U27134 ( .I(n18156), .ZN(n20404) );
  XOR2_X1 U27136 ( .A1(Plaintext[5]), .A2(Key[5]), .Z(n18157) );
  XOR2_X1 U27139 ( .A1(Plaintext[63]), .A2(Key[63]), .Z(n18722) );
  XNOR2_X1 U27140 ( .A1(n23879), .A2(n24014), .ZN(n18179) );
  XOR2_X1 U27145 ( .A1(n23730), .A2(n18172), .Z(n21316) );
  XOR2_X1 U27147 ( .A1(n18404), .A2(n18403), .Z(n18178) );
  INV_X2 U27150 ( .I(n18183), .ZN(n26751) );
  XOR2_X1 U27152 ( .A1(n18184), .A2(n29707), .Z(Ciphertext[90]) );
  OAI22_X1 U27153 ( .A1(n29706), .A2(n29722), .B1(n29705), .B2(n29712), .ZN(
        n18184) );
  NAND2_X1 U27156 ( .A1(n18952), .A2(n18951), .ZN(n18950) );
  NAND3_X2 U27159 ( .A1(n22014), .A2(n22012), .A3(n22013), .ZN(n22790) );
  NOR2_X1 U27162 ( .A1(n19367), .A2(n25558), .ZN(n19236) );
  XNOR2_X1 U27163 ( .A1(n19983), .A2(n19984), .ZN(n19714) );
  NAND2_X2 U27164 ( .A1(n18208), .A2(n28903), .ZN(n29548) );
  NAND3_X1 U27165 ( .A1(n28902), .A2(n18720), .A3(n29491), .ZN(n18208) );
  XOR2_X1 U27170 ( .A1(n26403), .A2(n26407), .Z(n25986) );
  AND2_X1 U27171 ( .A1(n23484), .A2(n22493), .Z(n20992) );
  OR2_X1 U27179 ( .A1(n29682), .A2(n33128), .Z(n18945) );
  XOR2_X1 U27182 ( .A1(n18243), .A2(n1724), .Z(Ciphertext[81]) );
  XOR2_X1 U27185 ( .A1(n22699), .A2(n22715), .Z(n18255) );
  NOR2_X1 U27189 ( .A1(n19347), .A2(n29717), .ZN(n29706) );
  BUF_X2 U27190 ( .I(n21753), .Z(n18266) );
  XOR2_X1 U27191 ( .A1(n26366), .A2(n26398), .Z(n18267) );
  NAND2_X1 U27192 ( .A1(n21698), .A2(n19709), .ZN(n19036) );
  OAI22_X1 U27196 ( .A1(n27584), .A2(n27585), .B1(n31955), .B2(n27586), .ZN(
        n27591) );
  XOR2_X1 U27198 ( .A1(n5836), .A2(n22418), .Z(n22421) );
  XNOR2_X1 U27201 ( .A1(n24011), .A2(n29718), .ZN(n20973) );
  XOR2_X1 U27203 ( .A1(n29042), .A2(n38290), .Z(n18319) );
  NAND2_X2 U27205 ( .A1(n24438), .A2(n24437), .ZN(n25290) );
  XOR2_X1 U27207 ( .A1(n36886), .A2(n19152), .Z(n22495) );
  NAND2_X1 U27211 ( .A1(n29617), .A2(n29612), .ZN(n18306) );
  OAI21_X1 U27214 ( .A1(n30031), .A2(n30030), .B(n18313), .ZN(Ciphertext[142])
         );
  XOR2_X1 U27219 ( .A1(n25166), .A2(n24697), .Z(n18327) );
  XOR2_X1 U27222 ( .A1(n26142), .A2(n17551), .Z(n18335) );
  INV_X2 U27226 ( .I(n18345), .ZN(n24465) );
  INV_X2 U27228 ( .I(n7705), .ZN(n25647) );
  XOR2_X1 U27231 ( .A1(n26508), .A2(n18367), .Z(n18366) );
  NAND2_X1 U27233 ( .A1(n13336), .A2(n12392), .ZN(n18386) );
  NOR3_X1 U27235 ( .A1(n39574), .A2(n28233), .A3(n18392), .ZN(n27062) );
  NAND2_X1 U27236 ( .A1(n24504), .A2(n6977), .ZN(n18394) );
  NAND2_X2 U27238 ( .A1(n25458), .A2(n25457), .ZN(n26020) );
  XOR2_X1 U27239 ( .A1(n23937), .A2(n23330), .Z(n18403) );
  XOR2_X1 U27240 ( .A1(n14638), .A2(n29299), .Z(n18405) );
  XOR2_X1 U27242 ( .A1(n23985), .A2(n18410), .Z(n18427) );
  XOR2_X1 U27243 ( .A1(n18422), .A2(n25044), .Z(n18421) );
  XOR2_X1 U27244 ( .A1(n13342), .A2(n24927), .Z(n18422) );
  XOR2_X1 U27245 ( .A1(n25043), .A2(n25042), .Z(n18423) );
  INV_X2 U27248 ( .I(n24202), .ZN(n18907) );
  XOR2_X1 U27253 ( .A1(n27042), .A2(n760), .Z(n18449) );
  XOR2_X1 U27256 ( .A1(n39631), .A2(n28953), .Z(n28954) );
  NAND2_X1 U27259 ( .A1(n18484), .A2(n24229), .ZN(n24230) );
  OAI21_X1 U27260 ( .A1(n20133), .A2(n11820), .B(n18488), .ZN(n27185) );
  XOR2_X1 U27263 ( .A1(n31941), .A2(n26541), .Z(n26431) );
  XOR2_X1 U27265 ( .A1(n18526), .A2(n28806), .Z(n18491) );
  OAI21_X1 U27267 ( .A1(n27951), .A2(n12303), .B(n18497), .ZN(n27868) );
  XOR2_X1 U27272 ( .A1(n24930), .A2(n19742), .Z(n25720) );
  XOR2_X1 U27273 ( .A1(n9930), .A2(n18523), .Z(n18522) );
  INV_X2 U27274 ( .I(n18542), .ZN(n19397) );
  XOR2_X1 U27277 ( .A1(n5021), .A2(n33569), .Z(n18546) );
  NOR2_X1 U27280 ( .A1(n19203), .A2(n18549), .ZN(n26273) );
  XOR2_X1 U27282 ( .A1(n18554), .A2(n20329), .Z(Ciphertext[158]) );
  XOR2_X1 U27285 ( .A1(n25317), .A2(n25028), .Z(n18557) );
  XOR2_X1 U27287 ( .A1(Plaintext[75]), .A2(Key[75]), .Z(n19496) );
  XOR2_X1 U27291 ( .A1(n12690), .A2(n18579), .Z(n18578) );
  XNOR2_X1 U27295 ( .A1(Plaintext[51]), .A2(Key[51]), .ZN(n18585) );
  XOR2_X1 U27304 ( .A1(n26532), .A2(n19721), .Z(n18609) );
  NOR2_X1 U27305 ( .A1(n38142), .A2(n29284), .ZN(n18610) );
  XOR2_X1 U27308 ( .A1(n23778), .A2(n29920), .Z(n18612) );
  XOR2_X1 U27310 ( .A1(n14386), .A2(n23834), .Z(n18620) );
  XOR2_X1 U27313 ( .A1(n22500), .A2(n18635), .Z(n18634) );
  XOR2_X1 U27315 ( .A1(n25208), .A2(n18643), .Z(n18642) );
  NOR2_X1 U27316 ( .A1(n11411), .A2(n4116), .ZN(n18645) );
  NAND2_X1 U27318 ( .A1(n18659), .A2(n29581), .ZN(n18658) );
  NAND2_X1 U27319 ( .A1(n28843), .A2(n39830), .ZN(n18659) );
  NAND2_X1 U27320 ( .A1(n13508), .A2(n28758), .ZN(n19796) );
  NAND2_X1 U27323 ( .A1(n23006), .A2(n18679), .ZN(n23007) );
  XOR2_X1 U27324 ( .A1(n18692), .A2(n18690), .Z(n19954) );
  XOR2_X1 U27325 ( .A1(n22728), .A2(n18691), .Z(n18690) );
  XOR2_X1 U27326 ( .A1(n20335), .A2(n22580), .Z(n18692) );
  XOR2_X1 U27328 ( .A1(n20976), .A2(n19720), .Z(n27161) );
  XOR2_X1 U27330 ( .A1(Plaintext[62]), .A2(Key[62]), .Z(n18723) );
  XOR2_X1 U27331 ( .A1(n27556), .A2(n27853), .Z(n18709) );
  INV_X1 U27332 ( .I(n26804), .ZN(n18719) );
  INV_X2 U27333 ( .I(n18723), .ZN(n20266) );
  NAND2_X2 U27334 ( .A1(n18726), .A2(n18725), .ZN(n29574) );
  XOR2_X1 U27336 ( .A1(n18738), .A2(n18735), .Z(n18741) );
  XOR2_X1 U27337 ( .A1(n18737), .A2(n18736), .Z(n18735) );
  NOR2_X1 U27343 ( .A1(n22797), .A2(n18750), .ZN(n20109) );
  XOR2_X1 U27345 ( .A1(n20698), .A2(n29394), .Z(n18764) );
  XOR2_X1 U27347 ( .A1(Plaintext[48]), .A2(Key[48]), .Z(n18774) );
  INV_X2 U27348 ( .I(n18774), .ZN(n21684) );
  OAI21_X1 U27350 ( .A1(n19434), .A2(n21882), .B(n18784), .ZN(n21884) );
  AND2_X1 U27356 ( .A1(n29672), .A2(n29684), .Z(n18793) );
  XOR2_X1 U27358 ( .A1(n26254), .A2(n18797), .Z(n18796) );
  XOR2_X1 U27359 ( .A1(n26244), .A2(n26349), .Z(n18797) );
  XOR2_X1 U27360 ( .A1(n27802), .A2(n30085), .Z(n18800) );
  NAND3_X1 U27361 ( .A1(n39048), .A2(n31626), .A3(n17791), .ZN(n25705) );
  NAND2_X1 U27362 ( .A1(n27247), .A2(n7973), .ZN(n20455) );
  XOR2_X1 U27363 ( .A1(n18811), .A2(n14571), .Z(n20196) );
  XOR2_X1 U27364 ( .A1(n7549), .A2(n30063), .Z(n18817) );
  XOR2_X1 U27366 ( .A1(n23829), .A2(n29003), .Z(n18828) );
  MUX2_X1 U27367 ( .I0(n10118), .I1(n30117), .S(n30109), .Z(n30118) );
  XOR2_X1 U27369 ( .A1(n22700), .A2(n18834), .Z(n18833) );
  XOR2_X1 U27376 ( .A1(n18846), .A2(n18847), .Z(n28132) );
  XOR2_X1 U27378 ( .A1(n844), .A2(n1237), .Z(n18852) );
  XOR2_X1 U27380 ( .A1(Plaintext[188]), .A2(Key[188]), .Z(n21722) );
  XOR2_X1 U27388 ( .A1(n33194), .A2(n29399), .Z(n18887) );
  MUX2_X1 U27389 ( .I0(n23295), .I1(n23294), .S(n35001), .Z(n18890) );
  XOR2_X1 U27390 ( .A1(n39348), .A2(n13639), .Z(n28876) );
  NAND2_X1 U27393 ( .A1(n18897), .A2(n29981), .ZN(n29965) );
  AOI21_X1 U27395 ( .A1(n31512), .A2(n29980), .B(n18897), .ZN(n19143) );
  XOR2_X1 U27397 ( .A1(n17653), .A2(n29808), .Z(n18898) );
  XOR2_X1 U27401 ( .A1(n28982), .A2(n19583), .Z(n18905) );
  XOR2_X1 U27402 ( .A1(n18211), .A2(n19681), .Z(n24711) );
  XOR2_X1 U27403 ( .A1(n18914), .A2(n18911), .Z(n23102) );
  XOR2_X1 U27404 ( .A1(n18913), .A2(n18912), .Z(n18911) );
  XOR2_X1 U27405 ( .A1(n22443), .A2(n22453), .Z(n18913) );
  XOR2_X1 U27409 ( .A1(n23734), .A2(n23733), .Z(n18921) );
  XOR2_X1 U27413 ( .A1(n25009), .A2(n20592), .Z(n18930) );
  XOR2_X1 U27414 ( .A1(n26163), .A2(n29325), .Z(n18934) );
  XOR2_X1 U27415 ( .A1(n23813), .A2(n23915), .Z(n18935) );
  XOR2_X1 U27416 ( .A1(n20753), .A2(n18943), .Z(n18942) );
  NAND2_X1 U27420 ( .A1(n23532), .A2(n6217), .ZN(n23222) );
  INV_X2 U27424 ( .I(n18968), .ZN(n21928) );
  XOR2_X1 U27427 ( .A1(n23598), .A2(n18977), .Z(n18976) );
  XOR2_X1 U27428 ( .A1(n37701), .A2(n30203), .Z(n18977) );
  MUX2_X1 U27429 ( .I0(n1299), .I1(n23516), .S(n12396), .Z(n23520) );
  NOR2_X1 U27430 ( .A1(n18985), .A2(n37758), .ZN(n18984) );
  NAND2_X1 U27431 ( .A1(n31663), .A2(n28661), .ZN(n18985) );
  XOR2_X1 U27434 ( .A1(n15930), .A2(n18993), .Z(n18992) );
  INV_X2 U27436 ( .I(n19001), .ZN(n23149) );
  INV_X2 U27437 ( .I(n19008), .ZN(n19599) );
  XOR2_X1 U27438 ( .A1(n28858), .A2(n28859), .Z(n19008) );
  XOR2_X1 U27442 ( .A1(n21201), .A2(n22579), .Z(n19015) );
  XOR2_X1 U27446 ( .A1(n26370), .A2(n19019), .Z(n19018) );
  XOR2_X1 U27449 ( .A1(n25240), .A2(n29920), .Z(n19022) );
  XOR2_X1 U27450 ( .A1(n334), .A2(n19940), .Z(n19025) );
  XOR2_X1 U27452 ( .A1(n19031), .A2(n30120), .Z(Ciphertext[160]) );
  NAND2_X1 U27453 ( .A1(n19709), .A2(n18266), .ZN(n21392) );
  NOR2_X1 U27454 ( .A1(n19416), .A2(n18266), .ZN(n21541) );
  NAND2_X1 U27455 ( .A1(n26988), .A2(n19045), .ZN(n26991) );
  XOR2_X1 U27457 ( .A1(n34564), .A2(n19613), .Z(n20069) );
  XOR2_X1 U27459 ( .A1(n518), .A2(n37357), .Z(n19155) );
  XOR2_X1 U27464 ( .A1(n19067), .A2(n28898), .Z(n19066) );
  XOR2_X1 U27465 ( .A1(n29242), .A2(n1719), .Z(n19078) );
  NAND2_X1 U27467 ( .A1(n19084), .A2(n21770), .ZN(n21771) );
  NOR2_X1 U27469 ( .A1(n38142), .A2(n19085), .ZN(n29267) );
  NAND3_X1 U27470 ( .A1(n19091), .A2(n21465), .A3(n34922), .ZN(n20750) );
  XOR2_X1 U27472 ( .A1(n24061), .A2(n14668), .Z(n24063) );
  XOR2_X1 U27473 ( .A1(n24005), .A2(n14668), .Z(n24007) );
  NAND2_X1 U27474 ( .A1(n19097), .A2(n29929), .ZN(n29918) );
  XOR2_X1 U27476 ( .A1(n26224), .A2(n26207), .Z(n19099) );
  XOR2_X1 U27478 ( .A1(n24068), .A2(n19101), .Z(n19100) );
  XOR2_X1 U27479 ( .A1(n24064), .A2(n19102), .Z(n19101) );
  MUX2_X1 U27482 ( .I0(n24704), .I1(n24705), .S(n38674), .Z(n24706) );
  XOR2_X1 U27486 ( .A1(n29254), .A2(n19721), .Z(n19126) );
  NAND2_X2 U27487 ( .A1(n19129), .A2(n19130), .ZN(n29339) );
  NAND2_X1 U27488 ( .A1(n21285), .A2(n105), .ZN(n19312) );
  XOR2_X1 U27490 ( .A1(n19138), .A2(n1735), .Z(Ciphertext[126]) );
  XOR2_X1 U27491 ( .A1(n11974), .A2(n29295), .Z(n19145) );
  XOR2_X1 U27495 ( .A1(n25315), .A2(n19155), .Z(n19154) );
  NOR2_X1 U27496 ( .A1(n19157), .A2(n29410), .ZN(n20132) );
  XOR2_X1 U27497 ( .A1(n29818), .A2(n1737), .Z(n19160) );
  AOI21_X1 U27498 ( .A1(n19164), .A2(n30252), .B(n31529), .ZN(n19163) );
  INV_X2 U27500 ( .I(n19170), .ZN(n28237) );
  XOR2_X1 U27502 ( .A1(n19185), .A2(n19182), .Z(n27964) );
  XOR2_X1 U27503 ( .A1(n19184), .A2(n19183), .Z(n19182) );
  XOR2_X1 U27504 ( .A1(n34332), .A2(n27862), .Z(n19184) );
  XOR2_X1 U27505 ( .A1(n27565), .A2(n27500), .Z(n19185) );
  XOR2_X1 U27506 ( .A1(n11923), .A2(n16618), .Z(n19186) );
  XOR2_X1 U27507 ( .A1(n9701), .A2(n25196), .Z(n19187) );
  INV_X2 U27509 ( .I(n19955), .ZN(n25606) );
  XOR2_X1 U27510 ( .A1(n22713), .A2(n19201), .Z(n19200) );
  NAND2_X1 U27514 ( .A1(n27272), .A2(n35228), .ZN(n19300) );
  XOR2_X1 U27515 ( .A1(n27532), .A2(n35229), .Z(n19213) );
  NOR2_X1 U27518 ( .A1(n12672), .A2(n25048), .ZN(n25049) );
  XOR2_X1 U27519 ( .A1(n19824), .A2(n4348), .Z(n19220) );
  NAND2_X1 U27521 ( .A1(n20276), .A2(n33786), .ZN(n23414) );
  NAND2_X2 U27522 ( .A1(n20059), .A2(n20062), .ZN(n26594) );
  NOR2_X1 U27529 ( .A1(n27279), .A2(n21144), .ZN(n19456) );
  NOR2_X1 U27530 ( .A1(n33538), .A2(n23516), .ZN(n19249) );
  XOR2_X1 U27531 ( .A1(n22693), .A2(n21994), .Z(n22004) );
  XOR2_X1 U27532 ( .A1(n38641), .A2(n38993), .Z(n24858) );
  XOR2_X1 U27533 ( .A1(n25097), .A2(n25096), .Z(n25099) );
  INV_X1 U27534 ( .I(n34914), .ZN(n29583) );
  INV_X2 U27535 ( .I(n19266), .ZN(n20053) );
  XOR2_X1 U27538 ( .A1(n28542), .A2(n19277), .Z(n28883) );
  XOR2_X1 U27539 ( .A1(n28540), .A2(n28541), .Z(n19277) );
  XOR2_X1 U27541 ( .A1(n29140), .A2(n29119), .Z(n20447) );
  NOR2_X1 U27542 ( .A1(n13410), .A2(n25611), .ZN(n25412) );
  NOR2_X1 U27544 ( .A1(n26564), .A2(n26905), .ZN(n19285) );
  XOR2_X1 U27547 ( .A1(n22624), .A2(n22773), .Z(n22514) );
  NAND2_X1 U27548 ( .A1(n37230), .A2(n24241), .ZN(n24242) );
  NAND2_X1 U27551 ( .A1(n15509), .A2(n920), .ZN(n19303) );
  NOR2_X2 U27552 ( .A1(n19305), .A2(n19304), .ZN(n19741) );
  OR2_X1 U27555 ( .A1(n29764), .A2(n19568), .Z(n28862) );
  XOR2_X1 U27556 ( .A1(n28983), .A2(n1375), .Z(n19309) );
  XOR2_X1 U27557 ( .A1(Key[149]), .A2(Plaintext[149]), .Z(n19313) );
  XOR2_X1 U27559 ( .A1(n19316), .A2(n1697), .Z(Ciphertext[140]) );
  NOR2_X1 U27560 ( .A1(n30013), .A2(n30012), .ZN(n19316) );
  BUF_X2 U27563 ( .I(n21735), .Z(n19323) );
  XOR2_X1 U27565 ( .A1(n22676), .A2(n30126), .Z(n20980) );
  NOR2_X1 U27568 ( .A1(n21734), .A2(n21919), .ZN(n19335) );
  BUF_X2 U27569 ( .I(n21875), .Z(n19337) );
  OR2_X1 U27572 ( .A1(n22135), .A2(n11044), .Z(n22018) );
  NOR2_X1 U27573 ( .A1(n29708), .A2(n29721), .ZN(n19347) );
  XOR2_X1 U27579 ( .A1(n22569), .A2(n22449), .Z(n22413) );
  NAND2_X2 U27582 ( .A1(n25344), .A2(n25343), .ZN(n25941) );
  XOR2_X1 U27586 ( .A1(n23693), .A2(n23692), .Z(n24095) );
  BUF_X2 U27589 ( .I(n26921), .Z(n19371) );
  OAI21_X1 U27592 ( .A1(n11171), .A2(n1672), .B(n19385), .ZN(n22010) );
  INV_X1 U27597 ( .I(n29419), .ZN(n19404) );
  NOR2_X1 U27598 ( .A1(n29652), .A2(n17382), .ZN(n19411) );
  OAI21_X2 U27601 ( .A1(n25439), .A2(n19400), .B(n25438), .ZN(n26041) );
  XOR2_X1 U27604 ( .A1(n20747), .A2(n27573), .Z(n19421) );
  NAND2_X1 U27607 ( .A1(n24842), .A2(n24733), .ZN(n19595) );
  INV_X1 U27609 ( .I(n27197), .ZN(n27279) );
  OAI21_X1 U27611 ( .A1(n1240), .A2(n33237), .B(n19439), .ZN(n26095) );
  XOR2_X1 U27613 ( .A1(n21186), .A2(n19445), .Z(n19444) );
  XOR2_X1 U27614 ( .A1(n19446), .A2(n20822), .Z(n20821) );
  INV_X2 U27620 ( .I(n19459), .ZN(n26695) );
  XOR2_X1 U27625 ( .A1(n21381), .A2(Key[140]), .Z(n21608) );
  BUF_X2 U27630 ( .I(n21777), .Z(n19479) );
  XOR2_X1 U27631 ( .A1(n19744), .A2(n19493), .Z(n19492) );
  XOR2_X1 U27633 ( .A1(n18273), .A2(n29808), .Z(n26285) );
  AOI22_X2 U27641 ( .A1(n21543), .A2(n21542), .B1(n21541), .B2(n21540), .ZN(
        n21973) );
  INV_X2 U27643 ( .I(n29721), .ZN(n29712) );
  OAI21_X1 U27645 ( .A1(n25647), .A2(n25429), .B(n19532), .ZN(n25430) );
  XOR2_X1 U27646 ( .A1(n19533), .A2(n26230), .Z(n19867) );
  NOR2_X1 U27647 ( .A1(n7725), .A2(n9188), .ZN(n21256) );
  OAI21_X1 U27648 ( .A1(n17568), .A2(n36839), .B(n14561), .ZN(n22684) );
  OR2_X1 U27649 ( .A1(n30212), .A2(n39083), .Z(n30205) );
  NAND2_X1 U27650 ( .A1(n21812), .A2(n21683), .ZN(n19552) );
  AOI21_X1 U27655 ( .A1(n20725), .A2(n27201), .B(n35895), .ZN(n27076) );
  XOR2_X1 U27656 ( .A1(n16897), .A2(n25086), .Z(n25088) );
  INV_X1 U27657 ( .I(n28546), .ZN(n28322) );
  INV_X2 U27658 ( .I(n19576), .ZN(n24433) );
  XOR2_X1 U27664 ( .A1(n26518), .A2(n26402), .Z(n20260) );
  OR2_X1 U27668 ( .A1(n37183), .A2(n18545), .Z(n20644) );
  XOR2_X1 U27674 ( .A1(n19617), .A2(n15181), .Z(Ciphertext[42]) );
  XOR2_X1 U27676 ( .A1(n26561), .A2(n26562), .Z(n19632) );
  XOR2_X1 U27677 ( .A1(n11721), .A2(n28815), .Z(n19640) );
  XOR2_X1 U27683 ( .A1(n19652), .A2(n20096), .Z(n20095) );
  INV_X1 U27684 ( .I(n12410), .ZN(n20570) );
  INV_X1 U27688 ( .I(n25555), .ZN(n20237) );
  NOR2_X1 U27689 ( .A1(n14453), .A2(n26614), .ZN(n26851) );
  XOR2_X1 U27695 ( .A1(Plaintext[118]), .A2(Key[118]), .Z(n19822) );
  AND2_X1 U27697 ( .A1(n33073), .A2(n35116), .Z(n21661) );
  INV_X1 U27698 ( .I(n24420), .ZN(n24442) );
  INV_X2 U27699 ( .I(n21752), .ZN(n19709) );
  OAI21_X1 U27701 ( .A1(n452), .A2(n10120), .B(n7278), .ZN(n21626) );
  XOR2_X1 U27702 ( .A1(Key[135]), .A2(Plaintext[135]), .Z(n21790) );
  NAND2_X1 U27704 ( .A1(n28381), .A2(n28382), .ZN(n28385) );
  XOR2_X1 U27705 ( .A1(n27687), .A2(n19775), .Z(n20096) );
  XOR2_X1 U27709 ( .A1(n26481), .A2(n26438), .Z(n19744) );
  NOR2_X2 U27710 ( .A1(n19747), .A2(n20473), .ZN(n29684) );
  INV_X2 U27712 ( .I(n19764), .ZN(n27969) );
  XOR2_X1 U27716 ( .A1(n19784), .A2(n29476), .Z(Ciphertext[52]) );
  NAND2_X1 U27717 ( .A1(n20809), .A2(n20808), .ZN(n23289) );
  XOR2_X1 U27718 ( .A1(n23691), .A2(n19792), .Z(n23693) );
  XOR2_X1 U27719 ( .A1(n23690), .A2(n39073), .Z(n19792) );
  XOR2_X1 U27720 ( .A1(n26223), .A2(n19799), .Z(n19798) );
  XOR2_X1 U27722 ( .A1(n27829), .A2(n29808), .Z(n20796) );
  XOR2_X1 U27724 ( .A1(n25188), .A2(n25190), .Z(n19809) );
  OAI21_X1 U27727 ( .A1(n22110), .A2(n22111), .B(n133), .ZN(n19812) );
  XOR2_X1 U27728 ( .A1(n27564), .A2(n27799), .Z(n27769) );
  INV_X1 U27729 ( .I(n21875), .ZN(n21696) );
  INV_X2 U27733 ( .I(n19838), .ZN(n20830) );
  INV_X1 U27736 ( .I(n29837), .ZN(n28819) );
  NOR2_X1 U27737 ( .A1(n22184), .A2(n1048), .ZN(n22186) );
  INV_X1 U27740 ( .I(n24683), .ZN(n24774) );
  INV_X2 U27743 ( .I(n21630), .ZN(n21775) );
  OAI21_X2 U27746 ( .A1(n27742), .A2(n27743), .B(n27741), .ZN(n28753) );
  INV_X2 U27747 ( .I(n19867), .ZN(n26974) );
  XOR2_X1 U27749 ( .A1(n9246), .A2(n29680), .Z(n19983) );
  XOR2_X1 U27751 ( .A1(n21142), .A2(n19882), .Z(n19881) );
  XOR2_X1 U27755 ( .A1(n26210), .A2(n26209), .Z(n19900) );
  NAND2_X1 U27756 ( .A1(n20833), .A2(n25945), .ZN(n25946) );
  XOR2_X1 U27757 ( .A1(n18273), .A2(n30150), .Z(n25947) );
  INV_X2 U27762 ( .I(n19920), .ZN(n29642) );
  OAI21_X1 U27765 ( .A1(n13767), .A2(n19924), .B(n1308), .ZN(n19923) );
  BUF_X2 U27766 ( .I(Key[54]), .Z(n19933) );
  OR2_X1 U27770 ( .A1(n21933), .A2(n20476), .Z(n19985) );
  XOR2_X1 U27772 ( .A1(n22433), .A2(n19954), .Z(n22973) );
  INV_X2 U27777 ( .I(n18576), .ZN(n21820) );
  INV_X1 U27778 ( .I(n29624), .ZN(n29608) );
  XOR2_X1 U27779 ( .A1(n27806), .A2(n19988), .Z(n19987) );
  XOR2_X1 U27780 ( .A1(n27749), .A2(n29320), .Z(n19988) );
  NAND2_X2 U27784 ( .A1(n20008), .A2(n20007), .ZN(n25814) );
  NOR3_X1 U27785 ( .A1(n15350), .A2(n22341), .A3(n22342), .ZN(n22343) );
  XOR2_X1 U27786 ( .A1(n29167), .A2(n28868), .Z(n20033) );
  XOR2_X1 U27789 ( .A1(n23876), .A2(n20045), .Z(n20044) );
  INV_X1 U27792 ( .I(n19676), .ZN(n20489) );
  XOR2_X1 U27793 ( .A1(n24047), .A2(n19676), .Z(n23690) );
  INV_X2 U27795 ( .I(n20063), .ZN(n26852) );
  XOR2_X1 U27796 ( .A1(n26254), .A2(n14670), .Z(n20065) );
  INV_X2 U27799 ( .I(n24224), .ZN(n24432) );
  NAND2_X2 U27800 ( .A1(n20090), .A2(n20089), .ZN(n22503) );
  XOR2_X1 U27801 ( .A1(n27800), .A2(n27797), .Z(n20093) );
  XOR2_X1 U27802 ( .A1(n20098), .A2(n20097), .Z(n20858) );
  XOR2_X1 U27803 ( .A1(n26401), .A2(n749), .Z(n20097) );
  XOR2_X1 U27804 ( .A1(n26593), .A2(n26261), .Z(n20101) );
  XOR2_X1 U27807 ( .A1(n26347), .A2(n14568), .Z(n20107) );
  OAI21_X1 U27809 ( .A1(n29491), .A2(n29418), .B(n20113), .ZN(n29419) );
  XOR2_X1 U27810 ( .A1(n26073), .A2(n26059), .Z(n20117) );
  INV_X1 U27811 ( .I(n35273), .ZN(n29604) );
  XOR2_X1 U27812 ( .A1(n20129), .A2(n17275), .Z(Ciphertext[39]) );
  XOR2_X1 U27816 ( .A1(n27607), .A2(n35270), .Z(n20167) );
  INV_X1 U27817 ( .I(n24728), .ZN(n24727) );
  INV_X2 U27819 ( .I(n20194), .ZN(n25695) );
  INV_X2 U27820 ( .I(n20196), .ZN(n24381) );
  XOR2_X1 U27821 ( .A1(Plaintext[110]), .A2(Key[110]), .Z(n21330) );
  XOR2_X1 U27822 ( .A1(n24047), .A2(n20205), .Z(n23871) );
  XOR2_X1 U27823 ( .A1(n23968), .A2(n20205), .Z(n23720) );
  INV_X1 U27824 ( .I(n26207), .ZN(n26472) );
  MUX2_X1 U27828 ( .I0(n22098), .I1(n22099), .S(n32609), .Z(n22105) );
  XOR2_X1 U27834 ( .A1(n20261), .A2(n20262), .Z(n20257) );
  XOR2_X1 U27836 ( .A1(n26487), .A2(n26520), .Z(n20262) );
  XOR2_X1 U27840 ( .A1(n26263), .A2(n25511), .Z(n20268) );
  INV_X2 U27843 ( .I(n33999), .ZN(n21712) );
  XOR2_X1 U27846 ( .A1(n26461), .A2(n26464), .Z(n20279) );
  XOR2_X1 U27847 ( .A1(n18133), .A2(n28776), .Z(n28777) );
  INV_X2 U27852 ( .I(n20300), .ZN(n21506) );
  NOR2_X1 U27855 ( .A1(n30145), .A2(n18588), .ZN(n30147) );
  AOI21_X1 U27856 ( .A1(n30145), .A2(n18588), .B(n34177), .ZN(n30138) );
  NOR2_X2 U27857 ( .A1(n26733), .A2(n26732), .ZN(n27267) );
  XOR2_X1 U27860 ( .A1(n20325), .A2(n20323), .Z(n29941) );
  XOR2_X1 U27861 ( .A1(n29072), .A2(n29003), .Z(n20324) );
  NOR2_X1 U27863 ( .A1(n11851), .A2(n21762), .ZN(n20332) );
  XOR2_X1 U27864 ( .A1(n20333), .A2(n25278), .Z(n25120) );
  INV_X2 U27865 ( .I(n26931), .ZN(n26564) );
  INV_X1 U27869 ( .I(n23861), .ZN(n24020) );
  NAND2_X1 U27870 ( .A1(n20544), .A2(n21779), .ZN(n20348) );
  XOR2_X1 U27871 ( .A1(n16639), .A2(n30065), .Z(n28318) );
  XOR2_X1 U27872 ( .A1(n18180), .A2(n29522), .Z(n26241) );
  INV_X2 U27873 ( .I(n20361), .ZN(n21808) );
  XOR2_X1 U27876 ( .A1(n20365), .A2(n24973), .Z(n25418) );
  XOR2_X1 U27881 ( .A1(n20392), .A2(n30090), .Z(n22501) );
  XOR2_X1 U27883 ( .A1(n27490), .A2(n27819), .Z(n20400) );
  XOR2_X1 U27884 ( .A1(n39295), .A2(n19936), .Z(n20409) );
  XOR2_X1 U27892 ( .A1(n28895), .A2(n28894), .Z(n29344) );
  XOR2_X1 U27894 ( .A1(n38150), .A2(n31548), .Z(n20446) );
  XOR2_X1 U27895 ( .A1(n21284), .A2(n27550), .Z(n20448) );
  XOR2_X1 U27897 ( .A1(n20452), .A2(n18432), .Z(n29132) );
  XOR2_X1 U27898 ( .A1(n20452), .A2(n30170), .Z(n28853) );
  XOR2_X1 U27900 ( .A1(n20452), .A2(n19815), .Z(n28973) );
  NAND2_X1 U27902 ( .A1(n25336), .A2(n25337), .ZN(n20463) );
  XOR2_X1 U27906 ( .A1(Plaintext[24]), .A2(Key[24]), .Z(n21849) );
  XOR2_X1 U27909 ( .A1(n26349), .A2(n20489), .Z(n26526) );
  NAND2_X1 U27910 ( .A1(n37776), .A2(n28380), .ZN(n20497) );
  XOR2_X1 U27911 ( .A1(n21225), .A2(n22673), .Z(n20502) );
  XOR2_X1 U27916 ( .A1(Plaintext[121]), .A2(Key[121]), .Z(n21740) );
  OAI21_X1 U27918 ( .A1(n28028), .A2(n33331), .B(n33307), .ZN(n28029) );
  INV_X2 U27919 ( .I(n20526), .ZN(n24408) );
  XOR2_X1 U27926 ( .A1(n22420), .A2(n22421), .Z(n20555) );
  INV_X2 U27927 ( .I(n20555), .ZN(n23089) );
  XOR2_X1 U27929 ( .A1(Plaintext[136]), .A2(Key[136]), .Z(n21791) );
  XOR2_X1 U27931 ( .A1(n20559), .A2(n19925), .Z(Ciphertext[13]) );
  XOR2_X1 U27933 ( .A1(n25191), .A2(n662), .Z(n20571) );
  NAND2_X1 U27935 ( .A1(n547), .A2(n21571), .ZN(n20593) );
  XOR2_X1 U27936 ( .A1(Plaintext[70]), .A2(Key[70]), .Z(n20694) );
  XNOR2_X1 U27938 ( .A1(n21426), .A2(Key[1]), .ZN(n20596) );
  INV_X2 U27939 ( .I(n20601), .ZN(n24241) );
  NAND2_X1 U27947 ( .A1(n23075), .A2(n23076), .ZN(n20625) );
  NAND2_X1 U27949 ( .A1(n23210), .A2(n20408), .ZN(n20741) );
  XOR2_X1 U27950 ( .A1(n33470), .A2(n27829), .Z(n20641) );
  XOR2_X1 U27953 ( .A1(n20656), .A2(n26377), .Z(n21277) );
  NAND2_X1 U27955 ( .A1(n26607), .A2(n20666), .ZN(n26608) );
  XOR2_X1 U27956 ( .A1(n20675), .A2(n28579), .Z(n20674) );
  INV_X2 U27957 ( .I(n20677), .ZN(n29598) );
  XOR2_X1 U27958 ( .A1(n28829), .A2(n28828), .Z(n20684) );
  INV_X2 U27959 ( .I(n20685), .ZN(n21924) );
  INV_X2 U27961 ( .I(n20694), .ZN(n21810) );
  INV_X2 U27963 ( .I(n20702), .ZN(n21023) );
  XOR2_X1 U27964 ( .A1(n20707), .A2(n29671), .Z(n25143) );
  XOR2_X1 U27965 ( .A1(n17758), .A2(n18700), .Z(n20713) );
  XOR2_X1 U27966 ( .A1(n24063), .A2(n20717), .Z(n20716) );
  XOR2_X1 U27967 ( .A1(n24059), .A2(n19751), .Z(n20717) );
  XOR2_X1 U27969 ( .A1(n27724), .A2(n27766), .Z(n20723) );
  INV_X2 U27970 ( .I(n20726), .ZN(n29455) );
  BUF_X2 U27973 ( .I(n25351), .Z(n25616) );
  OAI21_X2 U27978 ( .A1(n5059), .A2(n27405), .B(n27083), .ZN(n27799) );
  XOR2_X1 U27979 ( .A1(n19770), .A2(n27754), .Z(n20747) );
  OR2_X1 U27983 ( .A1(n26355), .A2(n26354), .Z(n20764) );
  XOR2_X1 U27984 ( .A1(n37044), .A2(n23950), .Z(n20767) );
  MUX2_X1 U27985 ( .I0(n26023), .I1(n20771), .S(n1105), .Z(n20770) );
  XOR2_X1 U27986 ( .A1(Plaintext[81]), .A2(Key[81]), .Z(n21488) );
  XOR2_X1 U27988 ( .A1(n25178), .A2(n20780), .Z(n20779) );
  XOR2_X1 U27989 ( .A1(n25301), .A2(n20781), .Z(n20780) );
  XOR2_X1 U27990 ( .A1(n22490), .A2(n22633), .Z(n20794) );
  XOR2_X1 U27992 ( .A1(n38201), .A2(n20804), .Z(n20803) );
  XNOR2_X1 U27993 ( .A1(Plaintext[58]), .A2(Key[58]), .ZN(n20810) );
  INV_X2 U27995 ( .I(n20821), .ZN(n30049) );
  XOR2_X1 U27996 ( .A1(n29830), .A2(n29834), .Z(n20822) );
  XOR2_X1 U27997 ( .A1(n30733), .A2(n20483), .Z(n20824) );
  NAND3_X1 U27998 ( .A1(n21422), .A2(n275), .A3(n21843), .ZN(n20825) );
  XOR2_X1 U27999 ( .A1(n6727), .A2(n18981), .Z(n20828) );
  XOR2_X1 U28000 ( .A1(n20836), .A2(n22753), .Z(n23129) );
  OAI21_X1 U28001 ( .A1(n21635), .A2(n21942), .B(n19546), .ZN(n21638) );
  INV_X2 U28005 ( .I(n20866), .ZN(n29777) );
  INV_X1 U28006 ( .I(n27389), .ZN(n27291) );
  XOR2_X1 U28008 ( .A1(Plaintext[84]), .A2(Key[84]), .Z(n21880) );
  XOR2_X1 U28009 ( .A1(n26436), .A2(n26435), .Z(n20886) );
  XNOR2_X1 U28010 ( .A1(Plaintext[156]), .A2(Key[156]), .ZN(n20887) );
  XOR2_X1 U28014 ( .A1(Plaintext[158]), .A2(Key[158]), .Z(n21496) );
  XOR2_X1 U28015 ( .A1(n24561), .A2(n20893), .Z(n20892) );
  XOR2_X1 U28016 ( .A1(n7247), .A2(n25274), .Z(n20893) );
  NAND2_X1 U28017 ( .A1(n1404), .A2(n14417), .ZN(n20901) );
  NOR2_X1 U28018 ( .A1(n24419), .A2(n1596), .ZN(n20903) );
  XOR2_X1 U28026 ( .A1(n20939), .A2(n1719), .Z(Ciphertext[105]) );
  INV_X2 U28027 ( .I(n29797), .ZN(n29788) );
  NAND2_X1 U28032 ( .A1(n29797), .A2(n20963), .ZN(n20962) );
  NOR2_X1 U28034 ( .A1(n26800), .A2(n20120), .ZN(n26801) );
  XOR2_X1 U28037 ( .A1(n21009), .A2(n1723), .Z(Ciphertext[102]) );
  INV_X2 U28038 ( .I(n28132), .ZN(n28229) );
  XOR2_X1 U28039 ( .A1(Plaintext[45]), .A2(Key[45]), .Z(n21674) );
  XOR2_X1 U28042 ( .A1(n10560), .A2(n23838), .Z(n23839) );
  XOR2_X1 U28043 ( .A1(n27863), .A2(n29974), .Z(n21044) );
  XOR2_X1 U28045 ( .A1(n25133), .A2(n33208), .Z(n25134) );
  OR2_X1 U28046 ( .A1(n272), .A2(n22875), .Z(n21063) );
  MUX2_X1 U28047 ( .I0(n21065), .I1(n22769), .S(n32228), .Z(n21064) );
  XOR2_X1 U28050 ( .A1(n29125), .A2(n17039), .Z(n21076) );
  XOR2_X1 U28052 ( .A1(n39032), .A2(n37882), .Z(n21086) );
  XOR2_X1 U28053 ( .A1(n36905), .A2(n19903), .Z(n21095) );
  XOR2_X1 U28054 ( .A1(n29145), .A2(n29146), .Z(n21097) );
  INV_X1 U28055 ( .I(n9151), .ZN(n21100) );
  XOR2_X1 U28059 ( .A1(n21134), .A2(n22414), .Z(n21133) );
  NOR2_X1 U28060 ( .A1(n2799), .A2(n954), .ZN(n21135) );
  NOR2_X1 U28061 ( .A1(n29732), .A2(n29754), .ZN(n21146) );
  NAND2_X1 U28062 ( .A1(n29741), .A2(n29754), .ZN(n21147) );
  XOR2_X1 U28065 ( .A1(n21158), .A2(n32218), .Z(Ciphertext[65]) );
  XOR2_X1 U28067 ( .A1(n21162), .A2(n21161), .Z(n29586) );
  XOR2_X1 U28068 ( .A1(n28767), .A2(n28762), .Z(n21161) );
  XOR2_X1 U28074 ( .A1(n29833), .A2(n19758), .Z(n21172) );
  XOR2_X1 U28076 ( .A1(n24417), .A2(n24932), .Z(n21174) );
  XOR2_X1 U28077 ( .A1(n27000), .A2(n27650), .Z(n21176) );
  NAND3_X1 U28080 ( .A1(n37102), .A2(n26695), .A3(n946), .ZN(n21191) );
  XOR2_X1 U28082 ( .A1(n359), .A2(n19649), .Z(n21197) );
  XOR2_X1 U28084 ( .A1(n9074), .A2(n22445), .Z(n21206) );
  NOR2_X1 U28086 ( .A1(n28569), .A2(n3900), .ZN(n28665) );
  XOR2_X1 U28087 ( .A1(n21215), .A2(n22025), .Z(n21217) );
  XOR2_X1 U28088 ( .A1(n21217), .A2(n14673), .Z(n21216) );
  XOR2_X1 U28089 ( .A1(n22462), .A2(n21219), .Z(n21218) );
  XOR2_X1 U28090 ( .A1(n22566), .A2(n22670), .Z(n21219) );
  XOR2_X1 U28091 ( .A1(Plaintext[56]), .A2(Key[56]), .Z(n21805) );
  NAND2_X1 U28093 ( .A1(n7693), .A2(n21231), .ZN(n24621) );
  NAND2_X1 U28094 ( .A1(n24852), .A2(n21231), .ZN(n24854) );
  INV_X2 U28096 ( .I(n21234), .ZN(n30000) );
  XOR2_X1 U28098 ( .A1(n29282), .A2(n25303), .Z(n21252) );
  INV_X1 U28099 ( .I(n22783), .ZN(n22818) );
  XOR2_X1 U28102 ( .A1(n25113), .A2(n21280), .Z(n21279) );
  NAND2_X1 U28103 ( .A1(n21698), .A2(n1353), .ZN(n21701) );
  AOI21_X1 U28105 ( .A1(n21393), .A2(n1353), .B(n19709), .ZN(n21394) );
  NOR2_X1 U28114 ( .A1(n30134), .A2(n37117), .ZN(n30146) );
  OR2_X1 U28115 ( .A1(n29202), .A2(n6938), .Z(n28789) );
  NAND3_X1 U28120 ( .A1(n28191), .A2(n28189), .A3(n16325), .ZN(n27874) );
  NAND2_X1 U28128 ( .A1(n23344), .A2(n23430), .ZN(n23345) );
  INV_X1 U28129 ( .I(n24104), .ZN(n24174) );
  NAND2_X1 U28130 ( .A1(n25726), .A2(n16168), .ZN(n25732) );
  INV_X1 U28131 ( .I(n26172), .ZN(n26173) );
  NOR2_X1 U28132 ( .A1(n21272), .A2(n27165), .ZN(n27166) );
  INV_X1 U28133 ( .I(n8875), .ZN(n27493) );
  XOR2_X1 U28137 ( .A1(Key[119]), .A2(Plaintext[119]), .Z(n21754) );
  XOR2_X1 U28138 ( .A1(Key[115]), .A2(Plaintext[115]), .Z(n21753) );
  XOR2_X1 U28139 ( .A1(Key[117]), .A2(Plaintext[117]), .Z(n21752) );
  XOR2_X1 U28140 ( .A1(Key[87]), .A2(Plaintext[87]), .Z(n21577) );
  INV_X1 U28141 ( .I(Plaintext[85]), .ZN(n21326) );
  XOR2_X1 U28142 ( .A1(n21326), .A2(Key[85]), .Z(n21575) );
  NAND3_X1 U28143 ( .A1(n21593), .A2(n21507), .A3(n21594), .ZN(n21327) );
  XOR2_X1 U28147 ( .A1(Key[111]), .A2(Plaintext[111]), .Z(n21875) );
  XOR2_X1 U28148 ( .A1(Key[113]), .A2(Plaintext[113]), .Z(n21871) );
  INV_X1 U28150 ( .I(n21330), .ZN(n21876) );
  INV_X1 U28151 ( .I(Plaintext[112]), .ZN(n21329) );
  XOR2_X1 U28152 ( .A1(n21329), .A2(Key[112]), .Z(n21872) );
  OAI21_X1 U28153 ( .A1(n21546), .A2(n19395), .B(n21697), .ZN(n21331) );
  XOR2_X1 U28154 ( .A1(Key[107]), .A2(Plaintext[107]), .Z(n21750) );
  INV_X1 U28155 ( .I(Plaintext[102]), .ZN(n21332) );
  INV_X1 U28158 ( .I(Plaintext[40]), .ZN(n21340) );
  XOR2_X1 U28159 ( .A1(n21340), .A2(Key[40]), .Z(n21688) );
  XOR2_X1 U28160 ( .A1(Plaintext[47]), .A2(Key[47]), .Z(n21432) );
  INV_X1 U28161 ( .I(Plaintext[42]), .ZN(n21341) );
  XOR2_X1 U28162 ( .A1(n21341), .A2(Key[42]), .Z(n21857) );
  OAI21_X1 U28163 ( .A1(n33053), .A2(n18174), .B(n21860), .ZN(n21345) );
  XOR2_X1 U28164 ( .A1(Key[43]), .A2(Plaintext[43]), .Z(n21823) );
  INV_X1 U28167 ( .I(Plaintext[25]), .ZN(n21346) );
  INV_X1 U28169 ( .I(Plaintext[27]), .ZN(n21347) );
  XOR2_X1 U28170 ( .A1(n21347), .A2(Key[27]), .Z(n21848) );
  INV_X1 U28174 ( .I(Plaintext[26]), .ZN(n21350) );
  XOR2_X1 U28175 ( .A1(n21350), .A2(Key[26]), .Z(n21846) );
  XOR2_X1 U28176 ( .A1(Key[19]), .A2(Plaintext[19]), .Z(n21841) );
  INV_X1 U28177 ( .I(Plaintext[50]), .ZN(n21351) );
  XOR2_X1 U28178 ( .A1(n21351), .A2(Key[50]), .Z(n21352) );
  XOR2_X1 U28179 ( .A1(Key[53]), .A2(Plaintext[53]), .Z(n21814) );
  XOR2_X1 U28180 ( .A1(Key[52]), .A2(Plaintext[52]), .Z(n21428) );
  INV_X1 U28183 ( .I(Plaintext[35]), .ZN(n21357) );
  XOR2_X1 U28184 ( .A1(n21357), .A2(Key[35]), .Z(n21358) );
  XOR2_X1 U28185 ( .A1(Key[32]), .A2(Plaintext[32]), .Z(n21835) );
  XOR2_X1 U28186 ( .A1(Key[34]), .A2(Plaintext[34]), .Z(n21628) );
  NOR2_X1 U28188 ( .A1(n21665), .A2(n21837), .ZN(n21360) );
  INV_X1 U28189 ( .I(Plaintext[60]), .ZN(n21366) );
  XOR2_X1 U28190 ( .A1(n21366), .A2(Key[60]), .Z(n21818) );
  XOR2_X1 U28191 ( .A1(Key[78]), .A2(Plaintext[78]), .Z(n21368) );
  INV_X1 U28192 ( .I(n21368), .ZN(n21568) );
  INV_X1 U28193 ( .I(Plaintext[83]), .ZN(n21367) );
  XOR2_X1 U28194 ( .A1(n21367), .A2(Key[83]), .Z(n21567) );
  NAND2_X1 U28197 ( .A1(n1350), .A2(n14373), .ZN(n21373) );
  INV_X1 U28198 ( .I(Plaintext[68]), .ZN(n21376) );
  INV_X1 U28200 ( .I(Plaintext[67]), .ZN(n21378) );
  INV_X1 U28201 ( .I(Plaintext[130]), .ZN(n21380) );
  XOR2_X1 U28202 ( .A1(Key[141]), .A2(Plaintext[141]), .Z(n21655) );
  INV_X1 U28203 ( .I(Plaintext[140]), .ZN(n21381) );
  INV_X1 U28204 ( .I(Plaintext[137]), .ZN(n21382) );
  XOR2_X1 U28205 ( .A1(n21382), .A2(Key[137]), .Z(n21792) );
  OAI21_X1 U28207 ( .A1(n7062), .A2(n21787), .B(n18205), .ZN(n21383) );
  INV_X1 U28209 ( .I(Plaintext[125]), .ZN(n21386) );
  XOR2_X1 U28211 ( .A1(Key[122]), .A2(Plaintext[122]), .Z(n21743) );
  INV_X1 U28212 ( .I(Plaintext[124]), .ZN(n21389) );
  XOR2_X1 U28213 ( .A1(n21389), .A2(Key[124]), .Z(n21742) );
  INV_X1 U28214 ( .I(Plaintext[123]), .ZN(n21390) );
  XOR2_X1 U28215 ( .A1(n21390), .A2(Key[123]), .Z(n21741) );
  AOI21_X1 U28216 ( .A1(n21542), .A2(n21392), .B(n19822), .ZN(n21395) );
  XOR2_X1 U28218 ( .A1(Key[170]), .A2(Plaintext[170]), .Z(n21927) );
  INV_X1 U28220 ( .I(Plaintext[181]), .ZN(n21398) );
  XOR2_X1 U28221 ( .A1(n21398), .A2(Key[181]), .Z(n21905) );
  INV_X1 U28222 ( .I(Plaintext[183]), .ZN(n21399) );
  XOR2_X1 U28225 ( .A1(Key[182]), .A2(Plaintext[182]), .Z(n21721) );
  XOR2_X1 U28228 ( .A1(Key[184]), .A2(Plaintext[184]), .Z(n21641) );
  NAND2_X1 U28229 ( .A1(n21782), .A2(n35116), .ZN(n21402) );
  INV_X1 U28230 ( .I(Plaintext[152]), .ZN(n21403) );
  XOR2_X1 U28231 ( .A1(n21403), .A2(Key[152]), .Z(n21602) );
  XOR2_X1 U28232 ( .A1(Key[154]), .A2(Plaintext[154]), .Z(n21951) );
  INV_X1 U28233 ( .I(n32664), .ZN(n21405) );
  NAND2_X1 U28236 ( .A1(n21782), .A2(n32664), .ZN(n21406) );
  INV_X1 U28237 ( .I(Plaintext[162]), .ZN(n21407) );
  XOR2_X1 U28238 ( .A1(n21407), .A2(Key[162]), .Z(n21630) );
  XOR2_X1 U28239 ( .A1(Key[165]), .A2(Plaintext[165]), .Z(n21777) );
  INV_X1 U28240 ( .I(Plaintext[163]), .ZN(n21408) );
  INV_X1 U28241 ( .I(Plaintext[167]), .ZN(n21409) );
  XOR2_X1 U28242 ( .A1(n21409), .A2(Key[167]), .Z(n21937) );
  XOR2_X1 U28243 ( .A1(Key[166]), .A2(Plaintext[166]), .Z(n21776) );
  NAND2_X1 U28246 ( .A1(n21862), .A2(n18143), .ZN(n21417) );
  INV_X1 U28250 ( .I(Plaintext[1]), .ZN(n21426) );
  XOR2_X1 U28251 ( .A1(Key[0]), .A2(Plaintext[0]), .Z(n21735) );
  AOI21_X1 U28254 ( .A1(n21808), .A2(n21692), .B(n38241), .ZN(n21438) );
  INV_X1 U28257 ( .I(n21460), .ZN(n22118) );
  INV_X1 U28258 ( .I(n21459), .ZN(n22117) );
  NOR2_X1 U28259 ( .A1(n21756), .A2(n19337), .ZN(n21454) );
  NOR2_X1 U28260 ( .A1(n21546), .A2(n21756), .ZN(n21457) );
  NOR2_X1 U28261 ( .A1(n21697), .A2(n19650), .ZN(n21456) );
  NOR2_X1 U28262 ( .A1(n19647), .A2(n21401), .ZN(n21464) );
  NOR2_X1 U28263 ( .A1(n21644), .A2(n21462), .ZN(n21463) );
  NOR2_X1 U28264 ( .A1(n14837), .A2(n21923), .ZN(n21468) );
  NOR2_X1 U28265 ( .A1(n37612), .A2(n21724), .ZN(n21467) );
  NAND2_X1 U28269 ( .A1(n21485), .A2(n32544), .ZN(n21486) );
  MUX2_X1 U28270 ( .I0(n17209), .I1(n21893), .S(n21892), .Z(n21491) );
  NAND2_X1 U28272 ( .A1(n21806), .A2(n21492), .ZN(n21493) );
  INV_X2 U28273 ( .I(n21496), .ZN(n21944) );
  INV_X1 U28274 ( .I(n21770), .ZN(n21635) );
  NOR2_X1 U28276 ( .A1(n21507), .A2(n19434), .ZN(n21508) );
  NAND2_X1 U28279 ( .A1(n21476), .A2(n19543), .ZN(n21519) );
  NAND2_X1 U28280 ( .A1(n1157), .A2(n39192), .ZN(n21532) );
  MUX2_X1 U28282 ( .I0(n21532), .I1(n21531), .S(n18417), .Z(n21534) );
  NAND2_X1 U28283 ( .A1(n21539), .A2(n21699), .ZN(n21540) );
  OAI22_X1 U28285 ( .A1(n21872), .A2(n21756), .B1(n21546), .B2(n19337), .ZN(
        n21548) );
  NAND2_X1 U28286 ( .A1(n21696), .A2(n21695), .ZN(n21547) );
  OAI21_X2 U28287 ( .A1(n21549), .A2(n21548), .B(n21547), .ZN(n22047) );
  NAND2_X1 U28288 ( .A1(n293), .A2(n21111), .ZN(n21556) );
  NOR2_X1 U28289 ( .A1(n21575), .A2(n21883), .ZN(n21881) );
  OAI21_X2 U28290 ( .A1(n21598), .A2(n21597), .B(n21596), .ZN(n22170) );
  NOR2_X1 U28292 ( .A1(n21782), .A2(n35116), .ZN(n21604) );
  NOR2_X1 U28293 ( .A1(n4342), .A2(n15697), .ZN(n21616) );
  INV_X1 U28294 ( .I(n21612), .ZN(n21610) );
  AOI22_X1 U28299 ( .A1(n21624), .A2(n21900), .B1(n21623), .B2(n21840), .ZN(
        n21625) );
  OAI21_X1 U28300 ( .A1(n21939), .A2(n19350), .B(n21632), .ZN(n21633) );
  NOR2_X1 U28301 ( .A1(n16128), .A2(n21770), .ZN(n21639) );
  NAND2_X1 U28303 ( .A1(n21401), .A2(n39650), .ZN(n21642) );
  NOR2_X1 U28305 ( .A1(n21645), .A2(n21909), .ZN(n21646) );
  OAI21_X1 U28306 ( .A1(n21720), .A2(n21646), .B(n21910), .ZN(n21647) );
  NOR2_X1 U28315 ( .A1(n21813), .A2(n21684), .ZN(n21685) );
  NAND2_X1 U28318 ( .A1(n21699), .A2(n19822), .ZN(n21700) );
  MUX2_X1 U28319 ( .I0(n21701), .I1(n21700), .S(n21702), .Z(n21705) );
  NAND2_X1 U28320 ( .A1(n21886), .A2(n15338), .ZN(n21706) );
  OAI21_X1 U28321 ( .A1(n21748), .A2(n1157), .B(n39192), .ZN(n21711) );
  NAND2_X1 U28322 ( .A1(n21711), .A2(n19542), .ZN(n21717) );
  NOR2_X1 U28323 ( .A1(n21748), .A2(n21712), .ZN(n21714) );
  INV_X1 U28325 ( .I(n21732), .ZN(n21733) );
  NAND2_X1 U28326 ( .A1(n670), .A2(n21111), .ZN(n21737) );
  OAI22_X1 U28327 ( .A1(n21737), .A2(n18412), .B1(n21736), .B2(n19323), .ZN(
        n21738) );
  NOR2_X1 U28328 ( .A1(n1157), .A2(n19287), .ZN(n21745) );
  MUX2_X1 U28329 ( .I0(n694), .I1(n18266), .S(n19416), .Z(n21755) );
  NAND2_X1 U28330 ( .A1(n21874), .A2(n21756), .ZN(n21760) );
  NOR2_X1 U28331 ( .A1(n1692), .A2(n19337), .ZN(n21758) );
  NAND2_X1 U28332 ( .A1(n21872), .A2(n21756), .ZN(n21757) );
  NAND2_X1 U28335 ( .A1(n20923), .A2(n32138), .ZN(n21772) );
  MUX2_X1 U28336 ( .I0(n21772), .I1(n21771), .S(n21944), .Z(n21773) );
  NAND2_X1 U28339 ( .A1(n9759), .A2(n18205), .ZN(n21793) );
  AOI21_X1 U28340 ( .A1(n21794), .A2(n21793), .B(n16945), .ZN(n21795) );
  INV_X1 U28341 ( .I(n22034), .ZN(n21799) );
  NOR2_X1 U28342 ( .A1(n21799), .A2(n22246), .ZN(n21800) );
  NAND2_X1 U28343 ( .A1(n21980), .A2(n22300), .ZN(n21801) );
  NAND2_X1 U28344 ( .A1(n22039), .A2(n22038), .ZN(n21803) );
  NAND2_X1 U28346 ( .A1(n1345), .A2(n1693), .ZN(n21809) );
  OAI21_X1 U28347 ( .A1(n13632), .A2(n21816), .B(n21815), .ZN(n21829) );
  NAND2_X1 U28348 ( .A1(n21821), .A2(n22146), .ZN(n21827) );
  NAND2_X1 U28350 ( .A1(n21830), .A2(n11344), .ZN(n21831) );
  NOR2_X1 U28354 ( .A1(n21857), .A2(n21861), .ZN(n21859) );
  OAI21_X1 U28355 ( .A1(n21862), .A2(n21861), .B(n21860), .ZN(n21863) );
  NAND2_X1 U28356 ( .A1(n22241), .A2(n1047), .ZN(n21865) );
  XOR2_X1 U28357 ( .A1(n7055), .A2(n22528), .Z(n21866) );
  AOI21_X1 U28361 ( .A1(n21877), .A2(n19395), .B(n21876), .ZN(n21878) );
  NOR2_X1 U28362 ( .A1(n2533), .A2(n21889), .ZN(n21890) );
  NOR2_X1 U28363 ( .A1(n19647), .A2(n21909), .ZN(n21906) );
  NOR2_X1 U28364 ( .A1(n21908), .A2(n21401), .ZN(n21911) );
  NAND2_X1 U28367 ( .A1(n32164), .A2(n20003), .ZN(n21931) );
  NOR2_X1 U28368 ( .A1(n14769), .A2(n20003), .ZN(n21934) );
  OAI21_X1 U28369 ( .A1(n6722), .A2(n22130), .B(n22282), .ZN(n21957) );
  INV_X1 U28370 ( .I(n21945), .ZN(n21947) );
  NAND2_X2 U28371 ( .A1(n21953), .A2(n21952), .ZN(n22281) );
  NOR2_X1 U28372 ( .A1(n22282), .A2(n19486), .ZN(n21954) );
  INV_X1 U28374 ( .I(n21963), .ZN(n21960) );
  NAND2_X1 U28375 ( .A1(n22281), .A2(n22189), .ZN(n21964) );
  NOR2_X1 U28378 ( .A1(n22344), .A2(n22342), .ZN(n21986) );
  NAND3_X1 U28380 ( .A1(n19471), .A2(n21990), .A3(n32313), .ZN(n21993) );
  NAND3_X1 U28381 ( .A1(n22265), .A2(n33623), .A3(n22266), .ZN(n21998) );
  NOR2_X1 U28382 ( .A1(n32259), .A2(n22267), .ZN(n21997) );
  INV_X1 U28383 ( .I(n22644), .ZN(n21999) );
  XOR2_X1 U28385 ( .A1(n22002), .A2(n22001), .Z(n22003) );
  NAND3_X1 U28389 ( .A1(n22204), .A2(n9685), .A3(n19837), .ZN(n22013) );
  NAND2_X1 U28391 ( .A1(n9736), .A2(n22100), .ZN(n22060) );
  NOR2_X1 U28392 ( .A1(n22268), .A2(n22266), .ZN(n22072) );
  OAI21_X1 U28393 ( .A1(n22140), .A2(n18854), .B(n9265), .ZN(n22078) );
  NOR2_X1 U28394 ( .A1(n22246), .A2(n37938), .ZN(n22077) );
  NAND2_X1 U28395 ( .A1(n19471), .A2(n14139), .ZN(n22081) );
  XOR2_X1 U28396 ( .A1(n22583), .A2(n29562), .Z(n22082) );
  NOR2_X1 U28398 ( .A1(n22356), .A2(n22353), .ZN(n22093) );
  NAND2_X1 U28399 ( .A1(n22334), .A2(n22100), .ZN(n22099) );
  NAND2_X1 U28401 ( .A1(n22172), .A2(n19873), .ZN(n22106) );
  NOR2_X1 U28402 ( .A1(n22108), .A2(n22184), .ZN(n22110) );
  NAND2_X1 U28403 ( .A1(n1049), .A2(n1334), .ZN(n22115) );
  NAND3_X1 U28404 ( .A1(n22118), .A2(n22117), .A3(n22116), .ZN(n22121) );
  INV_X1 U28405 ( .I(n22119), .ZN(n22120) );
  OAI22_X1 U28406 ( .A1(n22265), .A2(n22122), .B1(n22121), .B2(n22120), .ZN(
        n22123) );
  NAND2_X1 U28411 ( .A1(n22985), .A2(n35288), .ZN(n22168) );
  NAND3_X1 U28412 ( .A1(n22225), .A2(n35618), .A3(n22365), .ZN(n22159) );
  NOR2_X1 U28414 ( .A1(n22165), .A2(n196), .ZN(n22166) );
  XOR2_X1 U28415 ( .A1(n22485), .A2(n29399), .Z(n22167) );
  XOR2_X1 U28417 ( .A1(n22610), .A2(n31576), .Z(n22195) );
  NOR2_X1 U28418 ( .A1(n22282), .A2(n22281), .ZN(n22192) );
  XOR2_X1 U28419 ( .A1(n22459), .A2(n3953), .Z(n22201) );
  NAND2_X1 U28423 ( .A1(n22216), .A2(n9938), .ZN(n22217) );
  XOR2_X1 U28424 ( .A1(n22439), .A2(n28910), .Z(n22231) );
  XOR2_X1 U28425 ( .A1(n22452), .A2(n22231), .Z(n22232) );
  XOR2_X1 U28427 ( .A1(n22391), .A2(n22761), .Z(n22279) );
  MUX2_X1 U28430 ( .I0(n22309), .I1(n22308), .S(n14024), .Z(n22312) );
  NAND3_X1 U28431 ( .A1(n1335), .A2(n22310), .A3(n31651), .ZN(n22311) );
  XOR2_X1 U28433 ( .A1(n22634), .A2(n29805), .Z(n22370) );
  INV_X1 U28434 ( .I(n22376), .ZN(n22374) );
  INV_X1 U28435 ( .I(n22375), .ZN(n22373) );
  NAND3_X1 U28436 ( .A1(n22374), .A2(n18270), .A3(n22373), .ZN(n22378) );
  OAI21_X1 U28437 ( .A1(n22376), .A2(n22375), .B(n23591), .ZN(n22377) );
  NAND2_X1 U28438 ( .A1(n22378), .A2(n22377), .ZN(n22379) );
  XOR2_X1 U28439 ( .A1(n359), .A2(n30114), .Z(n22383) );
  XOR2_X1 U28440 ( .A1(n22729), .A2(n22749), .Z(n22384) );
  XOR2_X1 U28441 ( .A1(n22567), .A2(n22384), .Z(n22385) );
  XOR2_X1 U28442 ( .A1(n22715), .A2(n29206), .Z(n22393) );
  XOR2_X1 U28444 ( .A1(n34678), .A2(n19875), .Z(n22394) );
  INV_X1 U28447 ( .I(n22398), .ZN(n22404) );
  OAI22_X1 U28448 ( .A1(n22404), .A2(n22403), .B1(n22402), .B2(n22401), .ZN(
        n22405) );
  NAND3_X1 U28449 ( .A1(n23103), .A2(n23104), .A3(n903), .ZN(n22407) );
  XOR2_X1 U28450 ( .A1(n11541), .A2(n19825), .Z(n22409) );
  XOR2_X1 U28453 ( .A1(n22700), .A2(n22550), .Z(n22415) );
  XOR2_X1 U28454 ( .A1(n9874), .A2(n28821), .Z(n22414) );
  XOR2_X1 U28455 ( .A1(n9116), .A2(n19874), .Z(n22417) );
  XOR2_X1 U28456 ( .A1(n16226), .A2(n19721), .Z(n22418) );
  XOR2_X1 U28458 ( .A1(n31863), .A2(n30950), .Z(n22422) );
  XOR2_X1 U28459 ( .A1(n22422), .A2(n22755), .Z(n22425) );
  XOR2_X1 U28462 ( .A1(n31576), .A2(n22563), .Z(n22426) );
  XOR2_X1 U28464 ( .A1(n22566), .A2(n21215), .Z(n22431) );
  XOR2_X1 U28465 ( .A1(n22432), .A2(n22431), .Z(n22433) );
  XOR2_X1 U28466 ( .A1(n34678), .A2(n29319), .Z(n22436) );
  XOR2_X1 U28467 ( .A1(n39804), .A2(n29003), .Z(n22442) );
  XOR2_X1 U28468 ( .A1(n36596), .A2(n19903), .Z(n22446) );
  XOR2_X1 U28469 ( .A1(n22643), .A2(n22763), .Z(n22451) );
  XOR2_X1 U28472 ( .A1(n22509), .A2(n19774), .Z(n22469) );
  XOR2_X1 U28473 ( .A1(n18568), .A2(n22580), .Z(n22470) );
  XOR2_X1 U28477 ( .A1(n31339), .A2(n9874), .Z(n22474) );
  XOR2_X1 U28478 ( .A1(n39682), .A2(n19947), .Z(n22478) );
  XOR2_X1 U28479 ( .A1(n9982), .A2(n19897), .Z(n22487) );
  XOR2_X1 U28481 ( .A1(n22575), .A2(n19624), .Z(n22494) );
  MUX2_X1 U28482 ( .I0(n22496), .I1(n36245), .S(n20376), .Z(n22498) );
  XOR2_X1 U28483 ( .A1(n15439), .A2(n29442), .Z(n22505) );
  XOR2_X1 U28484 ( .A1(n34718), .A2(n22562), .Z(n22519) );
  XOR2_X1 U28485 ( .A1(n22583), .A2(n29801), .Z(n22521) );
  XOR2_X1 U28486 ( .A1(n22522), .A2(n22521), .Z(n22523) );
  NAND2_X1 U28487 ( .A1(n15770), .A2(n22890), .ZN(n22526) );
  XOR2_X1 U28490 ( .A1(n37428), .A2(n22582), .Z(n22537) );
  XOR2_X1 U28491 ( .A1(n17195), .A2(n29964), .Z(n22536) );
  XOR2_X1 U28492 ( .A1(n22536), .A2(n22537), .Z(n22538) );
  XOR2_X1 U28494 ( .A1(n20294), .A2(n22544), .Z(n22548) );
  XOR2_X1 U28495 ( .A1(n22546), .A2(n22545), .Z(n22547) );
  XOR2_X1 U28496 ( .A1(n22548), .A2(n22547), .Z(n22853) );
  NAND2_X1 U28498 ( .A1(n19288), .A2(n22928), .ZN(n22558) );
  XOR2_X1 U28499 ( .A1(n22647), .A2(n22621), .Z(n22560) );
  XOR2_X1 U28500 ( .A1(n22610), .A2(n19887), .Z(n22564) );
  XOR2_X1 U28503 ( .A1(n35920), .A2(n19622), .Z(n22576) );
  XOR2_X1 U28504 ( .A1(n22668), .A2(n14309), .Z(n22579) );
  XOR2_X1 U28505 ( .A1(n16798), .A2(n22582), .Z(n22584) );
  XOR2_X1 U28507 ( .A1(n22601), .A2(n2383), .Z(n22602) );
  XOR2_X1 U28508 ( .A1(n36867), .A2(n22610), .Z(n22611) );
  XOR2_X1 U28509 ( .A1(n39804), .A2(n19722), .Z(n22613) );
  XOR2_X1 U28510 ( .A1(n38330), .A2(n19933), .Z(n22617) );
  XOR2_X1 U28511 ( .A1(n19094), .A2(n19894), .Z(n22618) );
  XOR2_X1 U28512 ( .A1(n22629), .A2(n22749), .Z(n22630) );
  XOR2_X1 U28514 ( .A1(n22634), .A2(n19833), .Z(n22636) );
  XOR2_X1 U28515 ( .A1(n39682), .A2(n19913), .Z(n22641) );
  XOR2_X1 U28516 ( .A1(n22645), .A2(n19808), .Z(n22646) );
  XOR2_X1 U28517 ( .A1(n22648), .A2(n29554), .Z(n22649) );
  XOR2_X1 U28518 ( .A1(n17195), .A2(n29538), .Z(n22653) );
  XOR2_X1 U28519 ( .A1(n22659), .A2(n19820), .Z(n22660) );
  XOR2_X1 U28520 ( .A1(n22671), .A2(n22670), .Z(n22673) );
  XOR2_X1 U28524 ( .A1(n3475), .A2(n19910), .Z(n22704) );
  NAND2_X1 U28527 ( .A1(n23012), .A2(n33972), .ZN(n22708) );
  XOR2_X1 U28528 ( .A1(n22715), .A2(n30016), .Z(n22716) );
  XOR2_X1 U28529 ( .A1(n22717), .A2(n22716), .Z(n22718) );
  XOR2_X1 U28530 ( .A1(n22718), .A2(n22719), .Z(n23140) );
  XOR2_X1 U28532 ( .A1(n22778), .A2(n22761), .Z(n22726) );
  XOR2_X1 U28533 ( .A1(n22724), .A2(n19758), .Z(n22725) );
  XOR2_X1 U28534 ( .A1(n22726), .A2(n22725), .Z(n22727) );
  XOR2_X1 U28535 ( .A1(n35559), .A2(n19780), .Z(n22734) );
  XOR2_X1 U28537 ( .A1(n1657), .A2(n30094), .Z(n22737) );
  NAND2_X1 U28540 ( .A1(n23034), .A2(n4682), .ZN(n22746) );
  XOR2_X1 U28541 ( .A1(n38838), .A2(n29463), .Z(n22751) );
  XOR2_X1 U28542 ( .A1(n22752), .A2(n22751), .Z(n22753) );
  XOR2_X1 U28544 ( .A1(n22763), .A2(n19817), .Z(n22764) );
  XOR2_X1 U28545 ( .A1(n22766), .A2(n29476), .Z(n22768) );
  XOR2_X1 U28549 ( .A1(n39682), .A2(n19831), .Z(n22782) );
  NAND2_X1 U28552 ( .A1(n9050), .A2(n59), .ZN(n22797) );
  OAI21_X1 U28554 ( .A1(n22903), .A2(n906), .B(n20872), .ZN(n22815) );
  NAND2_X1 U28555 ( .A1(n19307), .A2(n23028), .ZN(n22817) );
  NAND3_X1 U28560 ( .A1(n23149), .A2(n31838), .A3(n14556), .ZN(n22831) );
  NAND3_X1 U28563 ( .A1(n5702), .A2(n4573), .A3(n22931), .ZN(n22846) );
  NAND2_X1 U28564 ( .A1(n31906), .A2(n17090), .ZN(n22852) );
  NOR2_X1 U28566 ( .A1(n22875), .A2(n19840), .ZN(n22876) );
  INV_X1 U28567 ( .I(n23123), .ZN(n22877) );
  OAI21_X1 U28568 ( .A1(n45), .A2(n23034), .B(n35994), .ZN(n22881) );
  NOR2_X1 U28569 ( .A1(n38173), .A2(n1642), .ZN(n22911) );
  NOR2_X1 U28573 ( .A1(n23189), .A2(n23188), .ZN(n22977) );
  NAND2_X1 U28574 ( .A1(n34419), .A2(n23188), .ZN(n22978) );
  NAND2_X1 U28580 ( .A1(n36829), .A2(n23456), .ZN(n22986) );
  NAND2_X1 U28581 ( .A1(n18762), .A2(n30574), .ZN(n22988) );
  MUX2_X1 U28585 ( .I0(n23071), .I1(n23005), .S(n5976), .Z(n23006) );
  INV_X1 U28587 ( .I(n23479), .ZN(n23017) );
  INV_X1 U28590 ( .I(n121), .ZN(n23026) );
  NAND2_X1 U28593 ( .A1(n18284), .A2(n23458), .ZN(n23040) );
  NAND2_X1 U28595 ( .A1(n23045), .A2(n11658), .ZN(n23046) );
  NAND2_X1 U28596 ( .A1(n9854), .A2(n38542), .ZN(n23049) );
  NAND2_X1 U28597 ( .A1(n33817), .A2(n23159), .ZN(n23050) );
  INV_X1 U28598 ( .I(n23054), .ZN(n23055) );
  NOR2_X1 U28607 ( .A1(n14556), .A2(n31838), .ZN(n23151) );
  NAND2_X1 U28608 ( .A1(n16963), .A2(n36095), .ZN(n23431) );
  AOI21_X1 U28610 ( .A1(n38524), .A2(n23189), .B(n23188), .ZN(n23193) );
  XOR2_X1 U28613 ( .A1(n19649), .A2(n23911), .Z(n23220) );
  NAND3_X1 U28615 ( .A1(n32351), .A2(n17556), .A3(n31644), .ZN(n23218) );
  NAND2_X1 U28617 ( .A1(n23277), .A2(n1629), .ZN(n23228) );
  NAND3_X1 U28620 ( .A1(n23462), .A2(n23458), .A3(n5083), .ZN(n23240) );
  NAND2_X1 U28621 ( .A1(n23420), .A2(n23602), .ZN(n23252) );
  NAND2_X1 U28624 ( .A1(n39001), .A2(n10024), .ZN(n23267) );
  NAND2_X1 U28625 ( .A1(n12093), .A2(n32158), .ZN(n23271) );
  NAND2_X1 U28626 ( .A1(n31332), .A2(n23539), .ZN(n23276) );
  MUX2_X1 U28627 ( .I0(n23534), .I1(n23276), .S(n23538), .Z(n23279) );
  XOR2_X1 U28628 ( .A1(n23846), .A2(n29983), .Z(n23280) );
  NAND3_X1 U28633 ( .A1(n23450), .A2(n38173), .A3(n1642), .ZN(n23291) );
  NAND2_X1 U28635 ( .A1(n18762), .A2(n31586), .ZN(n23295) );
  NAND2_X1 U28636 ( .A1(n1135), .A2(n23293), .ZN(n23294) );
  XOR2_X1 U28639 ( .A1(n23783), .A2(n29879), .Z(n23330) );
  OAI21_X1 U28646 ( .A1(n39214), .A2(n7485), .B(n23367), .ZN(n23368) );
  NAND2_X1 U28649 ( .A1(n39300), .A2(n23502), .ZN(n23375) );
  XOR2_X1 U28650 ( .A1(n33452), .A2(n19735), .Z(n23378) );
  XOR2_X1 U28651 ( .A1(n32122), .A2(n17462), .Z(n23382) );
  INV_X1 U28653 ( .I(n23548), .ZN(n23386) );
  NOR2_X1 U28659 ( .A1(n30499), .A2(n23401), .ZN(n23403) );
  XOR2_X1 U28660 ( .A1(n23888), .A2(n29666), .Z(n23409) );
  XOR2_X1 U28661 ( .A1(n23734), .A2(n23409), .Z(n23410) );
  XOR2_X1 U28664 ( .A1(n23755), .A2(n29808), .Z(n23428) );
  NAND3_X1 U28665 ( .A1(n33287), .A2(n31661), .A3(n32930), .ZN(n23427) );
  XOR2_X1 U28666 ( .A1(n23717), .A2(n23428), .Z(n23429) );
  AOI21_X1 U28667 ( .A1(n1628), .A2(n3496), .B(n23624), .ZN(n23435) );
  NAND3_X1 U28671 ( .A1(n23484), .A2(n23483), .A3(n9078), .ZN(n23485) );
  NAND2_X1 U28672 ( .A1(n23251), .A2(n23496), .ZN(n23494) );
  NAND4_X1 U28675 ( .A1(n23511), .A2(n11245), .A3(n23510), .A4(n23509), .ZN(
        n23512) );
  XOR2_X1 U28677 ( .A1(n19608), .A2(n30179), .Z(n23549) );
  NAND2_X1 U28678 ( .A1(n23583), .A2(n23582), .ZN(n23584) );
  NOR2_X1 U28680 ( .A1(n12597), .A2(n23602), .ZN(n23603) );
  NAND2_X1 U28683 ( .A1(n35506), .A2(n13305), .ZN(n23630) );
  XOR2_X1 U28685 ( .A1(n32122), .A2(n29831), .Z(n23649) );
  XOR2_X1 U28686 ( .A1(n24070), .A2(n19804), .Z(n23653) );
  XOR2_X1 U28687 ( .A1(n23886), .A2(n19527), .Z(n23656) );
  XOR2_X1 U28690 ( .A1(n24017), .A2(n23665), .Z(n23666) );
  XOR2_X1 U28691 ( .A1(n23955), .A2(n19913), .Z(n23668) );
  XOR2_X1 U28692 ( .A1(n24025), .A2(n19817), .Z(n23672) );
  XOR2_X1 U28694 ( .A1(n238), .A2(n29801), .Z(n23687) );
  XOR2_X1 U28695 ( .A1(n18279), .A2(n29325), .Z(n23689) );
  XOR2_X1 U28696 ( .A1(n18310), .A2(n23728), .Z(n23692) );
  XOR2_X1 U28698 ( .A1(n23698), .A2(n28910), .Z(n23699) );
  XOR2_X1 U28701 ( .A1(n24005), .A2(n19592), .Z(n23713) );
  XOR2_X1 U28702 ( .A1(n24077), .A2(n29474), .Z(n23719) );
  XOR2_X1 U28705 ( .A1(n35942), .A2(n29538), .Z(n23727) );
  XOR2_X1 U28706 ( .A1(n1617), .A2(n23728), .Z(n23813) );
  INV_X1 U28707 ( .I(n24079), .ZN(n23792) );
  XOR2_X1 U28709 ( .A1(n23769), .A2(n19583), .Z(n23733) );
  XOR2_X1 U28710 ( .A1(n23884), .A2(n29707), .Z(n23738) );
  INV_X1 U28712 ( .I(n23972), .ZN(n23742) );
  INV_X1 U28714 ( .I(n23746), .ZN(n23747) );
  INV_X1 U28715 ( .I(n23748), .ZN(n23750) );
  NAND2_X1 U28716 ( .A1(n23750), .A2(n23749), .ZN(n23751) );
  XOR2_X1 U28717 ( .A1(n23757), .A2(n23814), .Z(n23758) );
  XOR2_X1 U28718 ( .A1(n23850), .A2(n23759), .Z(n23760) );
  XOR2_X1 U28719 ( .A1(n23808), .A2(n19877), .Z(n23763) );
  NAND4_X1 U28720 ( .A1(n23767), .A2(n23766), .A3(n23796), .A4(n23765), .ZN(
        n23768) );
  XOR2_X1 U28721 ( .A1(n23769), .A2(n29442), .Z(n23770) );
  XOR2_X1 U28722 ( .A1(n23771), .A2(n23770), .Z(n23772) );
  XOR2_X1 U28723 ( .A1(n23933), .A2(n35942), .Z(n23795) );
  MUX2_X1 U28724 ( .I0(n9822), .I1(n23799), .S(n1125), .Z(n23800) );
  XOR2_X1 U28725 ( .A1(n39209), .A2(n33866), .Z(n23803) );
  NAND2_X1 U28728 ( .A1(n9844), .A2(n12771), .ZN(n23821) );
  OR2_X1 U28729 ( .A1(n23821), .A2(n11265), .Z(n23822) );
  NAND2_X1 U28731 ( .A1(n545), .A2(n19915), .ZN(n23828) );
  XOR2_X1 U28732 ( .A1(n23851), .A2(n30016), .Z(n23834) );
  XOR2_X1 U28733 ( .A1(n35561), .A2(n19831), .Z(n23836) );
  NOR2_X1 U28734 ( .A1(n19880), .A2(n39467), .ZN(n23845) );
  INV_X1 U28735 ( .I(n24061), .ZN(n23838) );
  XOR2_X1 U28736 ( .A1(n23866), .A2(n23842), .Z(n23843) );
  XOR2_X1 U28738 ( .A1(n23846), .A2(n29238), .Z(n23847) );
  XOR2_X1 U28739 ( .A1(n23890), .A2(n19952), .Z(n23849) );
  XOR2_X1 U28740 ( .A1(n19608), .A2(n29206), .Z(n23853) );
  XOR2_X1 U28742 ( .A1(n23861), .A2(n19839), .Z(n23862) );
  XOR2_X1 U28743 ( .A1(n23863), .A2(n23862), .Z(n23864) );
  XOR2_X1 U28744 ( .A1(n33452), .A2(n35702), .Z(n23867) );
  XOR2_X1 U28745 ( .A1(n24075), .A2(n29221), .Z(n23870) );
  XOR2_X1 U28748 ( .A1(n23970), .A2(n19866), .Z(n23879) );
  XOR2_X1 U28749 ( .A1(n24077), .A2(n33672), .Z(n24014) );
  XOR2_X1 U28751 ( .A1(n23988), .A2(n23893), .Z(n23925) );
  XOR2_X1 U28752 ( .A1(n23894), .A2(n19736), .Z(n23895) );
  XOR2_X1 U28753 ( .A1(n23925), .A2(n23895), .Z(n23896) );
  XOR2_X1 U28754 ( .A1(n23897), .A2(n23896), .Z(n23907) );
  XOR2_X1 U28756 ( .A1(n23900), .A2(n30170), .Z(n23901) );
  XOR2_X1 U28757 ( .A1(n23905), .A2(n29319), .Z(n23906) );
  XOR2_X1 U28760 ( .A1(n23609), .A2(n29689), .Z(n23927) );
  XOR2_X1 U28761 ( .A1(n23944), .A2(n23945), .Z(n23949) );
  XOR2_X1 U28762 ( .A1(n23609), .A2(n19780), .Z(n23946) );
  XOR2_X1 U28764 ( .A1(n23973), .A2(n19908), .Z(n23974) );
  XOR2_X1 U28765 ( .A1(n23976), .A2(n29602), .Z(n23977) );
  MUX2_X1 U28766 ( .I0(n24444), .I1(n23983), .S(n24311), .Z(n23994) );
  XOR2_X1 U28769 ( .A1(n23988), .A2(n23987), .Z(n23989) );
  XOR2_X1 U28770 ( .A1(n23989), .A2(n20594), .Z(n23990) );
  XOR2_X1 U28771 ( .A1(n23991), .A2(n23990), .Z(n24420) );
  XOR2_X1 U28776 ( .A1(n24030), .A2(n19885), .Z(n24032) );
  XOR2_X1 U28777 ( .A1(n24036), .A2(n6561), .Z(n24037) );
  XOR2_X1 U28779 ( .A1(n30321), .A2(n19721), .Z(n24042) );
  XOR2_X1 U28780 ( .A1(n24047), .A2(n29295), .Z(n24048) );
  XOR2_X1 U28781 ( .A1(n24052), .A2(n19616), .Z(n24054) );
  INV_X1 U28782 ( .I(n24133), .ZN(n24072) );
  XOR2_X1 U28783 ( .A1(n24076), .A2(n29363), .Z(n24078) );
  NOR3_X1 U28787 ( .A1(n16917), .A2(n24311), .A3(n253), .ZN(n24091) );
  MUX2_X1 U28790 ( .I0(n277), .I1(n24398), .S(n24396), .Z(n24105) );
  INV_X1 U28791 ( .I(n19880), .ZN(n24170) );
  NAND2_X1 U28792 ( .A1(n24105), .A2(n24170), .ZN(n24109) );
  NOR2_X1 U28794 ( .A1(n24168), .A2(n24395), .ZN(n24107) );
  INV_X1 U28797 ( .I(n24410), .ZN(n24111) );
  INV_X1 U28798 ( .I(n24161), .ZN(n24117) );
  MUX2_X1 U28802 ( .I0(n24129), .I1(n24157), .S(n13653), .Z(n24131) );
  NAND2_X1 U28805 ( .A1(n24271), .A2(n18697), .ZN(n24148) );
  XOR2_X1 U28806 ( .A1(n38714), .A2(n19648), .Z(n24150) );
  NOR2_X1 U28807 ( .A1(n6849), .A2(n20537), .ZN(n24163) );
  OAI21_X1 U28808 ( .A1(n19942), .A2(n30897), .B(n802), .ZN(n24193) );
  NAND2_X1 U28809 ( .A1(n35890), .A2(n31452), .ZN(n24194) );
  NAND2_X1 U28813 ( .A1(n24221), .A2(n6839), .ZN(n24222) );
  NAND3_X1 U28823 ( .A1(n19745), .A2(n24267), .A3(n24266), .ZN(n24268) );
  NAND2_X1 U28827 ( .A1(n24300), .A2(n37045), .ZN(n24298) );
  NOR2_X1 U28828 ( .A1(n37267), .A2(n24463), .ZN(n24302) );
  NAND2_X1 U28831 ( .A1(n24419), .A2(n24311), .ZN(n24312) );
  XOR2_X1 U28835 ( .A1(n19817), .A2(n25086), .Z(n24325) );
  NAND4_X1 U28836 ( .A1(n24342), .A2(n24341), .A3(n24339), .A4(n24340), .ZN(
        n24343) );
  NOR2_X1 U28838 ( .A1(n36082), .A2(n4008), .ZN(n24363) );
  NAND3_X1 U28840 ( .A1(n14167), .A2(n24818), .A3(n24824), .ZN(n24388) );
  NAND2_X1 U28841 ( .A1(n24392), .A2(n1283), .ZN(n24393) );
  XOR2_X1 U28845 ( .A1(n39756), .A2(n19761), .Z(n24436) );
  NAND2_X1 U28846 ( .A1(n24606), .A2(n20696), .ZN(n24437) );
  NAND2_X1 U28848 ( .A1(n14491), .A2(n24449), .ZN(n24452) );
  MUX2_X1 U28850 ( .I0(n24452), .I1(n24451), .S(n17871), .Z(n24456) );
  NAND2_X1 U28856 ( .A1(n34123), .A2(n31684), .ZN(n24498) );
  NOR2_X1 U28858 ( .A1(n24876), .A2(n1580), .ZN(n24504) );
  INV_X1 U28862 ( .I(n24530), .ZN(n24531) );
  XOR2_X1 U28866 ( .A1(n24944), .A2(n30248), .Z(n24541) );
  XOR2_X1 U28867 ( .A1(n24542), .A2(n24541), .Z(n24543) );
  XOR2_X1 U28868 ( .A1(n24544), .A2(n24543), .Z(n25395) );
  XOR2_X1 U28869 ( .A1(n9701), .A2(n24942), .Z(n24551) );
  XOR2_X1 U28871 ( .A1(n25218), .A2(n29689), .Z(n24550) );
  XOR2_X1 U28872 ( .A1(n24551), .A2(n24550), .Z(n24552) );
  XOR2_X1 U28875 ( .A1(n17184), .A2(n28910), .Z(n24563) );
  NAND2_X1 U28879 ( .A1(n18788), .A2(n24753), .ZN(n24577) );
  NAND4_X1 U28882 ( .A1(n24585), .A2(n24584), .A3(n24583), .A4(n24582), .ZN(
        n24586) );
  INV_X1 U28888 ( .I(n24625), .ZN(n24626) );
  XOR2_X1 U28889 ( .A1(n1260), .A2(n19583), .Z(n24632) );
  XOR2_X1 U28891 ( .A1(n25247), .A2(n25280), .Z(n24641) );
  XOR2_X1 U28898 ( .A1(n24678), .A2(n19816), .Z(n24679) );
  INV_X1 U28899 ( .I(n24687), .ZN(n24690) );
  XOR2_X1 U28900 ( .A1(n10792), .A2(n18991), .Z(n24697) );
  NAND2_X1 U28901 ( .A1(n16502), .A2(n7769), .ZN(n24705) );
  AOI21_X1 U28902 ( .A1(n24723), .A2(n5056), .B(n24721), .ZN(n24725) );
  XOR2_X1 U28904 ( .A1(n38581), .A2(n25071), .Z(n24801) );
  NOR2_X1 U28905 ( .A1(n14939), .A2(n19868), .ZN(n24815) );
  NOR3_X1 U28906 ( .A1(n24821), .A2(n24820), .A3(n7529), .ZN(n24822) );
  INV_X1 U28910 ( .I(n24843), .ZN(n24844) );
  NAND2_X1 U28911 ( .A1(n24844), .A2(n4973), .ZN(n24845) );
  XOR2_X1 U28915 ( .A1(n24857), .A2(n24858), .Z(n24859) );
  XOR2_X1 U28916 ( .A1(n25030), .A2(n18270), .Z(n24860) );
  MUX2_X1 U28917 ( .I0(n37477), .I1(n24869), .S(n19901), .Z(n24871) );
  NAND2_X1 U28919 ( .A1(n24885), .A2(n24884), .ZN(n24886) );
  XOR2_X1 U28920 ( .A1(n25113), .A2(n19801), .Z(n24891) );
  INV_X1 U28922 ( .I(n24904), .ZN(n24905) );
  XOR2_X1 U28923 ( .A1(n6727), .A2(n19763), .Z(n24913) );
  XOR2_X1 U28924 ( .A1(n24914), .A2(n24913), .Z(n24915) );
  XOR2_X1 U28925 ( .A1(n25085), .A2(n29978), .Z(n24918) );
  XOR2_X1 U28926 ( .A1(n38950), .A2(n19890), .Z(n24919) );
  XOR2_X1 U28927 ( .A1(n16627), .A2(n19732), .Z(n24923) );
  XOR2_X1 U28929 ( .A1(n16864), .A2(n29970), .Z(n24940) );
  XOR2_X1 U28930 ( .A1(n25232), .A2(n24940), .Z(n24941) );
  XOR2_X1 U28931 ( .A1(n25238), .A2(n29875), .Z(n24945) );
  XOR2_X1 U28933 ( .A1(n25226), .A2(n19774), .Z(n24947) );
  XOR2_X1 U28935 ( .A1(n24953), .A2(n24952), .Z(n24954) );
  XOR2_X1 U28936 ( .A1(n24955), .A2(n24954), .Z(n25157) );
  XOR2_X1 U28938 ( .A1(n25203), .A2(n29887), .Z(n24960) );
  XOR2_X1 U28939 ( .A1(n10792), .A2(n29363), .Z(n24966) );
  OAI21_X2 U28940 ( .A1(n24968), .A2(n24967), .B(n19574), .ZN(n26388) );
  XOR2_X1 U28941 ( .A1(n25215), .A2(n19883), .Z(n24971) );
  XOR2_X1 U28942 ( .A1(n24972), .A2(n24971), .Z(n24973) );
  XOR2_X1 U28943 ( .A1(n25218), .A2(n29983), .Z(n24975) );
  XOR2_X1 U28944 ( .A1(n24976), .A2(n24975), .Z(n24977) );
  XOR2_X1 U28949 ( .A1(n25026), .A2(n30150), .Z(n24988) );
  XOR2_X1 U28950 ( .A1(n39146), .A2(n32195), .Z(n24989) );
  XOR2_X1 U28951 ( .A1(n25167), .A2(n24989), .Z(n24990) );
  INV_X1 U28952 ( .I(n25546), .ZN(n25482) );
  XOR2_X1 U28953 ( .A1(n24991), .A2(n19721), .Z(n24992) );
  XOR2_X1 U28954 ( .A1(n25237), .A2(n5208), .Z(n25004) );
  XOR2_X1 U28955 ( .A1(n33208), .A2(n25090), .Z(n25005) );
  MUX2_X1 U28956 ( .I0(n31580), .I1(n12825), .S(n18704), .Z(n25012) );
  XOR2_X1 U28957 ( .A1(n25014), .A2(n19903), .Z(n25015) );
  INV_X1 U28959 ( .I(n25018), .ZN(n25020) );
  NOR3_X1 U28960 ( .A1(n25020), .A2(n38631), .A3(n25019), .ZN(n25021) );
  XOR2_X1 U28961 ( .A1(n25104), .A2(n30114), .Z(n25023) );
  XOR2_X1 U28962 ( .A1(n25024), .A2(n30104), .Z(n25025) );
  XOR2_X1 U28963 ( .A1(n25026), .A2(n19866), .Z(n25027) );
  XOR2_X1 U28964 ( .A1(n25226), .A2(n19839), .Z(n25034) );
  NOR2_X1 U28965 ( .A1(n34010), .A2(n25307), .ZN(n25036) );
  XOR2_X1 U28966 ( .A1(n39491), .A2(n29506), .Z(n25041) );
  INV_X1 U28967 ( .I(n25047), .ZN(n25051) );
  AOI22_X1 U28968 ( .A1(n25051), .A2(n36634), .B1(n32488), .B2(n25049), .ZN(
        n25056) );
  INV_X1 U28969 ( .I(n25052), .ZN(n25054) );
  NAND2_X1 U28970 ( .A1(n25054), .A2(n25053), .ZN(n25055) );
  XOR2_X1 U28972 ( .A1(n25259), .A2(n19407), .Z(n25059) );
  XOR2_X1 U28973 ( .A1(n25060), .A2(n25059), .Z(n25061) );
  XOR2_X1 U28976 ( .A1(n36075), .A2(n29514), .Z(n25064) );
  XOR2_X1 U28977 ( .A1(n25326), .A2(n25064), .Z(n25065) );
  NOR2_X1 U28979 ( .A1(n21302), .A2(n955), .ZN(n25073) );
  XOR2_X1 U28980 ( .A1(n6185), .A2(n25175), .Z(n25078) );
  XOR2_X1 U28981 ( .A1(n25076), .A2(n29371), .Z(n25077) );
  XOR2_X1 U28983 ( .A1(n10199), .A2(n25090), .Z(n25092) );
  XOR2_X1 U28984 ( .A1(n35900), .A2(n19825), .Z(n25094) );
  XOR2_X1 U28985 ( .A1(n39491), .A2(n29357), .Z(n25098) );
  XOR2_X1 U28986 ( .A1(n25098), .A2(n25099), .Z(n25101) );
  INV_X1 U28987 ( .I(n25106), .ZN(n25582) );
  XOR2_X1 U28991 ( .A1(n29680), .A2(n38665), .Z(n25119) );
  XOR2_X1 U28992 ( .A1(n25120), .A2(n25119), .Z(n25121) );
  INV_X1 U28994 ( .I(n25123), .ZN(n25125) );
  XOR2_X1 U28995 ( .A1(n25283), .A2(n25149), .Z(n25129) );
  XOR2_X1 U28996 ( .A1(n25127), .A2(n19877), .Z(n25128) );
  XOR2_X1 U28998 ( .A1(n25155), .A2(n35996), .Z(n25135) );
  XOR2_X1 U28999 ( .A1(n25135), .A2(n25134), .Z(n25139) );
  XOR2_X1 U29000 ( .A1(n39756), .A2(n19738), .Z(n25137) );
  XOR2_X1 U29002 ( .A1(n30865), .A2(n33216), .Z(n25187) );
  XOR2_X1 U29003 ( .A1(n25189), .A2(n1561), .Z(n25190) );
  XOR2_X1 U29005 ( .A1(n35707), .A2(n30169), .Z(n25207) );
  XOR2_X1 U29006 ( .A1(n39491), .A2(n30203), .Z(n25213) );
  XOR2_X1 U29009 ( .A1(n25231), .A2(n25232), .Z(n25236) );
  XOR2_X1 U29010 ( .A1(n24417), .A2(n19860), .Z(n25233) );
  XOR2_X1 U29011 ( .A1(n25234), .A2(n25233), .Z(n25235) );
  XOR2_X1 U29012 ( .A1(n16900), .A2(n28968), .Z(n25276) );
  XOR2_X1 U29013 ( .A1(n25280), .A2(n30120), .Z(n25281) );
  XOR2_X1 U29014 ( .A1(n38714), .A2(n29522), .Z(n25304) );
  XOR2_X1 U29015 ( .A1(n39491), .A2(n29647), .Z(n25320) );
  OAI21_X1 U29016 ( .A1(n25552), .A2(n19478), .B(n18704), .ZN(n25336) );
  NOR2_X1 U29019 ( .A1(n12533), .A2(n31509), .ZN(n25341) );
  NAND2_X1 U29023 ( .A1(n25352), .A2(n25386), .ZN(n25354) );
  NAND3_X1 U29025 ( .A1(n14410), .A2(n6731), .A3(n9132), .ZN(n25358) );
  MUX2_X1 U29027 ( .I0(n25371), .I1(n25370), .S(n25886), .Z(n25377) );
  NAND2_X1 U29030 ( .A1(n25394), .A2(n19398), .ZN(n25397) );
  XOR2_X1 U29032 ( .A1(n3413), .A2(n29920), .Z(n25407) );
  NAND2_X1 U29036 ( .A1(n38183), .A2(n20614), .ZN(n25425) );
  NAND3_X1 U29038 ( .A1(n952), .A2(n15406), .A3(n17029), .ZN(n25428) );
  NAND2_X1 U29039 ( .A1(n8070), .A2(n1252), .ZN(n25776) );
  NAND2_X1 U29040 ( .A1(n25429), .A2(n33946), .ZN(n25431) );
  INV_X1 U29042 ( .I(n25717), .ZN(n25437) );
  NAND2_X1 U29043 ( .A1(n25869), .A2(n18162), .ZN(n25440) );
  NAND3_X1 U29045 ( .A1(n25614), .A2(n36816), .A3(n25575), .ZN(n25451) );
  NOR2_X1 U29047 ( .A1(n1109), .A2(n25577), .ZN(n25456) );
  OAI21_X1 U29048 ( .A1(n12404), .A2(n25381), .B(n1109), .ZN(n25457) );
  NOR2_X1 U29050 ( .A1(n25469), .A2(n1257), .ZN(n25471) );
  NAND2_X1 U29057 ( .A1(n19548), .A2(n4603), .ZN(n25503) );
  NOR2_X1 U29058 ( .A1(n26015), .A2(n25899), .ZN(n25507) );
  NAND2_X1 U29059 ( .A1(n25507), .A2(n1522), .ZN(n25508) );
  XOR2_X1 U29060 ( .A1(n26418), .A2(n19820), .Z(n25511) );
  NAND2_X1 U29067 ( .A1(n12825), .A2(n14602), .ZN(n25549) );
  AOI21_X1 U29069 ( .A1(n25554), .A2(n19581), .B(n12825), .ZN(n25555) );
  NOR3_X1 U29070 ( .A1(n14410), .A2(n6731), .A3(n9132), .ZN(n25560) );
  NOR2_X1 U29075 ( .A1(n37553), .A2(n1552), .ZN(n25592) );
  XOR2_X1 U29076 ( .A1(n26532), .A2(n19613), .Z(n25594) );
  NAND3_X1 U29084 ( .A1(n20856), .A2(n14082), .A3(n25642), .ZN(n25643) );
  NAND2_X1 U29087 ( .A1(n20456), .A2(n36226), .ZN(n25657) );
  NAND2_X1 U29088 ( .A1(n30436), .A2(n3356), .ZN(n25658) );
  NOR2_X1 U29091 ( .A1(n25677), .A2(n25674), .ZN(n25675) );
  NAND2_X1 U29095 ( .A1(n25712), .A2(n8304), .ZN(n25713) );
  MUX2_X1 U29098 ( .I0(n25730), .I1(n25729), .S(n5166), .Z(n25731) );
  XOR2_X1 U29099 ( .A1(n25734), .A2(n25735), .Z(n25736) );
  NAND2_X1 U29100 ( .A1(n9530), .A2(n19793), .ZN(n25741) );
  NAND2_X1 U29104 ( .A1(n11807), .A2(n25760), .ZN(n25762) );
  NAND3_X1 U29105 ( .A1(n9855), .A2(n37683), .A3(n1012), .ZN(n25761) );
  INV_X1 U29106 ( .I(n25775), .ZN(n25780) );
  NAND3_X1 U29107 ( .A1(n25778), .A2(n25777), .A3(n25776), .ZN(n25779) );
  NAND2_X1 U29109 ( .A1(n25747), .A2(n26020), .ZN(n25787) );
  AOI21_X1 U29113 ( .A1(n25966), .A2(n25804), .B(n25803), .ZN(n25805) );
  INV_X1 U29114 ( .I(n26186), .ZN(n25810) );
  NOR2_X1 U29115 ( .A1(n25814), .A2(n25813), .ZN(n25815) );
  NAND2_X1 U29119 ( .A1(n25830), .A2(n31340), .ZN(n25831) );
  NOR2_X1 U29123 ( .A1(n34898), .A2(n26075), .ZN(n25840) );
  NAND2_X1 U29128 ( .A1(n1522), .A2(n1098), .ZN(n25902) );
  NAND2_X1 U29129 ( .A1(n26015), .A2(n25899), .ZN(n25901) );
  MUX2_X1 U29130 ( .I0(n25902), .I1(n25901), .S(n33327), .Z(n25907) );
  MUX2_X1 U29134 ( .I0(n25911), .I1(n25910), .S(n26004), .Z(n25914) );
  XOR2_X1 U29135 ( .A1(n5084), .A2(n29661), .Z(n25930) );
  NOR3_X1 U29137 ( .A1(n25345), .A2(n26063), .A3(n25941), .ZN(n25942) );
  NAND3_X1 U29138 ( .A1(n11807), .A2(n15283), .A3(n9883), .ZN(n25950) );
  NAND3_X1 U29139 ( .A1(n37683), .A2(n34898), .A3(n15283), .ZN(n25949) );
  NAND2_X1 U29141 ( .A1(n25961), .A2(n25965), .ZN(n25964) );
  NAND2_X1 U29144 ( .A1(n25966), .A2(n26028), .ZN(n25967) );
  INV_X1 U29146 ( .I(n26034), .ZN(n25982) );
  NOR2_X1 U29149 ( .A1(n26237), .A2(n30883), .ZN(n26036) );
  NOR2_X1 U29150 ( .A1(n1100), .A2(n26034), .ZN(n26239) );
  XOR2_X1 U29151 ( .A1(n26259), .A2(n26548), .Z(n26085) );
  XOR2_X1 U29154 ( .A1(n26319), .A2(n30253), .Z(n26141) );
  NOR2_X1 U29155 ( .A1(n37524), .A2(n12066), .ZN(n26149) );
  XOR2_X1 U29156 ( .A1(n1502), .A2(n19780), .Z(n26144) );
  XOR2_X1 U29157 ( .A1(n26411), .A2(n26144), .Z(n26147) );
  AOI21_X1 U29159 ( .A1(n36262), .A2(n10902), .B(n26151), .ZN(n26152) );
  XOR2_X1 U29161 ( .A1(n4622), .A2(n19947), .Z(n26156) );
  XOR2_X1 U29162 ( .A1(n2150), .A2(n19860), .Z(n26162) );
  INV_X1 U29163 ( .I(n26995), .ZN(n26878) );
  NAND2_X1 U29164 ( .A1(n20981), .A2(n27081), .ZN(n26195) );
  XOR2_X1 U29165 ( .A1(n26568), .A2(n35202), .Z(n26168) );
  XOR2_X1 U29166 ( .A1(n38279), .A2(n26168), .Z(n26171) );
  XOR2_X1 U29168 ( .A1(n26568), .A2(n26231), .Z(n26192) );
  XOR2_X1 U29169 ( .A1(n38896), .A2(n18270), .Z(n26191) );
  NAND2_X1 U29170 ( .A1(n33254), .A2(n37201), .ZN(n26196) );
  XOR2_X1 U29172 ( .A1(n26198), .A2(n26567), .Z(n26200) );
  XOR2_X1 U29176 ( .A1(n26291), .A2(n29319), .Z(n26206) );
  XOR2_X1 U29177 ( .A1(n26531), .A2(n19534), .Z(n26209) );
  NAND2_X1 U29178 ( .A1(n26212), .A2(n5908), .ZN(n26217) );
  NAND3_X1 U29179 ( .A1(n9868), .A2(n26214), .A3(n26213), .ZN(n26216) );
  XOR2_X1 U29182 ( .A1(n26388), .A2(n30120), .Z(n26232) );
  XOR2_X1 U29185 ( .A1(n39129), .A2(n19616), .Z(n26243) );
  MUX2_X1 U29186 ( .I0(n13181), .I1(n38483), .S(n26876), .Z(n26251) );
  XOR2_X1 U29187 ( .A1(n26404), .A2(n19890), .Z(n26260) );
  NOR2_X1 U29188 ( .A1(n948), .A2(n26269), .ZN(n26268) );
  XOR2_X1 U29189 ( .A1(n36958), .A2(n29657), .Z(n26277) );
  INV_X1 U29190 ( .I(n26379), .ZN(n26280) );
  XOR2_X1 U29191 ( .A1(n334), .A2(n26476), .Z(n26282) );
  XOR2_X1 U29192 ( .A1(n12839), .A2(n19770), .Z(n26281) );
  XOR2_X1 U29194 ( .A1(n2150), .A2(n19839), .Z(n26289) );
  NAND2_X1 U29195 ( .A1(n13392), .A2(n26764), .ZN(n26299) );
  XOR2_X1 U29196 ( .A1(n12649), .A2(n29394), .Z(n26292) );
  XOR2_X1 U29197 ( .A1(n26293), .A2(n26292), .Z(n26294) );
  XOR2_X1 U29200 ( .A1(n26386), .A2(n26465), .Z(n26297) );
  XOR2_X1 U29201 ( .A1(n26591), .A2(n19527), .Z(n26301) );
  XOR2_X1 U29205 ( .A1(n26510), .A2(n19950), .Z(n26310) );
  XOR2_X1 U29206 ( .A1(n26311), .A2(n26310), .Z(n26312) );
  NAND2_X1 U29208 ( .A1(n36424), .A2(n14377), .ZN(n26316) );
  XOR2_X1 U29210 ( .A1(n9989), .A2(n26504), .Z(n26317) );
  XOR2_X1 U29211 ( .A1(n26438), .A2(n26584), .Z(n26574) );
  XOR2_X1 U29212 ( .A1(n26319), .A2(n29295), .Z(n26320) );
  XOR2_X1 U29213 ( .A1(n26320), .A2(n26574), .Z(n26321) );
  NAND2_X1 U29215 ( .A1(n26331), .A2(n7460), .ZN(n26327) );
  NAND4_X1 U29216 ( .A1(n19574), .A2(n19775), .A3(n26327), .A4(n26326), .ZN(
        n26333) );
  NAND3_X1 U29217 ( .A1(n26331), .A2(n26330), .A3(n7460), .ZN(n26332) );
  XOR2_X1 U29218 ( .A1(n26441), .A2(n9085), .Z(n26336) );
  XOR2_X1 U29221 ( .A1(n29554), .A2(n1010), .Z(n26343) );
  XOR2_X1 U29222 ( .A1(n30090), .A2(n34148), .Z(n26350) );
  NAND2_X1 U29224 ( .A1(n1091), .A2(n26804), .ZN(n26355) );
  XOR2_X1 U29225 ( .A1(n26359), .A2(n29879), .Z(n26360) );
  XOR2_X1 U29229 ( .A1(n26456), .A2(n26404), .Z(n26371) );
  XOR2_X1 U29231 ( .A1(n26380), .A2(n26518), .Z(n26383) );
  XOR2_X1 U29232 ( .A1(n26381), .A2(n26542), .Z(n26382) );
  XOR2_X1 U29233 ( .A1(n26383), .A2(n26382), .Z(n26384) );
  INV_X1 U29234 ( .I(n26389), .ZN(n26390) );
  XOR2_X1 U29235 ( .A1(n26391), .A2(n35702), .Z(n26392) );
  XOR2_X1 U29236 ( .A1(n26404), .A2(n19936), .Z(n26405) );
  XOR2_X1 U29238 ( .A1(n26456), .A2(n26407), .Z(n26409) );
  NAND2_X1 U29243 ( .A1(n26424), .A2(n19762), .ZN(n26426) );
  XOR2_X1 U29249 ( .A1(n35251), .A2(n26460), .Z(n26461) );
  XOR2_X1 U29250 ( .A1(n1238), .A2(n29538), .Z(n26464) );
  XOR2_X1 U29252 ( .A1(n34469), .A2(n19804), .Z(n26473) );
  XOR2_X1 U29253 ( .A1(n19450), .A2(n19622), .Z(n26493) );
  XOR2_X1 U29254 ( .A1(n35251), .A2(n19801), .Z(n26496) );
  NAND2_X1 U29256 ( .A1(n26936), .A2(n26937), .ZN(n26515) );
  XOR2_X1 U29257 ( .A1(n11105), .A2(n19774), .Z(n26536) );
  XOR2_X1 U29258 ( .A1(n39793), .A2(n26542), .Z(n26544) );
  XOR2_X1 U29260 ( .A1(n32464), .A2(n19732), .Z(n26562) );
  INV_X1 U29261 ( .I(n26560), .ZN(n26561) );
  XOR2_X1 U29267 ( .A1(n26599), .A2(n19908), .Z(n26600) );
  INV_X1 U29268 ( .I(n26989), .ZN(n26607) );
  NAND2_X1 U29270 ( .A1(n26692), .A2(n26879), .ZN(n26610) );
  NOR2_X1 U29274 ( .A1(n20223), .A2(n26780), .ZN(n26621) );
  INV_X1 U29280 ( .I(n26929), .ZN(n26636) );
  OAI21_X1 U29288 ( .A1(n35197), .A2(n19442), .B(n14488), .ZN(n26675) );
  MUX2_X1 U29289 ( .I0(n20021), .I1(n26675), .S(n26674), .Z(n26678) );
  NOR2_X1 U29299 ( .A1(n33858), .A2(n26961), .ZN(n26721) );
  NOR2_X1 U29301 ( .A1(n26948), .A2(n39595), .ZN(n26730) );
  NOR3_X1 U29302 ( .A1(n26951), .A2(n26731), .A3(n26730), .ZN(n26732) );
  NAND3_X1 U29304 ( .A1(n17047), .A2(n26740), .A3(n1235), .ZN(n26741) );
  OAI21_X1 U29308 ( .A1(n12755), .A2(n19179), .B(n26760), .ZN(n26762) );
  NOR2_X1 U29310 ( .A1(n26934), .A2(n17993), .ZN(n26776) );
  NAND2_X1 U29313 ( .A1(n866), .A2(n17712), .ZN(n26783) );
  NAND2_X1 U29314 ( .A1(n39564), .A2(n9147), .ZN(n26793) );
  NAND2_X1 U29318 ( .A1(n39823), .A2(n20321), .ZN(n26842) );
  OAI21_X1 U29320 ( .A1(n26849), .A2(n26945), .B(n26848), .ZN(n26850) );
  MUX2_X1 U29321 ( .I0(n26851), .I1(n26850), .S(n20660), .Z(n26853) );
  NAND2_X1 U29325 ( .A1(n30429), .A2(n27138), .ZN(n26887) );
  NOR2_X1 U29326 ( .A1(n26923), .A2(n26922), .ZN(n26897) );
  XOR2_X1 U29327 ( .A1(n19612), .A2(n29474), .Z(n26916) );
  AOI21_X1 U29330 ( .A1(n859), .A2(n26936), .B(n26935), .ZN(n26939) );
  NAND2_X1 U29331 ( .A1(n36477), .A2(n26937), .ZN(n26938) );
  INV_X1 U29334 ( .I(n26955), .ZN(n26956) );
  NAND2_X1 U29335 ( .A1(n26957), .A2(n8103), .ZN(n26958) );
  NAND3_X1 U29336 ( .A1(n27508), .A2(n31287), .A3(n19529), .ZN(n26965) );
  NAND2_X1 U29338 ( .A1(n26981), .A2(n26980), .ZN(n26985) );
  NAND2_X1 U29340 ( .A1(n26992), .A2(n13111), .ZN(n26993) );
  NAND2_X1 U29341 ( .A1(n27108), .A2(n18246), .ZN(n26998) );
  NOR2_X1 U29346 ( .A1(n27044), .A2(n27043), .ZN(n27048) );
  INV_X1 U29347 ( .I(n27045), .ZN(n27047) );
  NOR2_X1 U29349 ( .A1(n27059), .A2(n38571), .ZN(n27060) );
  XOR2_X1 U29351 ( .A1(n38937), .A2(n16613), .Z(n27080) );
  XOR2_X1 U29354 ( .A1(n27362), .A2(n27087), .Z(n27088) );
  XOR2_X1 U29355 ( .A1(n27089), .A2(n27088), .Z(n27481) );
  NAND2_X1 U29357 ( .A1(n27092), .A2(n15276), .ZN(n27094) );
  NAND3_X1 U29358 ( .A1(n20092), .A2(n13992), .A3(n27098), .ZN(n27099) );
  NAND3_X1 U29362 ( .A1(n32697), .A2(n19334), .A3(n18717), .ZN(n27106) );
  NAND3_X1 U29363 ( .A1(n27180), .A2(n1085), .A3(n1478), .ZN(n27109) );
  NAND2_X1 U29364 ( .A1(n27430), .A2(n30986), .ZN(n27121) );
  INV_X1 U29366 ( .I(n27124), .ZN(n27127) );
  INV_X1 U29367 ( .I(n27125), .ZN(n27126) );
  INV_X1 U29368 ( .I(n27139), .ZN(n27143) );
  INV_X1 U29369 ( .I(n27140), .ZN(n27142) );
  NAND4_X1 U29370 ( .A1(n27144), .A2(n27143), .A3(n27142), .A4(n9593), .ZN(
        n27145) );
  NAND2_X1 U29374 ( .A1(n27175), .A2(n33369), .ZN(n27176) );
  NAND3_X1 U29380 ( .A1(n27391), .A2(n35895), .A3(n13699), .ZN(n27203) );
  OAI21_X1 U29383 ( .A1(n37), .A2(n38579), .B(n1448), .ZN(n27215) );
  AOI21_X1 U29385 ( .A1(n28495), .A2(n1427), .B(n7454), .ZN(n27458) );
  INV_X1 U29387 ( .I(n27224), .ZN(n27225) );
  XOR2_X1 U29388 ( .A1(n27592), .A2(n19883), .Z(n27229) );
  XOR2_X1 U29394 ( .A1(n37812), .A2(n30065), .Z(n27302) );
  NAND3_X1 U29395 ( .A1(n14614), .A2(n4434), .A3(n27409), .ZN(n27316) );
  INV_X1 U29398 ( .I(n27334), .ZN(n27335) );
  NAND2_X1 U29401 ( .A1(n19455), .A2(n38571), .ZN(n27353) );
  NAND2_X1 U29403 ( .A1(n33050), .A2(n35228), .ZN(n27369) );
  NAND2_X1 U29407 ( .A1(n27384), .A2(n33336), .ZN(n27386) );
  NOR2_X1 U29408 ( .A1(n27417), .A2(n27416), .ZN(n27419) );
  NAND2_X1 U29413 ( .A1(n4847), .A2(n27449), .ZN(n27451) );
  NAND3_X1 U29414 ( .A1(n27452), .A2(n2923), .A3(n27451), .ZN(n27453) );
  XOR2_X1 U29415 ( .A1(n13289), .A2(n27849), .Z(n27461) );
  XOR2_X1 U29416 ( .A1(n27594), .A2(n27766), .Z(n27463) );
  XOR2_X1 U29417 ( .A1(n27540), .A2(n29970), .Z(n27467) );
  XNOR2_X1 U29418 ( .A1(n27663), .A2(n29711), .ZN(n27471) );
  XOR2_X1 U29420 ( .A1(n29319), .A2(n27815), .Z(n27479) );
  NAND2_X1 U29421 ( .A1(n28124), .A2(n14404), .ZN(n27482) );
  MUX2_X1 U29422 ( .I0(n27486), .I1(n27485), .S(n33335), .Z(n27489) );
  INV_X1 U29423 ( .I(n27487), .ZN(n27488) );
  XOR2_X1 U29424 ( .A1(n4934), .A2(n29879), .Z(n27491) );
  INV_X1 U29425 ( .I(Key[184]), .ZN(n29017) );
  XOR2_X1 U29428 ( .A1(n38205), .A2(n27525), .Z(n27514) );
  INV_X1 U29429 ( .I(n27592), .ZN(n27517) );
  XOR2_X1 U29430 ( .A1(n19612), .A2(n27517), .Z(n27518) );
  XOR2_X1 U29431 ( .A1(n27661), .A2(n29978), .Z(n27521) );
  XOR2_X1 U29432 ( .A1(n7549), .A2(n29432), .Z(n27522) );
  XOR2_X1 U29433 ( .A1(n38228), .A2(n29689), .Z(n27529) );
  XOR2_X1 U29435 ( .A1(n4934), .A2(n19929), .Z(n27533) );
  XOR2_X1 U29436 ( .A1(n27738), .A2(n19804), .Z(n27536) );
  XOR2_X1 U29438 ( .A1(n27661), .A2(n29371), .Z(n27548) );
  XOR2_X1 U29440 ( .A1(n16320), .A2(n4934), .Z(n27551) );
  NAND2_X1 U29441 ( .A1(n27553), .A2(n38860), .ZN(n27572) );
  XOR2_X1 U29442 ( .A1(n27786), .A2(n19721), .Z(n27568) );
  XOR2_X1 U29443 ( .A1(n37499), .A2(n19735), .Z(n27577) );
  XOR2_X1 U29444 ( .A1(n27735), .A2(n19498), .Z(n27578) );
  NOR2_X1 U29446 ( .A1(n27589), .A2(n27588), .ZN(n27590) );
  XOR2_X1 U29448 ( .A1(n29223), .A2(n27758), .Z(n27600) );
  XOR2_X1 U29449 ( .A1(n27601), .A2(n27600), .Z(n27602) );
  XOR2_X1 U29450 ( .A1(n27603), .A2(n27602), .Z(n27604) );
  XOR2_X1 U29451 ( .A1(n27609), .A2(n27608), .Z(n27614) );
  XOR2_X1 U29452 ( .A1(n34829), .A2(n29801), .Z(n27611) );
  XOR2_X1 U29453 ( .A1(n27612), .A2(n27611), .Z(n27613) );
  XOR2_X1 U29456 ( .A1(n35177), .A2(n30248), .Z(n27627) );
  XOR2_X1 U29457 ( .A1(n27633), .A2(n27828), .Z(n27634) );
  XOR2_X1 U29458 ( .A1(n17418), .A2(n27637), .Z(n27639) );
  XOR2_X1 U29459 ( .A1(n19355), .A2(n19613), .Z(n27638) );
  XOR2_X1 U29460 ( .A1(n27640), .A2(n29141), .Z(n27641) );
  INV_X1 U29461 ( .I(n28074), .ZN(n27652) );
  XOR2_X1 U29462 ( .A1(n900), .A2(n27823), .Z(n27649) );
  XOR2_X1 U29463 ( .A1(n4934), .A2(n19738), .Z(n27651) );
  XOR2_X1 U29464 ( .A1(n19913), .A2(n27724), .Z(n27658) );
  XOR2_X1 U29466 ( .A1(n27679), .A2(n19612), .Z(n27681) );
  XOR2_X1 U29471 ( .A1(n27703), .A2(n31602), .Z(n27704) );
  XOR2_X1 U29472 ( .A1(n27754), .A2(n27705), .Z(n27706) );
  XOR2_X1 U29473 ( .A1(n27848), .A2(n19937), .Z(n27720) );
  XOR2_X1 U29474 ( .A1(n38207), .A2(n27739), .Z(n27740) );
  INV_X1 U29475 ( .I(n27870), .ZN(n27741) );
  XOR2_X1 U29478 ( .A1(n27761), .A2(n29399), .Z(n27762) );
  XOR2_X1 U29479 ( .A1(n27860), .A2(n29363), .Z(n27764) );
  XOR2_X1 U29480 ( .A1(n27765), .A2(n27764), .Z(n27771) );
  XOR2_X1 U29481 ( .A1(n27767), .A2(n27766), .Z(n27768) );
  XOR2_X1 U29482 ( .A1(n27769), .A2(n27768), .Z(n27770) );
  XOR2_X1 U29484 ( .A1(n27786), .A2(n27787), .Z(n27789) );
  XOR2_X1 U29485 ( .A1(n27796), .A2(n19648), .Z(n27797) );
  XOR2_X1 U29486 ( .A1(n35190), .A2(n30068), .Z(n27803) );
  XOR2_X1 U29487 ( .A1(n31585), .A2(n29282), .Z(n27812) );
  MUX2_X1 U29489 ( .I0(n3989), .I1(n28255), .S(n19601), .Z(n27822) );
  XOR2_X1 U29490 ( .A1(n37338), .A2(n27834), .Z(n27836) );
  XOR2_X1 U29491 ( .A1(n4934), .A2(n19833), .Z(n27839) );
  NOR2_X1 U29495 ( .A1(n28727), .A2(n38230), .ZN(n27879) );
  XOR2_X1 U29496 ( .A1(n28874), .A2(n19902), .Z(n27880) );
  NAND3_X1 U29499 ( .A1(n28103), .A2(n17314), .A3(n32352), .ZN(n27889) );
  NAND2_X2 U29500 ( .A1(n27890), .A2(n27889), .ZN(n28696) );
  INV_X1 U29501 ( .I(n28066), .ZN(n27892) );
  NAND3_X1 U29505 ( .A1(n28224), .A2(n39112), .A3(n28229), .ZN(n27913) );
  NOR2_X1 U29507 ( .A1(n28715), .A2(n31015), .ZN(n27927) );
  NOR2_X1 U29509 ( .A1(n33460), .A2(n31015), .ZN(n27926) );
  XOR2_X1 U29511 ( .A1(n36913), .A2(n28827), .Z(n27943) );
  XOR2_X1 U29514 ( .A1(n19774), .A2(n29833), .Z(n27942) );
  NAND2_X1 U29522 ( .A1(n28256), .A2(n28260), .ZN(n27982) );
  NAND2_X1 U29523 ( .A1(n1420), .A2(n13379), .ZN(n27984) );
  NAND3_X1 U29524 ( .A1(n38365), .A2(n11375), .A3(n879), .ZN(n27983) );
  NAND2_X1 U29525 ( .A1(n8522), .A2(n5266), .ZN(n27986) );
  NAND3_X1 U29527 ( .A1(n28238), .A2(n28103), .A3(n1453), .ZN(n27992) );
  NAND2_X1 U29530 ( .A1(n32783), .A2(n1450), .ZN(n28007) );
  NAND2_X1 U29531 ( .A1(n34120), .A2(n13714), .ZN(n28006) );
  NAND2_X1 U29532 ( .A1(n28008), .A2(n1447), .ZN(n28009) );
  NAND2_X1 U29533 ( .A1(n28011), .A2(n28012), .ZN(n28014) );
  NAND2_X1 U29537 ( .A1(n20739), .A2(n4803), .ZN(n28021) );
  NAND2_X1 U29538 ( .A1(n28025), .A2(n28024), .ZN(n28026) );
  NAND2_X1 U29539 ( .A1(n28027), .A2(n28026), .ZN(n28030) );
  OAI21_X1 U29540 ( .A1(n28035), .A2(n28034), .B(n36979), .ZN(n28039) );
  NAND2_X1 U29545 ( .A1(n19280), .A2(n1205), .ZN(n28057) );
  NOR3_X1 U29546 ( .A1(n1072), .A2(n34008), .A3(n28054), .ZN(n28056) );
  NAND2_X1 U29548 ( .A1(n28064), .A2(n28155), .ZN(n28065) );
  XOR2_X1 U29555 ( .A1(n29689), .A2(n28982), .Z(n28100) );
  NAND2_X1 U29556 ( .A1(n7325), .A2(n984), .ZN(n28107) );
  NAND3_X1 U29558 ( .A1(n19946), .A2(n28133), .A3(n28131), .ZN(n28134) );
  MUX2_X1 U29564 ( .I0(n28228), .I1(n28229), .S(n28224), .Z(n28226) );
  NAND2_X1 U29568 ( .A1(n28257), .A2(n28256), .ZN(n28259) );
  NAND2_X1 U29570 ( .A1(n37329), .A2(n28157), .ZN(n28270) );
  NAND2_X1 U29573 ( .A1(n28307), .A2(n9599), .ZN(n28308) );
  AOI21_X1 U29574 ( .A1(n28632), .A2(n14209), .B(n28635), .ZN(n28317) );
  INV_X1 U29575 ( .I(n28634), .ZN(n28316) );
  INV_X1 U29576 ( .I(n28633), .ZN(n28315) );
  XOR2_X1 U29577 ( .A1(n28319), .A2(n28318), .Z(n28320) );
  NAND4_X1 U29578 ( .A1(n28326), .A2(n19038), .A3(n28325), .A4(n30389), .ZN(
        n28328) );
  XOR2_X1 U29579 ( .A1(n4816), .A2(n19879), .Z(n28332) );
  NAND2_X1 U29581 ( .A1(n11413), .A2(n1433), .ZN(n28337) );
  NAND2_X1 U29583 ( .A1(n28350), .A2(n28349), .ZN(n28354) );
  NAND2_X1 U29586 ( .A1(n28509), .A2(n33460), .ZN(n28364) );
  XOR2_X1 U29595 ( .A1(n29221), .A2(n19035), .Z(n28411) );
  XOR2_X1 U29596 ( .A1(n29001), .A2(n28411), .Z(n28412) );
  INV_X1 U29598 ( .I(n28418), .ZN(n28421) );
  NAND3_X1 U29599 ( .A1(n28421), .A2(n28420), .A3(n28419), .ZN(n28424) );
  NAND2_X1 U29600 ( .A1(n28422), .A2(n35694), .ZN(n28423) );
  NOR3_X1 U29601 ( .A1(n18871), .A2(n31045), .A3(n1429), .ZN(n28426) );
  MUX2_X1 U29602 ( .I0(n18875), .I1(n28437), .S(n28554), .Z(n28429) );
  NAND2_X1 U29608 ( .A1(n17735), .A2(n32002), .ZN(n28475) );
  MUX2_X1 U29610 ( .I0(n28486), .I1(n28485), .S(n28484), .Z(n28487) );
  NAND2_X1 U29611 ( .A1(n28487), .A2(n19893), .ZN(n28488) );
  NAND2_X1 U29618 ( .A1(n28745), .A2(n34244), .ZN(n28524) );
  AOI21_X1 U29620 ( .A1(n28530), .A2(n12527), .B(n39435), .ZN(n28531) );
  XOR2_X1 U29622 ( .A1(n7288), .A2(n29832), .Z(n28534) );
  XOR2_X1 U29623 ( .A1(n29076), .A2(n28534), .Z(n28542) );
  XOR2_X1 U29624 ( .A1(n29247), .A2(n19860), .Z(n28541) );
  XOR2_X1 U29626 ( .A1(n28783), .A2(n10794), .Z(n28540) );
  XOR2_X1 U29627 ( .A1(n28791), .A2(n19770), .Z(n28549) );
  NAND2_X1 U29631 ( .A1(n1404), .A2(n29486), .ZN(n28583) );
  AOI21_X1 U29632 ( .A1(n29596), .A2(n33482), .B(n28583), .ZN(n28584) );
  NAND3_X1 U29634 ( .A1(n9599), .A2(n35199), .A3(n35888), .ZN(n28592) );
  XOR2_X1 U29637 ( .A1(n28891), .A2(n28783), .Z(n28630) );
  XOR2_X1 U29646 ( .A1(n29303), .A2(n29145), .Z(n28763) );
  XOR2_X1 U29647 ( .A1(n29058), .A2(n19894), .Z(n28762) );
  XOR2_X1 U29649 ( .A1(n38189), .A2(n29647), .Z(n28775) );
  INV_X1 U29650 ( .I(n19592), .ZN(n28776) );
  XOR2_X1 U29651 ( .A1(n18242), .A2(n29122), .Z(n28779) );
  XOR2_X1 U29652 ( .A1(n29121), .A2(n19936), .Z(n28778) );
  XOR2_X1 U29653 ( .A1(n28779), .A2(n28778), .Z(n28782) );
  XOR2_X1 U29654 ( .A1(n28991), .A2(n5130), .Z(n28786) );
  XOR2_X1 U29655 ( .A1(n28786), .A2(n28785), .Z(n28787) );
  XOR2_X1 U29656 ( .A1(n28842), .A2(n28794), .Z(n28795) );
  NAND3_X1 U29657 ( .A1(n28798), .A2(n28799), .A3(n15273), .ZN(n28797) );
  OAI21_X1 U29658 ( .A1(n28800), .A2(n28798), .B(n28797), .ZN(n28802) );
  NOR2_X1 U29659 ( .A1(n28802), .A2(n28801), .ZN(n28803) );
  XOR2_X1 U29660 ( .A1(n28990), .A2(n28803), .Z(n28804) );
  XOR2_X1 U29661 ( .A1(n296), .A2(n30114), .Z(n28806) );
  AOI21_X1 U29662 ( .A1(n28808), .A2(n33577), .B(n976), .ZN(n28811) );
  XOR2_X1 U29663 ( .A1(n28813), .A2(n30888), .Z(n28814) );
  XOR2_X1 U29664 ( .A1(n29824), .A2(n19760), .Z(n28815) );
  XOR2_X1 U29666 ( .A1(n28865), .A2(n27465), .Z(n28820) );
  NAND2_X1 U29668 ( .A1(n30161), .A2(n29185), .ZN(n28825) );
  XOR2_X1 U29669 ( .A1(n36913), .A2(n5130), .Z(n28828) );
  XOR2_X1 U29670 ( .A1(n29142), .A2(n29718), .Z(n28844) );
  XOR2_X1 U29673 ( .A1(n29837), .A2(n19780), .Z(n28849) );
  XOR2_X1 U29674 ( .A1(n28851), .A2(n28852), .Z(n29099) );
  XOR2_X1 U29675 ( .A1(n28855), .A2(n28854), .Z(n28859) );
  XOR2_X1 U29676 ( .A1(n29030), .A2(n28857), .Z(n28858) );
  NAND3_X1 U29677 ( .A1(n28962), .A2(n28862), .A3(n1178), .ZN(n28863) );
  XOR2_X1 U29678 ( .A1(n29063), .A2(n28865), .Z(n28866) );
  INV_X1 U29683 ( .I(n28883), .ZN(n29592) );
  INV_X1 U29684 ( .I(n29483), .ZN(n29645) );
  NOR2_X1 U29685 ( .A1(n29642), .A2(n29643), .ZN(n29578) );
  XOR2_X1 U29688 ( .A1(n19952), .A2(n28891), .Z(n28892) );
  XOR2_X1 U29689 ( .A1(n28893), .A2(n28892), .Z(n28894) );
  XOR2_X1 U29690 ( .A1(n39220), .A2(n19933), .Z(n28898) );
  NAND2_X1 U29693 ( .A1(n28901), .A2(n28900), .ZN(n28903) );
  NAND2_X1 U29694 ( .A1(n29548), .A2(n35176), .ZN(n29556) );
  NAND2_X1 U29695 ( .A1(n28904), .A2(n29556), .ZN(n28905) );
  XOR2_X1 U29696 ( .A1(n29058), .A2(n19732), .Z(n28912) );
  XOR2_X1 U29697 ( .A1(n34848), .A2(n31127), .Z(n28915) );
  XOR2_X1 U29698 ( .A1(n28916), .A2(n28915), .Z(n28919) );
  XOR2_X1 U29699 ( .A1(n16336), .A2(n28917), .Z(n28918) );
  XOR2_X1 U29700 ( .A1(n31396), .A2(n9930), .Z(n28930) );
  XOR2_X1 U29702 ( .A1(n29306), .A2(n35140), .Z(n28935) );
  XOR2_X1 U29704 ( .A1(n32022), .A2(n19943), .Z(n28944) );
  XOR2_X1 U29707 ( .A1(n29115), .A2(n29146), .Z(n28951) );
  AND2_X1 U29711 ( .A1(n28963), .A2(n28962), .Z(n28964) );
  XOR2_X1 U29712 ( .A1(n29023), .A2(n29123), .Z(n28976) );
  OAI21_X1 U29715 ( .A1(n9649), .A2(n29863), .B(n19878), .ZN(n28980) );
  XOR2_X1 U29718 ( .A1(n9106), .A2(n10794), .Z(n28993) );
  XOR2_X1 U29719 ( .A1(n28991), .A2(n16320), .Z(n28992) );
  XOR2_X1 U29720 ( .A1(n28993), .A2(n28992), .Z(n28994) );
  NAND2_X1 U29721 ( .A1(n29940), .A2(n34179), .ZN(n28996) );
  XOR2_X1 U29722 ( .A1(n28997), .A2(n37112), .Z(n28998) );
  NAND2_X1 U29726 ( .A1(n30134), .A2(n37117), .ZN(n29014) );
  NAND2_X1 U29727 ( .A1(n29014), .A2(n30136), .ZN(n29016) );
  XOR2_X1 U29728 ( .A1(n29019), .A2(n31249), .Z(Ciphertext[61]) );
  XOR2_X1 U29729 ( .A1(n29837), .A2(n29034), .Z(n29035) );
  XOR2_X1 U29730 ( .A1(n29824), .A2(n29320), .Z(n29046) );
  XOR2_X1 U29731 ( .A1(n29801), .A2(n6661), .Z(n29055) );
  XOR2_X1 U29732 ( .A1(n19513), .A2(n29063), .Z(n29064) );
  XOR2_X1 U29734 ( .A1(n17039), .A2(n29805), .Z(n29075) );
  XOR2_X1 U29735 ( .A1(n29076), .A2(n29075), .Z(n29077) );
  XOR2_X1 U29736 ( .A1(n29970), .A2(n29082), .Z(n29083) );
  XOR2_X1 U29738 ( .A1(n29088), .A2(n30253), .Z(n29089) );
  XOR2_X1 U29739 ( .A1(n29090), .A2(n29089), .Z(n29091) );
  XOR2_X1 U29740 ( .A1(n19622), .A2(n29096), .Z(n29097) );
  XOR2_X1 U29743 ( .A1(n19937), .A2(n16357), .Z(n29107) );
  XOR2_X1 U29744 ( .A1(n15581), .A2(n29109), .Z(n29110) );
  XOR2_X1 U29746 ( .A1(n29133), .A2(n29132), .Z(n29134) );
  XOR2_X1 U29747 ( .A1(n31522), .A2(n18242), .Z(n29156) );
  XOR2_X1 U29748 ( .A1(n29155), .A2(n29156), .Z(n29157) );
  NOR2_X1 U29751 ( .A1(n30093), .A2(n35175), .ZN(n29176) );
  NAND2_X1 U29756 ( .A1(n29843), .A2(n773), .ZN(n29190) );
  MUX2_X1 U29757 ( .I0(n29190), .I1(n29871), .S(n29869), .Z(n29193) );
  NAND2_X1 U29758 ( .A1(n29692), .A2(n28), .ZN(n29191) );
  NAND3_X1 U29759 ( .A1(n29871), .A2(n37936), .A3(n29191), .ZN(n29192) );
  NOR2_X1 U29762 ( .A1(n29241), .A2(n29346), .ZN(n29212) );
  INV_X1 U29764 ( .I(n30238), .ZN(n29214) );
  XOR2_X1 U29766 ( .A1(n29217), .A2(n30803), .Z(Ciphertext[8]) );
  NOR2_X1 U29768 ( .A1(n29231), .A2(n29236), .ZN(n29232) );
  XOR2_X1 U29770 ( .A1(n1410), .A2(n29357), .Z(n29244) );
  XOR2_X1 U29773 ( .A1(n38221), .A2(n29290), .Z(n29293) );
  XOR2_X1 U29774 ( .A1(n29829), .A2(n1697), .Z(n29291) );
  NOR2_X1 U29776 ( .A1(n771), .A2(n37100), .ZN(n29314) );
  NOR3_X1 U29777 ( .A1(n14400), .A2(n29446), .A3(n29445), .ZN(n29313) );
  XOR2_X1 U29780 ( .A1(n29338), .A2(n1718), .Z(n29323) );
  NAND3_X1 U29781 ( .A1(n29323), .A2(n29335), .A3(n1391), .ZN(n29332) );
  NAND3_X1 U29782 ( .A1(n29324), .A2(n29338), .A3(n32790), .ZN(n29331) );
  XOR2_X1 U29783 ( .A1(n29325), .A2(n29339), .Z(n29326) );
  NAND3_X1 U29784 ( .A1(n29326), .A2(n20481), .A3(n38156), .ZN(n29330) );
  XOR2_X1 U29785 ( .A1(n16889), .A2(n1718), .Z(n29327) );
  NAND2_X1 U29786 ( .A1(n29328), .A2(n29327), .ZN(n29329) );
  NAND4_X1 U29787 ( .A1(n29332), .A2(n29331), .A3(n29330), .A4(n29329), .ZN(
        Ciphertext[26]) );
  INV_X1 U29788 ( .I(Key[81]), .ZN(n29337) );
  NAND2_X1 U29790 ( .A1(n29361), .A2(n31307), .ZN(n29356) );
  NOR2_X1 U29793 ( .A1(n29373), .A2(n37096), .ZN(n29359) );
  INV_X1 U29794 ( .I(n19933), .ZN(n29360) );
  NAND3_X1 U29798 ( .A1(n29410), .A2(n29413), .A3(n9790), .ZN(n29393) );
  NAND3_X1 U29803 ( .A1(n29390), .A2(n29413), .A3(n17849), .ZN(n29391) );
  NAND2_X1 U29805 ( .A1(n29413), .A2(n29409), .ZN(n29396) );
  INV_X1 U29807 ( .I(n17849), .ZN(n29407) );
  INV_X1 U29808 ( .I(n29413), .ZN(n29408) );
  AOI21_X1 U29809 ( .A1(n35272), .A2(n17849), .B(n29412), .ZN(n29415) );
  XOR2_X1 U29810 ( .A1(n29417), .A2(n19732), .Z(Ciphertext[41]) );
  OAI21_X1 U29812 ( .A1(n1392), .A2(n29438), .B(n29434), .ZN(n29431) );
  NOR3_X1 U29813 ( .A1(n771), .A2(n14400), .A3(n29446), .ZN(n29447) );
  INV_X1 U29814 ( .I(n29461), .ZN(n29469) );
  XOR2_X1 U29815 ( .A1(n29467), .A2(n19839), .Z(Ciphertext[50]) );
  OAI21_X1 U29817 ( .A1(n9636), .A2(n39178), .B(n29490), .ZN(n29505) );
  NAND2_X1 U29818 ( .A1(n29527), .A2(n33427), .ZN(n29504) );
  XOR2_X1 U29821 ( .A1(n29510), .A2(n29509), .Z(Ciphertext[55]) );
  MUX2_X1 U29822 ( .I0(n19362), .I1(n35180), .S(n18384), .Z(n29513) );
  AOI21_X1 U29824 ( .A1(n29513), .A2(n29517), .B(n29512), .ZN(n29515) );
  XOR2_X1 U29825 ( .A1(n29515), .A2(n29514), .Z(Ciphertext[56]) );
  NAND2_X1 U29828 ( .A1(n29519), .A2(n32317), .ZN(n29520) );
  XOR2_X1 U29829 ( .A1(n29523), .A2(n29522), .Z(Ciphertext[57]) );
  OAI21_X1 U29830 ( .A1(n33427), .A2(n35180), .B(n29524), .ZN(n29526) );
  XOR2_X1 U29831 ( .A1(n29529), .A2(n29528), .Z(Ciphertext[58]) );
  AOI21_X1 U29832 ( .A1(n39178), .A2(n29531), .B(n19362), .ZN(n29533) );
  XOR2_X1 U29835 ( .A1(n29539), .A2(n1698), .Z(Ciphertext[60]) );
  MUX2_X1 U29837 ( .I0(n29548), .I1(n35176), .S(n29555), .Z(n29549) );
  NAND2_X1 U29838 ( .A1(n29556), .A2(n29555), .ZN(n29557) );
  NOR2_X1 U29840 ( .A1(n29565), .A2(n29570), .ZN(n29569) );
  XOR2_X1 U29841 ( .A1(n29573), .A2(n35140), .Z(Ciphertext[70]) );
  NOR2_X1 U29842 ( .A1(n20979), .A2(n19147), .ZN(n29580) );
  INV_X1 U29843 ( .I(n29578), .ZN(n29579) );
  NOR2_X1 U29848 ( .A1(n29597), .A2(n29596), .ZN(n29599) );
  AOI21_X1 U29850 ( .A1(n35405), .A2(n29618), .B(n29616), .ZN(n29605) );
  OAI21_X1 U29853 ( .A1(n29616), .A2(n31540), .B(n29617), .ZN(n29607) );
  XOR2_X1 U29854 ( .A1(n29610), .A2(n1733), .Z(Ciphertext[74]) );
  MUX2_X1 U29855 ( .I0(n29616), .I1(n29617), .S(n29619), .Z(n29613) );
  XOR2_X1 U29856 ( .A1(n29615), .A2(n29614), .Z(Ciphertext[75]) );
  NAND2_X1 U29857 ( .A1(n31540), .A2(n29619), .ZN(n29621) );
  NAND2_X1 U29858 ( .A1(n29624), .A2(n29623), .ZN(n29628) );
  INV_X1 U29859 ( .I(n29630), .ZN(n29631) );
  NOR3_X1 U29862 ( .A1(n481), .A2(n29776), .A3(n34914), .ZN(n29640) );
  NAND2_X1 U29867 ( .A1(n19297), .A2(n29641), .ZN(n29652) );
  OAI21_X1 U29868 ( .A1(n29662), .A2(n19297), .B(n17382), .ZN(n29663) );
  NAND2_X1 U29873 ( .A1(n29712), .A2(n29708), .ZN(n29710) );
  NAND3_X1 U29875 ( .A1(n14337), .A2(n29720), .A3(n29721), .ZN(n29715) );
  AOI21_X1 U29877 ( .A1(n29726), .A2(n19348), .B(n29725), .ZN(n29727) );
  XOR2_X1 U29878 ( .A1(n29727), .A2(n1369), .Z(Ciphertext[96]) );
  NOR2_X1 U29880 ( .A1(n29729), .A2(n29752), .ZN(n29731) );
  XOR2_X1 U29881 ( .A1(n29731), .A2(n29730), .Z(Ciphertext[97]) );
  NOR3_X1 U29883 ( .A1(n38143), .A2(n29732), .A3(n29754), .ZN(n29733) );
  XOR2_X1 U29893 ( .A1(n29759), .A2(n19583), .Z(Ciphertext[101]) );
  AOI21_X1 U29896 ( .A1(n1407), .A2(n29815), .B(n29902), .ZN(n29775) );
  NAND2_X1 U29898 ( .A1(n29788), .A2(n19716), .ZN(n29784) );
  NOR2_X1 U29901 ( .A1(n29794), .A2(n29792), .ZN(n29793) );
  NAND2_X1 U29902 ( .A1(n29795), .A2(n29794), .ZN(n29796) );
  NAND3_X1 U29904 ( .A1(n29811), .A2(n6652), .A3(n39018), .ZN(n29807) );
  XOR2_X1 U29905 ( .A1(n29809), .A2(n29808), .Z(Ciphertext[111]) );
  INV_X1 U29906 ( .I(n14403), .ZN(n29900) );
  XOR2_X1 U29907 ( .A1(n11923), .A2(n19885), .Z(n29821) );
  INV_X1 U29908 ( .I(n19890), .ZN(n29825) );
  XOR2_X1 U29909 ( .A1(n39348), .A2(n29825), .Z(n29827) );
  XOR2_X1 U29910 ( .A1(n29828), .A2(n5130), .Z(n29830) );
  INV_X1 U29911 ( .I(n11861), .ZN(n29842) );
  NAND2_X1 U29914 ( .A1(n29883), .A2(n38217), .ZN(n29874) );
  INV_X1 U29915 ( .I(n29883), .ZN(n29888) );
  NOR2_X1 U29919 ( .A1(n30057), .A2(n16353), .ZN(n29896) );
  NAND2_X1 U29920 ( .A1(n1407), .A2(n29900), .ZN(n29901) );
  NOR2_X1 U29922 ( .A1(n29905), .A2(n29954), .ZN(n29910) );
  OAI21_X1 U29923 ( .A1(n29908), .A2(n19878), .B(n29906), .ZN(n29909) );
  AOI21_X1 U29925 ( .A1(n29922), .A2(n1174), .B(n29912), .ZN(n29914) );
  XOR2_X1 U29926 ( .A1(n29915), .A2(n16320), .Z(Ciphertext[128]) );
  INV_X1 U29928 ( .I(n29927), .ZN(n29928) );
  OAI21_X1 U29929 ( .A1(n29929), .A2(n31570), .B(n29928), .ZN(n29933) );
  NAND2_X1 U29930 ( .A1(n21285), .A2(n17240), .ZN(n29947) );
  OAI21_X1 U29931 ( .A1(n29960), .A2(n29955), .B(n29954), .ZN(n29959) );
  OAI21_X1 U29932 ( .A1(n29957), .A2(n18104), .B(n29956), .ZN(n29958) );
  NAND2_X1 U29933 ( .A1(n18104), .A2(n29960), .ZN(n29961) );
  AOI21_X1 U29934 ( .A1(n13705), .A2(n29977), .B(n31512), .ZN(n29962) );
  OAI21_X1 U29936 ( .A1(n29982), .A2(n29973), .B(n29966), .ZN(n29967) );
  XOR2_X1 U29937 ( .A1(n29967), .A2(n19897), .Z(Ciphertext[133]) );
  NAND2_X1 U29939 ( .A1(n9918), .A2(n19909), .ZN(n29985) );
  NAND2_X1 U29940 ( .A1(n29986), .A2(n29985), .ZN(n29988) );
  NOR3_X1 U29943 ( .A1(n15643), .A2(n30038), .A3(n30024), .ZN(n30004) );
  NAND3_X1 U29944 ( .A1(n8529), .A2(n32628), .A3(n36850), .ZN(n30002) );
  XOR2_X1 U29946 ( .A1(n30008), .A2(n30007), .Z(Ciphertext[138]) );
  AOI21_X1 U29947 ( .A1(n30037), .A2(n30024), .B(n30011), .ZN(n30012) );
  AOI21_X1 U29949 ( .A1(n30025), .A2(n39407), .B(n33311), .ZN(n30021) );
  INV_X1 U29950 ( .I(n30017), .ZN(n30019) );
  NOR2_X1 U29951 ( .A1(n30033), .A2(n30022), .ZN(n30018) );
  OAI21_X1 U29952 ( .A1(n30019), .A2(n30018), .B(n30037), .ZN(n30020) );
  NAND2_X1 U29953 ( .A1(n30021), .A2(n30020), .ZN(n30030) );
  OAI21_X1 U29954 ( .A1(n30035), .A2(n30033), .B(n33311), .ZN(n30023) );
  AOI21_X1 U29955 ( .A1(n30025), .A2(n30024), .B(n30023), .ZN(n30028) );
  NAND2_X1 U29956 ( .A1(n30026), .A2(n15643), .ZN(n30027) );
  OAI21_X1 U29957 ( .A1(n30035), .A2(n30034), .B(n30033), .ZN(n30036) );
  XOR2_X1 U29959 ( .A1(n30040), .A2(n16332), .Z(Ciphertext[143]) );
  XOR2_X1 U29964 ( .A1(n30091), .A2(n30090), .Z(Ciphertext[153]) );
  NOR2_X1 U29967 ( .A1(n10118), .A2(n30117), .ZN(n30102) );
  XOR2_X1 U29968 ( .A1(n30105), .A2(n1163), .Z(Ciphertext[157]) );
  MUX2_X1 U29969 ( .I0(n10118), .I1(n35187), .S(n30117), .Z(n30113) );
  NAND2_X1 U29970 ( .A1(n30109), .A2(n35186), .ZN(n30110) );
  XOR2_X1 U29971 ( .A1(n30116), .A2(n30115), .Z(Ciphertext[159]) );
  INV_X1 U29974 ( .I(n19721), .ZN(n30130) );
  XOR2_X1 U29976 ( .A1(n30140), .A2(n17463), .Z(Ciphertext[170]) );
  NAND2_X1 U29977 ( .A1(n34177), .A2(n30141), .ZN(n30143) );
  NAND3_X1 U29980 ( .A1(n30183), .A2(n16676), .A3(n17997), .ZN(n30168) );
  INV_X1 U29981 ( .I(n30162), .ZN(n30163) );
  NAND2_X1 U29982 ( .A1(n30193), .A2(n35210), .ZN(n30194) );
  NOR2_X1 U29984 ( .A1(n31549), .A2(n30210), .ZN(n30204) );
  OAI21_X1 U29986 ( .A1(n30215), .A2(n30214), .B(n30213), .ZN(n30216) );
  NOR2_X1 U29987 ( .A1(n1399), .A2(n30220), .ZN(n30223) );
  NAND3_X1 U29988 ( .A1(n10590), .A2(n17238), .A3(n29210), .ZN(n30231) );
  MUX2_X1 U29990 ( .I0(n30260), .I1(n30259), .S(n30257), .Z(n30255) );
  XOR2_X1 U29991 ( .A1(n30256), .A2(n965), .Z(Ciphertext[190]) );
  OAI21_X1 U29993 ( .A1(n30260), .A2(n30259), .B(n30258), .ZN(n30261) );
  OAI21_X2 U6354 ( .A1(n1042), .A2(n1320), .B(n5111), .ZN(n23056) );
  INV_X2 U1533 ( .I(n7304), .ZN(n21900) );
  AOI21_X2 U8697 ( .A1(n9809), .A2(n19397), .B(n21588), .ZN(n18559) );
  AOI21_X2 U10139 ( .A1(n37216), .A2(n20238), .B(n1840), .ZN(n1839) );
  INV_X4 U357 ( .I(n18689), .ZN(n1206) );
  INV_X2 U1348 ( .I(n17169), .ZN(n13995) );
  INV_X2 U478 ( .I(n7757), .ZN(n27378) );
  NAND2_X2 U6816 ( .A1(n25819), .A2(n32924), .ZN(n12252) );
  INV_X4 U1322 ( .I(n19586), .ZN(n1314) );
  OAI21_X2 U10040 ( .A1(n8720), .A2(n23095), .B(n39356), .ZN(n8719) );
  INV_X4 U1540 ( .I(n3562), .ZN(n21599) );
  INV_X2 U5940 ( .I(n728), .ZN(n9161) );
  NAND2_X2 U2360 ( .A1(n29426), .A2(n29454), .ZN(n29453) );
  AOI21_X2 U2417 ( .A1(n38580), .A2(n28744), .B(n10081), .ZN(n13671) );
  INV_X2 U578 ( .I(n17217), .ZN(n18534) );
  NAND2_X2 U219 ( .A1(n28010), .A2(n28009), .ZN(n28569) );
  INV_X2 U625 ( .I(n26278), .ZN(n26456) );
  INV_X2 U481 ( .I(n27267), .ZN(n27266) );
  OAI21_X2 U801 ( .A1(n25753), .A2(n579), .B(n38300), .ZN(n2316) );
  INV_X2 U6553 ( .I(n8919), .ZN(n29421) );
  INV_X2 U6099 ( .I(n12055), .ZN(n8919) );
  AOI21_X2 U22329 ( .A1(n20308), .A2(n12077), .B(n10242), .ZN(n20961) );
  INV_X2 U6566 ( .I(n30186), .ZN(n30159) );
  INV_X2 U5570 ( .I(n29341), .ZN(n1391) );
  NAND2_X2 U1446 ( .A1(n15382), .A2(n15380), .ZN(n22132) );
  INV_X2 U6323 ( .I(n10635), .ZN(n1613) );
  INV_X2 U1346 ( .I(n13694), .ZN(n23142) );
  INV_X2 U753 ( .I(n18987), .ZN(n25770) );
  INV_X2 U1454 ( .I(n9970), .ZN(n1151) );
  NAND2_X2 U10923 ( .A1(n3965), .A2(n6435), .ZN(n3964) );
  AOI21_X2 U13851 ( .A1(n21694), .A2(n15910), .B(n15812), .ZN(n15811) );
  BUF_X2 U8778 ( .I(Key[30]), .Z(n29509) );
  AOI21_X2 U1300 ( .A1(n1043), .A2(n19000), .B(n14556), .ZN(n23155) );
  NAND2_X2 U50 ( .A1(n29272), .A2(n29273), .ZN(n29277) );
  AOI22_X2 U8104 ( .A1(n25427), .A2(n19296), .B1(n15180), .B2(n14515), .ZN(
        n4595) );
  NAND2_X2 U785 ( .A1(n17471), .A2(n4046), .ZN(n26019) );
  INV_X2 U586 ( .I(n19225), .ZN(n7752) );
  NAND2_X2 U414 ( .A1(n21248), .A2(n31287), .ZN(n27507) );
  NOR2_X2 U1074 ( .A1(n24184), .A2(n24300), .ZN(n13881) );
  NAND2_X2 U6076 ( .A1(n33404), .A2(n18720), .ZN(n16074) );
  INV_X2 U1244 ( .I(n4618), .ZN(n23569) );
  INV_X2 U897 ( .I(n7967), .ZN(n25116) );
  NAND2_X1 U3017 ( .A1(n22829), .A2(n23042), .ZN(n20911) );
  BUF_X2 U10480 ( .I(Key[9]), .Z(n19498) );
  INV_X2 U1124 ( .I(n14709), .ZN(n24266) );
  INV_X4 U18608 ( .I(n20793), .ZN(n29869) );
  NOR2_X2 U5813 ( .A1(n3293), .A2(n21895), .ZN(n13421) );
  AOI21_X2 U7500 ( .A1(n9017), .A2(n34915), .B(n33841), .ZN(n9016) );
  NAND2_X2 U13839 ( .A1(n14920), .A2(n14919), .ZN(n21370) );
  NAND2_X2 U25076 ( .A1(n7613), .A2(n133), .ZN(n22187) );
  INV_X2 U2474 ( .I(n19844), .ZN(n28311) );
  AOI22_X2 U26764 ( .A1(n31359), .A2(n25468), .B1(n25609), .B2(n17332), .ZN(
        n17331) );
  AOI21_X2 U1402 ( .A1(n11277), .A2(n15229), .B(n11276), .ZN(n11275) );
  NAND2_X2 U8055 ( .A1(n5098), .A2(n4516), .ZN(n19241) );
  NOR2_X2 U2487 ( .A1(n28772), .A2(n17771), .ZN(n28293) );
  NAND2_X2 U9923 ( .A1(n4207), .A2(n31931), .ZN(n10709) );
  NAND2_X2 U9639 ( .A1(n24770), .A2(n8173), .ZN(n24772) );
  INV_X2 U100 ( .I(n37060), .ZN(n6851) );
  AOI21_X2 U7065 ( .A1(n20998), .A2(n10709), .B(n23444), .ZN(n9347) );
  NOR2_X2 U2467 ( .A1(n11658), .A2(n30443), .ZN(n13642) );
  INV_X2 U8623 ( .I(n22178), .ZN(n1148) );
  INV_X1 U10677 ( .I(n29437), .ZN(n1389) );
  INV_X2 U6137 ( .I(n16327), .ZN(n28191) );
  INV_X2 U1441 ( .I(n22155), .ZN(n15004) );
  NOR2_X2 U163 ( .A1(n20737), .A2(n20736), .ZN(n20735) );
  INV_X2 U1093 ( .I(n802), .ZN(n24221) );
  INV_X4 U1104 ( .I(n17911), .ZN(n1125) );
  NAND2_X2 U8455 ( .A1(n14305), .A2(n19614), .ZN(n8721) );
  NOR2_X2 U11632 ( .A1(n27270), .A2(n33050), .ZN(n16479) );
  AOI21_X2 U15569 ( .A1(n13337), .A2(n3119), .B(n13336), .ZN(n13335) );
  INV_X2 U5680 ( .I(n833), .ZN(n18734) );
  INV_X2 U1442 ( .I(n8493), .ZN(n15493) );
  NAND2_X2 U5518 ( .A1(n1300), .A2(n6218), .ZN(n23553) );
  INV_X1 U3123 ( .I(n26876), .ZN(n4218) );
  INV_X2 U346 ( .I(n27910), .ZN(n15704) );
  INV_X2 U9998 ( .I(n22923), .ZN(n15770) );
  INV_X2 U7213 ( .I(n9422), .ZN(n18999) );
  INV_X2 U7110 ( .I(n23390), .ZN(n1644) );
  AOI21_X2 U13228 ( .A1(n37196), .A2(n23355), .B(n32158), .ZN(n19006) );
  AOI21_X2 U821 ( .A1(n25472), .A2(n31359), .B(n25409), .ZN(n15404) );
  INV_X4 U5938 ( .I(n18164), .ZN(n25359) );
  INV_X2 U356 ( .I(n5525), .ZN(n28286) );
  AOI22_X2 U8930 ( .A1(n17115), .A2(n3532), .B1(n1419), .B2(n28683), .ZN(
        n18191) );
  NAND2_X2 U6933 ( .A1(n19678), .A2(n25261), .ZN(n15459) );
  AOI22_X2 U14233 ( .A1(n4697), .A2(n9141), .B1(n1881), .B2(n33591), .ZN(n4076) );
  NAND2_X1 U1769 ( .A1(n25396), .A2(n25397), .ZN(n12995) );
  AND2_X1 U5449 ( .A1(n27985), .A2(n34008), .Z(n6050) );
  NOR2_X2 U1391 ( .A1(n22126), .A2(n12077), .ZN(n22255) );
  AOI21_X2 U7111 ( .A1(n23027), .A2(n23026), .B(n23025), .ZN(n23542) );
  AOI22_X2 U18300 ( .A1(n37146), .A2(n17225), .B1(n20508), .B2(n5384), .ZN(
        n15710) );
  AOI21_X2 U2260 ( .A1(n6045), .A2(n19693), .B(n36225), .ZN(n6044) );
  NAND2_X2 U10043 ( .A1(n22928), .A2(n14817), .ZN(n23066) );
  NAND2_X2 U1461 ( .A1(n3618), .A2(n1990), .ZN(n2190) );
  NAND2_X2 U8251 ( .A1(n24696), .A2(n39196), .ZN(n24695) );
  CLKBUF_X4 U2025 ( .I(n4179), .Z(n26) );
  INV_X2 U324 ( .I(n27903), .ZN(n28181) );
  OAI21_X2 U13768 ( .A1(n20773), .A2(n21664), .B(n1344), .ZN(n4917) );
  OAI21_X2 U16088 ( .A1(n1300), .A2(n6218), .B(n31685), .ZN(n4606) );
  INV_X2 U8169 ( .I(n25380), .ZN(n10674) );
  NAND2_X2 U12321 ( .A1(n25702), .A2(n19296), .ZN(n11889) );
  NAND2_X2 U1383 ( .A1(n1658), .A2(n10037), .ZN(n3025) );
  OAI21_X2 U279 ( .A1(n14585), .A2(n4306), .B(n33612), .ZN(n20201) );
  OAI21_X2 U12783 ( .A1(n14154), .A2(n36757), .B(n6298), .ZN(n24277) );
  OAI22_X2 U25154 ( .A1(n23262), .A2(n23263), .B1(n20867), .B2(n961), .ZN(
        n16758) );
  INV_X4 U841 ( .I(n10414), .ZN(n14410) );
  INV_X2 U1833 ( .I(n33263), .ZN(n25939) );
  INV_X2 U5849 ( .I(n29307), .ZN(n29389) );
  AOI22_X2 U5862 ( .A1(n27887), .A2(n39789), .B1(n18687), .B2(n28175), .ZN(
        n28595) );
  INV_X2 U1094 ( .I(n7319), .ZN(n17871) );
  INV_X2 U6005 ( .I(n22599), .ZN(n1656) );
  INV_X2 U5959 ( .I(n24696), .ZN(n24806) );
  INV_X4 U6930 ( .I(n19863), .ZN(n1117) );
  INV_X2 U134 ( .I(n39443), .ZN(n29459) );
  NAND2_X2 U6745 ( .A1(n18904), .A2(n18902), .ZN(n26822) );
  NAND2_X2 U9835 ( .A1(n7399), .A2(n11167), .ZN(n23655) );
  OAI21_X2 U9043 ( .A1(n28282), .A2(n16544), .B(n10827), .ZN(n28069) );
  NAND2_X2 U16181 ( .A1(n13421), .A2(n3670), .ZN(n14920) );
  NOR2_X2 U12098 ( .A1(n25977), .A2(n7258), .ZN(n11032) );
  NAND2_X2 U6391 ( .A1(n22356), .A2(n22353), .ZN(n22352) );
  AOI21_X2 U24827 ( .A1(n22880), .A2(n23034), .B(n23035), .ZN(n22882) );
  NAND2_X2 U25819 ( .A1(n21579), .A2(n11274), .ZN(n21707) );
  INV_X2 U5857 ( .I(n28621), .ZN(n974) );
  INV_X2 U1497 ( .I(n21506), .ZN(n21551) );
  NOR2_X2 U7221 ( .A1(n22267), .A2(n19515), .ZN(n22071) );
  INV_X2 U22122 ( .I(n16500), .ZN(n17114) );
  NAND2_X2 U6501 ( .A1(n8147), .A2(n20720), .ZN(n29472) );
  INV_X4 U6283 ( .I(n24874), .ZN(n1580) );
  INV_X2 U6061 ( .I(n29475), .ZN(n29478) );
  NAND2_X2 U21805 ( .A1(n17485), .A2(n39666), .ZN(n17484) );
  OAI22_X2 U24501 ( .A1(n12144), .A2(n36887), .B1(n17938), .B2(n17233), .ZN(
        n17485) );
  CLKBUF_X4 U5588 ( .I(n29495), .Z(n18720) );
  INV_X2 U558 ( .I(n38591), .ZN(n1500) );
  INV_X4 U12741 ( .I(n10667), .ZN(n2731) );
  INV_X4 U15485 ( .I(n3158), .ZN(n28246) );
  NOR2_X2 U1728 ( .A1(n12540), .A2(n12538), .ZN(n20642) );
  NAND2_X2 U5892 ( .A1(n9240), .A2(n9239), .ZN(n27131) );
  NAND2_X2 U1382 ( .A1(n1663), .A2(n3236), .ZN(n3237) );
  INV_X2 U615 ( .I(n302), .ZN(n5960) );
  NAND2_X2 U265 ( .A1(n28030), .A2(n28029), .ZN(n28390) );
  INV_X2 U25429 ( .I(n21937), .ZN(n21939) );
  OAI21_X2 U18209 ( .A1(n23405), .A2(n5258), .B(n9190), .ZN(n23407) );
  OAI21_X2 U1281 ( .A1(n16892), .A2(n32878), .B(n21143), .ZN(n22814) );
  NOR2_X2 U2785 ( .A1(n4827), .A2(n4620), .ZN(n6830) );
  NAND2_X2 U8408 ( .A1(n23539), .A2(n23337), .ZN(n23116) );
  OAI21_X2 U915 ( .A1(n14168), .A2(n24740), .B(n14165), .ZN(n14164) );
  INV_X4 U7261 ( .I(n14493), .ZN(n21702) );
  INV_X2 U13356 ( .I(n23592), .ZN(n19232) );
  BUF_X4 U1245 ( .I(n23613), .Z(n4525) );
  BUF_X2 U10885 ( .I(n29865), .Z(n29937) );
  BUF_X4 U5566 ( .I(n20307), .Z(n18588) );
  OAI21_X2 U6624 ( .A1(n14103), .A2(n11876), .B(n11875), .ZN(n14760) );
  NAND2_X2 U6333 ( .A1(n12154), .A2(n6159), .ZN(n12153) );
  OAI21_X2 U25235 ( .A1(n14952), .A2(n25855), .B(n34961), .ZN(n16117) );
  BUF_X2 U14043 ( .I(Key[5]), .Z(n29602) );
  NAND2_X2 U2309 ( .A1(n10003), .A2(n32258), .ZN(n8727) );
  OAI21_X2 U7194 ( .A1(n18566), .A2(n21449), .B(n3676), .ZN(n9225) );
  INV_X2 U1536 ( .I(n20596), .ZN(n18926) );
  OAI21_X2 U5900 ( .A1(n30348), .A2(n2929), .B(n36392), .ZN(n7282) );
  INV_X2 U6098 ( .I(n30154), .ZN(n30155) );
  OAI21_X2 U28816 ( .A1(n1288), .A2(n1593), .B(n32360), .ZN(n24240) );
  INV_X2 U616 ( .I(n20389), .ZN(n26992) );
  OAI21_X2 U12259 ( .A1(n14589), .A2(n15924), .B(n17029), .ZN(n16896) );
  INV_X4 U6538 ( .I(n892), .ZN(n9394) );
  NAND2_X2 U7156 ( .A1(n14560), .A2(n783), .ZN(n20518) );
  AOI21_X2 U283 ( .A1(n2664), .A2(n1206), .B(n2663), .ZN(n3192) );
  BUF_X2 U6371 ( .I(n8943), .Z(n5581) );
  NAND2_X2 U940 ( .A1(n24964), .A2(n3214), .ZN(n25022) );
  INV_X2 U126 ( .I(n20524), .ZN(n30242) );
  INV_X2 U1123 ( .I(n12758), .ZN(n5985) );
  BUF_X2 U8546 ( .I(n22943), .Z(n23167) );
  NAND2_X2 U6023 ( .A1(n11329), .A2(n8519), .ZN(n22288) );
  INV_X2 U8559 ( .I(n22676), .ZN(n1667) );
  INV_X2 U7476 ( .I(n17225), .ZN(n13762) );
  AOI22_X2 U13428 ( .A1(n23185), .A2(n19538), .B1(n14396), .B2(n11328), .ZN(
        n14017) );
  INV_X2 U96 ( .I(n20649), .ZN(n29940) );
  AOI21_X2 U7847 ( .A1(n12173), .A2(n31502), .B(n12172), .ZN(n12171) );
  INV_X1 U3209 ( .I(n27854), .ZN(n1461) );
  NOR2_X2 U7287 ( .A1(n18205), .A2(n21787), .ZN(n21499) );
  NAND2_X2 U8639 ( .A1(n22086), .A2(n36006), .ZN(n22022) );
  INV_X2 U393 ( .I(n20976), .ZN(n1077) );
  AOI22_X2 U24537 ( .A1(n37152), .A2(n17112), .B1(n21508), .B2(n33852), .ZN(
        n21513) );
  INV_X4 U28865 ( .I(n25048), .ZN(n24909) );
  INV_X2 U1350 ( .I(n12471), .ZN(n13650) );
  NAND2_X2 U756 ( .A1(n1098), .A2(n25899), .ZN(n10168) );
  NAND2_X2 U8016 ( .A1(n26016), .A2(n25899), .ZN(n26118) );
  INV_X4 U7241 ( .I(n11568), .ZN(n19873) );
  NOR2_X2 U11326 ( .A1(n4809), .A2(n14562), .ZN(n2663) );
  OAI22_X2 U13449 ( .A1(n22554), .A2(n19288), .B1(n22555), .B2(n22995), .ZN(
        n6970) );
  INV_X2 U475 ( .I(n9037), .ZN(n13471) );
  OAI21_X2 U6008 ( .A1(n4765), .A2(n22136), .B(n31412), .ZN(n16347) );
  AOI21_X2 U12289 ( .A1(n25471), .A2(n25472), .B(n2962), .ZN(n25473) );
  OAI21_X2 U5946 ( .A1(n1118), .A2(n16547), .B(n2747), .ZN(n2745) );
  OAI21_X1 U4157 ( .A1(n29918), .A2(n31570), .B(n29916), .ZN(n434) );
  NOR2_X2 U5941 ( .A1(n39289), .A2(n16246), .ZN(n10753) );
  BUF_X2 U10464 ( .I(Key[142]), .Z(n29838) );
  AOI21_X2 U2266 ( .A1(n27031), .A2(n27318), .B(n16101), .ZN(n27032) );
  INV_X1 U4597 ( .I(n529), .ZN(n528) );
  NAND2_X2 U24771 ( .A1(n37152), .A2(n32544), .ZN(n21596) );
  INV_X1 U8523 ( .I(n8628), .ZN(n19319) );
  INV_X2 U5943 ( .I(n15883), .ZN(n16246) );
  AOI21_X2 U9416 ( .A1(n19241), .A2(n4602), .B(n32979), .ZN(n4400) );
  INV_X2 U1352 ( .I(n30443), .ZN(n23045) );
  NAND2_X2 U7055 ( .A1(n23373), .A2(n23374), .ZN(n23376) );
  INV_X4 U7113 ( .I(n16528), .ZN(n1302) );
  INV_X2 U635 ( .I(n26252), .ZN(n26504) );
  AOI21_X2 U9634 ( .A1(n6770), .A2(n1565), .B(n11957), .ZN(n23826) );
  INV_X4 U112 ( .I(n29455), .ZN(n29426) );
  INV_X2 U1134 ( .I(n14290), .ZN(n16832) );
  INV_X2 U638 ( .I(n19847), .ZN(n1503) );
  INV_X4 U16530 ( .I(n4056), .ZN(n5077) );
  INV_X1 U12236 ( .I(n11148), .ZN(n1519) );
  NAND2_X2 U10119 ( .A1(n8744), .A2(n8745), .ZN(n9334) );
  INV_X4 U5673 ( .I(n9959), .ZN(n910) );
  INV_X2 U382 ( .I(n27674), .ZN(n18924) );
  NAND3_X2 U20219 ( .A1(n1203), .A2(n28419), .A3(n33902), .ZN(n28154) );
  BUF_X2 U6057 ( .I(Key[73]), .Z(n19937) );
  NOR2_X2 U27638 ( .A1(n20930), .A2(n20929), .ZN(n20928) );
  NOR2_X2 U27690 ( .A1(n3293), .A2(n19699), .ZN(n21489) );
  NOR2_X2 U8511 ( .A1(n4846), .A2(n23101), .ZN(n15638) );
  NAND2_X2 U1456 ( .A1(n6419), .A2(n6417), .ZN(n20351) );
  INV_X2 U6440 ( .I(n20703), .ZN(n21550) );
  INV_X2 U2045 ( .I(n33417), .ZN(n18374) );
  INV_X2 U1537 ( .I(n21575), .ZN(n21594) );
  OAI21_X1 U26110 ( .A1(n31412), .A2(n35771), .B(n16364), .ZN(n16621) );
  INV_X2 U1523 ( .I(n2533), .ZN(n17102) );
  OAI22_X2 U10142 ( .A1(n21985), .A2(n21986), .B1(n37216), .B2(n20238), .ZN(
        n14754) );
  NOR2_X2 U1043 ( .A1(n1606), .A2(n626), .ZN(n4475) );
  INV_X2 U7891 ( .I(n26994), .ZN(n19433) );
  INV_X4 U7088 ( .I(n37774), .ZN(n12597) );
  INV_X2 U6123 ( .I(n28595), .ZN(n28698) );
  NAND3_X2 U2734 ( .A1(n22021), .A2(n22020), .A3(n14181), .ZN(n22024) );
  AOI22_X2 U1464 ( .A1(n1349), .A2(n2280), .B1(n2279), .B2(n21820), .ZN(n237)
         );
  INV_X1 U7102 ( .I(n32616), .ZN(n1291) );
  INV_X1 U3833 ( .I(n35373), .ZN(n14939) );
  OAI22_X2 U29291 ( .A1(n26831), .A2(n38928), .B1(n38852), .B2(n7752), .ZN(
        n26682) );
  AOI21_X2 U2271 ( .A1(n12398), .A2(n39037), .B(n8036), .ZN(n5287) );
  AOI22_X2 U8644 ( .A1(n21719), .A2(n32704), .B1(n21720), .B2(n19647), .ZN(
        n13241) );
  AOI22_X2 U11769 ( .A1(n8815), .A2(n26951), .B1(n8816), .B2(n1236), .ZN(
        n16700) );
  NOR2_X2 U8378 ( .A1(n23508), .A2(n13150), .ZN(n13149) );
  BUF_X4 U8451 ( .I(n14856), .Z(n10174) );
  NAND2_X2 U10747 ( .A1(n7749), .A2(n32415), .ZN(n10731) );
  OAI21_X2 U5933 ( .A1(n20216), .A2(n25514), .B(n13129), .ZN(n19209) );
  NAND3_X1 U12551 ( .A1(n8648), .A2(n33412), .A3(n8647), .ZN(n11906) );
  INV_X2 U1127 ( .I(n39814), .ZN(n19895) );
  INV_X2 U1498 ( .I(n13473), .ZN(n6241) );
  INV_X2 U9758 ( .I(n37934), .ZN(n24411) );
  BUF_X2 U13974 ( .I(n21602), .Z(n21784) );
  INV_X2 U2342 ( .I(n7993), .ZN(n94) );
  NAND2_X2 U6757 ( .A1(n33952), .A2(n31157), .ZN(n26975) );
  NAND2_X2 U8712 ( .A1(n20544), .A2(n17938), .ZN(n21309) );
  AOI22_X2 U24454 ( .A1(n16448), .A2(n14705), .B1(n16447), .B2(n12771), .ZN(
        n16446) );
  INV_X2 U9500 ( .I(n31010), .ZN(n7853) );
  INV_X4 U19660 ( .I(n23467), .ZN(n6969) );
  NAND2_X2 U24804 ( .A1(n10174), .A2(n23582), .ZN(n23581) );
  NAND2_X2 U1436 ( .A1(n14027), .A2(n2839), .ZN(n14037) );
  OAI21_X2 U1413 ( .A1(n14251), .A2(n19471), .B(n22080), .ZN(n16623) );
  NAND2_X2 U8578 ( .A1(n36731), .A2(n4613), .ZN(n22059) );
  BUF_X4 U5984 ( .I(n23296), .Z(n23458) );
  INV_X2 U6446 ( .I(n21882), .ZN(n21507) );
  BUF_X4 U394 ( .I(n3963), .Z(n10653) );
  INV_X2 U8708 ( .I(n21640), .ZN(n11411) );
  NAND2_X2 U13358 ( .A1(n8144), .A2(n8143), .ZN(n22927) );
  INV_X1 U13597 ( .I(n1323), .ZN(n6473) );
  INV_X2 U10435 ( .I(n14418), .ZN(n20544) );
  OAI21_X2 U8030 ( .A1(n6543), .A2(n25835), .B(n31954), .ZN(n9461) );
  NAND2_X2 U8059 ( .A1(n1522), .A2(n25900), .ZN(n26119) );
  OAI22_X2 U24300 ( .A1(n17333), .A2(n17334), .B1(n17335), .B2(n14196), .ZN(
        n17942) );
  OR2_X2 U13963 ( .A1(n21387), .A2(n21743), .Z(n21749) );
  INV_X2 U10143 ( .I(n16487), .ZN(n5246) );
  NAND3_X2 U15522 ( .A1(n6345), .A2(n3077), .A3(n6346), .ZN(n23561) );
  INV_X1 U8034 ( .I(n603), .ZN(n21041) );
  NAND2_X2 U2980 ( .A1(n126), .A2(n16495), .ZN(n29249) );
  NOR2_X1 U11246 ( .A1(n27621), .A2(n28149), .ZN(n17753) );
  INV_X2 U6542 ( .I(n14179), .ZN(n29348) );
  INV_X2 U7222 ( .I(n21961), .ZN(n22190) );
  INV_X1 U307 ( .I(n11890), .ZN(n27962) );
  INV_X2 U5996 ( .I(n23132), .ZN(n23209) );
  NAND2_X1 U2117 ( .A1(n13268), .A2(n7403), .ZN(n13267) );
  AOI22_X2 U10726 ( .A1(n34070), .A2(n29059), .B1(n30187), .B2(n7989), .ZN(
        n8202) );
  OAI22_X2 U24133 ( .A1(n15788), .A2(n25512), .B1(n36991), .B2(n13744), .ZN(
        n15789) );
  INV_X1 U1741 ( .I(n21674), .ZN(n21862) );
  NAND2_X2 U24338 ( .A1(n14305), .A2(n16463), .ZN(n18227) );
  NAND2_X1 U2110 ( .A1(n22079), .A2(n16625), .ZN(n16624) );
  INV_X4 U2168 ( .I(n20309), .ZN(n1146) );
  AOI21_X2 U12260 ( .A1(n21136), .A2(n9161), .B(n21135), .ZN(n11251) );
  NAND2_X2 U7012 ( .A1(n1127), .A2(n24232), .ZN(n24332) );
  NAND2_X1 U17878 ( .A1(n12323), .A2(n11055), .ZN(n9313) );
  INV_X2 U1121 ( .I(n15873), .ZN(n16366) );
  INV_X2 U7597 ( .I(n28390), .ZN(n28486) );
  INV_X2 U22098 ( .I(n15165), .ZN(n13076) );
  INV_X2 U9561 ( .I(n30317), .ZN(n25512) );
  INV_X4 U11872 ( .I(n19712), .ZN(n2140) );
  INV_X1 U243 ( .I(n32535), .ZN(n1189) );
  INV_X4 U7282 ( .I(n670), .ZN(n21920) );
  AOI21_X2 U12261 ( .A1(n25383), .A2(n1117), .B(n25382), .ZN(n25384) );
  AOI21_X2 U9853 ( .A1(n23579), .A2(n23581), .B(n13831), .ZN(n20946) );
  OAI21_X2 U2666 ( .A1(n14634), .A2(n15276), .B(n40), .ZN(n15772) );
  OAI21_X2 U10000 ( .A1(n15638), .A2(n1824), .B(n13734), .ZN(n6469) );
  OAI21_X2 U6952 ( .A1(n24824), .A2(n24494), .B(n4351), .ZN(n24496) );
  INV_X1 U3177 ( .I(n2799), .ZN(n10104) );
  INV_X2 U16523 ( .I(n4048), .ZN(n10158) );
  OAI22_X2 U24440 ( .A1(n22839), .A2(n23103), .B1(n22838), .B2(n19788), .ZN(
        n22842) );
  AOI21_X1 U12095 ( .A1(n6783), .A2(n2349), .B(n2621), .ZN(n6785) );
  INV_X4 U13015 ( .I(n7834), .ZN(n5953) );
  AOI21_X2 U3171 ( .A1(n12387), .A2(n10019), .B(n10193), .ZN(n12364) );
  INV_X2 U5820 ( .I(n21668), .ZN(n21845) );
  BUF_X4 U8445 ( .I(n23478), .Z(n8692) );
  INV_X4 U6667 ( .I(n14389), .ZN(n1074) );
  INV_X2 U619 ( .I(n10523), .ZN(n26269) );
  INV_X4 U10102 ( .I(n6327), .ZN(n23060) );
  NAND2_X1 U949 ( .A1(n12385), .A2(n18110), .ZN(n4608) );
  NAND2_X1 U12055 ( .A1(n7677), .A2(n7678), .ZN(n4431) );
  AOI21_X2 U12846 ( .A1(n8360), .A2(n1279), .B(n8359), .ZN(n8358) );
  NAND2_X2 U10168 ( .A1(n22070), .A2(n34452), .ZN(n22381) );
  INV_X2 U9594 ( .I(n14164), .ZN(n25014) );
  INV_X4 U7836 ( .I(n614), .ZN(n15360) );
  OAI21_X2 U957 ( .A1(n24518), .A2(n39817), .B(n18114), .ZN(n12914) );
  INV_X2 U6565 ( .I(n21116), .ZN(n9918) );
  NAND3_X2 U22955 ( .A1(n11378), .A2(n13805), .A3(n39672), .ZN(n18594) );
  AOI22_X2 U9981 ( .A1(n22893), .A2(n20590), .B1(n22793), .B2(n9975), .ZN(
        n11671) );
  INV_X2 U5869 ( .I(n27523), .ZN(n27674) );
  INV_X1 U24388 ( .I(n10029), .ZN(n26672) );
  NAND2_X2 U12466 ( .A1(n4603), .A2(n5050), .ZN(n19965) );
  NAND2_X2 U29860 ( .A1(n31517), .A2(n29636), .ZN(n29638) );
  NAND2_X2 U916 ( .A1(n14826), .A2(n24845), .ZN(n25155) );
  INV_X2 U28 ( .I(n17996), .ZN(n30177) );
  INV_X4 U6121 ( .I(n17751), .ZN(n11164) );
  INV_X2 U335 ( .I(n34008), .ZN(n984) );
  OAI21_X2 U9740 ( .A1(n9386), .A2(n9519), .B(n1606), .ZN(n9381) );
  AOI22_X2 U9690 ( .A1(n24399), .A2(n1587), .B1(n35384), .B2(n24107), .ZN(
        n24108) );
  AOI22_X2 U11186 ( .A1(n12787), .A2(n38307), .B1(n12785), .B2(n12784), .ZN(
        n6926) );
  INV_X1 U6664 ( .I(n9775), .ZN(n18948) );
  NAND2_X2 U13477 ( .A1(n20564), .A2(n23088), .ZN(n17083) );
  NAND2_X1 U11196 ( .A1(n13847), .A2(n7586), .ZN(n10394) );
  OR2_X1 U14227 ( .A1(n14967), .A2(n1874), .Z(n2899) );
  INV_X4 U23616 ( .I(n17509), .ZN(n24359) );
  AOI21_X2 U2218 ( .A1(n18459), .A2(n31796), .B(n4845), .ZN(n18458) );
  INV_X1 U839 ( .I(n36019), .ZN(n7265) );
  NAND2_X2 U10135 ( .A1(n14036), .A2(n9843), .ZN(n22044) );
  INV_X2 U13806 ( .I(n22250), .ZN(n8496) );
  INV_X2 U898 ( .I(n25114), .ZN(n25267) );
  INV_X2 U7549 ( .I(n7429), .ZN(n28740) );
  INV_X2 U18790 ( .I(n5974), .ZN(n17464) );
  INV_X1 U9241 ( .I(n27165), .ZN(n1223) );
  NAND2_X2 U12293 ( .A1(n25335), .A2(n31809), .ZN(n20464) );
  INV_X4 U1455 ( .I(n7843), .ZN(n11329) );
  NAND2_X1 U20471 ( .A1(n13892), .A2(n38159), .ZN(n8734) );
  OAI21_X2 U7022 ( .A1(n13185), .A2(n12771), .B(n14705), .ZN(n12090) );
  NOR2_X2 U6274 ( .A1(n37105), .A2(n12672), .ZN(n12671) );
  AOI21_X2 U12265 ( .A1(n25476), .A2(n25512), .B(n16026), .ZN(n16024) );
  INV_X1 U24178 ( .I(n19085), .ZN(n29278) );
  INV_X1 U11399 ( .I(n31571), .ZN(n21160) );
  INV_X4 U23907 ( .I(n13316), .ZN(n16585) );
  INV_X2 U14157 ( .I(n20284), .ZN(n29870) );
  INV_X4 U1108 ( .I(n24244), .ZN(n959) );
  OAI21_X1 U24953 ( .A1(n1235), .A2(n26743), .B(n26741), .ZN(n26745) );
  INV_X2 U12154 ( .I(n25876), .ZN(n7079) );
  NAND2_X1 U24400 ( .A1(n24096), .A2(n24478), .ZN(n16430) );
  INV_X4 U20896 ( .I(n20359), .ZN(n17029) );
  NAND2_X1 U10678 ( .A1(n6803), .A2(n971), .ZN(n29895) );
  AOI21_X2 U13207 ( .A1(n23522), .A2(n34959), .B(n23521), .ZN(n17122) );
  NAND2_X2 U10049 ( .A1(n32515), .A2(n14409), .ZN(n18822) );
  OAI22_X2 U29409 ( .A1(n27421), .A2(n27420), .B1(n30544), .B2(n31518), .ZN(
        n27426) );
  AOI22_X2 U21478 ( .A1(n16236), .A2(n7426), .B1(n23318), .B2(n23317), .ZN(
        n16235) );
  INV_X2 U2608 ( .I(n19807), .ZN(n25) );
  INV_X8 U7001 ( .I(n16585), .ZN(n1029) );
  NAND2_X2 U17237 ( .A1(n31004), .A2(n8304), .ZN(n25400) );
  OR2_X1 U26387 ( .A1(n24265), .A2(n24086), .Z(n16311) );
  INV_X1 U7114 ( .I(n14856), .ZN(n23506) );
  INV_X2 U7127 ( .I(n23587), .ZN(n23325) );
  NOR2_X2 U10974 ( .A1(n28598), .A2(n39425), .ZN(n13718) );
  INV_X2 U2267 ( .I(n6285), .ZN(n1211) );
  AOI22_X2 U1467 ( .A1(n21760), .A2(n21759), .B1(n21758), .B2(n21757), .ZN(
        n22177) );
  NOR2_X2 U12661 ( .A1(n5431), .A2(n13495), .ZN(n24568) );
  INV_X2 U6316 ( .I(n11449), .ZN(n24403) );
  BUF_X2 U6000 ( .I(n23196), .Z(n12029) );
  OAI21_X2 U12080 ( .A1(n4248), .A2(n13885), .B(n30937), .ZN(n4247) );
  OAI21_X2 U13124 ( .A1(n20066), .A2(n21118), .B(n19665), .ZN(n7399) );
  INV_X1 U5555 ( .I(n7696), .ZN(n20535) );
  NAND2_X2 U8029 ( .A1(n930), .A2(n7258), .ZN(n9228) );
  INV_X1 U4472 ( .I(n29548), .ZN(n1394) );
  NAND2_X2 U8344 ( .A1(n17546), .A2(n19566), .ZN(n24129) );
  OAI22_X2 U12279 ( .A1(n8032), .A2(n12558), .B1(n8034), .B2(n12557), .ZN(
        n3343) );
  INV_X1 U29889 ( .I(n29750), .ZN(n29751) );
  AOI21_X2 U8672 ( .A1(n17126), .A2(n34021), .B(n21731), .ZN(n12511) );
  INV_X2 U6227 ( .I(n25961), .ZN(n8711) );
  INV_X2 U5614 ( .I(n19417), .ZN(n985) );
  OAI21_X1 U28730 ( .A1(n24819), .A2(n33412), .B(n23824), .ZN(n23825) );
  BUF_X2 U8783 ( .I(Key[180]), .Z(n30065) );
  NAND2_X2 U6030 ( .A1(n4242), .A2(n4241), .ZN(n22389) );
  INV_X2 U5692 ( .I(n25216), .ZN(n13531) );
  AOI21_X2 U8092 ( .A1(n37071), .A2(n39327), .B(n14316), .ZN(n16767) );
  NAND2_X2 U1796 ( .A1(n13202), .A2(n21053), .ZN(n13201) );
  INV_X2 U1519 ( .I(n21742), .ZN(n21713) );
  BUF_X2 U11402 ( .I(n27875), .Z(n28200) );
  NAND3_X1 U16672 ( .A1(n28456), .A2(n28099), .A3(n6405), .ZN(n4196) );
  INV_X1 U17947 ( .I(n9668), .ZN(n15580) );
  NAND2_X2 U6265 ( .A1(n1267), .A2(n19422), .ZN(n18573) );
  INV_X1 U13155 ( .I(n24051), .ZN(n1621) );
  INV_X1 U5751 ( .I(n39070), .ZN(n1308) );
  INV_X2 U11758 ( .I(n21101), .ZN(n1486) );
  OAI21_X2 U914 ( .A1(n24580), .A2(n9997), .B(n24885), .ZN(n24984) );
  OAI21_X2 U1194 ( .A1(n3363), .A2(n3366), .B(n17122), .ZN(n16488) );
  OAI21_X2 U13459 ( .A1(n14628), .A2(n16604), .B(n22996), .ZN(n8144) );
  NAND2_X2 U12568 ( .A1(n24568), .A2(n6822), .ZN(n21053) );
  NAND2_X2 U8404 ( .A1(n23488), .A2(n23487), .ZN(n23599) );
  BUF_X2 U10451 ( .I(Key[8]), .Z(n29718) );
  NAND2_X2 U12868 ( .A1(n11265), .A2(n10694), .ZN(n10693) );
  INV_X2 U18480 ( .I(n8395), .ZN(n28267) );
  BUF_X2 U10458 ( .I(Key[137]), .Z(n29394) );
  BUF_X2 U6454 ( .I(Key[108]), .Z(n29320) );
  BUF_X2 U14036 ( .I(Key[146]), .Z(n19648) );
  BUF_X2 U7319 ( .I(Key[151]), .Z(n29970) );
  BUF_X2 U10450 ( .I(Key[163]), .Z(n29325) );
  BUF_X2 U7311 ( .I(Key[96]), .Z(n19897) );
  BUF_X2 U6463 ( .I(Key[124]), .Z(n29983) );
  BUF_X2 U14047 ( .I(Key[110]), .Z(n19947) );
  BUF_X2 U5828 ( .I(Key[103]), .Z(n19908) );
  BUF_X2 U10476 ( .I(Key[154]), .Z(n19903) );
  BUF_X2 U8782 ( .I(Key[16]), .Z(n19407) );
  BUF_X2 U7321 ( .I(Key[160]), .Z(n19751) );
  BUF_X2 U8785 ( .I(Key[138]), .Z(n19890) );
  BUF_X2 U6472 ( .I(Key[70]), .Z(n19613) );
  BUF_X2 U6055 ( .I(Key[1]), .Z(n19758) );
  BUF_X2 U8786 ( .I(Key[42]), .Z(n30010) );
  BUF_X2 U20017 ( .I(Key[98]), .Z(n19866) );
  BUF_X2 U10456 ( .I(Key[165]), .Z(n29411) );
  BUF_X2 U6469 ( .I(Key[19]), .Z(n19860) );
  BUF_X2 U6457 ( .I(Key[82]), .Z(n19894) );
  BUF_X2 U6462 ( .I(Key[7]), .Z(n19952) );
  BUF_X2 U7322 ( .I(Key[162]), .Z(n19845) );
  BUF_X2 U8780 ( .I(Key[79]), .Z(n19681) );
  BUF_X2 U6470 ( .I(Key[190]), .Z(n19592) );
  BUF_X2 U14029 ( .I(Key[169]), .Z(n19820) );
  BUF_X2 U14027 ( .I(Key[13]), .Z(n19876) );
  BUF_X2 U14031 ( .I(Key[14]), .Z(n29974) );
  BUF_X2 U14040 ( .I(Key[127]), .Z(n19833) );
  BUF_X2 U10442 ( .I(Key[141]), .Z(n29554) );
  BUF_X2 U8791 ( .I(Key[120]), .Z(n19808) );
  BUF_X2 U8777 ( .I(Key[121]), .Z(n19774) );
  BUF_X2 U8788 ( .I(Key[50]), .Z(n29295) );
  BUF_X2 U6058 ( .I(Key[85]), .Z(n29514) );
  BUF_X2 U14033 ( .I(Key[170]), .Z(n19910) );
  BUF_X2 U10462 ( .I(Key[39]), .Z(n19874) );
  BUF_X2 U14026 ( .I(Key[84]), .Z(n19760) );
  BUF_X2 U14063 ( .I(Key[189]), .Z(n18270) );
  BUF_X2 U7316 ( .I(Key[46]), .Z(n19721) );
  BUF_X2 U8771 ( .I(Key[60]), .Z(n29003) );
  BUF_X2 U10468 ( .I(Key[76]), .Z(n19877) );
  BUF_X2 U14068 ( .I(Key[25]), .Z(n29269) );
  BUF_X2 U8770 ( .I(Key[88]), .Z(n19919) );
  BUF_X2 U8757 ( .I(Key[69]), .Z(n29978) );
  BUF_X2 U6455 ( .I(Key[130]), .Z(n19932) );
  BUF_X2 U10441 ( .I(Key[181]), .Z(n30085) );
  BUF_X2 U6471 ( .I(Key[40]), .Z(n19527) );
  INV_X1 U13991 ( .I(n29229), .ZN(n17705) );
  BUF_X2 U6046 ( .I(n21880), .Z(n17112) );
  INV_X1 U8736 ( .I(n19730), .ZN(n1362) );
  CLKBUF_X2 U4582 ( .I(n688), .Z(n526) );
  INV_X2 U3061 ( .I(n32370), .ZN(n19202) );
  INV_X1 U28713 ( .I(n19749), .ZN(n29934) );
  INV_X1 U14055 ( .I(n21791), .ZN(n1722) );
  BUF_X2 U6445 ( .I(n21368), .Z(n21892) );
  INV_X1 U1507 ( .I(n32820), .ZN(n918) );
  CLKBUF_X2 U4668 ( .I(n17964), .Z(n547) );
  INV_X2 U7278 ( .I(n21684), .ZN(n21681) );
  NAND2_X1 U24533 ( .A1(n21932), .A2(n21931), .ZN(n21936) );
  NAND2_X1 U10353 ( .A1(n6504), .A2(n21476), .ZN(n21522) );
  NOR3_X1 U28210 ( .A1(n21748), .A2(n21712), .A3(n21652), .ZN(n21388) );
  INV_X1 U13903 ( .I(n21718), .ZN(n5531) );
  OAI21_X1 U1472 ( .A1(n3943), .A2(n10961), .B(n261), .ZN(n3913) );
  CLKBUF_X4 U8637 ( .I(n22350), .Z(n19837) );
  INV_X1 U13670 ( .I(n17308), .ZN(n21996) );
  INV_X2 U16609 ( .I(n8882), .ZN(n9252) );
  AOI21_X1 U8596 ( .A1(n16266), .A2(n22356), .B(n30315), .ZN(n3971) );
  BUF_X2 U8541 ( .I(n22862), .Z(n9472) );
  INV_X1 U20559 ( .I(n2046), .ZN(n17131) );
  CLKBUF_X1 U10085 ( .I(n23131), .Z(n19859) );
  CLKBUF_X1 U13560 ( .I(n19692), .Z(n9975) );
  BUF_X2 U13529 ( .I(n18220), .Z(n16963) );
  CLKBUF_X2 U2720 ( .I(n3952), .Z(n59) );
  CLKBUF_X2 U5239 ( .I(n11643), .Z(n3310) );
  OR2_X1 U2089 ( .A1(n23100), .A2(n21094), .Z(n13137) );
  INV_X1 U13436 ( .I(n23146), .ZN(n5945) );
  NAND2_X1 U28604 ( .A1(n23134), .A2(n23133), .ZN(n23137) );
  NAND2_X1 U23379 ( .A1(n23191), .A2(n12163), .ZN(n18501) );
  NAND2_X1 U13350 ( .A1(n5749), .A2(n17917), .ZN(n5748) );
  NAND2_X1 U13363 ( .A1(n5039), .A2(n5038), .ZN(n6423) );
  INV_X2 U5746 ( .I(n30881), .ZN(n1038) );
  NOR2_X1 U22846 ( .A1(n23588), .A2(n1306), .ZN(n11168) );
  CLKBUF_X2 U3871 ( .I(n23685), .Z(n360) );
  INV_X2 U1097 ( .I(n37259), .ZN(n13653) );
  BUF_X2 U13034 ( .I(n19341), .Z(n9844) );
  CLKBUF_X2 U13036 ( .I(n24196), .Z(n19402) );
  INV_X1 U8332 ( .I(n38702), .ZN(n24357) );
  INV_X2 U12975 ( .I(n13453), .ZN(n8463) );
  CLKBUF_X2 U3744 ( .I(n17844), .Z(n326) );
  NOR2_X1 U28824 ( .A1(n24275), .A2(n17709), .ZN(n24278) );
  INV_X2 U5711 ( .I(n24764), .ZN(n1269) );
  NOR2_X1 U20984 ( .A1(n35813), .A2(n8430), .ZN(n9257) );
  NOR2_X1 U16273 ( .A1(n36955), .A2(n24638), .ZN(n3751) );
  INV_X2 U12525 ( .I(n24961), .ZN(n1555) );
  BUF_X2 U8199 ( .I(n11497), .Z(n4664) );
  BUF_X2 U12473 ( .I(n25392), .Z(n25689) );
  OAI21_X1 U2696 ( .A1(n21233), .A2(n9241), .B(n12675), .ZN(n25628) );
  NAND2_X1 U28874 ( .A1(n24553), .A2(n25394), .ZN(n24554) );
  NAND2_X1 U22764 ( .A1(n34583), .A2(n11018), .ZN(n14669) );
  INV_X1 U9437 ( .I(n37378), .ZN(n8883) );
  NOR2_X1 U17452 ( .A1(n9380), .A2(n9379), .ZN(n4776) );
  INV_X2 U591 ( .I(n861), .ZN(n1492) );
  INV_X1 U2119 ( .I(n13854), .ZN(n13952) );
  INV_X1 U11697 ( .I(n37245), .ZN(n27098) );
  INV_X1 U11491 ( .I(n6818), .ZN(n13270) );
  INV_X1 U1711 ( .I(n27407), .ZN(n1483) );
  OR2_X1 U21027 ( .A1(n26889), .A2(n36183), .Z(n8485) );
  NAND2_X1 U23096 ( .A1(n11638), .A2(n11637), .ZN(n11639) );
  INV_X1 U1651 ( .I(n37639), .ZN(n1459) );
  INV_X1 U11456 ( .I(n27537), .ZN(n8865) );
  CLKBUF_X2 U2863 ( .I(n11459), .Z(n99) );
  INV_X1 U11392 ( .I(n28101), .ZN(n11732) );
  OAI22_X1 U29493 ( .A1(n27996), .A2(n11461), .B1(n27876), .B2(n27998), .ZN(
        n27877) );
  INV_X1 U11280 ( .I(n28197), .ZN(n8880) );
  OAI21_X1 U23674 ( .A1(n12807), .A2(n30846), .B(n27980), .ZN(n12808) );
  INV_X1 U25498 ( .I(n28324), .ZN(n19038) );
  INV_X1 U10977 ( .I(n10305), .ZN(n28697) );
  INV_X1 U4165 ( .I(n28382), .ZN(n28457) );
  OAI21_X1 U4685 ( .A1(n552), .A2(n551), .B(n36775), .ZN(n28477) );
  NAND2_X1 U10999 ( .A1(n11163), .A2(n28337), .ZN(n28338) );
  INV_X1 U15169 ( .I(n3126), .ZN(n3127) );
  INV_X1 U26306 ( .I(n14525), .ZN(n29353) );
  INV_X1 U25319 ( .I(n35210), .ZN(n19193) );
  NAND2_X1 U10782 ( .A1(n29842), .A2(n21290), .ZN(n21289) );
  CLKBUF_X4 U6084 ( .I(n8919), .Z(n8918) );
  NOR2_X1 U10735 ( .A1(n21324), .A2(n3379), .ZN(n17877) );
  NAND2_X1 U10716 ( .A1(n7899), .A2(n18043), .ZN(n8228) );
  CLKBUF_X2 U10439 ( .I(Key[66]), .Z(n19763) );
  BUF_X2 U7314 ( .I(Key[147]), .Z(n19950) );
  BUF_X2 U10491 ( .I(Key[36]), .Z(n19817) );
  BUF_X2 U14054 ( .I(Key[176]), .Z(n29857) );
  BUF_X2 U6460 ( .I(Key[61]), .Z(n29051) );
  INV_X1 U25528 ( .I(n30253), .ZN(n20483) );
  INV_X1 U27951 ( .I(n21628), .ZN(n21435) );
  BUF_X2 U1506 ( .I(n18576), .Z(n1990) );
  INV_X1 U8533 ( .I(n23196), .ZN(n19645) );
  NOR2_X1 U9985 ( .A1(n22922), .A2(n5838), .ZN(n5749) );
  OAI21_X1 U13175 ( .A1(n20841), .A2(n35506), .B(n4968), .ZN(n11530) );
  INV_X1 U13121 ( .I(n23764), .ZN(n2044) );
  BUF_X2 U13047 ( .I(n16792), .Z(n9963) );
  INV_X2 U24173 ( .I(n13872), .ZN(n25261) );
  BUF_X2 U3643 ( .I(n33947), .Z(n299) );
  INV_X2 U12430 ( .I(n25695), .ZN(n13129) );
  OAI22_X1 U28873 ( .A1(n19398), .A2(n25681), .B1(n33946), .B2(n25647), .ZN(
        n24553) );
  NAND2_X1 U29062 ( .A1(n25515), .A2(n19767), .ZN(n25516) );
  NAND2_X1 U29049 ( .A1(n5886), .A2(n31311), .ZN(n25459) );
  NOR2_X1 U27213 ( .A1(n39112), .A2(n19891), .ZN(n20164) );
  CLKBUF_X2 U8916 ( .I(n9393), .Z(n5414) );
  BUF_X2 U5585 ( .I(n11348), .Z(n10590) );
  AOI22_X2 U9229 ( .A1(n26710), .A2(n26179), .B1(n11305), .B2(n1493), .ZN(
        n10595) );
  NOR2_X2 U10997 ( .A1(n12541), .A2(n11438), .ZN(n12540) );
  NAND2_X2 U1730 ( .A1(n34171), .A2(n11490), .ZN(n12541) );
  AOI21_X2 U7990 ( .A1(n9228), .A2(n25925), .B(n9227), .ZN(n9226) );
  INV_X2 U27135 ( .I(n18157), .ZN(n21111) );
  INV_X4 U8498 ( .I(n9677), .ZN(n13734) );
  OAI21_X2 U8663 ( .A1(n38438), .A2(n1355), .B(n5601), .ZN(n7964) );
  INV_X1 U6421 ( .I(n19387), .ZN(n21887) );
  NOR2_X1 U21688 ( .A1(n9552), .A2(n10629), .ZN(n21710) );
  NAND2_X1 U28360 ( .A1(n1692), .A2(n19337), .ZN(n21877) );
  NOR2_X1 U3733 ( .A1(n31604), .A2(n21667), .ZN(n20468) );
  AOI21_X1 U24722 ( .A1(n18417), .A2(n19542), .B(n1157), .ZN(n21533) );
  NAND2_X1 U10359 ( .A1(n1692), .A2(n19395), .ZN(n21874) );
  INV_X2 U1500 ( .I(n21436), .ZN(n919) );
  NOR2_X1 U10356 ( .A1(n21833), .A2(n19620), .ZN(n8436) );
  AOI22_X1 U13943 ( .A1(n19434), .A2(n21484), .B1(n21881), .B2(n17112), .ZN(
        n13856) );
  AOI21_X1 U28247 ( .A1(n21678), .A2(n21417), .B(n36351), .ZN(n21420) );
  NAND2_X1 U22030 ( .A1(n17792), .A2(n9809), .ZN(n19511) );
  AOI21_X1 U26135 ( .A1(n15338), .A2(n13855), .B(n21579), .ZN(n21580) );
  NOR2_X1 U26692 ( .A1(n21868), .A2(n15359), .ZN(n17992) );
  NOR2_X1 U22925 ( .A1(n21902), .A2(n35921), .ZN(n21623) );
  AOI21_X1 U24513 ( .A1(n15761), .A2(n21579), .B(n36754), .ZN(n15522) );
  NOR3_X1 U26737 ( .A1(n9642), .A2(n20332), .A3(n21308), .ZN(n20331) );
  NOR2_X1 U1491 ( .A1(n31604), .A2(n21668), .ZN(n21670) );
  AOI21_X1 U10336 ( .A1(n1158), .A2(n21666), .B(n8936), .ZN(n9318) );
  AOI21_X1 U2947 ( .A1(n3293), .A2(n21892), .B(n21894), .ZN(n119) );
  NAND2_X1 U1468 ( .A1(n10961), .A2(n587), .ZN(n6295) );
  NAND2_X1 U2562 ( .A1(n21834), .A2(n21837), .ZN(n9317) );
  NOR3_X1 U24511 ( .A1(n18417), .A2(n21712), .A3(n1157), .ZN(n19274) );
  NOR2_X1 U26230 ( .A1(n16302), .A2(n21751), .ZN(n15926) );
  NAND3_X1 U28275 ( .A1(n36728), .A2(n21784), .A3(n32664), .ZN(n21504) );
  NOR2_X1 U10281 ( .A1(n19037), .A2(n9425), .ZN(n21460) );
  AOI22_X1 U24540 ( .A1(n21621), .A2(n21917), .B1(n33141), .B2(n18412), .ZN(
        n18900) );
  INV_X1 U8613 ( .I(n22150), .ZN(n22151) );
  INV_X2 U14928 ( .I(n8431), .ZN(n18567) );
  INV_X2 U16434 ( .I(n39489), .ZN(n22327) );
  NAND2_X1 U5789 ( .A1(n38687), .A2(n22038), .ZN(n3835) );
  NAND2_X1 U4927 ( .A1(n18567), .A2(n8040), .ZN(n3682) );
  NOR2_X1 U18583 ( .A1(n33581), .A2(n915), .ZN(n5734) );
  NOR2_X1 U27848 ( .A1(n1335), .A2(n22310), .ZN(n20282) );
  INV_X1 U24538 ( .I(n32675), .ZN(n17411) );
  NOR2_X1 U10152 ( .A1(n22065), .A2(n12077), .ZN(n20299) );
  INV_X1 U4174 ( .I(n19773), .ZN(n22268) );
  AOI21_X1 U16723 ( .A1(n12230), .A2(n4240), .B(n19873), .ZN(n7815) );
  NAND2_X1 U13668 ( .A1(n34282), .A2(n13519), .ZN(n22309) );
  AOI21_X1 U20323 ( .A1(n37089), .A2(n22143), .B(n8029), .ZN(n8028) );
  INV_X1 U27346 ( .I(n22342), .ZN(n18766) );
  NAND3_X1 U28146 ( .A1(n22307), .A2(n33359), .A3(n1335), .ZN(n21335) );
  AOI21_X1 U13653 ( .A1(n16499), .A2(n22256), .B(n18567), .ZN(n15967) );
  INV_X2 U13601 ( .I(n10488), .ZN(n22668) );
  INV_X1 U13725 ( .I(n13704), .ZN(n3239) );
  INV_X1 U28349 ( .I(n22572), .ZN(n22559) );
  INV_X1 U13585 ( .I(n22508), .ZN(n7162) );
  INV_X1 U1699 ( .I(n34073), .ZN(n23005) );
  INV_X1 U1364 ( .I(n4997), .ZN(n19000) );
  NOR2_X1 U13546 ( .A1(n12925), .A2(n36369), .ZN(n22467) );
  NAND2_X1 U10064 ( .A1(n12315), .A2(n19645), .ZN(n23199) );
  OAI21_X1 U8487 ( .A1(n16963), .A2(n22915), .B(n3310), .ZN(n6712) );
  NOR2_X1 U10021 ( .A1(n20372), .A2(n5515), .ZN(n5785) );
  NAND2_X1 U25742 ( .A1(n22467), .A2(n22899), .ZN(n15201) );
  INV_X1 U1299 ( .I(n23190), .ZN(n10828) );
  NAND2_X1 U10024 ( .A1(n7960), .A2(n19293), .ZN(n22917) );
  NOR2_X1 U4706 ( .A1(n22709), .A2(n18415), .ZN(n22861) );
  INV_X2 U8524 ( .I(n33934), .ZN(n19538) );
  NAND3_X1 U5987 ( .A1(n14396), .A2(n17968), .A3(n23186), .ZN(n20302) );
  NAND3_X1 U13439 ( .A1(n22979), .A2(n22978), .A3(n38524), .ZN(n10471) );
  NOR2_X1 U13420 ( .A1(n23030), .A2(n5380), .ZN(n12509) );
  NAND2_X1 U18105 ( .A1(n23161), .A2(n5111), .ZN(n16887) );
  INV_X2 U1259 ( .I(n23607), .ZN(n1637) );
  OAI21_X1 U8394 ( .A1(n1302), .A2(n5492), .B(n5487), .ZN(n5491) );
  AOI21_X1 U7062 ( .A1(n10432), .A2(n13834), .B(n1138), .ZN(n9758) );
  NAND2_X1 U27907 ( .A1(n23576), .A2(n23577), .ZN(n20472) );
  NAND2_X1 U28676 ( .A1(n23567), .A2(n23566), .ZN(n23544) );
  NAND2_X1 U20053 ( .A1(n23324), .A2(n19481), .ZN(n7389) );
  NAND2_X1 U23342 ( .A1(n37523), .A2(n31906), .ZN(n12094) );
  NAND2_X1 U13200 ( .A1(n23638), .A2(n23637), .ZN(n3276) );
  INV_X1 U8416 ( .I(n31331), .ZN(n1629) );
  AOI22_X1 U13293 ( .A1(n14901), .A2(n34012), .B1(n23346), .B2(n35191), .ZN(
        n2814) );
  NAND3_X1 U28588 ( .A1(n23364), .A2(n9078), .A3(n23361), .ZN(n23018) );
  AOI21_X1 U28681 ( .A1(n23611), .A2(n23610), .B(n38611), .ZN(n23616) );
  NOR2_X1 U3543 ( .A1(n18866), .A2(n34959), .ZN(n3365) );
  INV_X2 U5976 ( .I(n2117), .ZN(n14491) );
  INV_X1 U6315 ( .I(n24369), .ZN(n24087) );
  INV_X1 U5539 ( .I(n24421), .ZN(n24419) );
  NAND2_X1 U1058 ( .A1(n24432), .A2(n24431), .ZN(n21125) );
  INV_X1 U9812 ( .I(n30320), .ZN(n24392) );
  OAI21_X1 U24855 ( .A1(n17546), .A2(n24465), .B(n24316), .ZN(n18346) );
  AOI21_X1 U5034 ( .A1(n1602), .A2(n16779), .B(n9922), .ZN(n14052) );
  NAND2_X1 U25804 ( .A1(n15320), .A2(n20312), .ZN(n15319) );
  AOI21_X1 U3529 ( .A1(n13453), .A2(n9066), .B(n12248), .ZN(n9068) );
  NAND2_X1 U5965 ( .A1(n24338), .A2(n12953), .ZN(n10421) );
  NOR2_X1 U5729 ( .A1(n18697), .A2(n20027), .ZN(n24147) );
  NAND2_X1 U1029 ( .A1(n24814), .A2(n24623), .ZN(n24734) );
  NOR2_X1 U970 ( .A1(n24529), .A2(n5897), .ZN(n24530) );
  INV_X1 U6278 ( .I(n33230), .ZN(n19431) );
  INV_X1 U5285 ( .I(n24735), .ZN(n24852) );
  NAND2_X1 U6982 ( .A1(n17618), .A2(n7529), .ZN(n24494) );
  NOR2_X1 U28884 ( .A1(n16238), .A2(n35981), .ZN(n24596) );
  NAND2_X1 U12611 ( .A1(n6822), .A2(n5431), .ZN(n9478) );
  NAND2_X1 U22153 ( .A1(n18845), .A2(n36376), .ZN(n18844) );
  NAND2_X1 U9660 ( .A1(n14267), .A2(n19431), .ZN(n14266) );
  NOR2_X1 U26524 ( .A1(n39681), .A2(n7552), .ZN(n24715) );
  NAND2_X1 U19083 ( .A1(n6337), .A2(n19484), .ZN(n6336) );
  NAND2_X1 U12642 ( .A1(n6186), .A2(n1026), .ZN(n6184) );
  INV_X1 U25204 ( .I(n24532), .ZN(n24618) );
  NAND3_X1 U17943 ( .A1(n38674), .A2(n38668), .A3(n5124), .ZN(n5122) );
  NOR2_X1 U9655 ( .A1(n31845), .A2(n1026), .ZN(n13583) );
  NAND2_X1 U9619 ( .A1(n37106), .A2(n5431), .ZN(n9500) );
  OAI22_X1 U23403 ( .A1(n20301), .A2(n19886), .B1(n24566), .B2(n12159), .ZN(
        n12208) );
  INV_X2 U19609 ( .I(n37052), .ZN(n13943) );
  INV_X1 U22529 ( .I(n10584), .ZN(n17774) );
  NOR2_X1 U25559 ( .A1(n18880), .A2(n20359), .ZN(n14778) );
  INV_X1 U9572 ( .I(n25631), .ZN(n25728) );
  NAND2_X1 U29068 ( .A1(n25550), .A2(n25549), .ZN(n25556) );
  NOR2_X1 U6896 ( .A1(n25550), .A2(n1537), .ZN(n11066) );
  NOR2_X1 U8118 ( .A1(n13943), .A2(n16264), .ZN(n14100) );
  NOR2_X1 U12385 ( .A1(n9800), .A2(n14460), .ZN(n9482) );
  NAND2_X1 U16100 ( .A1(n3602), .A2(n34755), .ZN(n25346) );
  INV_X1 U2599 ( .I(n25157), .ZN(n9915) );
  INV_X1 U2179 ( .I(n835), .ZN(n1543) );
  NOR2_X1 U2652 ( .A1(n33785), .A2(n25623), .ZN(n17075) );
  NAND2_X1 U1838 ( .A1(n7238), .A2(n19237), .ZN(n7237) );
  NAND3_X1 U21225 ( .A1(n20855), .A2(n1546), .A3(n19589), .ZN(n14262) );
  INV_X1 U757 ( .I(n25836), .ZN(n18375) );
  INV_X1 U739 ( .I(n21204), .ZN(n1512) );
  INV_X1 U15899 ( .I(n33644), .ZN(n25934) );
  NOR2_X1 U27387 ( .A1(n1528), .A2(n1245), .ZN(n20134) );
  INV_X1 U20192 ( .I(n25849), .ZN(n25888) );
  NAND2_X1 U744 ( .A1(n834), .A2(n1245), .ZN(n4769) );
  NAND2_X1 U9436 ( .A1(n1011), .A2(n6056), .ZN(n3838) );
  OR2_X1 U6206 ( .A1(n17008), .A2(n11533), .Z(n9892) );
  NAND3_X1 U19144 ( .A1(n25850), .A2(n25851), .A3(n928), .ZN(n6398) );
  NAND2_X1 U28988 ( .A1(n25996), .A2(n25994), .ZN(n25112) );
  OAI21_X1 U9421 ( .A1(n6056), .A2(n4382), .B(n4381), .ZN(n2124) );
  NOR2_X1 U26842 ( .A1(n7767), .A2(n33263), .ZN(n20611) );
  AOI21_X1 U4889 ( .A1(n26213), .A2(n9868), .B(n26212), .ZN(n14503) );
  INV_X1 U9345 ( .I(n26968), .ZN(n19338) );
  NAND2_X1 U2010 ( .A1(n36344), .A2(n860), .ZN(n26622) );
  NOR3_X1 U19421 ( .A1(n862), .A2(n26639), .A3(n17515), .ZN(n12177) );
  NOR2_X1 U24957 ( .A1(n26847), .A2(n10314), .ZN(n20316) );
  NOR2_X1 U570 ( .A1(n39823), .A2(n17237), .ZN(n17323) );
  NAND2_X1 U11851 ( .A1(n20699), .A2(n9179), .ZN(n16177) );
  INV_X1 U24962 ( .I(n19371), .ZN(n16222) );
  NOR2_X1 U9328 ( .A1(n26830), .A2(n26959), .ZN(n6909) );
  NAND2_X1 U26161 ( .A1(n19332), .A2(n26740), .ZN(n27014) );
  AOI21_X1 U24922 ( .A1(n11616), .A2(n26751), .B(n26752), .ZN(n17229) );
  NOR2_X1 U7852 ( .A1(n26898), .A2(n39287), .ZN(n27043) );
  NAND2_X1 U24997 ( .A1(n20575), .A2(n20576), .ZN(n20574) );
  NOR2_X1 U9290 ( .A1(n11707), .A2(n36391), .ZN(n12987) );
  OAI21_X1 U524 ( .A1(n11674), .A2(n16522), .B(n19425), .ZN(n10535) );
  INV_X1 U7832 ( .I(n8988), .ZN(n8830) );
  OAI21_X1 U3326 ( .A1(n31254), .A2(n20699), .B(n212), .ZN(n10796) );
  AOI21_X1 U29230 ( .A1(n26724), .A2(n16970), .B(n26627), .ZN(n26372) );
  INV_X2 U19038 ( .I(n9369), .ZN(n20133) );
  NAND2_X1 U22471 ( .A1(n10461), .A2(n12156), .ZN(n17720) );
  INV_X1 U441 ( .I(n18047), .ZN(n1085) );
  INV_X1 U2627 ( .I(n17072), .ZN(n27201) );
  INV_X1 U517 ( .I(n7424), .ZN(n16946) );
  NAND2_X1 U15504 ( .A1(n31518), .A2(n3059), .ZN(n26953) );
  NAND2_X1 U29411 ( .A1(n30412), .A2(n19719), .ZN(n27445) );
  NOR2_X1 U25318 ( .A1(n27092), .A2(n16043), .ZN(n19077) );
  NOR2_X1 U29112 ( .A1(n27069), .A2(n31433), .ZN(n26074) );
  NAND2_X1 U25259 ( .A1(n17720), .A2(n35427), .ZN(n17719) );
  INV_X2 U11731 ( .I(n997), .ZN(n1474) );
  OAI21_X1 U29389 ( .A1(n27436), .A2(n27235), .B(n27234), .ZN(n27236) );
  INV_X1 U11439 ( .I(n27776), .ZN(n27705) );
  INV_X2 U23394 ( .I(n12187), .ZN(n28114) );
  INV_X1 U26252 ( .I(n32932), .ZN(n28248) );
  NOR2_X1 U7695 ( .A1(n28024), .A2(n20739), .ZN(n28022) );
  NOR2_X1 U9052 ( .A1(n7690), .A2(n2877), .ZN(n2876) );
  NAND3_X1 U342 ( .A1(n8523), .A2(n27901), .A3(n27996), .ZN(n28403) );
  NAND3_X1 U20312 ( .A1(n39574), .A2(n99), .A3(n19366), .ZN(n7586) );
  NAND3_X1 U6642 ( .A1(n11283), .A2(n36854), .A3(n3662), .ZN(n2872) );
  AOI21_X1 U1737 ( .A1(n19366), .A2(n28230), .B(n12257), .ZN(n28232) );
  NOR2_X1 U9066 ( .A1(n28079), .A2(n1070), .ZN(n7431) );
  NOR3_X1 U9082 ( .A1(n3159), .A2(n28248), .A3(n28246), .ZN(n3065) );
  NAND2_X1 U24994 ( .A1(n28187), .A2(n16325), .ZN(n16063) );
  NAND2_X1 U11185 ( .A1(n33959), .A2(n6236), .ZN(n3794) );
  NOR2_X1 U29641 ( .A1(n30716), .A2(n180), .ZN(n28664) );
  INV_X2 U19163 ( .I(n6426), .ZN(n28759) );
  INV_X2 U204 ( .I(n28330), .ZN(n1186) );
  INV_X1 U2672 ( .I(n28478), .ZN(n3532) );
  INV_X1 U6631 ( .I(n36478), .ZN(n1427) );
  INV_X1 U11121 ( .I(n28580), .ZN(n13825) );
  NOR2_X1 U24106 ( .A1(n39724), .A2(n18871), .ZN(n14489) );
  INV_X1 U259 ( .I(n33100), .ZN(n1415) );
  AOI22_X1 U169 ( .A1(n17771), .A2(n31378), .B1(n12061), .B2(n9355), .ZN(n309)
         );
  AOI22_X1 U10973 ( .A1(n11488), .A2(n34007), .B1(n1189), .B2(n28528), .ZN(
        n8853) );
  NAND3_X1 U15257 ( .A1(n28501), .A2(n38145), .A3(n2790), .ZN(n2789) );
  NAND2_X1 U8961 ( .A1(n28515), .A2(n5093), .ZN(n4429) );
  NAND2_X1 U22712 ( .A1(n33318), .A2(n13508), .ZN(n11869) );
  OAI21_X1 U27685 ( .A1(n1420), .A2(n37204), .B(n19668), .ZN(n28568) );
  INV_X1 U4486 ( .I(n28463), .ZN(n28641) );
  NAND3_X1 U25301 ( .A1(n28495), .A2(n35173), .A3(n28356), .ZN(n28357) );
  INV_X1 U2247 ( .I(n29042), .ZN(n15480) );
  INV_X1 U2236 ( .I(n9393), .ZN(n21299) );
  INV_X1 U8921 ( .I(n14076), .ZN(n16116) );
  INV_X1 U8911 ( .I(n29344), .ZN(n29481) );
  INV_X1 U16871 ( .I(n4392), .ZN(n19693) );
  INV_X2 U7439 ( .I(n14400), .ZN(n1401) );
  INV_X2 U6572 ( .I(n14559), .ZN(n1181) );
  INV_X2 U20669 ( .I(n29195), .ZN(n29702) );
  INV_X1 U10828 ( .I(n9716), .ZN(n13136) );
  INV_X1 U4263 ( .I(n6163), .ZN(n29182) );
  OAI21_X1 U10789 ( .A1(n33784), .A2(n30241), .B(n6443), .ZN(n5306) );
  AOI21_X1 U23491 ( .A1(n29287), .A2(n29286), .B(n17225), .ZN(n12372) );
  NAND2_X1 U29742 ( .A1(n29102), .A2(n1175), .ZN(n29103) );
  INV_X2 U23554 ( .I(n30178), .ZN(n30183) );
  INV_X1 U25 ( .I(n18896), .ZN(n18897) );
  INV_X1 U8836 ( .I(n30184), .ZN(n16676) );
  INV_X1 U32 ( .I(n30097), .ZN(n1380) );
  INV_X1 U7379 ( .I(n29855), .ZN(n1171) );
  INV_X1 U5838 ( .I(n2858), .ZN(n3725) );
  NOR3_X1 U4996 ( .A1(n633), .A2(n1171), .A3(n32258), .ZN(n9676) );
  AND2_X1 U3 ( .A1(n12979), .A2(n29220), .Z(n9606) );
  INV_X1 U19 ( .I(n20538), .ZN(n30822) );
  INV_X1 U40 ( .I(n30079), .ZN(n30793) );
  INV_X1 U43 ( .I(n6205), .ZN(n1054) );
  NAND2_X1 U64 ( .A1(n31717), .A2(n14788), .ZN(n31532) );
  NOR2_X1 U82 ( .A1(n621), .A2(n20616), .ZN(n4075) );
  AND2_X1 U88 ( .A1(n29481), .A2(n29454), .Z(n29425) );
  OAI21_X1 U91 ( .A1(n39392), .A2(n12081), .B(n29061), .ZN(n400) );
  NAND3_X1 U92 ( .A1(n32894), .A2(n3986), .A3(n621), .ZN(n31170) );
  NAND2_X1 U135 ( .A1(n29445), .A2(n29446), .ZN(n5336) );
  NAND2_X1 U137 ( .A1(n8726), .A2(n29346), .ZN(n29349) );
  NAND2_X1 U139 ( .A1(n29384), .A2(n11084), .ZN(n31280) );
  AOI21_X1 U162 ( .A1(n29591), .A2(n29592), .B(n29598), .ZN(n31374) );
  NAND2_X1 U181 ( .A1(n11389), .A2(n9955), .ZN(n31550) );
  NAND2_X1 U191 ( .A1(n31313), .A2(n89), .ZN(n5543) );
  NAND2_X1 U269 ( .A1(n6405), .A2(n28434), .ZN(n31389) );
  NAND2_X1 U270 ( .A1(n7324), .A2(n28617), .ZN(n30857) );
  NOR2_X1 U274 ( .A1(n3014), .A2(n6426), .ZN(n32274) );
  AND2_X1 U362 ( .A1(n1446), .A2(n20577), .Z(n30357) );
  OR2_X1 U364 ( .A1(n28114), .A2(n28248), .Z(n30293) );
  NAND2_X1 U372 ( .A1(n32963), .A2(n33321), .ZN(n18341) );
  NAND3_X1 U391 ( .A1(n3983), .A2(n19996), .A3(n28279), .ZN(n7186) );
  NOR2_X1 U397 ( .A1(n5062), .A2(n28194), .ZN(n5910) );
  NAND2_X1 U398 ( .A1(n33669), .A2(n2877), .ZN(n33959) );
  NOR2_X1 U410 ( .A1(n28050), .A2(n11891), .ZN(n32479) );
  NAND3_X1 U422 ( .A1(n1453), .A2(n982), .A3(n2302), .ZN(n3097) );
  NOR2_X1 U429 ( .A1(n28246), .A2(n28247), .ZN(n32657) );
  NAND2_X1 U447 ( .A1(n27888), .A2(n28238), .ZN(n33199) );
  NOR2_X1 U452 ( .A1(n1072), .A2(n34008), .ZN(n14263) );
  INV_X1 U455 ( .I(n27948), .ZN(n33321) );
  NAND2_X1 U462 ( .A1(n1074), .A2(n28181), .ZN(n30799) );
  NOR2_X1 U466 ( .A1(n13081), .A2(n14399), .ZN(n12475) );
  NAND2_X1 U486 ( .A1(n1202), .A2(n11676), .ZN(n33931) );
  NAND2_X1 U500 ( .A1(n28102), .A2(n32352), .ZN(n33201) );
  INV_X1 U516 ( .I(n9470), .ZN(n8960) );
  NOR2_X1 U528 ( .A1(n28238), .A2(n1453), .ZN(n33202) );
  BUF_X2 U539 ( .I(n28153), .Z(n33481) );
  BUF_X2 U563 ( .I(n10009), .Z(n9534) );
  INV_X1 U581 ( .I(n27631), .ZN(n31218) );
  NAND2_X1 U654 ( .A1(n7606), .A2(n16520), .ZN(n16514) );
  NOR2_X1 U715 ( .A1(n31006), .A2(n17072), .ZN(n31399) );
  NOR2_X1 U723 ( .A1(n16482), .A2(n5772), .ZN(n31680) );
  AND2_X1 U767 ( .A1(n30986), .A2(n35427), .Z(n3605) );
  OR2_X1 U810 ( .A1(n26687), .A2(n17097), .Z(n30335) );
  OR2_X1 U812 ( .A1(n26979), .A2(n852), .Z(n30352) );
  OAI22_X1 U843 ( .A1(n27014), .A2(n11679), .B1(n27013), .B2(n38577), .ZN(
        n32549) );
  NAND2_X1 U846 ( .A1(n26815), .A2(n26973), .ZN(n26816) );
  AOI21_X1 U849 ( .A1(n20699), .A2(n849), .B(n7516), .ZN(n212) );
  NOR2_X1 U854 ( .A1(n26718), .A2(n735), .ZN(n33303) );
  NOR2_X1 U855 ( .A1(n13393), .A2(n26764), .ZN(n32669) );
  NOR2_X1 U868 ( .A1(n16160), .A2(n866), .ZN(n17279) );
  AOI21_X1 U902 ( .A1(n18226), .A2(n26833), .B(n26628), .ZN(n30983) );
  INV_X1 U942 ( .I(n26899), .ZN(n32016) );
  NOR2_X1 U963 ( .A1(n875), .A2(n26937), .ZN(n11325) );
  NAND2_X1 U964 ( .A1(n26752), .A2(n26751), .ZN(n33708) );
  OR2_X1 U979 ( .A1(n26818), .A2(n4599), .Z(n13219) );
  NAND2_X1 U1022 ( .A1(n31919), .A2(n4769), .ZN(n8295) );
  OAI21_X1 U1032 ( .A1(n10179), .A2(n10180), .B(n1101), .ZN(n20116) );
  AOI21_X1 U1049 ( .A1(n603), .A2(n34961), .B(n26005), .ZN(n33891) );
  NAND2_X2 U1059 ( .A1(n20849), .A2(n5236), .ZN(n2150) );
  NAND2_X1 U1075 ( .A1(n7767), .A2(n8481), .ZN(n31919) );
  NOR2_X1 U1083 ( .A1(n15085), .A2(n15121), .ZN(n10180) );
  NAND2_X1 U1096 ( .A1(n36546), .A2(n31192), .ZN(n30547) );
  NAND2_X1 U1106 ( .A1(n26063), .A2(n25345), .ZN(n25348) );
  NOR2_X1 U1110 ( .A1(n26063), .A2(n26061), .ZN(n33465) );
  NOR2_X1 U1113 ( .A1(n17212), .A2(n7767), .ZN(n25818) );
  NAND2_X1 U1119 ( .A1(n16407), .A2(n18320), .ZN(n25586) );
  NOR2_X1 U1126 ( .A1(n36666), .A2(n5126), .ZN(n4867) );
  NAND2_X1 U1169 ( .A1(n35138), .A2(n33514), .ZN(n2942) );
  NOR2_X1 U1182 ( .A1(n603), .A2(n12548), .ZN(n30695) );
  NAND2_X1 U1198 ( .A1(n30625), .A2(n6939), .ZN(n7136) );
  OAI21_X1 U1199 ( .A1(n31388), .A2(n31386), .B(n25755), .ZN(n25758) );
  OAI21_X1 U1207 ( .A1(n25008), .A2(n20052), .B(n10082), .ZN(n30625) );
  NOR2_X1 U1211 ( .A1(n25753), .A2(n38338), .ZN(n31388) );
  OAI21_X1 U1222 ( .A1(n31809), .A2(n25460), .B(n17183), .ZN(n31843) );
  NOR2_X1 U1233 ( .A1(n25337), .A2(n12828), .ZN(n31842) );
  NAND2_X1 U1263 ( .A1(n25469), .A2(n25468), .ZN(n30936) );
  NAND2_X1 U1266 ( .A1(n3568), .A2(n38661), .ZN(n11243) );
  NOR2_X1 U1280 ( .A1(n4384), .A2(n37795), .ZN(n25536) );
  NOR2_X1 U1307 ( .A1(n2250), .A2(n15515), .ZN(n33250) );
  NOR2_X1 U1308 ( .A1(n15422), .A2(n14779), .ZN(n3319) );
  AND2_X1 U1329 ( .A1(n3568), .A2(n5051), .Z(n30388) );
  NAND2_X1 U1373 ( .A1(n25615), .A2(n19264), .ZN(n33648) );
  BUF_X2 U1493 ( .I(n25132), .Z(n33208) );
  NAND2_X1 U1528 ( .A1(n37852), .A2(n24866), .ZN(n6934) );
  NOR2_X1 U1545 ( .A1(n30843), .A2(n31861), .ZN(n33125) );
  OAI21_X1 U1553 ( .A1(n30948), .A2(n30947), .B(n1271), .ZN(n24502) );
  NOR2_X1 U1557 ( .A1(n24759), .A2(n12633), .ZN(n32971) );
  NAND2_X1 U1559 ( .A1(n24621), .A2(n10116), .ZN(n32062) );
  AND2_X1 U1561 ( .A1(n8173), .A2(n30464), .Z(n24771) );
  NAND2_X1 U1563 ( .A1(n24824), .A2(n30845), .ZN(n24387) );
  AND2_X1 U1569 ( .A1(n36321), .A2(n7445), .Z(n8804) );
  NOR2_X1 U1584 ( .A1(n1581), .A2(n7770), .ZN(n12681) );
  AND2_X1 U1593 ( .A1(n31650), .A2(n17806), .Z(n31530) );
  NAND2_X1 U1594 ( .A1(n3076), .A2(n24668), .ZN(n30915) );
  INV_X2 U1595 ( .I(n2341), .ZN(n24664) );
  NOR2_X1 U1602 ( .A1(n24680), .A2(n24883), .ZN(n6707) );
  NAND2_X1 U1616 ( .A1(n19828), .A2(n30464), .ZN(n32618) );
  NAND3_X1 U1617 ( .A1(n38194), .A2(n36471), .A3(n35901), .ZN(n24574) );
  NAND2_X1 U1685 ( .A1(n23817), .A2(n37134), .ZN(n30766) );
  OAI21_X1 U1692 ( .A1(n17709), .A2(n14378), .B(n1586), .ZN(n11317) );
  NAND2_X1 U1701 ( .A1(n37732), .A2(n20083), .ZN(n31044) );
  OAI21_X1 U1702 ( .A1(n16366), .A2(n24406), .B(n18920), .ZN(n31175) );
  NAND2_X1 U1715 ( .A1(n21043), .A2(n32899), .ZN(n24424) );
  NAND2_X1 U1732 ( .A1(n32742), .A2(n4986), .ZN(n32741) );
  NAND2_X1 U1735 ( .A1(n16918), .A2(n30927), .ZN(n23993) );
  NAND2_X1 U1743 ( .A1(n24478), .A2(n24479), .ZN(n32784) );
  NAND2_X1 U1744 ( .A1(n12975), .A2(n24433), .ZN(n30646) );
  NOR2_X1 U1749 ( .A1(n1282), .A2(n20404), .ZN(n31921) );
  AOI21_X1 U1752 ( .A1(n626), .A2(n24245), .B(n959), .ZN(n24094) );
  NAND2_X1 U1754 ( .A1(n17546), .A2(n24465), .ZN(n33904) );
  NAND2_X1 U1755 ( .A1(n30463), .A2(n30580), .ZN(n31102) );
  AND2_X1 U1772 ( .A1(n10477), .A2(n30311), .Z(n32786) );
  BUF_X2 U1778 ( .I(n19295), .Z(n32899) );
  INV_X1 U1793 ( .I(n30280), .ZN(n30320) );
  OAI21_X1 U1856 ( .A1(n21019), .A2(n23467), .B(n31223), .ZN(n23422) );
  NAND3_X1 U1861 ( .A1(n1310), .A2(n35232), .A3(n14011), .ZN(n13580) );
  NAND3_X1 U1870 ( .A1(n35367), .A2(n23577), .A3(n20955), .ZN(n20954) );
  AND2_X1 U1874 ( .A1(n23631), .A2(n11342), .Z(n20841) );
  NAND2_X1 U1887 ( .A1(n23355), .A2(n31749), .ZN(n14576) );
  OAI21_X1 U1920 ( .A1(n32798), .A2(n23455), .B(n33080), .ZN(n20984) );
  AND2_X1 U1935 ( .A1(n33496), .A2(n23619), .Z(n30460) );
  OAI21_X1 U1946 ( .A1(n23552), .A2(n37814), .B(n14163), .ZN(n30548) );
  AOI21_X1 U1957 ( .A1(n22845), .A2(n22682), .B(n15242), .ZN(n15771) );
  INV_X1 U1963 ( .I(n3256), .ZN(n5492) );
  INV_X1 U1971 ( .I(n23121), .ZN(n9238) );
  NAND2_X1 U1974 ( .A1(n31351), .A2(n33247), .ZN(n19521) );
  NAND3_X1 U1979 ( .A1(n23175), .A2(n121), .A3(n3803), .ZN(n11472) );
  AOI22_X1 U1984 ( .A1(n23149), .A2(n1146), .B1(n14234), .B2(n38604), .ZN(
        n10699) );
  NAND2_X1 U1989 ( .A1(n22709), .A2(n1651), .ZN(n15344) );
  OAI21_X1 U1991 ( .A1(n14409), .A2(n32677), .B(n32676), .ZN(n23207) );
  NOR2_X1 U2016 ( .A1(n14396), .A2(n33745), .ZN(n9770) );
  NOR2_X1 U2017 ( .A1(n18515), .A2(n19945), .ZN(n32216) );
  NOR2_X1 U2018 ( .A1(n19698), .A2(n23101), .ZN(n33074) );
  NOR2_X1 U2035 ( .A1(n32636), .A2(n23149), .ZN(n12239) );
  OAI21_X1 U2036 ( .A1(n15033), .A2(n22932), .B(n39527), .ZN(n15032) );
  INV_X1 U2050 ( .I(n22559), .ZN(n33694) );
  INV_X1 U2051 ( .I(n12437), .ZN(n22575) );
  NOR2_X1 U2068 ( .A1(n22676), .A2(n1670), .ZN(n17341) );
  NAND3_X1 U2084 ( .A1(n22299), .A2(n22301), .A3(n22300), .ZN(n22302) );
  INV_X1 U2103 ( .I(n30818), .ZN(n30817) );
  INV_X1 U2108 ( .I(n22262), .ZN(n22125) );
  NOR2_X1 U2123 ( .A1(n3003), .A2(n22229), .ZN(n31859) );
  AOI21_X1 U2124 ( .A1(n22234), .A2(n20351), .B(n7497), .ZN(n33859) );
  INV_X1 U2130 ( .I(n33678), .ZN(n16635) );
  INV_X2 U2139 ( .I(n22234), .ZN(n33860) );
  AOI21_X1 U2164 ( .A1(n19377), .A2(n19376), .B(n21894), .ZN(n21369) );
  NOR2_X1 U2166 ( .A1(n21670), .A2(n6198), .ZN(n33636) );
  AND2_X1 U2167 ( .A1(n35921), .A2(n21903), .Z(n30397) );
  NOR2_X1 U2171 ( .A1(n14424), .A2(n21788), .ZN(n32857) );
  NOR2_X1 U2181 ( .A1(n18417), .A2(n30731), .ZN(n31975) );
  NOR2_X1 U2188 ( .A1(n31335), .A2(n21888), .ZN(n21333) );
  NAND2_X1 U2197 ( .A1(n35921), .A2(n18152), .ZN(n33731) );
  NOR2_X2 U2211 ( .A1(n38782), .A2(n16677), .ZN(n17816) );
  INV_X2 U2220 ( .I(n5871), .ZN(n24738) );
  NAND2_X2 U2230 ( .A1(n16990), .A2(n5871), .ZN(n7847) );
  INV_X2 U2232 ( .I(n15350), .ZN(n21987) );
  NAND2_X2 U2262 ( .A1(n18831), .A2(n25557), .ZN(n13988) );
  NOR2_X2 U2265 ( .A1(n30851), .A2(n35904), .ZN(n19569) );
  INV_X2 U2270 ( .I(n25718), .ZN(n25563) );
  INV_X2 U2281 ( .I(n14350), .ZN(n25009) );
  BUF_X4 U2308 ( .I(n21445), .Z(n21847) );
  OAI21_X2 U2317 ( .A1(n10374), .A2(n12671), .B(n25048), .ZN(n10373) );
  CLKBUF_X4 U2330 ( .I(n30095), .Z(n6147) );
  NAND2_X1 U2377 ( .A1(n14076), .A2(n29493), .ZN(n29451) );
  NAND2_X1 U2387 ( .A1(n4083), .A2(n30195), .ZN(n1757) );
  AOI21_X1 U2405 ( .A1(n12320), .A2(n29441), .B(n12317), .ZN(n12316) );
  NOR2_X1 U2422 ( .A1(n28089), .A2(n288), .ZN(n8206) );
  AOI22_X1 U2431 ( .A1(n26826), .A2(n26825), .B1(n19442), .B2(n19762), .ZN(
        n20022) );
  OAI21_X1 U2435 ( .A1(n31283), .A2(n9249), .B(n3700), .ZN(n9248) );
  NAND2_X1 U2445 ( .A1(n9716), .A2(n1061), .ZN(n32649) );
  NAND3_X1 U2453 ( .A1(n6818), .A2(n1798), .A3(n33803), .ZN(n13292) );
  AOI21_X1 U2485 ( .A1(n3860), .A2(n29927), .B(n19097), .ZN(n29925) );
  NAND2_X1 U2490 ( .A1(n14949), .A2(n17072), .ZN(n17298) );
  AOI21_X1 U2499 ( .A1(n16917), .A2(n24443), .B(n1596), .ZN(n30927) );
  AOI21_X1 U2516 ( .A1(n6684), .A2(n6421), .B(n1637), .ZN(n23216) );
  BUF_X2 U2524 ( .I(Key[41]), .Z(n29964) );
  OAI21_X1 U2536 ( .A1(n31516), .A2(n29761), .B(n19599), .ZN(n7001) );
  NAND2_X1 U2592 ( .A1(n31889), .A2(n31888), .ZN(n31887) );
  CLKBUF_X2 U2601 ( .I(n15153), .Z(n31788) );
  AOI21_X1 U2611 ( .A1(n12303), .A2(n12302), .B(n9534), .ZN(n18497) );
  NOR2_X1 U2623 ( .A1(n982), .A2(n28236), .ZN(n27991) );
  OAI21_X1 U2629 ( .A1(n6181), .A2(n19318), .B(n39689), .ZN(n29646) );
  AND2_X1 U2645 ( .A1(n37085), .A2(n25421), .Z(n25612) );
  OR2_X1 U2647 ( .A1(n28962), .A2(n19599), .Z(n30391) );
  NAND2_X1 U2669 ( .A1(n25540), .A2(n30317), .ZN(n25474) );
  NOR2_X1 U2674 ( .A1(n14418), .A2(n19202), .ZN(n21536) );
  NOR2_X1 U2675 ( .A1(n19202), .A2(n13285), .ZN(n32372) );
  OR2_X1 U2701 ( .A1(n5348), .A2(n19458), .Z(n4169) );
  INV_X1 U2705 ( .I(n38584), .ZN(n1502) );
  INV_X1 U2721 ( .I(n7335), .ZN(n1628) );
  NAND2_X1 U2757 ( .A1(n33307), .A2(n28021), .ZN(n32963) );
  INV_X1 U2760 ( .I(n28676), .ZN(n28671) );
  CLKBUF_X4 U2771 ( .I(n17876), .Z(n14337) );
  NAND2_X1 U2804 ( .A1(n2717), .A2(n15925), .ZN(n30955) );
  NAND2_X1 U2808 ( .A1(n11125), .A2(n30165), .ZN(n30166) );
  NOR2_X1 U2840 ( .A1(n30716), .A2(n28454), .ZN(n32236) );
  NAND2_X1 U2850 ( .A1(n31307), .A2(n29367), .ZN(n29368) );
  NAND2_X1 U2857 ( .A1(n29412), .A2(n17849), .ZN(n15043) );
  NAND3_X1 U2886 ( .A1(n15345), .A2(n15344), .A3(n39034), .ZN(n15343) );
  NAND2_X1 U2898 ( .A1(n982), .A2(n17314), .ZN(n16851) );
  INV_X2 U2902 ( .I(n29660), .ZN(n1390) );
  INV_X1 U2907 ( .I(n2296), .ZN(n29593) );
  AOI21_X1 U2921 ( .A1(n27292), .A2(n27221), .B(n39546), .ZN(n27018) );
  NOR2_X1 U2926 ( .A1(n13981), .A2(n12943), .ZN(n12942) );
  AOI21_X1 U2934 ( .A1(n6036), .A2(n22156), .B(n37199), .ZN(n667) );
  OAI22_X1 U2936 ( .A1(n22048), .A2(n16935), .B1(n36151), .B2(n6036), .ZN(
        n14957) );
  NOR2_X1 U2945 ( .A1(n1178), .A2(n17105), .ZN(n7002) );
  AOI22_X1 U2946 ( .A1(n29762), .A2(n29764), .B1(n29696), .B2(n17105), .ZN(
        n7003) );
  NAND3_X1 U2949 ( .A1(n30793), .A2(n30078), .A3(n30077), .ZN(n30075) );
  OAI22_X1 U3046 ( .A1(n19945), .A2(n17080), .B1(n17918), .B2(n17021), .ZN(
        n22845) );
  NOR2_X1 U3065 ( .A1(n9329), .A2(n38162), .ZN(n9352) );
  NAND2_X1 U3074 ( .A1(n32601), .A2(n23473), .ZN(n32630) );
  CLKBUF_X1 U3079 ( .I(n37632), .Z(n31160) );
  INV_X2 U3080 ( .I(n13799), .ZN(n14400) );
  INV_X1 U3089 ( .I(n26713), .ZN(n26849) );
  INV_X1 U3092 ( .I(n18711), .ZN(n22245) );
  INV_X1 U3100 ( .I(n36798), .ZN(n18801) );
  NAND2_X1 U3129 ( .A1(n22204), .A2(n16265), .ZN(n22206) );
  NAND2_X1 U3130 ( .A1(n22204), .A2(n16265), .ZN(n16262) );
  NOR2_X1 U3151 ( .A1(n36340), .A2(n19901), .ZN(n7154) );
  INV_X2 U3155 ( .I(n35443), .ZN(n24792) );
  NAND2_X1 U3160 ( .A1(n14400), .A2(n9733), .ZN(n18140) );
  OAI21_X1 U3161 ( .A1(n30144), .A2(n30132), .B(n35234), .ZN(n30133) );
  NOR2_X1 U3168 ( .A1(n29975), .A2(n29980), .ZN(n19041) );
  INV_X2 U3176 ( .I(n10907), .ZN(n10906) );
  INV_X1 U3199 ( .I(n7485), .ZN(n10494) );
  NOR2_X1 U3200 ( .A1(n35367), .A2(n7485), .ZN(n32363) );
  AOI21_X1 U3203 ( .A1(n23572), .A2(n7485), .B(n23571), .ZN(n23367) );
  OAI21_X1 U3220 ( .A1(n13805), .A2(n21684), .B(n21431), .ZN(n21416) );
  NAND2_X1 U3229 ( .A1(n26702), .A2(n6190), .ZN(n32261) );
  NAND2_X1 U3244 ( .A1(n24759), .A2(n10054), .ZN(n24762) );
  NAND2_X1 U3248 ( .A1(n14404), .A2(n11891), .ZN(n32059) );
  NAND2_X1 U3272 ( .A1(n28237), .A2(n14462), .ZN(n3779) );
  NAND2_X1 U3282 ( .A1(n306), .A2(n28677), .ZN(n28575) );
  OR2_X1 U3298 ( .A1(n27919), .A2(n20860), .Z(n27920) );
  NOR2_X1 U3305 ( .A1(n17989), .A2(n35755), .ZN(n7108) );
  INV_X1 U3332 ( .I(n3760), .ZN(n24685) );
  NAND2_X1 U3348 ( .A1(n25727), .A2(n16264), .ZN(n25730) );
  NOR2_X1 U3365 ( .A1(n4524), .A2(n37088), .ZN(n23253) );
  NOR2_X1 U3420 ( .A1(n18415), .A2(n18707), .ZN(n5437) );
  AOI22_X1 U3437 ( .A1(n12115), .A2(n1527), .B1(n31263), .B2(n38185), .ZN(
        n13280) );
  INV_X1 U3438 ( .I(n32243), .ZN(n13065) );
  AND2_X1 U3450 ( .A1(n36369), .A2(n2350), .Z(n30272) );
  INV_X2 U3453 ( .I(n8452), .ZN(n9854) );
  OR2_X1 U3456 ( .A1(n23531), .A2(n36539), .Z(n30275) );
  NOR2_X2 U3461 ( .A1(n23078), .A2(n23076), .ZN(n32878) );
  INV_X2 U3472 ( .I(n38749), .ZN(n32391) );
  XNOR2_X1 U3474 ( .A1(n23773), .A2(n23772), .ZN(n30280) );
  AND2_X1 U3493 ( .A1(n27181), .A2(n27180), .Z(n30288) );
  OR2_X1 U3533 ( .A1(n29641), .A2(n29660), .Z(n30295) );
  OR2_X2 U3539 ( .A1(n2047), .A2(n17169), .Z(n9651) );
  INV_X1 U3561 ( .I(n734), .ZN(n2366) );
  NAND2_X1 U3565 ( .A1(n28431), .A2(n28728), .ZN(n31889) );
  NAND2_X1 U3575 ( .A1(n8537), .A2(n19998), .ZN(n19997) );
  AND2_X2 U3602 ( .A1(n7666), .A2(n13794), .Z(n14525) );
  NAND2_X1 U3611 ( .A1(n36569), .A2(n11729), .ZN(n27415) );
  NOR2_X1 U3614 ( .A1(n6686), .A2(n11729), .ZN(n11728) );
  NOR2_X1 U3617 ( .A1(n9290), .A2(n38162), .ZN(n9353) );
  NAND3_X1 U3638 ( .A1(n28671), .A2(n36685), .A3(n1068), .ZN(n28678) );
  NOR2_X1 U3645 ( .A1(n3992), .A2(n2451), .ZN(n30825) );
  INV_X1 U3689 ( .I(n10621), .ZN(n10622) );
  INV_X2 U3700 ( .I(n4803), .ZN(n27951) );
  NOR2_X1 U3709 ( .A1(n11020), .A2(n27306), .ZN(n12214) );
  NAND2_X1 U3714 ( .A1(n9751), .A2(n19746), .ZN(n18880) );
  INV_X1 U3749 ( .I(n26115), .ZN(n25927) );
  NOR2_X1 U3750 ( .A1(n2561), .A2(n26115), .ZN(n2423) );
  AND2_X2 U3781 ( .A1(n8628), .A2(n16174), .Z(n17226) );
  NAND2_X1 U3805 ( .A1(n3313), .A2(n35198), .ZN(n27067) );
  NAND2_X1 U3808 ( .A1(n8173), .A2(n5957), .ZN(n14838) );
  AOI21_X1 U3840 ( .A1(n12952), .A2(n1145), .B(n35994), .ZN(n4895) );
  NAND2_X1 U3844 ( .A1(n257), .A2(n7810), .ZN(n24669) );
  CLKBUF_X1 U3895 ( .I(n34175), .Z(n33358) );
  BUF_X2 U3896 ( .I(n1418), .Z(n32014) );
  NAND2_X1 U3902 ( .A1(n274), .A2(n28278), .ZN(n31116) );
  OR2_X1 U3905 ( .A1(n33553), .A2(n10817), .Z(n10827) );
  CLKBUF_X1 U3910 ( .I(n19982), .Z(n30846) );
  NAND2_X1 U3937 ( .A1(n1008), .A2(n36873), .ZN(n32006) );
  NOR2_X1 U3938 ( .A1(n32170), .A2(n19338), .ZN(n32169) );
  OAI21_X1 U3943 ( .A1(n21041), .A2(n25912), .B(n32689), .ZN(n16952) );
  INV_X2 U3949 ( .I(n5356), .ZN(n1514) );
  NAND2_X1 U3959 ( .A1(n826), .A2(n9893), .ZN(n5860) );
  BUF_X2 U3960 ( .I(n15883), .Z(n10882) );
  INV_X1 U4004 ( .I(n23199), .ZN(n32872) );
  INV_X1 U4013 ( .I(n4846), .ZN(n33075) );
  BUF_X2 U4016 ( .I(n22925), .Z(n19535) );
  NAND2_X1 U4028 ( .A1(n1683), .A2(n17781), .ZN(n32803) );
  NOR2_X1 U4043 ( .A1(n11149), .A2(n17307), .ZN(n30826) );
  CLKBUF_X4 U4046 ( .I(n133), .Z(n32640) );
  NAND2_X1 U4047 ( .A1(n21751), .A2(n33876), .ZN(n31365) );
  NAND2_X1 U4059 ( .A1(n21676), .A2(n33053), .ZN(n33052) );
  NOR2_X1 U4062 ( .A1(n19641), .A2(n18143), .ZN(n31034) );
  INV_X1 U4066 ( .I(n29964), .ZN(n30324) );
  BUF_X2 U4067 ( .I(Key[58]), .Z(n19624) );
  NAND2_X1 U4076 ( .A1(n3465), .A2(n31160), .ZN(n31495) );
  INV_X2 U4084 ( .I(n29754), .ZN(n30555) );
  NAND2_X1 U4085 ( .A1(n31549), .A2(n30210), .ZN(n33520) );
  NAND2_X1 U4086 ( .A1(n20078), .A2(n30793), .ZN(n20949) );
  NAND2_X1 U4087 ( .A1(n20437), .A2(n29568), .ZN(n30496) );
  AOI22_X1 U4089 ( .A1(n4445), .A2(n5471), .B1(n19508), .B2(n2121), .ZN(n32192) );
  NOR2_X1 U4095 ( .A1(n34175), .A2(n19994), .ZN(n5001) );
  OR2_X1 U4103 ( .A1(n30160), .A2(n29185), .Z(n3958) );
  NAND2_X1 U4110 ( .A1(n29768), .A2(n29769), .ZN(n5762) );
  CLKBUF_X2 U4118 ( .I(n29941), .Z(n31629) );
  INV_X1 U4128 ( .I(n29249), .ZN(n31173) );
  NOR2_X1 U4149 ( .A1(n11028), .A2(n9141), .ZN(n30714) );
  NOR2_X1 U4158 ( .A1(n28749), .A2(n28748), .ZN(n33123) );
  NOR2_X1 U4166 ( .A1(n4228), .A2(n28356), .ZN(n5926) );
  NAND2_X1 U4172 ( .A1(n28443), .A2(n28444), .ZN(n33472) );
  NOR2_X1 U4176 ( .A1(n10305), .A2(n1418), .ZN(n32314) );
  INV_X1 U4179 ( .I(n20621), .ZN(n33555) );
  INV_X1 U4198 ( .I(n4232), .ZN(n33353) );
  OR2_X1 U4200 ( .A1(n11413), .A2(n20662), .Z(n11613) );
  CLKBUF_X2 U4205 ( .I(n28689), .Z(n31418) );
  NAND2_X1 U4207 ( .A1(n31118), .A2(n31116), .ZN(n13179) );
  NAND2_X1 U4219 ( .A1(n35827), .A2(n30955), .ZN(n5938) );
  NAND2_X1 U4234 ( .A1(n13623), .A2(n1069), .ZN(n31002) );
  INV_X1 U4238 ( .I(n31119), .ZN(n31118) );
  INV_X1 U4246 ( .I(n28247), .ZN(n31616) );
  NOR2_X1 U4248 ( .A1(n28123), .A2(n10836), .ZN(n32480) );
  CLKBUF_X2 U4260 ( .I(n28017), .Z(n18150) );
  CLKBUF_X2 U4284 ( .I(n15287), .Z(n31438) );
  CLKBUF_X4 U4285 ( .I(n27755), .Z(n33587) );
  AND3_X2 U4295 ( .A1(n17151), .A2(n15277), .A3(n15275), .Z(n31602) );
  NAND2_X1 U4304 ( .A1(n15748), .A2(n33017), .ZN(n33016) );
  NAND2_X1 U4314 ( .A1(n27113), .A2(n1481), .ZN(n32756) );
  INV_X1 U4324 ( .I(n26889), .ZN(n11432) );
  CLKBUF_X2 U4340 ( .I(n7632), .Z(n32020) );
  BUF_X2 U4349 ( .I(n37245), .Z(n5035) );
  NAND2_X1 U4365 ( .A1(n32006), .A2(n32005), .ZN(n9654) );
  NOR2_X1 U4372 ( .A1(n33802), .A2(n10754), .ZN(n21317) );
  NAND2_X1 U4374 ( .A1(n17449), .A2(n8010), .ZN(n17448) );
  INV_X1 U4377 ( .I(n26149), .ZN(n33026) );
  AND2_X1 U4388 ( .A1(n26918), .A2(n13393), .Z(n30363) );
  BUF_X2 U4396 ( .I(n10029), .Z(n15411) );
  CLKBUF_X2 U4417 ( .I(n755), .Z(n30942) );
  CLKBUF_X2 U4419 ( .I(n18210), .Z(n32009) );
  NAND2_X1 U4447 ( .A1(n25905), .A2(n25904), .ZN(n33630) );
  OR2_X1 U4459 ( .A1(n26005), .A2(n25856), .Z(n30468) );
  NOR2_X1 U4462 ( .A1(n17791), .A2(n31133), .ZN(n14680) );
  OR2_X1 U4464 ( .A1(n38548), .A2(n34217), .Z(n30425) );
  NOR2_X1 U4481 ( .A1(n26019), .A2(n5859), .ZN(n26022) );
  INV_X1 U4495 ( .I(n25108), .ZN(n31416) );
  NAND2_X1 U4498 ( .A1(n3278), .A2(n34087), .ZN(n31963) );
  NAND2_X1 U4503 ( .A1(n18145), .A2(n32355), .ZN(n20007) );
  OAI21_X1 U4505 ( .A1(n32291), .A2(n32279), .B(n32278), .ZN(n19501) );
  OR2_X1 U4507 ( .A1(n21254), .A2(n33242), .Z(n25724) );
  OR2_X1 U4513 ( .A1(n31895), .A2(n31587), .Z(n25444) );
  BUF_X2 U4520 ( .I(n25683), .Z(n30633) );
  OR2_X1 U4531 ( .A1(n10563), .A2(n25754), .Z(n30399) );
  BUF_X2 U4550 ( .I(n10686), .Z(n4467) );
  INV_X1 U4555 ( .I(n25239), .ZN(n32613) );
  CLKBUF_X4 U4562 ( .I(n25292), .Z(n30865) );
  BUF_X1 U4565 ( .I(n15186), .Z(n33439) );
  CLKBUF_X2 U4584 ( .I(n19691), .Z(n30733) );
  NAND2_X1 U4586 ( .A1(n7830), .A2(n5607), .ZN(n32368) );
  NAND2_X1 U4587 ( .A1(n31361), .A2(n31360), .ZN(n6081) );
  NAND2_X1 U4595 ( .A1(n32641), .A2(n24800), .ZN(n32644) );
  INV_X1 U4596 ( .I(n32641), .ZN(n24656) );
  INV_X1 U4620 ( .I(n8173), .ZN(n31713) );
  INV_X2 U4622 ( .I(n10931), .ZN(n33409) );
  CLKBUF_X2 U4624 ( .I(n24673), .Z(n33042) );
  NAND2_X1 U4631 ( .A1(n14283), .A2(n1028), .ZN(n16854) );
  OR2_X1 U4656 ( .A1(n37732), .A2(n21125), .Z(n30414) );
  INV_X1 U4672 ( .I(n7406), .ZN(n30647) );
  INV_X1 U4687 ( .I(n24483), .ZN(n33442) );
  NAND2_X1 U4691 ( .A1(n24100), .A2(n37467), .ZN(n24101) );
  CLKBUF_X2 U4704 ( .I(n19846), .Z(n32973) );
  INV_X1 U4709 ( .I(n23724), .ZN(n31178) );
  CLKBUF_X4 U4711 ( .I(n10638), .Z(n32776) );
  INV_X1 U4715 ( .I(n23911), .ZN(n1619) );
  INV_X1 U4716 ( .I(n2656), .ZN(n31927) );
  OR2_X1 U4725 ( .A1(n20817), .A2(n23516), .Z(n23265) );
  NAND2_X1 U4727 ( .A1(n2601), .A2(n17556), .ZN(n2598) );
  NAND2_X1 U4728 ( .A1(n33721), .A2(n23571), .ZN(n33720) );
  AND2_X1 U4736 ( .A1(n31586), .A2(n23456), .Z(n30440) );
  NOR2_X1 U4741 ( .A1(n20972), .A2(n23483), .ZN(n20991) );
  AND2_X1 U4742 ( .A1(n38535), .A2(n23516), .Z(n14649) );
  CLKBUF_X2 U4743 ( .I(n33703), .Z(n30499) );
  AND2_X1 U4751 ( .A1(n18199), .A2(n31906), .Z(n31949) );
  CLKBUF_X2 U4752 ( .I(n23607), .Z(n32246) );
  BUF_X2 U4753 ( .I(n23568), .Z(n31644) );
  OR2_X1 U4756 ( .A1(n16197), .A2(n14429), .Z(n30340) );
  NAND2_X1 U4768 ( .A1(n21292), .A2(n33414), .ZN(n22984) );
  OR2_X1 U4770 ( .A1(n23022), .A2(n1655), .Z(n7751) );
  CLKBUF_X2 U4774 ( .I(n4862), .Z(n32270) );
  INV_X1 U4778 ( .I(n22932), .ZN(n33554) );
  AND2_X1 U4783 ( .A1(n19134), .A2(n23124), .Z(n30360) );
  INV_X1 U4788 ( .I(n22990), .ZN(n17930) );
  CLKBUF_X2 U4792 ( .I(n17464), .Z(n31019) );
  CLKBUF_X2 U4793 ( .I(n782), .Z(n31093) );
  CLKBUF_X2 U4800 ( .I(n4997), .Z(n31838) );
  CLKBUF_X2 U4806 ( .I(n4291), .Z(n32796) );
  BUF_X2 U4809 ( .I(n23129), .Z(n19621) );
  INV_X1 U4818 ( .I(n10382), .ZN(n33273) );
  NOR2_X1 U4826 ( .A1(n16453), .A2(n16452), .ZN(n30798) );
  INV_X2 U4831 ( .I(n17942), .ZN(n30323) );
  INV_X1 U4832 ( .I(n33781), .ZN(n33780) );
  AOI21_X1 U4834 ( .A1(n31458), .A2(n17529), .B(n22289), .ZN(n2384) );
  NAND2_X1 U4837 ( .A1(n22266), .A2(n33282), .ZN(n21458) );
  NAND2_X1 U4840 ( .A1(n22050), .A2(n4200), .ZN(n30615) );
  INV_X2 U4844 ( .I(n22274), .ZN(n1676) );
  CLKBUF_X2 U4846 ( .I(n22219), .Z(n32408) );
  CLKBUF_X2 U4854 ( .I(n19518), .Z(n33489) );
  NOR2_X1 U4856 ( .A1(n21671), .A2(n6197), .ZN(n31972) );
  NAND2_X1 U4862 ( .A1(n33363), .A2(n21545), .ZN(n33700) );
  NAND2_X1 U4863 ( .A1(n21675), .A2(n19641), .ZN(n33054) );
  OAI21_X1 U4865 ( .A1(n18174), .A2(n36351), .B(n31034), .ZN(n6269) );
  CLKBUF_X2 U4869 ( .I(n21818), .Z(n19388) );
  CLKBUF_X2 U4873 ( .I(n18027), .Z(n32525) );
  CLKBUF_X2 U4877 ( .I(n21740), .Z(n19287) );
  INV_X1 U4878 ( .I(n19932), .ZN(n33515) );
  CLKBUF_X2 U4885 ( .I(n20887), .Z(n32138) );
  CLKBUF_X2 U4886 ( .I(n21823), .Z(n18143) );
  CLKBUF_X2 U4887 ( .I(n16333), .Z(n33280) );
  NAND2_X1 U4903 ( .A1(n15891), .A2(n21887), .ZN(n33876) );
  NOR2_X1 U4905 ( .A1(n14493), .A2(n19709), .ZN(n19708) );
  NOR2_X1 U4908 ( .A1(n19287), .A2(n38546), .ZN(n21391) );
  INV_X1 U4912 ( .I(n21814), .ZN(n21429) );
  NOR2_X1 U4921 ( .A1(n17265), .A2(n19274), .ZN(n12025) );
  NOR3_X1 U4928 ( .A1(n21681), .A2(n19262), .A3(n19768), .ZN(n18593) );
  NOR2_X1 U4937 ( .A1(n10961), .A2(n21810), .ZN(n36) );
  INV_X1 U4945 ( .I(n20368), .ZN(n15053) );
  NAND2_X1 U4955 ( .A1(n20996), .A2(n22047), .ZN(n21971) );
  INV_X1 U4960 ( .I(n19655), .ZN(n3001) );
  OR2_X1 U4998 ( .A1(n22298), .A2(n19778), .Z(n4280) );
  INV_X2 U5015 ( .I(n22067), .ZN(n10242) );
  INV_X1 U5018 ( .I(n22569), .ZN(n31012) );
  INV_X1 U5028 ( .I(n22463), .ZN(n9187) );
  CLKBUF_X1 U5045 ( .I(n33990), .Z(n32993) );
  NAND2_X1 U5055 ( .A1(n17021), .A2(n22682), .ZN(n18515) );
  INV_X1 U5068 ( .I(n23106), .ZN(n31947) );
  CLKBUF_X2 U5077 ( .I(n22837), .Z(n19788) );
  NOR2_X1 U5078 ( .A1(n12163), .A2(n23188), .ZN(n12699) );
  AOI21_X1 U5082 ( .A1(n11307), .A2(n23107), .B(n23111), .ZN(n33414) );
  NAND2_X1 U5104 ( .A1(n32042), .A2(n23060), .ZN(n32041) );
  NAND2_X1 U5109 ( .A1(n12083), .A2(n12028), .ZN(n31611) );
  NOR2_X1 U5188 ( .A1(n35689), .A2(n1642), .ZN(n21250) );
  AND3_X1 U5190 ( .A1(n1138), .A2(n10174), .A3(n23582), .Z(n30445) );
  AND3_X1 U5235 ( .A1(n17931), .A2(n23352), .A3(n13217), .Z(n30456) );
  OAI22_X1 U5249 ( .A1(n13150), .A2(n23578), .B1(n23506), .B2(n23580), .ZN(
        n20947) );
  AND3_X1 U5250 ( .A1(n15981), .A2(n17556), .A3(n1137), .Z(n789) );
  OAI21_X1 U5256 ( .A1(n13602), .A2(n23390), .B(n23452), .ZN(n4543) );
  AND2_X1 U5262 ( .A1(n18747), .A2(n23531), .Z(n30457) );
  AOI22_X1 U5268 ( .A1(n16716), .A2(n8692), .B1(n6176), .B2(n22513), .ZN(n6139) );
  INV_X1 U5276 ( .I(n20777), .ZN(n33573) );
  INV_X1 U5284 ( .I(n23841), .ZN(n23788) );
  INV_X1 U5286 ( .I(n23812), .ZN(n32097) );
  NAND2_X1 U5304 ( .A1(n24114), .A2(n30320), .ZN(n32742) );
  NOR2_X1 U5310 ( .A1(n24371), .A2(n18466), .ZN(n4784) );
  INV_X1 U5316 ( .I(n12975), .ZN(n20339) );
  INV_X1 U5353 ( .I(n24863), .ZN(n1566) );
  NAND2_X1 U5376 ( .A1(n1909), .A2(n38626), .ZN(n30635) );
  NOR2_X1 U5384 ( .A1(n24692), .A2(n24576), .ZN(n30642) );
  NAND2_X1 U5390 ( .A1(n16196), .A2(n30699), .ZN(n30698) );
  NAND2_X1 U5404 ( .A1(n12633), .A2(n24759), .ZN(n14267) );
  NOR2_X1 U5410 ( .A1(n8127), .A2(n12124), .ZN(n13638) );
  NAND2_X1 U5419 ( .A1(n958), .A2(n30642), .ZN(n6837) );
  INV_X1 U5433 ( .I(n33439), .ZN(n30649) );
  CLKBUF_X2 U5476 ( .I(n21254), .Z(n560) );
  INV_X2 U5482 ( .I(n13943), .ZN(n18294) );
  NOR2_X1 U5485 ( .A1(n31780), .A2(n19696), .ZN(n11268) );
  NOR2_X1 U5487 ( .A1(n25409), .A2(n25470), .ZN(n25410) );
  NAND2_X1 U5491 ( .A1(n4603), .A2(n31557), .ZN(n32355) );
  NAND3_X1 U5500 ( .A1(n9161), .A2(n17353), .A3(n32085), .ZN(n11847) );
  INV_X2 U5515 ( .I(n35828), .ZN(n26056) );
  INV_X1 U5596 ( .I(n19498), .ZN(n33216) );
  INV_X1 U5611 ( .I(n21098), .ZN(n17360) );
  INV_X1 U5619 ( .I(n33486), .ZN(n26308) );
  OAI21_X1 U5622 ( .A1(n31473), .A2(n1852), .B(n18801), .ZN(n1851) );
  NAND2_X1 U5632 ( .A1(n26708), .A2(n36355), .ZN(n32005) );
  NAND2_X1 U5636 ( .A1(n26700), .A2(n14636), .ZN(n17449) );
  NAND2_X1 U5639 ( .A1(n26645), .A2(n34005), .ZN(n19673) );
  NAND2_X1 U5643 ( .A1(n14412), .A2(n17158), .ZN(n32280) );
  INV_X1 U5645 ( .I(n26987), .ZN(n13949) );
  AND3_X1 U5647 ( .A1(n11864), .A2(n852), .A3(n26978), .Z(n30356) );
  NAND2_X1 U5660 ( .A1(n26831), .A2(n2882), .ZN(n3091) );
  INV_X1 U5712 ( .I(n15433), .ZN(n30811) );
  AOI21_X1 U5720 ( .A1(n31518), .A2(n21248), .B(n35265), .ZN(n27422) );
  NAND2_X1 U5731 ( .A1(n32169), .A2(n32167), .ZN(n32166) );
  NOR2_X1 U5737 ( .A1(n27372), .A2(n27269), .ZN(n3469) );
  INV_X1 U5797 ( .I(n3604), .ZN(n32021) );
  INV_X1 U5840 ( .I(n38213), .ZN(n31304) );
  INV_X1 U5851 ( .I(n33584), .ZN(n11947) );
  OAI21_X1 U5863 ( .A1(n37418), .A2(n36197), .B(n1076), .ZN(n31119) );
  NAND2_X1 U5875 ( .A1(n27877), .A2(n28001), .ZN(n27878) );
  INV_X1 U5904 ( .I(n28739), .ZN(n30581) );
  NAND2_X1 U5909 ( .A1(n30370), .A2(n28138), .ZN(n27966) );
  AOI21_X1 U5932 ( .A1(n4284), .A2(n1196), .B(n32575), .ZN(n30741) );
  NAND2_X1 U5947 ( .A1(n37204), .A2(n9668), .ZN(n19668) );
  NAND2_X1 U5983 ( .A1(n30741), .A2(n28682), .ZN(n33610) );
  INV_X1 U6016 ( .I(n28888), .ZN(n31398) );
  INV_X1 U6019 ( .I(n29099), .ZN(n31692) );
  NAND2_X1 U6025 ( .A1(n31699), .A2(n30380), .ZN(n7030) );
  NAND2_X1 U6068 ( .A1(n6443), .A2(n30242), .ZN(n29009) );
  AOI21_X1 U6070 ( .A1(n1175), .A2(n10590), .B(n29210), .ZN(n7899) );
  NAND2_X1 U6082 ( .A1(n9508), .A2(n5570), .ZN(n2861) );
  NOR2_X1 U6083 ( .A1(n7141), .A2(n3986), .ZN(n3170) );
  INV_X1 U6086 ( .I(n4169), .ZN(n18413) );
  OAI21_X1 U6090 ( .A1(n29699), .A2(n29701), .B(n29700), .ZN(n8345) );
  NAND2_X1 U6093 ( .A1(n775), .A2(n34652), .ZN(n33071) );
  CLKBUF_X1 U6101 ( .I(n29885), .Z(n31598) );
  INV_X1 U6103 ( .I(n10848), .ZN(n32706) );
  INV_X1 U6106 ( .I(n31532), .ZN(n31211) );
  NOR2_X1 U6109 ( .A1(n35176), .A2(n6252), .ZN(n29540) );
  OAI21_X1 U6114 ( .A1(n29732), .A2(n29755), .B(n29756), .ZN(n33766) );
  NAND2_X1 U6134 ( .A1(n6622), .A2(n29968), .ZN(n30709) );
  XNOR2_X1 U6166 ( .A1(n36750), .A2(n19908), .ZN(n30329) );
  XNOR2_X1 U6169 ( .A1(n35241), .A2(n27576), .ZN(n30333) );
  NOR2_X1 U6173 ( .A1(n26687), .A2(n26978), .ZN(n30336) );
  AND2_X1 U6179 ( .A1(n18186), .A2(n17598), .Z(n30339) );
  AND2_X1 U6191 ( .A1(n18197), .A2(n18198), .Z(n30342) );
  AND2_X1 U6194 ( .A1(n31594), .A2(n23380), .Z(n30345) );
  OR2_X1 U6207 ( .A1(n22051), .A2(n35755), .Z(n30354) );
  AND2_X1 U6215 ( .A1(n26973), .A2(n26974), .Z(n30355) );
  AND2_X1 U6234 ( .A1(n1212), .A2(n15357), .Z(n30369) );
  XNOR2_X1 U6236 ( .A1(n9611), .A2(n1358), .ZN(n30371) );
  AND2_X1 U6244 ( .A1(n19415), .A2(n12235), .Z(n30378) );
  NOR2_X1 U6264 ( .A1(n37067), .A2(n9197), .ZN(n30385) );
  OR2_X1 U6284 ( .A1(n18417), .A2(n19287), .Z(n30393) );
  AND2_X1 U6285 ( .A1(n14880), .A2(n33925), .Z(n30394) );
  XNOR2_X1 U6297 ( .A1(n22665), .A2(n28968), .ZN(n30402) );
  XNOR2_X1 U6302 ( .A1(n23880), .A2(n30120), .ZN(n30403) );
  XNOR2_X1 U6307 ( .A1(n13569), .A2(n37109), .ZN(n30404) );
  XNOR2_X1 U6309 ( .A1(n29831), .A2(n25160), .ZN(n30405) );
  XNOR2_X1 U6310 ( .A1(n22651), .A2(n29298), .ZN(n30406) );
  XNOR2_X1 U6322 ( .A1(n11923), .A2(n28831), .ZN(n30408) );
  XNOR2_X1 U6327 ( .A1(n19221), .A2(n965), .ZN(n30409) );
  AND3_X1 U6342 ( .A1(n1472), .A2(n32926), .A3(n27447), .Z(n30416) );
  OR2_X1 U6359 ( .A1(n23570), .A2(n17556), .Z(n30420) );
  INV_X1 U6364 ( .I(n21818), .ZN(n21817) );
  XOR2_X1 U6370 ( .A1(n20340), .A2(n20016), .Z(n30423) );
  INV_X1 U6375 ( .I(n30629), .ZN(n21039) );
  AND3_X2 U6380 ( .A1(n19470), .A2(n34016), .A3(n20694), .Z(n30427) );
  INV_X1 U6384 ( .I(n31473), .ZN(n9320) );
  INV_X2 U6386 ( .I(n23542), .ZN(n12154) );
  INV_X2 U6393 ( .I(n13442), .ZN(n15209) );
  AND2_X1 U6400 ( .A1(n28708), .A2(n28716), .Z(n30431) );
  AND2_X1 U6403 ( .A1(n16224), .A2(n29935), .Z(n30432) );
  NAND2_X1 U6410 ( .A1(n18077), .A2(n9781), .ZN(n31358) );
  XOR2_X1 U6431 ( .A1(n25279), .A2(n25281), .Z(n30433) );
  INV_X1 U6434 ( .I(n30117), .ZN(n30100) );
  XNOR2_X1 U6448 ( .A1(n25189), .A2(n35379), .ZN(n30435) );
  INV_X1 U6450 ( .I(n8745), .ZN(n3109) );
  INV_X1 U6486 ( .I(n21571), .ZN(n19271) );
  XNOR2_X1 U6496 ( .A1(n22630), .A2(n36362), .ZN(n30442) );
  INV_X2 U6499 ( .I(n5891), .ZN(n12952) );
  XNOR2_X1 U6506 ( .A1(n9982), .A2(n19902), .ZN(n30444) );
  XNOR2_X1 U6508 ( .A1(n23720), .A2(n23719), .ZN(n30446) );
  XNOR2_X1 U6511 ( .A1(n18582), .A2(n16893), .ZN(n30447) );
  INV_X1 U6512 ( .I(n4291), .ZN(n19698) );
  XNOR2_X1 U6514 ( .A1(n15608), .A2(n15607), .ZN(n30448) );
  XOR2_X1 U6519 ( .A1(n22479), .A2(n22478), .Z(n30450) );
  XOR2_X1 U6521 ( .A1(n23739), .A2(n23738), .Z(n30451) );
  XNOR2_X1 U6522 ( .A1(n23915), .A2(n23914), .ZN(n30452) );
  INV_X1 U6523 ( .I(n25683), .ZN(n25649) );
  OR3_X1 U6527 ( .A1(n4525), .A2(n20788), .A3(n37088), .Z(n30453) );
  INV_X1 U6534 ( .I(n23610), .ZN(n23292) );
  XNOR2_X1 U6541 ( .A1(n23715), .A2(n14220), .ZN(n30458) );
  XOR2_X1 U6549 ( .A1(n19775), .A2(n6185), .Z(n30459) );
  XOR2_X1 U6552 ( .A1(n15679), .A2(n19875), .Z(n30461) );
  INV_X1 U6568 ( .I(n25553), .ZN(n18704) );
  XNOR2_X1 U6573 ( .A1(n26520), .A2(n26551), .ZN(n30469) );
  XNOR2_X1 U6584 ( .A1(n8833), .A2(n30101), .ZN(n30471) );
  XNOR2_X1 U6592 ( .A1(n18399), .A2(n29238), .ZN(n30473) );
  XNOR2_X1 U6599 ( .A1(n35227), .A2(n15700), .ZN(n30478) );
  XNOR2_X1 U6600 ( .A1(n34332), .A2(n11994), .ZN(n30479) );
  XNOR2_X1 U6602 ( .A1(n1358), .A2(n9757), .ZN(n30480) );
  XNOR2_X1 U6605 ( .A1(n14566), .A2(n27578), .ZN(n30481) );
  XNOR2_X1 U6606 ( .A1(n27683), .A2(n19624), .ZN(n30482) );
  XNOR2_X1 U6610 ( .A1(n27683), .A2(n19583), .ZN(n30483) );
  XNOR2_X1 U6632 ( .A1(n38153), .A2(n31017), .ZN(n30487) );
  XNOR2_X1 U6635 ( .A1(n12430), .A2(n30094), .ZN(n30488) );
  INV_X2 U6636 ( .I(n20010), .ZN(n28149) );
  XNOR2_X1 U6641 ( .A1(n29087), .A2(n28834), .ZN(n30489) );
  OAI22_X1 U6659 ( .A1(n14075), .A2(n29571), .B1(n31899), .B2(n30496), .ZN(
        n14072) );
  NAND2_X2 U6676 ( .A1(n5424), .A2(n19771), .ZN(n28739) );
  XOR2_X1 U6683 ( .A1(n31370), .A2(n30433), .Z(n19582) );
  NAND2_X1 U6686 ( .A1(n6181), .A2(n19318), .ZN(n29648) );
  INV_X2 U6720 ( .I(n30503), .ZN(n12682) );
  AND2_X1 U6734 ( .A1(n2882), .A2(n7527), .Z(n26726) );
  INV_X2 U6737 ( .I(n33966), .ZN(n11898) );
  AOI21_X2 U6739 ( .A1(n37138), .A2(n22890), .B(n33361), .ZN(n30701) );
  NAND3_X2 U6789 ( .A1(n4484), .A2(n4483), .A3(n26547), .ZN(n4034) );
  AOI22_X2 U6791 ( .A1(n1746), .A2(n17530), .B1(n18303), .B2(n22042), .ZN(
        n22182) );
  XNOR2_X1 U6797 ( .A1(n3521), .A2(n30207), .ZN(n31830) );
  NAND2_X1 U6802 ( .A1(n3581), .A2(n7921), .ZN(n31302) );
  XOR2_X1 U6814 ( .A1(n30509), .A2(n12016), .Z(n10162) );
  XOR2_X1 U6815 ( .A1(n7582), .A2(n10163), .Z(n30509) );
  XOR2_X1 U6832 ( .A1(n23661), .A2(n31247), .Z(n722) );
  XOR2_X1 U6841 ( .A1(n30512), .A2(n19866), .Z(Ciphertext[147]) );
  OAI21_X2 U6880 ( .A1(n13398), .A2(n19670), .B(n30520), .ZN(n19807) );
  NAND2_X2 U6903 ( .A1(n24666), .A2(n24665), .ZN(n2653) );
  NOR2_X1 U6914 ( .A1(n12625), .A2(n16933), .ZN(n33251) );
  INV_X2 U6928 ( .I(n23352), .ZN(n31906) );
  XOR2_X1 U6934 ( .A1(n27524), .A2(n27204), .Z(n7061) );
  OR2_X1 U6951 ( .A1(n27969), .A2(n876), .Z(n18440) );
  XOR2_X1 U6958 ( .A1(n29095), .A2(n17880), .Z(n29835) );
  AOI21_X2 U6961 ( .A1(n28059), .A2(n28548), .B(n19354), .ZN(n29095) );
  NOR2_X1 U6964 ( .A1(n19891), .A2(n19605), .ZN(n15569) );
  OAI21_X2 U6967 ( .A1(n10626), .A2(n1588), .B(n30529), .ZN(n20326) );
  NAND2_X2 U7015 ( .A1(n10254), .A2(n19750), .ZN(n28052) );
  NAND2_X1 U7024 ( .A1(n38198), .A2(n39140), .ZN(n30611) );
  XOR2_X1 U7025 ( .A1(n26253), .A2(n26026), .Z(n26154) );
  OR2_X1 U7064 ( .A1(n29346), .A2(n29241), .Z(n13738) );
  XOR2_X1 U7122 ( .A1(n18642), .A2(n30541), .Z(n13410) );
  XOR2_X1 U7124 ( .A1(n25028), .A2(n25029), .Z(n30541) );
  XOR2_X1 U7165 ( .A1(n27651), .A2(n27649), .Z(n8281) );
  AOI21_X2 U7216 ( .A1(n30547), .A2(n30546), .B(n33795), .ZN(n20491) );
  XOR2_X1 U7240 ( .A1(n26227), .A2(n7602), .Z(n26145) );
  AND2_X1 U7285 ( .A1(n33147), .A2(n114), .Z(n3784) );
  XOR2_X1 U7326 ( .A1(n30551), .A2(n1980), .Z(n1978) );
  XOR2_X1 U7330 ( .A1(n31565), .A2(n10558), .Z(n13383) );
  AND2_X1 U7338 ( .A1(n23404), .A2(n2273), .Z(n2274) );
  XOR2_X1 U7343 ( .A1(n27769), .A2(n2582), .Z(n20341) );
  NOR2_X2 U7364 ( .A1(n33135), .A2(n13335), .ZN(n31944) );
  OR2_X1 U7367 ( .A1(n19941), .A2(n25581), .Z(n32172) );
  NAND2_X1 U7393 ( .A1(n4240), .A2(n32107), .ZN(n30558) );
  AOI21_X2 U7395 ( .A1(n18603), .A2(n20896), .B(n19242), .ZN(n15014) );
  XOR2_X1 U7397 ( .A1(n20586), .A2(n19936), .Z(n6768) );
  OAI21_X2 U7403 ( .A1(n31825), .A2(n30457), .B(n6611), .ZN(n20586) );
  XOR2_X1 U7425 ( .A1(n4476), .A2(n27847), .Z(n30560) );
  XOR2_X1 U7427 ( .A1(n30561), .A2(n14221), .Z(n2372) );
  XOR2_X1 U7428 ( .A1(n12741), .A2(n7489), .Z(n30561) );
  XOR2_X1 U7440 ( .A1(n30562), .A2(n13575), .Z(n24741) );
  XOR2_X1 U7462 ( .A1(n1504), .A2(n2150), .Z(n8075) );
  NOR3_X2 U7498 ( .A1(n19042), .A2(n31416), .A3(n18407), .ZN(n25111) );
  NAND2_X2 U7521 ( .A1(n10787), .A2(n10785), .ZN(n33440) );
  NAND2_X1 U7525 ( .A1(n24903), .A2(n37097), .ZN(n24906) );
  NOR2_X2 U7534 ( .A1(n2260), .A2(n2258), .ZN(n27828) );
  OAI21_X2 U7543 ( .A1(n5834), .A2(n9928), .B(n4713), .ZN(n11588) );
  XOR2_X1 U7556 ( .A1(n7089), .A2(n29246), .Z(n30578) );
  NAND2_X2 U7561 ( .A1(n18257), .A2(n3096), .ZN(n29789) );
  OAI22_X2 U7562 ( .A1(n3245), .A2(n3246), .B1(n3247), .B2(n19508), .ZN(n3096)
         );
  NOR2_X1 U7614 ( .A1(n32046), .A2(n32566), .ZN(n30582) );
  XOR2_X1 U7616 ( .A1(n29021), .A2(n18931), .Z(n29000) );
  AND2_X1 U7655 ( .A1(n21822), .A2(n21857), .Z(n21676) );
  INV_X2 U7656 ( .I(n19945), .ZN(n33361) );
  NOR3_X1 U7658 ( .A1(n1211), .A2(n31571), .A3(n30484), .ZN(n31808) );
  NAND2_X2 U7665 ( .A1(n17745), .A2(n17742), .ZN(n24011) );
  NAND2_X2 U7677 ( .A1(n24476), .A2(n24475), .ZN(n24784) );
  XOR2_X1 U7678 ( .A1(n3748), .A2(n3747), .Z(n13124) );
  NAND3_X1 U7682 ( .A1(n2861), .A2(n2859), .A3(n2860), .ZN(n30664) );
  OR2_X1 U7691 ( .A1(n840), .A2(n35828), .Z(n5680) );
  NAND3_X1 U7697 ( .A1(n25056), .A2(n37215), .A3(n25055), .ZN(n33176) );
  NAND2_X2 U7701 ( .A1(n32077), .A2(n6264), .ZN(n28695) );
  XOR2_X1 U7709 ( .A1(n30727), .A2(n29301), .Z(n30602) );
  XOR2_X1 U7711 ( .A1(n17567), .A2(n29054), .Z(n29301) );
  INV_X2 U7718 ( .I(n28660), .ZN(n28551) );
  AOI21_X2 U7744 ( .A1(n28743), .A2(n28742), .B(n30596), .ZN(n12430) );
  OAI22_X2 U7745 ( .A1(n30949), .A2(n31269), .B1(n28740), .B2(n28739), .ZN(
        n30596) );
  AOI22_X2 U7752 ( .A1(n13843), .A2(n24912), .B1(n30598), .B2(n36752), .ZN(
        n25026) );
  AOI21_X2 U7763 ( .A1(n8576), .A2(n17351), .B(n8575), .ZN(n12233) );
  AOI22_X2 U7764 ( .A1(n30599), .A2(n22882), .B1(n22881), .B2(n14402), .ZN(
        n23237) );
  XOR2_X1 U7770 ( .A1(n31535), .A2(n1365), .Z(n9164) );
  XOR2_X1 U7785 ( .A1(n30602), .A2(n18405), .Z(n4850) );
  NOR2_X2 U7801 ( .A1(n9178), .A2(n9188), .ZN(n18773) );
  NAND3_X1 U7805 ( .A1(n6569), .A2(n24381), .A3(n6570), .ZN(n30603) );
  XOR2_X1 U7834 ( .A1(n3557), .A2(n31304), .Z(n2159) );
  XOR2_X1 U7842 ( .A1(n32646), .A2(n29522), .Z(n33037) );
  OR2_X1 U7870 ( .A1(n31164), .A2(n31661), .Z(n11286) );
  XOR2_X1 U7872 ( .A1(n35053), .A2(n14374), .Z(n16190) );
  INV_X2 U7877 ( .I(n30607), .ZN(n31809) );
  NAND2_X2 U7914 ( .A1(n17214), .A2(n30608), .ZN(n7063) );
  XOR2_X1 U7921 ( .A1(n26523), .A2(n26526), .Z(n30609) );
  XOR2_X1 U7922 ( .A1(n38177), .A2(n16665), .Z(n30610) );
  AOI22_X1 U7932 ( .A1(n29577), .A2(n29565), .B1(n29566), .B2(n29563), .ZN(
        n31197) );
  OR2_X1 U7933 ( .A1(n13038), .A2(n39070), .Z(n31235) );
  XOR2_X1 U7949 ( .A1(n9947), .A2(n30482), .Z(n30781) );
  NAND3_X1 U7966 ( .A1(n29965), .A2(n1170), .A3(n29975), .ZN(n29966) );
  NAND2_X1 U7975 ( .A1(n31310), .A2(n1242), .ZN(n25454) );
  OAI21_X1 U7982 ( .A1(n29852), .A2(n11898), .B(n11897), .ZN(n30616) );
  XOR2_X1 U8002 ( .A1(n2825), .A2(n20446), .Z(n2824) );
  NAND2_X2 U8006 ( .A1(n15023), .A2(n14513), .ZN(n30894) );
  XOR2_X1 U8021 ( .A1(n22774), .A2(n706), .Z(n10237) );
  INV_X4 U8024 ( .I(n19828), .ZN(n24770) );
  XOR2_X1 U8032 ( .A1(n30619), .A2(n4616), .Z(n1794) );
  OAI21_X2 U8075 ( .A1(n13666), .A2(n8139), .B(n13664), .ZN(n25296) );
  XOR2_X1 U8084 ( .A1(n27835), .A2(n27836), .Z(n30626) );
  XNOR2_X1 U8093 ( .A1(n27697), .A2(n12999), .ZN(n32137) );
  OAI21_X2 U8152 ( .A1(n30353), .A2(n30886), .B(n29342), .ZN(n15768) );
  INV_X1 U8156 ( .I(n792), .ZN(n30632) );
  OAI22_X2 U8164 ( .A1(n8446), .A2(n8445), .B1(n32548), .B2(n39828), .ZN(
        n29885) );
  AND2_X1 U8176 ( .A1(n27198), .A2(n13973), .Z(n27031) );
  NAND2_X1 U8226 ( .A1(n32670), .A2(n29375), .ZN(n29315) );
  NAND3_X1 U8230 ( .A1(n30643), .A2(n26643), .A3(n6606), .ZN(n4484) );
  INV_X1 U8235 ( .I(n16466), .ZN(n30988) );
  XOR2_X1 U8245 ( .A1(n30645), .A2(n19624), .Z(Ciphertext[59]) );
  OAI21_X2 U8259 ( .A1(n33422), .A2(n29973), .B(n29971), .ZN(n32570) );
  OR2_X1 U8272 ( .A1(n23071), .A2(n14390), .Z(n32626) );
  XOR2_X1 U8278 ( .A1(n25009), .A2(n30649), .Z(n30648) );
  NOR2_X2 U8308 ( .A1(n30652), .A2(n16744), .ZN(n17101) );
  XOR2_X1 U8314 ( .A1(n28839), .A2(n28871), .Z(n27944) );
  NAND2_X2 U8334 ( .A1(n19661), .A2(n19360), .ZN(n18682) );
  NAND2_X1 U8359 ( .A1(n3218), .A2(n3217), .ZN(n30653) );
  XOR2_X1 U8401 ( .A1(n30657), .A2(n1365), .Z(Ciphertext[73]) );
  XOR2_X1 U8424 ( .A1(n24933), .A2(n25197), .Z(n25314) );
  NAND2_X2 U8425 ( .A1(n17962), .A2(n17963), .ZN(n24933) );
  XOR2_X1 U8462 ( .A1(n19374), .A2(n14221), .Z(n10156) );
  AOI21_X2 U8478 ( .A1(n30360), .A2(n272), .B(n30663), .ZN(n3047) );
  NAND2_X2 U8483 ( .A1(n30664), .A2(n2856), .ZN(n2858) );
  OAI21_X2 U8528 ( .A1(n27445), .A2(n27444), .B(n30667), .ZN(n27852) );
  XNOR2_X1 U8531 ( .A1(n23658), .A2(n23910), .ZN(n23740) );
  OAI21_X2 U8539 ( .A1(n13776), .A2(n5427), .B(n28269), .ZN(n30668) );
  NOR2_X1 U8572 ( .A1(n1470), .A2(n34279), .ZN(n7922) );
  NAND2_X2 U8577 ( .A1(n8506), .A2(n12510), .ZN(n27288) );
  XOR2_X1 U8611 ( .A1(n31782), .A2(n29022), .Z(n32604) );
  NOR2_X1 U8748 ( .A1(n29578), .A2(n28885), .ZN(n30675) );
  AND2_X1 U8749 ( .A1(n22407), .A2(n30676), .Z(n18166) );
  NAND2_X2 U8755 ( .A1(n4952), .A2(n30677), .ZN(n15085) );
  OR2_X1 U8799 ( .A1(n18519), .A2(n12162), .Z(n7235) );
  XNOR2_X1 U8803 ( .A1(n7247), .A2(n38184), .ZN(n30819) );
  NAND2_X1 U8820 ( .A1(n30454), .A2(n33734), .ZN(n24216) );
  INV_X1 U8840 ( .I(n16657), .ZN(n16655) );
  XOR2_X1 U8842 ( .A1(n31778), .A2(n19213), .Z(n31777) );
  XOR2_X1 U8846 ( .A1(n29257), .A2(n29031), .Z(n28041) );
  XOR2_X1 U8858 ( .A1(n12399), .A2(n12402), .Z(n12414) );
  XOR2_X1 U8862 ( .A1(n32795), .A2(n30682), .Z(n679) );
  AOI21_X2 U8892 ( .A1(n20863), .A2(n31270), .B(n30684), .ZN(n4670) );
  XOR2_X1 U8913 ( .A1(n8400), .A2(n30688), .Z(n30687) );
  XOR2_X1 U8918 ( .A1(n25156), .A2(n25043), .Z(n8702) );
  NAND2_X2 U8922 ( .A1(n3654), .A2(n3653), .ZN(n25043) );
  INV_X2 U8960 ( .I(n18480), .ZN(n2639) );
  INV_X1 U8962 ( .I(n32620), .ZN(n17426) );
  NAND2_X2 U8978 ( .A1(n19873), .A2(n34813), .ZN(n7768) );
  INV_X2 U8979 ( .I(n30701), .ZN(n71) );
  NOR2_X1 U8981 ( .A1(n2868), .A2(n19888), .ZN(n30702) );
  NAND2_X2 U8989 ( .A1(n30704), .A2(n11847), .ZN(n17212) );
  OAI21_X2 U8991 ( .A1(n16317), .A2(n16316), .B(n16315), .ZN(n30704) );
  INV_X1 U8992 ( .I(n31984), .ZN(n25362) );
  INV_X2 U8995 ( .I(n1666), .ZN(n22459) );
  XOR2_X1 U8998 ( .A1(n1666), .A2(n22503), .Z(n20753) );
  NOR2_X2 U8999 ( .A1(n30424), .A2(n30706), .ZN(n1666) );
  XOR2_X1 U9024 ( .A1(n27817), .A2(n18182), .Z(n32698) );
  XOR2_X1 U9038 ( .A1(n32621), .A2(n14872), .Z(n29500) );
  NOR2_X2 U9046 ( .A1(n20533), .A2(n30980), .ZN(n28715) );
  OAI22_X1 U9050 ( .A1(n5677), .A2(n19143), .B1(n30711), .B2(n30709), .ZN(
        n17030) );
  NOR2_X1 U9051 ( .A1(n1170), .A2(n6623), .ZN(n30711) );
  NAND3_X1 U9055 ( .A1(n5019), .A2(n13705), .A3(n5018), .ZN(n19252) );
  NOR2_X1 U9056 ( .A1(n35265), .A2(n27424), .ZN(n30712) );
  NOR2_X1 U9070 ( .A1(n19294), .A2(n24812), .ZN(n24615) );
  XOR2_X1 U9074 ( .A1(n22732), .A2(n4819), .Z(n4896) );
  OR2_X2 U9079 ( .A1(n9501), .A2(n9338), .Z(n9441) );
  XOR2_X1 U9080 ( .A1(n3028), .A2(n3029), .Z(n9501) );
  XNOR2_X1 U9107 ( .A1(n38181), .A2(n35249), .ZN(n10183) );
  OAI21_X1 U9125 ( .A1(n25469), .A2(n10004), .B(n25606), .ZN(n18249) );
  OR2_X1 U9143 ( .A1(n39489), .A2(n22250), .Z(n21090) );
  OR2_X1 U9178 ( .A1(n3369), .A2(n26691), .Z(n30726) );
  XOR2_X1 U9198 ( .A1(n15271), .A2(n29300), .Z(n30727) );
  XOR2_X1 U9217 ( .A1(n30730), .A2(n30065), .Z(Ciphertext[145]) );
  NAND2_X1 U9219 ( .A1(n33677), .A2(n33679), .ZN(n31379) );
  INV_X1 U9226 ( .I(n21387), .ZN(n21652) );
  NAND2_X1 U9232 ( .A1(n30731), .A2(n18417), .ZN(n14587) );
  XOR2_X1 U9233 ( .A1(n21386), .A2(Key[125]), .Z(n21387) );
  AOI21_X2 U9238 ( .A1(n30392), .A2(n18298), .B(n17182), .ZN(n2167) );
  NAND2_X2 U9240 ( .A1(n16289), .A2(n16290), .ZN(n22274) );
  INV_X2 U9262 ( .I(n2457), .ZN(n20749) );
  NAND2_X2 U9266 ( .A1(n27895), .A2(n28290), .ZN(n2457) );
  NAND2_X1 U9267 ( .A1(n231), .A2(n26268), .ZN(n33142) );
  XOR2_X1 U9270 ( .A1(n16334), .A2(n30734), .Z(n19639) );
  XOR2_X1 U9272 ( .A1(n19405), .A2(n29131), .Z(n30734) );
  NAND2_X2 U9284 ( .A1(n37245), .A2(n27211), .ZN(n27259) );
  INV_X2 U9289 ( .I(n30736), .ZN(n18721) );
  NAND2_X2 U9299 ( .A1(n30738), .A2(n16137), .ZN(n26009) );
  NAND2_X1 U9305 ( .A1(n25740), .A2(n12624), .ZN(n30738) );
  AND2_X1 U9317 ( .A1(n1131), .A2(n12064), .Z(n9460) );
  XOR2_X1 U9329 ( .A1(n5434), .A2(n11321), .Z(n32349) );
  NAND2_X1 U9358 ( .A1(n29762), .A2(n29761), .ZN(n30745) );
  XOR2_X1 U9404 ( .A1(Plaintext[89]), .A2(Key[89]), .Z(n21883) );
  NAND2_X2 U9428 ( .A1(n11148), .A2(n15575), .ZN(n25829) );
  INV_X4 U9444 ( .I(n33955), .ZN(n1446) );
  OAI21_X2 U9504 ( .A1(n1551), .A2(n15180), .B(n16234), .ZN(n25702) );
  XOR2_X1 U9512 ( .A1(n25285), .A2(n13530), .Z(n30756) );
  NAND2_X2 U9559 ( .A1(n17118), .A2(n1151), .ZN(n22178) );
  NAND2_X2 U9563 ( .A1(n19907), .A2(n19906), .ZN(n17118) );
  NOR2_X2 U9577 ( .A1(n24833), .A2(n31385), .ZN(n24755) );
  AOI21_X1 U9618 ( .A1(n39065), .A2(n27069), .B(n39417), .ZN(n3581) );
  INV_X1 U9657 ( .I(n34166), .ZN(n33842) );
  NAND2_X2 U9675 ( .A1(n1951), .A2(n4416), .ZN(n23931) );
  XOR2_X1 U9691 ( .A1(n24064), .A2(n23658), .Z(n23598) );
  XOR2_X1 U9700 ( .A1(n4896), .A2(n15311), .Z(n5540) );
  NAND2_X2 U9704 ( .A1(n3025), .A2(n3024), .ZN(n15311) );
  NAND2_X2 U9736 ( .A1(n12523), .A2(n12524), .ZN(n17455) );
  OAI21_X2 U9746 ( .A1(n28377), .A2(n28665), .B(n4002), .ZN(n9112) );
  XOR2_X1 U9747 ( .A1(n27759), .A2(n30771), .Z(n33373) );
  XOR2_X1 U9748 ( .A1(n27537), .A2(n37443), .Z(n30771) );
  NAND2_X2 U9769 ( .A1(n11083), .A2(n33662), .ZN(n27273) );
  AOI21_X2 U9777 ( .A1(n31130), .A2(n32725), .B(n13159), .ZN(n33662) );
  XOR2_X1 U9818 ( .A1(n26167), .A2(n19798), .Z(n30776) );
  XOR2_X1 U9827 ( .A1(n39723), .A2(n19676), .Z(n28958) );
  AOI21_X2 U9840 ( .A1(n6065), .A2(n13033), .B(n24963), .ZN(n30778) );
  OAI21_X2 U9856 ( .A1(n13469), .A2(n12475), .B(n28165), .ZN(n30780) );
  NAND2_X1 U9895 ( .A1(n26706), .A2(n26705), .ZN(n32347) );
  NAND2_X2 U9900 ( .A1(n3319), .A2(n30945), .ZN(n26115) );
  XOR2_X1 U9904 ( .A1(n10483), .A2(n31983), .Z(n4841) );
  NOR2_X1 U9920 ( .A1(n31755), .A2(n36623), .ZN(n30952) );
  OR2_X1 U9934 ( .A1(n29236), .A2(n8728), .Z(n14198) );
  AOI21_X1 U9942 ( .A1(n23467), .A2(n3256), .B(n18682), .ZN(n31223) );
  OAI22_X1 U9946 ( .A1(n5418), .A2(n28209), .B1(n28210), .B2(n28313), .ZN(
        n30785) );
  OR2_X1 U9969 ( .A1(n30764), .A2(n24719), .Z(n6540) );
  BUF_X4 U9986 ( .I(n20326), .Z(n6822) );
  OAI21_X2 U9990 ( .A1(n3600), .A2(n3671), .B(n3599), .ZN(n20078) );
  NAND2_X2 U9997 ( .A1(n30794), .A2(n10263), .ZN(n12892) );
  NAND2_X2 U10008 ( .A1(n17126), .A2(n13959), .ZN(n30794) );
  NOR2_X2 U10016 ( .A1(n30808), .A2(n5325), .ZN(n12667) );
  NOR2_X2 U10039 ( .A1(n30798), .A2(n16454), .ZN(n17605) );
  NAND2_X2 U10042 ( .A1(n21705), .A2(n21704), .ZN(n22204) );
  INV_X4 U10057 ( .I(n30800), .ZN(n22287) );
  XOR2_X1 U10112 ( .A1(n27464), .A2(n30803), .Z(n27029) );
  INV_X1 U10116 ( .I(n19816), .ZN(n30803) );
  NAND2_X2 U10125 ( .A1(n28539), .A2(n28495), .ZN(n11129) );
  XOR2_X1 U10145 ( .A1(n30806), .A2(n27816), .Z(n31996) );
  NAND2_X2 U10151 ( .A1(n26264), .A2(n15429), .ZN(n15434) );
  NAND2_X1 U10192 ( .A1(n19173), .A2(n29565), .ZN(n31284) );
  OAI22_X2 U10228 ( .A1(n15771), .A2(n15770), .B1(n18518), .B2(n22923), .ZN(
        n23354) );
  OAI21_X2 U10274 ( .A1(n32335), .A2(n2559), .B(n29583), .ZN(n2557) );
  XOR2_X1 U10300 ( .A1(n26274), .A2(n26223), .Z(n31627) );
  NOR2_X2 U10301 ( .A1(n16344), .A2(n19048), .ZN(n26274) );
  INV_X2 U10363 ( .I(n19746), .ZN(n15443) );
  XOR2_X1 U10398 ( .A1(n22625), .A2(n15610), .Z(n15609) );
  AOI22_X1 U10495 ( .A1(n29625), .A2(n29626), .B1(n29628), .B2(n29627), .ZN(
        n31366) );
  NAND2_X2 U10500 ( .A1(n1350), .A2(n39716), .ZN(n11378) );
  INV_X2 U10507 ( .I(n32474), .ZN(n19601) );
  NOR2_X2 U10514 ( .A1(n24495), .A2(n24496), .ZN(n24931) );
  XOR2_X1 U10572 ( .A1(n5252), .A2(n5251), .Z(n30831) );
  OAI21_X2 U10613 ( .A1(n12062), .A2(n19452), .B(n11860), .ZN(n26070) );
  NOR2_X1 U10639 ( .A1(n29498), .A2(n37614), .ZN(n29302) );
  XOR2_X1 U10646 ( .A1(n30318), .A2(n1260), .Z(n30838) );
  OAI21_X2 U10650 ( .A1(n27360), .A2(n32557), .B(n30840), .ZN(n2260) );
  XOR2_X1 U10668 ( .A1(n23917), .A2(n23953), .Z(n2120) );
  AOI21_X2 U10680 ( .A1(n29633), .A2(n20816), .B(n30847), .ZN(n19297) );
  OAI22_X2 U10682 ( .A1(n34089), .A2(n29632), .B1(n16385), .B2(n20982), .ZN(
        n30847) );
  XOR2_X1 U10683 ( .A1(n37699), .A2(n963), .Z(n10163) );
  OR2_X1 U10759 ( .A1(n23983), .A2(n16917), .Z(n12646) );
  OAI21_X1 U10761 ( .A1(n16502), .A2(n37640), .B(n30854), .ZN(n5123) );
  NAND2_X2 U10767 ( .A1(n22227), .A2(n7357), .ZN(n4316) );
  INV_X2 U10801 ( .I(n17984), .ZN(n30859) );
  INV_X4 U10803 ( .I(n22238), .ZN(n9546) );
  XOR2_X1 U10869 ( .A1(n4592), .A2(n9518), .Z(n16858) );
  OR2_X1 U10898 ( .A1(n12302), .A2(n4803), .Z(n11353) );
  INV_X1 U10908 ( .I(n36371), .ZN(n1334) );
  XOR2_X1 U10931 ( .A1(n16897), .A2(n18395), .Z(n15450) );
  NOR2_X2 U10932 ( .A1(n14935), .A2(n14934), .ZN(n18395) );
  XOR2_X1 U10943 ( .A1(n8775), .A2(n8773), .Z(n28843) );
  OR2_X1 U10954 ( .A1(n12331), .A2(n20449), .Z(n22554) );
  NAND2_X1 U10971 ( .A1(n15928), .A2(n21029), .ZN(n32663) );
  NAND2_X2 U10979 ( .A1(n20387), .A2(n20386), .ZN(n22776) );
  AOI21_X2 U10998 ( .A1(n29503), .A2(n29502), .B(n37374), .ZN(n29530) );
  NOR2_X1 U11000 ( .A1(n29501), .A2(n18190), .ZN(n30886) );
  XOR2_X1 U11012 ( .A1(n1259), .A2(n19359), .Z(n14639) );
  INV_X2 U11024 ( .I(n30890), .ZN(n826) );
  XOR2_X1 U11025 ( .A1(n13936), .A2(n13937), .Z(n30890) );
  NAND2_X2 U11028 ( .A1(n30323), .A2(n17943), .ZN(n22772) );
  XOR2_X1 U11031 ( .A1(n30891), .A2(n8631), .Z(n8824) );
  XOR2_X1 U11049 ( .A1(n33272), .A2(n30895), .Z(n33244) );
  XOR2_X1 U11050 ( .A1(n22321), .A2(n16531), .Z(n30895) );
  BUF_X2 U11052 ( .I(n24192), .Z(n30897) );
  NAND2_X1 U11078 ( .A1(n27411), .A2(n6355), .ZN(n10359) );
  INV_X2 U11117 ( .I(n30905), .ZN(n10817) );
  XOR2_X1 U11119 ( .A1(n10818), .A2(n10819), .Z(n30905) );
  NOR2_X1 U11123 ( .A1(n28396), .A2(n9848), .ZN(n28298) );
  XOR2_X1 U11162 ( .A1(n27675), .A2(n5697), .Z(n30907) );
  OAI21_X1 U11164 ( .A1(n1028), .A2(n24782), .B(n24545), .ZN(n16948) );
  NAND2_X2 U11172 ( .A1(n30908), .A2(n4568), .ZN(n11694) );
  INV_X1 U11180 ( .I(n13155), .ZN(n26509) );
  XOR2_X1 U11181 ( .A1(n19289), .A2(n13155), .Z(n12860) );
  XOR2_X1 U11190 ( .A1(n25144), .A2(n25299), .Z(n30910) );
  NAND2_X2 U11212 ( .A1(n30914), .A2(n24131), .ZN(n24887) );
  XOR2_X1 U11248 ( .A1(n1462), .A2(n17418), .Z(n18633) );
  NAND2_X2 U11315 ( .A1(n28573), .A2(n30928), .ZN(n29837) );
  NAND3_X1 U11318 ( .A1(n19321), .A2(n19322), .A3(n28666), .ZN(n30928) );
  OR2_X1 U11334 ( .A1(n691), .A2(n29548), .Z(n15174) );
  AOI21_X2 U11348 ( .A1(n27328), .A2(n27325), .B(n32555), .ZN(n30933) );
  XOR2_X1 U11373 ( .A1(n13969), .A2(n12775), .Z(n13332) );
  XOR2_X1 U11376 ( .A1(n11358), .A2(n30938), .Z(n9958) );
  XOR2_X1 U11378 ( .A1(n17621), .A2(n30487), .Z(n30938) );
  NAND2_X2 U11383 ( .A1(n30939), .A2(n27324), .ZN(n27735) );
  INV_X2 U11397 ( .I(n29441), .ZN(n29435) );
  NAND2_X2 U11398 ( .A1(n12261), .A2(n18494), .ZN(n29441) );
  AOI21_X1 U11435 ( .A1(n18518), .A2(n7537), .B(n33361), .ZN(n18516) );
  INV_X2 U11444 ( .I(n30946), .ZN(n875) );
  NOR2_X1 U11458 ( .A1(n1579), .A2(n19420), .ZN(n30948) );
  XOR2_X1 U11473 ( .A1(n28373), .A2(n28372), .Z(n30956) );
  XOR2_X1 U11520 ( .A1(n24013), .A2(n17725), .Z(n16109) );
  XOR2_X1 U11533 ( .A1(n23755), .A2(n18301), .Z(n23736) );
  OAI22_X2 U11535 ( .A1(n10612), .A2(n13560), .B1(n10614), .B2(n10613), .ZN(
        n18301) );
  NAND2_X2 U11550 ( .A1(n30962), .A2(n27925), .ZN(n5418) );
  XOR2_X1 U11555 ( .A1(n24068), .A2(n5842), .Z(n30963) );
  NAND2_X2 U11583 ( .A1(n30965), .A2(n28477), .ZN(n29093) );
  OAI21_X2 U11584 ( .A1(n9674), .A2(n31088), .B(n9673), .ZN(n30965) );
  OAI21_X2 U11594 ( .A1(n31452), .A2(n24283), .B(n24284), .ZN(n24120) );
  NOR2_X1 U11601 ( .A1(n38367), .A2(n32472), .ZN(n17867) );
  XOR2_X1 U11622 ( .A1(n23813), .A2(n34851), .Z(n30976) );
  AOI22_X2 U11630 ( .A1(n1673), .A2(n30306), .B1(n12077), .B2(n22126), .ZN(
        n32667) );
  XOR2_X1 U11631 ( .A1(n27731), .A2(n19943), .Z(n27079) );
  XOR2_X1 U11639 ( .A1(n30971), .A2(n30169), .Z(Ciphertext[174]) );
  AOI21_X2 U11647 ( .A1(n20947), .A2(n14855), .B(n20946), .ZN(n23762) );
  XOR2_X1 U11650 ( .A1(n30972), .A2(n27518), .Z(n7729) );
  XOR2_X1 U11651 ( .A1(n27640), .A2(n30973), .Z(n30972) );
  INV_X1 U11656 ( .I(n29718), .ZN(n30973) );
  NOR2_X2 U11657 ( .A1(n8385), .A2(n14261), .ZN(n10508) );
  XNOR2_X1 U11662 ( .A1(n5688), .A2(n34513), .ZN(n33486) );
  XOR2_X1 U11663 ( .A1(n26369), .A2(n26371), .Z(n19021) );
  NOR2_X1 U11672 ( .A1(n21445), .A2(n16496), .ZN(n21671) );
  OR2_X1 U11686 ( .A1(n7424), .A2(n14949), .Z(n27321) );
  NAND2_X1 U11699 ( .A1(n1382), .A2(n35175), .ZN(n2490) );
  OR2_X2 U11730 ( .A1(n17767), .A2(n7281), .Z(n6777) );
  INV_X2 U11748 ( .I(n30982), .ZN(n33949) );
  NOR2_X1 U11763 ( .A1(n23435), .A2(n34494), .ZN(n31798) );
  OR2_X1 U11785 ( .A1(n30986), .A2(n9369), .Z(n9415) );
  XOR2_X1 U11796 ( .A1(n30990), .A2(n8975), .Z(n13595) );
  XOR2_X1 U11798 ( .A1(n27727), .A2(n8974), .Z(n30990) );
  OAI21_X2 U11814 ( .A1(n10467), .A2(n10468), .B(n9683), .ZN(n31181) );
  XOR2_X1 U11819 ( .A1(n26530), .A2(n26559), .Z(n32386) );
  AND3_X1 U11827 ( .A1(n1755), .A2(n4083), .A3(n20405), .Z(n30197) );
  XOR2_X1 U11842 ( .A1(n34091), .A2(n8283), .Z(n30994) );
  NAND2_X2 U11845 ( .A1(n10261), .A2(n12892), .ZN(n22194) );
  NAND2_X2 U11854 ( .A1(n16024), .A2(n13743), .ZN(n25860) );
  OR2_X1 U11876 ( .A1(n7424), .A2(n31006), .Z(n20725) );
  XOR2_X1 U11887 ( .A1(n10860), .A2(n10858), .Z(n17169) );
  NAND2_X1 U11891 ( .A1(n31002), .A2(n31001), .ZN(n13621) );
  NOR2_X1 U11902 ( .A1(n20655), .A2(n24433), .ZN(n20654) );
  NOR2_X1 U11903 ( .A1(n24444), .A2(n24443), .ZN(n31003) );
  NAND2_X1 U11908 ( .A1(n20873), .A2(n22813), .ZN(n23075) );
  NOR2_X1 U11909 ( .A1(n12790), .A2(n17887), .ZN(n22967) );
  AOI22_X2 U11918 ( .A1(n31475), .A2(n33864), .B1(n3884), .B2(n8757), .ZN(
        n32506) );
  OR3_X1 U11953 ( .A1(n9790), .A2(n35272), .A3(n16260), .Z(n31997) );
  INV_X2 U11985 ( .I(n14949), .ZN(n31006) );
  NAND2_X2 U12011 ( .A1(n20663), .A2(n14232), .ZN(n11875) );
  AOI22_X2 U12020 ( .A1(n18645), .A2(n21469), .B1(n2628), .B2(n12314), .ZN(
        n2736) );
  OAI21_X2 U12031 ( .A1(n23571), .A2(n23577), .B(n12153), .ZN(n23540) );
  NAND2_X1 U12088 ( .A1(n33905), .A2(n33904), .ZN(n32057) );
  XOR2_X1 U12090 ( .A1(n19428), .A2(n31016), .Z(n32621) );
  XOR2_X1 U12104 ( .A1(n29303), .A2(n31017), .Z(n31016) );
  INV_X1 U12110 ( .I(n19534), .ZN(n31017) );
  AOI21_X2 U12123 ( .A1(n14103), .A2(n11875), .B(n11876), .ZN(n7428) );
  XOR2_X1 U12152 ( .A1(n15450), .A2(n21259), .Z(n13936) );
  XOR2_X1 U12159 ( .A1(n19072), .A2(n3589), .Z(n437) );
  XOR2_X1 U12166 ( .A1(n17486), .A2(n17487), .Z(n7371) );
  NAND3_X1 U12172 ( .A1(n4864), .A2(n4865), .A3(n1047), .ZN(n6032) );
  NAND2_X2 U12185 ( .A1(n28557), .A2(n28558), .ZN(n9930) );
  OAI21_X1 U12199 ( .A1(n24784), .A2(n37411), .B(n31023), .ZN(n15878) );
  XOR2_X1 U12222 ( .A1(n32646), .A2(n19800), .Z(n22532) );
  AND2_X1 U12253 ( .A1(n29361), .A2(n13804), .Z(n32767) );
  AOI22_X1 U12263 ( .A1(n21618), .A2(n3907), .B1(n38673), .B2(n38448), .ZN(
        n3909) );
  XOR2_X1 U12277 ( .A1(n31031), .A2(n33434), .Z(n20284) );
  XOR2_X1 U12329 ( .A1(n25077), .A2(n25078), .Z(n33044) );
  NAND2_X1 U12331 ( .A1(n21282), .A2(n21283), .ZN(n31726) );
  INV_X2 U12393 ( .I(n28025), .ZN(n27948) );
  OR2_X1 U12406 ( .A1(n19863), .A2(n19153), .Z(n12463) );
  XOR2_X1 U12439 ( .A1(n447), .A2(n31046), .Z(n3852) );
  XOR2_X1 U12451 ( .A1(n3855), .A2(n29029), .Z(n31046) );
  OR2_X1 U12454 ( .A1(n31278), .A2(n13144), .Z(n24114) );
  INV_X2 U12462 ( .I(n31507), .ZN(n21401) );
  NAND3_X2 U12464 ( .A1(n18341), .A2(n19038), .A3(n19039), .ZN(n28434) );
  XOR2_X1 U12470 ( .A1(n3645), .A2(n31047), .Z(n25669) );
  XOR2_X1 U12489 ( .A1(n25202), .A2(n30459), .Z(n31047) );
  XOR2_X1 U12494 ( .A1(n26155), .A2(n25947), .Z(n5965) );
  NOR2_X2 U12510 ( .A1(n30131), .A2(n18588), .ZN(n12350) );
  XOR2_X1 U12535 ( .A1(n8132), .A2(n14102), .Z(n14101) );
  NOR2_X2 U12559 ( .A1(n10420), .A2(n37056), .ZN(n28418) );
  AOI21_X1 U12563 ( .A1(n28546), .A2(n3944), .B(n36623), .ZN(n31699) );
  XNOR2_X1 U12596 ( .A1(n15671), .A2(n11253), .ZN(n31352) );
  NAND3_X1 U12624 ( .A1(n29763), .A2(n29764), .A3(n19599), .ZN(n31059) );
  INV_X4 U12630 ( .I(n2242), .ZN(n9105) );
  AOI21_X2 U12633 ( .A1(n6332), .A2(n19147), .B(n2243), .ZN(n2242) );
  NAND3_X1 U12638 ( .A1(n15737), .A2(n35224), .A3(n15224), .ZN(n28466) );
  XOR2_X1 U12643 ( .A1(n269), .A2(n31062), .Z(n31061) );
  INV_X1 U12645 ( .I(n19843), .ZN(n31062) );
  XOR2_X1 U12682 ( .A1(n24959), .A2(n30682), .Z(n1819) );
  XOR2_X1 U12696 ( .A1(n31070), .A2(n31585), .Z(n27473) );
  NOR2_X1 U12710 ( .A1(n32318), .A2(n17685), .ZN(n22253) );
  NAND2_X1 U12730 ( .A1(n4889), .A2(n5938), .ZN(n3193) );
  AOI21_X2 U12742 ( .A1(n11056), .A2(n29422), .B(n907), .ZN(n29354) );
  NAND2_X2 U12747 ( .A1(n18550), .A2(n18552), .ZN(n18148) );
  XOR2_X1 U12752 ( .A1(n8110), .A2(n11935), .Z(n26225) );
  NOR2_X1 U12754 ( .A1(n21747), .A2(n38546), .ZN(n32808) );
  NAND3_X1 U12775 ( .A1(n29384), .A2(n10422), .A3(n11084), .ZN(n6262) );
  XOR2_X1 U12786 ( .A1(n11074), .A2(n11076), .Z(n13417) );
  AOI21_X2 U12819 ( .A1(n23331), .A2(n32226), .B(n20118), .ZN(n24070) );
  AOI21_X2 U12821 ( .A1(n20438), .A2(n4601), .B(n5245), .ZN(n25247) );
  INV_X2 U12825 ( .I(n31078), .ZN(n12064) );
  OAI21_X2 U12832 ( .A1(n16224), .A2(n29935), .B(n8593), .ZN(n8592) );
  INV_X2 U12833 ( .I(n18910), .ZN(n18972) );
  NAND2_X2 U12864 ( .A1(n31082), .A2(n25628), .ZN(n11033) );
  NAND2_X2 U12881 ( .A1(n35618), .A2(n8275), .ZN(n5527) );
  NOR2_X2 U12892 ( .A1(n3685), .A2(n38886), .ZN(n12665) );
  XOR2_X1 U12910 ( .A1(n31086), .A2(n29934), .Z(Ciphertext[131]) );
  AOI22_X1 U12930 ( .A1(n29931), .A2(n9591), .B1(n29933), .B2(n29932), .ZN(
        n31086) );
  NAND2_X2 U12944 ( .A1(n24243), .A2(n17591), .ZN(n7520) );
  OAI22_X2 U12964 ( .A1(n13762), .A2(n34064), .B1(n29287), .B2(n29348), .ZN(
        n12371) );
  XOR2_X1 U12972 ( .A1(n31089), .A2(n7382), .Z(n10816) );
  NAND2_X2 U13005 ( .A1(n14017), .A2(n31090), .ZN(n23619) );
  OR2_X1 U13009 ( .A1(n23186), .A2(n11197), .Z(n31090) );
  NAND2_X1 U13011 ( .A1(n20835), .A2(n23390), .ZN(n31091) );
  BUF_X2 U13013 ( .I(n14349), .Z(n31092) );
  XOR2_X1 U13017 ( .A1(n7358), .A2(n22614), .Z(n4279) );
  NAND2_X2 U13037 ( .A1(n31094), .A2(n16543), .ZN(n33707) );
  AOI21_X2 U13042 ( .A1(n28699), .A2(n16494), .B(n13718), .ZN(n126) );
  NAND2_X2 U13059 ( .A1(n2725), .A2(n32918), .ZN(n20276) );
  XOR2_X1 U13064 ( .A1(n22748), .A2(n7200), .Z(n7199) );
  XOR2_X1 U13079 ( .A1(n13871), .A2(n14104), .Z(n24369) );
  XOR2_X1 U13086 ( .A1(n2135), .A2(n2136), .Z(n2134) );
  NAND2_X2 U13131 ( .A1(n22043), .A2(n22044), .ZN(n22634) );
  NOR2_X2 U13134 ( .A1(n9667), .A2(n26008), .ZN(n33892) );
  NOR2_X2 U13151 ( .A1(n32183), .A2(n31102), .ZN(n33286) );
  AND2_X2 U13156 ( .A1(n32838), .A2(n16832), .Z(n13884) );
  XOR2_X1 U13157 ( .A1(n3240), .A2(n31103), .Z(n11643) );
  XOR2_X1 U13158 ( .A1(n22530), .A2(n18969), .Z(n31103) );
  XOR2_X1 U13163 ( .A1(n31628), .A2(n25271), .Z(n21154) );
  INV_X4 U13172 ( .I(n12064), .ZN(n15049) );
  XOR2_X1 U13189 ( .A1(n6388), .A2(n31108), .Z(n10810) );
  XOR2_X1 U13196 ( .A1(n20695), .A2(n6387), .Z(n31108) );
  OR2_X1 U13220 ( .A1(n27009), .A2(n12156), .Z(n31110) );
  NAND2_X2 U13224 ( .A1(n4988), .A2(n4989), .ZN(n33293) );
  NAND2_X2 U13225 ( .A1(n31115), .A2(n31114), .ZN(n18987) );
  XOR2_X1 U13236 ( .A1(n25226), .A2(n14385), .Z(n25289) );
  OR2_X1 U13245 ( .A1(n12408), .A2(n16547), .Z(n32430) );
  INV_X2 U13247 ( .I(n31121), .ZN(n28152) );
  NOR3_X2 U13255 ( .A1(n4578), .A2(n31123), .A3(n31122), .ZN(n24961) );
  NAND2_X2 U13259 ( .A1(n31124), .A2(n33042), .ZN(n3214) );
  AOI22_X1 U13265 ( .A1(n29665), .A2(n30295), .B1(n29648), .B2(n29654), .ZN(
        n32288) );
  INV_X2 U13279 ( .I(n9113), .ZN(n9114) );
  XOR2_X1 U13302 ( .A1(n31129), .A2(n33466), .Z(n12315) );
  XOR2_X1 U13306 ( .A1(n19118), .A2(n22602), .Z(n31129) );
  XOR2_X1 U13309 ( .A1(n20668), .A2(n22532), .Z(n11750) );
  XOR2_X1 U13319 ( .A1(n9121), .A2(n9123), .Z(n9458) );
  XOR2_X1 U13335 ( .A1(n15164), .A2(n27719), .Z(n17138) );
  NAND2_X2 U13378 ( .A1(n24120), .A2(n32891), .ZN(n23766) );
  XOR2_X1 U13382 ( .A1(n26420), .A2(n3710), .Z(n33751) );
  XOR2_X1 U13406 ( .A1(n31138), .A2(n27229), .Z(n342) );
  XOR2_X1 U13410 ( .A1(n24994), .A2(n31139), .Z(n14350) );
  INV_X2 U13415 ( .I(n36992), .ZN(n4880) );
  INV_X4 U13430 ( .I(n23523), .ZN(n23522) );
  XOR2_X1 U13432 ( .A1(n4305), .A2(n1819), .Z(n33188) );
  XOR2_X1 U13435 ( .A1(n31149), .A2(n1361), .Z(Ciphertext[83]) );
  AOI22_X1 U13445 ( .A1(n29665), .A2(n29664), .B1(n29663), .B2(n1390), .ZN(
        n31149) );
  NAND2_X2 U13454 ( .A1(n992), .A2(n32557), .ZN(n31150) );
  NAND2_X2 U13458 ( .A1(n13228), .A2(n13227), .ZN(n24250) );
  XOR2_X1 U13491 ( .A1(n16587), .A2(n31152), .Z(n6834) );
  XOR2_X1 U13493 ( .A1(n29071), .A2(n19814), .Z(n31152) );
  XOR2_X1 U13500 ( .A1(n2864), .A2(n39172), .Z(n31154) );
  NAND2_X1 U13562 ( .A1(n35828), .A2(n9743), .ZN(n5681) );
  XOR2_X1 U13578 ( .A1(n21197), .A2(n22614), .Z(n5703) );
  XOR2_X1 U13581 ( .A1(n22711), .A2(n22475), .Z(n22614) );
  XOR2_X1 U13646 ( .A1(n29111), .A2(n13933), .Z(n31162) );
  XOR2_X1 U13704 ( .A1(n27714), .A2(n7345), .Z(n4783) );
  XOR2_X1 U13790 ( .A1(n35529), .A2(n31173), .Z(n20006) );
  NAND2_X2 U13803 ( .A1(n18281), .A2(n7905), .ZN(n28516) );
  AND2_X1 U13810 ( .A1(n39504), .A2(n8735), .Z(n31177) );
  XOR2_X1 U13819 ( .A1(n9122), .A2(n31178), .Z(n8300) );
  OR2_X1 U13828 ( .A1(n15854), .A2(n10959), .Z(n29892) );
  XOR2_X1 U13836 ( .A1(n2161), .A2(n2162), .Z(n29865) );
  XOR2_X1 U13841 ( .A1(n12850), .A2(n33165), .Z(n11562) );
  NAND2_X2 U13876 ( .A1(n1102), .A2(n25966), .ZN(n19340) );
  OAI22_X2 U13902 ( .A1(n20287), .A2(n29634), .B1(n20286), .B2(n20289), .ZN(
        n29660) );
  XOR2_X1 U13982 ( .A1(n31191), .A2(n27695), .Z(n27696) );
  XOR2_X1 U13983 ( .A1(n13569), .A2(n34963), .Z(n31191) );
  NAND2_X1 U14073 ( .A1(n16778), .A2(n9405), .ZN(n9404) );
  NAND2_X1 U14076 ( .A1(n16778), .A2(n13880), .ZN(n31194) );
  INV_X2 U14094 ( .I(n31196), .ZN(n2799) );
  XOR2_X1 U14096 ( .A1(n2800), .A2(n4129), .Z(n31196) );
  XOR2_X1 U14102 ( .A1(n31197), .A2(n33661), .Z(Ciphertext[67]) );
  XOR2_X1 U14104 ( .A1(n27777), .A2(n27707), .Z(n27204) );
  NOR3_X1 U14124 ( .A1(n30859), .A2(n37104), .A3(n33561), .ZN(n5481) );
  INV_X2 U14139 ( .I(n31204), .ZN(n27790) );
  XOR2_X1 U14141 ( .A1(n22447), .A2(n700), .Z(n7932) );
  INV_X2 U14149 ( .I(n31207), .ZN(n10383) );
  NAND2_X2 U14156 ( .A1(n31132), .A2(n24416), .ZN(n17496) );
  AOI21_X1 U14173 ( .A1(n31212), .A2(n31211), .B(n29338), .ZN(n3285) );
  NAND2_X1 U14174 ( .A1(n29339), .A2(n29336), .ZN(n31212) );
  INV_X4 U14175 ( .I(n10383), .ZN(n33745) );
  XOR2_X1 U14196 ( .A1(n11374), .A2(n746), .Z(n31215) );
  NAND2_X2 U14211 ( .A1(n32813), .A2(n2363), .ZN(n27408) );
  OAI21_X1 U14217 ( .A1(n19972), .A2(n1234), .B(n31220), .ZN(n2364) );
  XOR2_X1 U14246 ( .A1(n6470), .A2(n31230), .Z(n9516) );
  XOR2_X1 U14247 ( .A1(n27555), .A2(n18709), .Z(n31230) );
  OR2_X1 U14248 ( .A1(n29810), .A2(n13192), .Z(n31231) );
  XOR2_X1 U14265 ( .A1(n8908), .A2(n38225), .Z(n31233) );
  AOI22_X2 U14273 ( .A1(n13259), .A2(n13019), .B1(n25204), .B2(n24944), .ZN(
        n25299) );
  NAND2_X2 U14278 ( .A1(n31236), .A2(n5299), .ZN(n30178) );
  AND2_X1 U14305 ( .A1(n39814), .A2(n17509), .Z(n2975) );
  INV_X1 U14318 ( .I(n23768), .ZN(n31245) );
  NOR2_X1 U14319 ( .A1(n31245), .A2(n5897), .ZN(n31360) );
  XOR2_X1 U14320 ( .A1(n15930), .A2(n25275), .Z(n25007) );
  NOR2_X1 U14330 ( .A1(n24283), .A2(n24284), .ZN(n20732) );
  BUF_X2 U14338 ( .I(n23775), .Z(n31247) );
  XOR2_X1 U14344 ( .A1(n37812), .A2(n31249), .Z(n31248) );
  XOR2_X1 U14347 ( .A1(n17245), .A2(n31689), .Z(n31688) );
  INV_X2 U14353 ( .I(n31250), .ZN(n733) );
  XOR2_X1 U14354 ( .A1(n3579), .A2(n3577), .Z(n31250) );
  AND2_X1 U14357 ( .A1(n32146), .A2(n28620), .Z(n13404) );
  AOI21_X2 U14361 ( .A1(n25433), .A2(n36086), .B(n18565), .ZN(n26106) );
  AOI22_X2 U14367 ( .A1(n31252), .A2(n14371), .B1(n4128), .B2(n32899), .ZN(
        n20728) );
  INV_X2 U14369 ( .I(n14422), .ZN(n1055) );
  NAND2_X1 U14383 ( .A1(n31258), .A2(n19098), .ZN(n10031) );
  NAND2_X2 U14391 ( .A1(n33317), .A2(n20158), .ZN(n24713) );
  AND2_X1 U14406 ( .A1(n21671), .A2(n21672), .Z(n6046) );
  AND2_X1 U14407 ( .A1(n38886), .A2(n17509), .Z(n2971) );
  NAND2_X1 U14422 ( .A1(n10590), .A2(n16786), .ZN(n30228) );
  NOR2_X1 U14425 ( .A1(n15794), .A2(n10383), .ZN(n11197) );
  NAND2_X2 U14443 ( .A1(n31447), .A2(n10186), .ZN(n27275) );
  NAND2_X2 U14444 ( .A1(n30193), .A2(n35870), .ZN(n15267) );
  XOR2_X1 U14447 ( .A1(n12903), .A2(n1902), .Z(n12850) );
  OAI21_X1 U14468 ( .A1(n14968), .A2(n31269), .B(n31268), .ZN(n7478) );
  NAND2_X1 U14470 ( .A1(n14968), .A2(n1186), .ZN(n31268) );
  INV_X2 U14472 ( .I(n14987), .ZN(n31269) );
  XOR2_X1 U14479 ( .A1(n26521), .A2(n9301), .Z(n9300) );
  INV_X2 U14485 ( .I(n20864), .ZN(n31270) );
  INV_X2 U14504 ( .I(n31272), .ZN(n31494) );
  NAND2_X2 U14511 ( .A1(n31274), .A2(n16220), .ZN(n27292) );
  BUF_X2 U14520 ( .I(n37661), .Z(n31275) );
  NAND2_X2 U14560 ( .A1(n2955), .A2(n13466), .ZN(n17008) );
  XNOR2_X1 U14561 ( .A1(n28997), .A2(n38222), .ZN(n29139) );
  INV_X2 U14565 ( .I(n31278), .ZN(n14704) );
  XOR2_X1 U14567 ( .A1(n25296), .A2(n30761), .Z(n24976) );
  XOR2_X1 U14582 ( .A1(n2959), .A2(n24920), .Z(n15195) );
  XOR2_X1 U14583 ( .A1(n31281), .A2(n24977), .Z(n20514) );
  OR2_X1 U14601 ( .A1(n28114), .A2(n13457), .Z(n32485) );
  AOI21_X2 U14603 ( .A1(n3527), .A2(n19476), .B(n6044), .ZN(n9828) );
  OR2_X1 U14619 ( .A1(n19085), .A2(n5530), .Z(n11398) );
  NOR2_X2 U14639 ( .A1(n26001), .A2(n5753), .ZN(n25897) );
  XOR2_X1 U14658 ( .A1(n25159), .A2(n30405), .Z(n31289) );
  NAND2_X2 U14661 ( .A1(n16883), .A2(n16031), .ZN(n23808) );
  INV_X2 U14673 ( .I(n31294), .ZN(n17509) );
  NOR2_X1 U14680 ( .A1(n8165), .A2(n993), .ZN(n31806) );
  XOR2_X1 U14681 ( .A1(n33041), .A2(n31295), .Z(n32306) );
  INV_X1 U14683 ( .I(n29051), .ZN(n31295) );
  INV_X2 U14688 ( .I(n32536), .ZN(n13744) );
  AND2_X1 U14693 ( .A1(n19233), .A2(n17509), .Z(n4053) );
  XOR2_X1 U14695 ( .A1(n35350), .A2(n1215), .Z(n7345) );
  XOR2_X1 U14709 ( .A1(n25146), .A2(n24928), .Z(n25172) );
  NAND2_X2 U14722 ( .A1(n6019), .A2(n30052), .ZN(n30054) );
  XOR2_X1 U14729 ( .A1(n129), .A2(n11661), .Z(n11663) );
  NAND2_X2 U14747 ( .A1(n21445), .A2(n21845), .ZN(n14868) );
  NAND2_X2 U14751 ( .A1(n2765), .A2(n21864), .ZN(n13055) );
  NOR2_X1 U14755 ( .A1(n14635), .A2(n19955), .ZN(n18234) );
  XOR2_X1 U14756 ( .A1(n9154), .A2(n38291), .Z(n599) );
  AND2_X1 U14774 ( .A1(n23516), .A2(n23518), .Z(n18388) );
  AND2_X2 U14775 ( .A1(n24285), .A2(n24287), .Z(n9922) );
  XOR2_X1 U14786 ( .A1(n26357), .A2(n38219), .Z(n16082) );
  NAND2_X2 U14804 ( .A1(n5474), .A2(n25787), .ZN(n26520) );
  NAND2_X2 U14813 ( .A1(n9125), .A2(n9124), .ZN(n22492) );
  XOR2_X1 U14834 ( .A1(n1463), .A2(n19860), .Z(n31314) );
  NAND2_X1 U14856 ( .A1(n26093), .A2(n33258), .ZN(n31318) );
  NAND2_X2 U14867 ( .A1(n20236), .A2(n20237), .ZN(n33644) );
  OR2_X1 U14873 ( .A1(n1676), .A2(n36214), .Z(n33679) );
  XOR2_X1 U14878 ( .A1(n19103), .A2(n19100), .Z(n24463) );
  NAND2_X2 U14879 ( .A1(n7323), .A2(n31322), .ZN(n25867) );
  NOR2_X1 U14880 ( .A1(n7528), .A2(n12673), .ZN(n12785) );
  NOR2_X2 U14892 ( .A1(n36752), .A2(n37105), .ZN(n5653) );
  INV_X4 U14906 ( .I(n2765), .ZN(n12080) );
  XOR2_X1 U14912 ( .A1(n10129), .A2(n31327), .Z(n10132) );
  XOR2_X1 U14917 ( .A1(n27819), .A2(n1938), .Z(n31327) );
  NAND2_X2 U14924 ( .A1(n4329), .A2(n11912), .ZN(n33316) );
  INV_X2 U14925 ( .I(n31329), .ZN(n5112) );
  NOR2_X2 U14947 ( .A1(n31871), .A2(n6713), .ZN(n11413) );
  INV_X2 U14948 ( .I(n29591), .ZN(n29597) );
  AOI21_X1 U14954 ( .A1(n20041), .A2(n20517), .B(n11449), .ZN(n33264) );
  XOR2_X1 U14966 ( .A1(n17879), .A2(n31334), .Z(n17878) );
  XOR2_X1 U14968 ( .A1(n24927), .A2(n33311), .Z(n31334) );
  INV_X2 U14975 ( .I(n31335), .ZN(n2532) );
  XOR2_X1 U14976 ( .A1(Plaintext[104]), .A2(Key[104]), .Z(n31335) );
  NAND2_X2 U14985 ( .A1(n12130), .A2(n31343), .ZN(n2553) );
  AND2_X1 U14991 ( .A1(n775), .A2(n20616), .Z(n14127) );
  INV_X2 U14992 ( .I(n31341), .ZN(n10314) );
  XOR2_X1 U14993 ( .A1(n10316), .A2(n10315), .Z(n31341) );
  AND2_X1 U15008 ( .A1(n26031), .A2(n35903), .Z(n5981) );
  OR2_X2 U15028 ( .A1(n20171), .A2(n14000), .Z(n26674) );
  XOR2_X1 U15029 ( .A1(n17957), .A2(n29248), .Z(n13800) );
  NOR2_X1 U15050 ( .A1(n7445), .A2(n35981), .ZN(n31346) );
  AOI22_X2 U15069 ( .A1(n24374), .A2(n31349), .B1(n13070), .B2(n24430), .ZN(
        n24864) );
  NAND2_X1 U15074 ( .A1(n38609), .A2(n16081), .ZN(n31349) );
  NAND2_X2 U15084 ( .A1(n14553), .A2(n138), .ZN(n31984) );
  NAND2_X1 U15087 ( .A1(n31350), .A2(n1192), .ZN(n20487) );
  NAND2_X1 U15115 ( .A1(n9821), .A2(n9822), .ZN(n14169) );
  XOR2_X1 U15123 ( .A1(n11899), .A2(n25293), .Z(n9007) );
  XOR2_X1 U15127 ( .A1(n20333), .A2(n13342), .Z(n25293) );
  OAI21_X2 U15146 ( .A1(n6491), .A2(n24710), .B(n13046), .ZN(n24701) );
  OR2_X1 U15150 ( .A1(n14404), .A2(n28123), .Z(n27107) );
  XOR2_X1 U15154 ( .A1(n7137), .A2(n22587), .Z(n22605) );
  INV_X2 U15157 ( .I(n20541), .ZN(n19050) );
  NOR2_X1 U15168 ( .A1(n23958), .A2(n24469), .ZN(n17789) );
  NAND2_X2 U15185 ( .A1(n11065), .A2(n11064), .ZN(n17400) );
  NOR2_X2 U15186 ( .A1(n11066), .A2(n10719), .ZN(n11065) );
  NAND3_X2 U15199 ( .A1(n31735), .A2(n27135), .A3(n31734), .ZN(n12551) );
  XOR2_X1 U15206 ( .A1(n19536), .A2(n23939), .Z(n23972) );
  INV_X1 U15222 ( .I(n30095), .ZN(n30086) );
  AND2_X1 U15223 ( .A1(n15085), .A2(n5753), .Z(n10179) );
  NAND2_X2 U15240 ( .A1(n31365), .A2(n7551), .ZN(n10632) );
  XOR2_X1 U15242 ( .A1(n31366), .A2(n38962), .Z(Ciphertext[77]) );
  NOR2_X2 U15252 ( .A1(n31369), .A2(n9904), .ZN(n12661) );
  XOR2_X1 U15296 ( .A1(n31377), .A2(n893), .Z(n32251) );
  XOR2_X1 U15299 ( .A1(n29242), .A2(n12707), .Z(n12939) );
  AND2_X1 U15303 ( .A1(n28559), .A2(n31353), .Z(n7615) );
  NOR2_X1 U15305 ( .A1(n31378), .A2(n28402), .ZN(n9355) );
  AOI21_X1 U15307 ( .A1(n36827), .A2(n10544), .B(n37804), .ZN(n11680) );
  OAI22_X1 U15308 ( .A1(n24162), .A2(n914), .B1(n124), .B2(n10152), .ZN(n2674)
         );
  OR2_X1 U15309 ( .A1(n28152), .A2(n28153), .Z(n9168) );
  XOR2_X1 U15322 ( .A1(Plaintext[16]), .A2(Key[16]), .Z(n31381) );
  AND2_X1 U15323 ( .A1(n25460), .A2(n31809), .Z(n25008) );
  XOR2_X1 U15336 ( .A1(n16062), .A2(n8482), .Z(n32165) );
  OAI22_X2 U15337 ( .A1(n15706), .A2(n6670), .B1(n6671), .B2(n6672), .ZN(
        n33678) );
  XOR2_X1 U15345 ( .A1(n27579), .A2(n3891), .Z(n3887) );
  XOR2_X1 U15353 ( .A1(n3953), .A2(n39804), .Z(n17910) );
  OAI21_X1 U15359 ( .A1(n37748), .A2(n39226), .B(n38300), .ZN(n31386) );
  INV_X4 U15401 ( .I(n5112), .ZN(n14472) );
  AND2_X1 U15411 ( .A1(n25820), .A2(n17791), .Z(n11633) );
  NOR3_X1 U15414 ( .A1(n39083), .A2(n31549), .A3(n30213), .ZN(n7792) );
  NAND2_X2 U15419 ( .A1(n12617), .A2(n1630), .ZN(n23397) );
  OAI21_X2 U15427 ( .A1(n31400), .A2(n31399), .B(n27391), .ZN(n18171) );
  XOR2_X1 U15436 ( .A1(n507), .A2(n25298), .Z(n13919) );
  XOR2_X1 U15443 ( .A1(n10385), .A2(n34126), .Z(n31401) );
  XOR2_X1 U15453 ( .A1(n6641), .A2(n27696), .Z(n20531) );
  NAND2_X2 U15459 ( .A1(n18289), .A2(n7660), .ZN(n25991) );
  AND2_X1 U15463 ( .A1(n22320), .A2(n22319), .Z(n33594) );
  NOR2_X1 U15470 ( .A1(n23173), .A2(n34757), .ZN(n22939) );
  NAND2_X2 U15494 ( .A1(n1454), .A2(n18689), .ZN(n4809) );
  XOR2_X1 U15520 ( .A1(n33083), .A2(n26158), .Z(n31414) );
  NAND2_X2 U15526 ( .A1(n32091), .A2(n24753), .ZN(n5888) );
  OAI21_X2 U15543 ( .A1(n18456), .A2(n18455), .B(n18454), .ZN(n24694) );
  INV_X2 U15544 ( .I(n20512), .ZN(n28023) );
  XOR2_X1 U15547 ( .A1(n20511), .A2(n14641), .Z(n20512) );
  NAND2_X1 U15548 ( .A1(n33291), .A2(n8745), .ZN(n3107) );
  NAND2_X1 U15553 ( .A1(n38762), .A2(n4649), .ZN(n13769) );
  XOR2_X1 U15578 ( .A1(n12244), .A2(n29144), .Z(n29037) );
  NAND3_X2 U15584 ( .A1(n28359), .A2(n28357), .A3(n28358), .ZN(n12244) );
  NOR2_X1 U15595 ( .A1(n5926), .A2(n5927), .ZN(n31424) );
  INV_X2 U15596 ( .I(n31426), .ZN(n28231) );
  NAND2_X1 U15605 ( .A1(n30311), .A2(n3869), .ZN(n7773) );
  XOR2_X1 U15609 ( .A1(n31427), .A2(n28412), .Z(n28414) );
  XOR2_X1 U15610 ( .A1(n28406), .A2(n28959), .Z(n31427) );
  OAI22_X2 U15611 ( .A1(n39706), .A2(n10477), .B1(n1609), .B2(n15751), .ZN(
        n24353) );
  XNOR2_X1 U15612 ( .A1(n1659), .A2(n15513), .ZN(n32331) );
  AOI22_X2 U15620 ( .A1(n21336), .A2(n21599), .B1(n20535), .B2(n17992), .ZN(
        n17991) );
  NOR2_X2 U15643 ( .A1(n29909), .A2(n29910), .ZN(n29929) );
  OAI21_X2 U15645 ( .A1(n17145), .A2(n18656), .B(n31407), .ZN(n17154) );
  AOI22_X1 U15660 ( .A1(n30119), .A2(n16275), .B1(n16277), .B2(n30107), .ZN(
        n31430) );
  XOR2_X1 U15668 ( .A1(n11791), .A2(n33622), .Z(n17021) );
  NAND3_X1 U15669 ( .A1(n4986), .A2(n24393), .A3(n15018), .ZN(n16450) );
  NAND2_X2 U15676 ( .A1(n32404), .A2(n18050), .ZN(n27773) );
  AOI21_X2 U15687 ( .A1(n23441), .A2(n1290), .B(n17960), .ZN(n23442) );
  NAND2_X2 U15726 ( .A1(n16932), .A2(n11026), .ZN(n29144) );
  XOR2_X1 U15738 ( .A1(n25039), .A2(n25318), .Z(n4501) );
  AOI21_X2 U15762 ( .A1(n5490), .A2(n1302), .B(n31441), .ZN(n5488) );
  NOR2_X2 U15763 ( .A1(n18989), .A2(n23468), .ZN(n31441) );
  OAI21_X1 U15768 ( .A1(n31912), .A2(n31911), .B(n968), .ZN(n2569) );
  XOR2_X1 U15770 ( .A1(n31442), .A2(n870), .Z(n15774) );
  INV_X1 U15772 ( .I(n29903), .ZN(n31444) );
  OR2_X1 U15779 ( .A1(n35207), .A2(n18827), .Z(n16071) );
  NAND2_X2 U15780 ( .A1(n1295), .A2(n33840), .ZN(n11453) );
  XOR2_X1 U15816 ( .A1(n27722), .A2(n27753), .Z(n19231) );
  NAND2_X2 U15837 ( .A1(n1597), .A2(n37377), .ZN(n6298) );
  XOR2_X1 U15843 ( .A1(n29094), .A2(n29164), .Z(n6537) );
  XOR2_X1 U15844 ( .A1(n29058), .A2(n17880), .Z(n29164) );
  NAND2_X2 U15861 ( .A1(n14027), .A2(n1338), .ZN(n2841) );
  NOR2_X2 U15885 ( .A1(n19700), .A2(n26879), .ZN(n26994) );
  NOR2_X2 U15905 ( .A1(n32575), .A2(n38629), .ZN(n28683) );
  NOR2_X1 U15910 ( .A1(n24146), .A2(n1123), .ZN(n31464) );
  INV_X2 U15912 ( .I(n1230), .ZN(n20399) );
  XOR2_X1 U15936 ( .A1(n24079), .A2(n20340), .Z(n31466) );
  XOR2_X1 U15937 ( .A1(n14309), .A2(n31576), .Z(n2988) );
  NAND2_X2 U15951 ( .A1(n1418), .A2(n28695), .ZN(n28598) );
  OR2_X1 U15973 ( .A1(n33786), .A2(n20276), .Z(n23054) );
  NAND3_X2 U16028 ( .A1(n3746), .A2(n23385), .A3(n3743), .ZN(n9518) );
  NAND3_X1 U16037 ( .A1(n33608), .A2(n33607), .A3(n29732), .ZN(n31477) );
  NAND2_X2 U16067 ( .A1(n3681), .A2(n3682), .ZN(n22064) );
  NOR2_X1 U16070 ( .A1(n3452), .A2(n31019), .ZN(n19660) );
  NAND2_X2 U16076 ( .A1(n31484), .A2(n20250), .ZN(n19828) );
  NAND2_X2 U16082 ( .A1(n6089), .A2(n6088), .ZN(n9395) );
  XOR2_X1 U16084 ( .A1(n5241), .A2(n19833), .Z(n1880) );
  INV_X2 U16086 ( .I(n22350), .ZN(n21288) );
  NAND2_X1 U16093 ( .A1(n22350), .A2(n30315), .ZN(n16267) );
  NAND2_X2 U16094 ( .A1(n21716), .A2(n21717), .ZN(n22350) );
  XOR2_X1 U16095 ( .A1(n22570), .A2(n29657), .Z(n644) );
  NAND2_X2 U16130 ( .A1(n3513), .A2(n4034), .ZN(n27299) );
  NAND3_X2 U16142 ( .A1(n34117), .A2(n25790), .A3(n1019), .ZN(n18463) );
  INV_X1 U16144 ( .I(n33267), .ZN(n33266) );
  XOR2_X1 U16165 ( .A1(n19221), .A2(n29285), .Z(n31492) );
  AOI21_X2 U16176 ( .A1(n34064), .A2(n13349), .B(n29348), .ZN(n13000) );
  AND2_X1 U16183 ( .A1(n9775), .A2(n9791), .Z(n28101) );
  XOR2_X1 U16201 ( .A1(n31500), .A2(n29130), .Z(n13052) );
  XOR2_X1 U16202 ( .A1(n29124), .A2(n35255), .Z(n31500) );
  NAND3_X2 U16208 ( .A1(n15881), .A2(n15882), .A3(n37238), .ZN(n25778) );
  AOI21_X2 U16226 ( .A1(n3912), .A2(n2690), .B(n30427), .ZN(n32) );
  XOR2_X1 U16240 ( .A1(n31505), .A2(n30452), .Z(n32310) );
  OAI21_X2 U16272 ( .A1(n16252), .A2(n29421), .B(n13153), .ZN(n1820) );
  NAND2_X2 U16276 ( .A1(n9914), .A2(n6002), .ZN(n29218) );
  NAND2_X2 U16294 ( .A1(n38143), .A2(n29756), .ZN(n29737) );
  BUF_X2 U16305 ( .I(n28848), .Z(n31516) );
  CLKBUF_X4 U16318 ( .I(n12410), .Z(n11658) );
  INV_X1 U16323 ( .I(n32477), .ZN(n24270) );
  OAI21_X1 U16344 ( .A1(n14093), .A2(n4640), .B(n19435), .ZN(n13726) );
  AOI22_X1 U16347 ( .A1(n28773), .A2(n5662), .B1(n32286), .B2(n9353), .ZN(
        n20430) );
  XOR2_X1 U16361 ( .A1(Plaintext[185]), .A2(Key[185]), .Z(n31507) );
  XOR2_X1 U16363 ( .A1(n22754), .A2(n31508), .Z(n31559) );
  XOR2_X1 U16367 ( .A1(n22570), .A2(n29221), .Z(n31508) );
  XNOR2_X1 U16368 ( .A1(n5816), .A2(n5815), .ZN(n31509) );
  INV_X1 U16374 ( .I(n8475), .ZN(n1409) );
  OR2_X1 U16379 ( .A1(n33368), .A2(n31511), .Z(n19111) );
  AND2_X1 U16385 ( .A1(n17983), .A2(n29961), .Z(n31512) );
  OAI21_X1 U16386 ( .A1(n32480), .A2(n32479), .B(n19750), .ZN(n5665) );
  NAND2_X1 U16416 ( .A1(n2823), .A2(n14209), .ZN(n2774) );
  NAND2_X1 U16420 ( .A1(n252), .A2(n6657), .ZN(n6656) );
  INV_X2 U16422 ( .I(n15853), .ZN(n16510) );
  NAND2_X1 U16426 ( .A1(n16510), .A2(n21285), .ZN(n10147) );
  NOR2_X1 U16450 ( .A1(n20491), .A2(n20490), .ZN(n26349) );
  AOI21_X1 U16459 ( .A1(n13004), .A2(n10355), .B(n37955), .ZN(n32388) );
  NAND2_X2 U16467 ( .A1(n31516), .A2(n29760), .ZN(n31517) );
  NAND2_X1 U16493 ( .A1(n2364), .A2(n735), .ZN(n2363) );
  NAND3_X1 U16509 ( .A1(n29416), .A2(n29408), .A3(n29409), .ZN(n15042) );
  NOR2_X1 U16535 ( .A1(n27404), .A2(n27390), .ZN(n33888) );
  AOI22_X1 U16539 ( .A1(n10293), .A2(n31968), .B1(n10292), .B2(n29888), .ZN(
        n32470) );
  NAND2_X1 U16556 ( .A1(n3538), .A2(n28330), .ZN(n17522) );
  AND2_X2 U16557 ( .A1(n16700), .A2(n31638), .Z(n31518) );
  NAND3_X1 U16579 ( .A1(n29997), .A2(n30042), .A3(n16328), .ZN(n19196) );
  NOR2_X1 U16583 ( .A1(n7583), .A2(n33346), .ZN(n31660) );
  NOR2_X1 U16610 ( .A1(n35023), .A2(n28366), .ZN(n32315) );
  NAND2_X1 U16616 ( .A1(n30129), .A2(n17192), .ZN(n31693) );
  INV_X1 U16623 ( .I(n33324), .ZN(n938) );
  AND2_X1 U16631 ( .A1(n16542), .A2(n9528), .Z(n31520) );
  NAND2_X1 U16640 ( .A1(n9534), .A2(n12302), .ZN(n10351) );
  INV_X2 U16665 ( .I(n13054), .ZN(n27557) );
  AND2_X1 U16666 ( .A1(n30260), .A2(n30259), .Z(n14512) );
  NAND2_X1 U16670 ( .A1(n8659), .A2(n14237), .ZN(n31522) );
  BUF_X2 U16675 ( .I(n20207), .Z(n7949) );
  INV_X2 U16679 ( .I(n28578), .ZN(n3598) );
  NAND3_X1 U16684 ( .A1(n26972), .A2(n15980), .A3(n26973), .ZN(n15979) );
  NAND3_X1 U16686 ( .A1(n26974), .A2(n26972), .A3(n32427), .ZN(n16573) );
  NAND2_X1 U16705 ( .A1(n29338), .A2(n38151), .ZN(n3288) );
  NOR2_X1 U16712 ( .A1(n1173), .A2(n18042), .ZN(n29670) );
  OAI21_X1 U16727 ( .A1(n1178), .A2(n29763), .B(n17105), .ZN(n17539) );
  NAND2_X1 U16728 ( .A1(n13196), .A2(n13194), .ZN(n31523) );
  NOR2_X1 U16754 ( .A1(n28733), .A2(n13151), .ZN(n8036) );
  NOR2_X1 U16758 ( .A1(n16123), .A2(n18667), .ZN(n18616) );
  AND2_X1 U16763 ( .A1(n29403), .A2(n20159), .Z(n13850) );
  INV_X2 U16774 ( .I(n20522), .ZN(n1059) );
  AND2_X1 U16780 ( .A1(n15601), .A2(n3462), .Z(n3465) );
  NAND3_X1 U16781 ( .A1(n5525), .A2(n19541), .A3(n11375), .ZN(n28162) );
  OAI21_X2 U16799 ( .A1(n28419), .A2(n8960), .B(n7365), .ZN(n7483) );
  NAND2_X1 U16807 ( .A1(n33207), .A2(n13384), .ZN(n32079) );
  NOR2_X1 U16811 ( .A1(n1055), .A2(n771), .ZN(n13263) );
  NOR2_X2 U16822 ( .A1(n33548), .A2(n33547), .ZN(n33546) );
  XOR2_X1 U16825 ( .A1(n6536), .A2(n31525), .Z(n33674) );
  XOR2_X1 U16827 ( .A1(n19735), .A2(n29058), .Z(n31525) );
  XOR2_X1 U16834 ( .A1(n15077), .A2(n15453), .Z(n31526) );
  NOR2_X1 U16837 ( .A1(n139), .A2(n32925), .ZN(n31527) );
  INV_X1 U16844 ( .I(n17347), .ZN(n29546) );
  NAND2_X1 U16852 ( .A1(n28577), .A2(n28578), .ZN(n33195) );
  CLKBUF_X4 U16859 ( .I(n18806), .Z(n3631) );
  AOI21_X2 U16876 ( .A1(n4528), .A2(n1132), .B(n4526), .ZN(n31528) );
  NAND2_X1 U16905 ( .A1(n26876), .A2(n32168), .ZN(n32167) );
  NOR2_X1 U16906 ( .A1(n26876), .A2(n36801), .ZN(n32170) );
  OR2_X1 U16928 ( .A1(n12428), .A2(n18720), .Z(n29470) );
  NOR2_X1 U16935 ( .A1(n28220), .A2(n4649), .ZN(n31774) );
  NAND2_X1 U16936 ( .A1(n31774), .A2(n1436), .ZN(n9236) );
  NAND2_X1 U16943 ( .A1(n15981), .A2(n17017), .ZN(n23570) );
  NOR2_X1 U16966 ( .A1(n11334), .A2(n26935), .ZN(n32958) );
  NAND3_X1 U16992 ( .A1(n30051), .A2(n9918), .A3(n1057), .ZN(n20170) );
  INV_X1 U16996 ( .I(n9918), .ZN(n30053) );
  OAI21_X1 U16998 ( .A1(n12156), .A2(n27009), .B(n5983), .ZN(n27558) );
  XNOR2_X1 U17000 ( .A1(n33243), .A2(n26448), .ZN(n31537) );
  CLKBUF_X2 U17005 ( .I(n27737), .Z(n32795) );
  OAI21_X1 U17006 ( .A1(n33006), .A2(n26974), .B(n5935), .ZN(n15708) );
  AND2_X1 U17027 ( .A1(n29600), .A2(n33746), .Z(n31540) );
  NAND2_X1 U17032 ( .A1(n20427), .A2(n19896), .ZN(n20426) );
  NAND2_X1 U17035 ( .A1(n29511), .A2(n29516), .ZN(n33428) );
  NAND2_X1 U17039 ( .A1(n19260), .A2(n29535), .ZN(n29511) );
  NAND4_X1 U17047 ( .A1(n2450), .A2(n2448), .A3(n9104), .A4(n29479), .ZN(
        n33463) );
  AOI21_X2 U17054 ( .A1(n23024), .A2(n23177), .B(n14130), .ZN(n23025) );
  XNOR2_X1 U17055 ( .A1(n34545), .A2(n22615), .ZN(n31541) );
  INV_X1 U17060 ( .I(n4604), .ZN(n32185) );
  NAND2_X1 U17062 ( .A1(n20288), .A2(n33358), .ZN(n20287) );
  INV_X2 U17067 ( .I(n6287), .ZN(n28453) );
  NAND2_X1 U17079 ( .A1(n1052), .A2(n18829), .ZN(n33565) );
  INV_X1 U17091 ( .I(n30432), .ZN(n31545) );
  INV_X1 U17092 ( .I(n8275), .ZN(n20623) );
  NOR2_X1 U17093 ( .A1(n22364), .A2(n8275), .ZN(n22226) );
  NAND2_X1 U17094 ( .A1(n29870), .A2(n773), .ZN(n18477) );
  NAND3_X1 U17100 ( .A1(n31624), .A2(n2029), .A3(n25927), .ZN(n11771) );
  INV_X1 U17103 ( .I(n2029), .ZN(n3277) );
  INV_X2 U17107 ( .I(n22264), .ZN(n14251) );
  NAND2_X1 U17109 ( .A1(n32759), .A2(n16108), .ZN(n11028) );
  NOR2_X1 U17110 ( .A1(n8166), .A2(n8798), .ZN(n31805) );
  NAND2_X1 U17120 ( .A1(n38749), .A2(n24515), .ZN(n32389) );
  INV_X1 U17127 ( .I(n5880), .ZN(n32467) );
  NAND2_X1 U17136 ( .A1(n8253), .A2(n5675), .ZN(n8251) );
  XOR2_X1 U17153 ( .A1(n18738), .A2(n18735), .Z(n31546) );
  NAND2_X1 U17160 ( .A1(n29413), .A2(n29410), .ZN(n32234) );
  OAI21_X1 U17169 ( .A1(n2335), .A2(n2334), .B(n33649), .ZN(n31548) );
  NAND2_X2 U17170 ( .A1(n21300), .A2(n33651), .ZN(n31549) );
  NAND3_X2 U17178 ( .A1(n10998), .A2(n10999), .A3(n27059), .ZN(n31551) );
  INV_X2 U17200 ( .I(n37632), .ZN(n18039) );
  AOI22_X1 U17202 ( .A1(n16596), .A2(n16597), .B1(n16595), .B2(n17369), .ZN(
        n32353) );
  AOI21_X1 U17208 ( .A1(n19272), .A2(n29555), .B(n29546), .ZN(n28904) );
  AND3_X2 U17209 ( .A1(n6408), .A2(n9500), .A3(n6409), .Z(n31552) );
  AND2_X1 U17216 ( .A1(n19700), .A2(n14459), .Z(n31555) );
  NOR2_X1 U17218 ( .A1(n10764), .A2(n26098), .ZN(n10765) );
  OAI22_X1 U17224 ( .A1(n33023), .A2(n18140), .B1(n14400), .B2(n29445), .ZN(
        n29448) );
  NAND2_X1 U17225 ( .A1(n32671), .A2(n29445), .ZN(n32670) );
  NOR2_X1 U17226 ( .A1(n16295), .A2(n33707), .ZN(n16494) );
  NAND2_X1 U17244 ( .A1(n14891), .A2(n18667), .ZN(n29262) );
  NAND2_X1 U17254 ( .A1(n33555), .A2(n28738), .ZN(n5968) );
  NAND2_X1 U17294 ( .A1(n7529), .A2(n8646), .ZN(n251) );
  NAND2_X1 U17303 ( .A1(n15649), .A2(n5028), .ZN(n31755) );
  NAND2_X1 U17309 ( .A1(n13730), .A2(n1226), .ZN(n6818) );
  NOR2_X1 U17314 ( .A1(n29980), .A2(n29968), .ZN(n32130) );
  INV_X1 U17330 ( .I(n9939), .ZN(n10385) );
  XOR2_X1 U17363 ( .A1(n16942), .A2(n20767), .Z(n31564) );
  NAND3_X2 U17366 ( .A1(n34116), .A2(n1781), .A3(n1777), .ZN(n31566) );
  INV_X1 U17374 ( .I(n29033), .ZN(n31720) );
  NAND2_X2 U17376 ( .A1(n16050), .A2(n16051), .ZN(n31568) );
  NOR2_X1 U17391 ( .A1(n5921), .A2(n29721), .ZN(n566) );
  XNOR2_X1 U17413 ( .A1(n8502), .A2(n26570), .ZN(n33165) );
  NAND2_X1 U17415 ( .A1(n1036), .A2(n12966), .ZN(n3048) );
  AND3_X2 U17423 ( .A1(n8591), .A2(n8590), .A3(n31980), .Z(n31569) );
  AND3_X2 U17424 ( .A1(n8591), .A2(n8590), .A3(n31980), .Z(n31570) );
  NAND2_X1 U17426 ( .A1(n13094), .A2(n13414), .ZN(n23440) );
  XOR2_X1 U17428 ( .A1(n5566), .A2(n5565), .Z(n31571) );
  INV_X1 U17432 ( .I(n13055), .ZN(n22399) );
  AOI21_X2 U17437 ( .A1(n1799), .A2(n4225), .B(n24862), .ZN(n1802) );
  XNOR2_X1 U17443 ( .A1(n9151), .A2(n33504), .ZN(n31575) );
  INV_X1 U17444 ( .I(n22968), .ZN(n23035) );
  INV_X1 U17454 ( .I(n27697), .ZN(n32811) );
  AND2_X2 U17459 ( .A1(n16699), .A2(n11092), .Z(n14947) );
  INV_X2 U17466 ( .I(n12892), .ZN(n9987) );
  NOR2_X1 U17469 ( .A1(n24432), .A2(n24431), .ZN(n15828) );
  OAI22_X2 U17486 ( .A1(n2842), .A2(n2841), .B1(n1671), .B2(n22182), .ZN(
        n31576) );
  INV_X1 U17504 ( .I(n22490), .ZN(n7118) );
  NAND2_X1 U17518 ( .A1(n9329), .A2(n15540), .ZN(n32284) );
  XOR2_X1 U17531 ( .A1(n20303), .A2(n24949), .Z(n31587) );
  AOI21_X1 U17543 ( .A1(n13952), .A2(n17022), .B(n13951), .ZN(n13950) );
  NOR2_X2 U17573 ( .A1(n12772), .A2(n24394), .ZN(n11213) );
  NOR2_X1 U17577 ( .A1(n29220), .A2(n10429), .ZN(n13106) );
  XOR2_X1 U17578 ( .A1(n4898), .A2(n6158), .Z(n31595) );
  XOR2_X1 U17580 ( .A1(n11017), .A2(n33850), .Z(n31596) );
  NAND2_X1 U17604 ( .A1(n23516), .A2(n19671), .ZN(n4737) );
  AOI21_X1 U17612 ( .A1(n23356), .A2(n39534), .B(n33696), .ZN(n24051) );
  OAI21_X1 U17630 ( .A1(n25860), .A2(n33997), .B(n33558), .ZN(n3807) );
  INV_X1 U17646 ( .I(n9862), .ZN(n15123) );
  XOR2_X1 U17648 ( .A1(n21346), .A2(Key[25]), .Z(n31604) );
  XOR2_X1 U17653 ( .A1(n10225), .A2(n10221), .Z(n31605) );
  NOR2_X1 U17664 ( .A1(n37632), .A2(n3462), .ZN(n31911) );
  AND2_X2 U17667 ( .A1(n17833), .A2(n6484), .Z(n21475) );
  INV_X1 U17669 ( .I(n17833), .ZN(n21476) );
  NAND2_X2 U17692 ( .A1(n28749), .A2(n28622), .ZN(n18990) );
  INV_X1 U17709 ( .I(n19478), .ZN(n14602) );
  NAND2_X1 U17714 ( .A1(n27936), .A2(n28109), .ZN(n33613) );
  NOR2_X1 U17721 ( .A1(n19768), .A2(n35973), .ZN(n21414) );
  XOR2_X1 U17736 ( .A1(n22200), .A2(n22201), .Z(n31617) );
  XOR2_X1 U17743 ( .A1(n31618), .A2(n18296), .Z(Ciphertext[186]) );
  AOI22_X1 U17746 ( .A1(n20074), .A2(n11701), .B1(n30247), .B2(n19663), .ZN(
        n31618) );
  NOR2_X1 U17747 ( .A1(n13258), .A2(n1722), .ZN(n21659) );
  XOR2_X1 U17748 ( .A1(n6447), .A2(Plaintext[134]), .Z(n13258) );
  INV_X1 U17756 ( .I(n29120), .ZN(n1061) );
  OAI21_X2 U17757 ( .A1(n24263), .A2(n31621), .B(n16645), .ZN(n24634) );
  NAND2_X2 U17764 ( .A1(n14766), .A2(n33552), .ZN(n28330) );
  XOR2_X1 U17767 ( .A1(n15114), .A2(n31622), .Z(n24247) );
  XOR2_X1 U17768 ( .A1(n23870), .A2(n23871), .Z(n31622) );
  NOR2_X2 U17789 ( .A1(n7324), .A2(n15792), .ZN(n28442) );
  NAND2_X2 U17791 ( .A1(n24672), .A2(n12418), .ZN(n25271) );
  XOR2_X1 U17839 ( .A1(n31636), .A2(n672), .Z(n4118) );
  NAND2_X2 U17844 ( .A1(n31637), .A2(n12124), .ZN(n15943) );
  XOR2_X1 U17852 ( .A1(n27579), .A2(n18650), .Z(n7829) );
  XOR2_X1 U17855 ( .A1(n1938), .A2(n27557), .Z(n27579) );
  OR2_X1 U17874 ( .A1(n7847), .A2(n24538), .Z(n32699) );
  OAI22_X1 U17879 ( .A1(n29552), .A2(n29551), .B1(n29549), .B2(n29550), .ZN(
        n29553) );
  NAND2_X1 U17888 ( .A1(n3979), .A2(n27401), .ZN(n31812) );
  AND2_X1 U17889 ( .A1(n16252), .A2(n32946), .Z(n31958) );
  AOI21_X2 U17899 ( .A1(n5686), .A2(n1103), .B(n5684), .ZN(n9576) );
  OR2_X1 U17908 ( .A1(n22499), .A2(n31649), .Z(n31648) );
  OAI21_X2 U17912 ( .A1(n16615), .A2(n7130), .B(n23154), .ZN(n23434) );
  BUF_X2 U17927 ( .I(n17499), .Z(n31651) );
  XOR2_X1 U17942 ( .A1(n31655), .A2(n23790), .Z(n19577) );
  NAND2_X2 U17949 ( .A1(n31656), .A2(n7799), .ZN(n29045) );
  XOR2_X1 U17952 ( .A1(n17417), .A2(n38228), .Z(n27807) );
  NOR3_X1 U17971 ( .A1(n15172), .A2(n14553), .A3(n9751), .ZN(n14779) );
  NAND2_X2 U17982 ( .A1(n6810), .A2(n17732), .ZN(n18785) );
  XNOR2_X1 U17991 ( .A1(n25181), .A2(n25086), .ZN(n15779) );
  NAND2_X2 U17999 ( .A1(n31665), .A2(n25889), .ZN(n17309) );
  OR2_X1 U18024 ( .A1(n27252), .A2(n36840), .Z(n31668) );
  OR2_X1 U18030 ( .A1(n2257), .A2(n22085), .Z(n5345) );
  NOR2_X2 U18032 ( .A1(n21481), .A2(n21480), .ZN(n2257) );
  NAND2_X2 U18042 ( .A1(n18591), .A2(n18594), .ZN(n22263) );
  XOR2_X1 U18047 ( .A1(n3655), .A2(n12233), .Z(n4556) );
  AOI22_X2 U18101 ( .A1(n29427), .A2(n1176), .B1(n15864), .B2(n357), .ZN(
        n29284) );
  OAI22_X2 U18102 ( .A1(n32671), .A2(n29445), .B1(n29446), .B2(n14422), .ZN(
        n29427) );
  NAND2_X2 U18106 ( .A1(n24646), .A2(n16238), .ZN(n24793) );
  XOR2_X1 U18116 ( .A1(n27001), .A2(n21176), .Z(n31682) );
  XOR2_X1 U18126 ( .A1(n31688), .A2(n16010), .Z(n16009) );
  NAND2_X1 U18150 ( .A1(n31693), .A2(n30127), .ZN(n11446) );
  NAND3_X1 U18170 ( .A1(n25756), .A2(n10563), .A3(n25754), .ZN(n31695) );
  XOR2_X1 U18179 ( .A1(n16336), .A2(n8654), .Z(n13189) );
  XOR2_X1 U18195 ( .A1(n29139), .A2(n28834), .Z(n10365) );
  NAND2_X1 U18206 ( .A1(n344), .A2(n21023), .ZN(n20290) );
  NAND2_X2 U18213 ( .A1(n16777), .A2(n30894), .ZN(n15015) );
  OR2_X1 U18217 ( .A1(n39815), .A2(n37045), .Z(n33217) );
  AOI21_X2 U18230 ( .A1(n31713), .A2(n31711), .B(n13428), .ZN(n7968) );
  AND2_X1 U18233 ( .A1(n29925), .A2(n29924), .Z(n31727) );
  NAND2_X2 U18241 ( .A1(n45), .A2(n23034), .ZN(n23119) );
  XOR2_X1 U18243 ( .A1(n8873), .A2(n31718), .Z(n31824) );
  XOR2_X1 U18244 ( .A1(n27678), .A2(n30404), .Z(n31718) );
  NAND2_X2 U18247 ( .A1(n5458), .A2(n5459), .ZN(n27687) );
  AOI22_X2 U18250 ( .A1(n2971), .A2(n1031), .B1(n2972), .B2(n2439), .ZN(n33730) );
  XOR2_X1 U18262 ( .A1(n27592), .A2(n12613), .Z(n27813) );
  NAND2_X2 U18263 ( .A1(n53), .A2(n9739), .ZN(n12613) );
  NAND2_X1 U18272 ( .A1(n31595), .A2(n30000), .ZN(n15328) );
  OAI21_X2 U18276 ( .A1(n12706), .A2(n2340), .B(n31723), .ZN(n16050) );
  XOR2_X1 U18280 ( .A1(n31725), .A2(n3666), .Z(n21235) );
  NOR2_X2 U18293 ( .A1(n5093), .A2(n16108), .ZN(n4697) );
  INV_X2 U18310 ( .I(n31731), .ZN(n4201) );
  XOR2_X1 U18319 ( .A1(n25255), .A2(n25001), .Z(n7958) );
  XOR2_X1 U18320 ( .A1(n25278), .A2(n6759), .Z(n25255) );
  NAND2_X2 U18342 ( .A1(n31736), .A2(n22526), .ZN(n23484) );
  NAND2_X2 U18346 ( .A1(n31737), .A2(n18608), .ZN(n24883) );
  NAND2_X1 U18348 ( .A1(n24125), .A2(n38812), .ZN(n31737) );
  XOR2_X1 U18352 ( .A1(n7958), .A2(n7957), .Z(n25683) );
  XOR2_X1 U18353 ( .A1(n27779), .A2(n4709), .Z(n11564) );
  NOR2_X1 U18398 ( .A1(n19893), .A2(n35172), .ZN(n31743) );
  XNOR2_X1 U18415 ( .A1(n16565), .A2(n27715), .ZN(n32181) );
  NOR2_X1 U18420 ( .A1(n13217), .A2(n13029), .ZN(n31749) );
  XOR2_X1 U18439 ( .A1(n31752), .A2(n10955), .Z(n14395) );
  INV_X2 U18445 ( .I(n39484), .ZN(n1222) );
  AOI22_X2 U18451 ( .A1(n5374), .A2(n27037), .B1(n13895), .B2(n5035), .ZN(
        n27566) );
  AOI22_X2 U18458 ( .A1(n23652), .A2(n36556), .B1(n32937), .B2(n31759), .ZN(
        n18983) );
  NAND2_X2 U18472 ( .A1(n9342), .A2(n9343), .ZN(n8026) );
  INV_X2 U18482 ( .I(n31760), .ZN(n32989) );
  XOR2_X1 U18485 ( .A1(n2695), .A2(n31762), .Z(n7993) );
  XOR2_X1 U18486 ( .A1(n18655), .A2(n23689), .Z(n31762) );
  OAI22_X1 U18487 ( .A1(n8691), .A2(n11701), .B1(n30250), .B2(n11700), .ZN(
        n32204) );
  NAND2_X2 U18490 ( .A1(n11700), .A2(n30262), .ZN(n8691) );
  XOR2_X1 U18515 ( .A1(n10430), .A2(n3140), .Z(n10390) );
  XOR2_X1 U18523 ( .A1(n16898), .A2(n31771), .Z(n22450) );
  INV_X2 U18525 ( .I(n10429), .ZN(n31772) );
  NAND2_X2 U18550 ( .A1(n32482), .A2(n17448), .ZN(n27284) );
  NAND2_X1 U18572 ( .A1(n7317), .A2(n692), .ZN(n11257) );
  XOR2_X1 U18585 ( .A1(n31779), .A2(n19407), .Z(Ciphertext[149]) );
  OAI22_X1 U18586 ( .A1(n30080), .A2(n30081), .B1(n19551), .B2(n19550), .ZN(
        n31779) );
  XOR2_X1 U18598 ( .A1(n19642), .A2(n35318), .Z(n11612) );
  OAI22_X2 U18625 ( .A1(n11639), .A2(n7494), .B1(n8411), .B2(n26623), .ZN(
        n10301) );
  INV_X2 U18626 ( .I(n31784), .ZN(n28279) );
  XOR2_X1 U18662 ( .A1(n13931), .A2(n26280), .Z(n31790) );
  NAND2_X2 U18673 ( .A1(n28387), .A2(n18259), .ZN(n28891) );
  XOR2_X1 U18686 ( .A1(n27861), .A2(n2138), .Z(n31794) );
  OAI21_X2 U18700 ( .A1(n25563), .A2(n25716), .B(n9132), .ZN(n25564) );
  NOR2_X2 U18707 ( .A1(n8693), .A2(n22468), .ZN(n23478) );
  NAND2_X1 U18714 ( .A1(n33457), .A2(n33456), .ZN(n3593) );
  XOR2_X1 U18717 ( .A1(n31801), .A2(n29321), .Z(Ciphertext[25]) );
  NAND2_X2 U18719 ( .A1(n13947), .A2(n13950), .ZN(n27404) );
  XOR2_X1 U18721 ( .A1(n828), .A2(n14644), .Z(n19830) );
  NOR3_X2 U18731 ( .A1(n31806), .A2(n31805), .A3(n37241), .ZN(n8169) );
  INV_X2 U18737 ( .I(n27810), .ZN(n31807) );
  OAI22_X2 U18754 ( .A1(n1183), .A2(n29815), .B1(n18222), .B2(n8677), .ZN(
        n14216) );
  NAND2_X1 U18759 ( .A1(n7173), .A2(n25379), .ZN(n32826) );
  XOR2_X1 U18773 ( .A1(n17627), .A2(n29092), .Z(n31811) );
  OR2_X1 U18775 ( .A1(n17032), .A2(n8604), .Z(n28042) );
  NAND3_X2 U18782 ( .A1(n11877), .A2(n22998), .A3(n20214), .ZN(n3256) );
  XOR2_X1 U18787 ( .A1(n7942), .A2(n22476), .Z(n31815) );
  NAND3_X2 U18803 ( .A1(n3070), .A2(n28134), .A3(n3069), .ZN(n28685) );
  XOR2_X1 U18818 ( .A1(n27501), .A2(n17349), .Z(n27678) );
  XOR2_X1 U18823 ( .A1(n31823), .A2(n38176), .Z(n12824) );
  INV_X2 U18824 ( .I(n26582), .ZN(n31823) );
  NOR3_X1 U18839 ( .A1(n28105), .A2(n1205), .A3(n5352), .ZN(n28106) );
  INV_X2 U18846 ( .I(n31824), .ZN(n20056) );
  NAND2_X2 U18866 ( .A1(n3861), .A2(n5579), .ZN(n29855) );
  NOR2_X2 U18867 ( .A1(n2346), .A2(n11830), .ZN(n3861) );
  XOR2_X1 U18869 ( .A1(n10371), .A2(n23743), .Z(n6388) );
  XOR2_X1 U18876 ( .A1(n19188), .A2(n31830), .Z(n33809) );
  NAND2_X2 U18879 ( .A1(n23219), .A2(n23218), .ZN(n23899) );
  NAND2_X1 U18889 ( .A1(n30041), .A2(n5348), .ZN(n7208) );
  XOR2_X1 U18908 ( .A1(n27687), .A2(n27736), .Z(n15548) );
  NAND2_X2 U18910 ( .A1(n6875), .A2(n6874), .ZN(n27736) );
  NAND2_X2 U18922 ( .A1(n31835), .A2(n23158), .ZN(n23430) );
  AND2_X1 U18927 ( .A1(n19768), .A2(n35973), .Z(n18592) );
  NOR2_X1 U18930 ( .A1(n2688), .A2(n9321), .ZN(n31836) );
  XOR2_X1 U18932 ( .A1(n1666), .A2(n1323), .Z(n6546) );
  NAND2_X2 U18951 ( .A1(n32851), .A2(n8019), .ZN(n27153) );
  OAI22_X2 U18952 ( .A1(n27350), .A2(n8830), .B1(n993), .B2(n19477), .ZN(
        n26749) );
  INV_X2 U18953 ( .I(n31840), .ZN(n26459) );
  XOR2_X1 U18954 ( .A1(n31841), .A2(n29152), .Z(n4354) );
  AOI22_X2 U18972 ( .A1(n17856), .A2(n14176), .B1(n31848), .B2(n31847), .ZN(
        n17751) );
  XOR2_X1 U18978 ( .A1(n31851), .A2(n23565), .Z(n18811) );
  NAND2_X2 U18979 ( .A1(n31852), .A2(n9280), .ZN(n24623) );
  XOR2_X1 U18981 ( .A1(n19807), .A2(n25171), .Z(n317) );
  NAND2_X2 U18985 ( .A1(n13161), .A2(n19158), .ZN(n22624) );
  AND2_X1 U18998 ( .A1(n8688), .A2(n8679), .Z(n31857) );
  NAND2_X2 U19001 ( .A1(n33163), .A2(n16301), .ZN(n32471) );
  XOR2_X1 U19004 ( .A1(n32528), .A2(n26517), .Z(n9301) );
  XOR2_X1 U19084 ( .A1(Plaintext[142]), .A2(Key[142]), .Z(n32370) );
  OAI22_X2 U19089 ( .A1(n6217), .A2(n23531), .B1(n23528), .B2(n6218), .ZN(
        n23554) );
  XOR2_X1 U19090 ( .A1(n17659), .A2(n31867), .Z(n14254) );
  XOR2_X1 U19097 ( .A1(n5520), .A2(n27733), .Z(n32361) );
  XOR2_X1 U19103 ( .A1(n23835), .A2(n7919), .Z(n31869) );
  INV_X1 U19109 ( .I(n21249), .ZN(n33547) );
  XOR2_X1 U19122 ( .A1(n19081), .A2(n26542), .Z(n26369) );
  NAND2_X2 U19125 ( .A1(n25972), .A2(n9811), .ZN(n26542) );
  XOR2_X1 U19129 ( .A1(n22457), .A2(n3622), .Z(n3621) );
  OAI22_X2 U19145 ( .A1(n1440), .A2(n27940), .B1(n11732), .B2(n2717), .ZN(
        n31876) );
  XOR2_X1 U19158 ( .A1(n31880), .A2(n32842), .Z(n2264) );
  AND2_X1 U19190 ( .A1(n16224), .A2(n14557), .Z(n12276) );
  XOR2_X1 U19211 ( .A1(n5177), .A2(n5176), .Z(n11617) );
  NAND2_X2 U19230 ( .A1(n16006), .A2(n16007), .ZN(n7485) );
  OAI21_X2 U19258 ( .A1(n37169), .A2(n31893), .B(n38317), .ZN(n19356) );
  XOR2_X1 U19271 ( .A1(n29090), .A2(n14099), .Z(n6164) );
  XOR2_X1 U19282 ( .A1(n1669), .A2(n22371), .Z(n22597) );
  INV_X2 U19297 ( .I(n31897), .ZN(n852) );
  XOR2_X1 U19302 ( .A1(n26373), .A2(n5444), .Z(n31897) );
  XNOR2_X1 U19308 ( .A1(n10811), .A2(n15384), .ZN(n29696) );
  XOR2_X1 U19318 ( .A1(n14039), .A2(n31898), .Z(n3552) );
  XOR2_X1 U19324 ( .A1(n32092), .A2(n2996), .Z(n29942) );
  NAND2_X2 U19325 ( .A1(n9197), .A2(n24879), .ZN(n18744) );
  AOI21_X2 U19329 ( .A1(n39321), .A2(n3101), .B(n31900), .ZN(n3175) );
  INV_X2 U19346 ( .I(n37105), .ZN(n32488) );
  XOR2_X1 U19369 ( .A1(n33178), .A2(n18577), .Z(n31909) );
  NOR2_X2 U19377 ( .A1(n5817), .A2(n10713), .ZN(n5871) );
  XOR2_X1 U19380 ( .A1(n2229), .A2(n33676), .Z(n33734) );
  XOR2_X1 U19394 ( .A1(n31914), .A2(n29690), .Z(Ciphertext[89]) );
  AOI22_X2 U19407 ( .A1(n32247), .A2(n1126), .B1(n31916), .B2(n17076), .ZN(
        n32956) );
  XOR2_X1 U19408 ( .A1(n8183), .A2(n25274), .Z(n4238) );
  NAND2_X2 U19420 ( .A1(n32089), .A2(n20972), .ZN(n6141) );
  XOR2_X1 U19436 ( .A1(n10225), .A2(n10221), .Z(n26494) );
  NAND2_X2 U19446 ( .A1(n20264), .A2(n31918), .ZN(n31948) );
  INV_X2 U19456 ( .I(n31920), .ZN(n12729) );
  NOR2_X1 U19481 ( .A1(n27278), .A2(n27279), .ZN(n31925) );
  NOR2_X1 U19485 ( .A1(n35217), .A2(n12049), .ZN(n10451) );
  AND2_X1 U19492 ( .A1(n23515), .A2(n38292), .Z(n2853) );
  XOR2_X1 U19498 ( .A1(n31927), .A2(n23888), .Z(n2806) );
  NAND3_X1 U19539 ( .A1(n33656), .A2(n21160), .A3(n30484), .ZN(n31932) );
  XOR2_X1 U19560 ( .A1(n27466), .A2(n27858), .Z(n12971) );
  INV_X1 U19564 ( .I(n23928), .ZN(n32383) );
  XOR2_X1 U19574 ( .A1(n22778), .A2(n31933), .Z(n22780) );
  OAI21_X2 U19604 ( .A1(n33281), .A2(n18962), .B(n12232), .ZN(n30184) );
  AOI22_X2 U19621 ( .A1(n21925), .A2(n21469), .B1(n4057), .B2(n11411), .ZN(
        n4056) );
  INV_X1 U19646 ( .I(n16610), .ZN(n1510) );
  NAND2_X2 U19655 ( .A1(n31940), .A2(n31939), .ZN(n22161) );
  INV_X2 U19658 ( .I(n22008), .ZN(n31939) );
  XOR2_X1 U19661 ( .A1(n26588), .A2(n16294), .Z(n26296) );
  XOR2_X1 U19662 ( .A1(n22687), .A2(n12730), .Z(n22490) );
  NAND2_X2 U19686 ( .A1(n4903), .A2(n31946), .ZN(n17094) );
  AOI21_X2 U19693 ( .A1(n13774), .A2(n18244), .B(n31947), .ZN(n31946) );
  INV_X4 U19696 ( .I(n21099), .ZN(n32168) );
  XOR2_X1 U19709 ( .A1(n22391), .A2(n22510), .Z(n8547) );
  AND3_X1 U19713 ( .A1(n13233), .A2(n12924), .A3(n21270), .Z(n13722) );
  XOR2_X1 U19732 ( .A1(n4624), .A2(n22598), .Z(n22392) );
  OAI22_X2 U19733 ( .A1(n7132), .A2(n20375), .B1(n22499), .B2(n7131), .ZN(
        n22598) );
  AND2_X1 U19740 ( .A1(n29365), .A2(n37096), .Z(n13274) );
  INV_X4 U19749 ( .I(n33140), .ZN(n14423) );
  AOI21_X1 U19751 ( .A1(n1473), .A2(n17142), .B(n35500), .ZN(n4089) );
  NOR2_X1 U19756 ( .A1(n85), .A2(n2242), .ZN(n12148) );
  NAND2_X2 U19776 ( .A1(n13500), .A2(n13498), .ZN(n27959) );
  NAND2_X1 U19788 ( .A1(n21446), .A2(n21445), .ZN(n21349) );
  NAND2_X1 U19802 ( .A1(n31967), .A2(n19252), .ZN(n33484) );
  OAI21_X1 U19805 ( .A1(n32129), .A2(n32130), .B(n18897), .ZN(n31967) );
  XOR2_X1 U19838 ( .A1(n27774), .A2(n27570), .Z(n27539) );
  XNOR2_X1 U19843 ( .A1(n12494), .A2(n12491), .ZN(n31971) );
  OAI21_X2 U19845 ( .A1(n31972), .A2(n33636), .B(n21673), .ZN(n11044) );
  XOR2_X1 U19847 ( .A1(n32106), .A2(n19897), .Z(n32766) );
  OR2_X1 U19850 ( .A1(n25114), .A2(n25097), .Z(n33896) );
  OAI21_X2 U19851 ( .A1(n20927), .A2(n20928), .B(n20925), .ZN(n25114) );
  INV_X2 U19855 ( .I(n31976), .ZN(n8529) );
  INV_X2 U19856 ( .I(n20960), .ZN(n10231) );
  INV_X2 U19859 ( .I(n31978), .ZN(n876) );
  XOR2_X1 U19885 ( .A1(n13954), .A2(n32022), .Z(n32678) );
  NOR2_X1 U19894 ( .A1(n17412), .A2(n32304), .ZN(n11677) );
  XOR2_X1 U19895 ( .A1(n8516), .A2(n8514), .Z(n32304) );
  INV_X2 U19913 ( .I(n3873), .ZN(n31982) );
  XOR2_X1 U19919 ( .A1(n17272), .A2(n30480), .Z(n31983) );
  NAND3_X2 U19920 ( .A1(n31985), .A2(n26659), .A3(n30352), .ZN(n27249) );
  NAND2_X1 U19922 ( .A1(n32142), .A2(n11864), .ZN(n31985) );
  OR2_X1 U19929 ( .A1(n2147), .A2(n28745), .Z(n18201) );
  NOR2_X2 U19935 ( .A1(n2347), .A2(n3861), .ZN(n29858) );
  INV_X2 U19951 ( .I(n27919), .ZN(n28215) );
  NOR2_X1 U19961 ( .A1(n6217), .A2(n23532), .ZN(n8269) );
  XOR2_X1 U19971 ( .A1(n23910), .A2(n23884), .Z(n23979) );
  OAI22_X2 U19989 ( .A1(n23200), .A2(n11354), .B1(n13527), .B2(n33247), .ZN(
        n33453) );
  NAND2_X1 U19990 ( .A1(n13181), .A2(n26876), .ZN(n13182) );
  AND2_X1 U19994 ( .A1(n4947), .A2(n5112), .Z(n32076) );
  AOI21_X1 U20005 ( .A1(n5681), .A2(n5680), .B(n927), .ZN(n4677) );
  XOR2_X1 U20010 ( .A1(n33812), .A2(n1510), .Z(n31999) );
  OR2_X1 U20011 ( .A1(n24597), .A2(n36321), .Z(n10056) );
  INV_X2 U20012 ( .I(n32001), .ZN(n167) );
  NAND3_X2 U20018 ( .A1(n18859), .A2(n32004), .A3(n33841), .ZN(n11534) );
  XOR2_X1 U20021 ( .A1(n12341), .A2(n29649), .Z(n2997) );
  XOR2_X1 U20026 ( .A1(n26518), .A2(n32003), .Z(n5765) );
  NAND2_X2 U20038 ( .A1(n28666), .A2(n33995), .ZN(n4120) );
  AOI21_X2 U20039 ( .A1(n10753), .A2(n953), .B(n32011), .ZN(n6965) );
  NAND2_X2 U20043 ( .A1(n32926), .A2(n36496), .ZN(n27244) );
  AND2_X1 U20067 ( .A1(n32881), .A2(n15257), .Z(n32018) );
  NAND2_X2 U20071 ( .A1(n28184), .A2(n28185), .ZN(n17397) );
  XOR2_X1 U20076 ( .A1(n8742), .A2(n27558), .Z(n3604) );
  XOR2_X1 U20090 ( .A1(n11919), .A2(n30483), .Z(n18580) );
  XOR2_X1 U20091 ( .A1(n27786), .A2(n15401), .Z(n11919) );
  XOR2_X1 U20094 ( .A1(n23784), .A2(n6091), .Z(n6090) );
  XOR2_X1 U20095 ( .A1(n24070), .A2(n23903), .Z(n23784) );
  OR2_X1 U20102 ( .A1(n38822), .A2(n20566), .Z(n13739) );
  XOR2_X1 U20108 ( .A1(n25222), .A2(n32033), .Z(n821) );
  XOR2_X1 U20111 ( .A1(n25076), .A2(n31552), .Z(n32033) );
  OR2_X1 U20114 ( .A1(n15350), .A2(n10632), .Z(n22340) );
  OR2_X1 U20130 ( .A1(n5282), .A2(n32391), .Z(n12946) );
  XOR2_X1 U20144 ( .A1(n23722), .A2(n30446), .Z(n24279) );
  XOR2_X1 U20156 ( .A1(n14359), .A2(n32049), .Z(n33958) );
  OR2_X1 U20161 ( .A1(n28463), .A2(n28464), .Z(n15709) );
  AOI21_X2 U20181 ( .A1(n32916), .A2(n6469), .B(n14578), .ZN(n3116) );
  XOR2_X1 U20182 ( .A1(n7944), .A2(n30775), .Z(n6142) );
  NAND2_X2 U20183 ( .A1(n7150), .A2(n7149), .ZN(n7944) );
  OAI21_X2 U20194 ( .A1(n4868), .A2(n4867), .B(n32052), .ZN(n32051) );
  XOR2_X1 U20196 ( .A1(n16356), .A2(n29514), .Z(n3299) );
  NAND2_X2 U20197 ( .A1(n16256), .A2(n16272), .ZN(n16356) );
  OAI22_X2 U20200 ( .A1(n15952), .A2(n919), .B1(n15951), .B2(n32412), .ZN(
        n22264) );
  XOR2_X1 U20226 ( .A1(n32387), .A2(n9976), .Z(n18345) );
  XOR2_X1 U20227 ( .A1(n4587), .A2(n4588), .Z(n21152) );
  XOR2_X1 U20269 ( .A1(n32071), .A2(n13327), .Z(n15598) );
  XOR2_X1 U20275 ( .A1(n27547), .A2(n15548), .Z(n32071) );
  OR2_X1 U20276 ( .A1(n32535), .A2(n28621), .Z(n9107) );
  XOR2_X1 U20282 ( .A1(n8559), .A2(n8558), .Z(n8557) );
  XOR2_X1 U20283 ( .A1(n26544), .A2(n17051), .Z(n33357) );
  NAND2_X2 U20292 ( .A1(n26948), .A2(n20223), .ZN(n26950) );
  NAND2_X2 U20295 ( .A1(n16896), .A2(n13210), .ZN(n10834) );
  XOR2_X1 U20297 ( .A1(n36595), .A2(n29602), .Z(n32073) );
  XOR2_X1 U20313 ( .A1(n11571), .A2(n5002), .Z(n11569) );
  XOR2_X1 U20315 ( .A1(n13630), .A2(n13234), .Z(n4671) );
  XOR2_X1 U20322 ( .A1(n22760), .A2(n30329), .Z(n32083) );
  INV_X2 U20332 ( .I(n7090), .ZN(n20774) );
  NAND2_X1 U20334 ( .A1(n18651), .A2(n18652), .ZN(n18420) );
  NAND2_X2 U20338 ( .A1(n32087), .A2(n15846), .ZN(n25136) );
  XOR2_X1 U20355 ( .A1(n24024), .A2(n12972), .Z(n32090) );
  XOR2_X1 U20383 ( .A1(n2995), .A2(n29161), .Z(n32092) );
  XOR2_X1 U20403 ( .A1(n23982), .A2(n13978), .Z(n23801) );
  NAND3_X1 U20408 ( .A1(n23161), .A2(n7071), .A3(n10436), .ZN(n10438) );
  AND2_X1 U20415 ( .A1(n13029), .A2(n23352), .Z(n16456) );
  XOR2_X1 U20423 ( .A1(n32097), .A2(n713), .Z(n32096) );
  AND3_X1 U20431 ( .A1(n13584), .A2(n1285), .A3(n32838), .Z(n14291) );
  NAND2_X1 U20432 ( .A1(n25068), .A2(n32101), .ZN(n25070) );
  XOR2_X1 U20451 ( .A1(n32103), .A2(n17402), .Z(n10375) );
  XOR2_X1 U20452 ( .A1(n13844), .A2(n22278), .Z(n17402) );
  NAND2_X1 U20458 ( .A1(n7955), .A2(n14423), .ZN(n20869) );
  NAND2_X1 U20466 ( .A1(n7778), .A2(n32388), .ZN(n2239) );
  XOR2_X1 U20468 ( .A1(n3638), .A2(n32110), .Z(n11784) );
  XOR2_X1 U20469 ( .A1(n3641), .A2(n20886), .Z(n32110) );
  XOR2_X1 U20482 ( .A1(n26205), .A2(n13324), .Z(n33039) );
  XOR2_X1 U20491 ( .A1(n32118), .A2(n12132), .Z(n32486) );
  XOR2_X1 U20501 ( .A1(n29071), .A2(n32120), .Z(n18159) );
  INV_X1 U20502 ( .I(n29371), .ZN(n32120) );
  XOR2_X1 U20511 ( .A1(n38226), .A2(n19845), .Z(n18510) );
  BUF_X2 U20520 ( .I(n33073), .Z(n32123) );
  OAI21_X1 U20530 ( .A1(n28049), .A2(n19410), .B(n19435), .ZN(n7409) );
  XOR2_X1 U20540 ( .A1(n32126), .A2(n32125), .Z(n8219) );
  XOR2_X1 U20541 ( .A1(n8199), .A2(n20678), .Z(n32125) );
  XOR2_X1 U20547 ( .A1(n27648), .A2(n27819), .Z(n32127) );
  XOR2_X1 U20555 ( .A1(n32128), .A2(n30442), .Z(n22887) );
  OAI22_X2 U20592 ( .A1(n34459), .A2(n28669), .B1(n33337), .B2(n14209), .ZN(
        n28798) );
  XOR2_X1 U20593 ( .A1(n27698), .A2(n32137), .Z(n17110) );
  INV_X2 U20597 ( .I(n755), .ZN(n14458) );
  XOR2_X1 U20605 ( .A1(n6124), .A2(n22670), .Z(n32972) );
  INV_X4 U20618 ( .I(n32141), .ZN(n9197) );
  NOR2_X2 U20621 ( .A1(n15069), .A2(n298), .ZN(n32141) );
  XOR2_X1 U20643 ( .A1(n6930), .A2(n14307), .Z(n28373) );
  XOR2_X1 U20652 ( .A1(n32149), .A2(n27721), .Z(n18447) );
  OAI22_X2 U20660 ( .A1(n8017), .A2(n32039), .B1(n8792), .B2(n11044), .ZN(
        n32151) );
  AOI22_X2 U20679 ( .A1(n32152), .A2(n19007), .B1(n24403), .B2(n13412), .ZN(
        n12307) );
  NAND2_X2 U20686 ( .A1(n25767), .A2(n9379), .ZN(n11293) );
  NAND2_X2 U20688 ( .A1(n35015), .A2(n5753), .ZN(n25767) );
  XOR2_X1 U20689 ( .A1(n32154), .A2(n15400), .Z(n32446) );
  XOR2_X1 U20694 ( .A1(n27636), .A2(n5650), .Z(n5649) );
  NOR2_X1 U20697 ( .A1(n29267), .A2(n29276), .ZN(n29268) );
  INV_X1 U20699 ( .I(n32176), .ZN(n33668) );
  NOR2_X1 U20700 ( .A1(n25585), .A2(n16867), .ZN(n32156) );
  NOR2_X1 U20703 ( .A1(n19609), .A2(n21823), .ZN(n21675) );
  XNOR2_X1 U20712 ( .A1(n23884), .A2(n1725), .ZN(n33232) );
  AOI21_X1 U20713 ( .A1(n15597), .A2(n18383), .B(n15598), .ZN(n17248) );
  INV_X2 U20742 ( .I(n32161), .ZN(n15359) );
  XOR2_X1 U20746 ( .A1(Plaintext[98]), .A2(Key[98]), .Z(n32161) );
  AOI21_X2 U20750 ( .A1(n21797), .A2(n1354), .B(n32162), .ZN(n16659) );
  NOR2_X2 U20752 ( .A1(n1354), .A2(n32163), .ZN(n32162) );
  INV_X2 U20754 ( .I(n15619), .ZN(n32164) );
  AOI21_X1 U20755 ( .A1(n34166), .A2(n27895), .B(n28290), .ZN(n14176) );
  NAND2_X2 U20770 ( .A1(n19687), .A2(n32166), .ZN(n27108) );
  XOR2_X1 U20799 ( .A1(n33243), .A2(n26448), .Z(n5639) );
  XOR2_X1 U20809 ( .A1(n183), .A2(n32181), .Z(n6285) );
  XOR2_X1 U20810 ( .A1(n3393), .A2(n3392), .Z(n15187) );
  NAND2_X1 U20819 ( .A1(n32234), .A2(n32423), .ZN(n32303) );
  XOR2_X1 U20845 ( .A1(n18310), .A2(n7113), .Z(n7112) );
  NAND2_X2 U20846 ( .A1(n7114), .A2(n8023), .ZN(n18310) );
  NAND2_X2 U20850 ( .A1(n4297), .A2(n4296), .ZN(n14139) );
  XOR2_X1 U20852 ( .A1(n25105), .A2(n5058), .Z(n25351) );
  BUF_X2 U20865 ( .I(n9470), .Z(n32186) );
  XOR2_X1 U20874 ( .A1(n32188), .A2(n20479), .Z(Ciphertext[28]) );
  AOI21_X1 U20875 ( .A1(n32303), .A2(n29406), .B(n32302), .ZN(n13329) );
  NAND3_X1 U20880 ( .A1(n18071), .A2(n17578), .A3(n14524), .ZN(n23133) );
  XOR2_X1 U20882 ( .A1(n33718), .A2(n8900), .Z(n15913) );
  XOR2_X1 U20894 ( .A1(n8163), .A2(n19932), .Z(n25150) );
  OR2_X2 U20913 ( .A1(n19226), .A2(n26921), .Z(n26920) );
  NAND2_X1 U20914 ( .A1(n4957), .A2(n14558), .ZN(n2675) );
  XOR2_X1 U20924 ( .A1(n29835), .A2(n29305), .Z(n32203) );
  INV_X4 U20929 ( .I(n32956), .ZN(n25048) );
  NOR2_X2 U20939 ( .A1(n28532), .A2(n11413), .ZN(n11412) );
  OAI21_X2 U20944 ( .A1(n32208), .A2(n11008), .B(n3438), .ZN(n8519) );
  XOR2_X1 U20954 ( .A1(n32308), .A2(n2529), .Z(n2527) );
  XOR2_X1 U20959 ( .A1(n32210), .A2(n2025), .Z(n15907) );
  OAI22_X2 U20963 ( .A1(n6517), .A2(n33864), .B1(n6519), .B2(n6518), .ZN(
        n32230) );
  XOR2_X1 U20973 ( .A1(n32211), .A2(n9446), .Z(n2297) );
  XOR2_X1 U20974 ( .A1(n23382), .A2(n23387), .Z(n32211) );
  NAND2_X2 U20998 ( .A1(n6506), .A2(n8683), .ZN(n8120) );
  NAND2_X2 U20999 ( .A1(n6171), .A2(n8121), .ZN(n6506) );
  XOR2_X1 U21001 ( .A1(n27782), .A2(n32217), .Z(n9401) );
  XOR2_X1 U21007 ( .A1(n27542), .A2(n32218), .Z(n32217) );
  XOR2_X1 U21024 ( .A1(n11880), .A2(n15010), .Z(n32219) );
  BUF_X2 U21046 ( .I(n23639), .Z(n32226) );
  XOR2_X1 U21053 ( .A1(n32227), .A2(n25201), .Z(n3645) );
  XOR2_X1 U21056 ( .A1(n3647), .A2(n25203), .Z(n32227) );
  INV_X1 U21059 ( .I(n28188), .ZN(n14376) );
  MUX2_X1 U21064 ( .I0(n13492), .I1(n28036), .S(n28188), .Z(n16567) );
  XOR2_X1 U21101 ( .A1(n27617), .A2(n31163), .Z(n27619) );
  NAND2_X1 U21106 ( .A1(n30793), .A2(n20078), .ZN(n6453) );
  NAND2_X2 U21109 ( .A1(n11676), .A2(n27910), .ZN(n15727) );
  XNOR2_X1 U21125 ( .A1(n36075), .A2(n16864), .ZN(n25264) );
  XOR2_X1 U21148 ( .A1(n8336), .A2(n8333), .Z(n13989) );
  MUX2_X1 U21168 ( .I0(n30210), .I1(n14387), .S(n30213), .Z(n15420) );
  XOR2_X1 U21172 ( .A1(n32354), .A2(n27710), .Z(n8335) );
  XNOR2_X1 U21173 ( .A1(n26538), .A2(n26339), .ZN(n5176) );
  NOR2_X1 U21183 ( .A1(n38732), .A2(n36991), .ZN(n25538) );
  AND2_X1 U21208 ( .A1(n5042), .A2(n32536), .Z(n13301) );
  XNOR2_X1 U21233 ( .A1(n14039), .A2(n29165), .ZN(n29022) );
  NAND3_X2 U21240 ( .A1(n12413), .A2(n3194), .A3(n3195), .ZN(n20509) );
  NOR2_X1 U21253 ( .A1(n23467), .A2(n23634), .ZN(n23421) );
  BUF_X2 U21258 ( .I(n6205), .Z(n32258) );
  OR2_X1 U21259 ( .A1(n25990), .A2(n38548), .Z(n32586) );
  OAI22_X1 U21270 ( .A1(n30214), .A2(n31549), .B1(n14869), .B2(n30211), .ZN(
        n32263) );
  NAND2_X1 U21272 ( .A1(n9445), .A2(n1379), .ZN(n11395) );
  INV_X4 U21301 ( .I(n12729), .ZN(n14409) );
  NAND2_X1 U21313 ( .A1(n32280), .A2(n26672), .ZN(n11220) );
  XOR2_X1 U21328 ( .A1(n14364), .A2(n32275), .Z(n10134) );
  XOR2_X1 U21329 ( .A1(n8940), .A2(n28500), .Z(n32275) );
  XOR2_X1 U21331 ( .A1(n39231), .A2(n30248), .Z(n13115) );
  XOR2_X1 U21333 ( .A1(n20609), .A2(n32276), .Z(n22904) );
  XOR2_X1 U21334 ( .A1(n20607), .A2(n22379), .Z(n32276) );
  NOR2_X1 U21337 ( .A1(n29654), .A2(n32290), .ZN(n19412) );
  XOR2_X1 U21349 ( .A1(n32106), .A2(n26402), .Z(n26433) );
  INV_X2 U21351 ( .I(n27417), .ZN(n1478) );
  XOR2_X1 U21353 ( .A1(n25079), .A2(n25283), .Z(n13596) );
  XOR2_X1 U21367 ( .A1(n7829), .A2(n30481), .Z(n7828) );
  NOR2_X1 U21375 ( .A1(n19563), .A2(n27180), .ZN(n32837) );
  NAND3_X1 U21382 ( .A1(n18832), .A2(n19743), .A3(n18144), .ZN(n20431) );
  XOR2_X1 U21413 ( .A1(n32288), .A2(n1708), .Z(Ciphertext[79]) );
  XOR2_X1 U21418 ( .A1(n635), .A2(n3241), .Z(n11219) );
  XOR2_X1 U21441 ( .A1(n32293), .A2(n6549), .Z(n6548) );
  AND3_X1 U21445 ( .A1(n14271), .A2(n1236), .A3(n26862), .Z(n32563) );
  XOR2_X1 U21451 ( .A1(n31591), .A2(n29411), .Z(n28950) );
  NAND2_X2 U21453 ( .A1(n9842), .A2(n32301), .ZN(n24782) );
  OAI21_X1 U21456 ( .A1(n32297), .A2(n11757), .B(n36272), .ZN(n32301) );
  INV_X2 U21474 ( .I(n26598), .ZN(n1504) );
  NAND2_X2 U21475 ( .A1(n26052), .A2(n26051), .ZN(n26598) );
  AND2_X1 U21481 ( .A1(n29405), .A2(n35272), .Z(n32302) );
  XOR2_X1 U21521 ( .A1(n38370), .A2(n35215), .Z(n32308) );
  INV_X1 U21540 ( .I(n22419), .ZN(n33806) );
  XOR2_X1 U21553 ( .A1(n32312), .A2(n15273), .Z(Ciphertext[104]) );
  OAI22_X1 U21554 ( .A1(n5468), .A2(n32050), .B1(n5467), .B2(n3377), .ZN(
        n32312) );
  INV_X2 U21556 ( .I(n33738), .ZN(n32313) );
  XOR2_X1 U21558 ( .A1(n15838), .A2(Plaintext[94]), .Z(n21885) );
  NOR2_X1 U21606 ( .A1(n25576), .A2(n25577), .ZN(n32325) );
  NOR2_X1 U21608 ( .A1(n23003), .A2(n19823), .ZN(n32327) );
  NAND2_X2 U21633 ( .A1(n32332), .A2(n13462), .ZN(n8059) );
  OR2_X1 U21645 ( .A1(n14500), .A2(n14426), .Z(n19290) );
  XOR2_X1 U21646 ( .A1(n25093), .A2(n25132), .Z(n20304) );
  NOR2_X2 U21647 ( .A1(n12208), .A2(n30410), .ZN(n25093) );
  XOR2_X1 U21662 ( .A1(n1324), .A2(n22615), .Z(n10797) );
  XOR2_X1 U21663 ( .A1(n32339), .A2(n850), .Z(n32986) );
  XOR2_X1 U21665 ( .A1(n32340), .A2(n19801), .Z(Ciphertext[18]) );
  OAI22_X1 U21667 ( .A1(n29268), .A2(n16233), .B1(n16232), .B2(n29278), .ZN(
        n32340) );
  NAND2_X2 U21679 ( .A1(n13741), .A2(n13742), .ZN(n24759) );
  XOR2_X1 U21680 ( .A1(n13383), .A2(n33037), .Z(n709) );
  OAI21_X2 U21690 ( .A1(n6270), .A2(n6271), .B(n21809), .ZN(n22238) );
  NOR3_X1 U21704 ( .A1(n32796), .A2(n13042), .A3(n23101), .ZN(n14578) );
  XOR2_X1 U21739 ( .A1(n32353), .A2(n29051), .Z(Ciphertext[80]) );
  XOR2_X1 U21748 ( .A1(n18004), .A2(n7028), .Z(n26442) );
  NAND2_X2 U21761 ( .A1(n2238), .A2(n2239), .ZN(n8537) );
  XOR2_X1 U21762 ( .A1(n32361), .A2(n5522), .Z(n12909) );
  OAI21_X2 U21771 ( .A1(n32584), .A2(n32585), .B(n28181), .ZN(n8087) );
  XOR2_X1 U21775 ( .A1(n32369), .A2(n27569), .Z(n11137) );
  XOR2_X1 U21776 ( .A1(n33587), .A2(n27676), .Z(n32369) );
  AOI21_X2 U21778 ( .A1(n17484), .A2(n17483), .B(n17482), .ZN(n32675) );
  INV_X4 U21781 ( .I(n3662), .ZN(n33669) );
  XOR2_X1 U21782 ( .A1(n25214), .A2(n35268), .Z(n3163) );
  XOR2_X1 U21788 ( .A1(n29044), .A2(n14820), .Z(n13177) );
  XOR2_X1 U21796 ( .A1(n32375), .A2(n16440), .Z(n16160) );
  XOR2_X1 U21815 ( .A1(n32382), .A2(n2474), .Z(n33193) );
  AOI22_X2 U21822 ( .A1(n20749), .A2(n33842), .B1(n28291), .B2(n5469), .ZN(
        n33059) );
  XOR2_X1 U21824 ( .A1(n24001), .A2(n24000), .Z(n32387) );
  XOR2_X1 U21825 ( .A1(n3525), .A2(n3522), .Z(n4352) );
  NOR2_X1 U21826 ( .A1(n7361), .A2(n13653), .ZN(n33905) );
  XOR2_X1 U21829 ( .A1(n32239), .A2(n4117), .Z(n23723) );
  NAND2_X1 U21838 ( .A1(n32390), .A2(n32389), .ZN(n12518) );
  AND2_X1 U21850 ( .A1(n23619), .A2(n10480), .Z(n15458) );
  NAND2_X2 U21854 ( .A1(n19537), .A2(n32394), .ZN(n13300) );
  XOR2_X1 U21867 ( .A1(n32396), .A2(n5719), .Z(n5012) );
  XOR2_X1 U21868 ( .A1(n23745), .A2(n30371), .Z(n32396) );
  XOR2_X1 U21869 ( .A1(n17006), .A2(n16004), .Z(n32890) );
  NAND2_X2 U21878 ( .A1(n4280), .A2(n17841), .ZN(n22711) );
  XNOR2_X1 U21913 ( .A1(n14888), .A2(n14887), .ZN(n32661) );
  AND2_X1 U21914 ( .A1(n23574), .A2(n12154), .Z(n5049) );
  XOR2_X1 U21915 ( .A1(n1923), .A2(n32402), .Z(n1921) );
  XOR2_X1 U21916 ( .A1(n14386), .A2(n30403), .Z(n32402) );
  NAND2_X2 U21919 ( .A1(n2701), .A2(n15959), .ZN(n15960) );
  AOI21_X1 U21925 ( .A1(n1654), .A2(n9472), .B(n39155), .ZN(n5436) );
  XOR2_X1 U21935 ( .A1(n1745), .A2(n29509), .Z(n9497) );
  XOR2_X1 U21940 ( .A1(n2651), .A2(n22616), .Z(n2650) );
  XOR2_X1 U21944 ( .A1(n12839), .A2(n35200), .Z(n18737) );
  INV_X2 U21946 ( .I(n1921), .ZN(n15461) );
  NAND2_X1 U21955 ( .A1(n21435), .A2(n21358), .ZN(n21665) );
  XOR2_X1 U21974 ( .A1(n20608), .A2(n33990), .Z(n20607) );
  NAND2_X1 U21983 ( .A1(n11515), .A2(n37098), .ZN(n8822) );
  NOR2_X2 U21994 ( .A1(n12443), .A2(n17314), .ZN(n9688) );
  XOR2_X1 U22016 ( .A1(n35196), .A2(n19805), .Z(n2119) );
  XOR2_X1 U22025 ( .A1(n6363), .A2(n22565), .Z(n32420) );
  XOR2_X1 U22034 ( .A1(n22608), .A2(n18446), .Z(n353) );
  AND2_X1 U22043 ( .A1(n32666), .A2(n29409), .Z(n32423) );
  INV_X1 U22046 ( .I(n37064), .ZN(n33926) );
  XOR2_X1 U22070 ( .A1(n17758), .A2(n26253), .Z(n26457) );
  NOR3_X2 U22076 ( .A1(n26035), .A2(n26036), .A3(n26239), .ZN(n17758) );
  XOR2_X1 U22081 ( .A1(n22609), .A2(n22733), .Z(n32431) );
  NOR2_X2 U22092 ( .A1(n25920), .A2(n25919), .ZN(n18862) );
  OAI21_X2 U22128 ( .A1(n1991), .A2(n1992), .B(n25332), .ZN(n4382) );
  NOR2_X2 U22146 ( .A1(n28551), .A2(n37758), .ZN(n8800) );
  XOR2_X1 U22156 ( .A1(n33559), .A2(n32440), .Z(n8116) );
  XOR2_X1 U22160 ( .A1(n33420), .A2(n30461), .Z(n32440) );
  XOR2_X1 U22161 ( .A1(n11887), .A2(n32441), .Z(n129) );
  XOR2_X1 U22166 ( .A1(n295), .A2(n32464), .Z(n32442) );
  XOR2_X1 U22168 ( .A1(n29151), .A2(n30488), .Z(n6158) );
  XOR2_X1 U22176 ( .A1(n12988), .A2(n32443), .Z(n11284) );
  XOR2_X1 U22180 ( .A1(n4419), .A2(n27754), .Z(n32443) );
  INV_X2 U22198 ( .I(n32446), .ZN(n33955) );
  XOR2_X1 U22200 ( .A1(n13791), .A2(n32447), .Z(n18688) );
  XOR2_X1 U22201 ( .A1(n27841), .A2(n18893), .Z(n32447) );
  NAND3_X1 U22208 ( .A1(n12259), .A2(n28147), .A3(n12258), .ZN(n17214) );
  BUF_X2 U22225 ( .I(n1722), .Z(n32456) );
  AOI21_X1 U22232 ( .A1(n19017), .A2(n9422), .B(n32457), .ZN(n21365) );
  XOR2_X1 U22250 ( .A1(n32460), .A2(n21294), .Z(Ciphertext[146]) );
  AOI21_X1 U22259 ( .A1(n20131), .A2(n20132), .B(n32462), .ZN(n20129) );
  OR2_X1 U22263 ( .A1(n27395), .A2(n9037), .Z(n32463) );
  XOR2_X1 U22274 ( .A1(n29023), .A2(n32465), .Z(n3938) );
  NOR2_X1 U22283 ( .A1(n38141), .A2(n39018), .ZN(n32466) );
  AOI22_X2 U22288 ( .A1(n4887), .A2(n18575), .B1(n9764), .B2(n9763), .ZN(n4886) );
  XOR2_X1 U22295 ( .A1(n32470), .A2(n29875), .Z(Ciphertext[120]) );
  OR3_X1 U22299 ( .A1(n17072), .A2(n14881), .A3(n31006), .Z(n26868) );
  NAND2_X1 U22311 ( .A1(n1403), .A2(n20102), .ZN(n15327) );
  NAND2_X2 U22312 ( .A1(n18113), .A2(n32481), .ZN(n26128) );
  XOR2_X1 U22317 ( .A1(n13439), .A2(n11098), .Z(n23852) );
  XOR2_X1 U22320 ( .A1(n24050), .A2(n39038), .Z(n33055) );
  INV_X2 U22365 ( .I(n32486), .ZN(n25639) );
  XOR2_X1 U22377 ( .A1(n32490), .A2(n19805), .Z(n3560) );
  OAI21_X2 U22378 ( .A1(n32495), .A2(n32494), .B(n39321), .ZN(n32871) );
  NOR2_X1 U22379 ( .A1(n1116), .A2(n21042), .ZN(n32494) );
  NAND2_X2 U22404 ( .A1(n17055), .A2(n18019), .ZN(n32535) );
  XOR2_X1 U22411 ( .A1(n16427), .A2(n25848), .Z(n32505) );
  INV_X2 U22418 ( .I(n20514), .ZN(n33491) );
  AOI21_X2 U22429 ( .A1(n17023), .A2(n17025), .B(n8989), .ZN(n8988) );
  XOR2_X1 U22441 ( .A1(n32512), .A2(n28631), .Z(n28899) );
  XOR2_X1 U22454 ( .A1(n8732), .A2(n32516), .Z(n19446) );
  XOR2_X1 U22459 ( .A1(n29039), .A2(n29159), .Z(n4223) );
  XOR2_X1 U22463 ( .A1(n10256), .A2(n7564), .Z(n28125) );
  XOR2_X1 U22466 ( .A1(n32519), .A2(n29711), .Z(Ciphertext[91]) );
  NAND3_X2 U22472 ( .A1(n20169), .A2(n10435), .A3(n20170), .ZN(n30079) );
  XOR2_X1 U22514 ( .A1(n23905), .A2(n16055), .Z(n8113) );
  AND2_X1 U22517 ( .A1(n15325), .A2(n23440), .Z(n32526) );
  MUX2_X1 U22526 ( .I0(n15867), .I1(n29797), .S(n3096), .Z(n5468) );
  XOR2_X1 U22562 ( .A1(n32532), .A2(n10447), .Z(n25700) );
  INV_X2 U22572 ( .I(n32534), .ZN(n33948) );
  XOR2_X1 U22581 ( .A1(n25243), .A2(n25218), .Z(n17606) );
  NAND2_X1 U22591 ( .A1(n19307), .A2(n15290), .ZN(n22791) );
  INV_X2 U22592 ( .I(n32537), .ZN(n15289) );
  XOR2_X1 U22610 ( .A1(n6211), .A2(n32540), .Z(n6550) );
  BUF_X2 U22619 ( .I(n21594), .Z(n32544) );
  AOI22_X2 U22631 ( .A1(n32546), .A2(n30544), .B1(n9268), .B2(n30768), .ZN(
        n27470) );
  XOR2_X1 U22639 ( .A1(n27767), .A2(n8059), .Z(n15736) );
  NOR2_X2 U22645 ( .A1(n27015), .A2(n32549), .ZN(n27221) );
  OR2_X1 U22651 ( .A1(n23234), .A2(n20788), .Z(n2953) );
  NOR2_X2 U22701 ( .A1(n14394), .A2(n26786), .ZN(n26720) );
  NAND2_X2 U22723 ( .A1(n3099), .A2(n3098), .ZN(n26194) );
  OR2_X1 U22724 ( .A1(n10338), .A2(n26695), .Z(n231) );
  NAND2_X2 U22725 ( .A1(n33142), .A2(n26270), .ZN(n18549) );
  INV_X2 U22745 ( .I(n32556), .ZN(n18077) );
  INV_X1 U22761 ( .I(n7742), .ZN(n32559) );
  XOR2_X1 U22769 ( .A1(n23911), .A2(n32562), .Z(n10771) );
  NAND2_X2 U22771 ( .A1(n18382), .A2(n18381), .ZN(n23911) );
  XOR2_X1 U22811 ( .A1(n32567), .A2(n4022), .Z(n14347) );
  XOR2_X1 U22813 ( .A1(n26324), .A2(n4021), .Z(n32567) );
  XOR2_X1 U22822 ( .A1(n19967), .A2(n34096), .Z(n13116) );
  XOR2_X1 U22826 ( .A1(n33176), .A2(n1262), .Z(n19967) );
  NAND2_X2 U22829 ( .A1(n16879), .A2(n14431), .ZN(n6180) );
  NAND3_X1 U22839 ( .A1(n29947), .A2(n29946), .A3(n39745), .ZN(n29948) );
  NAND3_X1 U22842 ( .A1(n11181), .A2(n17286), .A3(n31598), .ZN(n32572) );
  NAND2_X2 U22851 ( .A1(n4529), .A2(n6797), .ZN(n6795) );
  XOR2_X1 U22863 ( .A1(n19254), .A2(n29970), .Z(n33862) );
  NAND2_X2 U22870 ( .A1(n6808), .A2(n4917), .ZN(n19254) );
  INV_X4 U22875 ( .I(n25639), .ZN(n33130) );
  INV_X2 U22923 ( .I(n32579), .ZN(n9242) );
  XOR2_X1 U22927 ( .A1(n9400), .A2(n9401), .Z(n32579) );
  INV_X1 U22928 ( .I(n11353), .ZN(n28027) );
  XOR2_X1 U22938 ( .A1(n25193), .A2(n24932), .Z(n6306) );
  NAND2_X2 U22939 ( .A1(n15877), .A2(n24491), .ZN(n25193) );
  NOR2_X2 U22946 ( .A1(n33249), .A2(n34016), .ZN(n11703) );
  XOR2_X1 U22947 ( .A1(n32581), .A2(n8059), .Z(n13283) );
  INV_X2 U22949 ( .I(n33470), .ZN(n32581) );
  NAND2_X2 U22966 ( .A1(n4193), .A2(n3809), .ZN(n4192) );
  NOR2_X2 U22967 ( .A1(n18832), .A2(n12406), .ZN(n32584) );
  NAND2_X2 U22970 ( .A1(n8697), .A2(n32588), .ZN(n8742) );
  AND2_X1 U22997 ( .A1(n1627), .A2(n37088), .Z(n32594) );
  INV_X2 U22998 ( .I(n32599), .ZN(n9797) );
  INV_X2 U23021 ( .I(n22887), .ZN(n22804) );
  OAI21_X1 U23036 ( .A1(n29658), .A2(n29662), .B(n30295), .ZN(n17368) );
  XOR2_X1 U23139 ( .A1(n22642), .A2(n22441), .Z(n6610) );
  NAND2_X2 U23162 ( .A1(n17436), .A2(n17435), .ZN(n4613) );
  INV_X2 U23176 ( .I(n11702), .ZN(n32617) );
  NOR2_X1 U23178 ( .A1(n1816), .A2(n15839), .ZN(n21574) );
  NAND2_X2 U23179 ( .A1(n24339), .A2(n24340), .ZN(n8173) );
  NAND2_X1 U23183 ( .A1(n17424), .A2(n29500), .ZN(n32620) );
  NAND2_X1 U23203 ( .A1(n3452), .A2(n23071), .ZN(n32625) );
  OR2_X1 U23233 ( .A1(n5044), .A2(n6159), .Z(n11214) );
  XOR2_X1 U23246 ( .A1(n8281), .A2(n33158), .Z(n32638) );
  XOR2_X1 U23247 ( .A1(n32639), .A2(n32910), .Z(n20152) );
  NAND2_X2 U23252 ( .A1(n19694), .A2(n26977), .ZN(n27417) );
  OAI21_X2 U23257 ( .A1(n26250), .A2(n26251), .B(n20912), .ZN(n27361) );
  NAND3_X2 U23290 ( .A1(n32644), .A2(n17979), .A3(n32643), .ZN(n25218) );
  XOR2_X1 U23298 ( .A1(n30322), .A2(n4210), .Z(n17988) );
  AOI22_X2 U23325 ( .A1(n6058), .A2(n16363), .B1(n27979), .B2(n885), .ZN(
        n32650) );
  OAI21_X2 U23334 ( .A1(n17669), .A2(n17668), .B(n12243), .ZN(n12242) );
  NOR2_X1 U23374 ( .A1(n27213), .A2(n4847), .ZN(n11767) );
  NAND2_X2 U23380 ( .A1(n10723), .A2(n25728), .ZN(n32658) );
  INV_X2 U23388 ( .I(n17533), .ZN(n11283) );
  XOR2_X1 U23410 ( .A1(n9643), .A2(n36068), .Z(n32660) );
  XOR2_X1 U23416 ( .A1(n32662), .A2(n32661), .Z(n32708) );
  BUF_X2 U23424 ( .I(n21951), .Z(n32664) );
  NAND4_X1 U23455 ( .A1(n29403), .A2(n29401), .A3(n29402), .A4(n29400), .ZN(
        n32666) );
  NAND2_X2 U23456 ( .A1(n33468), .A2(n32667), .ZN(n22741) );
  AOI22_X2 U23462 ( .A1(n6081), .A2(n6083), .B1(n32477), .B2(n33986), .ZN(
        n24944) );
  OR2_X1 U23470 ( .A1(n1755), .A2(n20405), .Z(n33206) );
  XOR2_X1 U23510 ( .A1(n28780), .A2(n32678), .Z(n266) );
  OR2_X1 U23525 ( .A1(n24712), .A2(n7506), .Z(n24902) );
  XOR2_X1 U23537 ( .A1(n5836), .A2(n22735), .Z(n5835) );
  XOR2_X1 U23556 ( .A1(n25126), .A2(n606), .Z(n32685) );
  XOR2_X1 U23560 ( .A1(n33690), .A2(n27689), .Z(n32686) );
  NOR2_X2 U23571 ( .A1(n16945), .A2(n7062), .ZN(n6381) );
  XOR2_X1 U23572 ( .A1(n20706), .A2(n27745), .Z(n27791) );
  XOR2_X1 U23581 ( .A1(n27713), .A2(n27548), .Z(n13327) );
  NOR2_X1 U23604 ( .A1(n15280), .A2(n33678), .ZN(n33677) );
  XOR2_X1 U23610 ( .A1(n32698), .A2(n20166), .Z(n19605) );
  NAND2_X2 U23649 ( .A1(n4531), .A2(n28453), .ZN(n32702) );
  XOR2_X1 U23650 ( .A1(n27859), .A2(n11919), .Z(n12775) );
  INV_X2 U23652 ( .I(n32708), .ZN(n33431) );
  NAND2_X1 U23668 ( .A1(n17527), .A2(n17526), .ZN(n17525) );
  NOR2_X1 U23678 ( .A1(n22274), .A2(n15868), .ZN(n16364) );
  NOR2_X2 U23694 ( .A1(n5590), .A2(n5589), .ZN(n5588) );
  XOR2_X1 U23716 ( .A1(n32718), .A2(n19444), .Z(n21184) );
  NAND3_X1 U23728 ( .A1(n20597), .A2(n28758), .A3(n2022), .ZN(n104) );
  NOR2_X1 U23730 ( .A1(n18719), .A2(n37188), .ZN(n32719) );
  NAND2_X1 U23734 ( .A1(n6137), .A2(n26354), .ZN(n6136) );
  XOR2_X1 U23737 ( .A1(n17110), .A2(n9026), .Z(n17767) );
  OAI21_X1 U23811 ( .A1(n19398), .A2(n25429), .B(n25679), .ZN(n25396) );
  XOR2_X1 U23812 ( .A1(n39723), .A2(n29920), .Z(n14098) );
  XNOR2_X1 U23834 ( .A1(n4341), .A2(n28891), .ZN(n28838) );
  AOI21_X2 U23840 ( .A1(n37622), .A2(n1293), .B(n37064), .ZN(n2369) );
  NAND2_X1 U23845 ( .A1(n27137), .A2(n27347), .ZN(n8166) );
  NAND2_X2 U23877 ( .A1(n12077), .A2(n32675), .ZN(n22066) );
  XOR2_X1 U23883 ( .A1(n3117), .A2(n32746), .Z(n33967) );
  XOR2_X1 U23886 ( .A1(n29251), .A2(n29250), .Z(n32746) );
  INV_X2 U23890 ( .I(n32750), .ZN(n33963) );
  NAND2_X1 U23923 ( .A1(n902), .A2(n28772), .ZN(n515) );
  NAND2_X2 U23948 ( .A1(n17228), .A2(n17229), .ZN(n27046) );
  INV_X2 U23958 ( .I(n32760), .ZN(n293) );
  XOR2_X1 U23962 ( .A1(Key[3]), .A2(Plaintext[3]), .Z(n32760) );
  NOR2_X1 U23974 ( .A1(n24650), .A2(n36340), .ZN(n32761) );
  XOR2_X1 U24006 ( .A1(n3490), .A2(n3489), .Z(n13365) );
  XOR2_X1 U24009 ( .A1(Plaintext[150]), .A2(Key[150]), .Z(n33073) );
  NOR2_X1 U24026 ( .A1(n4631), .A2(n19059), .ZN(n32768) );
  XOR2_X1 U24033 ( .A1(n26489), .A2(n26338), .Z(n26538) );
  XOR2_X1 U24052 ( .A1(n16431), .A2(n13326), .Z(n32773) );
  NOR2_X2 U24069 ( .A1(n26863), .A2(n15037), .ZN(n14065) );
  NAND3_X2 U24071 ( .A1(n15137), .A2(n18771), .A3(n24663), .ZN(n24665) );
  NAND3_X2 U24073 ( .A1(n12646), .A2(n11104), .A3(n5066), .ZN(n32825) );
  XOR2_X1 U24075 ( .A1(n20107), .A2(n32779), .Z(n18183) );
  XOR2_X1 U24078 ( .A1(n26346), .A2(n15078), .Z(n32779) );
  XOR2_X1 U24079 ( .A1(n14393), .A2(n27739), .Z(n26169) );
  OR2_X1 U24090 ( .A1(n22256), .A2(n1342), .Z(n22258) );
  NAND2_X2 U24114 ( .A1(n14139), .A2(n22262), .ZN(n22080) );
  NAND2_X2 U24150 ( .A1(n22086), .A2(n2696), .ZN(n12964) );
  XOR2_X1 U24160 ( .A1(Plaintext[190]), .A2(Key[190]), .Z(n20685) );
  NOR2_X1 U24164 ( .A1(n20835), .A2(n33496), .ZN(n32798) );
  NAND2_X2 U24166 ( .A1(n32799), .A2(n2077), .ZN(n3540) );
  INV_X2 U24184 ( .I(n32805), .ZN(n19697) );
  XOR2_X1 U24187 ( .A1(n21218), .A2(n21216), .Z(n32805) );
  XOR2_X1 U24188 ( .A1(n23866), .A2(n23867), .Z(n2511) );
  INV_X2 U24192 ( .I(n32806), .ZN(n735) );
  XOR2_X1 U24194 ( .A1(n32807), .A2(n11947), .Z(n5103) );
  NAND3_X1 U24202 ( .A1(n22128), .A2(n3678), .A3(n15663), .ZN(n3677) );
  XOR2_X1 U24205 ( .A1(n7247), .A2(n24928), .Z(n9390) );
  XOR2_X1 U24210 ( .A1(n38816), .A2(n32811), .Z(n767) );
  NOR2_X2 U24214 ( .A1(n2362), .A2(n32814), .ZN(n32813) );
  AND2_X1 U24217 ( .A1(n26787), .A2(n26470), .Z(n32814) );
  XOR2_X1 U24224 ( .A1(n13193), .A2(n6561), .Z(n17680) );
  INV_X2 U24235 ( .I(n32821), .ZN(n33939) );
  INV_X2 U24240 ( .I(n32822), .ZN(n281) );
  NAND3_X1 U24251 ( .A1(n14132), .A2(n26134), .A3(n33909), .ZN(n14131) );
  OR2_X2 U24263 ( .A1(n37052), .A2(n13873), .Z(n25566) );
  OAI22_X2 U24268 ( .A1(n33586), .A2(n1591), .B1(n24244), .B2(n18329), .ZN(
        n15955) );
  OAI21_X2 U24272 ( .A1(n2333), .A2(n7539), .B(n28530), .ZN(n33649) );
  NAND2_X1 U24278 ( .A1(n34016), .A2(n7900), .ZN(n9287) );
  NAND2_X2 U24285 ( .A1(n7253), .A2(n7252), .ZN(n20156) );
  NOR2_X2 U24317 ( .A1(n17602), .A2(n17600), .ZN(n32829) );
  OR2_X1 U24327 ( .A1(n37093), .A2(n11678), .Z(n20808) );
  INV_X2 U24330 ( .I(n37086), .ZN(n19978) );
  OR2_X1 U24356 ( .A1(n8818), .A2(n33955), .Z(n8370) );
  OR2_X1 U24361 ( .A1(n29890), .A2(n6885), .Z(n17526) );
  AND2_X1 U24366 ( .A1(n17630), .A2(n23078), .Z(n32877) );
  NAND2_X1 U24368 ( .A1(n1424), .A2(n38860), .ZN(n32833) );
  OAI21_X2 U24383 ( .A1(n22275), .A2(n16351), .B(n17576), .ZN(n22761) );
  NAND2_X2 U24399 ( .A1(n19503), .A2(n19501), .ZN(n25900) );
  XOR2_X1 U24403 ( .A1(n35220), .A2(n32836), .Z(n14643) );
  INV_X1 U24405 ( .I(n29711), .ZN(n32836) );
  AOI22_X2 U24412 ( .A1(n17444), .A2(n16828), .B1(n14525), .B2(n29266), .ZN(
        n29271) );
  XOR2_X1 U24417 ( .A1(n35936), .A2(n38468), .Z(n24000) );
  XOR2_X1 U24435 ( .A1(n15450), .A2(n15220), .Z(n3028) );
  XOR2_X1 U24438 ( .A1(n6710), .A2(n33220), .Z(n8151) );
  AOI21_X1 U24453 ( .A1(n11181), .A2(n31533), .B(n15773), .ZN(n10831) );
  XOR2_X1 U24455 ( .A1(n29260), .A2(n28948), .Z(n28949) );
  NOR2_X1 U24496 ( .A1(n27964), .A2(n20157), .ZN(n14093) );
  NAND2_X1 U24515 ( .A1(n37064), .A2(n23256), .ZN(n2368) );
  AND2_X1 U24519 ( .A1(n15627), .A2(n31049), .Z(n32850) );
  OAI21_X1 U24531 ( .A1(n28380), .A2(n20494), .B(n37776), .ZN(n28381) );
  NAND2_X1 U24565 ( .A1(n18667), .A2(n30233), .ZN(n14789) );
  INV_X2 U24576 ( .I(n32855), .ZN(n14424) );
  XOR2_X1 U24580 ( .A1(Plaintext[133]), .A2(Key[133]), .Z(n32855) );
  INV_X2 U24589 ( .I(n32856), .ZN(n23125) );
  OAI21_X2 U24612 ( .A1(n32857), .A2(n21528), .B(n35071), .ZN(n2991) );
  NAND2_X2 U24615 ( .A1(n32860), .A2(n20629), .ZN(n24049) );
  AOI22_X2 U24616 ( .A1(n9621), .A2(n2692), .B1(n32616), .B2(n19119), .ZN(
        n32860) );
  OAI21_X2 U24629 ( .A1(n25497), .A2(n32867), .B(n14490), .ZN(n25899) );
  XOR2_X1 U24643 ( .A1(n29158), .A2(n17452), .Z(n6774) );
  NOR2_X1 U24645 ( .A1(n30069), .A2(n30071), .ZN(n30067) );
  XOR2_X1 U24649 ( .A1(n28971), .A2(n19904), .Z(n13954) );
  AOI21_X2 U24654 ( .A1(n33829), .A2(n33472), .B(n28445), .ZN(n28971) );
  NAND2_X2 U24666 ( .A1(n28140), .A2(n28119), .ZN(n28345) );
  OAI21_X2 U24740 ( .A1(n32878), .A2(n32877), .B(n23183), .ZN(n23349) );
  OAI21_X2 U24760 ( .A1(n23504), .A2(n1133), .B(n23505), .ZN(n32883) );
  XOR2_X1 U24762 ( .A1(n359), .A2(n22285), .Z(n18291) );
  XOR2_X1 U24785 ( .A1(n32884), .A2(n30122), .Z(Ciphertext[162]) );
  INV_X2 U24834 ( .I(n22131), .ZN(n32889) );
  INV_X2 U24843 ( .I(n1627), .ZN(n1132) );
  XOR2_X1 U24856 ( .A1(n36516), .A2(n10370), .Z(n16153) );
  INV_X2 U24868 ( .I(n32893), .ZN(n33933) );
  XOR2_X1 U24891 ( .A1(n33660), .A2(n26453), .Z(n17657) );
  XOR2_X1 U24903 ( .A1(n28979), .A2(n18522), .Z(n32895) );
  XOR2_X1 U24919 ( .A1(n38560), .A2(n32896), .Z(n3657) );
  XOR2_X1 U24920 ( .A1(n26537), .A2(n748), .Z(n8187) );
  OR2_X1 U24942 ( .A1(n20517), .A2(n35242), .Z(n15899) );
  XOR2_X1 U24951 ( .A1(n6477), .A2(n8409), .Z(n8408) );
  XOR2_X1 U24954 ( .A1(n32903), .A2(n37112), .Z(Ciphertext[183]) );
  XOR2_X1 U24970 ( .A1(n33399), .A2(n17134), .Z(n816) );
  AOI21_X2 U24980 ( .A1(n23546), .A2(n31644), .B(n23545), .ZN(n23880) );
  OAI22_X2 U25017 ( .A1(n21297), .A2(n1138), .B1(n21296), .B2(n23579), .ZN(
        n33698) );
  INV_X2 U25024 ( .I(n8372), .ZN(n27174) );
  XOR2_X1 U25035 ( .A1(n17493), .A2(n30408), .Z(n447) );
  XOR2_X1 U25039 ( .A1(n24038), .A2(n23808), .Z(n16030) );
  XOR2_X1 U25059 ( .A1(n23904), .A2(n24067), .Z(n19103) );
  NAND2_X2 U25071 ( .A1(n16636), .A2(n22868), .ZN(n33703) );
  XOR2_X1 U25077 ( .A1(n10012), .A2(n25323), .Z(n32910) );
  AOI21_X2 U25078 ( .A1(n32911), .A2(n25537), .B(n25536), .ZN(n17803) );
  AOI21_X2 U25095 ( .A1(n13149), .A2(n23578), .B(n23257), .ZN(n6054) );
  NAND3_X1 U25104 ( .A1(n1224), .A2(n27379), .A3(n27378), .ZN(n32913) );
  XOR2_X1 U25117 ( .A1(n20448), .A2(n33837), .Z(n14456) );
  XOR2_X1 U25119 ( .A1(n26528), .A2(n646), .Z(n32915) );
  MUX2_X1 U25149 ( .I0(n4306), .I1(n38419), .S(n33955), .Z(n8369) );
  OAI21_X2 U25176 ( .A1(n20469), .A2(n20468), .B(n21668), .ZN(n33929) );
  XOR2_X1 U25199 ( .A1(n7936), .A2(n680), .Z(n1986) );
  XOR2_X1 U25215 ( .A1(n12431), .A2(n12432), .Z(n6493) );
  NAND2_X2 U25229 ( .A1(n17502), .A2(n30595), .ZN(n33816) );
  NAND2_X2 U25255 ( .A1(n946), .A2(n948), .ZN(n32929) );
  AOI22_X2 U25267 ( .A1(n3543), .A2(n5380), .B1(n3542), .B2(n23032), .ZN(n3544) );
  XOR2_X1 U25276 ( .A1(n17129), .A2(n19198), .Z(n19955) );
  NAND2_X1 U25288 ( .A1(n30111), .A2(n35186), .ZN(n32933) );
  XOR2_X1 U25299 ( .A1(n26334), .A2(n16830), .Z(n32934) );
  AOI22_X2 U25317 ( .A1(n12080), .A2(n37089), .B1(n22244), .B2(n8679), .ZN(
        n2589) );
  OR3_X1 U25334 ( .A1(n21042), .A2(n25639), .A3(n841), .Z(n25360) );
  AOI21_X2 U25351 ( .A1(n22064), .A2(n1341), .B(n4045), .ZN(n4441) );
  NOR3_X2 U25370 ( .A1(n30340), .A2(n33453), .A3(n14606), .ZN(n18747) );
  NAND2_X2 U25381 ( .A1(n3993), .A2(n4324), .ZN(n9037) );
  AOI21_X1 U25393 ( .A1(n2211), .A2(n11344), .B(n22324), .ZN(n4619) );
  NAND2_X2 U25397 ( .A1(n18855), .A2(n4116), .ZN(n2008) );
  INV_X2 U25426 ( .I(n32951), .ZN(n14553) );
  OAI21_X2 U25427 ( .A1(n32953), .A2(n32952), .B(n28415), .ZN(n2270) );
  NOR2_X2 U25435 ( .A1(n9599), .A2(n1068), .ZN(n32953) );
  XOR2_X1 U25440 ( .A1(n33865), .A2(n17223), .Z(n8629) );
  NOR2_X1 U25448 ( .A1(n4682), .A2(n12952), .ZN(n9928) );
  XOR2_X1 U25450 ( .A1(n31822), .A2(n32955), .Z(n33372) );
  XOR2_X1 U25452 ( .A1(n15481), .A2(n15480), .Z(n32955) );
  AND2_X1 U25477 ( .A1(n29740), .A2(n29739), .Z(n33767) );
  XOR2_X1 U25508 ( .A1(n16296), .A2(n29269), .Z(n11525) );
  NAND2_X2 U25533 ( .A1(n28385), .A2(n28384), .ZN(n1775) );
  XOR2_X1 U25581 ( .A1(n33129), .A2(n22492), .Z(n11437) );
  NAND2_X2 U25597 ( .A1(n21534), .A2(n16930), .ZN(n133) );
  XNOR2_X1 U25599 ( .A1(n9858), .A2(n30085), .ZN(n33121) );
  NAND2_X1 U25614 ( .A1(n36548), .A2(n35273), .ZN(n32980) );
  XOR2_X1 U25617 ( .A1(n28837), .A2(n29301), .Z(n21084) );
  NAND3_X2 U25622 ( .A1(n37776), .A2(n6405), .A3(n28458), .ZN(n32983) );
  INV_X4 U25624 ( .I(n32984), .ZN(n27235) );
  INV_X2 U25625 ( .I(n32985), .ZN(n4083) );
  NAND2_X2 U25628 ( .A1(n20823), .A2(n27236), .ZN(n27829) );
  NAND2_X1 U25711 ( .A1(n25327), .A2(n25484), .ZN(n25374) );
  XOR2_X1 U25726 ( .A1(n27080), .A2(n27079), .Z(n7564) );
  OAI21_X2 U25727 ( .A1(n16283), .A2(n33004), .B(n584), .ZN(n20387) );
  NOR2_X1 U25728 ( .A1(n1151), .A2(n17118), .ZN(n33004) );
  XOR2_X1 U25739 ( .A1(n35404), .A2(n37112), .Z(n33005) );
  AND2_X1 U25755 ( .A1(n38198), .A2(n26055), .Z(n13731) );
  XOR2_X1 U25773 ( .A1(n5534), .A2(n20232), .Z(n33007) );
  NAND2_X1 U25778 ( .A1(n13522), .A2(n13521), .ZN(n33028) );
  INV_X2 U25784 ( .I(n33008), .ZN(n17097) );
  INV_X4 U25805 ( .I(n21308), .ZN(n33771) );
  OR2_X1 U25810 ( .A1(n10223), .A2(n3669), .Z(n33011) );
  NAND2_X2 U25821 ( .A1(n24630), .A2(n11271), .ZN(n24526) );
  XOR2_X1 U25829 ( .A1(n33013), .A2(n6049), .Z(n5350) );
  XOR2_X1 U25833 ( .A1(n10036), .A2(n30333), .Z(n33013) );
  OR2_X1 U25856 ( .A1(n16042), .A2(n27267), .Z(n33017) );
  INV_X2 U25881 ( .I(n33023), .ZN(n771) );
  NAND2_X1 U25886 ( .A1(n18439), .A2(n18440), .ZN(n20920) );
  NAND2_X2 U25905 ( .A1(n33028), .A2(n33700), .ZN(n13519) );
  XOR2_X1 U25914 ( .A1(n26146), .A2(n26147), .Z(n33029) );
  OAI21_X2 U25925 ( .A1(n11386), .A2(n7260), .B(n33030), .ZN(n26596) );
  NAND2_X2 U25929 ( .A1(n9111), .A2(n9112), .ZN(n9106) );
  NOR2_X2 U25930 ( .A1(n33034), .A2(n5810), .ZN(n5807) );
  OAI22_X1 U25931 ( .A1(n10747), .A2(n14379), .B1(n13584), .B2(n10659), .ZN(
        n11134) );
  XOR2_X1 U25941 ( .A1(n25267), .A2(n6411), .Z(n6410) );
  NOR2_X2 U25945 ( .A1(n37198), .A2(n7606), .ZN(n27010) );
  NAND2_X1 U25975 ( .A1(n28222), .A2(n200), .ZN(n33048) );
  XOR2_X1 U25978 ( .A1(n10957), .A2(n33049), .Z(n11266) );
  XOR2_X1 U25995 ( .A1(n24030), .A2(n19770), .Z(n33049) );
  INV_X1 U25996 ( .I(n26286), .ZN(n8558) );
  XOR2_X1 U25998 ( .A1(n26286), .A2(n26228), .Z(n26230) );
  NAND3_X2 U26005 ( .A1(n26869), .A2(n27393), .A3(n26868), .ZN(n27617) );
  BUF_X2 U26006 ( .I(n27365), .Z(n33050) );
  INV_X2 U26013 ( .I(n19605), .ZN(n28133) );
  NOR2_X1 U26018 ( .A1(n11013), .A2(n11044), .ZN(n11012) );
  INV_X2 U26027 ( .I(n33055), .ZN(n16523) );
  NAND2_X2 U26032 ( .A1(n24554), .A2(n33056), .ZN(n26075) );
  INV_X2 U26038 ( .I(n33057), .ZN(n2395) );
  NAND2_X2 U26077 ( .A1(n33092), .A2(n12879), .ZN(n10429) );
  XOR2_X1 U26093 ( .A1(n33067), .A2(n6057), .Z(n2000) );
  OAI21_X2 U26099 ( .A1(n13263), .A2(n17089), .B(n19244), .ZN(n29403) );
  NAND2_X2 U26103 ( .A1(n12684), .A2(n15708), .ZN(n6686) );
  AND2_X1 U26105 ( .A1(n26837), .A2(n13758), .Z(n15512) );
  XOR2_X1 U26116 ( .A1(n6307), .A2(n6304), .Z(n835) );
  OAI22_X2 U26128 ( .A1(n25510), .A2(n11834), .B1(n16247), .B2(n34574), .ZN(
        n26338) );
  OR2_X1 U26157 ( .A1(n33782), .A2(n22268), .Z(n33072) );
  OR2_X1 U26160 ( .A1(n12403), .A2(n8517), .Z(n17848) );
  OAI21_X2 U26184 ( .A1(n4473), .A2(n9155), .B(n15743), .ZN(n4159) );
  NAND2_X2 U26190 ( .A1(n3006), .A2(n23502), .ZN(n12822) );
  NAND2_X1 U26198 ( .A1(n2429), .A2(n5630), .ZN(n2428) );
  XOR2_X1 U26219 ( .A1(n28954), .A2(n29304), .Z(n28955) );
  XOR2_X1 U26228 ( .A1(n2511), .A2(n2510), .Z(n16816) );
  AND2_X1 U26231 ( .A1(n6652), .A2(n5970), .Z(n3612) );
  INV_X2 U26241 ( .I(n14318), .ZN(n26833) );
  XOR2_X1 U26247 ( .A1(n6007), .A2(n14319), .Z(n14318) );
  XOR2_X1 U26263 ( .A1(n21007), .A2(n2431), .Z(n20622) );
  INV_X2 U26265 ( .I(n4498), .ZN(n16328) );
  XNOR2_X1 U26270 ( .A1(n29134), .A2(n29135), .ZN(n4498) );
  XOR2_X1 U26273 ( .A1(n33385), .A2(n20117), .Z(n26747) );
  NOR2_X2 U26276 ( .A1(n33156), .A2(n3691), .ZN(n5449) );
  XOR2_X1 U26280 ( .A1(n9091), .A2(n7346), .Z(n13994) );
  NAND2_X2 U26287 ( .A1(n6669), .A2(n15707), .ZN(n22150) );
  XOR2_X1 U26294 ( .A1(n28867), .A2(n19160), .Z(n11017) );
  XOR2_X1 U26308 ( .A1(n18001), .A2(n30402), .Z(n22424) );
  XOR2_X1 U26319 ( .A1(n22174), .A2(n22567), .Z(n18597) );
  XOR2_X1 U26331 ( .A1(n7475), .A2(n17423), .Z(n23777) );
  NAND2_X2 U26334 ( .A1(n22914), .A2(n22913), .ZN(n17423) );
  OR2_X1 U26345 ( .A1(n13728), .A2(n21805), .Z(n10875) );
  XOR2_X1 U26346 ( .A1(n10929), .A2(Key[59]), .Z(n13728) );
  OR2_X1 U26381 ( .A1(n27854), .A2(n27498), .Z(n5695) );
  OAI21_X2 U26399 ( .A1(n18464), .A2(n14504), .B(n18463), .ZN(n11935) );
  NOR2_X1 U26400 ( .A1(n14011), .A2(n23637), .ZN(n7598) );
  XOR2_X1 U26404 ( .A1(Plaintext[57]), .A2(Key[57]), .Z(n7654) );
  XOR2_X1 U26405 ( .A1(n27765), .A2(n682), .Z(n33111) );
  XOR2_X1 U26438 ( .A1(n33118), .A2(n4589), .Z(n4588) );
  XOR2_X1 U26444 ( .A1(n7603), .A2(n20843), .Z(n33118) );
  OAI21_X1 U26459 ( .A1(n14708), .A2(n21302), .B(n15541), .ZN(n15542) );
  XOR2_X1 U26466 ( .A1(n13171), .A2(n33121), .Z(n33120) );
  XNOR2_X1 U26467 ( .A1(n26182), .A2(n25407), .ZN(n33131) );
  NOR2_X1 U26470 ( .A1(n33123), .A2(n30953), .ZN(n7384) );
  INV_X1 U26494 ( .I(n4306), .ZN(n898) );
  AND2_X1 U26496 ( .A1(n18261), .A2(n4306), .Z(n19139) );
  INV_X2 U26501 ( .I(n22566), .ZN(n33129) );
  NOR2_X2 U26503 ( .A1(n23600), .A2(n23601), .ZN(n23605) );
  XOR2_X1 U26530 ( .A1(n27840), .A2(n8896), .Z(n33133) );
  XNOR2_X1 U26536 ( .A1(n23661), .A2(n38350), .ZN(n33524) );
  XOR2_X1 U26545 ( .A1(n12411), .A2(n31575), .Z(n11903) );
  NAND2_X2 U26581 ( .A1(n7812), .A2(n7811), .ZN(n7810) );
  AOI22_X2 U26596 ( .A1(n10731), .A2(n19480), .B1(n30246), .B2(n39187), .ZN(
        n30257) );
  AND2_X1 U26599 ( .A1(n19341), .A2(n24394), .Z(n16448) );
  NOR2_X1 U26600 ( .A1(n38151), .A2(n14858), .ZN(n33139) );
  INV_X2 U26628 ( .I(n33144), .ZN(n862) );
  XOR2_X1 U26632 ( .A1(n29111), .A2(n8285), .Z(n8284) );
  NAND2_X2 U26633 ( .A1(n33145), .A2(n15817), .ZN(n22307) );
  NAND2_X2 U26634 ( .A1(n33413), .A2(n15816), .ZN(n33145) );
  NOR2_X1 U26635 ( .A1(n8165), .A2(n33146), .ZN(n12626) );
  NOR2_X2 U26640 ( .A1(n26744), .A2(n26745), .ZN(n27347) );
  INV_X2 U26642 ( .I(n33147), .ZN(n1816) );
  OAI22_X2 U26645 ( .A1(n1059), .A2(n20525), .B1(n30243), .B2(n30242), .ZN(
        n30191) );
  NAND2_X2 U26648 ( .A1(n17187), .A2(n17188), .ZN(n26559) );
  XOR2_X1 U26652 ( .A1(n23979), .A2(n11938), .Z(n11117) );
  NOR2_X2 U26665 ( .A1(n18087), .A2(n16934), .ZN(n22676) );
  NAND2_X2 U26672 ( .A1(n26833), .A2(n7527), .ZN(n26831) );
  NAND2_X2 U26674 ( .A1(n15184), .A2(n12923), .ZN(n4604) );
  XOR2_X1 U26706 ( .A1(n25193), .A2(n25090), .Z(n25265) );
  XOR2_X1 U26711 ( .A1(Plaintext[174]), .A2(Key[174]), .Z(n695) );
  XOR2_X1 U26715 ( .A1(n33153), .A2(n25150), .Z(n9557) );
  XOR2_X1 U26716 ( .A1(n24933), .A2(n16422), .Z(n33153) );
  OAI21_X1 U26720 ( .A1(n9668), .A2(n6287), .B(n38155), .ZN(n7296) );
  NOR2_X1 U26721 ( .A1(n6414), .A2(n6416), .ZN(n6776) );
  AND2_X1 U26733 ( .A1(n17249), .A2(n37351), .Z(n33156) );
  AND2_X1 U26736 ( .A1(n20026), .A2(n12829), .Z(n29385) );
  XOR2_X1 U26753 ( .A1(n28805), .A2(n28804), .Z(n30243) );
  XOR2_X1 U26755 ( .A1(n27650), .A2(n8280), .Z(n33158) );
  INV_X2 U26758 ( .I(n15718), .ZN(n20102) );
  XOR2_X1 U26759 ( .A1(n4898), .A2(n6158), .Z(n15718) );
  XOR2_X1 U26792 ( .A1(n16019), .A2(n29060), .Z(n8516) );
  XOR2_X1 U26824 ( .A1(n20618), .A2(n648), .Z(n33166) );
  INV_X2 U26839 ( .I(n33170), .ZN(n21546) );
  XOR2_X1 U26851 ( .A1(Key[109]), .A2(Plaintext[109]), .Z(n33170) );
  OR2_X1 U26871 ( .A1(n27385), .A2(n27064), .Z(n33340) );
  XOR2_X1 U26896 ( .A1(n20353), .A2(n20352), .Z(n22603) );
  XOR2_X1 U26912 ( .A1(n13634), .A2(n33400), .Z(n14191) );
  XOR2_X1 U26938 ( .A1(n23730), .A2(n23788), .Z(n33179) );
  XOR2_X1 U26942 ( .A1(Plaintext[7]), .A2(Key[7]), .Z(n33324) );
  NAND2_X2 U26945 ( .A1(n33180), .A2(n14572), .ZN(n1326) );
  NAND2_X2 U26958 ( .A1(n29473), .A2(n29470), .ZN(n7303) );
  XOR2_X1 U26969 ( .A1(n29168), .A2(n33183), .Z(n9707) );
  XOR2_X1 U26976 ( .A1(n15581), .A2(n33184), .Z(n33183) );
  NAND2_X1 U27006 ( .A1(n14946), .A2(n2189), .ZN(n33186) );
  XOR2_X1 U27011 ( .A1(n1817), .A2(n33188), .Z(n25569) );
  NOR3_X1 U27030 ( .A1(n1414), .A2(n28478), .A3(n38629), .ZN(n3056) );
  AOI22_X2 U27031 ( .A1(n21514), .A2(n21568), .B1(n15528), .B2(n33885), .ZN(
        n16961) );
  NOR2_X2 U27032 ( .A1(n3293), .A2(n3294), .ZN(n15528) );
  XOR2_X1 U27033 ( .A1(n38209), .A2(n26460), .Z(n11050) );
  XOR2_X1 U27057 ( .A1(n33192), .A2(n19775), .Z(Ciphertext[172]) );
  INV_X2 U27065 ( .I(n33193), .ZN(n2741) );
  XOR2_X1 U27069 ( .A1(n25166), .A2(n33198), .Z(n10971) );
  XOR2_X1 U27079 ( .A1(n25165), .A2(n25275), .Z(n33198) );
  XOR2_X1 U27127 ( .A1(n12988), .A2(n5744), .Z(n5743) );
  XOR2_X1 U27128 ( .A1(n2867), .A2(n27511), .Z(n12988) );
  XOR2_X1 U27133 ( .A1(n22458), .A2(n33215), .Z(n33936) );
  XOR2_X1 U27141 ( .A1(n22648), .A2(n33216), .Z(n33215) );
  NAND3_X2 U27148 ( .A1(n14206), .A2(n33217), .A3(n14392), .ZN(n14205) );
  XOR2_X1 U27158 ( .A1(n29822), .A2(n33219), .Z(n27881) );
  XOR2_X1 U27167 ( .A1(n31522), .A2(n15745), .Z(n33219) );
  XOR2_X1 U27172 ( .A1(n6709), .A2(n18604), .Z(n33220) );
  XOR2_X1 U27181 ( .A1(n26570), .A2(n33223), .Z(n14144) );
  XOR2_X1 U27183 ( .A1(n33812), .A2(n19432), .Z(n33223) );
  XNOR2_X1 U27184 ( .A1(n14272), .A2(n4117), .ZN(n792) );
  AND2_X1 U27186 ( .A1(n19978), .A2(n33384), .Z(n3011) );
  INV_X2 U27199 ( .I(n33227), .ZN(n22567) );
  OAI21_X2 U27202 ( .A1(n5576), .A2(n5577), .B(n33228), .ZN(n33227) );
  XOR2_X1 U27216 ( .A1(n18359), .A2(n17528), .Z(n12464) );
  XOR2_X1 U27225 ( .A1(n9932), .A2(n1509), .Z(n33233) );
  NAND2_X2 U27250 ( .A1(n23754), .A2(n5740), .ZN(n5897) );
  XOR2_X1 U27257 ( .A1(n5571), .A2(n30450), .Z(n2309) );
  XOR2_X1 U27264 ( .A1(n33239), .A2(n3346), .Z(n16284) );
  XOR2_X1 U27268 ( .A1(n34498), .A2(n23957), .Z(n33239) );
  XOR2_X1 U27271 ( .A1(n22697), .A2(n22698), .Z(n21163) );
  XOR2_X1 U27281 ( .A1(n4091), .A2(n4090), .Z(n33242) );
  NAND3_X2 U27309 ( .A1(n24608), .A2(n31161), .A3(n19255), .ZN(n18563) );
  NAND2_X2 U27377 ( .A1(n33246), .A2(n29697), .ZN(n29721) );
  XOR2_X1 U27386 ( .A1(n23890), .A2(n7833), .Z(n33248) );
  AND2_X1 U27391 ( .A1(n19349), .A2(n38669), .Z(n552) );
  BUF_X2 U27392 ( .I(n33506), .Z(n33249) );
  NAND2_X1 U27400 ( .A1(n4737), .A2(n7049), .ZN(n13005) );
  NAND3_X1 U27406 ( .A1(n15822), .A2(n15823), .A3(n20423), .ZN(n33567) );
  OAI22_X2 U27460 ( .A1(n33257), .A2(n2102), .B1(n23096), .B2(n1144), .ZN(
        n23516) );
  NAND2_X2 U27475 ( .A1(n9225), .A2(n9222), .ZN(n22542) );
  XOR2_X1 U27477 ( .A1(n21376), .A2(Key[68]), .Z(n33506) );
  NAND2_X1 U27508 ( .A1(n27158), .A2(n27159), .ZN(n33262) );
  OR2_X1 U27517 ( .A1(n23473), .A2(n32601), .Z(n15462) );
  BUF_X2 U27545 ( .I(n19644), .Z(n33268) );
  XOR2_X1 U27566 ( .A1(n15339), .A2(n33273), .Z(n33272) );
  OR2_X1 U27570 ( .A1(n13055), .A2(n22243), .Z(n2588) );
  AND2_X1 U27593 ( .A1(n22118), .A2(n22117), .Z(n33282) );
  NAND2_X2 U27616 ( .A1(n18216), .A2(n2954), .ZN(n33284) );
  INV_X4 U27623 ( .I(n33286), .ZN(n2341) );
  OR2_X1 U27639 ( .A1(n22035), .A2(n33288), .Z(n18953) );
  NOR2_X1 U27644 ( .A1(n9486), .A2(n9484), .ZN(n33291) );
  XOR2_X1 U27660 ( .A1(n28913), .A2(n33295), .Z(n17906) );
  XOR2_X1 U27661 ( .A1(n36905), .A2(n5862), .Z(n33295) );
  XOR2_X1 U27663 ( .A1(n29065), .A2(n33296), .Z(n17326) );
  XOR2_X1 U27671 ( .A1(n29144), .A2(n19624), .Z(n33296) );
  AOI21_X2 U27675 ( .A1(n29873), .A2(n29869), .B(n33297), .ZN(n29890) );
  AND2_X1 U27680 ( .A1(n15463), .A2(n16593), .Z(n22871) );
  XOR2_X1 U27715 ( .A1(n33300), .A2(n33299), .Z(n846) );
  INV_X1 U27721 ( .I(n9989), .ZN(n33299) );
  XOR2_X1 U27723 ( .A1(n19879), .A2(n1009), .Z(n33300) );
  NAND2_X2 U27731 ( .A1(n25874), .A2(n36546), .ZN(n25876) );
  OAI22_X2 U27735 ( .A1(n33303), .A2(n9156), .B1(n26788), .B2(n26720), .ZN(
        n27365) );
  OAI21_X2 U27739 ( .A1(n14002), .A2(n14003), .B(n14001), .ZN(n14941) );
  XOR2_X1 U27744 ( .A1(n22610), .A2(n32836), .Z(n14610) );
  NAND2_X2 U27758 ( .A1(n8662), .A2(n22398), .ZN(n22610) );
  XOR2_X1 U27769 ( .A1(n27645), .A2(n33310), .Z(n33309) );
  INV_X2 U27781 ( .I(n20829), .ZN(n33310) );
  XOR2_X1 U27787 ( .A1(n33398), .A2(n33311), .Z(n8748) );
  XOR2_X1 U27798 ( .A1(n27598), .A2(n16972), .Z(n33313) );
  XOR2_X1 U27805 ( .A1(n33315), .A2(n22550), .Z(n7120) );
  OR2_X1 U27808 ( .A1(n37043), .A2(n10334), .Z(n15230) );
  BUF_X2 U27841 ( .I(n6426), .Z(n33318) );
  OR2_X1 U27845 ( .A1(n25537), .A2(n25484), .Z(n25464) );
  XOR2_X1 U27851 ( .A1(n15056), .A2(n33319), .Z(n881) );
  XOR2_X1 U27854 ( .A1(n27672), .A2(n33320), .Z(n33319) );
  INV_X1 U27867 ( .I(n29562), .ZN(n33320) );
  XOR2_X1 U27887 ( .A1(n5553), .A2(n26605), .Z(n13544) );
  XOR2_X1 U27890 ( .A1(n15609), .A2(n30448), .Z(n407) );
  INV_X2 U27901 ( .I(n28456), .ZN(n33325) );
  NAND2_X2 U27913 ( .A1(n1823), .A2(n28434), .ZN(n28456) );
  INV_X2 U27932 ( .I(n33326), .ZN(n892) );
  INV_X1 U27940 ( .I(n1010), .ZN(n26142) );
  XOR2_X1 U27991 ( .A1(n18733), .A2(n17884), .Z(n33334) );
  XOR2_X1 U27994 ( .A1(n8920), .A2(n25329), .Z(n13012) );
  XOR2_X1 U28003 ( .A1(n39756), .A2(n38993), .Z(n24981) );
  MUX2_X1 U28004 ( .I0(n29662), .I1(n29659), .S(n19297), .Z(n16595) );
  XOR2_X1 U28022 ( .A1(n11137), .A2(n7353), .Z(n11136) );
  OR2_X1 U28030 ( .A1(n15281), .A2(n10667), .Z(n5934) );
  INV_X2 U28070 ( .I(n28596), .ZN(n1418) );
  NAND2_X2 U28071 ( .A1(n10150), .A2(n10151), .ZN(n28596) );
  INV_X1 U28109 ( .I(n8365), .ZN(n33346) );
  XOR2_X1 U28119 ( .A1(n33350), .A2(n37109), .Z(Ciphertext[7]) );
  OAI21_X1 U28166 ( .A1(n33946), .A2(n7705), .B(n25429), .ZN(n7956) );
  AOI21_X2 U28168 ( .A1(n4423), .A2(n10408), .B(n33355), .ZN(n12198) );
  OAI21_X2 U28172 ( .A1(n30225), .A2(n33963), .B(n33362), .ZN(n33355) );
  NOR2_X1 U28173 ( .A1(n19157), .A2(n29409), .ZN(n29397) );
  XOR2_X1 U28199 ( .A1(n24632), .A2(n24631), .Z(n24633) );
  NAND2_X1 U28227 ( .A1(n29980), .A2(n33360), .ZN(n7271) );
  NOR2_X1 U28245 ( .A1(n29979), .A2(n29968), .ZN(n33360) );
  INV_X1 U28268 ( .I(n21331), .ZN(n33363) );
  XOR2_X1 U28313 ( .A1(n27751), .A2(n18122), .Z(n33364) );
  OAI22_X2 U28390 ( .A1(n33366), .A2(n33365), .B1(n6220), .B2(n32974), .ZN(
        n2915) );
  XOR2_X1 U28426 ( .A1(n25122), .A2(n25121), .Z(n25490) );
  XNOR2_X1 U28452 ( .A1(n6527), .A2(n24025), .ZN(n10413) );
  XOR2_X1 U28461 ( .A1(n22571), .A2(n33371), .Z(n11498) );
  XOR2_X1 U28470 ( .A1(n22588), .A2(n11500), .Z(n33371) );
  XOR2_X1 U28475 ( .A1(n15118), .A2(n30455), .Z(n23214) );
  OAI21_X2 U28525 ( .A1(n31550), .A2(n8473), .B(n33375), .ZN(n14221) );
  NAND2_X2 U28551 ( .A1(n20910), .A2(n20911), .ZN(n23523) );
  AOI21_X1 U28571 ( .A1(n2846), .A2(n27167), .B(n6908), .ZN(n33380) );
  NAND3_X2 U28622 ( .A1(n23291), .A2(n23289), .A3(n23290), .ZN(n24047) );
  XOR2_X1 U28629 ( .A1(n11190), .A2(n19848), .Z(n22607) );
  XOR2_X1 U28643 ( .A1(n12613), .A2(n29334), .Z(n10057) );
  XOR2_X1 U28656 ( .A1(n36958), .A2(n26504), .Z(n33388) );
  OAI21_X2 U28657 ( .A1(n21639), .A2(n21638), .B(n33389), .ZN(n22362) );
  XOR2_X1 U28658 ( .A1(n25102), .A2(n25103), .Z(n25105) );
  XOR2_X1 U28668 ( .A1(n9036), .A2(n19648), .Z(n3668) );
  BUF_X2 U28708 ( .I(n26018), .Z(n33395) );
  NAND3_X2 U28750 ( .A1(n25530), .A2(n25528), .A3(n25529), .ZN(n25797) );
  BUF_X2 U28758 ( .I(n9185), .Z(n33398) );
  XOR2_X1 U28825 ( .A1(n10427), .A2(n10426), .Z(n10282) );
  AOI21_X2 U28830 ( .A1(n21543), .A2(n19822), .B(n33402), .ZN(n16760) );
  NOR2_X1 U28834 ( .A1(n16762), .A2(n21702), .ZN(n33402) );
  XOR2_X1 U28851 ( .A1(n11667), .A2(n7603), .Z(n26276) );
  XOR2_X1 U28864 ( .A1(n27810), .A2(n19649), .Z(n11997) );
  XOR2_X1 U28909 ( .A1(n5635), .A2(n33410), .Z(n13725) );
  XOR2_X1 U28912 ( .A1(n11883), .A2(n11882), .Z(n33410) );
  NAND2_X2 U28932 ( .A1(n18938), .A2(n18936), .ZN(n5056) );
  NAND2_X2 U28978 ( .A1(n21886), .A2(n547), .ZN(n1847) );
  XOR2_X1 U28993 ( .A1(n17310), .A2(n33415), .Z(n22693) );
  AOI21_X1 U29004 ( .A1(n29739), .A2(n29755), .B(n29756), .ZN(n33416) );
  OAI21_X2 U29007 ( .A1(n3199), .A2(n7635), .B(n33418), .ZN(n28620) );
  XOR2_X1 U29017 ( .A1(n33419), .A2(n29399), .Z(Ciphertext[37]) );
  AOI22_X1 U29020 ( .A1(n29398), .A2(n29414), .B1(n29397), .B2(n29410), .ZN(
        n33419) );
  XOR2_X1 U29022 ( .A1(n5841), .A2(n7917), .Z(n33420) );
  INV_X2 U29028 ( .I(n11136), .ZN(n12406) );
  XOR2_X1 U29037 ( .A1(n14385), .A2(n14374), .Z(n9567) );
  XOR2_X1 U29046 ( .A1(n18363), .A2(n18317), .Z(n18316) );
  XOR2_X1 U29052 ( .A1(n33426), .A2(n10823), .Z(n2196) );
  XOR2_X1 U29053 ( .A1(n9989), .A2(n26440), .Z(n33426) );
  OR2_X1 U29078 ( .A1(n2741), .A2(n12519), .Z(n13114) );
  XOR2_X1 U29083 ( .A1(n26227), .A2(n18399), .Z(n26492) );
  NAND2_X2 U29101 ( .A1(n25477), .A2(n25479), .ZN(n25335) );
  XOR2_X1 U29131 ( .A1(n3790), .A2(n3791), .Z(n33429) );
  INV_X2 U29132 ( .I(n37117), .ZN(n30145) );
  NOR2_X2 U29158 ( .A1(n23245), .A2(n23244), .ZN(n23695) );
  INV_X4 U29278 ( .I(n33512), .ZN(n15643) );
  INV_X2 U29300 ( .I(n33446), .ZN(n33950) );
  NAND2_X2 U29332 ( .A1(n21247), .A2(n11970), .ZN(n21246) );
  NAND2_X1 U29393 ( .A1(n1596), .A2(n30833), .ZN(n33456) );
  NAND2_X2 U29396 ( .A1(n10937), .A2(n24172), .ZN(n33459) );
  OR2_X1 U29410 ( .A1(n15044), .A2(n29409), .Z(n14517) );
  NAND2_X2 U29465 ( .A1(n33911), .A2(n33462), .ZN(n3601) );
  XOR2_X1 U29469 ( .A1(n33463), .A2(n19760), .Z(Ciphertext[49]) );
  INV_X1 U29477 ( .I(n26060), .ZN(n33464) );
  XOR2_X1 U29508 ( .A1(n27689), .A2(n29206), .Z(n3114) );
  XOR2_X1 U29519 ( .A1(n8037), .A2(n8038), .Z(n33466) );
  XOR2_X1 U29544 ( .A1(n762), .A2(n30478), .Z(n11814) );
  NAND2_X2 U29562 ( .A1(n29181), .A2(n33476), .ZN(n18829) );
  XOR2_X1 U29565 ( .A1(n21055), .A2(n29143), .Z(n33478) );
  NAND2_X1 U29566 ( .A1(n20184), .A2(n13499), .ZN(n13498) );
  INV_X2 U29567 ( .I(n33479), .ZN(n21099) );
  AOI22_X1 U29593 ( .A1(n30263), .A2(n13786), .B1(n30261), .B2(n31529), .ZN(
        n7681) );
  XOR2_X1 U29606 ( .A1(n33484), .A2(n1162), .Z(Ciphertext[134]) );
  NAND2_X2 U29639 ( .A1(n33487), .A2(n22163), .ZN(n16667) );
  NOR2_X2 U29642 ( .A1(n19195), .A2(n19197), .ZN(n29981) );
  NOR3_X2 U29709 ( .A1(n7610), .A2(n12388), .A3(n24850), .ZN(n14385) );
  CLKBUF_X12 U29723 ( .I(n15159), .Z(n33495) );
  OAI22_X1 U29765 ( .A1(n29007), .A2(n17192), .B1(n38164), .B2(n29008), .ZN(
        n29012) );
  XOR2_X1 U29792 ( .A1(n27770), .A2(n27771), .Z(n27772) );
  OAI21_X1 U29795 ( .A1(n21339), .A2(n1693), .B(n7962), .ZN(n6690) );
  XOR2_X1 U29827 ( .A1(n33659), .A2(n16149), .Z(n24421) );
  XOR2_X1 U29836 ( .A1(n12437), .A2(n33515), .Z(n22410) );
  OAI21_X1 U29864 ( .A1(n31549), .A2(n33521), .B(n33520), .ZN(n8231) );
  XOR2_X1 U29871 ( .A1(n25180), .A2(n25198), .Z(n2959) );
  NAND3_X2 U29886 ( .A1(n5895), .A2(n7130), .A3(n31019), .ZN(n33526) );
  XOR2_X1 U29887 ( .A1(n33527), .A2(n9557), .Z(n7492) );
  NOR2_X2 U29913 ( .A1(n13976), .A2(n33528), .ZN(n15540) );
  INV_X1 U29935 ( .I(n30454), .ZN(n33531) );
  OAI21_X2 U29962 ( .A1(n9286), .A2(n9102), .B(n33534), .ZN(n474) );
  XOR2_X1 U30002 ( .A1(n22412), .A2(n22413), .Z(n22946) );
  OAI22_X2 U30003 ( .A1(n7003), .A2(n19599), .B1(n7001), .B2(n7002), .ZN(
        n29756) );
  OAI21_X1 U30007 ( .A1(n33767), .A2(n29756), .B(n33766), .ZN(n29749) );
  OR2_X1 U30010 ( .A1(n22287), .A2(n8519), .Z(n33549) );
  INV_X2 U30011 ( .I(n33550), .ZN(n670) );
  XOR2_X1 U30012 ( .A1(Plaintext[2]), .A2(Key[2]), .Z(n33550) );
  NAND2_X1 U30013 ( .A1(n30959), .A2(n28069), .ZN(n33552) );
  INV_X2 U30015 ( .I(n33553), .ZN(n33957) );
  OAI22_X2 U30018 ( .A1(n124), .A2(n11004), .B1(n12953), .B2(n15320), .ZN(
        n24337) );
  NAND2_X2 U30021 ( .A1(n12206), .A2(n24502), .ZN(n25132) );
  OAI21_X1 U30028 ( .A1(n20147), .A2(n22226), .B(n20643), .ZN(n20146) );
  XOR2_X1 U30042 ( .A1(n26308), .A2(n33566), .Z(n11975) );
  XOR2_X1 U30043 ( .A1(n5690), .A2(n26307), .Z(n33566) );
  XOR2_X1 U30046 ( .A1(n33568), .A2(n21076), .Z(n4856) );
  XOR2_X1 U30047 ( .A1(n29127), .A2(n33569), .Z(n33568) );
  INV_X1 U30048 ( .I(n19908), .ZN(n33569) );
  XOR2_X1 U30051 ( .A1(n10549), .A2(n33572), .Z(n19341) );
  XOR2_X1 U30052 ( .A1(n33573), .A2(n10548), .Z(n33572) );
  XNOR2_X1 U30053 ( .A1(n26551), .A2(n26541), .ZN(n15819) );
  NAND2_X2 U30060 ( .A1(n20969), .A2(n7831), .ZN(n16542) );
  NAND3_X1 U30061 ( .A1(n38156), .A2(n29339), .A3(n1391), .ZN(n20480) );
  NAND2_X2 U30065 ( .A1(n9250), .A2(n9248), .ZN(n29678) );
  XOR2_X1 U30073 ( .A1(n23959), .A2(n17404), .Z(n9446) );
  BUF_X2 U30074 ( .I(n12341), .Z(n33584) );
  OAI21_X1 U30075 ( .A1(n18294), .A2(n5166), .B(n25725), .ZN(n25726) );
  NOR2_X2 U30077 ( .A1(n948), .A2(n12844), .ZN(n8963) );
  XOR2_X1 U30082 ( .A1(n23662), .A2(n7129), .Z(n7128) );
  XOR2_X1 U30086 ( .A1(n28988), .A2(n28989), .Z(n6835) );
  INV_X2 U30090 ( .I(n27932), .ZN(n1072) );
  XOR2_X1 U30091 ( .A1(n11154), .A2(n11152), .Z(n27932) );
  XOR2_X1 U30096 ( .A1(n33595), .A2(n1938), .Z(n1936) );
  NAND2_X1 U30099 ( .A1(n2488), .A2(n2490), .ZN(n2487) );
  OR2_X1 U30101 ( .A1(n30494), .A2(n30833), .Z(n24269) );
  NAND2_X1 U30104 ( .A1(n10314), .A2(n26852), .ZN(n21249) );
  XOR2_X1 U30107 ( .A1(n26585), .A2(n4622), .Z(n10319) );
  INV_X2 U30109 ( .I(n33604), .ZN(n8193) );
  XNOR2_X1 U30110 ( .A1(n11575), .A2(n5600), .ZN(n33604) );
  XOR2_X1 U30113 ( .A1(n3696), .A2(n3695), .Z(n8889) );
  OR2_X1 U30115 ( .A1(n30555), .A2(n38143), .Z(n33608) );
  AOI21_X2 U30117 ( .A1(n33610), .A2(n4665), .B(n28309), .ZN(n2269) );
  OAI21_X1 U30118 ( .A1(n898), .A2(n20577), .B(n33612), .ZN(n33611) );
  XOR2_X1 U30120 ( .A1(n29074), .A2(n33614), .Z(n20325) );
  XOR2_X1 U30121 ( .A1(n29131), .A2(n18430), .Z(n33614) );
  INV_X2 U30130 ( .I(n33621), .ZN(n4603) );
  XOR2_X1 U30131 ( .A1(n22516), .A2(n11793), .Z(n33622) );
  NAND2_X1 U30134 ( .A1(n29175), .A2(n18134), .ZN(n30089) );
  INV_X2 U30137 ( .I(n33625), .ZN(n12478) );
  XNOR2_X1 U30138 ( .A1(n317), .A2(n9094), .ZN(n33625) );
  NAND2_X2 U30141 ( .A1(n15634), .A2(n33628), .ZN(n18062) );
  NAND3_X2 U30142 ( .A1(n37184), .A2(n25503), .A3(n35611), .ZN(n33628) );
  NAND3_X1 U30144 ( .A1(n29365), .A2(n12943), .A3(n37096), .ZN(n29370) );
  INV_X2 U30145 ( .I(n17179), .ZN(n10140) );
  XOR2_X1 U30149 ( .A1(n26433), .A2(n8625), .Z(n33733) );
  XOR2_X1 U30150 ( .A1(n21346), .A2(Key[25]), .Z(n21669) );
  XOR2_X1 U30155 ( .A1(n16689), .A2(n16687), .Z(n22798) );
  XOR2_X1 U30156 ( .A1(n33777), .A2(n19066), .Z(n29456) );
  XOR2_X1 U30158 ( .A1(n33642), .A2(n9159), .Z(n14462) );
  AOI21_X2 U30159 ( .A1(n33643), .A2(n12167), .B(n17383), .ZN(n29659) );
  XOR2_X1 U30161 ( .A1(n14039), .A2(n19035), .Z(n28999) );
  OR2_X1 U30162 ( .A1(n8479), .A2(n2752), .Z(n6137) );
  INV_X2 U30163 ( .I(n25966), .ZN(n26030) );
  NAND2_X2 U30164 ( .A1(n20187), .A2(n20186), .ZN(n25966) );
  NAND2_X2 U30167 ( .A1(n11910), .A2(n17132), .ZN(n27326) );
  NAND2_X2 U30168 ( .A1(n17415), .A2(n17416), .ZN(n12327) );
  XOR2_X1 U30170 ( .A1(n9230), .A2(n12989), .Z(n33650) );
  AOI22_X2 U30173 ( .A1(n30190), .A2(n5414), .B1(n10628), .B2(n30238), .ZN(
        n33651) );
  OAI22_X2 U30174 ( .A1(n11213), .A2(n15237), .B1(n12090), .B2(n13186), .ZN(
        n10931) );
  NAND3_X2 U30179 ( .A1(n7013), .A2(n7012), .A3(n7014), .ZN(n7712) );
  XOR2_X1 U30181 ( .A1(n26387), .A2(n10878), .Z(n33653) );
  XOR2_X1 U30184 ( .A1(n22778), .A2(n22687), .Z(n22546) );
  NOR2_X2 U30187 ( .A1(n29488), .A2(n29489), .ZN(n29535) );
  XOR2_X1 U30191 ( .A1(n23966), .A2(n16153), .Z(n33659) );
  XOR2_X1 U30192 ( .A1(n7152), .A2(n7153), .Z(n25553) );
  XOR2_X1 U30193 ( .A1(n26602), .A2(n33661), .Z(n33660) );
  XOR2_X1 U30195 ( .A1(n32885), .A2(n6634), .Z(n6633) );
  AOI22_X1 U30196 ( .A1(n8062), .A2(n33664), .B1(n8064), .B2(n21147), .ZN(
        n8060) );
  NAND2_X1 U30197 ( .A1(n19348), .A2(n29756), .ZN(n33664) );
  INV_X2 U30198 ( .I(n33665), .ZN(n4879) );
  XOR2_X1 U30199 ( .A1(n5782), .A2(n5781), .Z(n33665) );
  INV_X2 U30200 ( .I(n30249), .ZN(n30260) );
  NAND3_X2 U30210 ( .A1(n33671), .A2(n18101), .A3(n17584), .ZN(n24805) );
  NAND3_X1 U30211 ( .A1(n17586), .A2(n37122), .A3(n19880), .ZN(n33671) );
  OR2_X1 U30220 ( .A1(n12218), .A2(n15038), .Z(n28271) );
  XOR2_X1 U30223 ( .A1(n28850), .A2(n16017), .Z(n29152) );
  XOR2_X1 U30225 ( .A1(n25271), .A2(n25155), .Z(n24948) );
  NOR2_X1 U30229 ( .A1(n1450), .A2(n15357), .ZN(n13053) );
  XOR2_X1 U30234 ( .A1(n19254), .A2(n22598), .Z(n18446) );
  XOR2_X1 U30235 ( .A1(n15673), .A2(n33687), .Z(n15672) );
  XOR2_X1 U30236 ( .A1(n26590), .A2(n19736), .Z(n33687) );
  XOR2_X1 U30237 ( .A1(n16216), .A2(n7854), .Z(n7780) );
  XOR2_X1 U30241 ( .A1(n15824), .A2(n33694), .Z(n33693) );
  NAND2_X2 U30246 ( .A1(n2766), .A2(n25650), .ZN(n18661) );
  XOR2_X1 U30247 ( .A1(n25011), .A2(n13596), .Z(n2896) );
  OAI22_X2 U30248 ( .A1(n37196), .A2(n36564), .B1(n23351), .B2(n32158), .ZN(
        n33696) );
  NAND2_X2 U30255 ( .A1(n19337), .A2(n19395), .ZN(n21545) );
  XOR2_X1 U30262 ( .A1(n26531), .A2(n26341), .Z(n26342) );
  NAND3_X1 U30264 ( .A1(n39425), .A2(n1418), .A3(n37081), .ZN(n12947) );
  NAND2_X2 U30265 ( .A1(n33760), .A2(n21038), .ZN(n29755) );
  XOR2_X1 U30266 ( .A1(n1456), .A2(n27828), .Z(n18662) );
  MUX2_X1 U30269 ( .I0(n36226), .I1(n378), .S(n4604), .Z(n15183) );
  NOR2_X1 U30273 ( .A1(n15880), .A2(n17194), .ZN(n33709) );
  NOR2_X2 U30276 ( .A1(n6977), .A2(n35560), .ZN(n10468) );
  NOR2_X2 U30280 ( .A1(n15981), .A2(n1137), .ZN(n2601) );
  XOR2_X1 U30283 ( .A1(n33716), .A2(n29169), .Z(n29897) );
  NAND2_X2 U30284 ( .A1(n37105), .A2(n12672), .ZN(n24728) );
  XOR2_X1 U30285 ( .A1(n28935), .A2(n33717), .Z(n33965) );
  XOR2_X1 U30286 ( .A1(n28500), .A2(n38195), .Z(n33717) );
  XOR2_X1 U30290 ( .A1(n26194), .A2(n20539), .Z(n33718) );
  XOR2_X1 U30292 ( .A1(n1825), .A2(n11559), .Z(n33722) );
  OAI21_X1 U30298 ( .A1(n35921), .A2(n9942), .B(n33731), .ZN(n21443) );
  XOR2_X1 U30300 ( .A1(n33733), .A2(n8626), .Z(n860) );
  OAI21_X2 U30308 ( .A1(n8175), .A2(n24338), .B(n8174), .ZN(n24339) );
  NAND2_X2 U30310 ( .A1(n33944), .A2(n370), .ZN(n33743) );
  MUX2_X1 U30314 ( .I0(n28555), .I1(n28556), .S(n37758), .Z(n28557) );
  XOR2_X1 U30315 ( .A1(n29130), .A2(n29129), .Z(n29135) );
  XNOR2_X1 U30316 ( .A1(n29121), .A2(n29122), .ZN(n29130) );
  NAND2_X2 U30317 ( .A1(n29600), .A2(n33746), .ZN(n29623) );
  NAND3_X1 U30319 ( .A1(n37213), .A2(n19259), .A3(n26103), .ZN(n26104) );
  XOR2_X1 U30320 ( .A1(n29147), .A2(n15960), .Z(n29086) );
  XOR2_X1 U30321 ( .A1(n33749), .A2(n33751), .Z(n2819) );
  XOR2_X1 U30322 ( .A1(n12145), .A2(n26417), .Z(n5849) );
  XOR2_X1 U30326 ( .A1(n33750), .A2(n3712), .Z(n33749) );
  INV_X1 U30327 ( .I(n24744), .ZN(n33754) );
  XOR2_X1 U30328 ( .A1(n33756), .A2(n22476), .Z(n6329) );
  XOR2_X1 U30331 ( .A1(n12480), .A2(n33757), .Z(n12840) );
  XOR2_X1 U30332 ( .A1(n1621), .A2(n12842), .Z(n33757) );
  XOR2_X1 U30333 ( .A1(n27490), .A2(n1936), .Z(n33758) );
  XOR2_X1 U30334 ( .A1(n33759), .A2(n10070), .Z(n11727) );
  OAI21_X2 U30341 ( .A1(n20330), .A2(n20331), .B(n7601), .ZN(n22067) );
  INV_X1 U30346 ( .I(n6732), .ZN(n11146) );
  BUF_X2 U30349 ( .I(n18047), .Z(n33773) );
  XOR2_X1 U30356 ( .A1(n5382), .A2(n33776), .Z(n855) );
  XOR2_X1 U30357 ( .A1(n12860), .A2(n12859), .Z(n33776) );
  XOR2_X1 U30359 ( .A1(n12736), .A2(n12735), .Z(n12788) );
  NAND2_X2 U30360 ( .A1(n6036), .A2(n22277), .ZN(n22048) );
  XOR2_X1 U30366 ( .A1(n16650), .A2(n494), .Z(n33789) );
  XOR2_X1 U30382 ( .A1(n23783), .A2(n23938), .Z(n8671) );
  NAND2_X2 U30383 ( .A1(n33799), .A2(n27426), .ZN(n13054) );
  NOR2_X1 U30391 ( .A1(n33561), .A2(n26606), .ZN(n33802) );
  XOR2_X1 U30396 ( .A1(n6741), .A2(n4883), .Z(n18209) );
  XOR2_X1 U30398 ( .A1(n38148), .A2(n5261), .Z(n33807) );
  INV_X2 U30399 ( .I(n33808), .ZN(n20793) );
  XOR2_X1 U30410 ( .A1(n727), .A2(n33810), .Z(n354) );
  XOR2_X1 U30411 ( .A1(n8163), .A2(n33811), .Z(n33810) );
  INV_X1 U30412 ( .I(n19735), .ZN(n33811) );
  NOR2_X2 U30414 ( .A1(n33813), .A2(n10832), .ZN(n6885) );
  AOI22_X2 U30422 ( .A1(n8928), .A2(n20978), .B1(n23554), .B2(n35039), .ZN(
        n13617) );
  INV_X4 U30425 ( .I(n18519), .ZN(n33826) );
  XOR2_X1 U30429 ( .A1(n6893), .A2(n20483), .Z(n33824) );
  OAI21_X2 U30430 ( .A1(n19237), .A2(n25557), .B(n33825), .ZN(n25777) );
  XOR2_X1 U30439 ( .A1(n4059), .A2(n4061), .Z(n4300) );
  XOR2_X1 U30447 ( .A1(n18662), .A2(n27832), .Z(n33831) );
  NAND2_X1 U30449 ( .A1(n20743), .A2(n23211), .ZN(n33832) );
  XOR2_X1 U30453 ( .A1(n27552), .A2(n27551), .Z(n33837) );
  XOR2_X1 U30454 ( .A1(n33839), .A2(n36529), .Z(n3257) );
  XOR2_X1 U30455 ( .A1(n3261), .A2(n9184), .Z(n33839) );
  INV_X1 U30456 ( .I(n7194), .ZN(n30230) );
  OAI21_X2 U30460 ( .A1(n2294), .A2(n2378), .B(n29592), .ZN(n33844) );
  BUF_X2 U30464 ( .I(n7090), .Z(n33845) );
  XOR2_X1 U30470 ( .A1(n14264), .A2(n20454), .Z(n9038) );
  XOR2_X1 U30472 ( .A1(n33848), .A2(n3872), .Z(n15754) );
  XOR2_X1 U30475 ( .A1(n11015), .A2(n11016), .Z(n33850) );
  XOR2_X1 U30479 ( .A1(n13102), .A2(n13101), .Z(n33851) );
  NAND2_X1 U30488 ( .A1(n16693), .A2(n19823), .ZN(n19661) );
  NAND2_X2 U30489 ( .A1(n29870), .A2(n10096), .ZN(n29871) );
  OR2_X1 U30490 ( .A1(n15852), .A2(n36661), .Z(n21979) );
  OAI21_X2 U30491 ( .A1(n19320), .A2(n1813), .B(n532), .ZN(n11344) );
  AOI22_X2 U30492 ( .A1(n26728), .A2(n14380), .B1(n26777), .B2(n31982), .ZN(
        n33853) );
  XOR2_X1 U30502 ( .A1(n22594), .A2(n33866), .Z(n33865) );
  XOR2_X1 U30505 ( .A1(n10413), .A2(n3316), .Z(n33868) );
  NAND3_X1 U30506 ( .A1(n1623), .A2(n38535), .A3(n10024), .ZN(n33869) );
  XOR2_X1 U30510 ( .A1(n27526), .A2(n27473), .Z(n33870) );
  INV_X1 U30511 ( .I(n2940), .ZN(n25844) );
  XOR2_X1 U30514 ( .A1(n26399), .A2(n26398), .Z(n7689) );
  NAND2_X2 U30520 ( .A1(n2932), .A2(n30420), .ZN(n23996) );
  INV_X2 U30523 ( .I(n31378), .ZN(n10618) );
  INV_X2 U30526 ( .I(n33890), .ZN(n773) );
  NAND2_X2 U30530 ( .A1(n14080), .A2(n5960), .ZN(n26794) );
  XOR2_X1 U30531 ( .A1(n14563), .A2(n24950), .Z(n3029) );
  NAND2_X2 U30534 ( .A1(n14822), .A2(n21739), .ZN(n7560) );
  XOR2_X1 U30536 ( .A1(n33906), .A2(n1725), .Z(Ciphertext[78]) );
  AOI22_X1 U30537 ( .A1(n17368), .A2(n19318), .B1(n29646), .B2(n29658), .ZN(
        n33906) );
  NAND2_X2 U30539 ( .A1(n6208), .A2(n6206), .ZN(n6205) );
  XOR2_X1 U30547 ( .A1(n5246), .A2(n22562), .Z(n22419) );
  OAI22_X1 U30548 ( .A1(n18070), .A2(n1387), .B1(n29228), .B2(n14933), .ZN(
        n14200) );
  BUF_X2 U30550 ( .I(n16487), .Z(n33916) );
  NAND2_X2 U30569 ( .A1(n25778), .A2(n25776), .ZN(n2830) );
  XOR2_X1 U30572 ( .A1(n11903), .A2(n7573), .Z(n26818) );
  INV_X2 U30577 ( .I(n7273), .ZN(n24142) );
  NOR2_X2 U30579 ( .A1(n5015), .A2(n5014), .ZN(n9276) );
  OAI22_X2 U30583 ( .A1(n16411), .A2(n16810), .B1(n16410), .B2(n16809), .ZN(
        n25962) );
  CLKBUF_X4 U30585 ( .I(n26995), .Z(n19364) );
  XOR2_X1 U30588 ( .A1(n16551), .A2(n16550), .Z(n33954) );
  XOR2_X1 U30590 ( .A1(n13751), .A2(n13749), .Z(n33956) );
  INV_X4 U30591 ( .I(n12685), .ZN(n18246) );
  XNOR2_X1 U30592 ( .A1(n8909), .A2(n29083), .ZN(n33962) );
  INV_X2 U30595 ( .I(n11896), .ZN(n14557) );
  OR2_X2 U30597 ( .A1(n10097), .A2(n18445), .Z(n33966) );
  AND2_X1 U30598 ( .A1(n29721), .A2(n14337), .Z(n33968) );
  INV_X2 U30599 ( .I(n28817), .ZN(n28925) );
  BUF_X2 U3421 ( .I(n12519), .Z(n3226) );
  INV_X2 U15475 ( .I(n3462), .ZN(n8955) );
  INV_X4 U9227 ( .I(n27403), .ZN(n1220) );
  INV_X2 U3911 ( .I(n2561), .ZN(n9175) );
  INV_X4 U5822 ( .I(n18293), .ZN(n917) );
  INV_X2 U5706 ( .I(n24912), .ZN(n1273) );
  OAI21_X2 U12087 ( .A1(n25792), .A2(n25975), .B(n17002), .ZN(n25795) );
  INV_X2 U1188 ( .I(n19580), .ZN(n25835) );
  INV_X2 U6510 ( .I(n15535), .ZN(n968) );
  INV_X2 U16873 ( .I(n3861), .ZN(n2944) );
  NOR2_X2 U10138 ( .A1(n14270), .A2(n4902), .ZN(n9392) );
  INV_X2 U6809 ( .I(n26274), .ZN(n1509) );
  INV_X2 U22777 ( .I(n11048), .ZN(n11890) );
  OAI21_X2 U380 ( .A1(n27959), .A2(n20185), .B(n10721), .ZN(n10720) );
  NAND2_X2 U5871 ( .A1(n17114), .A2(n33405), .ZN(n13500) );
  INV_X2 U25694 ( .I(n13457), .ZN(n21223) );
  NAND2_X2 U5048 ( .A1(n26134), .A2(n25936), .ZN(n26024) );
  AOI21_X2 U1221 ( .A1(n32654), .A2(n10753), .B(n20683), .ZN(n11860) );
  OAI22_X2 U7339 ( .A1(n36764), .A2(n11898), .B1(n2858), .B2(n5579), .ZN(
        n29860) );
  NAND2_X2 U3258 ( .A1(n2625), .A2(n17400), .ZN(n21040) );
  INV_X2 U10896 ( .I(n11406), .ZN(n16252) );
  INV_X2 U23384 ( .I(n19147), .ZN(n12167) );
  NAND2_X2 U16469 ( .A1(n29354), .A2(n12994), .ZN(n12993) );
  INV_X2 U1098 ( .I(n17790), .ZN(n20864) );
  INV_X2 U17113 ( .I(n16692), .ZN(n23071) );
  OAI21_X2 U1040 ( .A1(n9384), .A2(n4475), .B(n1591), .ZN(n9382) );
  INV_X4 U842 ( .I(n16836), .ZN(n953) );
  AOI21_X2 U16551 ( .A1(n24392), .A2(n11265), .B(n12771), .ZN(n15237) );
  INV_X2 U2358 ( .I(n28692), .ZN(n18453) );
  NAND2_X2 U3582 ( .A1(n15176), .A2(n36442), .ZN(n23338) );
  NAND2_X2 U27370 ( .A1(n18838), .A2(n25108), .ZN(n25993) );
  INV_X2 U13068 ( .I(n16524), .ZN(n16368) );
  OAI21_X2 U9696 ( .A1(n24209), .A2(n24207), .B(n24208), .ZN(n18938) );
  INV_X2 U1938 ( .I(n13370), .ZN(n23578) );
  INV_X2 U580 ( .I(n866), .ZN(n26862) );
  NAND2_X2 U5776 ( .A1(n20403), .A2(n9295), .ZN(n9726) );
  NAND2_X1 U15038 ( .A1(n22807), .A2(n23119), .ZN(n31345) );
  NAND2_X2 U1485 ( .A1(n18715), .A2(n24882), .ZN(n25211) );
  INV_X2 U27483 ( .I(n28651), .ZN(n28490) );
  NAND2_X2 U763 ( .A1(n8137), .A2(n27379), .ZN(n27300) );
  INV_X2 U22306 ( .I(n37045), .ZN(n24184) );
  INV_X2 U246 ( .I(n6932), .ZN(n28386) );
  NAND2_X2 U13 ( .A1(n15773), .A2(n29890), .ZN(n29881) );
  OAI21_X2 U1777 ( .A1(n30900), .A2(n31827), .B(n5276), .ZN(n5508) );
  OAI21_X2 U10705 ( .A1(n9818), .A2(n9817), .B(n1056), .ZN(n4916) );
  NOR2_X2 U13467 ( .A1(n22812), .A2(n22811), .ZN(n23587) );
  INV_X4 U2155 ( .I(n5077), .ZN(n31940) );
  BUF_X4 U6320 ( .I(n23761), .Z(n24300) );
  NAND2_X2 U5290 ( .A1(n37319), .A2(n37107), .ZN(n11796) );
  INV_X2 U5569 ( .I(n26403), .ZN(n10491) );
  AOI21_X2 U10669 ( .A1(n3156), .A2(n3155), .B(n3154), .ZN(n3153) );
  OAI21_X2 U2350 ( .A1(n1997), .A2(n7591), .B(n1440), .ZN(n7252) );
  INV_X2 U349 ( .I(n6640), .ZN(n1069) );
  BUF_X4 U3916 ( .I(n33533), .Z(n33178) );
  INV_X2 U300 ( .I(n16067), .ZN(n28485) );
  NAND2_X2 U9745 ( .A1(n24209), .A2(n18937), .ZN(n18936) );
  NAND2_X2 U9838 ( .A1(n3382), .A2(n1629), .ZN(n5186) );
  INV_X2 U3630 ( .I(n26779), .ZN(n26945) );
  INV_X2 U1412 ( .I(n25569), .ZN(n15180) );
  INV_X2 U2047 ( .I(n20679), .ZN(n1341) );
  INV_X2 U991 ( .I(n24864), .ZN(n1030) );
  INV_X2 U2472 ( .I(n36996), .ZN(n23166) );
  INV_X4 U732 ( .I(n16867), .ZN(n10062) );
  AND2_X1 U6294 ( .A1(n35216), .A2(n220), .Z(n30400) );
  INV_X2 U1386 ( .I(n34134), .ZN(n7075) );
  BUF_X4 U1825 ( .I(n14272), .Z(n32190) );
  OAI21_X2 U7190 ( .A1(n18566), .A2(n21451), .B(n18567), .ZN(n21452) );
  AOI21_X2 U14730 ( .A1(n2300), .A2(n21672), .B(n21847), .ZN(n8073) );
  AOI22_X2 U1648 ( .A1(n18376), .A2(n1520), .B1(n31954), .B2(n362), .ZN(n25837) );
  NAND2_X2 U327 ( .A1(n28742), .A2(n5424), .ZN(n16530) );
  NOR2_X2 U448 ( .A1(n11375), .A2(n28159), .ZN(n28287) );
  NAND2_X2 U131 ( .A1(n9708), .A2(n30159), .ZN(n33362) );
  NAND2_X2 U22212 ( .A1(n17329), .A2(n17331), .ZN(n17458) );
  OAI21_X2 U3138 ( .A1(n4225), .A2(n32093), .B(n35952), .ZN(n2164) );
  INV_X4 U1908 ( .I(n10736), .ZN(n946) );
  OAI21_X2 U11661 ( .A1(n23350), .A2(n37523), .B(n30974), .ZN(n23356) );
  NAND2_X2 U12678 ( .A1(n9578), .A2(n9583), .ZN(n15282) );
  NAND3_X2 U30416 ( .A1(n33816), .A2(n10224), .A3(n33815), .ZN(n9499) );
  NOR2_X2 U4514 ( .A1(n24649), .A2(n31796), .ZN(n4845) );
  NAND2_X2 U3141 ( .A1(n24648), .A2(n36340), .ZN(n24649) );
  NOR2_X2 U6036 ( .A1(n15149), .A2(n33771), .ZN(n15148) );
  NAND2_X2 U2777 ( .A1(n30024), .A2(n30038), .ZN(n30015) );
  OAI21_X2 U5927 ( .A1(n27946), .A2(n12406), .B(n20431), .ZN(n33528) );
  BUF_X4 U3921 ( .I(n16692), .Z(n9954) );
  INV_X2 U1141 ( .I(n16296), .ZN(n16342) );
  BUF_X2 U1956 ( .I(n8668), .Z(n605) );
  OAI21_X2 U81 ( .A1(n29302), .A2(n29461), .B(n38051), .ZN(n21195) );
  NAND2_X2 U17554 ( .A1(n33190), .A2(n5287), .ZN(n31591) );
  INV_X2 U3433 ( .I(n21126), .ZN(n18603) );
  INV_X4 U3794 ( .I(n38220), .ZN(n7905) );
  AOI22_X2 U12600 ( .A1(n6229), .A2(n24910), .B1(n12671), .B2(n24909), .ZN(
        n6228) );
  INV_X2 U27338 ( .I(n18739), .ZN(n19091) );
  INV_X2 U15360 ( .I(n3713), .ZN(n17556) );
  NAND2_X2 U8386 ( .A1(n8757), .A2(n33864), .ZN(n23360) );
  AOI21_X2 U9389 ( .A1(n9962), .A2(n9961), .B(n1527), .ZN(n16344) );
  INV_X2 U5654 ( .I(n35543), .ZN(n20578) );
  NAND2_X2 U1551 ( .A1(n8139), .A2(n18654), .ZN(n30929) );
  OAI21_X2 U14862 ( .A1(n1823), .A2(n7555), .B(n28378), .ZN(n20496) );
  NOR2_X2 U6836 ( .A1(n3013), .A2(n35855), .ZN(n26190) );
  NAND2_X2 U2879 ( .A1(n28704), .A2(n38220), .ZN(n28700) );
  INV_X2 U1068 ( .I(n31917), .ZN(n9568) );
  NAND2_X2 U3240 ( .A1(n32338), .A2(n34559), .ZN(n28765) );
  INV_X4 U5561 ( .I(n15575), .ZN(n1021) );
  INV_X2 U12634 ( .I(n24724), .ZN(n6542) );
  NOR3_X1 U3693 ( .A1(n33925), .A2(n36422), .A3(n8809), .ZN(n14879) );
  INV_X4 U10098 ( .I(n23142), .ZN(n1652) );
  NOR2_X2 U7266 ( .A1(n5391), .A2(n36912), .ZN(n5551) );
  NAND2_X2 U2976 ( .A1(n16619), .A2(n11120), .ZN(n28650) );
  OAI21_X1 U7466 ( .A1(n28283), .A2(n27980), .B(n30565), .ZN(n16543) );
  NAND2_X1 U9288 ( .A1(n11968), .A2(n30180), .ZN(n30185) );
  INV_X2 U2099 ( .I(n22066), .ZN(n1673) );
  OAI21_X2 U17989 ( .A1(n30400), .A2(n31660), .B(n38013), .ZN(n31904) );
  INV_X2 U16704 ( .I(n26516), .ZN(n19081) );
  INV_X2 U18292 ( .I(n29532), .ZN(n29517) );
  NOR2_X2 U2657 ( .A1(n19546), .A2(n20923), .ZN(n4373) );
  NOR2_X2 U2703 ( .A1(n34114), .A2(n54), .ZN(n53) );
  AOI21_X2 U4988 ( .A1(n502), .A2(n34128), .B(n36443), .ZN(n32551) );
  NAND2_X2 U11773 ( .A1(n37074), .A2(n106), .ZN(n9239) );
  INV_X4 U7874 ( .I(n1006), .ZN(n3388) );
  INV_X2 U574 ( .I(n10314), .ZN(n20660) );
  NAND3_X2 U22525 ( .A1(n25534), .A2(n25535), .A3(n37795), .ZN(n32911) );
  INV_X2 U1814 ( .I(n33483), .ZN(n802) );
  INV_X2 U6604 ( .I(n28376), .ZN(n28377) );
  AOI21_X2 U13721 ( .A1(n9903), .A2(n22238), .B(n13632), .ZN(n9838) );
  NOR2_X2 U3196 ( .A1(n35580), .A2(n26354), .ZN(n14521) );
  OAI21_X2 U407 ( .A1(n19456), .A2(n16127), .B(n20561), .ZN(n27061) );
  BUF_X4 U7168 ( .I(n14395), .Z(n14396) );
  INV_X2 U542 ( .I(n31682), .ZN(n14480) );
  NAND2_X2 U17177 ( .A1(n38448), .A2(n1049), .ZN(n21983) );
  NAND2_X2 U1997 ( .A1(n23099), .A2(n13650), .ZN(n8337) );
  NAND2_X2 U12502 ( .A1(n2848), .A2(n2847), .ZN(n10646) );
  NAND2_X2 U2064 ( .A1(n12079), .A2(n22131), .ZN(n13615) );
  NOR2_X2 U252 ( .A1(n33424), .A2(n36165), .ZN(n14398) );
  NAND2_X2 U435 ( .A1(n33957), .A2(n10817), .ZN(n30959) );
  NOR2_X2 U119 ( .A1(n39322), .A2(n18667), .ZN(n14773) );
  INV_X2 U4989 ( .I(n9987), .ZN(n21001) );
  NAND3_X2 U5695 ( .A1(n18115), .A2(n24161), .A3(n13128), .ZN(n11768) );
  NOR2_X2 U337 ( .A1(n1190), .A2(n14209), .ZN(n2822) );
  INV_X4 U3109 ( .I(n14553), .ZN(n1108) );
  INV_X2 U3859 ( .I(n5888), .ZN(n355) );
  INV_X2 U8441 ( .I(n18762), .ZN(n20620) );
  OAI21_X1 U9367 ( .A1(n13971), .A2(n26000), .B(n2310), .ZN(n13387) );
  NAND2_X1 U5520 ( .A1(n2311), .A2(n25998), .ZN(n2310) );
  INV_X2 U24518 ( .I(n36728), .ZN(n21950) );
  NAND2_X2 U14186 ( .A1(n34485), .A2(n15677), .ZN(n21266) );
  OAI21_X1 U21593 ( .A1(n10345), .A2(n21783), .B(n21504), .ZN(n32319) );
  NAND2_X2 U16969 ( .A1(n4508), .A2(n4506), .ZN(n6932) );
  OAI21_X2 U16548 ( .A1(n14680), .A2(n15449), .B(n1018), .ZN(n25707) );
  OAI21_X2 U2158 ( .A1(n18372), .A2(n35822), .B(n6200), .ZN(n6199) );
  AOI21_X2 U12383 ( .A1(n30366), .A2(n21223), .B(n15087), .ZN(n31042) );
  INV_X4 U863 ( .I(n37051), .ZN(n1024) );
  INV_X2 U3797 ( .I(n17813), .ZN(n22055) );
  NAND2_X2 U1875 ( .A1(n32260), .A2(n23569), .ZN(n23365) );
  NOR2_X2 U21830 ( .A1(n22330), .A2(n22329), .ZN(n22671) );
  NAND2_X2 U4193 ( .A1(n13044), .A2(n19483), .ZN(n439) );
  NAND2_X1 U27166 ( .A1(n18214), .A2(n1015), .ZN(n18213) );
  INV_X2 U2427 ( .I(n13794), .ZN(n29384) );
  BUF_X2 U13970 ( .I(n21352), .Z(n21683) );
  AOI21_X2 U10685 ( .A1(n29991), .A2(n29992), .B(n29990), .ZN(n9233) );
  INV_X2 U26348 ( .I(n33980), .ZN(n28115) );
  NAND2_X2 U10350 ( .A1(n21920), .A2(n19323), .ZN(n7587) );
  INV_X2 U5772 ( .I(n22671), .ZN(n1662) );
  INV_X2 U23299 ( .I(n12012), .ZN(n20936) );
  OAI21_X2 U1273 ( .A1(n17930), .A2(n39518), .B(n39500), .ZN(n17929) );
  INV_X2 U16271 ( .I(n24637), .ZN(n11712) );
  NAND2_X2 U12302 ( .A1(n17271), .A2(n12500), .ZN(n14300) );
  NOR2_X2 U5409 ( .A1(n33042), .A2(n2731), .ZN(n16541) );
  NAND2_X2 U1872 ( .A1(n1301), .A2(n35915), .ZN(n2084) );
  INV_X4 U9732 ( .I(n17810), .ZN(n8041) );
  INV_X2 U5734 ( .I(n16271), .ZN(n18302) );
  OR2_X2 U17205 ( .A1(n24280), .A2(n19959), .Z(n24284) );
  NOR2_X2 U966 ( .A1(n13588), .A2(n14065), .ZN(n32948) );
  INV_X2 U29 ( .I(n29747), .ZN(n29739) );
  NAND2_X2 U9180 ( .A1(n26965), .A2(n27507), .ZN(n11462) );
  INV_X4 U1636 ( .I(n37097), .ZN(n20158) );
  BUF_X4 U4415 ( .I(n13543), .Z(n13393) );
  INV_X2 U582 ( .I(n26863), .ZN(n1089) );
  AOI21_X2 U6091 ( .A1(n14592), .A2(n39745), .B(n17633), .ZN(n6920) );
  INV_X2 U7080 ( .I(n13150), .ZN(n13831) );
  OAI21_X2 U9379 ( .A1(n26190), .A2(n32243), .B(n39507), .ZN(n19573) );
  AOI21_X2 U1556 ( .A1(n25674), .A2(n19589), .B(n6592), .ZN(n18058) );
  INV_X2 U5999 ( .I(n19692), .ZN(n16104) );
  OAI21_X2 U10329 ( .A1(n21423), .A2(n21667), .B(n21672), .ZN(n21424) );
  NAND2_X1 U978 ( .A1(n5389), .A2(n24852), .ZN(n199) );
  NAND2_X2 U6077 ( .A1(n13441), .A2(n29586), .ZN(n28864) );
  NAND2_X1 U11765 ( .A1(n3103), .A2(n30983), .ZN(n3102) );
  INV_X2 U4913 ( .I(n2008), .ZN(n2405) );
  AOI21_X2 U10314 ( .A1(n13956), .A2(n13044), .B(n18496), .ZN(n11174) );
  BUF_X2 U3027 ( .I(n32165), .Z(n138) );
  NAND2_X1 U5870 ( .A1(n28048), .A2(n28260), .ZN(n4975) );
  OAI21_X2 U8490 ( .A1(n1652), .A2(n1313), .B(n3906), .ZN(n8766) );
  NAND2_X2 U6043 ( .A1(n9863), .A2(n39495), .ZN(n13044) );
  INV_X4 U1378 ( .I(n2576), .ZN(n33114) );
  OAI21_X2 U13858 ( .A1(n21920), .A2(n21621), .B(n7587), .ZN(n6800) );
  NOR2_X2 U5593 ( .A1(n25934), .A2(n38185), .ZN(n25800) );
  NAND2_X2 U27627 ( .A1(n25556), .A2(n1537), .ZN(n20236) );
  AOI22_X2 U10365 ( .A1(n21455), .A2(n21695), .B1(n21454), .B2(n19395), .ZN(
        n13788) );
  NAND2_X2 U2774 ( .A1(n22891), .A2(n5838), .ZN(n70) );
  NAND2_X2 U5761 ( .A1(n33745), .A2(n31093), .ZN(n17968) );
  OAI21_X1 U10292 ( .A1(n15436), .A2(n15493), .B(n15435), .ZN(n30818) );
  NAND2_X2 U3829 ( .A1(n21101), .A2(n34001), .ZN(n27272) );
  NOR2_X2 U17108 ( .A1(n22264), .A2(n33738), .ZN(n14249) );
  INV_X2 U15764 ( .I(n39680), .ZN(n3294) );
  INV_X2 U1101 ( .I(n19341), .ZN(n16449) );
  BUF_X2 U2929 ( .I(n4392), .Z(n33861) );
  BUF_X4 U13968 ( .I(n21358), .Z(n21666) );
  INV_X2 U5392 ( .I(n24713), .ZN(n15193) );
  NOR2_X1 U6748 ( .A1(n26772), .A2(n18225), .ZN(n3103) );
  NAND2_X2 U4604 ( .A1(n10168), .A2(n25751), .ZN(n26014) );
  INV_X2 U27443 ( .I(n19016), .ZN(n19609) );
  INV_X1 U15765 ( .I(n39680), .ZN(n3670) );
  INV_X2 U1161 ( .I(n6302), .ZN(n32497) );
  INV_X1 U6001 ( .I(n22925), .ZN(n23058) );
  INV_X2 U24711 ( .I(n22137), .ZN(n16283) );
  NAND2_X2 U4892 ( .A1(n18417), .A2(n21712), .ZN(n21747) );
  INV_X2 U7184 ( .I(n22491), .ZN(n22025) );
  OAI22_X2 U25396 ( .A1(n2008), .A2(n21924), .B1(n11852), .B2(n9316), .ZN(
        n4913) );
  OAI22_X2 U19016 ( .A1(n1156), .A2(n21853), .B1(n1355), .B2(n21808), .ZN(
        n6271) );
  OAI21_X1 U201 ( .A1(n32274), .A2(n13508), .B(n32273), .ZN(n11536) );
  INV_X4 U27174 ( .I(n23089), .ZN(n23169) );
  NOR2_X2 U7996 ( .A1(n15021), .A2(n25898), .ZN(n10475) );
  INV_X4 U9771 ( .I(n24359), .ZN(n3685) );
  NOR2_X2 U6834 ( .A1(n34577), .A2(n26001), .ZN(n25898) );
  OAI21_X2 U1178 ( .A1(n23611), .A2(n4525), .B(n4527), .ZN(n4526) );
  NOR2_X2 U26636 ( .A1(n21266), .A2(n30900), .ZN(n16903) );
  OAI21_X2 U7724 ( .A1(n1442), .A2(n886), .B(n5239), .ZN(n7945) );
  INV_X4 U5825 ( .I(n7982), .ZN(n21339) );
  NOR2_X2 U2563 ( .A1(n13), .A2(n12), .ZN(n18454) );
  NAND2_X2 U8083 ( .A1(n7853), .A2(n38178), .ZN(n16373) );
  AOI21_X2 U1489 ( .A1(n18339), .A2(n20367), .B(n21950), .ZN(n18338) );
  INV_X4 U1659 ( .I(n17501), .ZN(n17502) );
  NAND2_X2 U5760 ( .A1(n7494), .A2(n27259), .ZN(n8411) );
  NAND2_X2 U10031 ( .A1(n121), .A2(n33045), .ZN(n23024) );
  OAI21_X2 U1621 ( .A1(n22246), .A2(n33571), .B(n37938), .ZN(n22247) );
  INV_X2 U11387 ( .I(n18148), .ZN(n24608) );
  INV_X2 U719 ( .I(n2830), .ZN(n26101) );
  INV_X2 U3742 ( .I(n36549), .ZN(n26866) );
  INV_X2 U865 ( .I(n733), .ZN(n25690) );
  NOR2_X2 U13656 ( .A1(n9838), .A2(n13633), .ZN(n13631) );
  OAI21_X2 U1530 ( .A1(n34040), .A2(n32761), .B(n31796), .ZN(n471) );
  OAI21_X2 U3792 ( .A1(n30475), .A2(n30712), .B(n27189), .ZN(n31421) );
  AOI21_X2 U9873 ( .A1(n10709), .A2(n35963), .B(n38894), .ZN(n10708) );
  AOI22_X2 U7390 ( .A1(n2907), .A2(n30558), .B1(n2909), .B2(n2910), .ZN(n8649)
         );
  NOR2_X2 U4055 ( .A1(n6864), .A2(n8892), .ZN(n29272) );
  NAND2_X2 U12347 ( .A1(n11589), .A2(n33268), .ZN(n4018) );
  INV_X4 U21346 ( .I(n7536), .ZN(n8971) );
  AOI22_X2 U17344 ( .A1(n22103), .A2(n20234), .B1(n22102), .B2(n22335), .ZN(
        n22104) );
  INV_X4 U18946 ( .I(n27153), .ZN(n5311) );
  NAND2_X1 U12109 ( .A1(n3837), .A2(n30629), .ZN(n11269) );
  INV_X4 U6042 ( .I(n19587), .ZN(n5391) );
  NAND2_X2 U13644 ( .A1(n15347), .A2(n36443), .ZN(n2587) );
  INV_X2 U19288 ( .I(n6581), .ZN(n19588) );
  INV_X2 U17467 ( .I(n8293), .ZN(n21692) );
  INV_X2 U5739 ( .I(n23623), .ZN(n23780) );
  NOR2_X2 U3314 ( .A1(n7485), .A2(n33747), .ZN(n23576) );
  NOR2_X1 U7262 ( .A1(n7962), .A2(n9964), .ZN(n5601) );
  INV_X2 U4665 ( .I(n15738), .ZN(n20321) );
  NAND2_X2 U336 ( .A1(n18144), .A2(n11136), .ZN(n28180) );
  OAI21_X2 U3963 ( .A1(n5215), .A2(n5214), .B(n36453), .ZN(n9504) );
  OAI21_X2 U2624 ( .A1(n16395), .A2(n16394), .B(n31331), .ZN(n16393) );
  INV_X4 U7155 ( .I(n23107), .ZN(n20782) );
  BUF_X2 U9578 ( .I(n25488), .Z(n6696) );
  NOR2_X2 U20510 ( .A1(n18174), .A2(n455), .ZN(n14541) );
  INV_X2 U6753 ( .I(n26269), .ZN(n26696) );
  AOI22_X2 U10185 ( .A1(n20374), .A2(n36245), .B1(n20375), .B2(n1154), .ZN(
        n9125) );
  NAND2_X2 U2071 ( .A1(n14027), .A2(n36428), .ZN(n31458) );
  OAI21_X2 U10170 ( .A1(n4110), .A2(n1681), .B(n6361), .ZN(n4109) );
  AOI22_X2 U3404 ( .A1(n16484), .A2(n23468), .B1(n21019), .B2(n32858), .ZN(
        n3194) );
  OR3_X2 U13961 ( .A1(n19549), .A2(n21870), .A3(n3562), .Z(n17665) );
  NAND2_X2 U1842 ( .A1(n18478), .A2(n23635), .ZN(n3195) );
  AND2_X2 U8549 ( .A1(n23080), .A2(n10962), .Z(n1824) );
  NAND2_X1 U7976 ( .A1(n8295), .A2(n34417), .ZN(n8294) );
  NAND2_X1 U14793 ( .A1(n9404), .A2(n13880), .ZN(n31313) );
  NAND2_X2 U6044 ( .A1(n21928), .A2(n19372), .ZN(n21727) );
  INV_X2 U27637 ( .I(n35290), .ZN(n33288) );
  OR2_X1 U4841 ( .A1(n22035), .A2(n35290), .Z(n20388) );
  INV_X2 U25129 ( .I(n23468), .ZN(n21019) );
  INV_X2 U15832 ( .I(n30897), .ZN(n6839) );
  AOI21_X2 U699 ( .A1(n8384), .A2(n26807), .B(n8382), .ZN(n8381) );
  AOI22_X2 U14590 ( .A1(n21379), .A2(n9102), .B1(n11703), .B2(n1346), .ZN(
        n5930) );
  AOI21_X2 U15138 ( .A1(n34016), .A2(n587), .B(n2690), .ZN(n21379) );
  AOI21_X2 U5246 ( .A1(n15462), .A2(n34823), .B(n9835), .ZN(n11560) );
  NAND2_X2 U6245 ( .A1(n5519), .A2(n14436), .ZN(n5672) );
  AOI21_X2 U408 ( .A1(n34387), .A2(n8642), .B(n1474), .ZN(n8641) );
  INV_X2 U16972 ( .I(n19891), .ZN(n28131) );
  INV_X2 U8655 ( .I(n22497), .ZN(n1154) );
  NAND2_X2 U534 ( .A1(n26708), .A2(n17034), .ZN(n15825) );
  BUF_X4 U2723 ( .I(n27392), .Z(n14881) );
  NAND2_X2 U3439 ( .A1(n7512), .A2(n33879), .ZN(n25799) );
  NAND2_X2 U13689 ( .A1(n7578), .A2(n22296), .ZN(n11144) );
  NAND2_X2 U409 ( .A1(n5239), .A2(n5352), .ZN(n7719) );
  INV_X1 U13056 ( .I(n12973), .ZN(n4563) );
  OAI21_X2 U1577 ( .A1(n933), .A2(n1271), .B(n13221), .ZN(n13220) );
  NOR2_X2 U6151 ( .A1(n34360), .A2(n37075), .ZN(n8383) );
  INV_X2 U5834 ( .I(n29720), .ZN(n29708) );
  BUF_X2 U10399 ( .I(n21937), .Z(n19375) );
  NOR2_X2 U17659 ( .A1(n3158), .A2(n3159), .ZN(n33292) );
  NAND2_X2 U1847 ( .A1(n23334), .A2(n23635), .ZN(n32573) );
  NAND2_X1 U8267 ( .A1(n12809), .A2(n12808), .ZN(n31094) );
  AOI21_X2 U10162 ( .A1(n14622), .A2(n22229), .B(n22230), .ZN(n20551) );
  OAI21_X1 U3346 ( .A1(n14100), .A2(n25727), .B(n19678), .ZN(n17740) );
  INV_X2 U836 ( .I(n37048), .ZN(n25337) );
  AOI21_X2 U12666 ( .A1(n18468), .A2(n15333), .B(n19630), .ZN(n7610) );
  NOR3_X2 U22344 ( .A1(n32938), .A2(n32937), .A3(n34044), .ZN(n32483) );
  AOI21_X2 U15178 ( .A1(n12407), .A2(n16547), .B(n2730), .ZN(n3253) );
  NAND2_X2 U1977 ( .A1(n14343), .A2(n14188), .ZN(n19168) );
  AOI22_X2 U4855 ( .A1(n21637), .A2(n21636), .B1(n21942), .B2(n19133), .ZN(
        n33389) );
  INV_X2 U20145 ( .I(n24733), .ZN(n24841) );
  INV_X2 U1505 ( .I(n16897), .ZN(n33400) );
  INV_X2 U2799 ( .I(n7225), .ZN(n15122) );
  NOR2_X1 U10686 ( .A1(n7363), .A2(n6372), .ZN(n10943) );
  INV_X1 U11710 ( .I(n19203), .ZN(n1471) );
  OAI21_X2 U16708 ( .A1(n18063), .A2(n24862), .B(n31684), .ZN(n4227) );
  NOR2_X1 U11109 ( .A1(n24424), .A2(n7658), .ZN(n7657) );
  AOI22_X2 U28579 ( .A1(n33196), .A2(n20782), .B1(n22982), .B2(n23111), .ZN(
        n22983) );
  INV_X2 U2460 ( .I(n6314), .ZN(n16580) );
  INV_X4 U16437 ( .I(n26837), .ZN(n20211) );
  NAND3_X2 U30293 ( .A1(n33724), .A2(n19591), .A3(n32014), .ZN(n16473) );
  OAI22_X2 U17082 ( .A1(n2746), .A2(n37202), .B1(n16541), .B2(n2745), .ZN(
        n16539) );
  NOR2_X2 U1046 ( .A1(n3228), .A2(n3227), .ZN(n10798) );
  CLKBUF_X2 U6464 ( .I(Key[164]), .Z(n29363) );
  INV_X2 U6439 ( .I(n10212), .ZN(n10211) );
  INV_X4 U4632 ( .I(n11710), .ZN(n19630) );
  NAND2_X2 U16536 ( .A1(n20634), .A2(n26219), .ZN(n13156) );
  AOI21_X2 U1458 ( .A1(n21936), .A2(n21935), .B(n21934), .ZN(n22130) );
  INV_X4 U26980 ( .I(n23567), .ZN(n15981) );
  NAND3_X2 U11225 ( .A1(n17647), .A2(n13955), .A3(n28276), .ZN(n11005) );
  OAI21_X2 U6956 ( .A1(n30528), .A2(n1490), .B(n26670), .ZN(n18879) );
  AOI22_X2 U6957 ( .A1(n19331), .A2(n26972), .B1(n32427), .B2(n5935), .ZN(
        n30528) );
  AOI21_X2 U12225 ( .A1(n15355), .A2(n8907), .B(n8905), .ZN(n16879) );
  INV_X1 U8543 ( .I(n8943), .ZN(n15911) );
  AOI22_X2 U3839 ( .A1(n5555), .A2(n12952), .B1(n23035), .B2(n7575), .ZN(n4972) );
  NOR2_X2 U2581 ( .A1(n26014), .A2(n26013), .ZN(n7517) );
  INV_X2 U249 ( .I(n16303), .ZN(n28756) );
  INV_X1 U6498 ( .I(n12952), .ZN(n14402) );
  INV_X4 U2338 ( .I(n29595), .ZN(n31667) );
  CLKBUF_X4 U9821 ( .I(n24318), .Z(n19566) );
  INV_X2 U5069 ( .I(n27884), .ZN(n28256) );
  OAI21_X2 U24679 ( .A1(n13081), .A2(n1437), .B(n28274), .ZN(n17647) );
  INV_X2 U7588 ( .I(n28659), .ZN(n28427) );
  NAND2_X2 U8366 ( .A1(n2087), .A2(n9011), .ZN(n2086) );
  INV_X2 U965 ( .I(n37235), .ZN(n6606) );
  NAND2_X2 U25997 ( .A1(n31595), .A2(n36166), .ZN(n30058) );
  OAI21_X2 U1038 ( .A1(n12984), .A2(n25989), .B(n30571), .ZN(n11423) );
  INV_X4 U17505 ( .I(n29885), .ZN(n15773) );
  NOR2_X2 U3676 ( .A1(n17013), .A2(n25410), .ZN(n9788) );
  INV_X2 U21744 ( .I(n3120), .ZN(n24592) );
  AOI21_X2 U18479 ( .A1(n23470), .A2(n1292), .B(n1310), .ZN(n15564) );
  NAND2_X2 U16639 ( .A1(n27370), .A2(n27369), .ZN(n32332) );
  AOI21_X2 U11586 ( .A1(n27366), .A2(n27364), .B(n16482), .ZN(n27370) );
  INV_X4 U2964 ( .I(n12430), .ZN(n29260) );
  NAND2_X2 U4361 ( .A1(n26822), .A2(n26823), .ZN(n4098) );
  NAND2_X1 U16237 ( .A1(n3723), .A2(n39418), .ZN(n3722) );
  NAND2_X1 U12614 ( .A1(n7806), .A2(n5167), .ZN(n7805) );
  INV_X2 U874 ( .I(n18966), .ZN(n25487) );
  AOI21_X2 U7072 ( .A1(n23493), .A2(n35130), .B(n23315), .ZN(n14129) );
  OAI22_X2 U29965 ( .A1(n5597), .A2(n25517), .B1(n5596), .B2(n25620), .ZN(
        n33535) );
  INV_X4 U15045 ( .I(n2597), .ZN(n10220) );
  BUF_X2 U5824 ( .I(n21927), .Z(n19372) );
  BUF_X4 U10279 ( .I(n18711), .Z(n9265) );
  OAI21_X2 U15546 ( .A1(n3377), .A2(n29793), .B(n36096), .ZN(n9456) );
  NAND2_X2 U24755 ( .A1(n1354), .A2(n18028), .ZN(n18026) );
  NOR2_X2 U5601 ( .A1(n33995), .A2(n39020), .ZN(n3389) );
  NAND2_X2 U13431 ( .A1(n8337), .A2(n11582), .ZN(n18499) );
  OAI21_X2 U22608 ( .A1(n18193), .A2(n2348), .B(n10747), .ZN(n24341) );
  INV_X4 U4384 ( .I(n20404), .ZN(n1593) );
  NAND2_X2 U9425 ( .A1(n2625), .A2(n6056), .ZN(n7292) );
  INV_X2 U3164 ( .I(n4209), .ZN(n22757) );
  INV_X2 U18075 ( .I(n18467), .ZN(n6604) );
  NAND2_X1 U14091 ( .A1(n17323), .A2(n1002), .ZN(n20575) );
  INV_X2 U1213 ( .I(n6263), .ZN(n23552) );
  NAND2_X2 U3303 ( .A1(n17989), .A2(n22310), .ZN(n22051) );
  BUF_X2 U4619 ( .I(n24694), .Z(n32398) );
  BUF_X2 U10103 ( .I(n23202), .Z(n2350) );
  INV_X4 U12942 ( .I(n35960), .ZN(n20411) );
  OAI21_X2 U5321 ( .A1(n7949), .A2(n24119), .B(n232), .ZN(n5853) );
  INV_X2 U647 ( .I(n38149), .ZN(n26568) );
  INV_X4 U1788 ( .I(n24432), .ZN(n1608) );
  NAND2_X1 U21795 ( .A1(n14876), .A2(n22804), .ZN(n14875) );
  INV_X4 U790 ( .I(n17029), .ZN(n19095) );
  NAND2_X2 U710 ( .A1(n9633), .A2(n27253), .ZN(n31716) );
  NAND2_X2 U5718 ( .A1(n12360), .A2(n13555), .ZN(n24098) );
  OAI21_X1 U12644 ( .A1(n957), .A2(n31845), .B(n10403), .ZN(n23858) );
  INV_X2 U1440 ( .I(n2696), .ZN(n18360) );
  INV_X1 U24648 ( .I(n26740), .ZN(n17786) );
  INV_X2 U5899 ( .I(n15371), .ZN(n1489) );
  BUF_X2 U3300 ( .I(n27919), .Z(n28079) );
  OAI21_X2 U8666 ( .A1(n6381), .A2(n21766), .B(n9759), .ZN(n5006) );
  NAND2_X2 U2579 ( .A1(n31038), .A2(n18809), .ZN(n6075) );
  OAI22_X2 U3642 ( .A1(n2451), .A2(n37289), .B1(n10479), .B2(n12373), .ZN(
        n31038) );
  INV_X2 U12240 ( .I(n19240), .ZN(n1522) );
  NAND2_X2 U9919 ( .A1(n14845), .A2(n35192), .ZN(n17521) );
  INV_X2 U1109 ( .I(n94), .ZN(n24235) );
  NAND2_X1 U8246 ( .A1(n11609), .A2(n5224), .ZN(n5223) );
  AOI21_X2 U23573 ( .A1(n13626), .A2(n34920), .B(n12628), .ZN(n13571) );
  INV_X1 U4950 ( .I(n4472), .ZN(n1312) );
  NOR2_X2 U6022 ( .A1(n22196), .A2(n38976), .ZN(n22286) );
  INV_X1 U2239 ( .I(n14784), .ZN(n6960) );
  INV_X2 U7179 ( .I(n14381), .ZN(n1046) );
  INV_X2 U7738 ( .I(n5350), .ZN(n5352) );
  NAND2_X2 U10250 ( .A1(n18360), .A2(n36006), .ZN(n5693) );
  BUF_X2 U2833 ( .I(n26795), .Z(n106) );
  AOI21_X2 U2337 ( .A1(n9688), .A2(n32352), .B(n17085), .ZN(n3945) );
  AOI21_X2 U3593 ( .A1(n5908), .A2(n35059), .B(n26039), .ZN(n9882) );
  AOI21_X2 U8454 ( .A1(n4890), .A2(n22905), .B(n23045), .ZN(n22906) );
  NAND2_X1 U9710 ( .A1(n24132), .A2(n39309), .ZN(n17259) );
  INV_X1 U5365 ( .I(n20891), .ZN(n26786) );
  OAI21_X2 U10778 ( .A1(n11410), .A2(n11409), .B(n17225), .ZN(n13134) );
  BUF_X4 U3306 ( .I(n13904), .Z(n13555) );
  AOI22_X2 U2127 ( .A1(n1340), .A2(n32478), .B1(n4200), .B2(n17499), .ZN(n7107) );
  NAND2_X2 U4362 ( .A1(n12162), .A2(n18519), .ZN(n13218) );
  OAI21_X2 U7774 ( .A1(n27115), .A2(n19334), .B(n9633), .ZN(n12744) );
  NOR2_X2 U18780 ( .A1(n9347), .A2(n9349), .ZN(n9344) );
  INV_X4 U22282 ( .I(n36422), .ZN(n14994) );
  INV_X4 U23214 ( .I(n11823), .ZN(n16576) );
  OAI21_X2 U12591 ( .A1(n12518), .A2(n37421), .B(n9826), .ZN(n24438) );
  INV_X2 U11544 ( .I(n27570), .ZN(n1468) );
  INV_X2 U25460 ( .I(n2348), .ZN(n24326) );
  NAND2_X1 U4226 ( .A1(n30991), .A2(n7409), .ZN(n27967) );
  INV_X2 U23288 ( .I(n32776), .ZN(n17580) );
  OAI21_X2 U12662 ( .A1(n18744), .A2(n35049), .B(n19643), .ZN(n15554) );
  INV_X4 U4292 ( .I(n28114), .ZN(n28249) );
  BUF_X2 U6407 ( .I(n33678), .Z(n2458) );
  AOI21_X2 U10041 ( .A1(n3119), .A2(n23110), .B(n33196), .ZN(n12121) );
  INV_X2 U27912 ( .I(n34013), .ZN(n23174) );
  INV_X2 U5777 ( .I(n32135), .ZN(n18568) );
  NOR2_X2 U2981 ( .A1(n27081), .A2(n35750), .ZN(n27163) );
  AOI21_X2 U1177 ( .A1(n23748), .A2(n13752), .B(n10763), .ZN(n6911) );
  NOR2_X2 U17298 ( .A1(n29426), .A2(n29454), .ZN(n29482) );
  OAI22_X2 U7144 ( .A1(n12123), .A2(n19697), .B1(n1142), .B2(n20230), .ZN(
        n12122) );
  OAI22_X2 U2537 ( .A1(n28525), .A2(n28736), .B1(n8050), .B2(n28735), .ZN(
        n19354) );
  INV_X2 U10095 ( .I(n22921), .ZN(n5838) );
  NAND2_X2 U5024 ( .A1(n9321), .A2(n23548), .ZN(n23229) );
  INV_X2 U26974 ( .I(n39830), .ZN(n29704) );
  NAND4_X2 U22555 ( .A1(n11065), .A2(n11064), .A3(n17331), .A4(n17329), .ZN(
        n25959) );
  INV_X2 U25909 ( .I(n33029), .ZN(n33952) );
  NAND2_X1 U4797 ( .A1(n20790), .A2(n35282), .ZN(n583) );
  BUF_X4 U18711 ( .I(n15426), .Z(n31796) );
  AOI21_X2 U1947 ( .A1(n35689), .A2(n30506), .B(n21130), .ZN(n15940) );
  NAND2_X2 U25817 ( .A1(n22344), .A2(n15350), .ZN(n21984) );
  AOI21_X2 U1306 ( .A1(n33826), .A2(n25557), .B(n19367), .ZN(n33825) );
  INV_X4 U3186 ( .I(n21822), .ZN(n18174) );
  INV_X2 U12014 ( .I(n31791), .ZN(n1879) );
  OAI22_X2 U13139 ( .A1(n5759), .A2(n23017), .B1(n8692), .B2(n9078), .ZN(
        n23019) );
  NAND2_X2 U21871 ( .A1(n11144), .A2(n22248), .ZN(n11143) );
  BUF_X2 U11568 ( .I(n7611), .Z(n4964) );
  AND2_X1 U3599 ( .A1(n27385), .A2(n18549), .Z(n5220) );
  INV_X4 U30384 ( .I(n9876), .ZN(n22344) );
  INV_X1 U18791 ( .I(n17464), .ZN(n18679) );
  INV_X2 U17549 ( .I(n17775), .ZN(n32441) );
  INV_X2 U5850 ( .I(n16116), .ZN(n29494) );
  OAI22_X2 U2595 ( .A1(n5669), .A2(n33081), .B1(n32777), .B2(n31788), .ZN(
        n30239) );
  OAI22_X2 U16617 ( .A1(n6720), .A2(n15773), .B1(n967), .B2(n38217), .ZN(
        n29889) );
  NOR2_X2 U44 ( .A1(n33813), .A2(n10832), .ZN(n31533) );
  AOI21_X2 U28432 ( .A1(n22345), .A2(n22344), .B(n22343), .ZN(n22346) );
  INV_X2 U21082 ( .I(n8544), .ZN(n9677) );
  INV_X2 U8721 ( .I(n21872), .ZN(n21695) );
  INV_X2 U5043 ( .I(n10705), .ZN(n22541) );
  NOR2_X2 U25106 ( .A1(n36227), .A2(n35685), .ZN(n16027) );
  INV_X2 U6444 ( .I(n21740), .ZN(n21748) );
  INV_X4 U8434 ( .I(n31931), .ZN(n1301) );
  OR2_X1 U2183 ( .A1(n21822), .A2(n19016), .Z(n21678) );
  INV_X4 U16378 ( .I(n31511), .ZN(n29587) );
  INV_X2 U13050 ( .I(n24318), .ZN(n18348) );
  NAND2_X2 U26149 ( .A1(n27959), .A2(n37671), .ZN(n18036) );
  NOR2_X2 U6149 ( .A1(n38900), .A2(n37075), .ZN(n27560) );
  AOI21_X2 U2032 ( .A1(n24390), .A2(n14292), .B(n14291), .ZN(n16068) );
  INV_X2 U10255 ( .I(n22223), .ZN(n22165) );
  NAND2_X1 U24504 ( .A1(n9670), .A2(n21576), .ZN(n20588) );
  AOI21_X2 U26286 ( .A1(n30306), .A2(n17685), .B(n22067), .ZN(n22068) );
  NAND3_X2 U651 ( .A1(n36528), .A2(n27244), .A3(n991), .ZN(n30678) );
  INV_X2 U4578 ( .I(n1326), .ZN(n8679) );
  INV_X2 U12763 ( .I(n19294), .ZN(n24811) );
  AOI21_X2 U22330 ( .A1(n937), .A2(n10242), .B(n17723), .ZN(n22127) );
  OAI21_X2 U9744 ( .A1(n24251), .A2(n24466), .B(n33379), .ZN(n13264) );
  AOI21_X2 U30004 ( .A1(n21482), .A2(n21483), .B(n5751), .ZN(n14125) );
  NAND2_X2 U1414 ( .A1(n7916), .A2(n22239), .ZN(n9903) );
  INV_X4 U2478 ( .I(n34016), .ZN(n5751) );
  CLKBUF_X4 U10429 ( .I(n21933), .Z(n20003) );
  INV_X2 U12459 ( .I(n18909), .ZN(n6894) );
  INV_X2 U3509 ( .I(n3014), .ZN(n1416) );
  INV_X2 U4984 ( .I(n22239), .ZN(n3181) );
  INV_X4 U6430 ( .I(n20266), .ZN(n1349) );
  OAI21_X2 U8036 ( .A1(n1521), .A2(n11033), .B(n7258), .ZN(n7260) );
  NAND2_X2 U3988 ( .A1(n4536), .A2(n36720), .ZN(n31446) );
  BUF_X2 U2466 ( .I(n29641), .Z(n6181) );
  OAI21_X2 U23304 ( .A1(n4600), .A2(n35525), .B(n12027), .ZN(n18123) );
  OAI21_X2 U28817 ( .A1(n33379), .A2(n19566), .B(n24467), .ZN(n24253) );
  INV_X4 U244 ( .I(n18875), .ZN(n1431) );
  NAND2_X1 U12820 ( .A1(n18532), .A2(n12146), .ZN(n2091) );
  INV_X4 U19566 ( .I(n12289), .ZN(n23533) );
  INV_X2 U19162 ( .I(n29937), .ZN(n16060) );
  INV_X2 U26468 ( .I(n19982), .ZN(n16544) );
  OAI22_X2 U8365 ( .A1(n1953), .A2(n2601), .B1(n31829), .B2(n1298), .ZN(n1951)
         );
  AOI22_X2 U11716 ( .A1(n10891), .A2(n10890), .B1(n7912), .B2(n35580), .ZN(
        n8506) );
  INV_X2 U16624 ( .I(n16186), .ZN(n4914) );
  INV_X1 U3204 ( .I(n25367), .ZN(n15791) );
  AOI22_X2 U8467 ( .A1(n22803), .A2(n12029), .B1(n10552), .B2(n1646), .ZN(
        n10551) );
  NAND2_X2 U1430 ( .A1(n2257), .A2(n6347), .ZN(n5894) );
  NAND3_X2 U1170 ( .A1(n6514), .A2(n36630), .A3(n4147), .ZN(n22971) );
  NAND2_X1 U975 ( .A1(n5387), .A2(n24853), .ZN(n198) );
  AOI21_X2 U5026 ( .A1(n17638), .A2(n22187), .B(n39607), .ZN(n17637) );
  NAND2_X2 U6547 ( .A1(n29937), .A2(n30049), .ZN(n2160) );
  CLKBUF_X4 U7270 ( .I(n21441), .Z(n21840) );
  OAI21_X2 U24420 ( .A1(n18253), .A2(n22322), .B(n22323), .ZN(n17970) );
  OAI21_X2 U11788 ( .A1(n20103), .A2(n18773), .B(n26734), .ZN(n21008) );
  INV_X4 U21247 ( .I(n15248), .ZN(n15389) );
  NOR2_X2 U341 ( .A1(n6115), .A2(n6114), .ZN(n30993) );
  INV_X1 U10409 ( .I(n21933), .ZN(n15696) );
  NAND2_X2 U8040 ( .A1(n29080), .A2(n1822), .ZN(n1821) );
  NAND2_X1 U18098 ( .A1(n20419), .A2(n35115), .ZN(n27333) );
  INV_X2 U16311 ( .I(n22765), .ZN(n19014) );
  NAND2_X2 U2993 ( .A1(n28115), .A2(n28246), .ZN(n21238) );
  OAI21_X1 U10502 ( .A1(n39656), .A2(n3562), .B(n31035), .ZN(n30824) );
  INV_X2 U1689 ( .I(n27895), .ZN(n981) );
  NOR2_X1 U1663 ( .A1(n815), .A2(n10089), .ZN(n8106) );
  NAND2_X2 U1230 ( .A1(n23533), .A2(n23535), .ZN(n5184) );
  INV_X2 U10268 ( .I(n22196), .ZN(n1327) );
  NAND2_X2 U12075 ( .A1(n9378), .A2(n7135), .ZN(n9377) );
  NAND2_X2 U14142 ( .A1(n31206), .A2(n14239), .ZN(n8659) );
  INV_X2 U25138 ( .I(n23955), .ZN(n21030) );
  NAND2_X2 U27678 ( .A1(n30396), .A2(n29871), .ZN(n33297) );
  AOI21_X2 U12917 ( .A1(n15899), .A2(n15968), .B(n13555), .ZN(n15898) );
  INV_X4 U26448 ( .I(n21137), .ZN(n28193) );
  INV_X2 U5259 ( .I(n24076), .ZN(n24075) );
  OAI21_X2 U1693 ( .A1(n37733), .A2(n5572), .B(n32507), .ZN(n2464) );
  BUF_X2 U4551 ( .I(n25553), .Z(n19581) );
  OAI22_X1 U7463 ( .A1(n3372), .A2(n12350), .B1(n3897), .B2(n3898), .ZN(n33192) );
  INV_X2 U3823 ( .I(n13728), .ZN(n7536) );
  INV_X2 U20477 ( .I(n22135), .ZN(n8017) );
  OAI21_X2 U9741 ( .A1(n35300), .A2(n24373), .B(n33937), .ZN(n12579) );
  NOR2_X2 U20083 ( .A1(n19530), .A2(n23085), .ZN(n19281) );
  NOR2_X1 U4183 ( .A1(n7615), .A2(n28442), .ZN(n33829) );
  INV_X2 U17937 ( .I(n19496), .ZN(n21587) );
  OAI21_X2 U12617 ( .A1(n1268), .A2(n20155), .B(n24712), .ZN(n1907) );
  OAI21_X2 U13267 ( .A1(n19119), .A2(n23281), .B(n1291), .ZN(n17443) );
  INV_X2 U5174 ( .I(n37218), .ZN(n23034) );
  INV_X2 U1933 ( .I(n23502), .ZN(n1294) );
  NOR2_X2 U3835 ( .A1(n24707), .A2(n34526), .ZN(n32477) );
  NAND3_X2 U2819 ( .A1(n25988), .A2(n25990), .A3(n38548), .ZN(n25766) );
  OR3_X1 U20728 ( .A1(n35586), .A2(n22996), .A3(n3310), .Z(n32159) );
  BUF_X2 U14044 ( .I(Key[156]), .Z(n19904) );
  OAI21_X2 U3002 ( .A1(n12392), .A2(n23111), .B(n23108), .ZN(n18527) );
  BUF_X4 U4790 ( .I(n19938), .Z(n15330) );
  INV_X2 U6251 ( .I(n32026), .ZN(n25545) );
  INV_X2 U945 ( .I(n12159), .ZN(n1843) );
  INV_X2 U23778 ( .I(n37084), .ZN(n14601) );
  AOI21_X1 U17359 ( .A1(n10846), .A2(n17885), .B(n10845), .ZN(n4739) );
  AOI22_X2 U1757 ( .A1(n12579), .A2(n24118), .B1(n12580), .B2(n14478), .ZN(
        n5139) );
  NAND2_X2 U11587 ( .A1(n27587), .A2(n12074), .ZN(n27039) );
  OAI22_X2 U1684 ( .A1(n21080), .A2(n9547), .B1(n21081), .B2(n18329), .ZN(
        n23908) );
  INV_X2 U17040 ( .I(n21152), .ZN(n10736) );
  INV_X2 U6986 ( .I(n24529), .ZN(n24710) );
  NOR2_X2 U6707 ( .A1(n9201), .A2(n13471), .ZN(n27319) );
  AOI22_X2 U21641 ( .A1(n11687), .A2(n34452), .B1(n33623), .B2(n13899), .ZN(
        n32337) );
  INV_X1 U4707 ( .I(n23944), .ZN(n30849) );
  AOI21_X2 U10309 ( .A1(n587), .A2(n13472), .B(n21565), .ZN(n3270) );
  INV_X2 U29789 ( .I(n29456), .ZN(n29377) );
  INV_X4 U1102 ( .I(n626), .ZN(n11673) );
  INV_X4 U7491 ( .I(n1962), .ZN(n29776) );
  INV_X4 U13988 ( .I(n14424), .ZN(n21787) );
  OAI21_X2 U16397 ( .A1(n38537), .A2(n28570), .B(n979), .ZN(n33663) );
  NOR2_X2 U10713 ( .A1(n16392), .A2(n16391), .ZN(n16390) );
  BUF_X4 U3242 ( .I(n10820), .Z(n196) );
  NAND2_X2 U1062 ( .A1(n26118), .A2(n1098), .ZN(n33485) );
  BUF_X2 U13564 ( .I(n22853), .Z(n22995) );
  INV_X2 U2843 ( .I(n9668), .ZN(n30716) );
  NAND2_X1 U4659 ( .A1(n24380), .A2(n32937), .ZN(n4178) );
  OAI21_X2 U12629 ( .A1(n35968), .A2(n35088), .B(n4176), .ZN(n17961) );
  NOR2_X2 U13357 ( .A1(n15373), .A2(n20076), .ZN(n7011) );
  AOI22_X1 U6940 ( .A1(n20030), .A2(n7445), .B1(n24794), .B2(n20029), .ZN(
        n20028) );
  INV_X2 U23583 ( .I(n17412), .ZN(n30240) );
  INV_X1 U7727 ( .I(n19667), .ZN(n28138) );
  INV_X4 U29551 ( .I(n39020), .ZN(n979) );
  INV_X2 U2818 ( .I(n20830), .ZN(n29378) );
  INV_X1 U2305 ( .I(n21445), .ZN(n21844) );
  NOR2_X2 U25212 ( .A1(n26118), .A2(n1098), .ZN(n20061) );
  NOR2_X2 U12287 ( .A1(n25506), .A2(n15635), .ZN(n15634) );
  NAND2_X2 U16759 ( .A1(n37544), .A2(n18667), .ZN(n11634) );
  OAI21_X2 U4030 ( .A1(n21954), .A2(n30996), .B(n22190), .ZN(n21956) );
  OAI21_X2 U1867 ( .A1(n25456), .A2(n25455), .B(n10674), .ZN(n25458) );
  NOR2_X2 U28118 ( .A1(n1117), .A2(n25379), .ZN(n25455) );
  INV_X1 U1745 ( .I(n9520), .ZN(n18329) );
  NAND2_X1 U14621 ( .A1(n29911), .A2(n7457), .ZN(n29931) );
  BUF_X2 U5896 ( .I(n20896), .Z(n31832) );
  INV_X1 U18046 ( .I(n5078), .ZN(n9899) );
  NAND2_X2 U5659 ( .A1(n26743), .A2(n11679), .ZN(n30722) );
  NOR2_X1 U22131 ( .A1(n23425), .A2(n10633), .ZN(n13579) );
  INV_X2 U5558 ( .I(n11834), .ZN(n25995) );
  NOR2_X2 U24808 ( .A1(n22833), .A2(n22937), .ZN(n15555) );
  BUF_X2 U8779 ( .I(Key[93]), .Z(n19804) );
  AOI21_X1 U15457 ( .A1(n22088), .A2(n31407), .B(n3002), .ZN(n22090) );
  NOR2_X2 U8576 ( .A1(n8749), .A2(n8679), .ZN(n22402) );
  BUF_X4 U8602 ( .I(n10463), .Z(n8749) );
  NAND2_X2 U8565 ( .A1(n21984), .A2(n20238), .ZN(n21985) );
  NOR2_X2 U8339 ( .A1(n3869), .A2(n24477), .ZN(n24234) );
  INV_X2 U7474 ( .I(n775), .ZN(n1058) );
  NOR2_X2 U13762 ( .A1(n4283), .A2(n6036), .ZN(n9904) );
  AND2_X1 U6615 ( .A1(n27066), .A2(n1000), .Z(n30485) );
  OAI21_X1 U12540 ( .A1(n24814), .A2(n9277), .B(n11121), .ZN(n12832) );
  INV_X1 U21094 ( .I(n3433), .ZN(n32232) );
  OAI22_X2 U12772 ( .A1(n11760), .A2(n7344), .B1(n17947), .B2(n14705), .ZN(
        n11759) );
  INV_X2 U5847 ( .I(n16252), .ZN(n29422) );
  BUF_X2 U4847 ( .I(n32675), .Z(n32318) );
  NOR2_X2 U20691 ( .A1(n8070), .A2(n7986), .ZN(n7987) );
  INV_X2 U6116 ( .I(n28473), .ZN(n9586) );
  AOI21_X2 U9708 ( .A1(n24332), .A2(n24336), .B(n19382), .ZN(n6955) );
  NAND2_X1 U4229 ( .A1(n8370), .A2(n8819), .ZN(n31781) );
  AOI21_X1 U18414 ( .A1(n5711), .A2(n5541), .B(n5710), .ZN(n6424) );
  NAND2_X2 U10167 ( .A1(n1671), .A2(n22289), .ZN(n1781) );
  CLKBUF_X2 U10454 ( .I(Key[20]), .Z(n19676) );
  NOR2_X1 U24457 ( .A1(n32843), .A2(n25815), .ZN(n193) );
  NOR2_X2 U29378 ( .A1(n25783), .A2(n10807), .ZN(n15552) );
  INV_X1 U16742 ( .I(n10071), .ZN(n17080) );
  NOR2_X2 U2935 ( .A1(n19136), .A2(n6036), .ZN(n15134) );
  NAND2_X1 U15164 ( .A1(n31353), .A2(n28656), .ZN(n10369) );
  INV_X1 U3528 ( .I(n29755), .ZN(n29741) );
  NAND3_X2 U22139 ( .A1(n1491), .A2(n19575), .A3(n14382), .ZN(n12220) );
  INV_X2 U8872 ( .I(n20113), .ZN(n29420) );
  OAI21_X2 U3412 ( .A1(n33442), .A2(n23704), .B(n24484), .ZN(n346) );
  NOR2_X2 U521 ( .A1(n7627), .A2(n7628), .ZN(n7397) );
  INV_X2 U4864 ( .I(n31664), .ZN(n17735) );
  NAND2_X2 U25446 ( .A1(n9288), .A2(n9287), .ZN(n33534) );
  NAND3_X2 U13506 ( .A1(n22746), .A2(n12032), .A3(n35040), .ZN(n11822) );
  NOR2_X1 U4670 ( .A1(n32787), .A2(n32786), .ZN(n32785) );
  NOR2_X2 U6398 ( .A1(n10418), .A2(n10417), .ZN(n22040) );
  NAND2_X2 U10811 ( .A1(n30166), .A2(n1181), .ZN(n30172) );
  INV_X2 U15604 ( .I(n319), .ZN(n16114) );
  CLKBUF_X4 U358 ( .I(n27772), .Z(n28282) );
  OAI21_X2 U16967 ( .A1(n24516), .A2(n38749), .B(n35801), .ZN(n24517) );
  OAI21_X2 U8117 ( .A1(n12629), .A2(n10055), .B(n1541), .ZN(n14025) );
  CLKBUF_X4 U19037 ( .I(n24878), .Z(n31861) );
  INV_X1 U17761 ( .I(n39112), .ZN(n8232) );
  INV_X2 U14769 ( .I(n19525), .ZN(n2338) );
  NAND2_X2 U29071 ( .A1(n25691), .A2(n18894), .ZN(n25568) );
  NAND3_X1 U14317 ( .A1(n14540), .A2(n17525), .A3(n32572), .ZN(n9953) );
  NAND2_X2 U20915 ( .A1(n7286), .A2(n19420), .ZN(n8318) );
  INV_X4 U10086 ( .I(n23028), .ZN(n1315) );
  INV_X2 U9350 ( .I(n26630), .ZN(n26761) );
  OAI21_X2 U4573 ( .A1(n38293), .A2(n24595), .B(n30960), .ZN(n25140) );
  NAND2_X2 U24510 ( .A1(n18412), .A2(n21920), .ZN(n21921) );
  NOR2_X2 U30287 ( .A1(n16107), .A2(n15112), .ZN(n5244) );
  OAI21_X2 U11882 ( .A1(n26922), .A2(n26764), .B(n26920), .ZN(n26737) );
  NAND2_X2 U2903 ( .A1(n2457), .A2(n5469), .ZN(n31847) );
  NAND2_X1 U8211 ( .A1(n7176), .A2(n9614), .ZN(n20030) );
  AOI22_X2 U16052 ( .A1(n32318), .A2(n17723), .B1(n12077), .B2(n30306), .ZN(
        n31481) );
  BUF_X2 U9138 ( .I(n27882), .Z(n28260) );
  AOI22_X2 U12158 ( .A1(n1243), .A2(n8377), .B1(n8376), .B2(n36404), .ZN(
        n11270) );
  OAI21_X2 U5886 ( .A1(n28034), .A2(n9969), .B(n7310), .ZN(n7309) );
  INV_X4 U2605 ( .I(n28191), .ZN(n28034) );
  OAI21_X1 U20503 ( .A1(n19017), .A2(n20376), .B(n21977), .ZN(n21978) );
  NAND2_X2 U6136 ( .A1(n1396), .A2(n9105), .ZN(n29479) );
  NAND2_X1 U17260 ( .A1(n16173), .A2(n27435), .ZN(n5998) );
  INV_X2 U16471 ( .I(n3974), .ZN(n14488) );
  NOR2_X1 U11795 ( .A1(n16402), .A2(n33396), .ZN(n16401) );
  AOI21_X1 U11306 ( .A1(n28272), .A2(n28012), .B(n8308), .ZN(n8307) );
  NOR2_X2 U2937 ( .A1(n6036), .A2(n4935), .ZN(n14925) );
  NAND2_X2 U7878 ( .A1(n26817), .A2(n20635), .ZN(n20634) );
  NOR2_X2 U10988 ( .A1(n5244), .A2(n5243), .ZN(n20845) );
  NAND2_X2 U12694 ( .A1(n24692), .A2(n30764), .ZN(n24693) );
  INV_X2 U8137 ( .I(n730), .ZN(n1530) );
  NAND3_X1 U24456 ( .A1(n24181), .A2(n277), .A3(n24398), .ZN(n18632) );
  NAND2_X1 U20015 ( .A1(n19028), .A2(n37377), .ZN(n11316) );
  NOR3_X2 U22904 ( .A1(n33843), .A2(n14209), .A3(n31597), .ZN(n12651) );
  INV_X1 U16532 ( .I(n14837), .ZN(n12314) );
  NAND2_X1 U11197 ( .A1(n20920), .A2(n39574), .ZN(n19414) );
  INV_X2 U6376 ( .I(n12015), .ZN(n963) );
  OAI22_X2 U23731 ( .A1(n29316), .A2(n38328), .B1(n29203), .B2(n39585), .ZN(
        n19706) );
  BUF_X2 U1645 ( .I(n18860), .Z(n8368) );
  INV_X2 U1496 ( .I(n20887), .ZN(n19133) );
  OAI21_X2 U9122 ( .A1(n10288), .A2(n16869), .B(n16950), .ZN(n10287) );
  INV_X2 U4929 ( .I(n13166), .ZN(n25422) );
  INV_X2 U7730 ( .I(n17410), .ZN(n1437) );
  INV_X2 U1534 ( .I(n4116), .ZN(n18657) );
  INV_X2 U27797 ( .I(n20070), .ZN(n28089) );
  NAND3_X2 U18036 ( .A1(n9456), .A2(n20962), .A3(n9457), .ZN(n5073) );
  AOI21_X2 U25153 ( .A1(n23262), .A2(n16047), .B(n23401), .ZN(n16757) );
  BUF_X2 U11448 ( .I(n27700), .Z(n19612) );
  NAND2_X2 U6578 ( .A1(n35248), .A2(n319), .ZN(n30470) );
  AOI21_X2 U13368 ( .A1(n23157), .A2(n23158), .B(n23156), .ZN(n6345) );
  NAND2_X1 U24061 ( .A1(n18814), .A2(n38145), .ZN(n20737) );
  BUF_X2 U4874 ( .I(n33324), .Z(n33154) );
  INV_X4 U10673 ( .I(n30844), .ZN(n6300) );
  INV_X4 U11422 ( .I(n988), .ZN(n28274) );
  NAND3_X2 U7053 ( .A1(n11214), .A2(n1134), .A3(n23383), .ZN(n3746) );
  NAND2_X1 U13862 ( .A1(n18954), .A2(n20003), .ZN(n3484) );
  AOI21_X1 U8661 ( .A1(n21522), .A2(n19511), .B(n21587), .ZN(n5104) );
  NAND3_X2 U1987 ( .A1(n32626), .A2(n7130), .A3(n32625), .ZN(n20907) );
  INV_X2 U23802 ( .I(n13091), .ZN(n28153) );
  BUF_X4 U4630 ( .I(n24759), .Z(n10019) );
  NOR2_X2 U12988 ( .A1(n914), .A2(n12953), .ZN(n4957) );
  INV_X2 U9950 ( .I(n19481), .ZN(n23588) );
  AOI21_X2 U2328 ( .A1(n28034), .A2(n36979), .B(n7309), .ZN(n11470) );
  INV_X1 U7568 ( .I(n1190), .ZN(n18098) );
  BUF_X4 U1776 ( .I(n14491), .Z(n32507) );
  INV_X2 U4337 ( .I(n21050), .ZN(n1218) );
  INV_X2 U6319 ( .I(n20484), .ZN(n24470) );
  AOI22_X2 U13723 ( .A1(n20280), .A2(n13519), .B1(n20282), .B2(n1340), .ZN(
        n19460) );
  INV_X2 U2770 ( .I(n38395), .ZN(n13632) );
  BUF_X2 U10423 ( .I(n21805), .Z(n19545) );
  BUF_X2 U8775 ( .I(Key[95]), .Z(n19885) );
  NAND2_X1 U8796 ( .A1(n20964), .A2(n29468), .ZN(n6343) );
  INV_X2 U10394 ( .I(n21111), .ZN(n8468) );
  AOI21_X2 U10045 ( .A1(n2350), .A2(n23201), .B(n33697), .ZN(n13527) );
  NAND2_X2 U6838 ( .A1(n4606), .A2(n30275), .ZN(n31825) );
  NOR2_X1 U3083 ( .A1(n6203), .A2(n6201), .ZN(n6208) );
  INV_X2 U10111 ( .I(n8197), .ZN(n23094) );
  NOR2_X2 U2779 ( .A1(n11090), .A2(n20528), .ZN(n11089) );
  INV_X2 U18543 ( .I(n27580), .ZN(n27532) );
  NAND2_X1 U24621 ( .A1(n25919), .A2(n16814), .ZN(n16813) );
  INV_X4 U7033 ( .I(n24461), .ZN(n1126) );
  BUF_X2 U30560 ( .I(n9861), .Z(n33921) );
  OAI21_X2 U22227 ( .A1(n31875), .A2(n997), .B(n13364), .ZN(n16248) );
  INV_X2 U3872 ( .I(n261), .ZN(n21565) );
  NAND2_X1 U20097 ( .A1(n18251), .A2(n18250), .ZN(n27324) );
  INV_X1 U17462 ( .I(n15159), .ZN(n1541) );
  INV_X2 U8904 ( .I(n8184), .ZN(n29497) );
  NAND3_X1 U2384 ( .A1(n26686), .A2(n18357), .A3(n33301), .ZN(n113) );
  INV_X4 U2737 ( .I(n15320), .ZN(n914) );
  BUF_X2 U14061 ( .I(Key[175]), .Z(n29805) );
  BUF_X2 U8774 ( .I(Key[4]), .Z(n19736) );
  BUF_X2 U6456 ( .I(Key[52]), .Z(n29238) );
  BUF_X2 U7315 ( .I(Key[0]), .Z(n29399) );
  BUF_X2 U6465 ( .I(Key[31]), .Z(n19843) );
  BUF_X2 U10465 ( .I(Key[45]), .Z(n30120) );
  BUF_X2 U14041 ( .I(Key[43]), .Z(n30068) );
  CLKBUF_X4 U10407 ( .I(n21743), .Z(n19542) );
  INV_X2 U6451 ( .I(n15354), .ZN(n13855) );
  BUF_X2 U7289 ( .I(n13679), .Z(n8597) );
  CLKBUF_X1 U14021 ( .I(n21722), .Z(n18855) );
  INV_X1 U14345 ( .I(n19902), .ZN(n31249) );
  INV_X1 U21020 ( .I(n19736), .ZN(n32218) );
  BUF_X2 U13990 ( .I(n21835), .Z(n19620) );
  INV_X1 U26614 ( .I(n33141), .ZN(n21620) );
  NOR2_X1 U13871 ( .A1(n21388), .A2(n21715), .ZN(n16290) );
  OAI21_X1 U13868 ( .A1(n21842), .A2(n21900), .B(n15031), .ZN(n12119) );
  NAND2_X1 U10345 ( .A1(n34021), .A2(n21554), .ZN(n10893) );
  NAND2_X1 U1476 ( .A1(n21622), .A2(n8467), .ZN(n2403) );
  INV_X2 U5794 ( .I(n22042), .ZN(n1338) );
  INV_X2 U27114 ( .I(n21980), .ZN(n22301) );
  NOR2_X1 U24738 ( .A1(n34488), .A2(n36303), .ZN(n19159) );
  INV_X2 U6396 ( .I(n22040), .ZN(n22289) );
  CLKBUF_X4 U10266 ( .I(n22294), .Z(n18854) );
  AOI22_X1 U10155 ( .A1(n21262), .A2(n22268), .B1(n21261), .B2(n32259), .ZN(
        n21260) );
  NOR2_X1 U13685 ( .A1(n20043), .A2(n21960), .ZN(n10025) );
  INV_X1 U13701 ( .I(n22213), .ZN(n12030) );
  NAND2_X1 U10134 ( .A1(n20146), .A2(n20148), .ZN(n19328) );
  INV_X1 U2097 ( .I(n17943), .ZN(n1670) );
  CLKBUF_X4 U2594 ( .I(n9873), .Z(n3475) );
  CLKBUF_X2 U2932 ( .I(n22744), .Z(n32863) );
  INV_X1 U13594 ( .I(n22604), .ZN(n11254) );
  INV_X1 U4391 ( .I(n1661), .ZN(n7158) );
  CLKBUF_X2 U5050 ( .I(n10962), .Z(n903) );
  BUF_X2 U2015 ( .I(n12925), .Z(n33247) );
  INV_X1 U14225 ( .I(n22974), .ZN(n1872) );
  BUF_X2 U4785 ( .I(n20840), .Z(n32032) );
  INV_X2 U19962 ( .I(n7327), .ZN(n14556) );
  NOR2_X1 U25722 ( .A1(n22974), .A2(n15163), .ZN(n16733) );
  INV_X2 U5992 ( .I(n14556), .ZN(n23114) );
  NOR2_X1 U16021 ( .A1(n18071), .A2(n20408), .ZN(n20743) );
  INV_X1 U12862 ( .I(n6827), .ZN(n31081) );
  OAI21_X1 U5100 ( .A1(n5786), .A2(n5785), .B(n19865), .ZN(n14352) );
  NAND2_X1 U21855 ( .A1(n23033), .A2(n16967), .ZN(n11435) );
  NOR2_X1 U21607 ( .A1(n23004), .A2(n23070), .ZN(n32326) );
  INV_X2 U13452 ( .I(n22512), .ZN(n4473) );
  AOI21_X1 U18343 ( .A1(n18516), .A2(n22924), .B(n32216), .ZN(n31736) );
  NAND2_X1 U1719 ( .A1(n11435), .A2(n23127), .ZN(n4597) );
  OAI21_X1 U13444 ( .A1(n22995), .A2(n23067), .B(n20024), .ZN(n8012) );
  AOI22_X1 U13399 ( .A1(n23112), .A2(n1142), .B1(n23113), .B2(n33196), .ZN(
        n18702) );
  NAND2_X1 U24392 ( .A1(n19361), .A2(n15503), .ZN(n15502) );
  INV_X2 U4217 ( .I(n17094), .ZN(n14845) );
  CLKBUF_X4 U6339 ( .I(n18682), .Z(n5487) );
  BUF_X2 U5750 ( .I(n34959), .Z(n3363) );
  CLKBUF_X4 U3997 ( .I(n31944), .Z(n30506) );
  INV_X2 U15838 ( .I(n33609), .ZN(n15787) );
  NAND2_X1 U1857 ( .A1(n18199), .A2(n37523), .ZN(n23274) );
  OAI21_X1 U5252 ( .A1(n22912), .A2(n22911), .B(n36191), .ZN(n22914) );
  INV_X1 U25263 ( .I(n23903), .ZN(n8704) );
  INV_X1 U1150 ( .I(n6527), .ZN(n5071) );
  INV_X1 U5279 ( .I(n23904), .ZN(n6051) );
  CLKBUF_X2 U13027 ( .I(n801), .Z(n7730) );
  CLKBUF_X4 U13048 ( .I(n23907), .Z(n24245) );
  CLKBUF_X2 U10602 ( .I(n24421), .Z(n30833) );
  CLKBUF_X4 U3722 ( .I(n36552), .Z(n6849) );
  CLKBUF_X4 U9810 ( .I(n10734), .Z(n2348) );
  OR2_X1 U6562 ( .A1(n15775), .A2(n16792), .Z(n30463) );
  NOR2_X1 U8340 ( .A1(n24446), .A2(n24445), .ZN(n13708) );
  OAI21_X1 U14495 ( .A1(n24426), .A2(n24258), .B(n2089), .ZN(n2088) );
  OR2_X1 U8319 ( .A1(n23958), .A2(n8193), .Z(n8194) );
  INV_X1 U1706 ( .I(n15018), .ZN(n16447) );
  NAND2_X1 U24881 ( .A1(n24474), .A2(n37916), .ZN(n24475) );
  NAND2_X1 U26417 ( .A1(n24386), .A2(n16375), .ZN(n16374) );
  BUF_X2 U1005 ( .I(n20728), .Z(n524) );
  BUF_X4 U3237 ( .I(n15266), .Z(n3120) );
  INV_X1 U4637 ( .I(n30530), .ZN(n30529) );
  OAI21_X1 U3664 ( .A1(n24794), .A2(n36321), .B(n24596), .ZN(n24598) );
  NAND2_X1 U1666 ( .A1(n31519), .A2(n32898), .ZN(n31328) );
  INV_X2 U5356 ( .I(n24623), .ZN(n21231) );
  BUF_X2 U4612 ( .I(n24614), .Z(n33821) );
  CLKBUF_X2 U4621 ( .I(n13966), .Z(n33480) );
  CLKBUF_X4 U6992 ( .I(n24623), .Z(n9277) );
  OAI21_X1 U3784 ( .A1(n15664), .A2(n34354), .B(n36471), .ZN(n13746) );
  NAND2_X1 U1658 ( .A1(n9277), .A2(n33818), .ZN(n14936) );
  INV_X1 U6963 ( .I(n24752), .ZN(n12706) );
  NAND2_X1 U951 ( .A1(n7342), .A2(n24659), .ZN(n24178) );
  INV_X1 U28785 ( .I(n24620), .ZN(n24084) );
  NAND2_X1 U20218 ( .A1(n24622), .A2(n32064), .ZN(n32063) );
  NOR2_X1 U12487 ( .A1(n16421), .A2(n16420), .ZN(n13398) );
  NOR2_X1 U2662 ( .A1(n9438), .A2(n2931), .ZN(n2930) );
  INV_X1 U1958 ( .I(n33038), .ZN(n6411) );
  INV_X1 U24864 ( .I(n24935), .ZN(n25024) );
  INV_X1 U24468 ( .I(n19418), .ZN(n25394) );
  INV_X1 U9564 ( .I(n39289), .ZN(n8879) );
  CLKBUF_X2 U12447 ( .I(n19418), .Z(n18298) );
  INV_X2 U6681 ( .I(n19582), .ZN(n6731) );
  CLKBUF_X4 U4506 ( .I(n11496), .Z(n32419) );
  OAI21_X1 U4501 ( .A1(n30377), .A2(n25341), .B(n1543), .ZN(n25344) );
  NAND2_X1 U12399 ( .A1(n25066), .A2(n35887), .ZN(n25067) );
  OAI21_X1 U1240 ( .A1(n5483), .A2(n7853), .B(n18810), .ZN(n31322) );
  OAI21_X1 U26900 ( .A1(n32419), .A2(n36249), .B(n17472), .ZN(n17471) );
  INV_X2 U21851 ( .I(n39140), .ZN(n1244) );
  NAND2_X1 U4497 ( .A1(n2958), .A2(n13465), .ZN(n32044) );
  INV_X2 U22287 ( .I(n26041), .ZN(n32469) );
  NAND2_X1 U25210 ( .A1(n18838), .A2(n25509), .ZN(n19042) );
  NAND2_X1 U15042 ( .A1(n6221), .A2(n3575), .ZN(n6220) );
  NAND2_X1 U12119 ( .A1(n25737), .A2(n9859), .ZN(n6153) );
  INV_X2 U17155 ( .I(n17212), .ZN(n8481) );
  INV_X1 U12175 ( .I(n26129), .ZN(n8543) );
  NAND2_X1 U9384 ( .A1(n6152), .A2(n6153), .ZN(n6150) );
  INV_X1 U25236 ( .I(n25854), .ZN(n14952) );
  NAND2_X1 U7985 ( .A1(n6478), .A2(n8255), .ZN(n6219) );
  INV_X1 U3446 ( .I(n35238), .ZN(n13147) );
  NAND2_X1 U12047 ( .A1(n25739), .A2(n30621), .ZN(n10509) );
  CLKBUF_X2 U18448 ( .I(n26520), .Z(n32528) );
  OR2_X1 U20616 ( .A1(n35269), .A2(n36392), .Z(n32693) );
  INV_X2 U17930 ( .I(n9081), .ZN(n8155) );
  INV_X2 U2795 ( .I(n14080), .ZN(n26708) );
  INV_X1 U7936 ( .I(n9899), .ZN(n9269) );
  NAND2_X1 U27161 ( .A1(n26266), .A2(n26655), .ZN(n19204) );
  INV_X2 U588 ( .I(n26688), .ZN(n26980) );
  NAND2_X1 U11750 ( .A1(n14485), .A2(n5405), .ZN(n4483) );
  INV_X1 U27574 ( .I(n26865), .ZN(n26775) );
  NAND2_X1 U20162 ( .A1(n20547), .A2(n20754), .ZN(n7469) );
  OAI21_X1 U29339 ( .A1(n26983), .A2(n852), .B(n17097), .ZN(n26984) );
  NAND2_X1 U23438 ( .A1(n26985), .A2(n26984), .ZN(n18047) );
  CLKBUF_X4 U25589 ( .I(n7974), .Z(n32976) );
  INV_X2 U22767 ( .I(n11020), .ZN(n17166) );
  INV_X2 U509 ( .I(n14153), .ZN(n27274) );
  INV_X1 U9186 ( .I(n10461), .ZN(n27429) );
  INV_X1 U5736 ( .I(n19061), .ZN(n32771) );
  NOR2_X1 U6711 ( .A1(n27084), .A2(n27274), .ZN(n5664) );
  OAI21_X1 U24035 ( .A1(n10677), .A2(n27410), .B(n32771), .ZN(n399) );
  OAI21_X1 U19671 ( .A1(n31943), .A2(n35299), .B(n9680), .ZN(n26447) );
  BUF_X4 U3690 ( .I(n10621), .Z(n33690) );
  INV_X1 U2088 ( .I(n12971), .ZN(n11502) );
  INV_X2 U29865 ( .I(n33522), .ZN(n3158) );
  INV_X2 U19902 ( .I(n7281), .ZN(n16065) );
  BUF_X4 U17161 ( .I(n27671), .Z(n28024) );
  BUF_X2 U4268 ( .I(n1455), .Z(n33405) );
  INV_X2 U5484 ( .I(n12218), .ZN(n14500) );
  NAND2_X1 U9044 ( .A1(n28257), .A2(n28258), .ZN(n11025) );
  CLKBUF_X2 U4259 ( .I(n12909), .Z(n33002) );
  NOR2_X1 U11388 ( .A1(n438), .A2(n28205), .ZN(n1753) );
  NAND2_X1 U9041 ( .A1(n20639), .A2(n27974), .ZN(n8265) );
  INV_X1 U11301 ( .I(n28004), .ZN(n7984) );
  NOR2_X1 U415 ( .A1(n3198), .A2(n32150), .ZN(n33418) );
  OAI22_X1 U11284 ( .A1(n8327), .A2(n4347), .B1(n8149), .B2(n8326), .ZN(n8325)
         );
  INV_X2 U27299 ( .I(n28685), .ZN(n1429) );
  INV_X2 U20101 ( .I(n7428), .ZN(n16778) );
  INV_X2 U11155 ( .I(n10544), .ZN(n3252) );
  INV_X2 U355 ( .I(n15792), .ZN(n17978) );
  NOR2_X1 U18074 ( .A1(n14516), .A2(n15631), .ZN(n15630) );
  NOR2_X1 U11074 ( .A1(n32315), .A2(n32314), .ZN(n10304) );
  OAI21_X1 U11072 ( .A1(n17073), .A2(n32595), .B(n3191), .ZN(n15323) );
  NAND2_X1 U16924 ( .A1(n28718), .A2(n16505), .ZN(n31608) );
  CLKBUF_X1 U6038 ( .I(n29146), .Z(n30888) );
  CLKBUF_X2 U20087 ( .I(n29121), .Z(n32022) );
  INV_X2 U18785 ( .I(n20460), .ZN(n29081) );
  INV_X2 U8903 ( .I(n771), .ZN(n1176) );
  CLKBUF_X2 U10848 ( .I(n29483), .Z(n19734) );
  INV_X2 U28063 ( .I(n29196), .ZN(n29701) );
  INV_X2 U1919 ( .I(n8529), .ZN(n14437) );
  NAND2_X1 U2471 ( .A1(n29702), .A2(n8941), .ZN(n7502) );
  OAI21_X1 U21889 ( .A1(n30051), .A2(n19909), .B(n10671), .ZN(n10670) );
  NAND2_X1 U27385 ( .A1(n17540), .A2(n17539), .ZN(n33246) );
  OAI21_X1 U8868 ( .A1(n1060), .A2(n29702), .B(n14511), .ZN(n16389) );
  NAND2_X1 U10734 ( .A1(n6207), .A2(n13573), .ZN(n6206) );
  CLKBUF_X2 U8787 ( .I(Key[166]), .Z(n29442) );
  CLKBUF_X2 U14034 ( .I(Key[107]), .Z(n19801) );
  CLKBUF_X2 U8769 ( .I(Key[167]), .Z(n29506) );
  BUF_X2 U14065 ( .I(Key[132]), .Z(n19887) );
  CLKBUF_X2 U7318 ( .I(Key[91]), .Z(n29831) );
  CLKBUF_X2 U5826 ( .I(Key[150]), .Z(n9981) );
  BUF_X2 U10489 ( .I(Key[92]), .Z(n19851) );
  BUF_X2 U6453 ( .I(Key[106]), .Z(n19780) );
  BUF_X2 U7317 ( .I(Key[33]), .Z(n19805) );
  BUF_X2 U8766 ( .I(Key[129]), .Z(n19775) );
  BUF_X2 U14016 ( .I(n21674), .Z(n19641) );
  INV_X1 U7293 ( .I(n29285), .ZN(n1160) );
  INV_X1 U13918 ( .I(n21749), .ZN(n21715) );
  INV_X2 U5786 ( .I(n22301), .ZN(n20357) );
  NAND2_X1 U2895 ( .A1(n10762), .A2(n11327), .ZN(n22213) );
  OAI22_X1 U19488 ( .A1(n11171), .A2(n35754), .B1(n34246), .B2(n22360), .ZN(
        n15488) );
  BUF_X2 U4021 ( .I(n11778), .Z(n33697) );
  BUF_X2 U13573 ( .I(n23089), .Z(n19488) );
  INV_X2 U19289 ( .I(n19588), .ZN(n22512) );
  BUF_X4 U1262 ( .I(n8660), .Z(n6684) );
  INV_X1 U2896 ( .I(n13217), .ZN(n17090) );
  INV_X1 U1904 ( .I(n23272), .ZN(n18939) );
  CLKBUF_X2 U13297 ( .I(n21068), .Z(n10024) );
  NOR2_X1 U24906 ( .A1(n18762), .A2(n1039), .ZN(n20997) );
  NOR2_X1 U29938 ( .A1(n4183), .A2(n37319), .ZN(n33532) );
  OAI21_X1 U12822 ( .A1(n12120), .A2(n24469), .B(n8200), .ZN(n10751) );
  AOI21_X1 U6970 ( .A1(n4666), .A2(n24132), .B(n1128), .ZN(n30530) );
  NAND2_X1 U5357 ( .A1(n24591), .A2(n24694), .ZN(n16079) );
  NAND2_X1 U17378 ( .A1(n16050), .A2(n16051), .ZN(n2931) );
  INV_X1 U12522 ( .I(n25040), .ZN(n11964) );
  NAND2_X1 U9554 ( .A1(n5541), .A2(n5519), .ZN(n8033) );
  INV_X2 U27774 ( .I(n33948), .ZN(n19963) );
  NOR2_X1 U5453 ( .A1(n299), .A2(n19495), .ZN(n25066) );
  CLKBUF_X4 U23372 ( .I(n16836), .Z(n32654) );
  OAI21_X1 U9476 ( .A1(n7956), .A2(n30633), .B(n19490), .ZN(n2766) );
  INV_X1 U12114 ( .I(n25933), .ZN(n12721) );
  OAI21_X1 U3763 ( .A1(n25737), .A2(n25887), .B(n26070), .ZN(n6152) );
  OAI21_X1 U1697 ( .A1(n8543), .A2(n34745), .B(n31827), .ZN(n25405) );
  NOR2_X1 U3893 ( .A1(n4138), .A2(n26797), .ZN(n9179) );
  NAND2_X1 U11800 ( .A1(n9731), .A2(n26951), .ZN(n4689) );
  INV_X2 U2126 ( .I(n12755), .ZN(n6891) );
  BUF_X1 U3928 ( .I(n31014), .Z(n30871) );
  NAND3_X1 U606 ( .A1(n1474), .A2(n16237), .A3(n16263), .ZN(n27312) );
  NAND2_X1 U29412 ( .A1(n4782), .A2(n3531), .ZN(n1939) );
  NAND2_X1 U9146 ( .A1(n10574), .A2(n16966), .ZN(n10580) );
  CLKBUF_X1 U26744 ( .I(n27779), .Z(n20772) );
  BUF_X2 U16281 ( .I(n5402), .Z(n4347) );
  BUF_X2 U30535 ( .I(n37056), .Z(n33902) );
  INV_X1 U7705 ( .I(n6990), .ZN(n8522) );
  INV_X2 U256 ( .I(n5237), .ZN(n9141) );
  INV_X1 U11131 ( .I(n14760), .ZN(n12717) );
  INV_X1 U7925 ( .I(n28301), .ZN(n21025) );
  INV_X1 U11122 ( .I(n28370), .ZN(n13824) );
  NAND2_X2 U158 ( .A1(n11665), .A2(n11664), .ZN(n28840) );
  AND2_X1 U10850 ( .A1(n21299), .A2(n15153), .Z(n10628) );
  CLKBUF_X2 U5832 ( .I(n29684), .Z(n19497) );
  NOR2_X2 U4433 ( .A1(n25939), .A2(n17915), .ZN(n20612) );
  BUF_X2 U2963 ( .I(n9001), .Z(n32309) );
  INV_X2 U28079 ( .I(n21184), .ZN(n29454) );
  INV_X2 U9636 ( .I(n24635), .ZN(n3125) );
  INV_X4 U4533 ( .I(n12246), .ZN(n13366) );
  BUF_X2 U13985 ( .I(n15370), .Z(n14783) );
  BUF_X2 U4228 ( .I(n18450), .Z(n452) );
  BUF_X2 U6424 ( .I(n19387), .Z(n4759) );
  INV_X1 U10412 ( .I(n21777), .ZN(n21465) );
  NOR2_X1 U4894 ( .A1(n35921), .A2(n1348), .ZN(n15456) );
  NAND2_X1 U8723 ( .A1(n10120), .A2(n8799), .ZN(n13701) );
  INV_X1 U6156 ( .I(n19641), .ZN(n33053) );
  NAND2_X1 U12309 ( .A1(n3562), .A2(n10629), .ZN(n31035) );
  NOR2_X1 U27471 ( .A1(n19479), .A2(n19091), .ZN(n21632) );
  INV_X1 U1517 ( .I(n35921), .ZN(n21440) );
  NOR2_X1 U2191 ( .A1(n35921), .A2(n18152), .ZN(n21842) );
  AOI21_X1 U24751 ( .A1(n21656), .A2(n17938), .B(n21780), .ZN(n18877) );
  OAI21_X1 U13916 ( .A1(n21465), .A2(n19091), .B(n21939), .ZN(n15437) );
  NAND2_X1 U30373 ( .A1(n8700), .A2(n21775), .ZN(n19075) );
  BUF_X2 U10406 ( .I(n13473), .Z(n13472) );
  NAND2_X1 U2200 ( .A1(n15696), .A2(n32164), .ZN(n32163) );
  NOR2_X1 U2007 ( .A1(n37111), .A2(n32123), .ZN(n20368) );
  NOR2_X1 U21947 ( .A1(n18412), .A2(n21111), .ZN(n21621) );
  INV_X1 U6418 ( .I(n18926), .ZN(n21557) );
  INV_X1 U20666 ( .I(n7935), .ZN(n14837) );
  NOR2_X1 U27340 ( .A1(n8700), .A2(n18710), .ZN(n21940) );
  NAND3_X1 U24532 ( .A1(n19517), .A2(n21672), .A3(n18219), .ZN(n16654) );
  AOI22_X1 U17769 ( .A1(n8700), .A2(n19479), .B1(n19350), .B2(n21775), .ZN(
        n18712) );
  NAND2_X1 U28253 ( .A1(n21666), .A2(n32412), .ZN(n21437) );
  AOI21_X1 U13874 ( .A1(n17679), .A2(n21309), .B(n17678), .ZN(n6669) );
  NOR2_X1 U24733 ( .A1(n15097), .A2(n21822), .ZN(n15096) );
  INV_X1 U24754 ( .I(n21932), .ZN(n21607) );
  OAI21_X1 U13932 ( .A1(n21333), .A2(n2531), .B(n21889), .ZN(n15814) );
  NOR2_X1 U1492 ( .A1(n13472), .A2(n5751), .ZN(n21377) );
  NOR2_X1 U5008 ( .A1(n20328), .A2(n21551), .ZN(n21653) );
  AOI21_X1 U25953 ( .A1(n21498), .A2(n20003), .B(n32164), .ZN(n16287) );
  OAI21_X1 U27341 ( .A1(n21775), .A2(n18710), .B(n8700), .ZN(n21609) );
  OAI22_X1 U26070 ( .A1(n21437), .A2(n19620), .B1(n20682), .B2(n21666), .ZN(
        n15490) );
  OAI21_X1 U13863 ( .A1(n21467), .A2(n21468), .B(n11411), .ZN(n2737) );
  INV_X2 U1976 ( .I(n21587), .ZN(n21588) );
  NOR2_X1 U8653 ( .A1(n16901), .A2(n3865), .ZN(n3864) );
  BUF_X2 U6401 ( .I(n22389), .Z(n4239) );
  NAND2_X1 U13759 ( .A1(n14027), .A2(n17086), .ZN(n17664) );
  NAND2_X1 U16601 ( .A1(n8496), .A2(n19373), .ZN(n22069) );
  NOR2_X1 U6395 ( .A1(n18303), .A2(n1746), .ZN(n3086) );
  INV_X1 U10273 ( .I(n11044), .ZN(n22220) );
  INV_X1 U14165 ( .I(n11344), .ZN(n22325) );
  INV_X1 U6394 ( .I(n22362), .ZN(n1672) );
  INV_X1 U6402 ( .I(n22389), .ZN(n4240) );
  NOR2_X1 U17243 ( .A1(n17074), .A2(n10632), .ZN(n10631) );
  NAND2_X1 U18844 ( .A1(n6036), .A2(n22315), .ZN(n18674) );
  INV_X1 U10275 ( .I(n19373), .ZN(n1681) );
  NAND2_X1 U26031 ( .A1(n7613), .A2(n22184), .ZN(n21974) );
  AOI21_X1 U10236 ( .A1(n6451), .A2(n1151), .B(n22177), .ZN(n16282) );
  NAND2_X1 U28377 ( .A1(n1048), .A2(n21973), .ZN(n21975) );
  NAND2_X1 U21861 ( .A1(n36563), .A2(n22332), .ZN(n22065) );
  INV_X1 U4979 ( .I(n22364), .ZN(n22366) );
  INV_X1 U4803 ( .I(n22315), .ZN(n22156) );
  INV_X1 U1408 ( .I(n3269), .ZN(n3268) );
  INV_X2 U5788 ( .I(n12077), .ZN(n17723) );
  INV_X1 U8581 ( .I(n22289), .ZN(n17531) );
  INV_X1 U18481 ( .I(n22215), .ZN(n22361) );
  INV_X1 U3131 ( .I(n20889), .ZN(n22140) );
  AOI21_X1 U20604 ( .A1(n164), .A2(n22293), .B(n22140), .ZN(n33792) );
  NOR2_X1 U9006 ( .A1(n8118), .A2(n22148), .ZN(n30706) );
  NAND2_X1 U1764 ( .A1(n22064), .A2(n3680), .ZN(n3679) );
  INV_X1 U5450 ( .I(n22332), .ZN(n22252) );
  NAND3_X1 U15641 ( .A1(n3181), .A2(n34407), .A3(n13632), .ZN(n21926) );
  NAND2_X1 U1406 ( .A1(n8348), .A2(n7613), .ZN(n20256) );
  AOI21_X1 U26544 ( .A1(n22140), .A2(n33713), .B(n18854), .ZN(n20354) );
  OAI21_X1 U17907 ( .A1(n22498), .A2(n1154), .B(n31648), .ZN(n18635) );
  INV_X1 U4982 ( .I(n22741), .ZN(n11500) );
  INV_X1 U6372 ( .I(n20353), .ZN(n22583) );
  INV_X1 U10122 ( .I(n22529), .ZN(n22515) );
  INV_X1 U26666 ( .I(n22699), .ZN(n17223) );
  INV_X1 U16458 ( .I(n22789), .ZN(n22601) );
  NOR2_X1 U2042 ( .A1(n1142), .A2(n12392), .ZN(n33763) );
  INV_X2 U2038 ( .I(n22929), .ZN(n22865) );
  INV_X1 U1318 ( .I(n3952), .ZN(n23032) );
  INV_X2 U17563 ( .I(n23078), .ZN(n23182) );
  INV_X1 U24005 ( .I(n782), .ZN(n23084) );
  NAND2_X1 U24829 ( .A1(n23169), .A2(n531), .ZN(n18147) );
  NAND2_X1 U13473 ( .A1(n1042), .A2(n1320), .ZN(n3200) );
  BUF_X2 U25972 ( .I(n21132), .Z(n33045) );
  INV_X1 U23498 ( .I(n301), .ZN(n32677) );
  INV_X1 U10106 ( .I(n23131), .ZN(n23211) );
  NAND2_X1 U5995 ( .A1(n23181), .A2(n23078), .ZN(n8673) );
  NOR2_X1 U27322 ( .A1(n9954), .A2(n18679), .ZN(n19659) );
  NOR2_X1 U28565 ( .A1(n22866), .A2(n22865), .ZN(n22867) );
  NAND3_X1 U8751 ( .A1(n18244), .A2(n13042), .A3(n23101), .ZN(n30676) );
  INV_X2 U8551 ( .I(n23125), .ZN(n23197) );
  NOR2_X1 U10052 ( .A1(n14396), .A2(n13719), .ZN(n14724) );
  INV_X1 U16597 ( .I(n23067), .ZN(n4107) );
  INV_X1 U1319 ( .I(n3273), .ZN(n22955) );
  NOR2_X1 U20186 ( .A1(n13734), .A2(n903), .ZN(n13775) );
  OR2_X1 U13541 ( .A1(n34014), .A2(n59), .Z(n23127) );
  OAI21_X1 U5110 ( .A1(n22867), .A2(n22991), .B(n39500), .ZN(n22868) );
  AOI21_X1 U8471 ( .A1(n272), .A2(n19351), .B(n9238), .ZN(n14189) );
  AOI21_X1 U10009 ( .A1(n36839), .A2(n23214), .B(n5569), .ZN(n2254) );
  AOI21_X1 U24432 ( .A1(n1316), .A2(n20174), .B(n1648), .ZN(n15503) );
  NAND2_X1 U15096 ( .A1(n22899), .A2(n36369), .ZN(n31351) );
  NOR2_X1 U13537 ( .A1(n3273), .A2(n19621), .ZN(n3542) );
  NAND2_X1 U21415 ( .A1(n23023), .A2(n9080), .ZN(n23027) );
  OAI21_X1 U4210 ( .A1(n13775), .A2(n23105), .B(n23104), .ZN(n4903) );
  NOR2_X1 U2752 ( .A1(n14882), .A2(n13408), .ZN(n13407) );
  NAND3_X1 U28609 ( .A1(n33045), .A2(n17691), .A3(n23178), .ZN(n23180) );
  OAI21_X1 U13370 ( .A1(n3547), .A2(n3546), .B(n19621), .ZN(n3545) );
  AOI21_X1 U15031 ( .A1(n6500), .A2(n1650), .B(n6498), .ZN(n6497) );
  INV_X2 U27628 ( .I(n32024), .ZN(n33287) );
  INV_X1 U3451 ( .I(n5357), .ZN(n12790) );
  CLKBUF_X2 U2100 ( .I(n17094), .Z(n14901) );
  INV_X1 U7118 ( .I(n23566), .ZN(n1643) );
  INV_X2 U13340 ( .I(n23496), .ZN(n23315) );
  AOI21_X1 U3863 ( .A1(n35068), .A2(n13305), .B(n35501), .ZN(n13304) );
  NAND2_X1 U18449 ( .A1(n33496), .A2(n10480), .ZN(n23284) );
  INV_X1 U2978 ( .I(n23308), .ZN(n1631) );
  NAND2_X1 U2552 ( .A1(n23307), .A2(n16182), .ZN(n23479) );
  INV_X1 U20667 ( .I(n23250), .ZN(n7939) );
  INV_X1 U1180 ( .I(n12154), .ZN(n20955) );
  AND2_X1 U17529 ( .A1(n71), .A2(n70), .Z(n31586) );
  NAND2_X1 U8379 ( .A1(n1290), .A2(n9862), .ZN(n23439) );
  NAND2_X1 U13130 ( .A1(n23439), .A2(n23440), .ZN(n9971) );
  NAND2_X1 U6326 ( .A1(n23575), .A2(n1134), .ZN(n3583) );
  NAND3_X1 U28619 ( .A1(n1134), .A2(n23571), .A3(n7485), .ZN(n23232) );
  INV_X1 U9964 ( .I(n17511), .ZN(n23474) );
  OAI21_X1 U13146 ( .A1(n22967), .A2(n23493), .B(n22966), .ZN(n22972) );
  NAND4_X1 U7115 ( .A1(n23432), .A2(n23433), .A3(n23434), .A4(n23431), .ZN(
        n23559) );
  NOR2_X1 U7094 ( .A1(n23624), .A2(n33894), .ZN(n23625) );
  NOR2_X1 U6674 ( .A1(n4600), .A2(n1310), .ZN(n21156) );
  NOR2_X1 U23776 ( .A1(n13305), .A2(n33349), .ZN(n23281) );
  AOI21_X1 U28647 ( .A1(n18284), .A2(n5083), .B(n23458), .ZN(n23372) );
  INV_X1 U13308 ( .I(n18989), .ZN(n16484) );
  AOI21_X1 U2517 ( .A1(n23312), .A2(n6421), .B(n1637), .ZN(n23313) );
  NAND3_X1 U5243 ( .A1(n33720), .A2(n33719), .A3(n12154), .ZN(n15495) );
  NAND2_X1 U9874 ( .A1(n35545), .A2(n36965), .ZN(n8054) );
  OAI21_X1 U21764 ( .A1(n32363), .A2(n33721), .B(n32362), .ZN(n23369) );
  OAI21_X1 U20233 ( .A1(n23282), .A2(n39194), .B(n32068), .ZN(n16883) );
  NAND2_X1 U28623 ( .A1(n36564), .A2(n36027), .ZN(n23259) );
  OAI21_X1 U25160 ( .A1(n12093), .A2(n36027), .B(n36564), .ZN(n14721) );
  NAND2_X1 U17484 ( .A1(n10989), .A2(n8054), .ZN(n8053) );
  INV_X1 U8364 ( .I(n23774), .ZN(n2221) );
  NAND3_X1 U9833 ( .A1(n36701), .A2(n36011), .A3(n1160), .ZN(n12819) );
  INV_X1 U1152 ( .I(n23899), .ZN(n20340) );
  INV_X1 U28795 ( .I(n24300), .ZN(n24110) );
  NAND2_X1 U18174 ( .A1(n12235), .A2(n16081), .ZN(n31697) );
  INV_X1 U14451 ( .I(n2052), .ZN(n24383) );
  INV_X1 U6321 ( .I(n16792), .ZN(n11585) );
  OAI21_X1 U9791 ( .A1(n19402), .A2(n37848), .B(n6515), .ZN(n24198) );
  NAND2_X1 U24276 ( .A1(n1597), .A2(n24143), .ZN(n14156) );
  NAND2_X1 U9766 ( .A1(n24359), .A2(n19895), .ZN(n4051) );
  NAND2_X1 U21506 ( .A1(n39605), .A2(n24282), .ZN(n32492) );
  INV_X1 U12895 ( .I(n19864), .ZN(n20396) );
  NAND2_X1 U9768 ( .A1(n17871), .A2(n33450), .ZN(n24152) );
  NAND2_X1 U1729 ( .A1(n24194), .A2(n6515), .ZN(n32491) );
  OAI21_X1 U1787 ( .A1(n1128), .A2(n1130), .B(n32069), .ZN(n24474) );
  NAND2_X1 U12849 ( .A1(n24473), .A2(n39309), .ZN(n2579) );
  NOR2_X1 U8328 ( .A1(n2348), .A2(n1285), .ZN(n14292) );
  NAND2_X1 U28812 ( .A1(n1599), .A2(n13453), .ZN(n24217) );
  NOR2_X1 U8299 ( .A1(n24390), .A2(n2348), .ZN(n16829) );
  NAND2_X1 U1712 ( .A1(n12481), .A2(n12202), .ZN(n32183) );
  NOR2_X1 U22917 ( .A1(n32891), .A2(n17911), .ZN(n5855) );
  INV_X1 U13004 ( .I(n33450), .ZN(n24449) );
  NOR2_X1 U3360 ( .A1(n10008), .A2(n17810), .ZN(n32938) );
  NOR2_X1 U9717 ( .A1(n24411), .A2(n37651), .ZN(n12423) );
  AOI21_X1 U17758 ( .A1(n18116), .A2(n33240), .B(n39373), .ZN(n31621) );
  OAI21_X1 U6999 ( .A1(n13881), .A2(n8581), .B(n14392), .ZN(n13742) );
  OAI21_X1 U9698 ( .A1(n24472), .A2(n24471), .B(n1130), .ZN(n24476) );
  NOR2_X1 U12965 ( .A1(n6839), .A2(n19942), .ZN(n9722) );
  NOR2_X1 U12959 ( .A1(n801), .A2(n24266), .ZN(n11194) );
  NAND2_X1 U6969 ( .A1(n10116), .A2(n17087), .ZN(n5388) );
  NAND2_X1 U12395 ( .A1(n31044), .A2(n24434), .ZN(n24511) );
  INV_X2 U24749 ( .I(n15467), .ZN(n32882) );
  AOI22_X1 U5964 ( .A1(n5358), .A2(n37264), .B1(n24147), .B2(n1604), .ZN(n5359) );
  INV_X1 U8253 ( .I(n35981), .ZN(n1583) );
  INV_X2 U26820 ( .I(n15426), .ZN(n19901) );
  NAND2_X1 U20158 ( .A1(n24620), .A2(n19868), .ZN(n24622) );
  NOR2_X1 U5379 ( .A1(n16210), .A2(n24782), .ZN(n7342) );
  NAND4_X1 U3832 ( .A1(n13045), .A2(n23796), .A3(n13048), .A4(n13047), .ZN(
        n13046) );
  AOI21_X1 U25202 ( .A1(n5056), .A2(n958), .B(n16077), .ZN(n16076) );
  NOR2_X1 U12524 ( .A1(n18168), .A2(n6037), .ZN(n8578) );
  NAND2_X1 U25206 ( .A1(n24695), .A2(n19565), .ZN(n24619) );
  INV_X1 U6990 ( .I(n24782), .ZN(n24660) );
  NAND2_X1 U981 ( .A1(n24698), .A2(n37097), .ZN(n24581) );
  AOI21_X1 U3667 ( .A1(n24794), .A2(n7445), .B(n36321), .ZN(n10141) );
  NAND2_X1 U12723 ( .A1(n31796), .A2(n37477), .ZN(n1948) );
  NAND2_X1 U20024 ( .A1(n24619), .A2(n11126), .ZN(n11258) );
  NOR2_X1 U20036 ( .A1(n24732), .A2(n24639), .ZN(n12782) );
  OAI21_X1 U1578 ( .A1(n14999), .A2(n1566), .B(n33480), .ZN(n30941) );
  NAND2_X1 U9651 ( .A1(n11712), .A2(n24592), .ZN(n3750) );
  INV_X1 U27708 ( .I(n39196), .ZN(n1574) );
  NAND2_X1 U28700 ( .A1(n35901), .A2(n34354), .ZN(n23705) );
  NAND2_X1 U28097 ( .A1(n33344), .A2(n7520), .ZN(n18468) );
  INV_X2 U972 ( .I(n1580), .ZN(n7831) );
  OR2_X1 U2659 ( .A1(n15266), .A2(n7520), .Z(n24849) );
  NOR2_X1 U3057 ( .A1(n11712), .A2(n24849), .ZN(n24850) );
  NAND2_X1 U1661 ( .A1(n37983), .A2(n39279), .ZN(n30700) );
  OAI21_X1 U10348 ( .A1(n7286), .A2(n8314), .B(n30554), .ZN(n24834) );
  OAI21_X1 U28883 ( .A1(n37396), .A2(n4973), .B(n24733), .ZN(n24595) );
  NOR2_X1 U3831 ( .A1(n5871), .A2(n31722), .ZN(n18504) );
  NAND3_X1 U12555 ( .A1(n24747), .A2(n24887), .A3(n13735), .ZN(n16195) );
  OAI21_X1 U9608 ( .A1(n4909), .A2(n24608), .B(n4908), .ZN(n7064) );
  NAND3_X1 U28855 ( .A1(n24691), .A2(n24765), .A3(n18324), .ZN(n24493) );
  NAND2_X1 U28847 ( .A1(n34138), .A2(n24795), .ZN(n24439) );
  NAND2_X1 U26131 ( .A1(n34138), .A2(n35981), .ZN(n17267) );
  NAND2_X1 U2012 ( .A1(n30764), .A2(n24717), .ZN(n24720) );
  NAND2_X1 U28886 ( .A1(n19886), .A2(n33821), .ZN(n24616) );
  AOI22_X1 U3967 ( .A1(n24671), .A2(n1119), .B1(n24670), .B2(n30843), .ZN(
        n12418) );
  NOR3_X1 U1554 ( .A1(n18570), .A2(n31346), .A3(n35521), .ZN(n18569) );
  NAND2_X1 U4601 ( .A1(n12672), .A2(n12654), .ZN(n30598) );
  NAND2_X1 U923 ( .A1(n6335), .A2(n442), .ZN(n11738) );
  OAI21_X1 U17496 ( .A1(n13340), .A2(n32019), .B(n17453), .ZN(n13342) );
  INV_X1 U869 ( .I(n25598), .ZN(n20515) );
  BUF_X2 U5312 ( .I(n20627), .Z(n16677) );
  INV_X1 U1395 ( .I(n2799), .ZN(n32085) );
  INV_X1 U21048 ( .I(n31669), .ZN(n14413) );
  NOR2_X1 U12377 ( .A1(n4664), .A2(n833), .ZN(n17472) );
  INV_X2 U6913 ( .I(n6300), .ZN(n12629) );
  INV_X1 U9584 ( .I(n11496), .ZN(n1256) );
  NAND2_X1 U14638 ( .A1(n3602), .A2(n33491), .ZN(n20746) );
  OAI21_X1 U30114 ( .A1(n34755), .A2(n3602), .B(n9815), .ZN(n17305) );
  NAND3_X1 U16478 ( .A1(n4467), .A2(n33268), .A3(n25361), .ZN(n4464) );
  NAND2_X1 U24878 ( .A1(n12309), .A2(n25574), .ZN(n18029) );
  OAI21_X1 U23218 ( .A1(n1543), .A2(n38178), .B(n7853), .ZN(n25342) );
  NAND2_X1 U12317 ( .A1(n11873), .A2(n1249), .ZN(n11549) );
  OAI21_X1 U786 ( .A1(n16316), .A2(n5455), .B(n6894), .ZN(n5454) );
  NAND2_X1 U16343 ( .A1(n541), .A2(n25620), .ZN(n11550) );
  NOR2_X1 U21721 ( .A1(n25620), .A2(n541), .ZN(n9602) );
  INV_X1 U6887 ( .I(n6448), .ZN(n20121) );
  INV_X1 U6559 ( .I(n4603), .ZN(n25688) );
  INV_X1 U6580 ( .I(n19589), .ZN(n20856) );
  AOI22_X1 U9498 ( .A1(n4664), .A2(n4047), .B1(n19637), .B2(n32419), .ZN(n4046) );
  NOR2_X1 U29066 ( .A1(n517), .A2(n16933), .ZN(n25547) );
  NAND2_X1 U18223 ( .A1(n9915), .A2(n25699), .ZN(n31707) );
  NAND3_X1 U14835 ( .A1(n14443), .A2(n25489), .A3(n38245), .ZN(n31820) );
  NAND2_X1 U29021 ( .A1(n25342), .A2(n12533), .ZN(n25343) );
  NAND2_X1 U12408 ( .A1(n25617), .A2(n25616), .ZN(n5248) );
  NAND2_X1 U9487 ( .A1(n7284), .A2(n7876), .ZN(n7875) );
  NAND2_X1 U12400 ( .A1(n12131), .A2(n32868), .ZN(n10313) );
  OAI21_X1 U8109 ( .A1(n25638), .A2(n25716), .B(n25637), .ZN(n18108) );
  NOR2_X1 U1223 ( .A1(n33491), .A2(n3602), .ZN(n31457) );
  NOR2_X1 U8132 ( .A1(n6573), .A2(n25416), .ZN(n14915) );
  AOI21_X1 U12358 ( .A1(n7875), .A2(n11495), .B(n1255), .ZN(n7874) );
  OAI21_X1 U8793 ( .A1(n25045), .A2(n17480), .B(n25467), .ZN(n30677) );
  INV_X2 U5597 ( .I(n4699), .ZN(n32747) );
  INV_X1 U1187 ( .I(n26020), .ZN(n31311) );
  INV_X2 U14300 ( .I(n31242), .ZN(n11834) );
  INV_X1 U9443 ( .I(n36922), .ZN(n26058) );
  NAND2_X1 U24887 ( .A1(n14793), .A2(n36226), .ZN(n18283) );
  NOR2_X1 U3475 ( .A1(n31192), .A2(n36546), .ZN(n2892) );
  CLKBUF_X2 U759 ( .I(n25956), .Z(n318) );
  INV_X2 U12202 ( .I(n25814), .ZN(n26131) );
  INV_X1 U5544 ( .I(n7660), .ZN(n11762) );
  OAI21_X1 U9402 ( .A1(n4602), .A2(n4516), .B(n929), .ZN(n12002) );
  OAI21_X1 U17281 ( .A1(n25928), .A2(n5356), .B(n30302), .ZN(n14774) );
  NAND2_X1 U12192 ( .A1(n1106), .A2(n14793), .ZN(n16432) );
  NOR2_X1 U1133 ( .A1(n25747), .A2(n1524), .ZN(n32782) );
  OAI21_X1 U8304 ( .A1(n2892), .A2(n2891), .B(n6390), .ZN(n30651) );
  NAND2_X1 U29102 ( .A1(n33348), .A2(n26020), .ZN(n25748) );
  OAI21_X1 U6837 ( .A1(n4382), .A2(n2625), .B(n25334), .ZN(n6105) );
  NAND2_X1 U2210 ( .A1(n16867), .A2(n25966), .ZN(n32333) );
  NAND2_X1 U2635 ( .A1(n6222), .A2(n6390), .ZN(n30546) );
  INV_X1 U2707 ( .I(n33909), .ZN(n26133) );
  INV_X2 U20195 ( .I(n15677), .ZN(n32052) );
  NOR2_X1 U23088 ( .A1(n19740), .A2(n11834), .ZN(n11624) );
  NOR2_X1 U9430 ( .A1(n25940), .A2(n1528), .ZN(n13524) );
  CLKBUF_X2 U8042 ( .I(n18176), .Z(n6578) );
  NAND2_X1 U662 ( .A1(n603), .A2(n25797), .ZN(n25911) );
  INV_X1 U6946 ( .I(n26093), .ZN(n931) );
  OAI22_X1 U15268 ( .A1(n10321), .A2(n25447), .B1(n17700), .B2(n31367), .ZN(
        n31831) );
  OAI21_X1 U12128 ( .A1(n13119), .A2(n25869), .B(n1017), .ZN(n13118) );
  NAND2_X1 U16062 ( .A1(n7961), .A2(n3575), .ZN(n25879) );
  OAI21_X1 U6824 ( .A1(n14573), .A2(n1106), .B(n25768), .ZN(n6103) );
  NOR2_X1 U17724 ( .A1(n13869), .A2(n446), .ZN(n12895) );
  AOI21_X1 U6843 ( .A1(n25993), .A2(n19740), .B(n12234), .ZN(n16397) );
  NAND2_X1 U4448 ( .A1(n3838), .A2(n21040), .ZN(n3837) );
  NAND2_X1 U669 ( .A1(n26065), .A2(n9530), .ZN(n26066) );
  NAND2_X1 U1028 ( .A1(n32109), .A2(n13732), .ZN(n5552) );
  INV_X1 U26122 ( .I(n9743), .ZN(n18002) );
  NOR2_X1 U7512 ( .A1(n32721), .A2(n30568), .ZN(n14286) );
  INV_X1 U12030 ( .I(n20600), .ZN(n7439) );
  NAND2_X1 U14563 ( .A1(n31654), .A2(n13391), .ZN(n13068) );
  INV_X1 U5664 ( .I(n26594), .ZN(n26484) );
  INV_X1 U7964 ( .I(n5848), .ZN(n26499) );
  INV_X1 U16652 ( .I(n7018), .ZN(n7028) );
  INV_X1 U3035 ( .I(n3781), .ZN(n19024) );
  INV_X1 U27261 ( .I(n18490), .ZN(n19217) );
  INV_X1 U637 ( .I(n5084), .ZN(n26588) );
  INV_X1 U12008 ( .I(n26334), .ZN(n8310) );
  INV_X2 U529 ( .I(n19951), .ZN(n1088) );
  BUF_X2 U20239 ( .I(n14347), .Z(n7527) );
  INV_X2 U6185 ( .I(n14962), .ZN(n13588) );
  NAND2_X1 U11805 ( .A1(n32168), .A2(n26970), .ZN(n17575) );
  INV_X1 U4526 ( .I(n37524), .ZN(n12549) );
  AOI21_X1 U2612 ( .A1(n14377), .A2(n19179), .B(n26811), .ZN(n26632) );
  INV_X1 U567 ( .I(n26665), .ZN(n26978) );
  NAND2_X1 U2763 ( .A1(n3369), .A2(n3368), .ZN(n30725) );
  NAND3_X1 U29296 ( .A1(n7978), .A2(n26703), .A3(n26702), .ZN(n26705) );
  NOR2_X1 U15959 ( .A1(n26934), .A2(n32745), .ZN(n4970) );
  NAND2_X1 U24655 ( .A1(n26952), .A2(n37055), .ZN(n15251) );
  OAI21_X1 U20942 ( .A1(n4138), .A2(n20699), .B(n26797), .ZN(n18792) );
  NOR2_X1 U27600 ( .A1(n7527), .A2(n35967), .ZN(n26628) );
  NAND2_X1 U18949 ( .A1(n6190), .A2(n26265), .ZN(n26266) );
  NOR2_X1 U9261 ( .A1(n14382), .A2(n10355), .ZN(n7392) );
  NOR2_X1 U29309 ( .A1(n13393), .A2(n26918), .ZN(n26766) );
  NOR2_X1 U30166 ( .A1(n26841), .A2(n20578), .ZN(n11708) );
  NAND2_X1 U2616 ( .A1(n19179), .A2(n12755), .ZN(n31647) );
  INV_X2 U7954 ( .I(n14355), .ZN(n26722) );
  BUF_X2 U4394 ( .I(n14459), .Z(n32797) );
  NAND2_X1 U15824 ( .A1(n19700), .A2(n14459), .ZN(n26691) );
  NAND2_X1 U856 ( .A1(n20575), .A2(n26612), .ZN(n11387) );
  AOI21_X1 U6766 ( .A1(n4138), .A2(n7516), .B(n26797), .ZN(n9764) );
  NOR2_X1 U24647 ( .A1(n38577), .A2(n6615), .ZN(n17785) );
  NAND2_X1 U11853 ( .A1(n26663), .A2(n15825), .ZN(n7005) );
  NAND2_X1 U9271 ( .A1(n33333), .A2(n26932), .ZN(n6605) );
  OAI21_X1 U6758 ( .A1(n20882), .A2(n26815), .B(n1497), .ZN(n18311) );
  NOR2_X1 U24956 ( .A1(n26803), .A2(n15594), .ZN(n19505) );
  NAND2_X1 U21006 ( .A1(n17237), .A2(n31526), .ZN(n8465) );
  NOR2_X1 U6833 ( .A1(n5480), .A2(n5481), .ZN(n5479) );
  NAND2_X1 U6171 ( .A1(n15763), .A2(n26975), .ZN(n19694) );
  OR2_X1 U29262 ( .A1(n26930), .A2(n26564), .Z(n26581) );
  INV_X2 U749 ( .I(n9956), .ZN(n27198) );
  INV_X2 U489 ( .I(n1487), .ZN(n27406) );
  INV_X1 U5884 ( .I(n3092), .ZN(n27401) );
  INV_X1 U7828 ( .I(n27449), .ZN(n27263) );
  INV_X1 U27417 ( .I(n27283), .ZN(n33254) );
  AOI21_X1 U7126 ( .A1(n27387), .A2(n35299), .B(n39826), .ZN(n30542) );
  INV_X1 U27373 ( .I(n27211), .ZN(n20092) );
  INV_X1 U1560 ( .I(n27397), .ZN(n2520) );
  BUF_X2 U4348 ( .I(n9956), .Z(n9201) );
  NAND2_X1 U9216 ( .A1(n27395), .A2(n9956), .ZN(n11805) );
  NAND2_X1 U29373 ( .A1(n27298), .A2(n27378), .ZN(n27171) );
  OAI21_X1 U24965 ( .A1(n27391), .A2(n35895), .B(n13699), .ZN(n18250) );
  NOR2_X1 U24381 ( .A1(n27438), .A2(n34977), .ZN(n14764) );
  OAI21_X1 U9172 ( .A1(n30986), .A2(n10051), .B(n12156), .ZN(n9454) );
  NAND2_X1 U10657 ( .A1(n15360), .A2(n1000), .ZN(n30840) );
  INV_X1 U425 ( .I(n27181), .ZN(n7418) );
  INV_X2 U6162 ( .I(n27484), .ZN(n11039) );
  NAND2_X1 U29344 ( .A1(n27358), .A2(n15360), .ZN(n27020) );
  NOR2_X1 U24563 ( .A1(n2949), .A2(n7606), .ZN(n32852) );
  NAND2_X1 U9203 ( .A1(n38060), .A2(n12485), .ZN(n27207) );
  NAND3_X1 U25253 ( .A1(n13471), .A2(n27199), .A3(n27198), .ZN(n26914) );
  NAND2_X1 U11507 ( .A1(n13793), .A2(n35897), .ZN(n13792) );
  NAND2_X1 U27576 ( .A1(n26999), .A2(n27054), .ZN(n19802) );
  NOR2_X1 U29361 ( .A1(n36911), .A2(n27455), .ZN(n27103) );
  AOI22_X1 U15938 ( .A1(n27055), .A2(n31672), .B1(n1475), .B2(n3466), .ZN(
        n3467) );
  NAND2_X1 U7762 ( .A1(n19077), .A2(n27265), .ZN(n18986) );
  NAND3_X1 U26138 ( .A1(n27154), .A2(n5311), .A3(n27406), .ZN(n26789) );
  INV_X2 U6733 ( .I(n2760), .ZN(n27388) );
  NAND2_X1 U17194 ( .A1(n7231), .A2(n27181), .ZN(n7230) );
  NAND2_X1 U14825 ( .A1(n14261), .A2(n38900), .ZN(n27559) );
  NAND2_X1 U15365 ( .A1(n15276), .A2(n36969), .ZN(n15275) );
  AOI22_X1 U5525 ( .A1(n11039), .A2(n11038), .B1(n27401), .B2(n11043), .ZN(
        n11037) );
  INV_X1 U2607 ( .I(n27735), .ZN(n27596) );
  INV_X1 U3501 ( .I(n5899), .ZN(n6990) );
  INV_X1 U16402 ( .I(n1455), .ZN(n20184) );
  NAND3_X1 U298 ( .A1(n28032), .A2(n8149), .A3(n1204), .ZN(n9663) );
  NAND2_X1 U25464 ( .A1(n989), .A2(n1069), .ZN(n14640) );
  INV_X2 U15718 ( .I(n11512), .ZN(n31942) );
  INV_X1 U14315 ( .I(n28093), .ZN(n16950) );
  AND2_X1 U12457 ( .A1(n33958), .A2(n19764), .Z(n28148) );
  NOR2_X1 U9092 ( .A1(n17032), .A2(n28267), .ZN(n3231) );
  NAND2_X1 U310 ( .A1(n3158), .A2(n28248), .ZN(n28251) );
  OAI21_X1 U3904 ( .A1(n33185), .A2(n16987), .B(n1071), .ZN(n30991) );
  NAND3_X1 U24111 ( .A1(n1442), .A2(n28054), .A3(n1205), .ZN(n13696) );
  NAND2_X1 U11286 ( .A1(n28035), .A2(n7310), .ZN(n13599) );
  NOR2_X1 U7625 ( .A1(n27934), .A2(n19435), .ZN(n10228) );
  OAI21_X1 U24995 ( .A1(n28193), .A2(n28194), .B(n27866), .ZN(n27906) );
  NAND2_X1 U24673 ( .A1(n17197), .A2(n17598), .ZN(n27930) );
  NOR2_X1 U30544 ( .A1(n18665), .A2(n28266), .ZN(n33912) );
  NAND2_X1 U11339 ( .A1(n17390), .A2(n28290), .ZN(n7190) );
  INV_X1 U7685 ( .I(n28267), .ZN(n20519) );
  INV_X1 U5395 ( .I(n14562), .ZN(n28265) );
  INV_X1 U21482 ( .I(n28152), .ZN(n9169) );
  AOI21_X1 U4015 ( .A1(n36844), .A2(n28248), .B(n37451), .ZN(n12531) );
  NOR2_X1 U15473 ( .A1(n33307), .A2(n28025), .ZN(n20967) );
  NAND2_X1 U7661 ( .A1(n5403), .A2(n21160), .ZN(n3843) );
  NAND3_X1 U7633 ( .A1(n28085), .A2(n6643), .A3(n989), .ZN(n28086) );
  NAND3_X1 U23235 ( .A1(n28283), .A2(n28067), .A3(n7528), .ZN(n32778) );
  OAI22_X1 U11250 ( .A1(n27929), .A2(n3511), .B1(n28193), .B2(n27930), .ZN(
        n5706) );
  NAND2_X1 U16910 ( .A1(n28024), .A2(n4803), .ZN(n27666) );
  NAND3_X1 U17699 ( .A1(n28251), .A2(n21223), .A3(n28249), .ZN(n31606) );
  OR2_X1 U3569 ( .A1(n15727), .A2(n28220), .Z(n11648) );
  OAI21_X1 U19496 ( .A1(n6643), .A2(n18841), .B(n6777), .ZN(n27917) );
  OR2_X1 U6198 ( .A1(n28047), .A2(n3990), .Z(n30350) );
  OAI22_X1 U9068 ( .A1(n15694), .A2(n21137), .B1(n15695), .B2(n28193), .ZN(
        n4504) );
  AOI21_X1 U14109 ( .A1(n28266), .A2(n14562), .B(n28267), .ZN(n28176) );
  NAND2_X1 U6649 ( .A1(n28223), .A2(n2868), .ZN(n3069) );
  NOR2_X1 U5926 ( .A1(n10166), .A2(n33185), .ZN(n3533) );
  NOR2_X1 U8521 ( .A1(n27917), .A2(n1069), .ZN(n30980) );
  INV_X1 U254 ( .I(n27908), .ZN(n28299) );
  INV_X1 U6621 ( .I(n28713), .ZN(n1425) );
  CLKBUF_X2 U4209 ( .I(n5237), .Z(n33591) );
  INV_X1 U6117 ( .I(n11296), .ZN(n15022) );
  INV_X1 U5855 ( .I(n28537), .ZN(n28495) );
  INV_X1 U3239 ( .I(n34559), .ZN(n1187) );
  NAND2_X1 U11142 ( .A1(n10618), .A2(n5662), .ZN(n18089) );
  AOI21_X1 U11079 ( .A1(n8800), .A2(n28553), .B(n18984), .ZN(n2327) );
  INV_X1 U11064 ( .I(n13598), .ZN(n16308) );
  INV_X1 U25306 ( .I(n32575), .ZN(n16038) );
  NOR2_X1 U11015 ( .A1(n18018), .A2(n13563), .ZN(n28693) );
  INV_X1 U4164 ( .I(n18990), .ZN(n33107) );
  OAI21_X1 U7501 ( .A1(n8759), .A2(n39147), .B(n28440), .ZN(n9783) );
  NAND3_X1 U21119 ( .A1(n16398), .A2(n8714), .A3(n13151), .ZN(n33190) );
  INV_X1 U222 ( .I(n16107), .ZN(n28499) );
  OAI21_X1 U29633 ( .A1(n28685), .A2(n18871), .B(n39724), .ZN(n28586) );
  NAND2_X1 U10982 ( .A1(n28428), .A2(n28661), .ZN(n12797) );
  INV_X2 U6550 ( .I(n30055), .ZN(n1057) );
  NAND2_X1 U10844 ( .A1(n29937), .A2(n14557), .ZN(n6692) );
  BUF_X2 U2380 ( .I(n28414), .Z(n29699) );
  INV_X1 U101 ( .I(n29769), .ZN(n1063) );
  NAND2_X1 U8874 ( .A1(n29815), .A2(n14600), .ZN(n13573) );
  INV_X1 U10843 ( .I(n29581), .ZN(n20085) );
  NAND2_X1 U2910 ( .A1(n2296), .A2(n31667), .ZN(n894) );
  OAI21_X1 U26264 ( .A1(n12878), .A2(n14525), .B(n16828), .ZN(n33092) );
  INV_X1 U29800 ( .I(n16828), .ZN(n29382) );
  INV_X2 U2359 ( .I(n29454), .ZN(n17295) );
  NOR2_X1 U2574 ( .A1(n8919), .A2(n37060), .ZN(n14755) );
  INV_X1 U104 ( .I(n30195), .ZN(n33394) );
  NOR2_X1 U1843 ( .A1(n1182), .A2(n29195), .ZN(n8346) );
  NAND2_X1 U25863 ( .A1(n29776), .A2(n29781), .ZN(n16790) );
  INV_X1 U5582 ( .I(n30153), .ZN(n19480) );
  NAND2_X1 U78 ( .A1(n29211), .A2(n17225), .ZN(n30655) );
  NAND2_X1 U14718 ( .A1(n31296), .A2(n19909), .ZN(n10435) );
  INV_X1 U25333 ( .I(n14773), .ZN(n29316) );
  OAI21_X1 U5578 ( .A1(n32671), .A2(n14400), .B(n31095), .ZN(n15864) );
  NOR2_X1 U20647 ( .A1(n29892), .A2(n971), .ZN(n10832) );
  NOR2_X1 U15237 ( .A1(n36207), .A2(n30198), .ZN(n2768) );
  NAND3_X1 U68 ( .A1(n1401), .A2(n37100), .A3(n9733), .ZN(n29400) );
  NAND2_X1 U5575 ( .A1(n7164), .A2(n7163), .ZN(n13384) );
  INV_X1 U7373 ( .I(n29339), .ZN(n29318) );
  NOR2_X1 U2381 ( .A1(n30071), .A2(n4377), .ZN(n30070) );
  INV_X2 U27745 ( .I(n15643), .ZN(n30037) );
  INV_X1 U12 ( .I(n1391), .ZN(n20481) );
  AND2_X1 U16973 ( .A1(n8399), .A2(n18457), .Z(n31534) );
  OAI21_X1 U22922 ( .A1(n30107), .A2(n35186), .B(n12203), .ZN(n18483) );
  NOR2_X1 U5 ( .A1(n30127), .A2(n17193), .ZN(n34706) );
  NAND2_X1 U17 ( .A1(n30022), .A2(n30034), .ZN(n30003) );
  OR2_X1 U35 ( .A1(n4377), .A2(n4378), .Z(n6489) );
  INV_X1 U53 ( .I(n30259), .ZN(n32865) );
  NOR2_X1 U63 ( .A1(n11596), .A2(n11594), .ZN(n35185) );
  NOR2_X1 U90 ( .A1(n1400), .A2(n30161), .ZN(n36607) );
  OAI21_X1 U98 ( .A1(n19050), .A2(n6938), .B(n34344), .ZN(n34589) );
  NAND2_X1 U106 ( .A1(n29896), .A2(n21167), .ZN(n36402) );
  NAND2_X1 U114 ( .A1(n482), .A2(n1181), .ZN(n36022) );
  NAND3_X1 U121 ( .A1(n7207), .A2(n12940), .A3(n29262), .ZN(n32189) );
  NOR2_X1 U132 ( .A1(n21287), .A2(n105), .ZN(n32498) );
  NAND2_X1 U147 ( .A1(n21270), .A2(n29586), .ZN(n34805) );
  NOR2_X1 U160 ( .A1(n37060), .A2(n20018), .ZN(n34761) );
  AND2_X1 U182 ( .A1(n16353), .A2(n20102), .Z(n34082) );
  INV_X1 U193 ( .I(n29643), .ZN(n34006) );
  INV_X1 U212 ( .I(n5289), .ZN(n36990) );
  AOI22_X1 U239 ( .A1(n2822), .A2(n30894), .B1(n16777), .B2(n28633), .ZN(
        n14929) );
  INV_X1 U240 ( .I(n34893), .ZN(n13422) );
  AND2_X1 U248 ( .A1(n11330), .A2(n39435), .Z(n12605) );
  OAI21_X1 U261 ( .A1(n36814), .A2(n16303), .B(n16304), .ZN(n28399) );
  NAND2_X1 U264 ( .A1(n36671), .A2(n1193), .ZN(n36567) );
  AND2_X1 U273 ( .A1(n35173), .A2(n28496), .Z(n34172) );
  NOR3_X1 U280 ( .A1(n36791), .A2(n15224), .A3(n13151), .ZN(n34893) );
  NAND2_X1 U289 ( .A1(n30894), .A2(n1190), .ZN(n28632) );
  OR2_X1 U292 ( .A1(n5418), .A2(n31015), .Z(n31077) );
  NAND2_X1 U295 ( .A1(n28505), .A2(n11164), .ZN(n34794) );
  NAND2_X1 U301 ( .A1(n31643), .A2(n34539), .ZN(n28467) );
  OR2_X1 U308 ( .A1(n17583), .A2(n5424), .Z(n30949) );
  NOR2_X1 U311 ( .A1(n28650), .A2(n18960), .ZN(n11469) );
  AOI21_X1 U320 ( .A1(n36993), .A2(n12653), .B(n15022), .ZN(n35935) );
  NAND3_X1 U323 ( .A1(n30716), .A2(n1420), .A3(n314), .ZN(n36124) );
  OR2_X1 U350 ( .A1(n31871), .A2(n6713), .Z(n35182) );
  BUF_X2 U363 ( .I(n28713), .Z(n36671) );
  NAND2_X1 U367 ( .A1(n30894), .A2(n28669), .ZN(n36993) );
  NAND2_X1 U388 ( .A1(n28544), .A2(n13133), .ZN(n34539) );
  NAND2_X1 U389 ( .A1(n32575), .A2(n36320), .ZN(n6819) );
  NAND2_X1 U402 ( .A1(n33707), .A2(n28695), .ZN(n10305) );
  NAND2_X1 U423 ( .A1(n1424), .A2(n36791), .ZN(n15235) );
  NAND2_X1 U431 ( .A1(n28724), .A2(n28723), .ZN(n18814) );
  NAND3_X1 U444 ( .A1(n33002), .A2(n889), .A3(n16325), .ZN(n34832) );
  NAND3_X1 U451 ( .A1(n35659), .A2(n35658), .A3(n35657), .ZN(n36236) );
  OAI21_X1 U458 ( .A1(n34442), .A2(n34441), .B(n20519), .ZN(n35570) );
  NAND2_X1 U472 ( .A1(n8232), .A2(n28224), .ZN(n35658) );
  AOI22_X1 U480 ( .A1(n12723), .A2(n3990), .B1(n28256), .B2(n28172), .ZN(
        n36936) );
  NAND2_X1 U483 ( .A1(n28151), .A2(n28152), .ZN(n37015) );
  INV_X1 U488 ( .I(n5239), .ZN(n19280) );
  OAI21_X1 U491 ( .A1(n28165), .A2(n37057), .B(n28274), .ZN(n36052) );
  NOR2_X1 U493 ( .A1(n15704), .A2(n33931), .ZN(n36689) );
  AND2_X1 U494 ( .A1(n17410), .A2(n28165), .Z(n34028) );
  NAND2_X1 U496 ( .A1(n34948), .A2(n34949), .ZN(n34470) );
  INV_X1 U499 ( .I(n4809), .ZN(n34442) );
  NOR2_X1 U520 ( .A1(n9514), .A2(n1438), .ZN(n28206) );
  AOI21_X1 U531 ( .A1(n28163), .A2(n7690), .B(n27979), .ZN(n6236) );
  NAND2_X1 U556 ( .A1(n28156), .A2(n28290), .ZN(n34186) );
  NOR2_X1 U564 ( .A1(n28290), .A2(n877), .ZN(n16513) );
  OR2_X1 U583 ( .A1(n988), .A2(n14399), .Z(n34069) );
  NAND2_X1 U597 ( .A1(n28260), .A2(n34410), .ZN(n34948) );
  BUF_X2 U602 ( .I(n21126), .Z(n13714) );
  AND2_X1 U617 ( .A1(n1445), .A2(n35225), .Z(n20188) );
  NOR2_X1 U630 ( .A1(n1204), .A2(n33656), .ZN(n18044) );
  NAND2_X1 U632 ( .A1(n4457), .A2(n14389), .ZN(n18530) );
  INV_X1 U661 ( .I(n27792), .ZN(n34812) );
  INV_X1 U670 ( .I(n27657), .ZN(n35853) );
  INV_X1 U673 ( .I(n27829), .ZN(n34531) );
  INV_X1 U681 ( .I(n9013), .ZN(n1464) );
  NOR2_X1 U683 ( .A1(n36234), .A2(n20740), .ZN(n15984) );
  NAND2_X1 U685 ( .A1(n4105), .A2(n4104), .ZN(n9739) );
  AND2_X1 U688 ( .A1(n34769), .A2(n27165), .Z(n18768) );
  OR2_X1 U690 ( .A1(n27403), .A2(n36865), .Z(n34111) );
  OR2_X1 U692 ( .A1(n27372), .A2(n37890), .Z(n27373) );
  NOR2_X1 U697 ( .A1(n35825), .A2(n33146), .ZN(n34777) );
  NAND2_X1 U702 ( .A1(n2306), .A2(n1891), .ZN(n34811) );
  AND2_X1 U703 ( .A1(n35904), .A2(n27284), .Z(n19570) );
  INV_X1 U726 ( .I(n36200), .ZN(n27311) );
  AND2_X1 U740 ( .A1(n9369), .A2(n30986), .Z(n18489) );
  CLKBUF_X1 U741 ( .I(n27383), .Z(n33336) );
  AND2_X1 U742 ( .A1(n6686), .A2(n11729), .Z(n27231) );
  NAND2_X1 U745 ( .A1(n27364), .A2(n5772), .ZN(n36073) );
  NAND3_X1 U751 ( .A1(n27131), .A2(n27343), .A3(n36183), .ZN(n26999) );
  AOI21_X1 U758 ( .A1(n39305), .A2(n33893), .B(n16043), .ZN(n34705) );
  AND2_X1 U779 ( .A1(n19477), .A2(n27349), .Z(n30429) );
  NOR2_X1 U795 ( .A1(n995), .A2(n1226), .ZN(n13266) );
  AOI21_X1 U820 ( .A1(n18246), .A2(n33773), .B(n27416), .ZN(n33235) );
  AND2_X1 U831 ( .A1(n10171), .A2(n27583), .Z(n8698) );
  INV_X1 U834 ( .I(n27284), .ZN(n1084) );
  NOR2_X1 U837 ( .A1(n27137), .A2(n8798), .ZN(n18652) );
  NAND2_X1 U859 ( .A1(n32602), .A2(n7978), .ZN(n36243) );
  NAND3_X1 U917 ( .A1(n35489), .A2(n34058), .A3(n1088), .ZN(n26657) );
  OR2_X1 U920 ( .A1(n26961), .A2(n20936), .Z(n8650) );
  AND2_X1 U921 ( .A1(n13111), .A2(n19364), .Z(n34071) );
  NAND2_X1 U935 ( .A1(n33302), .A2(n26619), .ZN(n36589) );
  NAND2_X1 U944 ( .A1(n3825), .A2(n11226), .ZN(n4195) );
  NAND3_X1 U961 ( .A1(n2100), .A2(n2101), .A3(n4211), .ZN(n30715) );
  NOR2_X1 U982 ( .A1(n20573), .A2(n17237), .ZN(n11709) );
  OR2_X1 U983 ( .A1(n26703), .A2(n10440), .Z(n34058) );
  NOR2_X1 U995 ( .A1(n3825), .A2(n11138), .ZN(n15314) );
  OAI21_X1 U1000 ( .A1(n26852), .A2(n14453), .B(n5537), .ZN(n35612) );
  AND2_X1 U1002 ( .A1(n26876), .A2(n14455), .Z(n2081) );
  INV_X1 U1009 ( .I(n26824), .ZN(n26424) );
  NAND2_X1 U1010 ( .A1(n18903), .A2(n19615), .ZN(n18902) );
  NOR2_X1 U1012 ( .A1(n26878), .A2(n26879), .ZN(n3369) );
  INV_X2 U1013 ( .I(n26619), .ZN(n26951) );
  CLKBUF_X2 U1019 ( .I(n26666), .Z(n19449) );
  NAND2_X1 U1026 ( .A1(n26849), .A2(n10314), .ZN(n34908) );
  OR2_X1 U1027 ( .A1(n13605), .A2(n5869), .Z(n4410) );
  AND2_X1 U1031 ( .A1(n26961), .A2(n35259), .Z(n34075) );
  CLKBUF_X2 U1067 ( .I(n26931), .Z(n19222) );
  OR2_X1 U1069 ( .A1(n32623), .A2(n15386), .Z(n26671) );
  BUF_X2 U1084 ( .I(n19436), .Z(n13111) );
  INV_X1 U1091 ( .I(n18012), .ZN(n33551) );
  OAI21_X1 U1103 ( .A1(n11386), .A2(n7260), .B(n33030), .ZN(n35240) );
  NAND2_X1 U1142 ( .A1(n16397), .A2(n25994), .ZN(n36951) );
  AND2_X1 U1153 ( .A1(n2561), .A2(n2029), .Z(n25846) );
  NAND2_X1 U1157 ( .A1(n15677), .A2(n36666), .ZN(n36665) );
  NAND2_X1 U1160 ( .A1(n18176), .A2(n25348), .ZN(n35891) );
  AND2_X1 U1167 ( .A1(n25742), .A2(n25770), .Z(n34018) );
  OR2_X1 U1173 ( .A1(n2865), .A2(n3642), .Z(n25926) );
  NAND3_X1 U1183 ( .A1(n586), .A2(n1020), .A3(n26018), .ZN(n15966) );
  NAND3_X1 U1201 ( .A1(n26121), .A2(n26123), .A3(n26122), .ZN(n8133) );
  NOR2_X1 U1202 ( .A1(n25945), .A2(n31523), .ZN(n26331) );
  NOR2_X1 U1203 ( .A1(n11834), .A2(n25956), .ZN(n34573) );
  OR2_X1 U1204 ( .A1(n26015), .A2(n31719), .Z(n12457) );
  NAND3_X1 U1235 ( .A1(n18283), .A2(n18282), .A3(n3356), .ZN(n18426) );
  AND2_X1 U1246 ( .A1(n33258), .A2(n26093), .Z(n8005) );
  NAND2_X1 U1250 ( .A1(n26070), .A2(n34685), .ZN(n15795) );
  OR2_X1 U1278 ( .A1(n9916), .A2(n26134), .Z(n32843) );
  INV_X1 U1298 ( .I(n834), .ZN(n36906) );
  NAND2_X1 U1315 ( .A1(n36451), .A2(n36449), .ZN(n17372) );
  NOR3_X1 U1335 ( .A1(n17915), .A2(n8481), .A3(n7767), .ZN(n8480) );
  CLKBUF_X4 U1357 ( .I(n35138), .Z(n365) );
  BUF_X4 U1385 ( .I(n25951), .Z(n34217) );
  OAI21_X1 U1398 ( .A1(n25525), .A2(n25526), .B(n517), .ZN(n25530) );
  OAI21_X1 U1411 ( .A1(n36941), .A2(n36940), .B(n19095), .ZN(n13210) );
  OAI21_X1 U1431 ( .A1(n35171), .A2(n25699), .B(n31721), .ZN(n24957) );
  NOR2_X1 U1437 ( .A1(n1536), .A2(n12368), .ZN(n35660) );
  NAND2_X1 U1438 ( .A1(n35763), .A2(n11550), .ZN(n11544) );
  INV_X1 U1459 ( .I(n7391), .ZN(n36411) );
  AND2_X1 U1462 ( .A1(n611), .A2(n25328), .Z(n14631) );
  OR2_X1 U1494 ( .A1(n14410), .A2(n6731), .Z(n34078) );
  NOR2_X1 U1501 ( .A1(n6300), .A2(n33495), .ZN(n34487) );
  NOR2_X1 U1503 ( .A1(n39599), .A2(n37993), .ZN(n25638) );
  NAND2_X1 U1510 ( .A1(n6731), .A2(n37051), .ZN(n35349) );
  NAND2_X1 U1515 ( .A1(n25603), .A2(n21302), .ZN(n25605) );
  NAND2_X1 U1543 ( .A1(n25462), .A2(n36133), .ZN(n36132) );
  CLKBUF_X2 U1588 ( .I(n25631), .Z(n5051) );
  NOR2_X1 U1589 ( .A1(n19548), .A2(n5050), .ZN(n25393) );
  AND2_X1 U1590 ( .A1(n13460), .A2(n25422), .Z(n34081) );
  NOR2_X1 U1596 ( .A1(n14708), .A2(n15541), .ZN(n36487) );
  OR2_X1 U1601 ( .A1(n33950), .A2(n25692), .Z(n12780) );
  INV_X1 U1603 ( .I(n15172), .ZN(n36524) );
  NOR2_X1 U1607 ( .A1(n25484), .A2(n3985), .ZN(n36135) );
  INV_X1 U1609 ( .I(n25486), .ZN(n19829) );
  OAI21_X1 U1622 ( .A1(n12533), .A2(n31010), .B(n14436), .ZN(n8034) );
  NAND2_X1 U1624 ( .A1(n841), .A2(n18164), .ZN(n9800) );
  NOR2_X1 U1626 ( .A1(n20888), .A2(n25614), .ZN(n10034) );
  CLKBUF_X1 U1630 ( .I(n14481), .Z(n36086) );
  NOR2_X1 U1634 ( .A1(n20515), .A2(n3602), .ZN(n25068) );
  AND2_X1 U1635 ( .A1(n252), .A2(n16931), .Z(n25495) );
  CLKBUF_X1 U1670 ( .I(n20153), .Z(n32904) );
  BUF_X2 U1674 ( .I(n25490), .Z(n25620) );
  INV_X1 U1723 ( .I(n8542), .ZN(n5434) );
  NOR2_X1 U1771 ( .A1(n13518), .A2(n8264), .ZN(n36786) );
  AND2_X1 U1774 ( .A1(n24728), .A2(n3510), .Z(n20180) );
  OR2_X1 U1783 ( .A1(n24900), .A2(n19279), .Z(n30419) );
  NOR2_X1 U1795 ( .A1(n24646), .A2(n24794), .ZN(n18570) );
  NOR2_X1 U1798 ( .A1(n24605), .A2(n24774), .ZN(n31122) );
  NOR2_X1 U1804 ( .A1(n24669), .A2(n24668), .ZN(n36787) );
  INV_X1 U1807 ( .I(n24749), .ZN(n24751) );
  AND2_X1 U1809 ( .A1(n24683), .A2(n36058), .Z(n18056) );
  CLKBUF_X2 U1813 ( .I(n36058), .Z(n35801) );
  OR2_X1 U1823 ( .A1(n16841), .A2(n24799), .Z(n11942) );
  NAND3_X1 U1828 ( .A1(n259), .A2(n24630), .A3(n24826), .ZN(n37017) );
  NOR2_X1 U1836 ( .A1(n24828), .A2(n9218), .ZN(n24816) );
  AND2_X1 U1853 ( .A1(n24416), .A2(n17351), .Z(n24507) );
  NAND2_X1 U1869 ( .A1(n9478), .A2(n34796), .ZN(n34904) );
  INV_X2 U1877 ( .I(n15332), .ZN(n33344) );
  OAI21_X1 U1878 ( .A1(n34039), .A2(n19566), .B(n34384), .ZN(n24324) );
  NAND2_X1 U1882 ( .A1(n31519), .A2(n24784), .ZN(n24613) );
  AND2_X1 U1895 ( .A1(n1600), .A2(n19782), .Z(n34039) );
  OAI21_X1 U1898 ( .A1(n33379), .A2(n13653), .B(n19566), .ZN(n34384) );
  OR2_X1 U1899 ( .A1(n39196), .A2(n24805), .Z(n24532) );
  INV_X1 U1901 ( .I(n24819), .ZN(n1565) );
  OAI21_X1 U1902 ( .A1(n24630), .A2(n9218), .B(n24826), .ZN(n34796) );
  NOR2_X1 U1903 ( .A1(n9197), .A2(n24879), .ZN(n35048) );
  NAND2_X1 U1926 ( .A1(n24819), .A2(n8646), .ZN(n14166) );
  NOR2_X1 U1929 ( .A1(n39818), .A2(n34758), .ZN(n34420) );
  NOR2_X1 U1937 ( .A1(n19653), .A2(n35712), .ZN(n35840) );
  NOR2_X1 U1950 ( .A1(n3133), .A2(n12953), .ZN(n36273) );
  NOR2_X1 U1953 ( .A1(n35150), .A2(n5855), .ZN(n5854) );
  NOR3_X1 U1964 ( .A1(n1125), .A2(n31452), .A3(n6515), .ZN(n35086) );
  NAND2_X1 U1983 ( .A1(n24459), .A2(n24457), .ZN(n36157) );
  NOR2_X1 U1993 ( .A1(n19782), .A2(n1600), .ZN(n35872) );
  CLKBUF_X1 U2001 ( .I(n23819), .Z(n35712) );
  CLKBUF_X2 U2002 ( .I(n16459), .Z(n609) );
  BUF_X2 U2004 ( .I(n24142), .Z(n36757) );
  NAND2_X1 U2013 ( .A1(n14491), .A2(n1605), .ZN(n35004) );
  NOR3_X1 U2014 ( .A1(n24443), .A2(n253), .A3(n30833), .ZN(n35815) );
  NAND2_X1 U2053 ( .A1(n24158), .A2(n1280), .ZN(n31852) );
  AND2_X1 U2060 ( .A1(n32899), .A2(n9193), .Z(n31490) );
  NOR2_X1 U2069 ( .A1(n6465), .A2(n1275), .ZN(n36622) );
  NOR2_X1 U2073 ( .A1(n19584), .A2(n24419), .ZN(n35814) );
  CLKBUF_X2 U2091 ( .I(n36500), .Z(n35761) );
  AND2_X1 U2095 ( .A1(n18302), .A2(n14378), .Z(n34074) );
  NAND2_X1 U2101 ( .A1(n1606), .A2(n24245), .ZN(n14662) );
  AND2_X1 U2113 ( .A1(n33057), .A2(n24104), .Z(n24331) );
  NOR2_X1 U2121 ( .A1(n24169), .A2(n277), .ZN(n34655) );
  BUF_X2 U2125 ( .I(n24308), .Z(n19745) );
  BUF_X2 U2128 ( .I(n24317), .Z(n19782) );
  INV_X1 U2147 ( .I(n23912), .ZN(n23957) );
  OAI21_X1 U2154 ( .A1(n34337), .A2(n34336), .B(n23560), .ZN(n14354) );
  AOI21_X1 U2160 ( .A1(n1301), .A2(n33316), .B(n23444), .ZN(n10989) );
  OR2_X1 U2162 ( .A1(n10143), .A2(n39401), .Z(n7819) );
  NAND2_X1 U2175 ( .A1(n34602), .A2(n36129), .ZN(n35355) );
  NAND3_X1 U2176 ( .A1(n37774), .A2(n23602), .A3(n35664), .ZN(n30276) );
  NAND2_X1 U2190 ( .A1(n35974), .A2(n35536), .ZN(n430) );
  AOI21_X1 U2202 ( .A1(n23522), .A2(n23521), .B(n36219), .ZN(n19227) );
  OAI21_X1 U2203 ( .A1(n3309), .A2(n5591), .B(n34635), .ZN(n3745) );
  OAI21_X1 U2205 ( .A1(n11468), .A2(n12851), .B(n15122), .ZN(n12982) );
  NOR2_X1 U2207 ( .A1(n35938), .A2(n7335), .ZN(n34337) );
  NAND3_X1 U2223 ( .A1(n35892), .A2(n23641), .A3(n1310), .ZN(n9609) );
  AOI21_X1 U2225 ( .A1(n11453), .A2(n23746), .B(n960), .ZN(n6910) );
  INV_X2 U2243 ( .I(n35331), .ZN(n23444) );
  NOR2_X1 U2261 ( .A1(n33840), .A2(n34506), .ZN(n2681) );
  NAND2_X1 U2263 ( .A1(n23494), .A2(n4147), .ZN(n36129) );
  OR2_X1 U2299 ( .A1(n33747), .A2(n35367), .Z(n23383) );
  BUF_X2 U2301 ( .I(n3496), .Z(n35938) );
  INV_X1 U2321 ( .I(n13038), .ZN(n35501) );
  OR2_X1 U2327 ( .A1(n8757), .A2(n19005), .Z(n34068) );
  NAND3_X1 U2334 ( .A1(n32032), .A2(n36185), .A3(n36184), .ZN(n11473) );
  NOR2_X1 U2336 ( .A1(n36422), .A2(n32515), .ZN(n34696) );
  INV_X1 U2341 ( .I(n33544), .ZN(n35955) );
  NAND2_X1 U2344 ( .A1(n34713), .A2(n1044), .ZN(n10553) );
  NOR2_X1 U2364 ( .A1(n19524), .A2(n22900), .ZN(n34401) );
  NAND2_X1 U2372 ( .A1(n19586), .A2(n23084), .ZN(n23186) );
  NOR2_X1 U2382 ( .A1(n1314), .A2(n23084), .ZN(n9769) );
  NOR3_X1 U2396 ( .A1(n14089), .A2(n1046), .A3(n20267), .ZN(n4773) );
  NAND2_X1 U2400 ( .A1(n22899), .A2(n23201), .ZN(n36638) );
  NAND2_X1 U2402 ( .A1(n32515), .A2(n33925), .ZN(n13945) );
  INV_X1 U2408 ( .I(n1831), .ZN(n35288) );
  INV_X1 U2410 ( .I(n5581), .ZN(n35591) );
  CLKBUF_X2 U2412 ( .I(n19966), .Z(n35918) );
  CLKBUF_X2 U2415 ( .I(n23122), .Z(n19351) );
  BUF_X2 U2434 ( .I(n13587), .Z(n1763) );
  NOR2_X1 U2440 ( .A1(n23165), .A2(n36554), .ZN(n36553) );
  INV_X1 U2456 ( .I(n12961), .ZN(n14439) );
  INV_X1 U2464 ( .I(n22443), .ZN(n35848) );
  NAND2_X1 U2473 ( .A1(n36466), .A2(n1329), .ZN(n7867) );
  INV_X1 U2476 ( .I(n19328), .ZN(n22687) );
  INV_X1 U2481 ( .I(n22665), .ZN(n34545) );
  AND2_X1 U2489 ( .A1(n2765), .A2(n34808), .Z(n2435) );
  INV_X1 U2495 ( .I(n37217), .ZN(n34015) );
  NAND2_X1 U2502 ( .A1(n22390), .A2(n19873), .ZN(n13778) );
  OR2_X1 U2506 ( .A1(n19655), .A2(n22160), .Z(n34023) );
  NAND3_X1 U2510 ( .A1(n22246), .A2(n33571), .A3(n20889), .ZN(n19080) );
  OAI21_X1 U2511 ( .A1(n22344), .A2(n21987), .B(n22341), .ZN(n1838) );
  INV_X1 U2521 ( .I(n3863), .ZN(n35822) );
  NAND2_X1 U2528 ( .A1(n22282), .A2(n22130), .ZN(n21963) );
  INV_X2 U2535 ( .I(n20376), .ZN(n36661) );
  AND2_X1 U2542 ( .A1(n9387), .A2(n22222), .Z(n19253) );
  INV_X1 U2543 ( .I(n15229), .ZN(n34925) );
  OR2_X1 U2546 ( .A1(n2765), .A2(n22243), .Z(n4864) );
  NAND2_X1 U2548 ( .A1(n22091), .A2(n19837), .ZN(n22097) );
  NOR2_X1 U2551 ( .A1(n22271), .A2(n22316), .ZN(n36139) );
  NAND2_X1 U2565 ( .A1(n1333), .A2(n18656), .ZN(n18730) );
  INV_X1 U2572 ( .I(n22067), .ZN(n36563) );
  NAND2_X1 U2575 ( .A1(n39489), .A2(n6947), .ZN(n6946) );
  NOR2_X2 U2582 ( .A1(n8442), .A2(n8440), .ZN(n22400) );
  NAND2_X1 U2588 ( .A1(n12927), .A2(n21932), .ZN(n16660) );
  AOI22_X1 U2593 ( .A1(n18742), .A2(n36519), .B1(n4084), .B2(n18710), .ZN(
        n35833) );
  OAI21_X1 U2596 ( .A1(n16163), .A2(n21601), .B(n17102), .ZN(n7551) );
  INV_X1 U2622 ( .I(n21743), .ZN(n17266) );
  AND2_X1 U2632 ( .A1(n12144), .A2(n1351), .Z(n12142) );
  NAND2_X1 U2634 ( .A1(n12332), .A2(n16305), .ZN(n35999) );
  INV_X1 U2636 ( .I(n21410), .ZN(n35043) );
  OAI22_X1 U2639 ( .A1(n21556), .A2(n19323), .B1(n21620), .B2(n18412), .ZN(
        n36353) );
  INV_X1 U2644 ( .I(n36062), .ZN(n14450) );
  NOR2_X1 U2649 ( .A1(n18710), .A2(n21630), .ZN(n21631) );
  INV_X1 U2653 ( .I(n21576), .ZN(n36781) );
  NOR2_X1 U2661 ( .A1(n21484), .A2(n21880), .ZN(n36780) );
  AND2_X1 U2673 ( .A1(n1454), .A2(n1206), .Z(n33981) );
  INV_X2 U2681 ( .I(n19658), .ZN(n24373) );
  BUF_X2 U2685 ( .I(n8219), .Z(n7866) );
  NAND2_X2 U2687 ( .A1(n19573), .A2(n4292), .ZN(n35454) );
  INV_X2 U2691 ( .I(n27882), .ZN(n28255) );
  NAND2_X2 U2704 ( .A1(n36685), .A2(n28677), .ZN(n28577) );
  NAND2_X2 U2708 ( .A1(n6075), .A2(n6077), .ZN(n32870) );
  BUF_X4 U2711 ( .I(n37378), .Z(n31626) );
  INV_X2 U2713 ( .I(n24759), .ZN(n14265) );
  NOR2_X2 U2722 ( .A1(n21583), .A2(n21893), .ZN(n21514) );
  OAI22_X2 U2724 ( .A1(n36673), .A2(n1578), .B1(n31213), .B2(n24799), .ZN(
        n8576) );
  OR2_X1 U2726 ( .A1(n33840), .A2(n14477), .Z(n2682) );
  OAI21_X1 U2741 ( .A1(n37783), .A2(n8149), .B(n28089), .ZN(n5403) );
  INV_X2 U2758 ( .I(n13151), .ZN(n1417) );
  AND2_X1 U2772 ( .A1(n8413), .A2(n11636), .Z(n11651) );
  NAND2_X1 U2783 ( .A1(n36348), .A2(n27974), .ZN(n27978) );
  AOI21_X1 U2793 ( .A1(n13081), .A2(n28273), .B(n10642), .ZN(n36348) );
  AOI21_X1 U2794 ( .A1(n29219), .A2(n31772), .B(n32209), .ZN(n122) );
  NAND2_X1 U2803 ( .A1(n6019), .A2(n9918), .ZN(n16490) );
  NAND3_X1 U2811 ( .A1(n18883), .A2(n28591), .A3(n306), .ZN(n15629) );
  NAND2_X1 U2837 ( .A1(n20274), .A2(n36421), .ZN(n36420) );
  NAND3_X1 U2841 ( .A1(n31120), .A2(n3818), .A3(n30076), .ZN(n34292) );
  NOR2_X1 U2848 ( .A1(n34592), .A2(n7637), .ZN(n9967) );
  NAND2_X1 U2849 ( .A1(n19884), .A2(n16874), .ZN(n29181) );
  OAI21_X1 U2856 ( .A1(n22149), .A2(n5821), .B(n18999), .ZN(n9124) );
  AOI22_X1 U2860 ( .A1(n32457), .A2(n8071), .B1(n20376), .B2(n1154), .ZN(n7212) );
  OR2_X1 U2861 ( .A1(n29884), .A2(n29883), .Z(n14540) );
  NAND2_X1 U2865 ( .A1(n8089), .A2(n14323), .ZN(n13616) );
  NOR2_X1 U2868 ( .A1(n20572), .A2(n38365), .ZN(n33725) );
  NOR2_X1 U2870 ( .A1(n38365), .A2(n20572), .ZN(n18013) );
  OAI21_X1 U2874 ( .A1(n15922), .A2(n20572), .B(n11166), .ZN(n11368) );
  NOR2_X1 U2882 ( .A1(n37040), .A2(n12685), .ZN(n14588) );
  NAND2_X1 U2887 ( .A1(n29635), .A2(n20290), .ZN(n20286) );
  NAND2_X1 U2892 ( .A1(n6001), .A2(n31772), .ZN(n36977) );
  NAND3_X1 U2905 ( .A1(n3818), .A2(n31120), .A3(n30077), .ZN(n30072) );
  NAND3_X1 U2913 ( .A1(n28723), .A2(n28724), .A3(n28722), .ZN(n18187) );
  INV_X2 U2957 ( .I(n20159), .ZN(n29409) );
  CLKBUF_X2 U2958 ( .I(n20159), .Z(n9790) );
  INV_X2 U2962 ( .I(n13545), .ZN(n2803) );
  NOR3_X1 U2972 ( .A1(n13446), .A2(n19007), .A3(n24403), .ZN(n7084) );
  NAND2_X1 U2973 ( .A1(n13446), .A2(n13555), .ZN(n34598) );
  AOI22_X1 U2975 ( .A1(n29400), .A2(n13850), .B1(n17849), .B2(n16260), .ZN(
        n29414) );
  NOR2_X1 U2982 ( .A1(n25481), .A2(n32026), .ZN(n25526) );
  NOR2_X1 U2984 ( .A1(n27887), .A2(n1454), .ZN(n33913) );
  NOR2_X1 U2986 ( .A1(n2989), .A2(n11361), .ZN(n3336) );
  NAND2_X1 U2998 ( .A1(n26780), .A2(n20223), .ZN(n32743) );
  NAND2_X1 U3001 ( .A1(n26780), .A2(n17712), .ZN(n35410) );
  CLKBUF_X4 U3009 ( .I(n23682), .Z(n1607) );
  NOR2_X1 U3010 ( .A1(n30003), .A2(n35103), .ZN(n35588) );
  AND2_X1 U3011 ( .A1(n19844), .A2(n28713), .Z(n8218) );
  NOR2_X1 U3028 ( .A1(n20274), .A2(n4768), .ZN(n34707) );
  NAND2_X1 U3029 ( .A1(n5270), .A2(n30032), .ZN(n30039) );
  OAI21_X1 U3030 ( .A1(n19458), .A2(n30042), .B(n30041), .ZN(n19884) );
  AOI21_X1 U3033 ( .A1(n24779), .A2(n16210), .B(n30421), .ZN(n3016) );
  NAND2_X1 U3071 ( .A1(n26578), .A2(n26564), .ZN(n26580) );
  NOR2_X1 U3085 ( .A1(n16889), .A2(n31532), .ZN(n12370) );
  AOI21_X1 U3102 ( .A1(n13014), .A2(n11981), .B(n29209), .ZN(n34592) );
  OR2_X1 U3108 ( .A1(n1404), .A2(n29592), .Z(n14433) );
  INV_X2 U3118 ( .I(n4945), .ZN(n27979) );
  NOR2_X1 U3137 ( .A1(n9751), .A2(n20359), .ZN(n14619) );
  NOR2_X1 U3143 ( .A1(n12829), .A2(n12876), .ZN(n29383) );
  NAND3_X1 U3144 ( .A1(n10422), .A2(n12876), .A3(n29310), .ZN(n29079) );
  NAND2_X1 U3167 ( .A1(n29367), .A2(n37095), .ZN(n19060) );
  NAND2_X1 U3173 ( .A1(n30117), .A2(n18829), .ZN(n12203) );
  OAI21_X1 U3179 ( .A1(n259), .A2(n33012), .B(n11081), .ZN(n11054) );
  NOR2_X1 U3184 ( .A1(n11081), .A2(n17986), .ZN(n11053) );
  NAND2_X1 U3185 ( .A1(n24826), .A2(n11081), .ZN(n14519) );
  NAND2_X1 U3189 ( .A1(n18743), .A2(n35051), .ZN(n12189) );
  NOR2_X1 U3194 ( .A1(n31557), .A2(n25689), .ZN(n36309) );
  NOR2_X1 U3202 ( .A1(n31557), .A2(n6448), .ZN(n25686) );
  NAND3_X1 U3206 ( .A1(n15038), .A2(n11628), .A3(n12218), .ZN(n27620) );
  NOR2_X1 U3215 ( .A1(n28012), .A2(n11628), .ZN(n15269) );
  OAI21_X1 U3219 ( .A1(n30128), .A2(n1385), .B(n10813), .ZN(n13298) );
  NAND2_X1 U3221 ( .A1(n1407), .A2(n31444), .ZN(n6202) );
  NOR2_X1 U3231 ( .A1(n1061), .A2(n14179), .ZN(n11410) );
  NAND2_X1 U3235 ( .A1(n9242), .A2(n20010), .ZN(n28150) );
  NOR2_X1 U3250 ( .A1(n14783), .A2(n20277), .ZN(n21472) );
  INV_X1 U3255 ( .I(n8605), .ZN(n14970) );
  NOR2_X1 U3263 ( .A1(n12717), .A2(n12718), .ZN(n33337) );
  INV_X1 U3268 ( .I(n19096), .ZN(n12442) );
  AOI21_X1 U3273 ( .A1(n2050), .A2(n14640), .B(n28222), .ZN(n436) );
  OAI22_X1 U3280 ( .A1(n16213), .A2(n21051), .B1(n7939), .B2(n23379), .ZN(
        n15969) );
  INV_X1 U3281 ( .I(n16213), .ZN(n35974) );
  CLKBUF_X1 U3283 ( .I(n18908), .Z(n34847) );
  OR2_X1 U3285 ( .A1(n25483), .A2(n25328), .Z(n18787) );
  AND2_X1 U3335 ( .A1(n19398), .A2(n25681), .Z(n30392) );
  BUF_X2 U3336 ( .I(n25395), .Z(n25681) );
  AOI21_X1 U3339 ( .A1(n31120), .A2(n30069), .B(n3815), .ZN(n19551) );
  NAND2_X1 U3340 ( .A1(n20535), .A2(n21869), .ZN(n9592) );
  NAND2_X1 U3341 ( .A1(n13594), .A2(n28680), .ZN(n28719) );
  NAND2_X1 U3369 ( .A1(n36996), .A2(n23165), .ZN(n22810) );
  NOR2_X1 U3383 ( .A1(n24473), .A2(n39074), .ZN(n24471) );
  AOI21_X1 U3386 ( .A1(n31494), .A2(n30484), .B(n288), .ZN(n5158) );
  NAND2_X1 U3397 ( .A1(n19366), .A2(n27969), .ZN(n18439) );
  NAND2_X1 U3406 ( .A1(n28048), .A2(n28255), .ZN(n34949) );
  NOR2_X1 U3413 ( .A1(n15518), .A2(n17477), .ZN(n36591) );
  INV_X1 U3415 ( .I(n15267), .ZN(n34618) );
  NOR3_X1 U3430 ( .A1(n5001), .A2(n21023), .A3(n8762), .ZN(n19747) );
  NAND3_X1 U3435 ( .A1(n32527), .A2(n15825), .A3(n31502), .ZN(n35436) );
  NOR3_X1 U3445 ( .A1(n31444), .A2(n14158), .A3(n19424), .ZN(n10605) );
  OR3_X2 U3449 ( .A1(n987), .A2(n1070), .A3(n7872), .Z(n16632) );
  INV_X2 U3477 ( .I(n29700), .ZN(n1060) );
  AOI21_X1 U3478 ( .A1(n1182), .A2(n5977), .B(n29700), .ZN(n20816) );
  CLKBUF_X2 U3480 ( .I(n29865), .Z(n33256) );
  AOI22_X1 U3504 ( .A1(n1398), .A2(n29701), .B1(n8941), .B2(n5977), .ZN(n8347)
         );
  NAND2_X1 U3510 ( .A1(n29430), .A2(n38051), .ZN(n29342) );
  NOR2_X1 U3517 ( .A1(n9677), .A2(n903), .ZN(n3410) );
  NAND2_X1 U3518 ( .A1(n35528), .A2(n9677), .ZN(n32916) );
  NOR2_X1 U3521 ( .A1(n9677), .A2(n19788), .ZN(n13774) );
  INV_X1 U3531 ( .I(n30054), .ZN(n31296) );
  NAND3_X1 U3534 ( .A1(n30054), .A2(n30053), .A3(n16468), .ZN(n20169) );
  NOR3_X1 U3551 ( .A1(n28222), .A2(n18841), .A3(n16065), .ZN(n35368) );
  OAI22_X1 U3556 ( .A1(n10803), .A2(n29222), .B1(n31772), .B2(n6002), .ZN(
        n12691) );
  NOR2_X1 U3572 ( .A1(n22245), .A2(n7046), .ZN(n22034) );
  NAND2_X1 U3573 ( .A1(n22245), .A2(n20889), .ZN(n22035) );
  NAND3_X1 U3588 ( .A1(n26234), .A2(n26066), .A3(n26067), .ZN(n8248) );
  NOR2_X1 U3594 ( .A1(n9020), .A2(n24309), .ZN(n13547) );
  OR2_X1 U3597 ( .A1(n29532), .A2(n29531), .Z(n17104) );
  NAND3_X1 U3615 ( .A1(n2348), .A2(n1285), .A3(n14379), .ZN(n12202) );
  AND2_X1 U3624 ( .A1(n33086), .A2(n14139), .Z(n34090) );
  AOI22_X1 U3627 ( .A1(n35526), .A2(n33086), .B1(n22263), .B2(n22262), .ZN(
        n14252) );
  AOI21_X1 U3637 ( .A1(n28615), .A2(n13379), .B(n37204), .ZN(n28455) );
  NOR3_X1 U3639 ( .A1(n28453), .A2(n13379), .A3(n180), .ZN(n2573) );
  NOR2_X1 U3644 ( .A1(n12626), .A2(n34777), .ZN(n18124) );
  NAND2_X1 U3673 ( .A1(n31263), .A2(n37502), .ZN(n9961) );
  NAND2_X1 U3677 ( .A1(n28578), .A2(n28591), .ZN(n34670) );
  NAND3_X1 U3683 ( .A1(n585), .A2(n1605), .A3(n33450), .ZN(n1875) );
  NOR2_X1 U3692 ( .A1(n36385), .A2(n24866), .ZN(n8315) );
  NAND2_X1 U3703 ( .A1(n26695), .A2(n10524), .ZN(n26699) );
  NAND2_X1 U3730 ( .A1(n13642), .A2(n21094), .ZN(n10123) );
  AOI22_X1 U3731 ( .A1(n13642), .A2(n11582), .B1(n38986), .B2(n2658), .ZN(
        n14066) );
  INV_X1 U3734 ( .I(n13642), .ZN(n34185) );
  INV_X1 U3736 ( .I(n19680), .ZN(n22129) );
  INV_X1 U3738 ( .I(n21291), .ZN(n21094) );
  NOR2_X1 U3739 ( .A1(n22161), .A2(n6576), .ZN(n36188) );
  NAND2_X1 U3740 ( .A1(n17066), .A2(n24382), .ZN(n16375) );
  NOR2_X1 U3760 ( .A1(n32537), .A2(n13124), .ZN(n33969) );
  INV_X2 U3771 ( .I(n17918), .ZN(n19945) );
  AND2_X1 U3772 ( .A1(n35955), .A2(n30326), .Z(n33973) );
  INV_X1 U3778 ( .I(n38173), .ZN(n1641) );
  INV_X2 U3789 ( .I(n8069), .ZN(n32450) );
  AND2_X1 U3795 ( .A1(n25484), .A2(n36162), .Z(n33976) );
  BUF_X4 U3809 ( .I(n38416), .Z(n3356) );
  INV_X4 U3810 ( .I(n3343), .ZN(n34265) );
  AND3_X1 U3814 ( .A1(n25931), .A2(n37378), .A3(n26135), .Z(n33978) );
  NAND2_X2 U3818 ( .A1(n6075), .A2(n6077), .ZN(n35228) );
  OR2_X1 U3825 ( .A1(n5675), .A2(n32191), .Z(n33979) );
  INV_X2 U3827 ( .I(n28179), .ZN(n36573) );
  AOI21_X2 U3848 ( .A1(n30786), .A2(n28311), .B(n30785), .ZN(n35249) );
  NAND2_X1 U3854 ( .A1(n28355), .A2(n28611), .ZN(n28358) );
  AND3_X1 U3864 ( .A1(n19886), .A2(n12159), .A3(n36296), .Z(n30410) );
  INV_X1 U3865 ( .I(n28186), .ZN(n15597) );
  AOI21_X1 U3867 ( .A1(n37209), .A2(n38724), .B(n11168), .ZN(n11167) );
  NAND2_X1 U3870 ( .A1(n38244), .A2(n38724), .ZN(n22822) );
  CLKBUF_X12 U3876 ( .I(n31558), .Z(n33817) );
  NAND2_X1 U3886 ( .A1(n3059), .A2(n31287), .ZN(n31744) );
  AOI21_X1 U3889 ( .A1(n35004), .A2(n7883), .B(n24314), .ZN(n7036) );
  OAI21_X1 U3891 ( .A1(n11512), .A2(n17447), .B(n28128), .ZN(n14118) );
  OR2_X2 U3901 ( .A1(n8824), .A2(n35233), .Z(n8825) );
  AOI21_X1 U3903 ( .A1(n1205), .A2(n5352), .B(n984), .ZN(n13251) );
  NAND2_X1 U3912 ( .A1(n37378), .A2(n18142), .ZN(n11888) );
  AOI22_X1 U3925 ( .A1(n4195), .A2(n17217), .B1(n36480), .B2(n4194), .ZN(n4193) );
  NAND2_X1 U3926 ( .A1(n15411), .A2(n17217), .ZN(n9060) );
  NOR2_X1 U3932 ( .A1(n23484), .A2(n6303), .ZN(n16716) );
  AOI21_X1 U3951 ( .A1(n924), .A2(n19449), .B(n1006), .ZN(n9099) );
  NAND2_X1 U3965 ( .A1(n27180), .A2(n6686), .ZN(n7231) );
  INV_X1 U3968 ( .I(n6686), .ZN(n36569) );
  NAND2_X1 U3994 ( .A1(n9956), .A2(n4353), .ZN(n2306) );
  INV_X1 U4000 ( .I(n25395), .ZN(n25429) );
  INV_X1 U4003 ( .I(n24753), .ZN(n24126) );
  NOR2_X2 U4006 ( .A1(n24404), .A2(n13904), .ZN(n13412) );
  INV_X2 U4009 ( .I(n16619), .ZN(n28653) );
  NAND2_X1 U4019 ( .A1(n2292), .A2(n26961), .ZN(n26962) );
  INV_X2 U4020 ( .I(n26961), .ZN(n4211) );
  INV_X1 U4038 ( .I(n24933), .ZN(n9324) );
  NAND2_X1 U4051 ( .A1(n26131), .A2(n9916), .ZN(n20771) );
  CLKBUF_X1 U4092 ( .I(n24761), .Z(n34458) );
  INV_X1 U4109 ( .I(n22517), .ZN(n36265) );
  INV_X1 U4113 ( .I(n22620), .ZN(n22724) );
  AND2_X2 U4117 ( .A1(n26668), .A2(n19867), .Z(n14922) );
  BUF_X4 U4145 ( .I(n22767), .Z(n33990) );
  INV_X2 U4148 ( .I(n21150), .ZN(n19637) );
  NOR3_X1 U4163 ( .A1(n9379), .A2(n33440), .A3(n5753), .ZN(n7111) );
  AOI22_X1 U4169 ( .A1(n21991), .A2(n22264), .B1(n22262), .B2(n22261), .ZN(
        n21992) );
  CLKBUF_X12 U4180 ( .I(n15261), .Z(n35248) );
  AOI21_X1 U4182 ( .A1(n38487), .A2(n24381), .B(n7210), .ZN(n24386) );
  NAND3_X2 U4184 ( .A1(n11328), .A2(n35567), .A3(n19586), .ZN(n7683) );
  NOR2_X1 U4187 ( .A1(n26041), .A2(n8407), .ZN(n25869) );
  NOR2_X1 U4191 ( .A1(n22154), .A2(n9824), .ZN(n35194) );
  NAND3_X1 U4192 ( .A1(n12814), .A2(n9824), .A3(n12793), .ZN(n6200) );
  NAND2_X1 U4202 ( .A1(n9824), .A2(n3863), .ZN(n22271) );
  AND3_X2 U4214 ( .A1(n1574), .A2(n24806), .A3(n7552), .Z(n18541) );
  INV_X2 U4216 ( .I(n7552), .ZN(n957) );
  OAI21_X1 U4231 ( .A1(n1643), .A2(n17017), .B(n23569), .ZN(n23217) );
  AND2_X2 U4242 ( .A1(n23132), .A2(n22674), .Z(n36783) );
  OAI22_X1 U4262 ( .A1(n6451), .A2(n33860), .B1(n22177), .B2(n17118), .ZN(
        n36466) );
  AND2_X2 U4269 ( .A1(n35859), .A2(n13745), .Z(n23085) );
  CLKBUF_X1 U4272 ( .I(n9876), .Z(n35685) );
  NAND2_X1 U4273 ( .A1(n22341), .A2(n9876), .ZN(n36176) );
  NOR2_X1 U4274 ( .A1(n22228), .A2(n22229), .ZN(n34256) );
  AND2_X2 U4300 ( .A1(n13572), .A2(n37218), .Z(n7575) );
  NAND2_X1 U4301 ( .A1(n35855), .A2(n7901), .ZN(n25933) );
  INV_X1 U4308 ( .I(n10792), .ZN(n6461) );
  NAND2_X1 U4313 ( .A1(n11081), .A2(n24817), .ZN(n24527) );
  NOR2_X1 U4335 ( .A1(n38996), .A2(n17032), .ZN(n34441) );
  NAND2_X1 U4382 ( .A1(n13872), .A2(n25631), .ZN(n5100) );
  INV_X1 U4402 ( .I(n23963), .ZN(n1622) );
  NOR2_X1 U4418 ( .A1(n11834), .A2(n9413), .ZN(n11833) );
  CLKBUF_X12 U4423 ( .I(n33645), .Z(n32003) );
  CLKBUF_X12 U4429 ( .I(n19658), .Z(n19415) );
  BUF_X4 U4431 ( .I(n3900), .Z(n33995) );
  OR2_X2 U4434 ( .A1(n5871), .A2(n31679), .Z(n18509) );
  NAND3_X1 U4440 ( .A1(n4192), .A2(n32926), .A3(n32566), .ZN(n4014) );
  NAND2_X1 U4451 ( .A1(n4232), .A2(n36827), .ZN(n10543) );
  NAND2_X2 U4452 ( .A1(n22326), .A2(n9165), .ZN(n22328) );
  INV_X1 U4484 ( .I(n5929), .ZN(n8204) );
  NOR2_X1 U4491 ( .A1(n20494), .A2(n39423), .ZN(n20495) );
  NAND2_X1 U4524 ( .A1(n18044), .A2(n28089), .ZN(n32182) );
  NAND2_X1 U4529 ( .A1(n33656), .A2(n28089), .ZN(n8326) );
  OR2_X2 U4535 ( .A1(n10379), .A2(n10375), .Z(n11913) );
  INV_X1 U4538 ( .I(n24070), .ZN(n19646) );
  NAND2_X1 U4549 ( .A1(n27098), .A2(n8412), .ZN(n13896) );
  NOR3_X1 U4569 ( .A1(n378), .A2(n1106), .A3(n36226), .ZN(n195) );
  OAI22_X1 U4591 ( .A1(n37213), .A2(n17624), .B1(n25866), .B2(n35207), .ZN(
        n30656) );
  INV_X1 U4606 ( .I(n9757), .ZN(n1462) );
  INV_X1 U4615 ( .I(n15540), .ZN(n32286) );
  NOR2_X1 U4616 ( .A1(n31418), .A2(n15540), .ZN(n36835) );
  INV_X1 U4625 ( .I(n16445), .ZN(n4986) );
  NOR2_X1 U4641 ( .A1(n25933), .A2(n38168), .ZN(n17954) );
  OR2_X2 U4643 ( .A1(n3092), .A2(n17095), .Z(n20419) );
  NAND3_X1 U4650 ( .A1(n33871), .A2(n25999), .A3(n9833), .ZN(n17994) );
  NAND2_X1 U4673 ( .A1(n26), .A2(n22317), .ZN(n18372) );
  INV_X1 U4675 ( .I(n22317), .ZN(n1679) );
  INV_X1 U4676 ( .I(n384), .ZN(n5405) );
  NOR2_X1 U4682 ( .A1(n15573), .A2(n33046), .ZN(n35789) );
  AOI21_X1 U4690 ( .A1(n19351), .A2(n1645), .B(n23124), .ZN(n23022) );
  NOR2_X1 U4714 ( .A1(n25769), .A2(n25943), .ZN(n6579) );
  INV_X1 U4744 ( .I(n35138), .ZN(n35098) );
  INV_X1 U4759 ( .I(n26092), .ZN(n25945) );
  NAND3_X1 U4794 ( .A1(n29266), .A2(n20026), .A3(n29384), .ZN(n30863) );
  AOI22_X1 U4795 ( .A1(n20099), .A2(n13559), .B1(n30087), .B2(n30093), .ZN(
        n36699) );
  NAND2_X1 U4796 ( .A1(n11940), .A2(n31534), .ZN(n34621) );
  CLKBUF_X2 U4823 ( .I(n29768), .Z(n10096) );
  INV_X1 U4829 ( .I(n28380), .ZN(n34638) );
  INV_X1 U4830 ( .I(n28679), .ZN(n34286) );
  CLKBUF_X2 U4842 ( .I(n16778), .Z(n34459) );
  INV_X2 U4851 ( .I(n28656), .ZN(n28617) );
  NOR2_X1 U4853 ( .A1(n36029), .A2(n10393), .ZN(n36478) );
  AOI21_X1 U4861 ( .A1(n14361), .A2(n9089), .B(n156), .ZN(n34212) );
  CLKBUF_X1 U4867 ( .I(n32474), .Z(n34410) );
  INV_X1 U4896 ( .I(n35617), .ZN(n34770) );
  CLKBUF_X1 U4907 ( .I(n27424), .Z(n35897) );
  CLKBUF_X2 U4914 ( .I(n12485), .Z(n36159) );
  CLKBUF_X2 U4951 ( .I(n9899), .Z(n36078) );
  AND2_X1 U4962 ( .A1(n30883), .A2(n25978), .Z(n25979) );
  NAND2_X1 U4967 ( .A1(n34745), .A2(n5126), .ZN(n34743) );
  CLKBUF_X2 U4993 ( .I(n34692), .Z(n34485) );
  BUF_X2 U4997 ( .I(n5859), .Z(n33348) );
  NAND2_X1 U5010 ( .A1(n15791), .A2(n34076), .ZN(n13743) );
  NAND2_X1 U5014 ( .A1(n12866), .A2(n34027), .ZN(n20337) );
  OR2_X1 U5035 ( .A1(n25637), .A2(n25716), .Z(n34027) );
  CLKBUF_X2 U5057 ( .I(n25581), .Z(n36794) );
  INV_X1 U5058 ( .I(n25290), .ZN(n35894) );
  OAI21_X1 U5061 ( .A1(n24793), .A2(n35981), .B(n35519), .ZN(n24647) );
  INV_X1 U5064 ( .I(n24869), .ZN(n36821) );
  NAND2_X1 U5071 ( .A1(n35521), .A2(n35520), .ZN(n35519) );
  INV_X1 U5073 ( .I(n35952), .ZN(n34694) );
  INV_X2 U5075 ( .I(n24745), .ZN(n16999) );
  BUF_X4 U5116 ( .I(n13045), .Z(n34526) );
  OR2_X1 U5173 ( .A1(n38886), .A2(n1129), .Z(n34077) );
  CLKBUF_X4 U5214 ( .I(n12822), .Z(n36701) );
  INV_X1 U5263 ( .I(n22836), .ZN(n34726) );
  INV_X1 U5265 ( .I(n12245), .ZN(n34772) );
  NOR2_X1 U5272 ( .A1(n8197), .A2(n31183), .ZN(n34727) );
  CLKBUF_X1 U5275 ( .I(n10375), .Z(n34190) );
  BUF_X4 U5297 ( .I(n22085), .Z(n36006) );
  AOI21_X1 U5299 ( .A1(n21947), .A2(n32123), .B(n21946), .ZN(n21953) );
  INV_X1 U5303 ( .I(n19780), .ZN(n34017) );
  BUF_X2 U5306 ( .I(Key[145]), .Z(n19738) );
  OAI21_X1 U5308 ( .A1(n30089), .A2(n1380), .B(n36699), .ZN(n30091) );
  NAND3_X1 U5328 ( .A1(n29559), .A2(n6252), .A3(n35176), .ZN(n35141) );
  NAND2_X1 U5333 ( .A1(n32865), .A2(n30260), .ZN(n36674) );
  INV_X1 U5338 ( .I(n3378), .ZN(n36676) );
  NOR2_X1 U5344 ( .A1(n36268), .A2(n34082), .ZN(n36172) );
  AND2_X1 U5351 ( .A1(n29531), .A2(n29535), .Z(n9636) );
  NAND2_X1 U5361 ( .A1(n20433), .A2(n21023), .ZN(n36126) );
  NAND2_X1 U5366 ( .A1(n29079), .A2(n18457), .ZN(n36997) );
  NAND2_X1 U5367 ( .A1(n29214), .A2(n10628), .ZN(n36694) );
  BUF_X2 U5377 ( .I(n16388), .Z(n5977) );
  OR2_X1 U5380 ( .A1(n16599), .A2(n16388), .Z(n29698) );
  INV_X1 U5394 ( .I(n29500), .ZN(n14873) );
  CLKBUF_X2 U5397 ( .I(n29943), .Z(n36166) );
  INV_X1 U5431 ( .I(n36742), .ZN(n30292) );
  INV_X1 U5445 ( .I(n28604), .ZN(n36248) );
  AND2_X1 U5448 ( .A1(n19893), .A2(n28484), .Z(n34047) );
  NAND2_X1 U5452 ( .A1(n2469), .A2(n19759), .ZN(n35805) );
  INV_X1 U5463 ( .I(n10680), .ZN(n34462) );
  CLKBUF_X1 U5470 ( .I(n13690), .Z(n36165) );
  NAND2_X1 U5493 ( .A1(n30293), .A2(n12531), .ZN(n36525) );
  NOR2_X1 U5495 ( .A1(n28164), .A2(n7690), .ZN(n34596) );
  INV_X1 U5506 ( .I(n34212), .ZN(n4978) );
  INV_X1 U5511 ( .I(n4155), .ZN(n28126) );
  NOR2_X1 U5517 ( .A1(n35469), .A2(n9242), .ZN(n27622) );
  BUF_X2 U5527 ( .I(n7828), .Z(n5469) );
  CLKBUF_X2 U5528 ( .I(n13332), .Z(n36877) );
  BUF_X4 U5530 ( .I(n8057), .Z(n34008) );
  INV_X1 U5532 ( .I(n32581), .ZN(n34313) );
  INV_X4 U5535 ( .I(n6847), .ZN(n900) );
  INV_X1 U5536 ( .I(n11487), .ZN(n11486) );
  NAND2_X1 U5542 ( .A1(n35107), .A2(n36679), .ZN(n27356) );
  NAND2_X1 U5545 ( .A1(n2563), .A2(n35730), .ZN(n35729) );
  INV_X1 U5559 ( .I(n30542), .ZN(n34889) );
  NAND2_X1 U5563 ( .A1(n27353), .A2(n7291), .ZN(n35107) );
  AND2_X1 U5571 ( .A1(n1481), .A2(n7716), .Z(n34114) );
  NAND2_X1 U5572 ( .A1(n19300), .A2(n36073), .ZN(n27057) );
  NOR2_X1 U5574 ( .A1(n35258), .A2(n13266), .ZN(n13268) );
  BUF_X4 U5579 ( .I(n5218), .Z(n34562) );
  NAND2_X1 U5589 ( .A1(n11765), .A2(n27449), .ZN(n34704) );
  CLKBUF_X1 U5595 ( .I(n13278), .Z(n35473) );
  NOR2_X1 U5613 ( .A1(n15616), .A2(n36984), .ZN(n26140) );
  BUF_X2 U5623 ( .I(n2722), .Z(n34853) );
  OAI21_X1 U5633 ( .A1(n26895), .A2(n16222), .B(n16221), .ZN(n16220) );
  NAND2_X1 U5635 ( .A1(n34003), .A2(n35410), .ZN(n35409) );
  AND2_X1 U5638 ( .A1(n8556), .A2(n20936), .Z(n34034) );
  OAI21_X2 U5646 ( .A1(n14485), .A2(n17394), .B(n26933), .ZN(n17393) );
  AND2_X1 U5650 ( .A1(n26707), .A2(n19951), .Z(n32348) );
  CLKBUF_X1 U5663 ( .I(n740), .Z(n35259) );
  INV_X1 U5676 ( .I(n26490), .ZN(n35637) );
  INV_X1 U5679 ( .I(n26233), .ZN(n35471) );
  INV_X1 U5685 ( .I(n26166), .ZN(n35639) );
  CLKBUF_X2 U5694 ( .I(n6130), .Z(n36544) );
  NOR2_X1 U5717 ( .A1(n4553), .A2(n34265), .ZN(n14564) );
  AOI21_X1 U5723 ( .A1(n26071), .A2(n11858), .B(n36896), .ZN(n36900) );
  NAND2_X1 U5730 ( .A1(n25970), .A2(n39015), .ZN(n34645) );
  NAND2_X1 U5735 ( .A1(n26058), .A2(n33293), .ZN(n36658) );
  CLKBUF_X4 U5756 ( .I(n8375), .Z(n36404) );
  BUF_X2 U5762 ( .I(n14212), .Z(n30937) );
  NAND2_X1 U5774 ( .A1(n36324), .A2(n35632), .ZN(n36163) );
  OAI21_X1 U5775 ( .A1(n611), .A2(n32904), .B(n36142), .ZN(n7488) );
  INV_X1 U5803 ( .I(n25068), .ZN(n36324) );
  AND2_X1 U5805 ( .A1(n6300), .A2(n9526), .Z(n34083) );
  BUF_X2 U5836 ( .I(n25481), .Z(n36083) );
  CLKBUF_X4 U5848 ( .I(n21031), .Z(n20052) );
  CLKBUF_X2 U5856 ( .I(n36075), .Z(n35996) );
  CLKBUF_X2 U5859 ( .I(n35900), .Z(n35053) );
  CLKBUF_X2 U5865 ( .I(n25040), .Z(n35379) );
  NOR2_X1 U5882 ( .A1(n24539), .A2(n16990), .ZN(n35118) );
  AOI21_X1 U5890 ( .A1(n24786), .A2(n7831), .B(n36697), .ZN(n30413) );
  NAND2_X1 U5902 ( .A1(n14275), .A2(n1565), .ZN(n35784) );
  OAI21_X1 U5919 ( .A1(n34694), .A2(n3697), .B(n2231), .ZN(n35886) );
  NAND2_X1 U5920 ( .A1(n24613), .A2(n37411), .ZN(n36697) );
  NAND2_X1 U5921 ( .A1(n24659), .A2(n19), .ZN(n36560) );
  INV_X1 U5929 ( .I(n21018), .ZN(n1799) );
  CLKBUF_X2 U5948 ( .I(n24732), .Z(n34662) );
  OAI21_X1 U5958 ( .A1(n17546), .A2(n24467), .B(n35774), .ZN(n24323) );
  BUF_X2 U5968 ( .I(n14999), .Z(n31684) );
  NAND2_X1 U5975 ( .A1(n24818), .A2(n24821), .ZN(n8647) );
  INV_X1 U5980 ( .I(n24821), .ZN(n36180) );
  NAND2_X1 U5993 ( .A1(n35503), .A2(n34043), .ZN(n35056) );
  INV_X2 U5998 ( .I(n8646), .ZN(n24824) );
  CLKBUF_X4 U6003 ( .I(n15467), .Z(n34011) );
  OR2_X1 U6004 ( .A1(n10065), .A2(n10439), .Z(n36542) );
  INV_X1 U6006 ( .I(n35504), .ZN(n35503) );
  NAND2_X2 U6017 ( .A1(n33743), .A2(n36740), .ZN(n30572) );
  CLKBUF_X2 U6035 ( .I(n24247), .Z(n19818) );
  OR2_X1 U6047 ( .A1(n24245), .A2(n24244), .Z(n21080) );
  CLKBUF_X2 U6059 ( .I(n16832), .Z(n36378) );
  CLKBUF_X1 U6065 ( .I(n24279), .Z(n35890) );
  CLKBUF_X2 U6078 ( .I(n24307), .Z(n305) );
  INV_X1 U6088 ( .I(n23960), .ZN(n36541) );
  NOR2_X1 U6094 ( .A1(n35812), .A2(n35811), .ZN(n11452) );
  INV_X1 U6107 ( .I(n9349), .ZN(n35278) );
  INV_X1 U6108 ( .I(n23752), .ZN(n35812) );
  NAND2_X1 U6111 ( .A1(n2274), .A2(n3363), .ZN(n23408) );
  NAND2_X1 U6113 ( .A1(n35007), .A2(n23229), .ZN(n21014) );
  INV_X1 U6115 ( .I(n10633), .ZN(n35892) );
  INV_X1 U6120 ( .I(n36888), .ZN(n23593) );
  NOR2_X1 U6122 ( .A1(n35068), .A2(n35501), .ZN(n13767) );
  CLKBUF_X4 U6153 ( .I(n32366), .Z(n36720) );
  CLKBUF_X2 U6180 ( .I(n11342), .Z(n35068) );
  NOR2_X1 U6183 ( .A1(n14429), .A2(n16197), .ZN(n32583) );
  INV_X1 U6186 ( .I(n34448), .ZN(n14606) );
  NAND2_X1 U6193 ( .A1(n16198), .A2(n23212), .ZN(n34448) );
  INV_X2 U6196 ( .I(n23423), .ZN(n34012) );
  NAND2_X1 U6202 ( .A1(n35806), .A2(n23211), .ZN(n20744) );
  CLKBUF_X2 U6217 ( .I(n33934), .Z(n35567) );
  INV_X1 U6243 ( .I(n18941), .ZN(n35148) );
  INV_X1 U6248 ( .I(n22616), .ZN(n34698) );
  INV_X1 U6269 ( .I(n22744), .ZN(n33863) );
  NAND2_X1 U6279 ( .A1(n34023), .A2(n34256), .ZN(n12568) );
  NOR2_X1 U6280 ( .A1(n22069), .A2(n4114), .ZN(n36084) );
  BUF_X2 U6290 ( .I(n22150), .Z(n31412) );
  CLKBUF_X2 U6295 ( .I(n16880), .Z(n34920) );
  CLKBUF_X4 U6317 ( .I(n36214), .Z(n35771) );
  CLKBUF_X1 U6329 ( .I(n16265), .Z(n35060) );
  NOR2_X1 U6330 ( .A1(n5733), .A2(n17242), .ZN(n3865) );
  INV_X1 U6337 ( .I(n28934), .ZN(n35140) );
  CLKBUF_X2 U6338 ( .I(n21428), .Z(n35973) );
  BUF_X4 U6340 ( .I(n21518), .Z(n34016) );
  NOR2_X1 U6347 ( .A1(n18293), .A2(n19372), .ZN(n37032) );
  INV_X1 U6355 ( .I(n32525), .ZN(n35651) );
  OAI21_X1 U6378 ( .A1(n17948), .A2(n21710), .B(n21868), .ZN(n21) );
  INV_X2 U6383 ( .I(n33249), .ZN(n2690) );
  NOR2_X1 U6389 ( .A1(n3484), .A2(n32410), .ZN(n34932) );
  AOI21_X1 U6406 ( .A1(n36781), .A2(n21484), .B(n36780), .ZN(n36779) );
  NAND2_X1 U6414 ( .A1(n10893), .A2(n36490), .ZN(n4242) );
  CLKBUF_X2 U6415 ( .I(n21791), .Z(n9759) );
  NAND2_X1 U6417 ( .A1(n17763), .A2(n21707), .ZN(n15817) );
  CLKBUF_X2 U6422 ( .I(n21484), .Z(n33852) );
  CLKBUF_X4 U6428 ( .I(n21741), .Z(n1157) );
  OAI22_X1 U6443 ( .A1(n21778), .A2(n34922), .B1(n21612), .B2(n36519), .ZN(
        n21614) );
  INV_X1 U6473 ( .I(n36397), .ZN(n10762) );
  OAI21_X1 U6474 ( .A1(n16536), .A2(n32164), .B(n15125), .ZN(n21658) );
  INV_X1 U6480 ( .I(n14139), .ZN(n22259) );
  INV_X1 U6484 ( .I(n22341), .ZN(n18558) );
  AOI21_X1 U6487 ( .A1(n21702), .A2(n19709), .B(n1353), .ZN(n21703) );
  AOI21_X1 U6490 ( .A1(n7357), .A2(n20646), .B(n20643), .ZN(n35943) );
  CLKBUF_X4 U6494 ( .I(n8899), .Z(n4388) );
  CLKBUF_X1 U6502 ( .I(n22250), .Z(n34488) );
  INV_X1 U6513 ( .I(n22214), .ZN(n22216) );
  INV_X2 U6528 ( .I(n1333), .ZN(n17359) );
  NOR2_X1 U6529 ( .A1(n22160), .A2(n18656), .ZN(n14622) );
  CLKBUF_X2 U6537 ( .I(n19373), .Z(n36303) );
  NAND3_X1 U6544 ( .A1(n21845), .A2(n21844), .A3(n21672), .ZN(n21673) );
  NAND2_X1 U6557 ( .A1(n30828), .A2(n30826), .ZN(n35675) );
  CLKBUF_X2 U6560 ( .I(n19515), .Z(n34452) );
  NOR2_X1 U6581 ( .A1(n22399), .A2(n31857), .ZN(n8662) );
  INV_X1 U6613 ( .I(n22702), .ZN(n22701) );
  INV_X1 U6614 ( .I(n22607), .ZN(n35078) );
  NAND2_X1 U6628 ( .A1(n3273), .A2(n23032), .ZN(n23033) );
  INV_X1 U6638 ( .I(n20449), .ZN(n22866) );
  NAND2_X1 U6639 ( .A1(n11582), .A2(n20570), .ZN(n4890) );
  NAND2_X1 U6640 ( .A1(n9954), .A2(n14390), .ZN(n23004) );
  NAND2_X1 U6662 ( .A1(n30594), .A2(n20372), .ZN(n3811) );
  NAND2_X1 U6663 ( .A1(n23013), .A2(n23012), .ZN(n5039) );
  INV_X1 U6665 ( .I(n14560), .ZN(n23000) );
  NOR2_X1 U6666 ( .A1(n12925), .A2(n36369), .ZN(n36368) );
  NAND2_X1 U6671 ( .A1(n13734), .A2(n19788), .ZN(n22839) );
  INV_X1 U6673 ( .I(n5337), .ZN(n15045) );
  AOI22_X1 U6699 ( .A1(n15885), .A2(n23128), .B1(n19621), .B2(n34014), .ZN(
        n15884) );
  NAND2_X1 U6700 ( .A1(n12621), .A2(n36763), .ZN(n12620) );
  NAND3_X1 U6702 ( .A1(n15163), .A2(n22810), .A3(n22809), .ZN(n16731) );
  NAND2_X1 U6708 ( .A1(n11108), .A2(n23423), .ZN(n1893) );
  NAND2_X1 U6716 ( .A1(n23358), .A2(n30299), .ZN(n36035) );
  NAND2_X1 U6724 ( .A1(n35130), .A2(n23315), .ZN(n33638) );
  NAND2_X1 U6742 ( .A1(n23749), .A2(n9321), .ZN(n35007) );
  OAI21_X1 U6768 ( .A1(n16094), .A2(n15176), .B(n35569), .ZN(n36785) );
  INV_X1 U6773 ( .I(n18849), .ZN(n13224) );
  INV_X1 U6781 ( .I(n7475), .ZN(n7185) );
  INV_X1 U6785 ( .I(n13395), .ZN(n23789) );
  NOR2_X1 U6799 ( .A1(n35253), .A2(n18907), .ZN(n31488) );
  INV_X1 U6801 ( .I(n23073), .ZN(n34900) );
  INV_X1 U6817 ( .I(n24457), .ZN(n2972) );
  NAND3_X1 U6831 ( .A1(n17711), .A2(n36757), .A3(n17709), .ZN(n17710) );
  NOR3_X1 U6839 ( .A1(n11361), .A2(n19895), .A3(n24359), .ZN(n23941) );
  AOI21_X1 U6846 ( .A1(n24087), .A2(n24433), .B(n1608), .ZN(n10023) );
  NAND3_X1 U6851 ( .A1(n1282), .A2(n20404), .A3(n24346), .ZN(n24347) );
  INV_X1 U6852 ( .I(n5955), .ZN(n24348) );
  NOR2_X1 U6856 ( .A1(n14704), .A2(n1283), .ZN(n13186) );
  NAND2_X1 U6861 ( .A1(n17259), .A2(n7240), .ZN(n3307) );
  OAI21_X1 U6874 ( .A1(n12423), .A2(n18920), .B(n1594), .ZN(n12422) );
  OR2_X1 U6875 ( .A1(n7693), .A2(n17087), .Z(n34115) );
  CLKBUF_X2 U6884 ( .I(n24492), .Z(n36090) );
  NAND2_X1 U6894 ( .A1(n18324), .A2(n24764), .ZN(n18325) );
  OR2_X1 U6901 ( .A1(n36471), .A2(n2018), .Z(n20064) );
  AOI21_X1 U6905 ( .A1(n11846), .A2(n19828), .B(n5957), .ZN(n7930) );
  NOR3_X1 U6919 ( .A1(n13128), .A2(n2747), .A3(n2731), .ZN(n2730) );
  NOR2_X1 U6922 ( .A1(n34935), .A2(n34934), .ZN(n34821) );
  INV_X1 U6931 ( .I(n38171), .ZN(n24978) );
  NOR3_X1 U6939 ( .A1(n35952), .A2(n3697), .A3(n14999), .ZN(n33945) );
  NAND2_X1 U6953 ( .A1(n11642), .A2(n31530), .ZN(n24882) );
  CLKBUF_X2 U6977 ( .I(n6759), .Z(n61) );
  INV_X1 U6980 ( .I(n25225), .ZN(n35511) );
  NOR2_X1 U6989 ( .A1(n4048), .A2(n18734), .ZN(n15356) );
  NOR2_X1 U6995 ( .A1(n36708), .A2(n36707), .ZN(n30705) );
  NAND2_X1 U6998 ( .A1(n33491), .A2(n20515), .ZN(n36323) );
  NAND2_X1 U7003 ( .A1(n36794), .A2(n25390), .ZN(n24894) );
  NAND2_X1 U7005 ( .A1(n1253), .A2(n16677), .ZN(n25388) );
  NOR2_X1 U7006 ( .A1(n15356), .A2(n19637), .ZN(n15355) );
  NAND2_X1 U7018 ( .A1(n1253), .A2(n19941), .ZN(n36793) );
  OR2_X1 U7020 ( .A1(n25261), .A2(n32989), .Z(n34103) );
  NOR2_X1 U7029 ( .A1(n25545), .A2(n25481), .ZN(n2247) );
  OR2_X1 U7032 ( .A1(n25680), .A2(n30633), .Z(n7540) );
  NAND2_X1 U7037 ( .A1(n25402), .A2(n5314), .ZN(n18113) );
  INV_X1 U7043 ( .I(n19264), .ZN(n12381) );
  NAND2_X1 U7046 ( .A1(n25547), .A2(n19701), .ZN(n18599) );
  NAND2_X1 U7048 ( .A1(n25416), .A2(n30377), .ZN(n14914) );
  OAI21_X1 U7049 ( .A1(n37049), .A2(n31457), .B(n32101), .ZN(n36277) );
  INV_X1 U7068 ( .I(n25111), .ZN(n25994) );
  NAND2_X1 U7070 ( .A1(n1101), .A2(n9380), .ZN(n8860) );
  INV_X2 U7089 ( .I(n16250), .ZN(n12199) );
  NAND2_X1 U7095 ( .A1(n34692), .A2(n36532), .ZN(n26129) );
  INV_X1 U7121 ( .I(n26340), .ZN(n26341) );
  NOR2_X1 U7125 ( .A1(n37073), .A2(n11858), .ZN(n17311) );
  INV_X1 U7130 ( .I(n26601), .ZN(n34478) );
  INV_X1 U7132 ( .I(n2594), .ZN(n5381) );
  NAND3_X1 U7142 ( .A1(n13391), .A2(n35744), .A3(n17008), .ZN(n26096) );
  INV_X1 U7158 ( .I(n26492), .ZN(n159) );
  INV_X1 U7163 ( .I(n5078), .ZN(n35967) );
  NAND2_X1 U7178 ( .A1(n30942), .A2(n1006), .ZN(n4651) );
  NAND3_X1 U7189 ( .A1(n1088), .A2(n26701), .A3(n26700), .ZN(n26706) );
  NAND2_X1 U7211 ( .A1(n3449), .A2(n13588), .ZN(n31226) );
  NAND2_X1 U7212 ( .A1(n21277), .A2(n20936), .ZN(n2101) );
  CLKBUF_X4 U7217 ( .I(n26747), .Z(n15594) );
  NAND2_X1 U7225 ( .A1(n34003), .A2(n34426), .ZN(n26785) );
  NAND2_X1 U7227 ( .A1(n6190), .A2(n10440), .ZN(n35489) );
  OAI21_X1 U7236 ( .A1(n14412), .A2(n15411), .B(n32892), .ZN(n36445) );
  NOR2_X1 U7242 ( .A1(n26632), .A2(n12755), .ZN(n19250) );
  NAND2_X1 U7249 ( .A1(n862), .A2(n2451), .ZN(n26892) );
  AOI21_X1 U7260 ( .A1(n925), .A2(n1008), .B(n15825), .ZN(n7007) );
  INV_X1 U7264 ( .I(n26264), .ZN(n34228) );
  NAND2_X1 U7273 ( .A1(n6605), .A2(n5720), .ZN(n7585) );
  NAND3_X1 U7276 ( .A1(n26722), .A2(n16970), .A3(n19225), .ZN(n8685) );
  NAND2_X1 U7299 ( .A1(n27214), .A2(n11765), .ZN(n27093) );
  INV_X1 U7337 ( .I(n27259), .ZN(n5365) );
  AOI21_X1 U7348 ( .A1(n10946), .A2(n27403), .B(n35258), .ZN(n31185) );
  NAND3_X1 U7365 ( .A1(n11805), .A2(n32463), .A3(n38907), .ZN(n576) );
  AOI22_X1 U7368 ( .A1(n27388), .A2(n14327), .B1(n39826), .B2(n2761), .ZN(
        n31943) );
  NAND2_X1 U7369 ( .A1(n34705), .A2(n34704), .ZN(n34493) );
  NAND2_X1 U7385 ( .A1(n27335), .A2(n2035), .ZN(n27487) );
  INV_X1 U7404 ( .I(n14808), .ZN(n35889) );
  NAND3_X1 U7418 ( .A1(n1086), .A2(n17166), .A3(n4781), .ZN(n12075) );
  INV_X1 U7420 ( .I(n27707), .ZN(n34708) );
  INV_X1 U7422 ( .I(n27678), .ZN(n34409) );
  INV_X1 U7426 ( .I(n886), .ZN(n36325) );
  INV_X1 U7429 ( .I(n4266), .ZN(n35089) );
  NOR2_X1 U7437 ( .A1(n28194), .A2(n17197), .ZN(n27928) );
  NOR2_X1 U7445 ( .A1(n27970), .A2(n28148), .ZN(n19969) );
  NAND2_X1 U7448 ( .A1(n28114), .A2(n28115), .ZN(n3066) );
  NOR2_X1 U7451 ( .A1(n580), .A2(n39571), .ZN(n7223) );
  NAND2_X1 U7458 ( .A1(n8207), .A2(n1204), .ZN(n8327) );
  NAND2_X1 U7472 ( .A1(n28172), .A2(n28258), .ZN(n18192) );
  OR2_X1 U7477 ( .A1(n28278), .A2(n19995), .Z(n27543) );
  NAND2_X1 U7484 ( .A1(n12260), .A2(n9845), .ZN(n13876) );
  NOR2_X1 U7511 ( .A1(n6819), .A2(n35911), .ZN(n3055) );
  NOR3_X1 U7516 ( .A1(n1195), .A2(n31542), .A3(n8131), .ZN(n32800) );
  NAND2_X1 U7523 ( .A1(n33046), .A2(n1815), .ZN(n28640) );
  NAND2_X1 U7536 ( .A1(n28409), .A2(n1426), .ZN(n28410) );
  INV_X1 U7538 ( .I(n5645), .ZN(n31615) );
  INV_X1 U7540 ( .I(n28997), .ZN(n1412) );
  INV_X1 U7541 ( .I(n28966), .ZN(n15682) );
  INV_X1 U7544 ( .I(n29152), .ZN(n36828) );
  CLKBUF_X2 U7547 ( .I(n28840), .Z(n7667) );
  CLKBUF_X2 U7553 ( .I(n29381), .Z(n32906) );
  CLKBUF_X1 U7570 ( .I(n29769), .Z(n28) );
  NAND2_X1 U7578 ( .A1(n5335), .A2(n1055), .ZN(n4790) );
  NOR2_X1 U7583 ( .A1(n18104), .A2(n29956), .ZN(n29905) );
  OR2_X1 U7584 ( .A1(n20524), .A2(n19224), .Z(n30152) );
  NAND2_X1 U7585 ( .A1(n38051), .A2(n2954), .ZN(n29502) );
  INV_X1 U7589 ( .I(n3430), .ZN(n35975) );
  AOI21_X1 U7593 ( .A1(n36550), .A2(n16828), .B(n29385), .ZN(n31180) );
  NAND2_X1 U7594 ( .A1(n28880), .A2(n31511), .ZN(n34806) );
  NAND3_X1 U7596 ( .A1(n29770), .A2(n29843), .A3(n29844), .ZN(n29771) );
  NAND3_X1 U7602 ( .A1(n30720), .A2(n1757), .A3(n11826), .ZN(n33557) );
  INV_X1 U7605 ( .I(n5530), .ZN(n3378) );
  INV_X1 U7606 ( .I(n15841), .ZN(n29440) );
  OAI22_X1 U7611 ( .A1(n29369), .A2(n11067), .B1(n13981), .B2(n16683), .ZN(
        n13277) );
  CLKBUF_X2 U7619 ( .I(n18257), .Z(n32050) );
  OAI22_X1 U7620 ( .A1(n10942), .A2(n30033), .B1(n30014), .B2(n15643), .ZN(
        n32531) );
  INV_X1 U7623 ( .I(n30203), .ZN(n1050) );
  AOI22_X1 U7624 ( .A1(n30039), .A2(n35103), .B1(n30036), .B2(n30037), .ZN(
        n30040) );
  OR2_X1 U7629 ( .A1(n22282), .A2(n22130), .Z(n34019) );
  XNOR2_X1 U7631 ( .A1(n4441), .A2(n10213), .ZN(n34020) );
  NAND2_X1 U7632 ( .A1(n9737), .A2(n12535), .ZN(n34021) );
  XNOR2_X1 U7634 ( .A1(n15413), .A2(n13356), .ZN(n34022) );
  XNOR2_X1 U7636 ( .A1(n26296), .A2(n26295), .ZN(n34024) );
  AND2_X1 U7644 ( .A1(n34014), .A2(n3273), .Z(n34030) );
  AND2_X1 U7645 ( .A1(n34080), .A2(n959), .Z(n34031) );
  XNOR2_X1 U7647 ( .A1(n25298), .A2(n30101), .ZN(n34032) );
  AND2_X1 U7649 ( .A1(n38163), .A2(n30128), .Z(n34033) );
  OR2_X1 U7654 ( .A1(n33888), .A2(n994), .Z(n34037) );
  XNOR2_X1 U7657 ( .A1(n28931), .A2(n28930), .ZN(n34038) );
  AND2_X1 U7659 ( .A1(n1432), .A2(n8349), .Z(n34041) );
  AND2_X1 U7663 ( .A1(n38317), .A2(n38668), .Z(n34042) );
  OR2_X1 U7667 ( .A1(n38303), .A2(n6849), .Z(n34043) );
  OR2_X1 U7676 ( .A1(n21860), .A2(n19641), .Z(n34048) );
  AND2_X1 U7681 ( .A1(n10120), .A2(n21839), .Z(n34049) );
  XOR2_X1 U7683 ( .A1(n18270), .A2(n32931), .Z(n34050) );
  XNOR2_X1 U7686 ( .A1(n3610), .A2(n19751), .ZN(n34052) );
  XNOR2_X1 U7688 ( .A1(n35376), .A2(n19613), .ZN(n34053) );
  XNOR2_X1 U7689 ( .A1(n13617), .A2(n29371), .ZN(n34054) );
  XNOR2_X1 U7693 ( .A1(n14907), .A2(n1459), .ZN(n34056) );
  AND2_X1 U7694 ( .A1(n32262), .A2(n32261), .Z(n34057) );
  AND2_X1 U7696 ( .A1(n14734), .A2(n14527), .Z(n34059) );
  XNOR2_X1 U7710 ( .A1(n7161), .A2(n7158), .ZN(n34062) );
  AND3_X1 U7715 ( .A1(n26764), .A2(n3606), .A3(n13393), .Z(n34063) );
  AND2_X1 U7721 ( .A1(n19647), .A2(n668), .Z(n34066) );
  OR2_X1 U7723 ( .A1(n13998), .A2(n13997), .Z(n34067) );
  AND2_X1 U7735 ( .A1(n9954), .A2(n19823), .Z(n34072) );
  INV_X1 U7739 ( .I(n8071), .ZN(n1339) );
  BUF_X2 U7740 ( .I(n8071), .Z(n5821) );
  AND2_X1 U7757 ( .A1(n25361), .A2(n12896), .Z(n34085) );
  OR2_X2 U7759 ( .A1(n16080), .A2(n14473), .Z(n34087) );
  XNOR2_X1 U7761 ( .A1(n17048), .A2(n33551), .ZN(n34088) );
  OR2_X1 U7766 ( .A1(n29701), .A2(n28414), .Z(n34089) );
  XNOR2_X1 U7769 ( .A1(n25256), .A2(n4556), .ZN(n34092) );
  XNOR2_X1 U7771 ( .A1(n29463), .A2(n27815), .ZN(n34094) );
  XNOR2_X1 U7776 ( .A1(n25229), .A2(n1710), .ZN(n34096) );
  OR2_X1 U7779 ( .A1(n34180), .A2(n29700), .Z(n34097) );
  XNOR2_X1 U7790 ( .A1(n22486), .A2(n22426), .ZN(n34104) );
  AND2_X1 U7793 ( .A1(n30843), .A2(n8264), .Z(n34105) );
  AND2_X1 U7804 ( .A1(n25677), .A2(n19589), .Z(n34112) );
  INV_X1 U7807 ( .I(n23792), .ZN(n34851) );
  INV_X1 U7809 ( .I(n29474), .ZN(n36040) );
  INV_X1 U7810 ( .I(n28807), .ZN(n28764) );
  INV_X1 U7818 ( .I(n29732), .ZN(n29753) );
  INV_X1 U7824 ( .I(n38217), .ZN(n11181) );
  XNOR2_X1 U7839 ( .A1(Key[189]), .A2(Plaintext[189]), .ZN(n34122) );
  AND2_X1 U7859 ( .A1(n3628), .A2(n16967), .Z(n34124) );
  INV_X2 U7861 ( .I(n4886), .ZN(n27069) );
  XNOR2_X1 U7863 ( .A1(n14374), .A2(n25193), .ZN(n34126) );
  OR2_X2 U7875 ( .A1(n22100), .A2(n22058), .Z(n34128) );
  AND2_X1 U7884 ( .A1(n23478), .A2(n23479), .Z(n34129) );
  INV_X1 U7888 ( .I(n37815), .ZN(n23159) );
  XNOR2_X1 U7892 ( .A1(n7475), .A2(n23880), .ZN(n34132) );
  XNOR2_X1 U7913 ( .A1(n39797), .A2(n29562), .ZN(n34135) );
  XOR2_X1 U7916 ( .A1(n33271), .A2(n25194), .Z(n34136) );
  XNOR2_X1 U7919 ( .A1(n25284), .A2(n25283), .ZN(n34137) );
  XNOR2_X1 U7935 ( .A1(n25006), .A2(n34945), .ZN(n34139) );
  XNOR2_X1 U7944 ( .A1(n25215), .A2(n29857), .ZN(n34142) );
  XNOR2_X1 U7947 ( .A1(n29707), .A2(n7481), .ZN(n34144) );
  XNOR2_X1 U7950 ( .A1(n19729), .A2(n26514), .ZN(n34145) );
  XNOR2_X1 U7951 ( .A1(n24985), .A2(n24984), .ZN(n34147) );
  OR2_X2 U7952 ( .A1(n20491), .A2(n20490), .Z(n34148) );
  XNOR2_X1 U7953 ( .A1(n37498), .A2(n35702), .ZN(n34149) );
  XNOR2_X1 U7961 ( .A1(n8340), .A2(n25853), .ZN(n34151) );
  XNOR2_X1 U7965 ( .A1(n26403), .A2(n15530), .ZN(n34152) );
  AND2_X2 U7967 ( .A1(n31362), .A2(n9833), .Z(n34154) );
  XNOR2_X1 U7971 ( .A1(n37476), .A2(n39559), .ZN(n34157) );
  INV_X1 U7977 ( .I(n18135), .ZN(n26220) );
  XNOR2_X1 U7983 ( .A1(n19450), .A2(n19733), .ZN(n34161) );
  INV_X1 U7984 ( .I(n7959), .ZN(n26702) );
  XOR2_X1 U7988 ( .A1(n27746), .A2(n19733), .Z(n34162) );
  NOR2_X1 U7991 ( .A1(n1093), .A2(n11334), .ZN(n34163) );
  XNOR2_X1 U8031 ( .A1(n21084), .A2(n30956), .ZN(n34175) );
  XNOR2_X1 U8035 ( .A1(n9786), .A2(n28994), .ZN(n34179) );
  XNOR2_X1 U8043 ( .A1(n29153), .A2(n14195), .ZN(n34181) );
  AND2_X1 U8044 ( .A1(n29755), .A2(n29754), .Z(n34182) );
  XNOR2_X1 U8045 ( .A1(n3941), .A2(n632), .ZN(n34183) );
  NAND2_X1 U8050 ( .A1(n34186), .A2(n5469), .ZN(n20306) );
  NAND2_X2 U8076 ( .A1(n36972), .A2(n28065), .ZN(n7429) );
  NAND2_X1 U8080 ( .A1(n6118), .A2(n6119), .ZN(n6117) );
  NOR2_X2 U8086 ( .A1(n34261), .A2(n25602), .ZN(n34260) );
  NAND2_X1 U8087 ( .A1(n36902), .A2(n26), .ZN(n20986) );
  XOR2_X1 U8102 ( .A1(n20025), .A2(n29072), .Z(n4616) );
  OAI21_X2 U8107 ( .A1(n28317), .A2(n28316), .B(n28315), .ZN(n29072) );
  NOR2_X2 U8120 ( .A1(n20319), .A2(n27879), .ZN(n28874) );
  AOI22_X2 U8124 ( .A1(n34193), .A2(n2603), .B1(n15623), .B2(n1076), .ZN(
        n15023) );
  AND2_X1 U8125 ( .A1(n28149), .A2(n2604), .Z(n34193) );
  XOR2_X1 U8130 ( .A1(n25210), .A2(n14214), .Z(n5721) );
  XOR2_X1 U8139 ( .A1(n135), .A2(n34196), .Z(n8365) );
  XOR2_X1 U8140 ( .A1(n6283), .A2(n650), .Z(n34196) );
  AOI21_X2 U8141 ( .A1(n16670), .A2(n16669), .B(n34197), .ZN(n16668) );
  XOR2_X1 U8150 ( .A1(n34178), .A2(n3082), .Z(n6316) );
  BUF_X4 U8158 ( .I(n35399), .Z(n35290) );
  OR2_X1 U8159 ( .A1(n12260), .A2(n12257), .Z(n12259) );
  INV_X2 U8161 ( .I(n16699), .ZN(n36105) );
  AOI21_X2 U8162 ( .A1(n7058), .A2(n12080), .B(n34201), .ZN(n22549) );
  OAI21_X2 U8163 ( .A1(n12080), .A2(n21865), .B(n36680), .ZN(n34201) );
  XOR2_X1 U8166 ( .A1(n3476), .A2(n34202), .Z(n7518) );
  NOR2_X1 U8173 ( .A1(n38487), .A2(n33314), .ZN(n6567) );
  INV_X1 U8182 ( .I(n25302), .ZN(n34208) );
  INV_X2 U8189 ( .I(n34203), .ZN(n30844) );
  XOR2_X1 U8191 ( .A1(n3185), .A2(n3186), .Z(n34203) );
  INV_X1 U8193 ( .I(n9059), .ZN(n34205) );
  AND2_X1 U8206 ( .A1(n15172), .A2(n11150), .Z(n14589) );
  NAND3_X2 U8217 ( .A1(n14748), .A2(n14747), .A3(n15238), .ZN(n4524) );
  NAND2_X1 U8219 ( .A1(n37003), .A2(n34521), .ZN(n10814) );
  AOI22_X2 U8221 ( .A1(n16016), .A2(n17102), .B1(n21029), .B2(n21601), .ZN(
        n16015) );
  NOR2_X2 U8222 ( .A1(n16302), .A2(n33280), .ZN(n16016) );
  XOR2_X1 U8223 ( .A1(n30632), .A2(n23850), .Z(n311) );
  XOR2_X1 U8227 ( .A1(n34208), .A2(n25329), .Z(n34414) );
  XOR2_X1 U8228 ( .A1(n17908), .A2(n19014), .Z(n17907) );
  NAND3_X2 U8241 ( .A1(n31704), .A2(n30863), .A3(n29353), .ZN(n29367) );
  XOR2_X1 U8268 ( .A1(n11563), .A2(n34213), .Z(n7090) );
  AND2_X1 U8270 ( .A1(n22229), .A2(n22228), .Z(n17145) );
  NAND2_X1 U8275 ( .A1(n13166), .A2(n34576), .ZN(n4726) );
  XOR2_X1 U8280 ( .A1(n17455), .A2(n26596), .Z(n34214) );
  XOR2_X1 U8303 ( .A1(Plaintext[66]), .A2(Key[66]), .Z(n261) );
  AOI22_X1 U8305 ( .A1(n29860), .A2(n29859), .B1(n34215), .B2(n36764), .ZN(
        n2070) );
  OR2_X1 U8306 ( .A1(n2073), .A2(n2858), .Z(n34215) );
  OAI22_X2 U8316 ( .A1(n21566), .A2(n7183), .B1(n35), .B2(n36), .ZN(n22038) );
  INV_X2 U8318 ( .I(n34218), .ZN(n889) );
  XOR2_X1 U8336 ( .A1(n34221), .A2(n12205), .Z(n36831) );
  XOR2_X1 U8337 ( .A1(n21866), .A2(n13591), .Z(n34221) );
  NOR2_X1 U8349 ( .A1(n29336), .A2(n14858), .ZN(n4520) );
  XOR2_X1 U8363 ( .A1(n9205), .A2(n22618), .Z(n12016) );
  AND2_X1 U8374 ( .A1(n24244), .A2(n9520), .Z(n9386) );
  NOR2_X2 U8392 ( .A1(n20211), .A2(n13757), .ZN(n34224) );
  NAND2_X1 U8402 ( .A1(n15430), .A2(n34225), .ZN(n35033) );
  NAND2_X1 U8403 ( .A1(n30811), .A2(n34226), .ZN(n34225) );
  NOR2_X1 U8405 ( .A1(n34228), .A2(n34227), .ZN(n34226) );
  NAND2_X1 U8406 ( .A1(n15429), .A2(n29602), .ZN(n34227) );
  MUX2_X1 U8413 ( .I0(n12527), .I1(n36588), .S(n5383), .Z(n2334) );
  NAND3_X2 U8417 ( .A1(n36460), .A2(n34501), .A3(n36459), .ZN(n3213) );
  OR2_X1 U8444 ( .A1(n25829), .A2(n32193), .Z(n1956) );
  OAI21_X2 U8446 ( .A1(n20222), .A2(n35230), .B(n20221), .ZN(n23829) );
  XOR2_X1 U8448 ( .A1(n21284), .A2(n34231), .Z(n8554) );
  XOR2_X1 U8456 ( .A1(n269), .A2(n35464), .Z(n34231) );
  XOR2_X1 U8463 ( .A1(n15871), .A2(n22621), .Z(n22714) );
  NAND2_X2 U8485 ( .A1(n6012), .A2(n35436), .ZN(n34279) );
  NAND2_X2 U8493 ( .A1(n34233), .A2(n12883), .ZN(n16309) );
  OAI21_X2 U8495 ( .A1(n12882), .A2(n32236), .B(n21073), .ZN(n34233) );
  INV_X2 U8505 ( .I(n34235), .ZN(n33964) );
  XOR2_X1 U8507 ( .A1(n12560), .A2(n12563), .Z(n34235) );
  NAND3_X1 U8515 ( .A1(n26217), .A2(n26216), .A3(n26218), .ZN(n34237) );
  NAND2_X1 U8516 ( .A1(n5670), .A2(n5525), .ZN(n34515) );
  AOI21_X1 U8522 ( .A1(n14928), .A2(n8493), .B(n19604), .ZN(n14927) );
  XOR2_X1 U8525 ( .A1(n10117), .A2(n34238), .Z(n32540) );
  XOR2_X1 U8529 ( .A1(n38207), .A2(n34239), .Z(n34238) );
  XOR2_X1 U8556 ( .A1(n22552), .A2(n14309), .Z(n7039) );
  NAND2_X2 U8558 ( .A1(n13766), .A2(n13765), .ZN(n14309) );
  BUF_X2 U8600 ( .I(n6263), .Z(n34245) );
  NAND2_X1 U8601 ( .A1(n30252), .A2(n30250), .ZN(n16167) );
  NAND2_X2 U8604 ( .A1(n19663), .A2(n30259), .ZN(n30252) );
  NOR2_X1 U8607 ( .A1(n21662), .A2(n36728), .ZN(n21946) );
  NAND2_X2 U8617 ( .A1(n35644), .A2(n32552), .ZN(n23548) );
  NAND2_X2 U8633 ( .A1(n18227), .A2(n21229), .ZN(n34962) );
  OR2_X1 U8642 ( .A1(n12078), .A2(n19371), .Z(n9204) );
  OAI21_X2 U8645 ( .A1(n26922), .A2(n19371), .B(n26764), .ZN(n12078) );
  XNOR2_X1 U8648 ( .A1(n11201), .A2(n30065), .ZN(n34274) );
  XOR2_X1 U8664 ( .A1(Plaintext[157]), .A2(Key[157]), .Z(n34247) );
  XOR2_X1 U8682 ( .A1(n12195), .A2(n18778), .Z(n15413) );
  NAND2_X2 U8684 ( .A1(n4630), .A2(n4629), .ZN(n12195) );
  XOR2_X1 U8695 ( .A1(n22747), .A2(n12194), .Z(n34250) );
  NAND3_X2 U8698 ( .A1(n7722), .A2(n18660), .A3(n22168), .ZN(n23472) );
  INV_X4 U8705 ( .I(n25328), .ZN(n36133) );
  XOR2_X1 U8711 ( .A1(n8181), .A2(n34251), .Z(n34594) );
  XOR2_X1 U8729 ( .A1(n12935), .A2(n12934), .Z(n12933) );
  XOR2_X1 U8743 ( .A1(n30831), .A2(n17043), .Z(n36034) );
  XOR2_X1 U8813 ( .A1(n25249), .A2(n25100), .Z(n24544) );
  NAND2_X2 U8817 ( .A1(n33896), .A2(n8606), .ZN(n25249) );
  XOR2_X1 U8824 ( .A1(n23928), .A2(n23965), .Z(n31851) );
  NAND2_X2 U8855 ( .A1(n34984), .A2(n12499), .ZN(n34559) );
  NOR2_X2 U8877 ( .A1(n14091), .A2(n28426), .ZN(n29167) );
  AOI21_X2 U8879 ( .A1(n35525), .A2(n12083), .B(n1292), .ZN(n12027) );
  INV_X2 U8880 ( .I(n14011), .ZN(n1292) );
  NAND2_X2 U8884 ( .A1(n7011), .A2(n15375), .ZN(n14011) );
  AOI21_X2 U8900 ( .A1(n11379), .A2(n34246), .B(n34259), .ZN(n22623) );
  OAI22_X2 U8915 ( .A1(n16580), .A2(n18290), .B1(n29482), .B2(n12479), .ZN(
        n29531) );
  AOI22_X2 U8925 ( .A1(n34868), .A2(n34262), .B1(n12590), .B2(n30335), .ZN(
        n27064) );
  NOR2_X1 U8933 ( .A1(n29841), .A2(n105), .ZN(n21236) );
  NAND2_X2 U8942 ( .A1(n33255), .A2(n13267), .ZN(n20706) );
  XOR2_X1 U8946 ( .A1(n7967), .A2(n24927), .Z(n25156) );
  NAND2_X2 U8949 ( .A1(n4224), .A2(n4227), .ZN(n24927) );
  NAND3_X2 U8957 ( .A1(n10003), .A2(n29851), .A3(n32258), .ZN(n34267) );
  XOR2_X1 U8970 ( .A1(n8702), .A2(n14507), .Z(n20627) );
  NOR2_X2 U8972 ( .A1(n7658), .A2(n9193), .ZN(n34268) );
  INV_X2 U8976 ( .I(n17095), .ZN(n13753) );
  NAND2_X2 U8977 ( .A1(n33631), .A2(n3095), .ZN(n17095) );
  XOR2_X1 U8985 ( .A1(n32433), .A2(n25175), .Z(n25254) );
  AOI21_X2 U8987 ( .A1(n33755), .A2(n33754), .B(n30385), .ZN(n32433) );
  INV_X2 U8988 ( .I(n33539), .ZN(n34857) );
  XOR2_X1 U8996 ( .A1(n26342), .A2(n26494), .Z(n10233) );
  NAND2_X2 U9010 ( .A1(n34270), .A2(n13134), .ZN(n5530) );
  OAI21_X2 U9011 ( .A1(n13136), .A2(n37146), .B(n13762), .ZN(n34270) );
  NAND2_X2 U9012 ( .A1(n34272), .A2(n39821), .ZN(n36535) );
  NAND3_X1 U9017 ( .A1(n17508), .A2(n32601), .A3(n17511), .ZN(n22680) );
  XOR2_X1 U9018 ( .A1(n20753), .A2(n34274), .Z(n10501) );
  NAND2_X2 U9035 ( .A1(n34275), .A2(n15795), .ZN(n2542) );
  OAI21_X2 U9040 ( .A1(n945), .A2(n15984), .B(n34276), .ZN(n15982) );
  NAND2_X2 U9042 ( .A1(n15983), .A2(n945), .ZN(n34276) );
  XOR2_X1 U9057 ( .A1(n14941), .A2(n28991), .Z(n29039) );
  NAND3_X2 U9059 ( .A1(n28471), .A2(n28470), .A3(n28730), .ZN(n28991) );
  XOR2_X1 U9062 ( .A1(n11541), .A2(n22761), .Z(n22543) );
  NAND2_X1 U9065 ( .A1(n25544), .A2(n15515), .ZN(n19702) );
  AOI21_X2 U9067 ( .A1(n28107), .A2(n28108), .B(n28106), .ZN(n34695) );
  AOI21_X2 U9076 ( .A1(n18312), .A2(n23333), .B(n12191), .ZN(n23245) );
  NAND2_X2 U9078 ( .A1(n6969), .A2(n3256), .ZN(n23333) );
  NOR2_X2 U9081 ( .A1(n37171), .A2(n34277), .ZN(n3112) );
  NAND2_X1 U9088 ( .A1(n24577), .A2(n19484), .ZN(n24578) );
  NAND2_X2 U9099 ( .A1(n8262), .A2(n27240), .ZN(n27102) );
  OR2_X1 U9105 ( .A1(n21111), .A2(n18926), .Z(n21558) );
  NAND2_X2 U9124 ( .A1(n17299), .A2(n17301), .ZN(n33230) );
  XOR2_X1 U9135 ( .A1(n10492), .A2(n10491), .Z(n9984) );
  XOR2_X1 U9139 ( .A1(n34284), .A2(n17428), .Z(Ciphertext[188]) );
  AOI22_X1 U9140 ( .A1(n16167), .A2(n11700), .B1(n13990), .B2(n13991), .ZN(
        n34284) );
  INV_X2 U9145 ( .I(n28036), .ZN(n28189) );
  XOR2_X1 U9150 ( .A1(n34287), .A2(n20483), .Z(Ciphertext[189]) );
  XOR2_X1 U9153 ( .A1(n36746), .A2(n34288), .Z(n404) );
  XOR2_X1 U9154 ( .A1(n3703), .A2(n4816), .Z(n34288) );
  INV_X2 U9162 ( .I(n26075), .ZN(n25992) );
  XOR2_X1 U9167 ( .A1(n34289), .A2(n34703), .Z(n9509) );
  XOR2_X1 U9175 ( .A1(n33058), .A2(n19220), .Z(n19418) );
  NOR2_X1 U9177 ( .A1(n3815), .A2(n20078), .ZN(n4379) );
  NAND2_X2 U9187 ( .A1(n6116), .A2(n30993), .ZN(n16559) );
  OAI22_X1 U9188 ( .A1(n1218), .A2(n17095), .B1(n21050), .B2(n3977), .ZN(n3979) );
  XOR2_X1 U9190 ( .A1(n27735), .A2(n34290), .Z(n27841) );
  NAND2_X1 U9192 ( .A1(n27336), .A2(n27487), .ZN(n34290) );
  NAND2_X2 U9193 ( .A1(n36709), .A2(n34291), .ZN(n29070) );
  XOR2_X1 U9195 ( .A1(n2627), .A2(n27504), .Z(n34986) );
  AND2_X1 U9204 ( .A1(n29810), .A2(n29803), .Z(n29812) );
  NAND2_X1 U9253 ( .A1(n8529), .A2(n30049), .ZN(n19108) );
  AND2_X1 U9254 ( .A1(n11453), .A2(n34506), .Z(n4960) );
  OAI21_X1 U9255 ( .A1(n1340), .A2(n32478), .B(n34296), .ZN(n22308) );
  NAND2_X1 U9260 ( .A1(n32478), .A2(n22307), .ZN(n34296) );
  NOR2_X2 U9273 ( .A1(n35660), .A2(n35117), .ZN(n34297) );
  NOR2_X2 U9283 ( .A1(n1432), .A2(n28690), .ZN(n34298) );
  NAND2_X1 U9293 ( .A1(n27137), .A2(n8798), .ZN(n34299) );
  AOI21_X2 U9309 ( .A1(n13403), .A2(n11488), .B(n13401), .ZN(n34301) );
  NAND2_X1 U9319 ( .A1(n1340), .A2(n4200), .ZN(n21337) );
  NOR2_X2 U9321 ( .A1(n20740), .A2(n12306), .ZN(n15986) );
  NOR2_X2 U9324 ( .A1(n18879), .A2(n18956), .ZN(n20740) );
  OAI21_X2 U9351 ( .A1(n34303), .A2(n1564), .B(n24630), .ZN(n14768) );
  XOR2_X1 U9394 ( .A1(n34306), .A2(n3802), .Z(n26265) );
  XOR2_X1 U9395 ( .A1(n26528), .A2(n36644), .Z(n34306) );
  OAI22_X2 U9396 ( .A1(n19364), .A2(n26992), .B1(n13110), .B2(n14459), .ZN(
        n26877) );
  NOR2_X1 U9417 ( .A1(n14502), .A2(n11778), .ZN(n6018) );
  NAND3_X1 U9435 ( .A1(n4171), .A2(n12328), .A3(n32168), .ZN(n34461) );
  NAND3_X1 U9446 ( .A1(n9913), .A2(n969), .A3(n29477), .ZN(n9104) );
  NAND2_X2 U9447 ( .A1(n34559), .A2(n35203), .ZN(n13170) );
  NOR2_X2 U9469 ( .A1(n30356), .A2(n30336), .ZN(n34311) );
  NAND2_X2 U9473 ( .A1(n36526), .A2(n27356), .ZN(n27766) );
  NAND2_X2 U9474 ( .A1(n34953), .A2(n36436), .ZN(n12437) );
  BUF_X2 U9477 ( .I(n19113), .Z(n34312) );
  INV_X4 U9483 ( .I(n16853), .ZN(n1424) );
  NOR2_X2 U9491 ( .A1(n32450), .A2(n5112), .ZN(n2149) );
  OR2_X1 U9502 ( .A1(n38395), .A2(n17864), .Z(n22148) );
  XOR2_X1 U9507 ( .A1(n26221), .A2(n16497), .Z(n15821) );
  OR2_X1 U9508 ( .A1(n858), .A2(n33895), .Z(n26872) );
  XOR2_X1 U9515 ( .A1(n34314), .A2(n34313), .Z(n36602) );
  XOR2_X1 U9518 ( .A1(n31585), .A2(n29857), .Z(n34314) );
  OAI21_X2 U9527 ( .A1(n15992), .A2(n37184), .B(n15991), .ZN(n34898) );
  NOR2_X2 U9531 ( .A1(n25433), .A2(n25685), .ZN(n15992) );
  XOR2_X1 U9537 ( .A1(n17478), .A2(n34315), .Z(n24039) );
  OAI21_X2 U9544 ( .A1(n16227), .A2(n16228), .B(n20943), .ZN(n34317) );
  OAI21_X2 U9549 ( .A1(n16306), .A2(n8933), .B(n8932), .ZN(n17417) );
  OAI21_X1 U9556 ( .A1(n30118), .A2(n30119), .B(n34319), .ZN(n19031) );
  AOI22_X1 U9557 ( .A1(n19032), .A2(n10118), .B1(n19033), .B2(n16180), .ZN(
        n34319) );
  XOR2_X1 U9560 ( .A1(n29063), .A2(n29115), .Z(n14388) );
  OAI21_X2 U9565 ( .A1(n36031), .A2(n36032), .B(n28587), .ZN(n29063) );
  NAND2_X2 U9567 ( .A1(n24639), .A2(n24732), .ZN(n24843) );
  NAND2_X2 U9579 ( .A1(n20378), .A2(n36267), .ZN(n24639) );
  OAI21_X1 U9585 ( .A1(n16060), .A2(n30047), .B(n8529), .ZN(n16059) );
  XOR2_X1 U9593 ( .A1(n27469), .A2(n10866), .Z(n35834) );
  NOR2_X2 U9613 ( .A1(n31205), .A2(n26131), .ZN(n26132) );
  INV_X2 U9629 ( .I(n17618), .ZN(n14167) );
  NAND2_X2 U9630 ( .A1(n36229), .A2(n23822), .ZN(n17618) );
  XOR2_X1 U9632 ( .A1(n34323), .A2(n19432), .Z(Ciphertext[84]) );
  NAND2_X2 U9644 ( .A1(n34324), .A2(n25678), .ZN(n33909) );
  OAI22_X2 U9648 ( .A1(n25676), .A2(n14273), .B1(n25675), .B2(n19589), .ZN(
        n34324) );
  OAI21_X2 U9650 ( .A1(n15110), .A2(n28756), .B(n15109), .ZN(n15270) );
  XOR2_X1 U9656 ( .A1(n13189), .A2(n13187), .Z(n34325) );
  NAND2_X1 U9661 ( .A1(n8014), .A2(n5227), .ZN(n24943) );
  AOI22_X1 U9680 ( .A1(n6629), .A2(n8082), .B1(n35172), .B2(n19893), .ZN(
        n34326) );
  OAI21_X2 U9693 ( .A1(n35514), .A2(n38337), .B(n35513), .ZN(n19976) );
  INV_X2 U9701 ( .I(n27499), .ZN(n34332) );
  AOI21_X2 U9729 ( .A1(n5751), .A2(n19470), .B(n34329), .ZN(n3271) );
  INV_X2 U9730 ( .I(n7900), .ZN(n34329) );
  NAND2_X2 U9733 ( .A1(n21517), .A2(n261), .ZN(n7900) );
  AND2_X1 U9770 ( .A1(n14793), .A2(n36922), .Z(n36575) );
  NAND2_X2 U9785 ( .A1(n34335), .A2(n32036), .ZN(n4771) );
  AND2_X1 U9790 ( .A1(n20359), .A2(n32951), .Z(n36707) );
  XOR2_X1 U9792 ( .A1(n5694), .A2(n30907), .Z(n15047) );
  INV_X2 U9793 ( .I(n23561), .ZN(n34336) );
  NOR2_X1 U9800 ( .A1(n31078), .A2(n36380), .ZN(n19140) );
  AOI21_X2 U9814 ( .A1(n28195), .A2(n9897), .B(n34342), .ZN(n15473) );
  NAND2_X2 U9822 ( .A1(n34343), .A2(n20665), .ZN(n25175) );
  NAND3_X2 U9824 ( .A1(n30419), .A2(n17377), .A3(n20158), .ZN(n34343) );
  AOI22_X2 U9830 ( .A1(n21915), .A2(n5391), .B1(n21913), .B2(n938), .ZN(n5303)
         );
  XNOR2_X1 U9842 ( .A1(n16526), .A2(n14164), .ZN(n25285) );
  NAND2_X2 U9849 ( .A1(n1898), .A2(n30572), .ZN(n19979) );
  NOR2_X2 U9850 ( .A1(n32633), .A2(n19465), .ZN(n35452) );
  NAND2_X2 U9852 ( .A1(n7305), .A2(n2140), .ZN(n32633) );
  INV_X2 U9854 ( .I(n34347), .ZN(n15592) );
  XOR2_X1 U9862 ( .A1(n26207), .A2(n20213), .Z(n26529) );
  AOI21_X2 U9864 ( .A1(n10139), .A2(n10138), .B(n10137), .ZN(n26207) );
  XOR2_X1 U9867 ( .A1(n7060), .A2(n12988), .Z(n7059) );
  OR2_X1 U9871 ( .A1(n1190), .A2(n11296), .Z(n28634) );
  XOR2_X1 U9888 ( .A1(n34352), .A2(n5279), .Z(n33856) );
  XOR2_X1 U9894 ( .A1(n22586), .A2(n33824), .Z(n34352) );
  NAND2_X2 U9909 ( .A1(n15618), .A2(n26099), .ZN(n26421) );
  NAND2_X2 U9910 ( .A1(n16118), .A2(n16117), .ZN(n26234) );
  OR2_X1 U9911 ( .A1(n38194), .A2(n34354), .Z(n18196) );
  NAND3_X2 U9932 ( .A1(n13571), .A2(n4662), .A3(n4661), .ZN(n9873) );
  XOR2_X1 U9939 ( .A1(n4783), .A2(n14174), .Z(n27575) );
  XOR2_X1 U9947 ( .A1(n22599), .A2(n12730), .Z(n6311) );
  NAND2_X2 U9952 ( .A1(n13480), .A2(n15487), .ZN(n12730) );
  NAND2_X1 U9959 ( .A1(n30304), .A2(n13601), .ZN(n28431) );
  XOR2_X1 U9961 ( .A1(n7068), .A2(n27820), .Z(n35871) );
  OR2_X1 U9965 ( .A1(n5112), .A2(n8069), .Z(n13033) );
  XOR2_X1 U9973 ( .A1(n34358), .A2(n30839), .Z(n31121) );
  XOR2_X1 U10015 ( .A1(n9085), .A2(n38176), .Z(n26397) );
  NAND2_X2 U10026 ( .A1(n31098), .A2(n3846), .ZN(n3845) );
  XOR2_X1 U10028 ( .A1(n1884), .A2(n1885), .Z(n1883) );
  NAND2_X2 U10054 ( .A1(n28264), .A2(n28263), .ZN(n28745) );
  XOR2_X1 U10055 ( .A1(n35209), .A2(n7402), .Z(n26537) );
  INV_X2 U10080 ( .I(n34365), .ZN(n871) );
  OR2_X1 U10089 ( .A1(n30859), .A2(n4599), .Z(n26882) );
  NOR2_X2 U10092 ( .A1(n34366), .A2(n17789), .ZN(n21242) );
  XOR2_X1 U10093 ( .A1(n3292), .A2(n25065), .Z(n9781) );
  INV_X2 U10120 ( .I(n34370), .ZN(n33960) );
  XOR2_X1 U10121 ( .A1(n20693), .A2(n10169), .Z(n34370) );
  NAND2_X2 U10123 ( .A1(n34371), .A2(n13334), .ZN(n17132) );
  NOR2_X2 U10124 ( .A1(n34372), .A2(n34123), .ZN(n2288) );
  NAND3_X1 U10126 ( .A1(n31280), .A2(n31279), .A3(n12876), .ZN(n31704) );
  NAND2_X2 U10130 ( .A1(n34904), .A2(n34905), .ZN(n11950) );
  NAND2_X2 U10140 ( .A1(n966), .A2(n13192), .ZN(n13986) );
  XOR2_X1 U10147 ( .A1(n467), .A2(n29025), .Z(n34375) );
  XOR2_X1 U10166 ( .A1(n34377), .A2(n23744), .Z(n36952) );
  XOR2_X1 U10172 ( .A1(n23846), .A2(n23987), .Z(n34377) );
  NAND2_X2 U10177 ( .A1(n10553), .A2(n10551), .ZN(n36442) );
  INV_X2 U10186 ( .I(n17864), .ZN(n34379) );
  OR2_X1 U10187 ( .A1(n22238), .A2(n34379), .Z(n9524) );
  NAND2_X2 U10215 ( .A1(n34383), .A2(n9993), .ZN(n36857) );
  OAI21_X2 U10217 ( .A1(n18720), .A2(n29491), .B(n29418), .ZN(n34383) );
  NOR2_X1 U10221 ( .A1(n19985), .A2(n32164), .ZN(n34931) );
  NAND3_X2 U10223 ( .A1(n1956), .A2(n1743), .A3(n1954), .ZN(n7402) );
  NAND2_X2 U10235 ( .A1(n30929), .A2(n30930), .ZN(n33271) );
  XOR2_X1 U10240 ( .A1(n23776), .A2(n16138), .Z(n4562) );
  AND2_X1 U10242 ( .A1(n15626), .A2(n12144), .Z(n13345) );
  NAND2_X2 U10248 ( .A1(n2191), .A2(n38629), .ZN(n28580) );
  XOR2_X1 U10259 ( .A1(n33921), .A2(n34017), .Z(n824) );
  INV_X2 U10260 ( .I(n31872), .ZN(n25214) );
  XOR2_X1 U10262 ( .A1(n31872), .A2(n34391), .Z(n17834) );
  INV_X1 U10263 ( .I(n29974), .ZN(n34391) );
  NAND2_X2 U10265 ( .A1(n35785), .A2(n35784), .ZN(n31872) );
  NOR2_X2 U10267 ( .A1(n193), .A2(n20451), .ZN(n34469) );
  NAND2_X2 U10269 ( .A1(n34392), .A2(n13589), .ZN(n26134) );
  XOR2_X1 U10277 ( .A1(n34394), .A2(n30207), .Z(Ciphertext[181]) );
  NAND3_X2 U10282 ( .A1(n30205), .A2(n16548), .A3(n30206), .ZN(n34394) );
  XOR2_X1 U10310 ( .A1(n34397), .A2(n354), .Z(n32951) );
  XOR2_X1 U10315 ( .A1(n34398), .A2(n391), .Z(n36292) );
  XOR2_X1 U10317 ( .A1(n4673), .A2(n34088), .Z(n34398) );
  INV_X4 U10333 ( .I(n11628), .ZN(n1198) );
  NAND2_X2 U10383 ( .A1(n17865), .A2(n6269), .ZN(n17864) );
  NAND2_X2 U10413 ( .A1(n34405), .A2(n34404), .ZN(n30424) );
  INV_X2 U10420 ( .I(n22145), .ZN(n34404) );
  NOR2_X2 U10496 ( .A1(n7916), .A2(n22238), .ZN(n34406) );
  XOR2_X1 U10501 ( .A1(n34408), .A2(n16103), .Z(n16102) );
  NAND3_X2 U10504 ( .A1(n36403), .A2(n32668), .A3(n36402), .ZN(n29930) );
  XOR2_X1 U10505 ( .A1(n10343), .A2(n14307), .Z(n5728) );
  NAND2_X2 U10537 ( .A1(n24364), .A2(n24365), .ZN(n25181) );
  XOR2_X1 U10547 ( .A1(n19072), .A2(n20618), .Z(n32210) );
  NAND2_X1 U10558 ( .A1(n15751), .A2(n24477), .ZN(n24479) );
  NOR2_X2 U10560 ( .A1(n31159), .A2(n31158), .ZN(n35828) );
  XOR2_X1 U10568 ( .A1(n8894), .A2(n31620), .Z(n18498) );
  OR2_X1 U10570 ( .A1(n20056), .A2(n35149), .Z(n28197) );
  AND2_X1 U10573 ( .A1(n5457), .A2(n14858), .Z(n5456) );
  AOI21_X2 U10578 ( .A1(n9135), .A2(n2192), .B(n33580), .ZN(n35924) );
  AOI22_X2 U10587 ( .A1(n34857), .A2(n26055), .B1(n26054), .B2(n25424), .ZN(
        n6784) );
  NAND2_X2 U10595 ( .A1(n34415), .A2(n27994), .ZN(n28659) );
  AND2_X1 U10596 ( .A1(n27993), .A2(n27992), .Z(n34415) );
  XOR2_X1 U10614 ( .A1(n15050), .A2(n34418), .Z(n15052) );
  XOR2_X1 U10617 ( .A1(n24987), .A2(n34147), .Z(n34418) );
  NAND2_X2 U10625 ( .A1(n34420), .A2(n16374), .ZN(n35952) );
  OAI22_X2 U10663 ( .A1(n18559), .A2(n21589), .B1(n18560), .B2(n18561), .ZN(
        n22341) );
  XOR2_X1 U10666 ( .A1(n14144), .A2(n34428), .Z(n26861) );
  XOR2_X1 U10671 ( .A1(n19051), .A2(n14143), .Z(n34428) );
  XOR2_X1 U10676 ( .A1(n2218), .A2(n2217), .Z(n20686) );
  NAND2_X1 U10688 ( .A1(n4986), .A2(n16449), .ZN(n34430) );
  XOR2_X1 U10696 ( .A1(n36041), .A2(n8100), .Z(n9374) );
  XOR2_X1 U10717 ( .A1(n24049), .A2(n23757), .Z(n34435) );
  XOR2_X1 U10732 ( .A1(n19989), .A2(n19987), .Z(n28174) );
  OR2_X1 U10739 ( .A1(n24470), .A2(n15461), .Z(n36789) );
  XOR2_X1 U10745 ( .A1(n22082), .A2(n696), .Z(n18434) );
  NAND2_X2 U10750 ( .A1(n34438), .A2(n34437), .ZN(n33919) );
  NAND2_X1 U10753 ( .A1(n32760), .A2(n18926), .ZN(n21559) );
  XOR2_X1 U10756 ( .A1(n34439), .A2(n4070), .Z(n31294) );
  INV_X2 U10768 ( .I(n22588), .ZN(n34440) );
  NAND3_X2 U10777 ( .A1(n28547), .A2(n14278), .A3(n28735), .ZN(n28627) );
  NOR2_X2 U10781 ( .A1(n1752), .A2(n34446), .ZN(n34503) );
  AOI21_X1 U10790 ( .A1(n36678), .A2(n1551), .B(n371), .ZN(n3278) );
  BUF_X2 U10798 ( .I(n19417), .Z(n34447) );
  NAND2_X2 U10804 ( .A1(n32132), .A2(n32413), .ZN(n32575) );
  NOR2_X2 U10812 ( .A1(n19373), .A2(n9165), .ZN(n11364) );
  NAND2_X2 U10819 ( .A1(n32583), .A2(n34448), .ZN(n23532) );
  XOR2_X1 U10825 ( .A1(n10771), .A2(n34450), .Z(n10770) );
  XOR2_X1 U10827 ( .A1(n23968), .A2(n34451), .Z(n34450) );
  XOR2_X1 U10838 ( .A1(n34453), .A2(n12912), .Z(n12951) );
  XOR2_X1 U10855 ( .A1(n4326), .A2(n22957), .Z(n34453) );
  XOR2_X1 U10857 ( .A1(n5724), .A2(n34454), .Z(n11896) );
  XOR2_X1 U10858 ( .A1(n29821), .A2(n5728), .Z(n34454) );
  OR2_X1 U10871 ( .A1(n17917), .A2(n22921), .Z(n32133) );
  NAND2_X2 U10920 ( .A1(n35453), .A2(n20644), .ZN(n8407) );
  NAND3_X2 U10930 ( .A1(n32752), .A2(n32650), .A3(n31882), .ZN(n15855) );
  AOI21_X2 U10937 ( .A1(n36850), .A2(n12273), .B(n12272), .ZN(n34460) );
  NAND2_X2 U10940 ( .A1(n34995), .A2(n20172), .ZN(n7044) );
  AOI22_X2 U10950 ( .A1(n11713), .A2(n11712), .B1(n11711), .B2(n10013), .ZN(
        n19156) );
  XOR2_X1 U10958 ( .A1(n25127), .A2(n25177), .Z(n25217) );
  OAI21_X1 U10964 ( .A1(n22975), .A2(n34467), .B(n34466), .ZN(n23087) );
  NAND2_X1 U10966 ( .A1(n34467), .A2(n23167), .ZN(n34466) );
  XOR2_X1 U10967 ( .A1(n34468), .A2(n34104), .Z(n35687) );
  AOI21_X2 U10985 ( .A1(n37279), .A2(n23559), .B(n34336), .ZN(n34472) );
  INV_X2 U10990 ( .I(n34473), .ZN(n33579) );
  INV_X2 U11005 ( .I(n17597), .ZN(n12940) );
  NAND3_X1 U11013 ( .A1(n15080), .A2(n15081), .A3(n19538), .ZN(n15079) );
  XOR2_X1 U11017 ( .A1(n17430), .A2(n34474), .Z(n17830) );
  XOR2_X1 U11018 ( .A1(n12125), .A2(n17429), .Z(n34474) );
  NAND2_X1 U11020 ( .A1(n19631), .A2(n1195), .ZN(n12336) );
  NAND2_X2 U11021 ( .A1(n11280), .A2(n11279), .ZN(n1195) );
  INV_X4 U11022 ( .I(n33579), .ZN(n35314) );
  INV_X4 U11023 ( .I(n34475), .ZN(n22324) );
  NAND2_X1 U11040 ( .A1(n20948), .A2(n20949), .ZN(n34476) );
  OAI22_X1 U11045 ( .A1(n21302), .A2(n17246), .B1(n955), .B2(n826), .ZN(n15543) );
  AND2_X1 U11046 ( .A1(n4377), .A2(n4378), .Z(n4168) );
  XOR2_X1 U11047 ( .A1(n34477), .A2(n32604), .Z(n28848) );
  XOR2_X1 U11058 ( .A1(n17797), .A2(n34478), .Z(n31261) );
  NAND2_X2 U11066 ( .A1(n34480), .A2(n4504), .ZN(n16619) );
  NAND2_X2 U11070 ( .A1(n6747), .A2(n20441), .ZN(n25435) );
  XNOR2_X1 U11073 ( .A1(n5816), .A2(n5815), .ZN(n34483) );
  XOR2_X1 U11076 ( .A1(n23926), .A2(n23925), .Z(n1929) );
  NAND3_X1 U11088 ( .A1(n32497), .A2(n6578), .A3(n9530), .ZN(n34486) );
  XOR2_X1 U11094 ( .A1(n21284), .A2(n27720), .Z(n18049) );
  XOR2_X1 U11096 ( .A1(n27773), .A2(n27503), .Z(n21284) );
  XOR2_X1 U11101 ( .A1(n26364), .A2(n26336), .Z(n9555) );
  XOR2_X1 U11104 ( .A1(n1009), .A2(n7133), .Z(n26364) );
  NAND2_X2 U11135 ( .A1(n28299), .A2(n16303), .ZN(n28301) );
  NOR2_X2 U11137 ( .A1(n13323), .A2(n13321), .ZN(n16303) );
  NOR2_X1 U11139 ( .A1(n34561), .A2(n24287), .ZN(n14684) );
  XOR2_X1 U11146 ( .A1(n5610), .A2(n26514), .Z(n34489) );
  OAI22_X1 U11149 ( .A1(n19564), .A2(n1478), .B1(n18246), .B2(n1085), .ZN(
        n7232) );
  NAND2_X1 U11150 ( .A1(n35881), .A2(n19587), .ZN(n5533) );
  NOR2_X2 U11154 ( .A1(n4317), .A2(n22157), .ZN(n6582) );
  XOR2_X1 U11168 ( .A1(n3376), .A2(n3375), .Z(n24192) );
  INV_X2 U11171 ( .I(n34490), .ZN(n30454) );
  XOR2_X1 U11173 ( .A1(n15860), .A2(n15859), .Z(n34490) );
  NAND2_X2 U11175 ( .A1(n36947), .A2(n28964), .ZN(n13192) );
  XOR2_X1 U11176 ( .A1(n15220), .A2(n25198), .Z(n3185) );
  AOI22_X2 U11177 ( .A1(n2930), .A2(n20168), .B1(n31568), .B2(n25242), .ZN(
        n15220) );
  XOR2_X1 U11191 ( .A1(n5347), .A2(n33478), .Z(n5348) );
  BUF_X2 U11193 ( .I(n33609), .Z(n34494) );
  XOR2_X1 U11194 ( .A1(n26335), .A2(n34495), .Z(n19533) );
  XOR2_X1 U11198 ( .A1(n26585), .A2(n34768), .Z(n26335) );
  NOR2_X2 U11203 ( .A1(n32853), .A2(n32852), .ZN(n27574) );
  NOR3_X1 U11207 ( .A1(n35588), .A2(n34622), .A3(n30004), .ZN(n30008) );
  INV_X2 U11217 ( .I(n34496), .ZN(n19891) );
  XNOR2_X1 U11219 ( .A1(n9039), .A2(n8781), .ZN(n34496) );
  XOR2_X1 U11221 ( .A1(n3773), .A2(n34497), .Z(n10620) );
  XOR2_X1 U11222 ( .A1(n33672), .A2(n34498), .Z(n34497) );
  NAND2_X2 U11228 ( .A1(n29237), .A2(n3263), .ZN(n29228) );
  NAND2_X2 U11231 ( .A1(n16839), .A2(n29079), .ZN(n29237) );
  XOR2_X1 U11238 ( .A1(n8474), .A2(n2371), .Z(n2370) );
  NAND2_X1 U11241 ( .A1(n6248), .A2(n25328), .ZN(n34501) );
  NAND2_X2 U11256 ( .A1(n34503), .A2(n14790), .ZN(n13151) );
  NAND2_X2 U11264 ( .A1(n13970), .A2(n1123), .ZN(n34504) );
  NOR2_X2 U11265 ( .A1(n36683), .A2(n26), .ZN(n16578) );
  NOR2_X2 U11267 ( .A1(n16407), .A2(n25961), .ZN(n25923) );
  INV_X2 U11282 ( .I(n9920), .ZN(n34506) );
  AOI22_X2 U11294 ( .A1(n38011), .A2(n5451), .B1(n17249), .B2(n938), .ZN(n5776) );
  NAND2_X2 U11298 ( .A1(n2566), .A2(n28693), .ZN(n31127) );
  XOR2_X1 U11305 ( .A1(n19766), .A2(n16362), .Z(n3890) );
  NAND2_X2 U11322 ( .A1(n35899), .A2(n17997), .ZN(n11968) );
  XOR2_X1 U11323 ( .A1(n476), .A2(n39575), .Z(n20016) );
  NAND2_X2 U11328 ( .A1(n35012), .A2(n23485), .ZN(n476) );
  XOR2_X1 U11332 ( .A1(n35227), .A2(n27845), .Z(n27605) );
  NAND2_X2 U11333 ( .A1(n22493), .A2(n6176), .ZN(n23480) );
  NOR2_X2 U11338 ( .A1(n28207), .A2(n7541), .ZN(n28720) );
  AOI22_X2 U11343 ( .A1(n16308), .A2(n19754), .B1(n5396), .B2(n34510), .ZN(
        n20319) );
  OAI21_X1 U11344 ( .A1(n1222), .A2(n15284), .B(n27197), .ZN(n6508) );
  XOR2_X1 U11349 ( .A1(n25310), .A2(n6232), .Z(n6231) );
  XOR2_X1 U11350 ( .A1(n34091), .A2(n3776), .Z(n35129) );
  AOI21_X2 U11357 ( .A1(n34512), .A2(n32333), .B(n37008), .ZN(n37007) );
  AOI21_X2 U11370 ( .A1(n16201), .A2(n36722), .B(n11668), .ZN(n26556) );
  XOR2_X1 U11372 ( .A1(n34514), .A2(n17707), .Z(n10039) );
  XOR2_X1 U11379 ( .A1(n30318), .A2(n24873), .Z(n34514) );
  XOR2_X1 U11390 ( .A1(n8284), .A2(n30994), .Z(n11782) );
  XOR2_X1 U11401 ( .A1(n34518), .A2(n30423), .Z(n32838) );
  NOR2_X1 U11404 ( .A1(n25957), .A2(n18406), .ZN(n34519) );
  OAI22_X2 U11407 ( .A1(n29782), .A2(n16682), .B1(n19716), .B2(n3096), .ZN(
        n29798) );
  XOR2_X1 U11421 ( .A1(n20065), .A2(n215), .Z(n35269) );
  XOR2_X1 U11426 ( .A1(n20540), .A2(n7474), .Z(n215) );
  INV_X2 U11436 ( .I(n34521), .ZN(n37050) );
  XNOR2_X1 U11437 ( .A1(n35510), .A2(n13938), .ZN(n34521) );
  NAND2_X2 U11440 ( .A1(n25593), .A2(n19401), .ZN(n25961) );
  NAND2_X2 U11461 ( .A1(n22919), .A2(n23072), .ZN(n34557) );
  NAND3_X2 U11464 ( .A1(n15836), .A2(n6450), .A3(n16259), .ZN(n9719) );
  INV_X1 U11466 ( .I(n34522), .ZN(n23143) );
  NOR2_X1 U11468 ( .A1(n8765), .A2(n34522), .ZN(n5628) );
  AOI21_X2 U11470 ( .A1(n32248), .A2(n12263), .B(n12427), .ZN(n8894) );
  NOR2_X2 U11472 ( .A1(n826), .A2(n37050), .ZN(n25602) );
  OAI21_X2 U11479 ( .A1(n33892), .A2(n33891), .B(n25911), .ZN(n34768) );
  AOI21_X1 U11480 ( .A1(n10479), .A2(n17515), .B(n9690), .ZN(n17514) );
  NOR2_X2 U11509 ( .A1(n32358), .A2(n31465), .ZN(n2600) );
  INV_X2 U11523 ( .I(n34532), .ZN(n26724) );
  XOR2_X1 U11527 ( .A1(n19021), .A2(n19018), .Z(n34532) );
  AOI22_X2 U11528 ( .A1(n34533), .A2(n1523), .B1(n5475), .B2(n5886), .ZN(n5474) );
  OAI22_X1 U11546 ( .A1(n29511), .A2(n35180), .B1(n29524), .B2(n29531), .ZN(
        n29512) );
  XOR2_X1 U11564 ( .A1(n35227), .A2(n14808), .Z(n27806) );
  AOI21_X2 U11565 ( .A1(n27073), .A2(n18228), .B(n30933), .ZN(n35227) );
  NAND2_X2 U11574 ( .A1(n6554), .A2(n34540), .ZN(n10461) );
  AOI22_X2 U11576 ( .A1(n6312), .A2(n441), .B1(n6313), .B2(n18809), .ZN(n34540) );
  INV_X2 U11607 ( .I(n34546), .ZN(n16692) );
  XNOR2_X1 U11608 ( .A1(n22605), .A2(n33856), .ZN(n34546) );
  INV_X4 U11610 ( .I(n9193), .ZN(n1034) );
  NAND2_X1 U11618 ( .A1(n692), .A2(n9833), .ZN(n16240) );
  BUF_X2 U11623 ( .I(n35233), .Z(n34547) );
  XOR2_X1 U11638 ( .A1(n18490), .A2(n26519), .Z(n12429) );
  INV_X2 U11648 ( .I(n34549), .ZN(n36197) );
  XOR2_X1 U11655 ( .A1(n33112), .A2(n33111), .Z(n34549) );
  AOI21_X1 U11667 ( .A1(n11111), .A2(n19108), .B(n29935), .ZN(n10097) );
  XOR2_X1 U11668 ( .A1(n34552), .A2(n29849), .Z(Ciphertext[114]) );
  NAND2_X2 U11673 ( .A1(n36555), .A2(n34554), .ZN(n7481) );
  XOR2_X1 U11676 ( .A1(n27847), .A2(n35678), .Z(n16607) );
  INV_X4 U11690 ( .I(n33952), .ZN(n36262) );
  OAI21_X2 U11691 ( .A1(n34072), .A2(n22919), .B(n34557), .ZN(n22828) );
  AOI21_X2 U11701 ( .A1(n6654), .A2(n13685), .B(n13684), .ZN(n13683) );
  XOR2_X1 U11703 ( .A1(n23830), .A2(n23804), .Z(n6530) );
  XOR2_X1 U11709 ( .A1(n26396), .A2(n3781), .Z(n26205) );
  NOR2_X1 U11717 ( .A1(n32682), .A2(n36935), .ZN(n34568) );
  AND2_X1 U11718 ( .A1(n36323), .A2(n25601), .Z(n35632) );
  NOR2_X1 U11728 ( .A1(n32059), .A2(n10254), .ZN(n34569) );
  XOR2_X1 U11738 ( .A1(n4223), .A2(n4221), .Z(n30233) );
  NAND2_X2 U11745 ( .A1(n31028), .A2(n34571), .ZN(n9413) );
  INV_X2 U11752 ( .I(n12234), .ZN(n34574) );
  XOR2_X1 U11755 ( .A1(n17593), .A2(n25087), .Z(n12311) );
  INV_X2 U11757 ( .I(n34957), .ZN(n26905) );
  AOI21_X2 U11767 ( .A1(n34575), .A2(n19402), .B(n9371), .ZN(n33108) );
  NAND2_X2 U11770 ( .A1(n6515), .A2(n33599), .ZN(n34575) );
  INV_X2 U11786 ( .I(n37085), .ZN(n13166) );
  NAND2_X1 U11787 ( .A1(n37085), .A2(n34576), .ZN(n19463) );
  XOR2_X1 U11790 ( .A1(n35645), .A2(n12293), .Z(n18507) );
  XNOR2_X1 U11794 ( .A1(n26566), .A2(n20139), .ZN(n34593) );
  AND2_X1 U11797 ( .A1(n26905), .A2(n39477), .Z(n9423) );
  NAND2_X1 U11806 ( .A1(n6415), .A2(n9267), .ZN(n6414) );
  NAND2_X2 U11808 ( .A1(n3918), .A2(n12887), .ZN(n9267) );
  XOR2_X1 U11820 ( .A1(n34580), .A2(n18852), .Z(n13127) );
  OAI21_X2 U11823 ( .A1(n14695), .A2(n3783), .B(n38305), .ZN(n21139) );
  XOR2_X1 U11828 ( .A1(n2431), .A2(n38167), .Z(n32512) );
  NOR3_X2 U11831 ( .A1(n1541), .A2(n6300), .A3(n34010), .ZN(n34581) );
  XOR2_X1 U11837 ( .A1(n32298), .A2(n35243), .Z(n4815) );
  NOR2_X2 U11870 ( .A1(n34801), .A2(n12651), .ZN(n12650) );
  XOR2_X1 U11885 ( .A1(n27864), .A2(n10653), .Z(n9160) );
  XOR2_X1 U11888 ( .A1(n34586), .A2(n23755), .Z(n12520) );
  INV_X2 U11922 ( .I(n34587), .ZN(n15922) );
  NAND2_X2 U11950 ( .A1(n13911), .A2(n13909), .ZN(n22511) );
  XOR2_X1 U11957 ( .A1(n3705), .A2(n3707), .Z(n4386) );
  XOR2_X1 U11958 ( .A1(n23734), .A2(n23662), .Z(n11724) );
  AOI22_X2 U11961 ( .A1(n34589), .A2(n30225), .B1(n30222), .B2(n30223), .ZN(
        n30259) );
  XOR2_X1 U11978 ( .A1(n23419), .A2(n9344), .Z(n23830) );
  OR2_X1 U11989 ( .A1(n10375), .A2(n10334), .Z(n10377) );
  NAND2_X1 U11994 ( .A1(n30647), .A2(n30646), .ZN(n34750) );
  XOR2_X1 U11996 ( .A1(n32844), .A2(n34593), .Z(n30989) );
  OR2_X1 U11998 ( .A1(n25923), .A2(n25922), .Z(n15378) );
  XOR2_X1 U11999 ( .A1(n16085), .A2(n27161), .Z(n4364) );
  AND2_X1 U12004 ( .A1(n24538), .A2(n35893), .Z(n35119) );
  NOR2_X2 U12035 ( .A1(n17476), .A2(n34596), .ZN(n28578) );
  INV_X2 U12044 ( .I(n34597), .ZN(n31010) );
  XNOR2_X1 U12050 ( .A1(n33044), .A2(n11103), .ZN(n34597) );
  NOR2_X1 U12057 ( .A1(n31010), .A2(n9740), .ZN(n8494) );
  INV_X2 U12058 ( .I(n36226), .ZN(n1097) );
  NAND2_X1 U12068 ( .A1(n8158), .A2(n8159), .ZN(n8157) );
  NAND2_X1 U12072 ( .A1(n35745), .A2(n34279), .ZN(n20143) );
  XOR2_X1 U12081 ( .A1(n33400), .A2(n39320), .Z(n33399) );
  OAI21_X2 U12103 ( .A1(n4466), .A2(n4465), .B(n4464), .ZN(n26090) );
  NOR2_X2 U12112 ( .A1(n34599), .A2(n35935), .ZN(n29166) );
  NAND2_X1 U12126 ( .A1(n13082), .A2(n32638), .ZN(n27974) );
  BUF_X2 U12132 ( .I(Key[67]), .Z(n29879) );
  AOI22_X1 U12144 ( .A1(n29890), .A2(n32706), .B1(n17286), .B2(n11182), .ZN(
        n11785) );
  AOI22_X2 U12149 ( .A1(n6703), .A2(n11412), .B1(n9443), .B2(n5890), .ZN(n9442) );
  BUF_X2 U12155 ( .I(n28616), .Z(n314) );
  XOR2_X1 U12164 ( .A1(n20447), .A2(n2824), .Z(n29120) );
  NAND2_X2 U12197 ( .A1(n36131), .A2(n36130), .ZN(n34602) );
  NAND2_X2 U12200 ( .A1(n11907), .A2(n20657), .ZN(n24938) );
  OR2_X2 U12214 ( .A1(n30853), .A2(n26832), .Z(n26835) );
  NAND2_X2 U12223 ( .A1(n25867), .A2(n26048), .ZN(n26021) );
  XOR2_X1 U12226 ( .A1(n6379), .A2(n34604), .Z(n2394) );
  XOR2_X1 U12227 ( .A1(n23669), .A2(n23668), .Z(n34604) );
  NOR2_X2 U12239 ( .A1(n27389), .A2(n21272), .ZN(n20871) );
  NAND2_X1 U12248 ( .A1(n20018), .A2(n35217), .ZN(n15712) );
  XOR2_X1 U12255 ( .A1(n27714), .A2(n184), .Z(n183) );
  XOR2_X1 U12256 ( .A1(n27525), .A2(n27834), .Z(n27714) );
  NAND3_X2 U12290 ( .A1(n7483), .A2(n28154), .A3(n17818), .ZN(n31597) );
  NAND2_X2 U12295 ( .A1(n33481), .A2(n18770), .ZN(n17818) );
  NOR2_X1 U12303 ( .A1(n35608), .A2(n39628), .ZN(n34608) );
  NAND2_X2 U12304 ( .A1(n10176), .A2(n399), .ZN(n27724) );
  INV_X2 U12332 ( .I(n34610), .ZN(n32080) );
  XOR2_X1 U12346 ( .A1(n13116), .A2(n34611), .Z(n19223) );
  NAND2_X1 U12363 ( .A1(n30588), .A2(n19334), .ZN(n30587) );
  NAND2_X2 U12379 ( .A1(n34615), .A2(n4690), .ZN(n23577) );
  XOR2_X1 U12387 ( .A1(n34616), .A2(n11503), .Z(n17210) );
  OAI22_X1 U12404 ( .A1(n30257), .A2(n30259), .B1(n30262), .B2(n38204), .ZN(
        n30263) );
  NAND2_X1 U12407 ( .A1(n28543), .A2(n28739), .ZN(n5969) );
  NAND2_X2 U12416 ( .A1(n16530), .A2(n17522), .ZN(n28543) );
  BUF_X2 U12421 ( .I(n18619), .Z(n34620) );
  XOR2_X1 U12426 ( .A1(n27527), .A2(n27567), .Z(n15400) );
  XOR2_X1 U12431 ( .A1(n15401), .A2(n8364), .Z(n27567) );
  NAND2_X2 U12453 ( .A1(n7469), .A2(n7468), .ZN(n36200) );
  NAND2_X2 U12463 ( .A1(n20768), .A2(n20770), .ZN(n26585) );
  AOI21_X1 U12479 ( .A1(n18780), .A2(n30014), .B(n30034), .ZN(n34622) );
  OAI22_X2 U12491 ( .A1(n33234), .A2(n33235), .B1(n35495), .B2(n27419), .ZN(
        n27737) );
  NOR2_X1 U12504 ( .A1(n17632), .A2(n17240), .ZN(n35063) );
  NAND2_X1 U12507 ( .A1(n19312), .A2(n35063), .ZN(n6921) );
  NAND2_X1 U12516 ( .A1(n21897), .A2(n11576), .ZN(n5733) );
  NOR2_X2 U12520 ( .A1(n34627), .A2(n8635), .ZN(n29044) );
  NAND2_X2 U12541 ( .A1(n8399), .A2(n18457), .ZN(n3263) );
  AOI22_X2 U12542 ( .A1(n1820), .A2(n15712), .B1(n8918), .B2(n34761), .ZN(
        n8399) );
  NAND3_X2 U12552 ( .A1(n9237), .A2(n9236), .A3(n15727), .ZN(n20445) );
  XOR2_X1 U12554 ( .A1(n254), .A2(n39691), .Z(n34630) );
  AND2_X1 U12557 ( .A1(n20056), .A2(n18186), .Z(n15694) );
  NAND2_X2 U12565 ( .A1(n12852), .A2(n11007), .ZN(n32208) );
  NAND2_X2 U12566 ( .A1(n1159), .A2(n17242), .ZN(n12852) );
  XOR2_X1 U12589 ( .A1(n27827), .A2(n34634), .Z(n19467) );
  XOR2_X1 U12593 ( .A1(n27826), .A2(n11031), .Z(n34634) );
  NOR2_X2 U12599 ( .A1(n34357), .A2(n39194), .ZN(n11468) );
  AOI22_X2 U12605 ( .A1(n34639), .A2(n34638), .B1(n28378), .B2(n28098), .ZN(
        n4197) );
  NAND2_X2 U12608 ( .A1(n29011), .A2(n20219), .ZN(n8287) );
  NOR2_X2 U12610 ( .A1(n7855), .A2(n34641), .ZN(n4847) );
  INV_X1 U12618 ( .I(n34642), .ZN(n34641) );
  NOR2_X2 U12622 ( .A1(n32326), .A2(n32327), .ZN(n35715) );
  NAND3_X1 U12625 ( .A1(n28246), .A2(n39399), .A3(n28115), .ZN(n32413) );
  XOR2_X1 U12627 ( .A1(n36379), .A2(n24009), .Z(n24316) );
  NAND2_X2 U12650 ( .A1(n6647), .A2(n1315), .ZN(n14006) );
  XOR2_X1 U12656 ( .A1(n29258), .A2(n34649), .Z(n13288) );
  XOR2_X1 U12664 ( .A1(n34650), .A2(n33313), .Z(n10255) );
  OR2_X1 U12670 ( .A1(n24383), .A2(n18402), .Z(n6569) );
  NAND3_X2 U12676 ( .A1(n18095), .A2(n1494), .A3(n20211), .ZN(n20217) );
  OAI21_X2 U12683 ( .A1(n979), .A2(n38075), .B(n28570), .ZN(n34651) );
  NAND2_X2 U12687 ( .A1(n3253), .A2(n32430), .ZN(n14374) );
  OAI22_X2 U12691 ( .A1(n5075), .A2(n36457), .B1(n8204), .B2(n32889), .ZN(
        n34654) );
  NOR2_X2 U12692 ( .A1(n37187), .A2(n34655), .ZN(n9581) );
  XOR2_X1 U12693 ( .A1(n15532), .A2(n8671), .Z(n8670) );
  XOR2_X1 U12695 ( .A1(n22588), .A2(n5242), .Z(n7137) );
  NAND2_X2 U12699 ( .A1(n4497), .A2(n35193), .ZN(n5242) );
  INV_X2 U12700 ( .I(n12718), .ZN(n1190) );
  OAI21_X2 U12701 ( .A1(n9850), .A2(n9684), .B(n12420), .ZN(n12718) );
  NAND2_X2 U12709 ( .A1(n23308), .A2(n23607), .ZN(n23413) );
  NAND2_X2 U12711 ( .A1(n35715), .A2(n23007), .ZN(n23308) );
  BUF_X2 U12716 ( .I(n11950), .Z(n35404) );
  NAND2_X2 U12731 ( .A1(n28427), .A2(n1194), .ZN(n28394) );
  OR2_X1 U12746 ( .A1(n1414), .A2(n2191), .Z(n30740) );
  XOR2_X1 U12749 ( .A1(n22723), .A2(n34663), .Z(n4738) );
  XOR2_X1 U12751 ( .A1(n15765), .A2(n22762), .Z(n34663) );
  NAND2_X2 U12769 ( .A1(n14924), .A2(n14926), .ZN(n36750) );
  AOI22_X1 U12776 ( .A1(n11022), .A2(n14512), .B1(n30263), .B2(n8691), .ZN(
        n34778) );
  BUF_X2 U12789 ( .I(n2052), .Z(n35253) );
  INV_X1 U12793 ( .I(n20865), .ZN(n35879) );
  NAND2_X2 U12804 ( .A1(n30689), .A2(n4485), .ZN(n34717) );
  NAND2_X2 U12808 ( .A1(n29885), .A2(n6720), .ZN(n29880) );
  INV_X4 U12823 ( .I(n28033), .ZN(n987) );
  AOI21_X2 U12826 ( .A1(n30285), .A2(n26882), .B(n37104), .ZN(n34669) );
  OAI21_X2 U12828 ( .A1(n34671), .A2(n34667), .B(n34670), .ZN(n28416) );
  INV_X1 U12829 ( .I(n28577), .ZN(n34671) );
  XOR2_X1 U12831 ( .A1(n20452), .A2(n34672), .Z(n35633) );
  INV_X1 U12835 ( .I(n29399), .ZN(n34672) );
  OR2_X1 U12856 ( .A1(n18619), .A2(n12138), .Z(n12801) );
  OAI22_X1 U12866 ( .A1(n16513), .A2(n5469), .B1(n5470), .B2(n21239), .ZN(
        n6588) );
  XOR2_X1 U12869 ( .A1(n5289), .A2(n8473), .Z(n12401) );
  OAI22_X2 U12874 ( .A1(n19588), .A2(n14561), .B1(n15388), .B2(n4472), .ZN(
        n15743) );
  XOR2_X1 U12877 ( .A1(n11383), .A2(n23829), .Z(n23943) );
  BUF_X2 U12885 ( .I(n22491), .Z(n34678) );
  XOR2_X1 U12886 ( .A1(n15448), .A2(n19717), .Z(n22466) );
  XOR2_X1 U12894 ( .A1(n30560), .A2(n34680), .Z(n5351) );
  XOR2_X1 U12896 ( .A1(n4266), .A2(n27825), .Z(n34680) );
  OR2_X1 U12897 ( .A1(n27624), .A2(n28153), .Z(n9721) );
  OAI21_X2 U12899 ( .A1(n16589), .A2(n30052), .B(n34681), .ZN(n18896) );
  XNOR2_X1 U12913 ( .A1(n1859), .A2(n27701), .ZN(n27089) );
  XOR2_X1 U12918 ( .A1(n27633), .A2(n27799), .Z(n27701) );
  NOR2_X2 U12922 ( .A1(n1220), .A2(n31683), .ZN(n34682) );
  AOI22_X1 U12932 ( .A1(n31326), .A2(n29990), .B1(n4011), .B2(n30045), .ZN(
        n30141) );
  NOR2_X2 U12941 ( .A1(n8423), .A2(n28740), .ZN(n1874) );
  XOR2_X1 U12947 ( .A1(n27605), .A2(n31248), .Z(n34686) );
  NAND2_X2 U12949 ( .A1(n29189), .A2(n34688), .ZN(n29754) );
  NAND2_X2 U12951 ( .A1(n3248), .A2(n3250), .ZN(n36913) );
  NOR2_X2 U12954 ( .A1(n36246), .A2(n13820), .ZN(n3248) );
  XOR2_X1 U12966 ( .A1(n34691), .A2(n9719), .Z(n22416) );
  OAI21_X2 U12979 ( .A1(n11735), .A2(n4463), .B(n4462), .ZN(n27710) );
  XOR2_X1 U12986 ( .A1(n23760), .A2(n16337), .Z(n23761) );
  INV_X2 U13010 ( .I(n10986), .ZN(n10724) );
  OAI21_X2 U13022 ( .A1(n33973), .A2(n34696), .B(n8806), .ZN(n7577) );
  XOR2_X1 U13028 ( .A1(n13840), .A2(n34697), .Z(n12961) );
  XOR2_X1 U13029 ( .A1(n13842), .A2(n34698), .Z(n34697) );
  OR2_X1 U13041 ( .A1(n690), .A2(n8736), .Z(n20682) );
  INV_X2 U13045 ( .I(n34699), .ZN(n15839) );
  XOR2_X1 U13046 ( .A1(Plaintext[92]), .A2(Key[92]), .Z(n34699) );
  NAND3_X2 U13049 ( .A1(n13137), .A2(n12473), .A3(n12472), .ZN(n23423) );
  OR2_X1 U13054 ( .A1(n22354), .A2(n22353), .Z(n22209) );
  NAND2_X2 U13062 ( .A1(n27004), .A2(n35914), .ZN(n27834) );
  NOR2_X1 U13072 ( .A1(n19364), .A2(n26879), .ZN(n26609) );
  NAND2_X2 U13082 ( .A1(n19413), .A2(n35124), .ZN(n4232) );
  NAND2_X1 U13094 ( .A1(n22051), .A2(n22307), .ZN(n30613) );
  XOR2_X1 U13101 ( .A1(n19355), .A2(n27729), .Z(n31204) );
  NAND2_X2 U13106 ( .A1(n18073), .A2(n18075), .ZN(n27729) );
  XOR2_X1 U13108 ( .A1(n9511), .A2(n22641), .Z(n34703) );
  INV_X1 U13109 ( .I(n39194), .ZN(n9924) );
  OR2_X1 U13110 ( .A1(n39194), .A2(n12966), .Z(n17958) );
  XOR2_X1 U13114 ( .A1(n10812), .A2(n10811), .Z(n29174) );
  XOR2_X1 U13115 ( .A1(n7004), .A2(n29082), .Z(n10811) );
  XOR2_X1 U13123 ( .A1(n34709), .A2(n34708), .Z(n14641) );
  XOR2_X1 U13125 ( .A1(n31438), .A2(n27815), .Z(n34709) );
  NAND2_X2 U13136 ( .A1(n34711), .A2(n34210), .ZN(n34820) );
  NAND2_X2 U13142 ( .A1(n23596), .A2(n23595), .ZN(n3006) );
  AOI21_X2 U13145 ( .A1(n36701), .A2(n36011), .B(n1160), .ZN(n12821) );
  XOR2_X1 U13148 ( .A1(n34712), .A2(n26417), .Z(n33473) );
  AOI21_X2 U13181 ( .A1(n22956), .A2(n34457), .B(n34716), .ZN(n5619) );
  BUF_X2 U13188 ( .I(n22561), .Z(n34718) );
  AOI22_X2 U13197 ( .A1(n11528), .A2(n1038), .B1(n17454), .B2(n23515), .ZN(
        n13978) );
  XOR2_X1 U13213 ( .A1(n14986), .A2(n8182), .Z(n8181) );
  XOR2_X1 U13227 ( .A1(n7402), .A2(n31791), .Z(n8902) );
  XOR2_X1 U13244 ( .A1(n26356), .A2(n18004), .Z(n14784) );
  OAI21_X2 U13248 ( .A1(n5508), .A2(n32052), .B(n32051), .ZN(n18004) );
  XOR2_X1 U13254 ( .A1(n6943), .A2(n6940), .Z(n35242) );
  NOR2_X2 U13257 ( .A1(n7423), .A2(n26120), .ZN(n26013) );
  XOR2_X1 U13262 ( .A1(n12383), .A2(n8310), .Z(n34722) );
  INV_X1 U13268 ( .I(n34723), .ZN(n24786) );
  NOR2_X1 U13270 ( .A1(n35686), .A2(n37016), .ZN(n34723) );
  XOR2_X1 U13290 ( .A1(n19342), .A2(n34724), .Z(n13694) );
  XOR2_X1 U13296 ( .A1(n13844), .A2(n32420), .Z(n34724) );
  XOR2_X1 U13321 ( .A1(n35554), .A2(n20684), .Z(n170) );
  NAND2_X2 U13322 ( .A1(n25900), .A2(n25801), .ZN(n25751) );
  XOR2_X1 U13324 ( .A1(n34728), .A2(n37129), .Z(n5520) );
  XOR2_X1 U13326 ( .A1(n27554), .A2(n1703), .Z(n34728) );
  NAND2_X2 U13333 ( .A1(n37031), .A2(n2883), .ZN(n3528) );
  NOR2_X1 U13347 ( .A1(n11658), .A2(n11582), .ZN(n11659) );
  XOR2_X1 U13348 ( .A1(n2594), .A2(n26395), .Z(n36719) );
  XOR2_X1 U13351 ( .A1(n39078), .A2(n7439), .Z(n26395) );
  OAI21_X2 U13384 ( .A1(n34747), .A2(n34746), .B(n24843), .ZN(n3629) );
  AOI21_X1 U13387 ( .A1(n16803), .A2(n29890), .B(n10848), .ZN(n17527) );
  INV_X2 U13388 ( .I(n6720), .ZN(n10848) );
  XOR2_X1 U13389 ( .A1(n10987), .A2(n30733), .Z(n6457) );
  NAND3_X1 U13407 ( .A1(n36789), .A2(n36790), .A3(n16377), .ZN(n36267) );
  XOR2_X1 U13409 ( .A1(n9979), .A2(n7185), .Z(n31773) );
  XOR2_X1 U13411 ( .A1(n11372), .A2(n29141), .Z(n562) );
  NAND2_X2 U13418 ( .A1(n24089), .A2(n34750), .ZN(n24879) );
  OAI21_X2 U13422 ( .A1(n34751), .A2(n19349), .B(n7480), .ZN(n18364) );
  XOR2_X1 U13429 ( .A1(n2096), .A2(n30489), .Z(n2094) );
  XOR2_X1 U13434 ( .A1(n38201), .A2(n19862), .Z(n30519) );
  BUF_X4 U13448 ( .I(n27575), .Z(n28290) );
  XOR2_X1 U13456 ( .A1(n26288), .A2(n26287), .Z(n34752) );
  NOR3_X1 U13482 ( .A1(n35253), .A2(n18402), .A3(n24382), .ZN(n34758) );
  XNOR2_X1 U13488 ( .A1(n15219), .A2(n27574), .ZN(n27677) );
  XOR2_X1 U13495 ( .A1(n34760), .A2(n34056), .Z(n33347) );
  XOR2_X1 U13497 ( .A1(n27643), .A2(n27497), .Z(n34760) );
  AND2_X1 U13504 ( .A1(n27341), .A2(n27338), .Z(n4668) );
  AOI22_X2 U13518 ( .A1(n27909), .A2(n28298), .B1(n28268), .B2(n28301), .ZN(
        n28790) );
  OAI22_X2 U13522 ( .A1(n27907), .A2(n28753), .B1(n16303), .B2(n27908), .ZN(
        n28268) );
  XOR2_X1 U13523 ( .A1(n20571), .A2(n19809), .Z(n25694) );
  XOR2_X1 U13525 ( .A1(n27769), .A2(n27798), .Z(n2758) );
  AOI22_X2 U13531 ( .A1(n35417), .A2(n35694), .B1(n37056), .B2(n28004), .ZN(
        n34762) );
  INV_X4 U13539 ( .I(n11867), .ZN(n5130) );
  XOR2_X1 U13542 ( .A1(n248), .A2(n15270), .Z(n28867) );
  NAND2_X2 U13545 ( .A1(n10148), .A2(n34763), .ZN(n33813) );
  INV_X2 U13548 ( .I(n34764), .ZN(n31669) );
  XOR2_X1 U13566 ( .A1(n3649), .A2(n34766), .Z(n9033) );
  OAI21_X1 U13569 ( .A1(n9032), .A2(n12846), .B(n9031), .ZN(n34766) );
  XOR2_X1 U13575 ( .A1(n26548), .A2(n26541), .Z(n34878) );
  AOI22_X2 U13586 ( .A1(n34767), .A2(n20423), .B1(n26973), .B2(n16000), .ZN(
        n15999) );
  XOR2_X1 U13612 ( .A1(n8364), .A2(n27781), .Z(n27718) );
  OR3_X1 U13638 ( .A1(n17410), .A2(n988), .A3(n13081), .Z(n27976) );
  NAND2_X1 U13640 ( .A1(n29396), .A2(n19157), .ZN(n29398) );
  OAI21_X2 U13652 ( .A1(n20651), .A2(n34772), .B(n23197), .ZN(n13982) );
  XOR2_X1 U13664 ( .A1(n28876), .A2(n35633), .Z(n34773) );
  OAI22_X2 U13669 ( .A1(n8347), .A2(n29700), .B1(n8346), .B2(n8345), .ZN(
        n18042) );
  XOR2_X1 U13671 ( .A1(n35637), .A2(n7714), .Z(n35636) );
  OAI21_X2 U13673 ( .A1(n10038), .A2(n5641), .B(n10906), .ZN(n34774) );
  XOR2_X1 U13680 ( .A1(n27804), .A2(n27802), .Z(n15994) );
  XOR2_X1 U13681 ( .A1(n1466), .A2(n36384), .Z(n27804) );
  NAND2_X1 U13697 ( .A1(n31647), .A2(n36424), .ZN(n8820) );
  XOR2_X1 U13698 ( .A1(n34778), .A2(n16562), .Z(Ciphertext[187]) );
  AOI21_X2 U13726 ( .A1(n37065), .A2(n24120), .B(n5854), .ZN(n24753) );
  XOR2_X1 U13727 ( .A1(n34780), .A2(n28973), .Z(n28975) );
  XOR2_X1 U13728 ( .A1(n28972), .A2(n39220), .Z(n34780) );
  OAI21_X2 U13735 ( .A1(n34105), .A2(n33125), .B(n33705), .ZN(n24672) );
  XOR2_X1 U13740 ( .A1(n10854), .A2(n10855), .Z(n853) );
  XOR2_X1 U13741 ( .A1(n28977), .A2(n29125), .Z(n16359) );
  AOI21_X2 U13767 ( .A1(n28314), .A2(n31045), .B(n4926), .ZN(n28972) );
  XOR2_X1 U13774 ( .A1(n22405), .A2(n7432), .Z(n6474) );
  NAND2_X1 U13787 ( .A1(n34357), .A2(n39194), .ZN(n32068) );
  NOR2_X2 U13795 ( .A1(n21725), .A2(n4913), .ZN(n36281) );
  INV_X2 U13800 ( .I(n20605), .ZN(n1564) );
  AOI22_X2 U13815 ( .A1(n23038), .A2(n23540), .B1(n6301), .B2(n18746), .ZN(
        n23686) );
  XOR2_X1 U13830 ( .A1(n32776), .A2(n24052), .Z(n18683) );
  NAND2_X1 U13833 ( .A1(n34842), .A2(n27081), .ZN(n34841) );
  XOR2_X1 U13866 ( .A1(n10540), .A2(n34785), .Z(n31978) );
  XOR2_X1 U13870 ( .A1(n10538), .A2(n10539), .Z(n34785) );
  NAND2_X2 U13881 ( .A1(n36425), .A2(n37775), .ZN(n15268) );
  INV_X2 U13882 ( .I(n9218), .ZN(n259) );
  XOR2_X1 U13908 ( .A1(n6719), .A2(n5542), .Z(n34787) );
  OR2_X1 U13922 ( .A1(n7387), .A2(n38724), .Z(n34924) );
  XOR2_X1 U13924 ( .A1(n16138), .A2(n23900), .Z(n18857) );
  OAI22_X2 U13927 ( .A1(n23508), .A2(n13829), .B1(n13832), .B2(n13831), .ZN(
        n16138) );
  XOR2_X1 U13931 ( .A1(n35987), .A2(n34999), .Z(n11230) );
  XOR2_X1 U13934 ( .A1(n34789), .A2(n35112), .Z(n34999) );
  NAND2_X1 U13938 ( .A1(n14428), .A2(n21270), .ZN(n19704) );
  NAND3_X2 U13957 ( .A1(n27873), .A2(n27872), .A3(n27871), .ZN(n13601) );
  XOR2_X1 U13973 ( .A1(n22742), .A2(n8312), .Z(n22551) );
  OAI21_X1 U13979 ( .A1(n5977), .A2(n29701), .B(n20982), .ZN(n34793) );
  AOI21_X2 U13981 ( .A1(n13780), .A2(n35182), .B(n11164), .ZN(n5757) );
  OAI21_X1 U13984 ( .A1(n29758), .A2(n19348), .B(n34795), .ZN(n29759) );
  OAI21_X1 U13992 ( .A1(n34182), .A2(n29753), .B(n29756), .ZN(n34795) );
  AOI22_X2 U14052 ( .A1(n3935), .A2(n37103), .B1(n3961), .B2(n1494), .ZN(
        n34799) );
  XOR2_X1 U14077 ( .A1(n31314), .A2(n10579), .Z(n34800) );
  AOI21_X2 U14080 ( .A1(n15024), .A2(n12653), .B(n89), .ZN(n34801) );
  XOR2_X1 U14081 ( .A1(n34802), .A2(n32773), .Z(n35896) );
  XNOR2_X1 U14093 ( .A1(n37593), .A2(n26599), .ZN(n26419) );
  AOI21_X2 U14098 ( .A1(n17144), .A2(n26975), .B(n17143), .ZN(n27325) );
  NAND2_X2 U14103 ( .A1(n2946), .A2(n35499), .ZN(n36555) );
  XOR2_X1 U14118 ( .A1(n19428), .A2(n21095), .Z(n34809) );
  NAND2_X1 U14119 ( .A1(n9169), .A2(n28004), .ZN(n27893) );
  NAND2_X2 U14121 ( .A1(n35666), .A2(n3307), .ZN(n15467) );
  NAND2_X2 U14143 ( .A1(n2341), .A2(n19422), .ZN(n24663) );
  NAND2_X2 U14144 ( .A1(n20229), .A2(n20227), .ZN(n19422) );
  XOR2_X1 U14162 ( .A1(n39536), .A2(n29838), .Z(n29839) );
  NAND2_X2 U14180 ( .A1(n5439), .A2(n5438), .ZN(n5089) );
  NOR2_X1 U14182 ( .A1(n2965), .A2(n32168), .ZN(n36682) );
  XOR2_X1 U14183 ( .A1(n33868), .A2(n34814), .Z(n36063) );
  XOR2_X1 U14184 ( .A1(n3317), .A2(n34815), .Z(n34814) );
  INV_X1 U14189 ( .I(n1612), .ZN(n34815) );
  NAND2_X2 U14195 ( .A1(n14916), .A2(n23329), .ZN(n23783) );
  XOR2_X1 U14199 ( .A1(n25039), .A2(n25213), .Z(n13920) );
  NAND2_X2 U14200 ( .A1(n26056), .A2(n26089), .ZN(n25882) );
  XOR2_X1 U14223 ( .A1(n33735), .A2(n6154), .Z(n2594) );
  INV_X2 U14224 ( .I(n36579), .ZN(n33735) );
  NAND2_X2 U14238 ( .A1(n927), .A2(n26090), .ZN(n13502) );
  AOI21_X2 U14244 ( .A1(n31345), .A2(n22969), .B(n13157), .ZN(n13370) );
  XOR2_X1 U14251 ( .A1(n4269), .A2(n4271), .Z(n10071) );
  XOR2_X1 U14258 ( .A1(n8909), .A2(n34825), .Z(n3297) );
  XOR2_X1 U14261 ( .A1(n3299), .A2(n9106), .Z(n34825) );
  NAND3_X2 U14263 ( .A1(n32586), .A2(n34826), .A3(n2418), .ZN(n11752) );
  NOR2_X2 U14270 ( .A1(n12329), .A2(n37166), .ZN(n14729) );
  INV_X2 U14272 ( .I(n34828), .ZN(n14080) );
  NAND2_X2 U14280 ( .A1(n1577), .A2(n8966), .ZN(n13221) );
  XOR2_X1 U14285 ( .A1(n22529), .A2(n22594), .Z(n22771) );
  NOR2_X2 U14286 ( .A1(n6199), .A2(n33594), .ZN(n22529) );
  OAI21_X2 U14289 ( .A1(n34830), .A2(n26822), .B(n14798), .ZN(n34969) );
  OR2_X1 U14303 ( .A1(n14377), .A2(n26761), .Z(n26758) );
  AND2_X1 U14304 ( .A1(n39112), .A2(n28224), .Z(n7326) );
  INV_X2 U14308 ( .I(n26224), .ZN(n17048) );
  NAND2_X2 U14309 ( .A1(n25112), .A2(n18864), .ZN(n26224) );
  OAI21_X1 U14310 ( .A1(n24607), .A2(n12846), .B(n29285), .ZN(n9031) );
  NOR2_X1 U14313 ( .A1(n17451), .A2(n37553), .ZN(n36488) );
  NAND2_X2 U14327 ( .A1(n11631), .A2(n11630), .ZN(n24745) );
  XOR2_X1 U14333 ( .A1(n6384), .A2(n8303), .Z(n28842) );
  NAND2_X2 U14337 ( .A1(n26678), .A2(n34837), .ZN(n27436) );
  NAND3_X1 U14339 ( .A1(n26823), .A2(n20021), .A3(n37643), .ZN(n34837) );
  NAND2_X2 U14342 ( .A1(n34838), .A2(n18350), .ZN(n14808) );
  OAI21_X2 U14343 ( .A1(n17390), .A2(n27973), .B(n28156), .ZN(n34871) );
  NOR2_X2 U14348 ( .A1(n21239), .A2(n28290), .ZN(n27973) );
  NOR2_X1 U14349 ( .A1(n34841), .A2(n34840), .ZN(n10336) );
  NOR2_X1 U14352 ( .A1(n27164), .A2(n35750), .ZN(n34840) );
  NAND2_X1 U14363 ( .A1(n25849), .A2(n34350), .ZN(n25851) );
  NAND2_X2 U14368 ( .A1(n35327), .A2(n25376), .ZN(n25849) );
  INV_X2 U14371 ( .I(n3863), .ZN(n36745) );
  INV_X2 U14375 ( .I(n20646), .ZN(n22365) );
  NAND4_X2 U14377 ( .A1(n14912), .A2(n16654), .A3(n16653), .A4(n34997), .ZN(
        n20646) );
  NAND3_X1 U14382 ( .A1(n19666), .A2(n39261), .A3(n34924), .ZN(n32487) );
  XOR2_X1 U14395 ( .A1(n38269), .A2(n34848), .Z(n744) );
  INV_X1 U14398 ( .I(n19925), .ZN(n34848) );
  OAI21_X2 U14401 ( .A1(n19215), .A2(n34402), .B(n19214), .ZN(n25659) );
  XOR2_X1 U14402 ( .A1(n3090), .A2(n35350), .Z(n36617) );
  XOR2_X1 U14411 ( .A1(n16284), .A2(n34849), .Z(n17084) );
  XOR2_X1 U14412 ( .A1(n23936), .A2(n35752), .Z(n34849) );
  XOR2_X1 U14417 ( .A1(n19577), .A2(n34850), .Z(n20207) );
  XOR2_X1 U14418 ( .A1(n23793), .A2(n34851), .Z(n34850) );
  XOR2_X1 U14431 ( .A1(n33693), .A2(n34854), .Z(n8628) );
  XOR2_X1 U14434 ( .A1(n8629), .A2(n22560), .Z(n34854) );
  NAND2_X2 U14435 ( .A1(n31325), .A2(n22826), .ZN(n34959) );
  NAND3_X1 U14440 ( .A1(n33565), .A2(n35187), .A3(n30106), .ZN(n34855) );
  XOR2_X1 U14456 ( .A1(n5586), .A2(n2543), .Z(n36884) );
  NAND2_X2 U14457 ( .A1(n4682), .A2(n12952), .ZN(n22880) );
  NOR2_X2 U14507 ( .A1(n20761), .A2(n15441), .ZN(n30800) );
  NAND2_X2 U14510 ( .A1(n38666), .A2(n18673), .ZN(n34863) );
  NAND2_X2 U14514 ( .A1(n580), .A2(n1202), .ZN(n34866) );
  INV_X1 U14530 ( .I(n21735), .ZN(n34867) );
  NAND2_X1 U14531 ( .A1(n34867), .A2(n293), .ZN(n20762) );
  XOR2_X1 U14532 ( .A1(n34869), .A2(n6739), .Z(n11948) );
  XOR2_X1 U14533 ( .A1(n35711), .A2(n26172), .Z(n34869) );
  XOR2_X1 U14534 ( .A1(n22595), .A2(n22594), .Z(n11190) );
  NOR2_X2 U14535 ( .A1(n13296), .A2(n22087), .ZN(n22595) );
  AOI22_X2 U14541 ( .A1(n34870), .A2(n11128), .B1(n8008), .B2(n1417), .ZN(
        n29819) );
  NAND3_X1 U14543 ( .A1(n21949), .A2(n21945), .A3(n21784), .ZN(n35623) );
  NAND2_X1 U14569 ( .A1(n36134), .A2(n36132), .ZN(n34877) );
  XOR2_X1 U14572 ( .A1(n26297), .A2(n34024), .Z(n36257) );
  NOR2_X1 U14573 ( .A1(n36296), .A2(n19886), .ZN(n3627) );
  INV_X4 U14574 ( .I(n24557), .ZN(n19886) );
  AOI21_X2 U14578 ( .A1(n36725), .A2(n16644), .B(n808), .ZN(n24557) );
  XOR2_X1 U14580 ( .A1(n21034), .A2(n26545), .Z(n13914) );
  XOR2_X1 U14586 ( .A1(n26455), .A2(n35627), .Z(n21034) );
  XOR2_X1 U14588 ( .A1(n10668), .A2(n34878), .Z(n3976) );
  AOI21_X2 U14602 ( .A1(n29866), .A2(n31545), .B(n34882), .ZN(n29883) );
  NOR2_X1 U14604 ( .A1(n15521), .A2(n16059), .ZN(n34882) );
  OAI21_X2 U14616 ( .A1(n32233), .A2(n32232), .B(n34885), .ZN(n26448) );
  NAND3_X2 U14622 ( .A1(n3434), .A2(n38168), .A3(n32243), .ZN(n34885) );
  NAND2_X2 U14625 ( .A1(n12650), .A2(n17541), .ZN(n16054) );
  NAND2_X2 U14628 ( .A1(n34886), .A2(n10972), .ZN(n25820) );
  AND2_X1 U14630 ( .A1(n23582), .A2(n23580), .Z(n22806) );
  NAND2_X2 U14632 ( .A1(n8460), .A2(n4698), .ZN(n23582) );
  NOR2_X1 U14633 ( .A1(n5541), .A2(n9740), .ZN(n12557) );
  INV_X2 U14634 ( .I(n5518), .ZN(n5541) );
  NAND2_X1 U14640 ( .A1(n3916), .A2(n39676), .ZN(n34939) );
  XOR2_X1 U14642 ( .A1(n9221), .A2(n9219), .Z(n14306) );
  NAND2_X2 U14662 ( .A1(n3076), .A2(n24877), .ZN(n24749) );
  NAND2_X2 U14676 ( .A1(n34890), .A2(n34889), .ZN(n6847) );
  NAND2_X2 U14677 ( .A1(n34891), .A2(n8087), .ZN(n36791) );
  NAND2_X1 U14701 ( .A1(n11306), .A2(n13801), .ZN(n34897) );
  XOR2_X1 U14724 ( .A1(n10253), .A2(n34900), .Z(n36264) );
  XOR2_X1 U14725 ( .A1(n23774), .A2(n23976), .Z(n10253) );
  NAND2_X2 U14728 ( .A1(n7882), .A2(n24246), .ZN(n34906) );
  XOR2_X1 U14739 ( .A1(n25256), .A2(n25116), .Z(n34901) );
  OAI21_X2 U14748 ( .A1(n33365), .A2(n25743), .B(n38899), .ZN(n14253) );
  XOR2_X1 U14762 ( .A1(n23884), .A2(n23774), .Z(n23696) );
  NAND2_X1 U14772 ( .A1(n30066), .A2(n30078), .ZN(n3947) );
  INV_X2 U14782 ( .I(n15697), .ZN(n36731) );
  XOR2_X1 U14789 ( .A1(n35998), .A2(n19760), .Z(n8908) );
  XOR2_X1 U14796 ( .A1(n19772), .A2(n8074), .Z(n26713) );
  AOI22_X2 U14798 ( .A1(n1872), .A2(n15163), .B1(n36553), .B2(n22944), .ZN(
        n10472) );
  OAI21_X2 U14806 ( .A1(n32795), .A2(n6689), .B(n34909), .ZN(n9184) );
  NAND3_X1 U14807 ( .A1(n27737), .A2(n27346), .A3(n27345), .ZN(n34909) );
  OAI22_X2 U14812 ( .A1(n6483), .A2(n33354), .B1(n34080), .B2(n18238), .ZN(
        n24585) );
  INV_X2 U14815 ( .I(n7317), .ZN(n33871) );
  INV_X2 U14829 ( .I(n14212), .ZN(n25764) );
  XOR2_X1 U14839 ( .A1(n10195), .A2(n34912), .Z(n25631) );
  XOR2_X1 U14841 ( .A1(n25264), .A2(n25265), .Z(n34912) );
  BUF_X2 U14846 ( .I(n26625), .Z(n26219) );
  NAND2_X1 U14859 ( .A1(n30636), .A2(n32769), .ZN(n36313) );
  AND2_X1 U14861 ( .A1(n23907), .A2(n24244), .Z(n9384) );
  NOR2_X2 U14865 ( .A1(n4973), .A2(n34906), .ZN(n3793) );
  XOR2_X1 U14874 ( .A1(n25270), .A2(n9624), .Z(n20416) );
  INV_X2 U14876 ( .I(n26807), .ZN(n34913) );
  BUF_X2 U14881 ( .I(n33964), .Z(n34914) );
  XOR2_X1 U14884 ( .A1(n26517), .A2(n26602), .Z(n26257) );
  NOR2_X2 U14885 ( .A1(n6400), .A2(n6401), .ZN(n26517) );
  OAI21_X2 U14896 ( .A1(n26937), .A2(n32745), .B(n34918), .ZN(n26940) );
  NAND2_X1 U14898 ( .A1(n10896), .A2(n17198), .ZN(n18120) );
  OAI21_X2 U14908 ( .A1(n6129), .A2(n1680), .B(n5232), .ZN(n5231) );
  NOR2_X2 U14910 ( .A1(n6128), .A2(n22295), .ZN(n6129) );
  OAI21_X2 U14914 ( .A1(n21941), .A2(n4084), .B(n36519), .ZN(n36518) );
  NOR2_X2 U14916 ( .A1(n34923), .A2(n34922), .ZN(n21941) );
  NOR2_X2 U14927 ( .A1(n34926), .A2(n34925), .ZN(n17882) );
  NOR2_X2 U14932 ( .A1(n17970), .A2(n33091), .ZN(n34926) );
  AOI22_X2 U14942 ( .A1(n20593), .A2(n15523), .B1(n15522), .B2(n17763), .ZN(
        n1812) );
  XOR2_X1 U14952 ( .A1(n35741), .A2(n12871), .Z(n36717) );
  XOR2_X1 U14953 ( .A1(n22004), .A2(n22003), .Z(n22005) );
  XOR2_X1 U14957 ( .A1(n29255), .A2(n6536), .Z(n4461) );
  NAND2_X1 U14960 ( .A1(n13579), .A2(n13578), .ZN(n35483) );
  NAND3_X2 U14979 ( .A1(n26979), .A2(n11864), .A3(n12290), .ZN(n34930) );
  NOR3_X2 U14983 ( .A1(n34932), .A2(n34931), .A3(n3480), .ZN(n35399) );
  XOR2_X1 U14995 ( .A1(n22615), .A2(n8552), .Z(n20668) );
  NOR2_X2 U14996 ( .A1(n9486), .A2(n9484), .ZN(n8552) );
  XOR2_X1 U15002 ( .A1(n3454), .A2(n23429), .Z(n36500) );
  AND2_X1 U15005 ( .A1(n5337), .A2(n12952), .Z(n5834) );
  NAND2_X2 U15006 ( .A1(n6576), .A2(n5077), .ZN(n22359) );
  OAI21_X2 U15014 ( .A1(n30272), .A2(n36368), .B(n37335), .ZN(n109) );
  NOR2_X1 U15016 ( .A1(n39405), .A2(n9197), .ZN(n34934) );
  NAND2_X1 U15017 ( .A1(n33541), .A2(n35137), .ZN(n34935) );
  NOR2_X2 U15025 ( .A1(n1962), .A2(n20673), .ZN(n2559) );
  BUF_X4 U15026 ( .I(n3927), .Z(n1823) );
  NAND2_X1 U15030 ( .A1(n24460), .A2(n19466), .ZN(n34938) );
  OR2_X1 U15032 ( .A1(n29755), .A2(n29754), .Z(n29735) );
  NOR2_X2 U15034 ( .A1(n23518), .A2(n23517), .ZN(n18475) );
  AOI21_X1 U15046 ( .A1(n12230), .A2(n4239), .B(n13778), .ZN(n35979) );
  NAND2_X2 U15049 ( .A1(n25400), .A2(n36678), .ZN(n34940) );
  XOR2_X1 U15051 ( .A1(n2582), .A2(n13883), .Z(n33112) );
  XOR2_X1 U15052 ( .A1(n34332), .A2(n27828), .Z(n2582) );
  AOI22_X2 U15059 ( .A1(n937), .A2(n30306), .B1(n17411), .B2(n12077), .ZN(
        n22333) );
  XOR2_X1 U15063 ( .A1(n12551), .A2(n31355), .Z(n15844) );
  XOR2_X1 U15088 ( .A1(n27823), .A2(n34945), .Z(n754) );
  INV_X1 U15092 ( .I(n19820), .ZN(n34945) );
  OAI21_X2 U15109 ( .A1(n21170), .A2(n21169), .B(n17697), .ZN(n27823) );
  XOR2_X1 U15112 ( .A1(n23755), .A2(n23728), .Z(n24013) );
  NAND2_X2 U15116 ( .A1(n23633), .A2(n23632), .ZN(n23728) );
  INV_X2 U15143 ( .I(n36500), .ZN(n18116) );
  OAI21_X2 U15145 ( .A1(n37163), .A2(n12435), .B(n12793), .ZN(n34953) );
  XOR2_X1 U15161 ( .A1(n22370), .A2(n22372), .Z(n34955) );
  INV_X1 U15167 ( .I(n17964), .ZN(n35073) );
  INV_X2 U15172 ( .I(n34956), .ZN(n10004) );
  NOR2_X2 U15188 ( .A1(n17041), .A2(n21800), .ZN(n22622) );
  INV_X1 U15190 ( .I(n18500), .ZN(n4748) );
  NAND2_X1 U15192 ( .A1(n34957), .A2(n18500), .ZN(n26930) );
  XOR2_X1 U15193 ( .A1(n4853), .A2(n26555), .Z(n18500) );
  INV_X2 U15200 ( .I(n8966), .ZN(n1579) );
  NAND2_X2 U15209 ( .A1(n34964), .A2(n35057), .ZN(n30174) );
  NAND2_X2 U15210 ( .A1(n31065), .A2(n30196), .ZN(n34964) );
  NOR2_X1 U15219 ( .A1(n16180), .A2(n35187), .ZN(n16277) );
  XOR2_X1 U15226 ( .A1(n21085), .A2(n34966), .Z(n26885) );
  NAND2_X2 U15230 ( .A1(n15082), .A2(n15079), .ZN(n10143) );
  XOR2_X1 U15232 ( .A1(n26376), .A2(n26490), .Z(n20656) );
  OR2_X1 U15238 ( .A1(n35693), .A2(n24735), .Z(n10115) );
  NAND2_X1 U15244 ( .A1(n34217), .A2(n35003), .ZN(n34967) );
  NOR2_X1 U15245 ( .A1(n9963), .A2(n14379), .ZN(n14630) );
  NAND2_X2 U15262 ( .A1(n34972), .A2(n12345), .ZN(n13564) );
  XOR2_X1 U15264 ( .A1(n16797), .A2(n23848), .Z(n16795) );
  INV_X2 U15289 ( .I(n29535), .ZN(n32317) );
  XOR2_X1 U15300 ( .A1(n22439), .A2(n31566), .Z(n35457) );
  NOR2_X1 U15311 ( .A1(n7804), .A2(n12630), .ZN(n34979) );
  NAND2_X2 U15326 ( .A1(n13785), .A2(n31379), .ZN(n22710) );
  NAND2_X2 U15332 ( .A1(n2900), .A2(n2899), .ZN(n18305) );
  XOR2_X1 U15342 ( .A1(n25238), .A2(n25298), .Z(n25028) );
  NOR2_X2 U15350 ( .A1(n36110), .A2(n33629), .ZN(n36109) );
  OAI21_X2 U15354 ( .A1(n35028), .A2(n1489), .B(n37955), .ZN(n34982) );
  INV_X4 U15355 ( .I(n12168), .ZN(n12237) );
  NOR2_X2 U15358 ( .A1(n11885), .A2(n15605), .ZN(n34983) );
  NOR2_X2 U15364 ( .A1(n12497), .A2(n12498), .ZN(n34984) );
  NAND3_X1 U15366 ( .A1(n1174), .A2(n31569), .A3(n29927), .ZN(n29916) );
  OAI22_X2 U15368 ( .A1(n34985), .A2(n8587), .B1(n37955), .B2(n15371), .ZN(
        n17795) );
  NOR2_X2 U15381 ( .A1(n9805), .A2(n7624), .ZN(n24819) );
  AOI21_X2 U15383 ( .A1(n37144), .A2(n1475), .B(n34990), .ZN(n34989) );
  XOR2_X1 U15389 ( .A1(n4315), .A2(n34993), .Z(n4392) );
  XOR2_X1 U15393 ( .A1(n4313), .A2(n29129), .Z(n34993) );
  AND2_X1 U15395 ( .A1(n28659), .A2(n8366), .Z(n6043) );
  NAND2_X2 U15409 ( .A1(n26075), .A2(n7660), .ZN(n26077) );
  NOR2_X2 U15412 ( .A1(n7874), .A2(n7877), .ZN(n7660) );
  NAND2_X1 U15418 ( .A1(n11497), .A2(n32419), .ZN(n11495) );
  BUF_X2 U15425 ( .I(n8972), .Z(n33083) );
  NOR2_X2 U15431 ( .A1(n35470), .A2(n789), .ZN(n5323) );
  OAI22_X2 U15440 ( .A1(n3359), .A2(n20456), .B1(n30644), .B2(n3356), .ZN(
        n35646) );
  XOR2_X1 U15447 ( .A1(n18557), .A2(n18556), .Z(n21150) );
  NAND2_X2 U15449 ( .A1(n6078), .A2(n2451), .ZN(n6077) );
  NAND3_X1 U15452 ( .A1(n21844), .A2(n6198), .A3(n18219), .ZN(n34997) );
  XOR2_X1 U15456 ( .A1(n34999), .A2(n11967), .Z(n34998) );
  NAND2_X1 U15468 ( .A1(n31799), .A2(n1435), .ZN(n3844) );
  NAND3_X2 U15482 ( .A1(n9204), .A2(n20792), .A3(n9203), .ZN(n4353) );
  NAND2_X2 U15487 ( .A1(n36094), .A2(n3813), .ZN(n21068) );
  AOI21_X2 U15498 ( .A1(n29150), .A2(n4858), .B(n29899), .ZN(n19539) );
  NAND3_X1 U15499 ( .A1(n34007), .A2(n32146), .A3(n974), .ZN(n4857) );
  INV_X2 U15503 ( .I(n36496), .ZN(n1472) );
  XOR2_X1 U15512 ( .A1(n18796), .A2(n33131), .Z(n26795) );
  NOR2_X2 U15518 ( .A1(n3010), .A2(n3011), .ZN(n36967) );
  XOR2_X1 U15533 ( .A1(n27592), .A2(n35334), .Z(n27593) );
  NOR2_X2 U15538 ( .A1(n35791), .A2(n35792), .ZN(n35006) );
  XOR2_X1 U15560 ( .A1(n5965), .A2(n35010), .Z(n302) );
  XOR2_X1 U15562 ( .A1(n9490), .A2(n33388), .Z(n35010) );
  AND2_X1 U15563 ( .A1(n39564), .A2(n5960), .Z(n10565) );
  AOI21_X2 U15577 ( .A1(n34129), .A2(n23480), .B(n35013), .ZN(n35012) );
  NAND2_X2 U15588 ( .A1(n1045), .A2(n16104), .ZN(n35016) );
  NAND2_X1 U15590 ( .A1(n35655), .A2(n20530), .ZN(n36598) );
  XOR2_X1 U15598 ( .A1(n6526), .A2(n6525), .Z(n35017) );
  NAND2_X1 U15602 ( .A1(n1400), .A2(n482), .ZN(n28823) );
  NAND2_X2 U15606 ( .A1(n19630), .A2(n33344), .ZN(n16749) );
  INV_X2 U15613 ( .I(n35021), .ZN(n20212) );
  XOR2_X1 U15614 ( .A1(n20210), .A2(n26009), .Z(n35021) );
  INV_X2 U15625 ( .I(n33707), .ZN(n35023) );
  OR2_X1 U15627 ( .A1(n28598), .A2(n35023), .Z(n28601) );
  NAND2_X2 U15630 ( .A1(n35025), .A2(n35336), .ZN(n15165) );
  NOR2_X2 U15631 ( .A1(n15169), .A2(n15168), .ZN(n35025) );
  OR2_X1 U15633 ( .A1(n10220), .A2(n35462), .Z(n36872) );
  XNOR2_X1 U15638 ( .A1(n4348), .A2(n19758), .ZN(n36494) );
  AOI22_X2 U15640 ( .A1(n35026), .A2(n14373), .B1(n19403), .B2(n19768), .ZN(
        n32292) );
  NAND2_X2 U15646 ( .A1(n19768), .A2(n19262), .ZN(n21813) );
  XOR2_X1 U15650 ( .A1(n10185), .A2(n10183), .Z(n35027) );
  INV_X2 U15654 ( .I(n28516), .ZN(n9674) );
  OAI21_X2 U15657 ( .A1(n24391), .A2(n9931), .B(n9840), .ZN(n24761) );
  XOR2_X1 U15663 ( .A1(n22572), .A2(n22595), .Z(n22717) );
  NOR2_X2 U15665 ( .A1(n21829), .A2(n21828), .ZN(n22572) );
  XOR2_X1 U15670 ( .A1(n37957), .A2(n29934), .Z(n23744) );
  OAI21_X2 U15689 ( .A1(n34041), .A2(n28691), .B(n33353), .ZN(n2566) );
  XOR2_X1 U15690 ( .A1(n28845), .A2(n28957), .Z(n13630) );
  XOR2_X1 U15697 ( .A1(n16776), .A2(n9977), .Z(n16775) );
  XOR2_X1 U15700 ( .A1(n8566), .A2(n34053), .Z(n24009) );
  XOR2_X1 U15701 ( .A1(n23762), .A2(n30321), .Z(n8566) );
  XOR2_X1 U15706 ( .A1(n35029), .A2(n19527), .Z(Ciphertext[125]) );
  NAND2_X1 U15716 ( .A1(n15174), .A2(n29542), .ZN(n7436) );
  NAND2_X1 U15717 ( .A1(n1497), .A2(n15996), .ZN(n26670) );
  NAND2_X1 U15720 ( .A1(n32558), .A2(n14229), .ZN(n25651) );
  OAI21_X2 U15740 ( .A1(n35031), .A2(n12987), .B(n7282), .ZN(n7632) );
  NAND2_X1 U15743 ( .A1(n12986), .A2(n1002), .ZN(n35031) );
  NAND2_X2 U15744 ( .A1(n36664), .A2(n36891), .ZN(n24416) );
  INV_X2 U15752 ( .I(n35032), .ZN(n30494) );
  XOR2_X1 U15753 ( .A1(n11117), .A2(n11114), .Z(n35032) );
  XOR2_X1 U15755 ( .A1(n35033), .A2(n27815), .Z(n30806) );
  OAI21_X2 U15756 ( .A1(n29899), .A2(n29898), .B(n29949), .ZN(n36843) );
  OAI22_X2 U15761 ( .A1(n9078), .A2(n22493), .B1(n8692), .B2(n6303), .ZN(
        n32089) );
  NAND2_X2 U15769 ( .A1(n36301), .A2(n24517), .ZN(n25215) );
  BUF_X4 U15778 ( .I(n28036), .Z(n36979) );
  OAI22_X2 U15788 ( .A1(n35733), .A2(n27996), .B1(n28002), .B2(n28001), .ZN(
        n3900) );
  NAND2_X1 U15790 ( .A1(n15232), .A2(n35034), .ZN(n4730) );
  NAND3_X1 U15794 ( .A1(n32317), .A2(n29534), .A3(n18384), .ZN(n35034) );
  OR2_X1 U15795 ( .A1(n29927), .A2(n29929), .Z(n7457) );
  AOI21_X2 U15796 ( .A1(n8666), .A2(n14600), .B(n31356), .ZN(n29927) );
  XOR2_X1 U15802 ( .A1(n27605), .A2(n35035), .Z(n10256) );
  XOR2_X1 U15804 ( .A1(n557), .A2(n32160), .Z(n35035) );
  NAND2_X1 U15820 ( .A1(n27304), .A2(n31955), .ZN(n35749) );
  BUF_X2 U15825 ( .I(n23532), .Z(n35039) );
  BUF_X2 U15828 ( .I(n1145), .Z(n35040) );
  NOR3_X1 U15830 ( .A1(n916), .A2(n14423), .A3(n19873), .ZN(n12377) );
  OAI21_X2 U15841 ( .A1(n7691), .A2(n15512), .B(n36112), .ZN(n16968) );
  NAND2_X2 U15855 ( .A1(n21804), .A2(n36735), .ZN(n35042) );
  XOR2_X1 U15874 ( .A1(n7786), .A2(n7785), .Z(n18574) );
  NAND2_X1 U15877 ( .A1(n36003), .A2(n232), .ZN(n35670) );
  NAND2_X2 U15879 ( .A1(n8332), .A2(n8331), .ZN(n35051) );
  OR2_X1 U15883 ( .A1(n10803), .A2(n29220), .Z(n12978) );
  NOR2_X2 U15888 ( .A1(n25361), .A2(n10686), .ZN(n25248) );
  XOR2_X1 U15893 ( .A1(n33372), .A2(n31720), .Z(n17597) );
  XOR2_X1 U15901 ( .A1(n7530), .A2(n17195), .Z(n17987) );
  OAI21_X2 U15906 ( .A1(n12815), .A2(n12813), .B(n12812), .ZN(n17195) );
  OAI21_X2 U15907 ( .A1(n19409), .A2(n28746), .B(n19408), .ZN(n35222) );
  NAND2_X2 U15908 ( .A1(n34244), .A2(n2147), .ZN(n18202) );
  OAI21_X2 U15920 ( .A1(n35863), .A2(n35045), .B(n1316), .ZN(n2796) );
  NOR2_X1 U15921 ( .A1(n9975), .A2(n20590), .ZN(n35045) );
  AOI22_X2 U15927 ( .A1(n35046), .A2(n35944), .B1(n9882), .B2(n1934), .ZN(
        n35821) );
  INV_X2 U15928 ( .I(n35047), .ZN(n22723) );
  XOR2_X1 U15929 ( .A1(n22599), .A2(n19819), .Z(n35047) );
  INV_X2 U15943 ( .I(n35137), .ZN(n35049) );
  XOR2_X1 U15945 ( .A1(n26598), .A2(n26325), .Z(n35656) );
  XOR2_X1 U15949 ( .A1(n27690), .A2(n33866), .Z(n33498) );
  AND2_X1 U15952 ( .A1(n34717), .A2(n6445), .Z(n3515) );
  INV_X2 U15972 ( .I(n22263), .ZN(n35526) );
  NAND3_X1 U15975 ( .A1(n35055), .A2(n1595), .A3(n35054), .ZN(n20250) );
  NAND2_X1 U15980 ( .A1(n5985), .A2(n1276), .ZN(n35054) );
  INV_X1 U15984 ( .I(n20068), .ZN(n35055) );
  NAND2_X2 U15994 ( .A1(n19630), .A2(n24635), .ZN(n11711) );
  NAND2_X2 U15997 ( .A1(n35056), .A2(n11577), .ZN(n11710) );
  AND2_X1 U16000 ( .A1(n28199), .A2(n18061), .Z(n35733) );
  NOR3_X2 U16001 ( .A1(n26014), .A2(n26013), .A3(n33474), .ZN(n20852) );
  XOR2_X1 U16012 ( .A1(n11899), .A2(n25311), .Z(n6233) );
  XOR2_X1 U16013 ( .A1(n25186), .A2(n19156), .Z(n25311) );
  NOR2_X1 U16029 ( .A1(n27894), .A2(n36253), .ZN(n35061) );
  AOI22_X2 U16031 ( .A1(n14398), .A2(n36663), .B1(n36076), .B2(n14489), .ZN(
        n6809) );
  NAND2_X2 U16035 ( .A1(n27180), .A2(n33773), .ZN(n31459) );
  OAI21_X2 U16036 ( .A1(n10699), .A2(n8569), .B(n10697), .ZN(n23550) );
  NOR2_X2 U16040 ( .A1(n24647), .A2(n18569), .ZN(n24935) );
  XOR2_X1 U16044 ( .A1(n35064), .A2(n18432), .Z(Ciphertext[127]) );
  OAI22_X1 U16045 ( .A1(n29914), .A2(n29931), .B1(n29913), .B2(n19097), .ZN(
        n35064) );
  XOR2_X1 U16058 ( .A1(n21087), .A2(n27844), .Z(n20140) );
  XOR2_X1 U16061 ( .A1(n27460), .A2(n1214), .Z(n27844) );
  OAI22_X2 U16064 ( .A1(n2300), .A2(n21845), .B1(n21349), .B2(n21667), .ZN(
        n37041) );
  NAND2_X2 U16066 ( .A1(n19517), .A2(n31222), .ZN(n2300) );
  XOR2_X1 U16083 ( .A1(n9028), .A2(n6475), .Z(n23080) );
  XOR2_X1 U16085 ( .A1(n6474), .A2(n6473), .Z(n6475) );
  OR2_X1 U16090 ( .A1(n9649), .A2(n10679), .Z(n29954) );
  NAND2_X2 U16102 ( .A1(n1688), .A2(n22222), .ZN(n22224) );
  NAND2_X2 U16103 ( .A1(n37105), .A2(n3510), .ZN(n25052) );
  XOR2_X1 U16106 ( .A1(n16254), .A2(n13254), .Z(n35070) );
  INV_X2 U16108 ( .I(n35072), .ZN(n31278) );
  XOR2_X1 U16109 ( .A1(n3167), .A2(n3166), .Z(n35072) );
  INV_X1 U16112 ( .I(n114), .ZN(n15337) );
  NAND2_X1 U16118 ( .A1(n35073), .A2(n114), .ZN(n15761) );
  XOR2_X1 U16119 ( .A1(Plaintext[90]), .A2(Key[90]), .Z(n114) );
  NOR2_X1 U16122 ( .A1(n32971), .A2(n34458), .ZN(n35281) );
  NAND2_X1 U16124 ( .A1(n38973), .A2(n35281), .ZN(n35280) );
  NAND4_X2 U16140 ( .A1(n18563), .A2(n10969), .A3(n17688), .A4(n18564), .ZN(
        n20987) );
  XOR2_X1 U16150 ( .A1(n5866), .A2(n23396), .Z(n35076) );
  INV_X2 U16151 ( .I(n35077), .ZN(n4048) );
  XOR2_X1 U16154 ( .A1(n35079), .A2(n35078), .Z(n32856) );
  XOR2_X1 U16156 ( .A1(n11192), .A2(n22606), .Z(n35079) );
  OAI22_X1 U16166 ( .A1(n36976), .A2(n36977), .B1(n10428), .B2(n14421), .ZN(
        n29217) );
  INV_X2 U16167 ( .I(n35080), .ZN(n783) );
  NAND2_X2 U16173 ( .A1(n31959), .A2(n18311), .ZN(n27399) );
  INV_X1 U16175 ( .I(n4761), .ZN(n35394) );
  XOR2_X1 U16178 ( .A1(n22604), .A2(n1161), .Z(n35081) );
  NOR2_X2 U16179 ( .A1(n35082), .A2(n12545), .ZN(n29253) );
  XOR2_X1 U16192 ( .A1(n8533), .A2(n8530), .Z(n31976) );
  XOR2_X1 U16193 ( .A1(n35084), .A2(n35511), .Z(n35842) );
  XOR2_X1 U16194 ( .A1(n25224), .A2(n16674), .Z(n35084) );
  XOR2_X1 U16195 ( .A1(n4461), .A2(n35085), .Z(n33023) );
  XOR2_X1 U16196 ( .A1(n14171), .A2(n19126), .Z(n35085) );
  NAND2_X2 U16198 ( .A1(n601), .A2(n27507), .ZN(n36639) );
  NAND2_X1 U16207 ( .A1(n9682), .A2(n17645), .ZN(n13756) );
  NOR2_X1 U16220 ( .A1(n36304), .A2(n9954), .ZN(n6005) );
  OR2_X2 U16224 ( .A1(n20830), .A2(n20726), .Z(n13261) );
  XOR2_X1 U16227 ( .A1(n1859), .A2(n14218), .Z(n35908) );
  XOR2_X1 U16234 ( .A1(n35087), .A2(n34022), .Z(n13352) );
  XOR2_X1 U16236 ( .A1(n13354), .A2(n22653), .Z(n35087) );
  OR2_X1 U16247 ( .A1(n24558), .A2(n35088), .Z(n10774) );
  XOR2_X1 U16249 ( .A1(n25032), .A2(n5026), .Z(n3187) );
  XOR2_X1 U16250 ( .A1(n25197), .A2(n25149), .Z(n5026) );
  AOI22_X2 U16254 ( .A1(n4713), .A2(n1145), .B1(n4682), .B2(n15045), .ZN(
        n22969) );
  NOR2_X2 U16261 ( .A1(n7429), .A2(n5424), .ZN(n20621) );
  NAND2_X2 U16266 ( .A1(n35092), .A2(n18702), .ZN(n6263) );
  NAND2_X2 U16268 ( .A1(n35093), .A2(n11893), .ZN(n33100) );
  OAI21_X2 U16274 ( .A1(n28126), .A2(n27482), .B(n11895), .ZN(n35093) );
  XOR2_X1 U16277 ( .A1(n3887), .A2(n3890), .Z(n21159) );
  AOI22_X1 U16288 ( .A1(n5821), .A2(n9422), .B1(n33168), .B2(n1339), .ZN(n7105) );
  NOR2_X2 U16289 ( .A1(n37041), .A2(n8073), .ZN(n33168) );
  NAND2_X2 U16292 ( .A1(n30174), .A2(n10101), .ZN(n20342) );
  NAND2_X2 U16295 ( .A1(n35096), .A2(n4799), .ZN(n30093) );
  XOR2_X1 U16303 ( .A1(n29819), .A2(n28817), .Z(n29245) );
  NOR2_X2 U16316 ( .A1(n22128), .A2(n4424), .ZN(n18566) );
  XOR2_X1 U16332 ( .A1(n12575), .A2(n35097), .Z(n4866) );
  XOR2_X1 U16334 ( .A1(n12574), .A2(n32306), .Z(n35097) );
  AOI22_X2 U16345 ( .A1(n31781), .A2(n42), .B1(n8369), .B2(n1444), .ZN(n8366)
         );
  XOR2_X1 U16346 ( .A1(n23725), .A2(n1993), .Z(n33559) );
  AOI21_X1 U16351 ( .A1(n38155), .A2(n6287), .B(n13379), .ZN(n10272) );
  OAI22_X1 U16372 ( .A1(n29735), .A2(n29728), .B1(n38143), .B2(n29750), .ZN(
        n29729) );
  NOR2_X2 U16388 ( .A1(n36071), .A2(n18786), .ZN(n2626) );
  NOR2_X1 U16414 ( .A1(n2035), .A2(n39296), .ZN(n27486) );
  XOR2_X1 U16419 ( .A1(n36867), .A2(n22644), .Z(n16254) );
  OAI21_X2 U16428 ( .A1(n2060), .A2(n28356), .B(n11129), .ZN(n28817) );
  BUF_X4 U16429 ( .I(n26177), .Z(n26700) );
  AOI21_X2 U16430 ( .A1(n1514), .A2(n9175), .B(n35102), .ZN(n3519) );
  INV_X2 U16431 ( .I(n26114), .ZN(n35102) );
  XOR2_X1 U16441 ( .A1(n27730), .A2(n27525), .Z(n12507) );
  XOR2_X1 U16443 ( .A1(n29128), .A2(n29126), .Z(n21077) );
  XOR2_X1 U16451 ( .A1(n26523), .A2(n2195), .Z(n35105) );
  NAND2_X1 U16455 ( .A1(n14739), .A2(n37088), .ZN(n14742) );
  NAND3_X2 U16460 ( .A1(n23069), .A2(n6000), .A3(n11366), .ZN(n31594) );
  XOR2_X1 U16466 ( .A1(n26565), .A2(n29476), .Z(n26198) );
  NAND2_X2 U16468 ( .A1(n33423), .A2(n21198), .ZN(n26565) );
  NAND2_X2 U16472 ( .A1(n20168), .A2(n16581), .ZN(n25242) );
  NAND2_X2 U16474 ( .A1(n24751), .A2(n24750), .ZN(n20168) );
  NAND2_X2 U16477 ( .A1(n37099), .A2(n29491), .ZN(n20209) );
  NAND2_X2 U16480 ( .A1(n35108), .A2(n24199), .ZN(n24719) );
  NAND3_X2 U16481 ( .A1(n37065), .A2(n32491), .A3(n32492), .ZN(n35108) );
  XOR2_X1 U16490 ( .A1(n19014), .A2(n14610), .Z(n31849) );
  INV_X4 U16491 ( .I(n32885), .ZN(n1323) );
  NAND2_X2 U16492 ( .A1(n5063), .A2(n5768), .ZN(n24704) );
  XOR2_X1 U16496 ( .A1(n28840), .A2(n29146), .Z(n36545) );
  OR2_X1 U16501 ( .A1(n9520), .A2(n23907), .Z(n10342) );
  OAI21_X2 U16511 ( .A1(n33725), .A2(n879), .B(n37623), .ZN(n6264) );
  BUF_X4 U16529 ( .I(n15933), .Z(n12771) );
  INV_X1 U16533 ( .I(n25851), .ZN(n36896) );
  XNOR2_X1 U16534 ( .A1(n9757), .A2(n15401), .ZN(n140) );
  XOR2_X1 U16540 ( .A1(n23777), .A2(n34054), .Z(n32610) );
  BUF_X2 U16545 ( .I(n6893), .Z(n35112) );
  NAND3_X2 U16547 ( .A1(n30584), .A2(n7227), .A3(n35113), .ZN(n32404) );
  INV_X2 U16560 ( .I(n1218), .ZN(n35114) );
  NOR2_X2 U16570 ( .A1(n22100), .A2(n9736), .ZN(n22176) );
  NAND3_X1 U16584 ( .A1(n1477), .A2(n997), .A3(n8537), .ZN(n27158) );
  XOR2_X1 U16605 ( .A1(n25249), .A2(n25299), .Z(n11519) );
  AND2_X1 U16606 ( .A1(n24425), .A2(n14371), .Z(n5254) );
  NAND2_X2 U16612 ( .A1(n14371), .A2(n10073), .ZN(n24425) );
  XOR2_X1 U16621 ( .A1(n34092), .A2(n35120), .Z(n36104) );
  XOR2_X1 U16634 ( .A1(n25156), .A2(n5829), .Z(n35120) );
  INV_X4 U16635 ( .I(n18028), .ZN(n12927) );
  OAI21_X2 U16636 ( .A1(n17098), .A2(n17099), .B(n35121), .ZN(n11020) );
  AOI22_X2 U16638 ( .A1(n14830), .A2(n26978), .B1(n14831), .B2(n33301), .ZN(
        n35121) );
  NAND2_X1 U16644 ( .A1(n8042), .A2(n10008), .ZN(n35122) );
  NOR2_X1 U16653 ( .A1(n978), .A2(n33100), .ZN(n30917) );
  NOR3_X1 U16655 ( .A1(n35979), .A2(n12377), .A3(n22388), .ZN(n36349) );
  AOI21_X2 U16657 ( .A1(n2028), .A2(n35822), .B(n35194), .ZN(n35193) );
  NAND2_X2 U16660 ( .A1(n12669), .A2(n8228), .ZN(n33437) );
  NOR2_X2 U16673 ( .A1(n21318), .A2(n19748), .ZN(n35124) );
  XOR2_X1 U16695 ( .A1(n36497), .A2(n2119), .Z(n36231) );
  NAND2_X1 U16717 ( .A1(n9211), .A2(n9213), .ZN(n36322) );
  AOI22_X2 U16724 ( .A1(n22950), .A2(n39752), .B1(n22951), .B2(n23020), .ZN(
        n22952) );
  NOR2_X1 U16729 ( .A1(n21609), .A2(n21610), .ZN(n36297) );
  NOR2_X2 U16730 ( .A1(n31437), .A2(n34031), .ZN(n35686) );
  XOR2_X1 U16734 ( .A1(n13917), .A2(n25211), .Z(n25039) );
  AOI21_X1 U16740 ( .A1(n22366), .A2(n22227), .B(n20623), .ZN(n21104) );
  NAND2_X2 U16748 ( .A1(n20643), .A2(n20646), .ZN(n22227) );
  INV_X2 U16789 ( .I(n38669), .ZN(n36777) );
  XOR2_X1 U16792 ( .A1(n22462), .A2(n6325), .Z(n7931) );
  XOR2_X1 U16793 ( .A1(n22582), .A2(n18778), .Z(n22462) );
  INV_X1 U16800 ( .I(n479), .ZN(n27433) );
  NOR3_X1 U16803 ( .A1(n29433), .A2(n14414), .A3(n18502), .ZN(n29436) );
  NAND2_X2 U16809 ( .A1(n28569), .A2(n33995), .ZN(n28448) );
  INV_X2 U16813 ( .I(n22586), .ZN(n1668) );
  NOR2_X1 U16835 ( .A1(n1313), .A2(n8942), .ZN(n10867) );
  INV_X2 U16841 ( .I(n5732), .ZN(n8942) );
  OR2_X1 U16843 ( .A1(n21445), .A2(n21669), .Z(n31292) );
  BUF_X4 U16858 ( .I(n19979), .Z(n36082) );
  NAND3_X1 U16868 ( .A1(n30071), .A2(n30076), .A3(n4377), .ZN(n30073) );
  OAI22_X1 U16874 ( .A1(n22840), .A2(n13042), .B1(n23106), .B2(n23104), .ZN(
        n22841) );
  XOR2_X1 U16882 ( .A1(n22391), .A2(n22656), .Z(n22457) );
  XOR2_X1 U16887 ( .A1(n18300), .A2(n8951), .Z(n15648) );
  XOR2_X1 U16892 ( .A1(n17775), .A2(n35139), .Z(n33676) );
  XOR2_X1 U16894 ( .A1(n9979), .A2(n35140), .Z(n35139) );
  NAND2_X1 U16902 ( .A1(n29547), .A2(n35141), .ZN(n21069) );
  INV_X2 U16907 ( .I(n19097), .ZN(n29932) );
  XOR2_X1 U16908 ( .A1(n11927), .A2(n11925), .Z(n15738) );
  INV_X2 U16917 ( .I(n35143), .ZN(n30853) );
  XOR2_X1 U16921 ( .A1(n29077), .A2(n20622), .Z(n29381) );
  NAND3_X2 U16929 ( .A1(n35144), .A2(n5294), .A3(n5295), .ZN(n36894) );
  NAND2_X1 U16940 ( .A1(n14127), .A2(n3693), .ZN(n35547) );
  OAI21_X2 U16942 ( .A1(n9292), .A2(n9293), .B(n25630), .ZN(n35145) );
  AOI21_X2 U16946 ( .A1(n35146), .A2(n5509), .B(n14642), .ZN(n5705) );
  NAND2_X2 U16953 ( .A1(n584), .A2(n33860), .ZN(n16281) );
  OAI21_X2 U16958 ( .A1(n17077), .A2(n28311), .B(n15211), .ZN(n8911) );
  XOR2_X1 U16970 ( .A1(n18942), .A2(n35147), .Z(n35868) );
  XOR2_X1 U16971 ( .A1(n35760), .A2(n35148), .Z(n35147) );
  INV_X2 U16977 ( .I(n35149), .ZN(n21137) );
  XNOR2_X1 U16978 ( .A1(n18578), .A2(n18580), .ZN(n35149) );
  AOI22_X2 U16981 ( .A1(n19146), .A2(n23321), .B1(n16047), .B2(n961), .ZN(
        n18485) );
  XOR2_X1 U16983 ( .A1(n7766), .A2(n28989), .Z(n20819) );
  XOR2_X1 U16984 ( .A1(n12741), .A2(n8939), .Z(n28989) );
  AND2_X1 U16986 ( .A1(n19667), .A2(n34370), .Z(n31913) );
  AOI21_X1 U16993 ( .A1(n33416), .A2(n29735), .B(n29733), .ZN(n29736) );
  NAND2_X2 U17003 ( .A1(n29486), .A2(n14417), .ZN(n29444) );
  NAND2_X2 U17019 ( .A1(n11952), .A2(n35155), .ZN(n18289) );
  AOI21_X1 U17031 ( .A1(n37050), .A2(n955), .B(n32105), .ZN(n35156) );
  XNOR2_X1 U17036 ( .A1(n29073), .A2(n18430), .ZN(n9994) );
  XNOR2_X1 U17041 ( .A1(n15595), .A2(n26397), .ZN(n36468) );
  NAND2_X1 U17045 ( .A1(n25883), .A2(n8006), .ZN(n35159) );
  XOR2_X1 U17059 ( .A1(n208), .A2(n23777), .Z(n5510) );
  BUF_X2 U17061 ( .I(n25427), .Z(n35160) );
  XOR2_X1 U17063 ( .A1(n27617), .A2(n27594), .Z(n35708) );
  NAND3_X2 U17065 ( .A1(n26846), .A2(n26844), .A3(n26845), .ZN(n27594) );
  INV_X2 U17066 ( .I(n35161), .ZN(n8293) );
  XOR2_X1 U17072 ( .A1(n35162), .A2(n35389), .Z(n32049) );
  XOR2_X1 U17073 ( .A1(n17349), .A2(n38174), .Z(n35162) );
  XOR2_X1 U17076 ( .A1(n3550), .A2(n3548), .Z(n9393) );
  XOR2_X1 U17080 ( .A1(n21030), .A2(n5116), .Z(n35163) );
  XOR2_X1 U17083 ( .A1(n7582), .A2(n34052), .Z(n32432) );
  OAI21_X2 U17105 ( .A1(n39829), .A2(n35165), .B(n28789), .ZN(n30131) );
  NOR2_X1 U17112 ( .A1(n28788), .A2(n38196), .ZN(n35165) );
  XOR2_X1 U17118 ( .A1(n8958), .A2(n35421), .Z(n9470) );
  XOR2_X1 U17121 ( .A1(n29086), .A2(n35168), .Z(n31867) );
  XOR2_X1 U17123 ( .A1(n8939), .A2(n35169), .Z(n35168) );
  INV_X1 U17125 ( .I(n29476), .ZN(n35169) );
  XOR2_X1 U17126 ( .A1(n36869), .A2(n6328), .Z(n36932) );
  AOI21_X1 U17131 ( .A1(n12189), .A2(n6648), .B(n35287), .ZN(n13721) );
  OAI22_X2 U17144 ( .A1(n17475), .A2(n39537), .B1(n20154), .B2(n35170), .ZN(
        n17474) );
  XOR2_X1 U17147 ( .A1(n25210), .A2(n25174), .Z(n5315) );
  AOI21_X2 U17157 ( .A1(n9997), .A2(n6337), .B(n24600), .ZN(n24128) );
  NOR3_X2 U17158 ( .A1(n11710), .A2(n3120), .A3(n15332), .ZN(n3124) );
  INV_X4 U17159 ( .I(n29862), .ZN(n29956) );
  OR2_X1 U17164 ( .A1(n35217), .A2(n37060), .Z(n19088) );
  INV_X2 U17165 ( .I(n27571), .ZN(n35417) );
  INV_X2 U17168 ( .I(n28961), .ZN(n29761) );
  NOR2_X2 U17173 ( .A1(n4322), .A2(n36546), .ZN(n25743) );
  NAND2_X2 U17176 ( .A1(n30260), .A2(n30257), .ZN(n30250) );
  OR2_X2 U17181 ( .A1(n11428), .A2(n39827), .Z(n11125) );
  INV_X2 U17188 ( .I(n482), .ZN(n30165) );
  NAND2_X1 U17189 ( .A1(n24235), .A2(n30311), .ZN(n8160) );
  NAND2_X2 U17201 ( .A1(n18873), .A2(n9105), .ZN(n20964) );
  NAND2_X2 U17204 ( .A1(n36859), .A2(n33316), .ZN(n13010) );
  NOR2_X1 U17207 ( .A1(n31587), .A2(n12931), .ZN(n35171) );
  INV_X1 U17210 ( .I(n25699), .ZN(n1110) );
  NOR2_X1 U17233 ( .A1(n38164), .A2(n8287), .ZN(n20922) );
  OAI22_X1 U17236 ( .A1(n981), .A2(n1207), .B1(n5469), .B2(n28290), .ZN(n30872) );
  AOI22_X1 U17242 ( .A1(n29605), .A2(n29604), .B1(n29625), .B2(n29611), .ZN(
        n30657) );
  NAND2_X1 U17245 ( .A1(n18306), .A2(n36382), .ZN(n29625) );
  NAND3_X1 U17247 ( .A1(n76), .A2(n17532), .A3(n2877), .ZN(n2666) );
  NOR2_X2 U17252 ( .A1(n36029), .A2(n10393), .ZN(n35173) );
  OR2_X1 U17263 ( .A1(n13442), .A2(n17262), .Z(n19173) );
  CLKBUF_X12 U17283 ( .I(n20512), .Z(n31022) );
  NAND2_X1 U17285 ( .A1(n31022), .A2(n6640), .ZN(n2050) );
  NAND2_X1 U17291 ( .A1(n9141), .A2(n28717), .ZN(n11009) );
  INV_X1 U17295 ( .I(n20454), .ZN(n20659) );
  NOR2_X1 U17301 ( .A1(n28490), .A2(n18960), .ZN(n12544) );
  NAND3_X1 U17304 ( .A1(n28490), .A2(n18960), .A3(n4950), .ZN(n28452) );
  NOR2_X1 U17307 ( .A1(n32781), .A2(n18626), .ZN(n18625) );
  AOI22_X1 U17320 ( .A1(n29688), .A2(n5067), .B1(n29685), .B2(n29686), .ZN(
        n31914) );
  INV_X1 U17321 ( .I(n18837), .ZN(n36767) );
  INV_X2 U17323 ( .I(n23307), .ZN(n22493) );
  NAND3_X1 U17324 ( .A1(n29392), .A2(n29393), .A3(n29391), .ZN(n35676) );
  NAND2_X1 U17338 ( .A1(n29232), .A2(n35185), .ZN(n36232) );
  NOR2_X1 U17339 ( .A1(n5955), .A2(n7834), .ZN(n5954) );
  OAI21_X1 U17351 ( .A1(n10763), .A2(n13752), .B(n11453), .ZN(n35811) );
  OR2_X1 U17355 ( .A1(n28585), .A2(n28584), .Z(n35179) );
  NAND2_X1 U17364 ( .A1(n30035), .A2(n8039), .ZN(n18783) );
  OAI21_X1 U17367 ( .A1(n20102), .A2(n37021), .B(n30059), .ZN(n36268) );
  AOI22_X1 U17381 ( .A1(n20922), .A2(n17192), .B1(n30129), .B2(n38164), .ZN(
        n20921) );
  NOR2_X1 U17392 ( .A1(n36964), .A2(n10708), .ZN(n24036) );
  AOI21_X2 U17393 ( .A1(n10711), .A2(n9011), .B(n36965), .ZN(n36964) );
  BUF_X2 U17397 ( .I(n26651), .Z(n4138) );
  NAND2_X1 U17400 ( .A1(n33203), .A2(n30986), .ZN(n31764) );
  INV_X2 U17401 ( .I(n29699), .ZN(n1182) );
  NAND2_X1 U17405 ( .A1(n38163), .A2(n20274), .ZN(n29007) );
  NAND2_X1 U17407 ( .A1(n1193), .A2(n28311), .ZN(n15211) );
  NOR2_X1 U17417 ( .A1(n28749), .A2(n28746), .ZN(n33106) );
  NAND2_X1 U17418 ( .A1(n4024), .A2(n28746), .ZN(n4023) );
  NAND2_X1 U17438 ( .A1(n9200), .A2(n38227), .ZN(n7797) );
  NOR2_X1 U17446 ( .A1(n28823), .A2(n30160), .ZN(n35183) );
  AND2_X1 U17448 ( .A1(n29979), .A2(n18896), .Z(n33422) );
  AOI22_X1 U17456 ( .A1(n1442), .A2(n14263), .B1(n1072), .B2(n28105), .ZN(
        n13249) );
  INV_X1 U17475 ( .I(n27249), .ZN(n19918) );
  AOI22_X1 U17479 ( .A1(n27027), .A2(n13213), .B1(n13212), .B2(n27247), .ZN(
        n13211) );
  AOI21_X1 U17482 ( .A1(n8651), .A2(n26961), .B(n8556), .ZN(n7607) );
  INV_X1 U17488 ( .I(n29137), .ZN(n36668) );
  AND2_X2 U17500 ( .A1(n9173), .A2(n35673), .Z(n35186) );
  NOR2_X1 U17503 ( .A1(n5825), .A2(n1379), .ZN(n36677) );
  NAND2_X1 U17506 ( .A1(n33963), .A2(n6938), .ZN(n30222) );
  NOR2_X1 U17514 ( .A1(n29310), .A2(n12876), .ZN(n12878) );
  NAND2_X1 U17546 ( .A1(n23159), .A2(n22935), .ZN(n18865) );
  AND2_X1 U17561 ( .A1(n18042), .A2(n29684), .Z(n18041) );
  NOR2_X1 U17567 ( .A1(n29747), .A2(n29740), .ZN(n29728) );
  NAND2_X1 U17568 ( .A1(n16889), .A2(n14858), .ZN(n36051) );
  NOR2_X1 U17574 ( .A1(n20184), .A2(n28143), .ZN(n20185) );
  NAND2_X1 U17582 ( .A1(n28375), .A2(n29635), .ZN(n36125) );
  INV_X1 U17583 ( .I(n30141), .ZN(n30136) );
  NOR2_X1 U17586 ( .A1(n28131), .A2(n28229), .ZN(n35819) );
  INV_X1 U17588 ( .I(n19891), .ZN(n35659) );
  NAND2_X1 U17591 ( .A1(n8592), .A2(n30047), .ZN(n8591) );
  XNOR2_X1 U17609 ( .A1(n26537), .A2(n26488), .ZN(n36077) );
  INV_X2 U17611 ( .I(n10803), .ZN(n32209) );
  INV_X2 U17613 ( .I(n18240), .ZN(n10803) );
  NAND2_X2 U17619 ( .A1(n53), .A2(n9739), .ZN(n35188) );
  NOR2_X1 U17625 ( .A1(n28224), .A2(n2868), .ZN(n35820) );
  OR2_X2 U17626 ( .A1(n33262), .A2(n33261), .Z(n35189) );
  OR2_X2 U17631 ( .A1(n33262), .A2(n33261), .Z(n35190) );
  INV_X1 U17633 ( .I(n17220), .ZN(n36260) );
  NOR2_X1 U17639 ( .A1(n3003), .A2(n22228), .ZN(n22089) );
  AOI22_X1 U17641 ( .A1(n10868), .A2(n29579), .B1(n10869), .B2(n29580), .ZN(
        n29619) );
  INV_X1 U17644 ( .I(n29815), .ZN(n13574) );
  INV_X2 U17655 ( .I(n4377), .ZN(n30078) );
  NAND2_X1 U17678 ( .A1(n15703), .A2(n26090), .ZN(n10511) );
  INV_X2 U17696 ( .I(n25601), .ZN(n1254) );
  INV_X1 U17698 ( .I(n26651), .ZN(n31254) );
  NAND2_X1 U17708 ( .A1(n11866), .A2(n35622), .ZN(n32142) );
  NAND2_X2 U17712 ( .A1(n8138), .A2(n32506), .ZN(n35196) );
  NOR2_X1 U17717 ( .A1(n9242), .A2(n35469), .ZN(n7839) );
  NAND3_X1 U17720 ( .A1(n7535), .A2(n7534), .A3(n1302), .ZN(n12269) );
  OAI21_X1 U17732 ( .A1(n31107), .A2(n11283), .B(n7690), .ZN(n35862) );
  INV_X1 U17749 ( .I(n26246), .ZN(n10776) );
  XNOR2_X1 U17750 ( .A1(n28830), .A2(n35320), .ZN(n28545) );
  INV_X2 U17759 ( .I(n20156), .ZN(n14278) );
  NAND2_X1 U17760 ( .A1(n4192), .A2(n32046), .ZN(n2429) );
  AND2_X1 U17770 ( .A1(n30173), .A2(n30172), .Z(n35254) );
  INV_X1 U17778 ( .I(n1403), .ZN(n36269) );
  NAND2_X1 U17780 ( .A1(n28720), .A2(n28722), .ZN(n4980) );
  NAND3_X1 U17784 ( .A1(n38073), .A2(n7044), .A3(n34011), .ZN(n18460) );
  OAI21_X1 U17786 ( .A1(n38073), .A2(n37983), .B(n32882), .ZN(n17862) );
  NAND2_X1 U17787 ( .A1(n38073), .A2(n34011), .ZN(n17857) );
  NAND2_X1 U17788 ( .A1(n31328), .A2(n24784), .ZN(n24506) );
  NOR2_X1 U17792 ( .A1(n24784), .A2(n24874), .ZN(n24643) );
  NAND2_X1 U17794 ( .A1(n24784), .A2(n31519), .ZN(n31023) );
  NAND3_X1 U17803 ( .A1(n30822), .A2(n16676), .A3(n20342), .ZN(n11264) );
  NAND3_X1 U17808 ( .A1(n11264), .A2(n11263), .A3(n30168), .ZN(n30971) );
  AND3_X1 U17809 ( .A1(n27338), .A2(n27053), .A3(n27341), .Z(n14692) );
  NOR2_X1 U17810 ( .A1(n20578), .A2(n14601), .ZN(n17466) );
  NAND2_X1 U17845 ( .A1(n28559), .A2(n15792), .ZN(n28561) );
  XNOR2_X1 U17850 ( .A1(n31215), .A2(n14802), .ZN(n35197) );
  AOI21_X1 U17851 ( .A1(n11421), .A2(n34484), .B(n35988), .ZN(n35198) );
  NOR2_X1 U17854 ( .A1(n27441), .A2(n27440), .ZN(n160) );
  INV_X1 U17865 ( .I(n28130), .ZN(n28228) );
  NAND2_X1 U17867 ( .A1(n30780), .A2(n36266), .ZN(n35199) );
  NAND2_X1 U17869 ( .A1(n1068), .A2(n28677), .ZN(n28675) );
  OAI21_X2 U17877 ( .A1(n18464), .A2(n14504), .B(n18463), .ZN(n35200) );
  INV_X1 U17880 ( .I(n33946), .ZN(n32291) );
  NOR2_X1 U17898 ( .A1(n910), .A2(n2678), .ZN(n33032) );
  NOR2_X1 U17904 ( .A1(n1100), .A2(n34265), .ZN(n14650) );
  NOR2_X1 U17911 ( .A1(n25688), .A2(n25587), .ZN(n36412) );
  NAND2_X1 U17913 ( .A1(n4603), .A2(n25587), .ZN(n36592) );
  CLKBUF_X12 U17919 ( .I(n27903), .Z(n19743) );
  NAND2_X1 U17924 ( .A1(n33254), .A2(n27284), .ZN(n35905) );
  OR2_X2 U17925 ( .A1(n7500), .A2(n8128), .Z(n16234) );
  OAI21_X2 U17926 ( .A1(n24968), .A2(n24967), .B(n19574), .ZN(n35202) );
  OAI21_X1 U17931 ( .A1(n29762), .A2(n19568), .B(n29764), .ZN(n29637) );
  CLKBUF_X4 U17939 ( .I(n29044), .Z(n30964) );
  INV_X1 U17940 ( .I(n3827), .ZN(n14412) );
  OAI21_X1 U17965 ( .A1(n31022), .A2(n20531), .B(n200), .ZN(n31001) );
  NAND2_X1 U17970 ( .A1(n14931), .A2(n89), .ZN(n35583) );
  NAND2_X1 U17986 ( .A1(n12288), .A2(n24158), .ZN(n12287) );
  NAND2_X1 U17998 ( .A1(n25978), .A2(n26031), .ZN(n16477) );
  NAND2_X2 U18008 ( .A1(n3248), .A2(n3250), .ZN(n35208) );
  AOI21_X1 U18012 ( .A1(n2629), .A2(n8393), .B(n1742), .ZN(n26275) );
  INV_X1 U18016 ( .I(n28591), .ZN(n28674) );
  XNOR2_X1 U18017 ( .A1(n33962), .A2(n16787), .ZN(n35210) );
  AOI21_X1 U18018 ( .A1(n30055), .A2(n34179), .B(n9918), .ZN(n10671) );
  BUF_X2 U18022 ( .I(n30055), .Z(n19909) );
  OAI21_X1 U18023 ( .A1(n12450), .A2(n29486), .B(n33425), .ZN(n10259) );
  NAND2_X1 U18029 ( .A1(n34006), .A2(n29642), .ZN(n36100) );
  OAI21_X1 U18037 ( .A1(n27349), .A2(n27347), .B(n35767), .ZN(n35766) );
  OAI22_X1 U18039 ( .A1(n30017), .A2(n30024), .B1(n30015), .B2(n15643), .ZN(
        n30013) );
  AOI22_X2 U18043 ( .A1(n36092), .A2(n34128), .B1(n22060), .B2(n8618), .ZN(
        n35211) );
  XOR2_X1 U18060 ( .A1(n16689), .A2(n16687), .Z(n35213) );
  NAND2_X1 U18062 ( .A1(n8235), .A2(n8234), .ZN(n35214) );
  AOI21_X1 U18067 ( .A1(n18406), .A2(n25993), .B(n37613), .ZN(n16247) );
  OAI21_X1 U18068 ( .A1(n23819), .A2(n24116), .B(n38224), .ZN(n14255) );
  AOI21_X2 U18069 ( .A1(n1830), .A2(n23340), .B(n1829), .ZN(n35215) );
  AOI21_X1 U18078 ( .A1(n1830), .A2(n23340), .B(n1829), .ZN(n3503) );
  NAND3_X1 U18082 ( .A1(n17224), .A2(n19559), .A3(n21246), .ZN(n20221) );
  NAND3_X1 U18090 ( .A1(n9591), .A2(n1174), .A3(n19097), .ZN(n21282) );
  NOR2_X1 U18094 ( .A1(n20510), .A2(n30128), .ZN(n35624) );
  INV_X2 U18095 ( .I(n26089), .ZN(n949) );
  XOR2_X1 U18096 ( .A1(n589), .A2(n14835), .Z(n35217) );
  OR3_X2 U18099 ( .A1(n33919), .A2(n20039), .A3(n8430), .Z(n10969) );
  INV_X1 U18109 ( .I(n20039), .ZN(n24787) );
  NAND2_X1 U18110 ( .A1(n21031), .A2(n37048), .ZN(n25479) );
  AOI21_X1 U18115 ( .A1(n33474), .A2(n1098), .B(n26123), .ZN(n26017) );
  INV_X1 U18127 ( .I(n16371), .ZN(n29263) );
  BUF_X2 U18134 ( .I(n16371), .Z(n16123) );
  OR2_X2 U18146 ( .A1(n17597), .A2(n16371), .Z(n19162) );
  INV_X1 U18147 ( .I(n10371), .ZN(n3932) );
  AOI21_X1 U18149 ( .A1(n20538), .A2(n12301), .B(n30176), .ZN(n11263) );
  NAND2_X1 U18151 ( .A1(n1481), .A2(n36840), .ZN(n30588) );
  INV_X1 U18153 ( .I(n27700), .ZN(n36566) );
  NOR2_X1 U18163 ( .A1(n39316), .A2(n33316), .ZN(n2085) );
  NAND2_X1 U18167 ( .A1(n33316), .A2(n35331), .ZN(n12212) );
  NAND2_X1 U18181 ( .A1(n31772), .A2(n13761), .ZN(n10685) );
  INV_X1 U18183 ( .I(n24700), .ZN(n35219) );
  AOI21_X2 U18184 ( .A1(n24531), .A2(n8389), .B(n8388), .ZN(n35220) );
  OAI22_X1 U18189 ( .A1(n36677), .A2(n36676), .B1(n17975), .B2(n17773), .ZN(
        n17974) );
  OR2_X1 U18196 ( .A1(n14800), .A2(n14801), .Z(n35221) );
  AND2_X2 U18204 ( .A1(n35928), .A2(n18378), .Z(n35224) );
  NOR2_X1 U18210 ( .A1(n378), .A2(n33293), .ZN(n14854) );
  NOR2_X1 U18211 ( .A1(n19448), .A2(n21277), .ZN(n20669) );
  NAND2_X1 U18212 ( .A1(n1823), .A2(n28460), .ZN(n32769) );
  XOR2_X1 U18218 ( .A1(n8403), .A2(n8404), .Z(n35225) );
  NAND2_X1 U18224 ( .A1(n35344), .A2(n10143), .ZN(n11776) );
  NAND2_X2 U18225 ( .A1(n19329), .A2(n8210), .ZN(n35229) );
  NAND2_X1 U18234 ( .A1(n10702), .A2(n19544), .ZN(n10703) );
  OAI21_X1 U18236 ( .A1(n5453), .A2(n2799), .B(n4914), .ZN(n5452) );
  AOI21_X1 U18237 ( .A1(n9161), .A2(n17353), .B(n4914), .ZN(n5354) );
  NAND3_X1 U18239 ( .A1(n4914), .A2(n2799), .A3(n728), .ZN(n13465) );
  NAND3_X1 U18240 ( .A1(n954), .A2(n4914), .A3(n10104), .ZN(n2958) );
  INV_X1 U18253 ( .I(n19436), .ZN(n26879) );
  CLKBUF_X4 U18255 ( .I(n5351), .Z(n5239) );
  INV_X1 U18264 ( .I(n23602), .ZN(n35230) );
  AND2_X2 U18271 ( .A1(n34160), .A2(n12836), .Z(n2966) );
  CLKBUF_X2 U18274 ( .I(n15332), .Z(n10013) );
  AND2_X2 U18295 ( .A1(n11296), .A2(n13880), .Z(n28633) );
  CLKBUF_X4 U18314 ( .I(n39489), .Z(n31383) );
  NAND2_X1 U18317 ( .A1(n25867), .A2(n26019), .ZN(n25868) );
  NAND3_X1 U18323 ( .A1(n856), .A2(n26672), .A3(n17217), .ZN(n11227) );
  AOI22_X1 U18328 ( .A1(n35274), .A2(n20357), .B1(n19778), .B2(n3833), .ZN(
        n35231) );
  NAND2_X2 U18344 ( .A1(n23210), .A2(n23209), .ZN(n7014) );
  NOR2_X1 U18347 ( .A1(n24309), .A2(n24446), .ZN(n8681) );
  INV_X2 U18349 ( .I(n24309), .ZN(n24086) );
  NOR2_X1 U18358 ( .A1(n29739), .A2(n29756), .ZN(n29752) );
  INV_X1 U18374 ( .I(n21669), .ZN(n21446) );
  INV_X2 U18384 ( .I(n23929), .ZN(n35235) );
  AOI21_X1 U18387 ( .A1(n7770), .A2(n7769), .B(n38674), .ZN(n30854) );
  NOR2_X1 U18390 ( .A1(n19065), .A2(n29481), .ZN(n16877) );
  INV_X2 U18391 ( .I(n9945), .ZN(n23819) );
  AOI21_X1 U18405 ( .A1(n28137), .A2(n33960), .B(n19667), .ZN(n10266) );
  XOR2_X1 U18412 ( .A1(n1259), .A2(n11698), .Z(n35237) );
  INV_X1 U18423 ( .I(n8407), .ZN(n19590) );
  NOR3_X1 U18430 ( .A1(n25661), .A2(n25660), .A3(n25379), .ZN(n25499) );
  AOI21_X1 U18440 ( .A1(n9277), .A2(n7693), .B(n17087), .ZN(n11121) );
  NAND2_X1 U18441 ( .A1(n10116), .A2(n7693), .ZN(n5390) );
  CLKBUF_X2 U18442 ( .I(n7693), .Z(n35373) );
  INV_X1 U18447 ( .I(n27213), .ZN(n31710) );
  NOR2_X1 U18455 ( .A1(n19580), .A2(n3213), .ZN(n33558) );
  CLKBUF_X4 U18456 ( .I(n25546), .Z(n19701) );
  NOR2_X1 U18467 ( .A1(n4232), .A2(n7023), .ZN(n36247) );
  NOR2_X1 U18468 ( .A1(n17469), .A2(n31527), .ZN(n36421) );
  NAND2_X1 U18473 ( .A1(n861), .A2(n19712), .ZN(n36261) );
  NOR2_X1 U18476 ( .A1(n36716), .A2(n5063), .ZN(n31893) );
  INV_X1 U18478 ( .I(n27357), .ZN(n13754) );
  NOR2_X1 U18484 ( .A1(n29534), .A2(n29531), .ZN(n15233) );
  XNOR2_X1 U18489 ( .A1(n35601), .A2(n32890), .ZN(n35244) );
  AND2_X2 U18493 ( .A1(n16445), .A2(n15933), .Z(n10690) );
  INV_X1 U18497 ( .I(n29616), .ZN(n36548) );
  XNOR2_X1 U18510 ( .A1(n22736), .A2(n4346), .ZN(n35247) );
  NAND2_X1 U18514 ( .A1(n29858), .A2(n29859), .ZN(n29847) );
  NAND2_X1 U18521 ( .A1(n28312), .A2(n5418), .ZN(n35479) );
  OAI22_X1 U18527 ( .A1(n29881), .A2(n17286), .B1(n29880), .B2(n29883), .ZN(
        n10845) );
  OR2_X1 U18531 ( .A1(n17198), .A2(n31596), .Z(n35572) );
  OAI21_X1 U18533 ( .A1(n18384), .A2(n29535), .B(n29532), .ZN(n29490) );
  NOR2_X1 U18538 ( .A1(n22316), .A2(n3863), .ZN(n37011) );
  OAI21_X1 U18551 ( .A1(n19497), .A2(n20672), .B(n29683), .ZN(n29685) );
  XNOR2_X1 U18557 ( .A1(n25146), .A2(n1895), .ZN(n25330) );
  NOR2_X1 U18562 ( .A1(n25539), .A2(n25540), .ZN(n25541) );
  AOI21_X1 U18578 ( .A1(n30786), .A2(n28311), .B(n30785), .ZN(n18931) );
  AOI21_X1 U18581 ( .A1(n841), .A2(n14460), .B(n18164), .ZN(n32867) );
  INV_X1 U18588 ( .I(n20536), .ZN(n36372) );
  INV_X1 U18595 ( .I(n22639), .ZN(n3203) );
  INV_X1 U18600 ( .I(n18920), .ZN(n24407) );
  NAND3_X1 U18615 ( .A1(n20578), .A2(n17237), .A3(n26841), .ZN(n26612) );
  NAND3_X1 U18622 ( .A1(n31161), .A2(n18148), .A3(n35813), .ZN(n17688) );
  NAND3_X2 U18623 ( .A1(n13165), .A2(n25796), .A3(n13164), .ZN(n35251) );
  XOR2_X1 U18624 ( .A1(n21084), .A2(n30956), .Z(n35252) );
  NAND3_X1 U18632 ( .A1(n13165), .A2(n25796), .A3(n13164), .ZN(n26495) );
  INV_X1 U18637 ( .I(n4671), .ZN(n13233) );
  NOR2_X1 U18639 ( .A1(n28655), .A2(n3664), .ZN(n28445) );
  INV_X1 U18647 ( .I(n7464), .ZN(n1915) );
  INV_X1 U18649 ( .I(n3687), .ZN(n30828) );
  NOR2_X1 U18650 ( .A1(n32259), .A2(n3687), .ZN(n11687) );
  OAI21_X1 U18658 ( .A1(n22265), .A2(n22266), .B(n3687), .ZN(n22070) );
  OAI21_X1 U18660 ( .A1(n12023), .A2(n3687), .B(n17307), .ZN(n21263) );
  XOR2_X1 U18666 ( .A1(n5849), .A2(n5851), .Z(n35256) );
  AND2_X2 U18676 ( .A1(n13156), .A2(n14757), .Z(n35258) );
  NAND2_X1 U18699 ( .A1(n29616), .A2(n29623), .ZN(n29622) );
  NAND2_X1 U18709 ( .A1(n29623), .A2(n35273), .ZN(n36382) );
  NOR2_X1 U18712 ( .A1(n29623), .A2(n29616), .ZN(n9046) );
  INV_X1 U18713 ( .I(n31547), .ZN(n31898) );
  INV_X2 U18724 ( .I(n1226), .ZN(n994) );
  NOR2_X1 U18733 ( .A1(n22222), .A2(n1688), .ZN(n17018) );
  NAND2_X1 U18739 ( .A1(n30872), .A2(n877), .ZN(n6978) );
  INV_X1 U18746 ( .I(n10582), .ZN(n9389) );
  NAND3_X1 U18752 ( .A1(n33591), .A2(n5093), .A3(n16108), .ZN(n28718) );
  AND2_X2 U18755 ( .A1(n33546), .A2(n15667), .Z(n35265) );
  OAI21_X1 U18769 ( .A1(n25812), .A2(n25813), .B(n35671), .ZN(n20451) );
  INV_X1 U18772 ( .I(n9267), .ZN(n9295) );
  OAI22_X2 U18776 ( .A1(n27559), .A2(n34360), .B1(n2381), .B2(n2380), .ZN(
        n35266) );
  OAI22_X1 U18779 ( .A1(n27559), .A2(n34360), .B1(n2381), .B2(n2380), .ZN(
        n27851) );
  AOI22_X1 U18784 ( .A1(n24701), .A2(n35219), .B1(n33986), .B2(n13049), .ZN(
        n35267) );
  AOI22_X1 U18793 ( .A1(n24701), .A2(n35219), .B1(n33986), .B2(n13049), .ZN(
        n35268) );
  AOI22_X1 U18795 ( .A1(n24701), .A2(n35219), .B1(n33986), .B2(n13049), .ZN(
        n25240) );
  OAI21_X2 U18799 ( .A1(n11486), .A2(n14667), .B(n26196), .ZN(n35270) );
  XNOR2_X1 U18805 ( .A1(n1886), .A2(n1883), .ZN(n35271) );
  NAND2_X1 U18808 ( .A1(n26134), .A2(n9916), .ZN(n17003) );
  NAND2_X1 U18809 ( .A1(n5311), .A2(n2947), .ZN(n32861) );
  NOR2_X1 U18826 ( .A1(n1478), .A2(n6686), .ZN(n37039) );
  AOI22_X2 U18833 ( .A1(n10868), .A2(n29579), .B1(n10869), .B2(n29580), .ZN(
        n35273) );
  NAND2_X1 U18852 ( .A1(n32691), .A2(n25798), .ZN(n36048) );
  NAND2_X1 U18853 ( .A1(n25797), .A2(n32691), .ZN(n26006) );
  NAND2_X1 U18854 ( .A1(n31899), .A2(n29568), .ZN(n17365) );
  NAND2_X1 U18860 ( .A1(n23625), .A2(n23430), .ZN(n36393) );
  INV_X1 U18862 ( .I(n22854), .ZN(n22928) );
  XOR2_X1 U18881 ( .A1(n36939), .A2(n29817), .Z(n11653) );
  XOR2_X1 U18885 ( .A1(n27663), .A2(n27785), .Z(n3320) );
  XOR2_X1 U18888 ( .A1(n7917), .A2(n11937), .Z(n11938) );
  AOI22_X2 U18895 ( .A1(n7820), .A2(n31787), .B1(n7819), .B2(n4634), .ZN(n7917) );
  OAI21_X1 U18898 ( .A1(n29618), .A2(n35405), .B(n31540), .ZN(n29601) );
  NAND2_X1 U18919 ( .A1(n27357), .A2(n7632), .ZN(n27021) );
  NOR2_X2 U18936 ( .A1(n10977), .A2(n10976), .ZN(n31821) );
  XOR2_X1 U18937 ( .A1(n10662), .A2(n36002), .Z(n2572) );
  AOI22_X2 U18958 ( .A1(n33663), .A2(n3390), .B1(n32012), .B2(n3389), .ZN(
        n36866) );
  NAND2_X2 U18973 ( .A1(n14548), .A2(n35280), .ZN(n11321) );
  XOR2_X1 U18977 ( .A1(n3387), .A2(n20718), .Z(n3386) );
  NAND2_X1 U18982 ( .A1(n1226), .A2(n995), .ZN(n8453) );
  NOR2_X2 U18986 ( .A1(n32444), .A2(n35573), .ZN(n1226) );
  NOR2_X2 U18996 ( .A1(n15465), .A2(n15464), .ZN(n27178) );
  XOR2_X1 U19002 ( .A1(n17703), .A2(n8602), .Z(n2615) );
  XOR2_X1 U19013 ( .A1(n6477), .A2(n16216), .Z(n8247) );
  XOR2_X1 U19029 ( .A1(n22733), .A2(n22734), .Z(n35286) );
  NAND2_X2 U19060 ( .A1(n24585), .A2(n24582), .ZN(n5063) );
  NAND2_X2 U19062 ( .A1(n35294), .A2(n35293), .ZN(n31355) );
  NAND2_X2 U19065 ( .A1(n36705), .A2(n7186), .ZN(n33765) );
  XOR2_X1 U19066 ( .A1(n35255), .A2(n31524), .Z(n19067) );
  NOR2_X2 U19075 ( .A1(n32866), .A2(n5535), .ZN(n7464) );
  NAND2_X1 U19079 ( .A1(n20830), .A2(n29481), .ZN(n18290) );
  NAND2_X2 U19091 ( .A1(n17929), .A2(n17928), .ZN(n13029) );
  NAND3_X1 U19099 ( .A1(n1755), .A2(n36207), .A3(n33861), .ZN(n35330) );
  INV_X2 U19106 ( .I(n2722), .ZN(n27583) );
  AOI22_X2 U19110 ( .A1(n8686), .A2(n7596), .B1(n15142), .B2(n9646), .ZN(n2722) );
  INV_X2 U19119 ( .I(n35300), .ZN(n800) );
  OR2_X2 U19151 ( .A1(n21933), .A2(n36062), .Z(n21932) );
  BUF_X2 U19152 ( .I(n27792), .Z(n35303) );
  OAI21_X2 U19156 ( .A1(n16282), .A2(n16283), .B(n16281), .ZN(n32886) );
  NAND2_X2 U19159 ( .A1(n22814), .A2(n22815), .ZN(n35534) );
  AOI21_X2 U19160 ( .A1(n4349), .A2(n4350), .B(n31714), .ZN(n24495) );
  XOR2_X1 U19166 ( .A1(n11236), .A2(n27204), .Z(n9196) );
  XOR2_X1 U19180 ( .A1(n18833), .A2(n21163), .Z(n33152) );
  XNOR2_X1 U19181 ( .A1(n26571), .A2(n12221), .ZN(n12903) );
  MUX2_X1 U19189 ( .I0(n12396), .I1(n39001), .S(n23517), .Z(n17788) );
  XOR2_X1 U19202 ( .A1(n18857), .A2(n24024), .Z(n17000) );
  AOI21_X2 U19205 ( .A1(n28202), .A2(n28203), .B(n35309), .ZN(n28680) );
  OAI21_X2 U19213 ( .A1(n4107), .A2(n14750), .B(n35310), .ZN(n23358) );
  XOR2_X1 U19214 ( .A1(n22735), .A2(n22663), .Z(n3800) );
  XOR2_X1 U19222 ( .A1(n2233), .A2(n19094), .Z(n22735) );
  AOI21_X2 U19244 ( .A1(n6381), .A2(n21787), .B(n35315), .ZN(n31960) );
  AND2_X1 U19245 ( .A1(n21659), .A2(n21660), .Z(n35315) );
  AOI21_X2 U19270 ( .A1(n11187), .A2(n23477), .B(n35322), .ZN(n11183) );
  XOR2_X1 U19283 ( .A1(n16191), .A2(n35323), .Z(n30607) );
  XOR2_X1 U19290 ( .A1(n16190), .A2(n34139), .Z(n35323) );
  NAND2_X2 U19301 ( .A1(n8106), .A2(n8107), .ZN(n35900) );
  XOR2_X1 U19303 ( .A1(n28870), .A2(n35324), .Z(n35857) );
  AOI22_X2 U19313 ( .A1(n35326), .A2(n16206), .B1(n4871), .B2(n28548), .ZN(
        n15780) );
  OAI21_X2 U19314 ( .A1(n14631), .A2(n25373), .B(n25327), .ZN(n35327) );
  NAND2_X2 U19348 ( .A1(n17739), .A2(n11388), .ZN(n8627) );
  XOR2_X1 U19352 ( .A1(n25184), .A2(n25176), .Z(n25310) );
  NAND2_X2 U19353 ( .A1(n17904), .A2(n24813), .ZN(n25184) );
  XOR2_X1 U19354 ( .A1(n20065), .A2(n215), .Z(n35543) );
  NOR2_X1 U19356 ( .A1(n27590), .A2(n27591), .ZN(n35334) );
  INV_X4 U19357 ( .I(n11678), .ZN(n35377) );
  AOI22_X2 U19358 ( .A1(n35335), .A2(n20815), .B1(n7052), .B2(n591), .ZN(
        n35448) );
  NOR2_X2 U19359 ( .A1(n6696), .A2(n2366), .ZN(n35335) );
  XOR2_X1 U19361 ( .A1(n2623), .A2(n2622), .Z(n25488) );
  XOR2_X1 U19362 ( .A1(n26211), .A2(n19900), .Z(n26836) );
  AOI22_X1 U19363 ( .A1(n11446), .A2(n11448), .B1(n32079), .B2(n32508), .ZN(
        n35340) );
  XOR2_X1 U19364 ( .A1(n29124), .A2(n28874), .Z(n28916) );
  NAND3_X1 U19370 ( .A1(n14519), .A2(n20605), .A3(n33012), .ZN(n35336) );
  AOI22_X2 U19376 ( .A1(n7908), .A2(n11803), .B1(n36328), .B2(n11429), .ZN(
        n7907) );
  XOR2_X1 U19392 ( .A1(n8922), .A2(n8923), .Z(n11780) );
  XOR2_X1 U19396 ( .A1(n24933), .A2(n34564), .Z(n24974) );
  NAND2_X1 U19399 ( .A1(n35500), .A2(n17132), .ZN(n8931) );
  XOR2_X1 U19410 ( .A1(n25262), .A2(n30519), .Z(n12749) );
  XOR2_X1 U19423 ( .A1(n35340), .A2(n30130), .Z(Ciphertext[167]) );
  INV_X2 U19426 ( .I(n33252), .ZN(n35627) );
  OAI21_X1 U19438 ( .A1(n29956), .A2(n29863), .B(n10679), .ZN(n35342) );
  XOR2_X1 U19439 ( .A1(n35343), .A2(n31815), .Z(n22942) );
  XOR2_X1 U19441 ( .A1(n11887), .A2(n34132), .Z(n36971) );
  NAND2_X2 U19443 ( .A1(n27198), .A2(n4353), .ZN(n27397) );
  INV_X2 U19444 ( .I(n26039), .ZN(n25830) );
  NAND2_X2 U19445 ( .A1(n35371), .A2(n2248), .ZN(n26039) );
  XOR2_X1 U19453 ( .A1(n5917), .A2(n9948), .Z(n32026) );
  NOR2_X2 U19457 ( .A1(n1129), .A2(n24360), .ZN(n11361) );
  AOI21_X2 U19467 ( .A1(n30355), .A2(n5935), .B(n35345), .ZN(n31959) );
  XOR2_X1 U19475 ( .A1(n12762), .A2(n12760), .Z(n14287) );
  NAND2_X2 U19486 ( .A1(n71), .A2(n70), .ZN(n30574) );
  INV_X2 U19500 ( .I(n16260), .ZN(n29412) );
  NAND2_X2 U19504 ( .A1(n12067), .A2(n35348), .ZN(n24877) );
  NAND2_X2 U19506 ( .A1(n17095), .A2(n31014), .ZN(n27402) );
  XOR2_X1 U19512 ( .A1(n13724), .A2(n21323), .Z(n13794) );
  NAND2_X2 U19513 ( .A1(n35353), .A2(n38168), .ZN(n32999) );
  XOR2_X1 U19523 ( .A1(n5918), .A2(n5920), .Z(n8250) );
  NAND2_X1 U19526 ( .A1(n35813), .A2(n8430), .ZN(n8426) );
  NAND2_X2 U19529 ( .A1(n35355), .A2(n23500), .ZN(n17937) );
  NAND2_X2 U19533 ( .A1(n11323), .A2(n11322), .ZN(n19759) );
  XOR2_X1 U19537 ( .A1(n29127), .A2(n29050), .Z(n29292) );
  NOR2_X1 U19555 ( .A1(n11296), .A2(n975), .ZN(n2823) );
  NAND2_X2 U19559 ( .A1(n6978), .A2(n6980), .ZN(n13880) );
  INV_X4 U19579 ( .I(n27349), .ZN(n993) );
  NAND2_X2 U19584 ( .A1(n583), .A2(n21008), .ZN(n27349) );
  XOR2_X1 U19595 ( .A1(Plaintext[8]), .A2(Key[8]), .Z(n35359) );
  XOR2_X1 U19597 ( .A1(n14110), .A2(n14109), .Z(n23189) );
  AOI22_X2 U19600 ( .A1(n29458), .A2(n19065), .B1(n29454), .B2(n29455), .ZN(
        n12479) );
  NAND2_X2 U19606 ( .A1(n12426), .A2(n12175), .ZN(n35376) );
  NAND2_X1 U19614 ( .A1(n14477), .A2(n33840), .ZN(n23547) );
  NAND2_X2 U19615 ( .A1(n12508), .A2(n36001), .ZN(n14477) );
  NOR2_X1 U19618 ( .A1(n31673), .A2(n35450), .ZN(n14509) );
  AOI22_X1 U19624 ( .A1(n30028), .A2(n30027), .B1(n33311), .B2(n30031), .ZN(
        n18313) );
  AND2_X1 U19630 ( .A1(n3092), .A2(n27484), .Z(n20528) );
  AOI22_X2 U19637 ( .A1(n6472), .A2(n35696), .B1(n8494), .B2(n18810), .ZN(
        n35362) );
  XOR2_X1 U19650 ( .A1(n4209), .A2(n35363), .Z(n36390) );
  XOR2_X1 U19651 ( .A1(n2126), .A2(n12437), .Z(n35363) );
  XOR2_X1 U19656 ( .A1(n27478), .A2(n27850), .Z(n27606) );
  NAND2_X2 U19657 ( .A1(n11040), .A2(n11037), .ZN(n27850) );
  XOR2_X1 U19663 ( .A1(n27495), .A2(n27833), .Z(n27646) );
  XNOR2_X1 U19664 ( .A1(n39161), .A2(n23996), .ZN(n6291) );
  NOR3_X1 U19682 ( .A1(n25498), .A2(n15036), .A3(n14401), .ZN(n25382) );
  XOR2_X1 U19695 ( .A1(n36971), .A2(n6880), .Z(n31078) );
  NOR2_X1 U19697 ( .A1(n28742), .A2(n17583), .ZN(n35370) );
  OAI21_X2 U19702 ( .A1(n35931), .A2(n33669), .B(n35374), .ZN(n33283) );
  NAND2_X2 U19723 ( .A1(n8656), .A2(n6694), .ZN(n8532) );
  XOR2_X1 U19734 ( .A1(n13001), .A2(n5284), .Z(n411) );
  AOI21_X2 U19735 ( .A1(n14588), .A2(n30434), .B(n27231), .ZN(n18641) );
  OAI22_X2 U19737 ( .A1(n27898), .A2(n28594), .B1(n7905), .B2(n31088), .ZN(
        n16357) );
  AOI21_X2 U19750 ( .A1(n14410), .A2(n1024), .B(n31574), .ZN(n2461) );
  NAND2_X2 U19752 ( .A1(n35467), .A2(n8737), .ZN(n8683) );
  AOI21_X2 U19762 ( .A1(n17744), .A2(n36210), .B(n35386), .ZN(n17742) );
  NOR3_X2 U19763 ( .A1(n14901), .A2(n23552), .A3(n34012), .ZN(n35386) );
  NAND2_X2 U19764 ( .A1(n35387), .A2(n6087), .ZN(n8668) );
  OAI21_X2 U19766 ( .A1(n22956), .A2(n22958), .B(n22955), .ZN(n35387) );
  XOR2_X1 U19769 ( .A1(n27834), .A2(n30104), .Z(n35389) );
  AND2_X1 U19772 ( .A1(n24866), .A2(n36385), .Z(n24499) );
  NAND2_X2 U19773 ( .A1(n24324), .A2(n24323), .ZN(n24866) );
  XOR2_X1 U19774 ( .A1(n6164), .A2(n35390), .Z(n11) );
  XOR2_X1 U19778 ( .A1(n14098), .A2(n3140), .Z(n35390) );
  OAI21_X2 U19781 ( .A1(n5306), .A2(n19480), .B(n35391), .ZN(n30210) );
  NAND3_X1 U19784 ( .A1(n17104), .A2(n35180), .A3(n17103), .ZN(n35392) );
  OAI21_X2 U19787 ( .A1(n10468), .A2(n34723), .B(n1580), .ZN(n9528) );
  AOI22_X2 U19789 ( .A1(n35394), .A2(n38303), .B1(n31270), .B2(n5), .ZN(n5613)
         );
  NAND2_X2 U19810 ( .A1(n18224), .A2(n18223), .ZN(n28560) );
  AND2_X1 U19813 ( .A1(n29880), .A2(n10294), .Z(n31968) );
  INV_X2 U19818 ( .I(n35395), .ZN(n20359) );
  AOI21_X2 U19832 ( .A1(n13010), .A2(n9350), .B(n39316), .ZN(n9349) );
  OAI21_X2 U19837 ( .A1(n14474), .A2(n17018), .B(n196), .ZN(n35400) );
  NAND2_X2 U19840 ( .A1(n33485), .A2(n35401), .ZN(n35992) );
  INV_X1 U19842 ( .I(n35402), .ZN(n1785) );
  AOI21_X1 U19846 ( .A1(n6274), .A2(n6491), .B(n6273), .ZN(n35402) );
  INV_X1 U19852 ( .I(n9360), .ZN(n35841) );
  OR2_X1 U19854 ( .A1(n33948), .A2(n31250), .Z(n19964) );
  OR2_X1 U19870 ( .A1(n29622), .A2(n35405), .Z(n17176) );
  XOR2_X1 U19897 ( .A1(n23887), .A2(n23713), .Z(n6277) );
  INV_X2 U19905 ( .I(n35407), .ZN(n8556) );
  XNOR2_X1 U19908 ( .A1(n8557), .A2(n26373), .ZN(n35407) );
  NAND2_X1 U19934 ( .A1(n11838), .A2(n38579), .ZN(n35414) );
  NAND2_X1 U19936 ( .A1(n7220), .A2(n7219), .ZN(n35415) );
  XNOR2_X1 U19940 ( .A1(n1669), .A2(n11541), .ZN(n35642) );
  XOR2_X1 U19942 ( .A1(n6572), .A2(n31791), .Z(n7787) );
  NAND2_X2 U19945 ( .A1(n1865), .A2(n1864), .ZN(n22620) );
  XOR2_X1 U19956 ( .A1(n6460), .A2(n24150), .Z(n31348) );
  NAND2_X1 U19960 ( .A1(n15301), .A2(n1403), .ZN(n36403) );
  XOR2_X1 U19963 ( .A1(n18886), .A2(n28933), .Z(n431) );
  NAND2_X2 U19965 ( .A1(n32186), .A2(n16576), .ZN(n27571) );
  NAND2_X2 U19970 ( .A1(n1351), .A2(n17938), .ZN(n21497) );
  NAND3_X1 U19974 ( .A1(n31184), .A2(n30368), .A3(n24406), .ZN(n30850) );
  AOI22_X2 U19979 ( .A1(n37257), .A2(n28246), .B1(n37451), .B2(n19003), .ZN(
        n35420) );
  XOR2_X1 U19980 ( .A1(n8957), .A2(n27569), .Z(n35421) );
  NAND3_X2 U19981 ( .A1(n1763), .A2(n23167), .A3(n22975), .ZN(n20564) );
  NAND3_X2 U19984 ( .A1(n1906), .A2(n35735), .A3(n30635), .ZN(n35422) );
  AOI22_X2 U19986 ( .A1(n35424), .A2(n19132), .B1(n35423), .B2(n1221), .ZN(
        n27785) );
  XOR2_X1 U19993 ( .A1(n24025), .A2(n19904), .Z(n11180) );
  NAND2_X2 U19995 ( .A1(n35600), .A2(n321), .ZN(n24025) );
  XOR2_X1 U19998 ( .A1(n11828), .A2(n16439), .Z(n35425) );
  NAND2_X1 U20013 ( .A1(n22928), .A2(n22994), .ZN(n22555) );
  NAND2_X1 U20014 ( .A1(n20616), .A2(n170), .ZN(n29993) );
  XOR2_X1 U20016 ( .A1(n9043), .A2(n18279), .Z(n33010) );
  NAND3_X2 U20020 ( .A1(n3275), .A2(n3276), .A3(n3274), .ZN(n9043) );
  BUF_X4 U20027 ( .I(n8267), .Z(n35921) );
  AOI21_X1 U20044 ( .A1(n18783), .A2(n18782), .B(n30037), .ZN(n36848) );
  NOR2_X1 U20048 ( .A1(n4964), .A2(n35427), .ZN(n32696) );
  OAI21_X2 U20059 ( .A1(n7212), .A2(n22496), .B(n36660), .ZN(n35920) );
  NAND2_X2 U20084 ( .A1(n12993), .A2(n12991), .ZN(n11067) );
  AND2_X1 U20088 ( .A1(n33980), .A2(n12187), .Z(n19003) );
  XOR2_X1 U20103 ( .A1(n35435), .A2(n14046), .Z(n35769) );
  NAND2_X2 U20110 ( .A1(n6252), .A2(n29558), .ZN(n29543) );
  NAND2_X2 U20112 ( .A1(n6253), .A2(n14850), .ZN(n29558) );
  XOR2_X1 U20131 ( .A1(n18106), .A2(n26605), .Z(n36915) );
  XOR2_X1 U20133 ( .A1(n8833), .A2(n17757), .Z(n26605) );
  XOR2_X1 U20137 ( .A1(n35746), .A2(n35747), .Z(n4256) );
  NAND2_X2 U20141 ( .A1(n35437), .A2(n14995), .ZN(n21864) );
  INV_X4 U20160 ( .I(n23350), .ZN(n36027) );
  XOR2_X1 U20170 ( .A1(n27837), .A2(n3207), .Z(n35438) );
  AOI21_X2 U20171 ( .A1(n16750), .A2(n16749), .B(n35439), .ZN(n7728) );
  OAI22_X2 U20185 ( .A1(n20414), .A2(n3120), .B1(n24849), .B2(n33344), .ZN(
        n35439) );
  NAND3_X2 U20187 ( .A1(n27124), .A2(n27125), .A3(n27129), .ZN(n16736) );
  NOR2_X1 U20189 ( .A1(n35679), .A2(n25770), .ZN(n30568) );
  NAND2_X1 U20203 ( .A1(n38395), .A2(n17864), .ZN(n64) );
  NOR2_X2 U20205 ( .A1(n10295), .A2(n35441), .ZN(n23634) );
  INV_X2 U20209 ( .I(n29005), .ZN(n4095) );
  XOR2_X1 U20211 ( .A1(n3938), .A2(n34183), .Z(n29005) );
  AOI22_X2 U20216 ( .A1(n12891), .A2(n12890), .B1(n36609), .B2(n34172), .ZN(
        n12889) );
  XOR2_X1 U20225 ( .A1(n12857), .A2(n7673), .Z(n35836) );
  XOR2_X1 U20229 ( .A1(n35446), .A2(n22438), .Z(n35445) );
  XOR2_X1 U20231 ( .A1(n29253), .A2(n9930), .Z(n16553) );
  NAND4_X2 U20232 ( .A1(n22820), .A2(n7683), .A3(n18856), .A4(n31748), .ZN(
        n18204) );
  NAND3_X2 U20235 ( .A1(n17971), .A2(n24778), .A3(n24777), .ZN(n16627) );
  NAND2_X2 U20241 ( .A1(n16700), .A2(n31638), .ZN(n31287) );
  INV_X2 U20250 ( .I(n35450), .ZN(n30279) );
  XNOR2_X1 U20251 ( .A1(n20516), .A2(n20716), .ZN(n35450) );
  NAND3_X2 U20273 ( .A1(n36785), .A2(n16098), .A3(n23338), .ZN(n23658) );
  INV_X1 U20274 ( .I(n32630), .ZN(n35569) );
  NOR2_X2 U20277 ( .A1(n35452), .A2(n7859), .ZN(n31862) );
  NOR2_X2 U20281 ( .A1(n20404), .A2(n33788), .ZN(n5955) );
  NAND2_X2 U20284 ( .A1(n35454), .A2(n25810), .ZN(n26437) );
  NAND2_X2 U20285 ( .A1(n3153), .A2(n3857), .ZN(n30076) );
  AOI21_X2 U20286 ( .A1(n22015), .A2(n20034), .B(n22165), .ZN(n35734) );
  INV_X2 U20299 ( .I(n35455), .ZN(n14418) );
  XOR2_X1 U20301 ( .A1(Plaintext[138]), .A2(Key[138]), .Z(n35455) );
  XOR2_X1 U20307 ( .A1(n35457), .A2(n22667), .Z(n10963) );
  INV_X2 U20333 ( .I(n35462), .ZN(n24155) );
  NOR2_X2 U20336 ( .A1(n12064), .A2(n19142), .ZN(n35462) );
  INV_X2 U20337 ( .I(n15047), .ZN(n17197) );
  NAND2_X1 U20342 ( .A1(n36623), .A2(n28729), .ZN(n15296) );
  XOR2_X1 U20343 ( .A1(n35463), .A2(n26480), .Z(n30551) );
  NAND2_X2 U20346 ( .A1(n9087), .A2(n9086), .ZN(n26480) );
  INV_X2 U20347 ( .I(n27532), .ZN(n35464) );
  NAND2_X1 U20348 ( .A1(n20724), .A2(n29410), .ZN(n35677) );
  XOR2_X1 U20365 ( .A1(n19064), .A2(n25007), .Z(n10717) );
  XOR2_X1 U20367 ( .A1(n12430), .A2(n3395), .Z(n35468) );
  INV_X2 U20370 ( .I(n31971), .ZN(n35469) );
  OAI22_X2 U20375 ( .A1(n3714), .A2(n32351), .B1(n2928), .B2(n3715), .ZN(
        n35470) );
  XOR2_X1 U20376 ( .A1(n3330), .A2(n35471), .Z(n36334) );
  XOR2_X1 U20378 ( .A1(n35472), .A2(n25033), .Z(n8713) );
  XOR2_X1 U20380 ( .A1(n24997), .A2(n25290), .Z(n25033) );
  XOR2_X1 U20387 ( .A1(n7337), .A2(n35532), .Z(n10380) );
  XOR2_X1 U20390 ( .A1(n22766), .A2(n22624), .Z(n7337) );
  NOR2_X1 U20391 ( .A1(n35474), .A2(n22253), .ZN(n17409) );
  NAND2_X1 U20393 ( .A1(n12930), .A2(n10242), .ZN(n35474) );
  INV_X2 U20396 ( .I(n35476), .ZN(n2752) );
  XOR2_X1 U20398 ( .A1(n2754), .A2(n2753), .Z(n35476) );
  XOR2_X1 U20410 ( .A1(n38191), .A2(n12480), .Z(n35480) );
  XOR2_X1 U20411 ( .A1(n24026), .A2(n5238), .Z(n35481) );
  NAND3_X2 U20414 ( .A1(n35483), .A2(n39813), .A3(n13580), .ZN(n10638) );
  XNOR2_X1 U20426 ( .A1(n17727), .A2(n22562), .ZN(n22733) );
  NAND2_X2 U20429 ( .A1(n6723), .A2(n6721), .ZN(n22562) );
  XNOR2_X1 U20436 ( .A1(n26455), .A2(n29785), .ZN(n36511) );
  NOR2_X2 U20450 ( .A1(n4147), .A2(n17887), .ZN(n4148) );
  INV_X2 U20457 ( .I(n31474), .ZN(n35705) );
  XOR2_X1 U20460 ( .A1(n4131), .A2(n36264), .Z(n31474) );
  XOR2_X1 U20461 ( .A1(n39161), .A2(n19629), .Z(n23924) );
  AOI21_X2 U20467 ( .A1(n24506), .A2(n9212), .B(n36017), .ZN(n18393) );
  NAND2_X1 U20479 ( .A1(n14396), .A2(n19586), .ZN(n15080) );
  NOR2_X2 U20480 ( .A1(n31037), .A2(n35487), .ZN(n23969) );
  OAI22_X2 U20481 ( .A1(n23621), .A2(n33496), .B1(n23284), .B2(n23452), .ZN(
        n35487) );
  XOR2_X1 U20487 ( .A1(n35490), .A2(n2743), .Z(n2742) );
  XOR2_X1 U20488 ( .A1(n33806), .A2(n22382), .Z(n35490) );
  OAI22_X2 U20489 ( .A1(n13306), .A2(n13304), .B1(n32616), .B2(n30274), .ZN(
        n23963) );
  NAND2_X2 U20490 ( .A1(n28345), .A2(n28347), .ZN(n28717) );
  XOR2_X1 U20505 ( .A1(n36863), .A2(n35494), .Z(n33553) );
  XOR2_X1 U20506 ( .A1(n27763), .A2(n27762), .Z(n35494) );
  XOR2_X1 U20513 ( .A1(n32200), .A2(n29247), .Z(n12853) );
  OR2_X1 U20516 ( .A1(n11728), .A2(n18246), .Z(n35495) );
  NAND2_X2 U20517 ( .A1(n28140), .A2(n28139), .ZN(n35496) );
  XOR2_X1 U20518 ( .A1(n26521), .A2(n35498), .Z(n11740) );
  XOR2_X1 U20519 ( .A1(n31941), .A2(n26407), .Z(n35498) );
  AND2_X1 U20521 ( .A1(n28586), .A2(n11030), .Z(n36031) );
  XOR2_X1 U20523 ( .A1(n18635), .A2(n5203), .Z(n31933) );
  XOR2_X1 U20525 ( .A1(n22784), .A2(n1710), .Z(n12516) );
  XOR2_X1 U20526 ( .A1(n14388), .A2(n16553), .Z(n16552) );
  NAND2_X1 U20529 ( .A1(n10171), .A2(n27304), .ZN(n35906) );
  INV_X2 U20543 ( .I(n32854), .ZN(n35506) );
  INV_X1 U20546 ( .I(n16203), .ZN(n35508) );
  NOR2_X1 U20551 ( .A1(n11030), .A2(n36076), .ZN(n36032) );
  OR2_X1 U20552 ( .A1(n8527), .A2(n38591), .Z(n26443) );
  XOR2_X1 U20564 ( .A1(n25293), .A2(n35511), .Z(n35510) );
  NAND2_X1 U20567 ( .A1(n33086), .A2(n22264), .ZN(n35513) );
  NAND3_X1 U20591 ( .A1(n15215), .A2(n9594), .A3(n16114), .ZN(n35763) );
  AOI21_X1 U20598 ( .A1(n29389), .A2(n29497), .B(n36275), .ZN(n35517) );
  NAND2_X2 U20599 ( .A1(n6954), .A2(n6953), .ZN(n7552) );
  NOR2_X1 U20614 ( .A1(n24795), .A2(n16238), .ZN(n35520) );
  XOR2_X1 U20615 ( .A1(n11207), .A2(n29306), .Z(n35728) );
  NOR2_X2 U20626 ( .A1(n20102), .A2(n30059), .ZN(n6496) );
  NAND2_X1 U20631 ( .A1(n39676), .A2(n26109), .ZN(n25790) );
  XOR2_X1 U20639 ( .A1(n8371), .A2(n36828), .Z(n4898) );
  AOI21_X2 U20668 ( .A1(n14355), .A2(n26833), .B(n7527), .ZN(n26772) );
  NAND2_X1 U20670 ( .A1(n39155), .A2(n18708), .ZN(n9507) );
  NAND2_X2 U20678 ( .A1(n35689), .A2(n1642), .ZN(n23392) );
  XOR2_X1 U20695 ( .A1(n21207), .A2(n7380), .Z(n25552) );
  NAND2_X2 U20704 ( .A1(n22119), .A2(n22116), .ZN(n3687) );
  AOI22_X2 U20705 ( .A1(n2164), .A2(n31198), .B1(n31257), .B2(n35968), .ZN(
        n25303) );
  NOR2_X1 U20726 ( .A1(n13555), .A2(n11449), .ZN(n6170) );
  NAND2_X1 U20729 ( .A1(n19204), .A2(n14636), .ZN(n35535) );
  BUF_X2 U20730 ( .I(n23250), .Z(n35536) );
  OAI21_X2 U20735 ( .A1(n10452), .A2(n31958), .B(n35541), .ZN(n17849) );
  XOR2_X1 U20737 ( .A1(n27538), .A2(n34094), .Z(n35542) );
  INV_X1 U20738 ( .I(n35233), .ZN(n12248) );
  NOR2_X2 U20748 ( .A1(n22396), .A2(n22397), .ZN(n22408) );
  XOR2_X1 U20766 ( .A1(n22517), .A2(n4123), .Z(n22382) );
  XOR2_X1 U20772 ( .A1(n35544), .A2(n27784), .Z(n33522) );
  XOR2_X1 U20786 ( .A1(n5153), .A2(n29145), .Z(n1740) );
  NAND2_X2 U20787 ( .A1(n28752), .A2(n28751), .ZN(n29145) );
  AND2_X1 U20791 ( .A1(n35550), .A2(n33538), .Z(n17787) );
  NAND2_X1 U20794 ( .A1(n23517), .A2(n19671), .ZN(n35550) );
  NAND3_X2 U20801 ( .A1(n31168), .A2(n16435), .A3(n35553), .ZN(n22728) );
  AOI22_X1 U20802 ( .A1(n10651), .A2(n9876), .B1(n22341), .B2(n15350), .ZN(
        n35553) );
  XOR2_X1 U20803 ( .A1(n8909), .A2(n774), .Z(n35554) );
  NAND2_X2 U20818 ( .A1(n17819), .A2(n17820), .ZN(n21802) );
  XOR2_X1 U20821 ( .A1(n4442), .A2(n35556), .Z(n10455) );
  XOR2_X1 U20822 ( .A1(n22609), .A2(n20350), .Z(n35556) );
  NAND2_X2 U20828 ( .A1(n28460), .A2(n28378), .ZN(n31390) );
  NAND2_X2 U20842 ( .A1(n10), .A2(n14066), .ZN(n33840) );
  NOR2_X1 U20858 ( .A1(n21914), .A2(n938), .ZN(n21915) );
  XOR2_X1 U20863 ( .A1(n19194), .A2(n10413), .Z(n10427) );
  NAND2_X1 U20887 ( .A1(n16832), .A2(n10733), .ZN(n36852) );
  NAND2_X2 U20889 ( .A1(n35563), .A2(n27938), .ZN(n16108) );
  NAND2_X1 U20890 ( .A1(n33613), .A2(n33611), .ZN(n35563) );
  NAND2_X2 U20918 ( .A1(n23355), .A2(n37523), .ZN(n23248) );
  XOR2_X1 U20925 ( .A1(n35566), .A2(n34062), .Z(n36454) );
  XOR2_X1 U20930 ( .A1(n6034), .A2(n5055), .Z(n35566) );
  XOR2_X1 U20931 ( .A1(n8183), .A2(n35267), .Z(n24702) );
  NOR2_X2 U20941 ( .A1(n33032), .A2(n7258), .ZN(n35568) );
  NOR2_X2 U20946 ( .A1(n21420), .A2(n21419), .ZN(n36371) );
  AOI21_X1 U20953 ( .A1(n29645), .A2(n35572), .B(n37879), .ZN(n17383) );
  NAND2_X2 U20958 ( .A1(n22000), .A2(n20298), .ZN(n17189) );
  NAND2_X2 U20962 ( .A1(n17882), .A2(n15652), .ZN(n22484) );
  XOR2_X1 U20982 ( .A1(n2387), .A2(n2388), .Z(n31403) );
  NOR2_X1 U20983 ( .A1(n7445), .A2(n36321), .ZN(n20029) );
  NAND2_X2 U20989 ( .A1(n35948), .A2(n16184), .ZN(n36321) );
  NAND2_X2 U21018 ( .A1(n24662), .A2(n35578), .ZN(n35577) );
  NOR2_X1 U21028 ( .A1(n18383), .A2(n14456), .ZN(n19242) );
  XOR2_X1 U21034 ( .A1(n3709), .A2(n5255), .Z(n33057) );
  XOR2_X1 U21042 ( .A1(n5652), .A2(n15960), .Z(n18886) );
  NAND2_X2 U21045 ( .A1(n6809), .A2(n30748), .ZN(n5652) );
  NAND2_X2 U21061 ( .A1(n6712), .A2(n35584), .ZN(n23433) );
  AOI21_X2 U21065 ( .A1(n22996), .A2(n35586), .B(n35585), .ZN(n35584) );
  NOR2_X2 U21076 ( .A1(n23163), .A2(n35586), .ZN(n35585) );
  INV_X2 U21079 ( .I(n23164), .ZN(n35586) );
  INV_X2 U21086 ( .I(n23530), .ZN(n23528) );
  NAND4_X2 U21088 ( .A1(n33832), .A2(n20741), .A3(n20744), .A4(n5464), .ZN(
        n23530) );
  XOR2_X1 U21090 ( .A1(n12853), .A2(n3297), .Z(n12055) );
  OR2_X1 U21100 ( .A1(n37230), .A2(n33788), .Z(n24483) );
  NOR2_X2 U21121 ( .A1(n8190), .A2(n23374), .ZN(n35594) );
  OAI21_X1 U21124 ( .A1(n16880), .A2(n5061), .B(n36425), .ZN(n9715) );
  NOR2_X2 U21126 ( .A1(n12511), .A2(n12512), .ZN(n16880) );
  XOR2_X1 U21134 ( .A1(n35595), .A2(n18255), .Z(n30455) );
  XOR2_X1 U21144 ( .A1(n37042), .A2(n35596), .Z(n35595) );
  INV_X2 U21153 ( .I(n22527), .ZN(n35596) );
  NAND2_X2 U21160 ( .A1(n12394), .A2(n7866), .ZN(n25691) );
  NAND2_X2 U21161 ( .A1(n35598), .A2(n5292), .ZN(n14890) );
  NAND2_X2 U21164 ( .A1(n25568), .A2(n25692), .ZN(n35598) );
  XOR2_X1 U21166 ( .A1(n35599), .A2(n26369), .Z(n19810) );
  XOR2_X1 U21167 ( .A1(n26432), .A2(n16169), .Z(n35599) );
  OR2_X2 U21169 ( .A1(n17464), .A2(n5975), .Z(n23072) );
  BUF_X4 U21175 ( .I(n7520), .Z(n35960) );
  AOI22_X2 U21178 ( .A1(n36137), .A2(n38244), .B1(n37209), .B2(n19686), .ZN(
        n35600) );
  XOR2_X1 U21181 ( .A1(n35601), .A2(n32890), .Z(n33788) );
  XOR2_X1 U21198 ( .A1(n11794), .A2(n5005), .Z(n36000) );
  NAND3_X2 U21201 ( .A1(n19670), .A2(n24965), .A3(n16819), .ZN(n30520) );
  XOR2_X1 U21221 ( .A1(n5463), .A2(n22667), .Z(n9137) );
  NAND2_X2 U21234 ( .A1(n12816), .A2(n22965), .ZN(n23496) );
  BUF_X2 U21241 ( .I(n27852), .Z(n35610) );
  XOR2_X1 U21245 ( .A1(n9449), .A2(n9448), .Z(n35614) );
  NOR2_X1 U21248 ( .A1(n38839), .A2(n17790), .ZN(n8201) );
  OAI21_X2 U21250 ( .A1(n14326), .A2(n2760), .B(n35616), .ZN(n2281) );
  NOR2_X2 U21257 ( .A1(n8927), .A2(n35619), .ZN(n33493) );
  NOR3_X2 U21262 ( .A1(n1125), .A2(n9371), .A3(n35890), .ZN(n35619) );
  XOR2_X1 U21267 ( .A1(n8469), .A2(n8471), .Z(n29149) );
  NAND2_X2 U21268 ( .A1(n21786), .A2(n35623), .ZN(n22294) );
  XOR2_X1 U21275 ( .A1(n27500), .A2(n26916), .Z(n35626) );
  XOR2_X1 U21288 ( .A1(n26593), .A2(n36383), .Z(n15674) );
  XOR2_X1 U21289 ( .A1(n26340), .A2(n6757), .Z(n26593) );
  OAI22_X1 U21291 ( .A1(n29414), .A2(n29413), .B1(n29415), .B2(n29416), .ZN(
        n29417) );
  XOR2_X1 U21298 ( .A1(n25237), .A2(n11964), .Z(n15011) );
  NAND2_X1 U21302 ( .A1(n19588), .A2(n14561), .ZN(n3039) );
  XOR2_X1 U21318 ( .A1(n24019), .A2(n35630), .Z(n16321) );
  XOR2_X1 U21325 ( .A1(n24020), .A2(n23890), .Z(n35630) );
  XOR2_X1 U21326 ( .A1(n35631), .A2(n24022), .Z(n13504) );
  XOR2_X1 U21338 ( .A1(n24023), .A2(n20317), .Z(n35631) );
  NOR3_X2 U21340 ( .A1(n12927), .A2(n14769), .A3(n1354), .ZN(n3480) );
  XOR2_X1 U21354 ( .A1(n35636), .A2(n848), .Z(n36283) );
  XOR2_X1 U21365 ( .A1(n24011), .A2(n30150), .Z(n35640) );
  INV_X1 U21400 ( .I(n32103), .ZN(n17403) );
  XOR2_X1 U21401 ( .A1(n35642), .A2(n22279), .Z(n32103) );
  NAND3_X2 U21420 ( .A1(n585), .A2(n32507), .A3(n609), .ZN(n35647) );
  OAI22_X2 U21455 ( .A1(n22333), .A2(n20308), .B1(n20961), .B2(n937), .ZN(
        n12267) );
  OR2_X1 U21458 ( .A1(n33786), .A2(n35932), .Z(n8416) );
  NAND3_X2 U21466 ( .A1(n38653), .A2(n34190), .A3(n13485), .ZN(n13406) );
  OAI21_X1 U21480 ( .A1(n30042), .A2(n30043), .B(n5348), .ZN(n35653) );
  NAND2_X1 U21483 ( .A1(n27213), .A2(n16043), .ZN(n17152) );
  NOR2_X2 U21485 ( .A1(n8627), .A2(n11387), .ZN(n27213) );
  NAND2_X2 U21491 ( .A1(n36672), .A2(n16570), .ZN(n24417) );
  OAI22_X1 U21492 ( .A1(n35744), .A2(n13391), .B1(n1240), .B2(n26093), .ZN(
        n35655) );
  NAND3_X2 U21493 ( .A1(n13695), .A2(n13697), .A3(n13696), .ZN(n18875) );
  NOR2_X1 U21496 ( .A1(n29946), .A2(n29996), .ZN(n6600) );
  INV_X2 U21497 ( .I(n29994), .ZN(n29946) );
  XOR2_X1 U21501 ( .A1(n5129), .A2(n10829), .Z(n29994) );
  XOR2_X1 U21511 ( .A1(n343), .A2(n35656), .Z(n33695) );
  NAND3_X1 U21514 ( .A1(n1403), .A2(n37368), .A3(n39828), .ZN(n32762) );
  NOR2_X2 U21518 ( .A1(n36387), .A2(n20850), .ZN(n20849) );
  INV_X2 U21523 ( .I(n5348), .ZN(n29997) );
  XOR2_X1 U21543 ( .A1(n10722), .A2(n38813), .Z(n3317) );
  AND2_X1 U21545 ( .A1(n36833), .A2(n27357), .Z(n21170) );
  XOR2_X1 U21555 ( .A1(n4440), .A2(n22530), .Z(n13514) );
  XOR2_X1 U21563 ( .A1(n12015), .A2(n3239), .Z(n22530) );
  XOR2_X1 U21580 ( .A1(n14346), .A2(n26163), .Z(n26401) );
  NAND2_X2 U21583 ( .A1(n8721), .A2(n8719), .ZN(n32366) );
  AND2_X1 U21589 ( .A1(n35667), .A2(n38282), .Z(n20651) );
  NOR2_X1 U21597 ( .A1(n21365), .A2(n21364), .ZN(n35668) );
  XOR2_X1 U21605 ( .A1(n5553), .A2(n34144), .Z(n16558) );
  XOR2_X1 U21610 ( .A1(n26498), .A2(n4875), .Z(n5553) );
  OAI21_X1 U21611 ( .A1(n10120), .A2(n21839), .B(n7278), .ZN(n3868) );
  OAI21_X2 U21619 ( .A1(n32415), .A2(n14520), .B(n20525), .ZN(n35673) );
  NAND3_X2 U21632 ( .A1(n35675), .A2(n11672), .A3(n8343), .ZN(n22604) );
  XOR2_X1 U21640 ( .A1(n19640), .A2(n19639), .Z(n20524) );
  XOR2_X1 U21653 ( .A1(n35676), .A2(n29394), .Z(Ciphertext[36]) );
  XOR2_X1 U21656 ( .A1(n33509), .A2(n29165), .Z(n29816) );
  NAND2_X2 U21658 ( .A1(n18191), .A2(n28122), .ZN(n29165) );
  NAND2_X1 U21659 ( .A1(n31997), .A2(n35677), .ZN(n32462) );
  XOR2_X1 U21670 ( .A1(n36384), .A2(n900), .Z(n35678) );
  XOR2_X1 U21681 ( .A1(n23886), .A2(n23808), .Z(n24060) );
  NAND2_X2 U21683 ( .A1(n17443), .A2(n17442), .ZN(n23886) );
  INV_X4 U21689 ( .I(n35686), .ZN(n6977) );
  NAND3_X2 U21692 ( .A1(n5408), .A2(n36271), .A3(n33581), .ZN(n6014) );
  INV_X2 U21717 ( .I(n35687), .ZN(n23165) );
  NAND2_X2 U21737 ( .A1(n13631), .A2(n21926), .ZN(n18595) );
  XOR2_X1 U21738 ( .A1(n26253), .A2(n26252), .Z(n26348) );
  NAND2_X2 U21742 ( .A1(n11625), .A2(n11623), .ZN(n26252) );
  AOI22_X2 U21745 ( .A1(n12680), .A2(n36716), .B1(n5063), .B2(n12681), .ZN(
        n35688) );
  XOR2_X1 U21746 ( .A1(n38021), .A2(n1620), .Z(n12026) );
  INV_X2 U21749 ( .I(n37092), .ZN(n35689) );
  OAI22_X1 U21759 ( .A1(n14662), .A2(n33712), .B1(n18238), .B2(n1606), .ZN(
        n23909) );
  INV_X2 U21793 ( .I(n35693), .ZN(n24855) );
  NAND2_X2 U21799 ( .A1(n15549), .A2(n15550), .ZN(n35895) );
  NAND2_X2 U21806 ( .A1(n28038), .A2(n28039), .ZN(n28484) );
  NAND2_X2 U21811 ( .A1(n13618), .A2(n13621), .ZN(n16067) );
  AOI21_X2 U21812 ( .A1(n35699), .A2(n19856), .B(n20832), .ZN(n20831) );
  NAND2_X2 U21820 ( .A1(n22856), .A2(n19945), .ZN(n17917) );
  XOR2_X1 U21823 ( .A1(n13235), .A2(n22466), .Z(n2200) );
  NAND2_X2 U21832 ( .A1(n4703), .A2(n13629), .ZN(n16897) );
  XOR2_X1 U21836 ( .A1(n18991), .A2(n8183), .Z(n24972) );
  NAND2_X1 U21843 ( .A1(n12119), .A2(n12118), .ZN(n33180) );
  NOR2_X1 U21844 ( .A1(n22222), .A2(n22221), .ZN(n15499) );
  XOR2_X1 U21853 ( .A1(n4201), .A2(n1077), .Z(n10396) );
  INV_X1 U21860 ( .I(n29017), .ZN(n35702) );
  NOR2_X2 U21879 ( .A1(n22223), .A2(n22221), .ZN(n22135) );
  NOR2_X2 U21881 ( .A1(n21686), .A2(n21685), .ZN(n22223) );
  XOR2_X1 U21882 ( .A1(n19096), .A2(n11950), .Z(n10215) );
  OAI21_X2 U21885 ( .A1(n30422), .A2(n31698), .B(n15208), .ZN(n19096) );
  XOR2_X1 U21891 ( .A1(n26263), .A2(n35704), .Z(n10854) );
  XOR2_X1 U21894 ( .A1(n26223), .A2(n343), .Z(n35704) );
  AOI21_X1 U21895 ( .A1(n4621), .A2(n9913), .B(n1396), .ZN(n6321) );
  XOR2_X1 U21896 ( .A1(n1929), .A2(n794), .Z(n16459) );
  OR2_X1 U21899 ( .A1(n35732), .A2(n9178), .Z(n10795) );
  XOR2_X1 U21900 ( .A1(n35706), .A2(n3422), .Z(n3973) );
  XOR2_X1 U21901 ( .A1(n31627), .A2(n36999), .Z(n35706) );
  XOR2_X1 U21905 ( .A1(n16378), .A2(n16380), .Z(n16388) );
  INV_X4 U21907 ( .I(n32829), .ZN(n21248) );
  INV_X2 U21921 ( .I(n35708), .ZN(n21036) );
  NOR2_X1 U21924 ( .A1(n29477), .A2(n7303), .ZN(n2449) );
  XOR2_X1 U21931 ( .A1(n35852), .A2(n27659), .Z(n36136) );
  OR2_X1 U21936 ( .A1(n17607), .A2(n2616), .Z(n24798) );
  XOR2_X1 U21943 ( .A1(n22566), .A2(n35824), .Z(n18359) );
  NAND2_X2 U21945 ( .A1(n9127), .A2(n9126), .ZN(n22566) );
  XOR2_X1 U21959 ( .A1(n15935), .A2(n32610), .Z(n15933) );
  NAND2_X2 U21970 ( .A1(n495), .A2(n1487), .ZN(n16520) );
  NAND2_X2 U21972 ( .A1(n35718), .A2(n16517), .ZN(n27607) );
  XOR2_X1 U21978 ( .A1(n4441), .A2(n22517), .Z(n4440) );
  NAND2_X2 U21981 ( .A1(n1839), .A2(n1837), .ZN(n22517) );
  OAI22_X2 U21995 ( .A1(n1265), .A2(n35893), .B1(n24737), .B2(n5871), .ZN(
        n24736) );
  NAND2_X2 U21999 ( .A1(n7845), .A2(n32699), .ZN(n25080) );
  NOR2_X2 U22003 ( .A1(n35723), .A2(n18979), .ZN(n36425) );
  INV_X1 U22006 ( .I(n25488), .ZN(n220) );
  INV_X2 U22011 ( .I(n35724), .ZN(n217) );
  AOI21_X2 U22013 ( .A1(n1399), .A2(n30220), .B(n30159), .ZN(n10568) );
  XOR2_X1 U22014 ( .A1(n35726), .A2(n15331), .Z(n19938) );
  XOR2_X1 U22015 ( .A1(n411), .A2(n19014), .Z(n35726) );
  NAND2_X1 U22042 ( .A1(n17364), .A2(n29567), .ZN(n35731) );
  NAND2_X2 U22050 ( .A1(n106), .A2(n4138), .ZN(n35732) );
  NAND3_X1 U22054 ( .A1(n35911), .A2(n32575), .A3(n2191), .ZN(n21188) );
  INV_X2 U22055 ( .I(n14213), .ZN(n15936) );
  NOR2_X2 U22057 ( .A1(n16841), .A2(n24416), .ZN(n14213) );
  XOR2_X1 U22058 ( .A1(n27833), .A2(n27731), .Z(n17043) );
  XOR2_X1 U22060 ( .A1(n25194), .A2(n25275), .Z(n25103) );
  NAND2_X2 U22061 ( .A1(n9999), .A2(n4608), .ZN(n25275) );
  AOI21_X2 U22066 ( .A1(n22018), .A2(n22017), .B(n35734), .ZN(n22430) );
  OAI21_X2 U22077 ( .A1(n2190), .A2(n14945), .B(n33186), .ZN(n35780) );
  XOR2_X1 U22099 ( .A1(n28865), .A2(n29252), .Z(n28979) );
  NOR2_X2 U22103 ( .A1(n6046), .A2(n35737), .ZN(n36700) );
  XOR2_X1 U22118 ( .A1(n25286), .A2(n34137), .Z(n35741) );
  XOR2_X1 U22123 ( .A1(n35743), .A2(n6927), .Z(n16339) );
  XOR2_X1 U22126 ( .A1(n27714), .A2(n27805), .Z(n35743) );
  INV_X4 U22127 ( .I(n17499), .ZN(n1340) );
  XOR2_X1 U22129 ( .A1(n22458), .A2(n9115), .Z(n8172) );
  XOR2_X1 U22130 ( .A1(n22443), .A2(n8026), .Z(n22458) );
  NOR2_X1 U22132 ( .A1(n15209), .A2(n35179), .ZN(n17364) );
  BUF_X2 U22135 ( .I(n33258), .Z(n35744) );
  OAI21_X2 U22147 ( .A1(n16373), .A2(n12533), .B(n16372), .ZN(n18407) );
  XOR2_X1 U22151 ( .A1(n38514), .A2(n36765), .Z(n35747) );
  INV_X1 U22159 ( .I(n35748), .ZN(n25408) );
  XOR2_X1 U22181 ( .A1(n27546), .A2(n19808), .Z(n5252) );
  XOR2_X1 U22187 ( .A1(n476), .A2(n5116), .Z(n35752) );
  XOR2_X1 U22194 ( .A1(n32839), .A2(n34151), .Z(n36858) );
  NOR2_X1 U22199 ( .A1(n35756), .A2(n35755), .ZN(n30878) );
  INV_X2 U22207 ( .I(n13519), .ZN(n35755) );
  NAND2_X1 U22209 ( .A1(n1335), .A2(n22307), .ZN(n35756) );
  INV_X2 U22210 ( .I(n35757), .ZN(n15248) );
  XOR2_X1 U22216 ( .A1(n35758), .A2(n26171), .Z(n26689) );
  XOR2_X1 U22219 ( .A1(n26173), .A2(n36270), .Z(n35758) );
  XOR2_X1 U22235 ( .A1(n1323), .A2(n35211), .Z(n35760) );
  INV_X2 U22244 ( .I(n35228), .ZN(n27364) );
  NOR2_X1 U22252 ( .A1(n859), .A2(n26936), .ZN(n11339) );
  OAI21_X2 U22255 ( .A1(n9951), .A2(n4833), .B(n306), .ZN(n28417) );
  NOR2_X2 U22257 ( .A1(n5908), .A2(n35333), .ZN(n25920) );
  NAND2_X1 U22262 ( .A1(n35764), .A2(n35259), .ZN(n6246) );
  XOR2_X1 U22264 ( .A1(n9408), .A2(n9409), .Z(n740) );
  XOR2_X1 U22271 ( .A1(n35765), .A2(n34038), .Z(n63) );
  XOR2_X1 U22272 ( .A1(n29094), .A2(n31811), .Z(n35765) );
  XNOR2_X1 U22273 ( .A1(n18813), .A2(n11722), .ZN(n36127) );
  XOR2_X1 U22275 ( .A1(n2269), .A2(n29122), .Z(n11722) );
  NOR2_X2 U22280 ( .A1(n31453), .A2(n18590), .ZN(n18241) );
  INV_X2 U22290 ( .I(n35769), .ZN(n730) );
  OAI22_X2 U22326 ( .A1(n11610), .A2(n5224), .B1(n5223), .B2(n20038), .ZN(
        n20707) );
  NAND2_X1 U22346 ( .A1(n28266), .A2(n38996), .ZN(n36059) );
  NAND2_X2 U22352 ( .A1(n10254), .A2(n28124), .ZN(n27963) );
  AND2_X1 U22357 ( .A1(n14075), .A2(n31899), .Z(n14073) );
  NOR2_X2 U22360 ( .A1(n6850), .A2(n5599), .ZN(n35779) );
  XOR2_X1 U22367 ( .A1(n25037), .A2(n9695), .Z(n24838) );
  XOR2_X1 U22380 ( .A1(n27809), .A2(n27529), .Z(n27530) );
  NAND2_X2 U22382 ( .A1(n11581), .A2(n35786), .ZN(n17179) );
  NAND2_X2 U22385 ( .A1(n17673), .A2(n36587), .ZN(n19608) );
  NAND2_X2 U22388 ( .A1(n31580), .A2(n12825), .ZN(n25478) );
  OAI22_X2 U22402 ( .A1(n15215), .A2(n34583), .B1(n20924), .B2(n541), .ZN(
        n5597) );
  INV_X2 U22403 ( .I(n15261), .ZN(n541) );
  NAND2_X2 U22408 ( .A1(n33535), .A2(n14669), .ZN(n35855) );
  XOR2_X1 U22417 ( .A1(n7659), .A2(n19839), .Z(n6363) );
  NOR2_X2 U22420 ( .A1(n8503), .A2(n8504), .ZN(n7659) );
  NOR2_X1 U22430 ( .A1(n38202), .A2(n36838), .ZN(n15695) );
  NOR2_X1 U22433 ( .A1(n17194), .A2(n13371), .ZN(n9366) );
  OAI21_X2 U22445 ( .A1(n6503), .A2(n26471), .B(n35794), .ZN(n7757) );
  XOR2_X1 U22449 ( .A1(n33498), .A2(n31020), .Z(n1825) );
  OAI21_X2 U22456 ( .A1(n23376), .A2(n23377), .B(n23375), .ZN(n33452) );
  NAND2_X2 U22460 ( .A1(n36866), .A2(n21212), .ZN(n16771) );
  NOR2_X2 U22465 ( .A1(n35795), .A2(n8257), .ZN(n27523) );
  XOR2_X1 U22485 ( .A1(n35796), .A2(n26374), .Z(n12012) );
  NAND2_X2 U22499 ( .A1(n6332), .A2(n29644), .ZN(n10868) );
  NAND2_X2 U22504 ( .A1(n29443), .A2(n10870), .ZN(n6332) );
  AOI21_X2 U22533 ( .A1(n21306), .A2(n25771), .B(n21305), .ZN(n10965) );
  AND2_X1 U22534 ( .A1(n9833), .A2(n25758), .Z(n16890) );
  XOR2_X1 U22536 ( .A1(n25215), .A2(n30973), .Z(n36259) );
  NAND2_X2 U22549 ( .A1(n3192), .A2(n36832), .ZN(n28729) );
  NAND2_X2 U22551 ( .A1(n14754), .A2(n21988), .ZN(n22476) );
  NOR2_X1 U22553 ( .A1(n3293), .A2(n21894), .ZN(n21515) );
  NAND2_X2 U22560 ( .A1(n35803), .A2(n13548), .ZN(n17087) );
  XOR2_X1 U22576 ( .A1(n26387), .A2(n26388), .Z(n26474) );
  XNOR2_X1 U22590 ( .A1(n5730), .A2(n25246), .ZN(n36339) );
  XOR2_X1 U22605 ( .A1(n35810), .A2(n22672), .Z(n36291) );
  XOR2_X1 U22607 ( .A1(n22582), .A2(n36290), .Z(n22672) );
  OAI21_X2 U22625 ( .A1(n13825), .A2(n13824), .B(n28682), .ZN(n13823) );
  INV_X2 U22628 ( .I(n35816), .ZN(n37043) );
  XOR2_X1 U22633 ( .A1(n30898), .A2(n784), .Z(n35816) );
  AOI22_X2 U22640 ( .A1(n35818), .A2(n34015), .B1(n8574), .B2(n21969), .ZN(
        n2193) );
  OAI21_X2 U22643 ( .A1(n21586), .A2(n119), .B(n21584), .ZN(n9876) );
  NAND2_X2 U22659 ( .A1(n21128), .A2(n36876), .ZN(n23900) );
  XOR2_X1 U22660 ( .A1(n33470), .A2(n990), .Z(n31138) );
  XOR2_X1 U22667 ( .A1(n22592), .A2(n22514), .Z(n20609) );
  NAND2_X1 U22670 ( .A1(n22317), .A2(n36745), .ZN(n7093) );
  AOI21_X2 U22678 ( .A1(n28370), .A2(n28580), .B(n16038), .ZN(n35823) );
  OR2_X1 U22684 ( .A1(n19477), .A2(n8798), .Z(n35825) );
  NAND2_X2 U22692 ( .A1(n35833), .A2(n36464), .ZN(n22282) );
  NAND3_X2 U22703 ( .A1(n33340), .A2(n33369), .A3(n12022), .ZN(n35826) );
  BUF_X2 U22716 ( .I(n35867), .Z(n35832) );
  XOR2_X1 U22718 ( .A1(n17890), .A2(n19758), .Z(n7763) );
  XOR2_X1 U22729 ( .A1(n35834), .A2(n10863), .Z(n11048) );
  INV_X2 U22732 ( .I(n35835), .ZN(n12101) );
  OAI22_X1 U22734 ( .A1(n13133), .A2(n13151), .B1(n35224), .B2(n14193), .ZN(
        n31350) );
  XOR2_X1 U22739 ( .A1(n35836), .A2(n12858), .Z(n12856) );
  XOR2_X1 U22741 ( .A1(n7250), .A2(n7247), .Z(n8199) );
  NAND2_X1 U22751 ( .A1(n307), .A2(n35837), .ZN(n19784) );
  AOI22_X1 U22753 ( .A1(n12369), .A2(n18873), .B1(n7303), .B2(n12148), .ZN(
        n35837) );
  XOR2_X1 U22754 ( .A1(n23948), .A2(n23949), .Z(n17790) );
  XOR2_X1 U22763 ( .A1(n7582), .A2(n34020), .Z(n36756) );
  OAI22_X2 U22779 ( .A1(n35841), .A2(n35840), .B1(n9362), .B2(n24290), .ZN(
        n24707) );
  AOI21_X2 U22783 ( .A1(n37118), .A2(n6668), .B(n35843), .ZN(n6875) );
  NOR3_X1 U22784 ( .A1(n5772), .A2(n35228), .A3(n34001), .ZN(n35843) );
  NAND2_X2 U22785 ( .A1(n35844), .A2(n1437), .ZN(n11006) );
  NOR2_X1 U22791 ( .A1(n27895), .A2(n1445), .ZN(n5470) );
  INV_X2 U22793 ( .I(n17755), .ZN(n27895) );
  INV_X1 U22823 ( .I(n35847), .ZN(n35846) );
  NAND2_X1 U22824 ( .A1(n39488), .A2(n28238), .ZN(n35847) );
  XOR2_X1 U22825 ( .A1(n22528), .A2(n35848), .Z(n494) );
  NAND2_X2 U22827 ( .A1(n21831), .A2(n21832), .ZN(n22528) );
  OAI21_X2 U22833 ( .A1(n36607), .A2(n35849), .B(n30163), .ZN(n30173) );
  XOR2_X1 U22847 ( .A1(n21036), .A2(n35853), .Z(n35852) );
  OR2_X1 U22850 ( .A1(n15218), .A2(n6581), .Z(n6827) );
  AOI21_X2 U22854 ( .A1(n3798), .A2(n3799), .B(n33519), .ZN(n35867) );
  XOR2_X1 U22855 ( .A1(n35856), .A2(n24942), .Z(n8277) );
  XOR2_X1 U22856 ( .A1(n25284), .A2(n19683), .Z(n35856) );
  XOR2_X1 U22859 ( .A1(n35857), .A2(n2031), .Z(n20866) );
  INV_X2 U22861 ( .I(n9900), .ZN(n3602) );
  XOR2_X1 U22862 ( .A1(n32959), .A2(n437), .Z(n9900) );
  XOR2_X1 U22864 ( .A1(n20485), .A2(n15471), .Z(n20484) );
  BUF_X2 U22865 ( .I(n29699), .Z(n35858) );
  NAND3_X2 U22873 ( .A1(n16195), .A2(n18460), .A3(n24748), .ZN(n25182) );
  XOR2_X1 U22874 ( .A1(n11312), .A2(n11309), .Z(n35859) );
  OAI22_X2 U22876 ( .A1(n3618), .A2(n1990), .B1(n18699), .B2(n20266), .ZN(
        n35860) );
  NOR2_X2 U22894 ( .A1(n1028), .A2(n18110), .ZN(n30421) );
  NAND2_X2 U22897 ( .A1(n16473), .A2(n17338), .ZN(n29034) );
  XOR2_X1 U22914 ( .A1(n2284), .A2(n13551), .Z(n12732) );
  CLKBUF_X4 U22921 ( .I(n21938), .Z(n35883) );
  XOR2_X1 U22932 ( .A1(n11999), .A2(n11998), .Z(n861) );
  XOR2_X1 U22935 ( .A1(n10971), .A2(n10970), .Z(n7923) );
  NAND2_X1 U22948 ( .A1(n2449), .A2(n18873), .ZN(n2448) );
  NAND3_X2 U22953 ( .A1(n9256), .A2(n10773), .A3(n19560), .ZN(n25149) );
  OR2_X1 U22962 ( .A1(n7303), .A2(n34534), .Z(n29480) );
  XOR2_X1 U22968 ( .A1(n22503), .A2(n21999), .Z(n22002) );
  NAND3_X2 U22982 ( .A1(n20751), .A2(n20750), .A3(n21612), .ZN(n19373) );
  NOR2_X1 U22991 ( .A1(n13927), .A2(n17378), .ZN(n27995) );
  XOR2_X1 U22993 ( .A1(n31777), .A2(n18060), .Z(n13927) );
  INV_X2 U22996 ( .I(n35868), .ZN(n20449) );
  NAND2_X2 U23004 ( .A1(n27988), .A2(n27987), .ZN(n28661) );
  OR2_X1 U23008 ( .A1(n12049), .A2(n36117), .Z(n32945) );
  XOR2_X1 U23023 ( .A1(n12231), .A2(n28987), .Z(n12215) );
  XOR2_X1 U23024 ( .A1(n35871), .A2(n2159), .Z(n5966) );
  XOR2_X1 U23026 ( .A1(n35908), .A2(n8540), .Z(n14217) );
  XOR2_X1 U23040 ( .A1(n8654), .A2(n35874), .Z(n4315) );
  XOR2_X1 U23043 ( .A1(n28851), .A2(n31524), .Z(n35874) );
  OAI22_X2 U23051 ( .A1(n16288), .A2(n14769), .B1(n16287), .B2(n12927), .ZN(
        n36214) );
  NAND2_X2 U23069 ( .A1(n26067), .A2(n26066), .ZN(n7602) );
  NAND3_X2 U23075 ( .A1(n15614), .A2(n17219), .A3(n15613), .ZN(n17440) );
  NAND2_X2 U23077 ( .A1(n1048), .A2(n22184), .ZN(n17793) );
  NAND2_X2 U23078 ( .A1(n23522), .A2(n2273), .ZN(n23525) );
  XOR2_X1 U23087 ( .A1(n22723), .A2(n35879), .Z(n35878) );
  NOR2_X2 U23095 ( .A1(n11646), .A2(n9481), .ZN(n35882) );
  AND2_X1 U23098 ( .A1(n4880), .A2(n34786), .Z(n30944) );
  NAND2_X2 U23103 ( .A1(n17499), .A2(n22307), .ZN(n36069) );
  XOR2_X1 U23104 ( .A1(n22787), .A2(n22672), .Z(n17277) );
  OR2_X1 U23106 ( .A1(n730), .A2(n8069), .Z(n8771) );
  NAND2_X2 U23112 ( .A1(n23065), .A2(n23064), .ZN(n23250) );
  NAND2_X2 U23117 ( .A1(n6213), .A2(n4760), .ZN(n23399) );
  NAND2_X2 U23118 ( .A1(n35886), .A2(n15001), .ZN(n25163) );
  BUF_X2 U23119 ( .I(n1254), .Z(n35887) );
  XNOR2_X1 U23131 ( .A1(n22622), .A2(n29223), .ZN(n36605) );
  XOR2_X1 U23140 ( .A1(n35889), .A2(n38226), .Z(n184) );
  AOI22_X2 U23146 ( .A1(n11878), .A2(n33489), .B1(n12169), .B2(n22367), .ZN(
        n13704) );
  OR2_X1 U23159 ( .A1(n20077), .A2(n15290), .Z(n22783) );
  NAND2_X2 U23160 ( .A1(n17132), .A2(n12327), .ZN(n27398) );
  NAND2_X2 U23163 ( .A1(n7010), .A2(n22730), .ZN(n23637) );
  XOR2_X1 U23190 ( .A1(n35996), .A2(n35894), .Z(n14672) );
  XNOR2_X1 U23191 ( .A1(n18807), .A2(n18279), .ZN(n35970) );
  NAND2_X1 U23197 ( .A1(n8495), .A2(n16039), .ZN(n15115) );
  XOR2_X1 U23199 ( .A1(n11901), .A2(Key[169]), .Z(n16039) );
  NAND2_X2 U23200 ( .A1(n32796), .A2(n13042), .ZN(n22838) );
  INV_X2 U23220 ( .I(n35896), .ZN(n17594) );
  OR2_X1 U23223 ( .A1(n7742), .A2(n26249), .Z(n2226) );
  AND2_X1 U23228 ( .A1(n30284), .A2(n14962), .Z(n36929) );
  BUF_X2 U23241 ( .I(n27283), .Z(n35904) );
  AOI21_X2 U23248 ( .A1(n27107), .A2(n28052), .B(n27962), .ZN(n36029) );
  NAND2_X1 U23250 ( .A1(n15224), .A2(n36791), .ZN(n28733) );
  AND2_X1 U23275 ( .A1(n30153), .A2(n20525), .Z(n8717) );
  XOR2_X1 U23278 ( .A1(n14425), .A2(n35909), .Z(n5002) );
  XOR2_X1 U23279 ( .A1(n15625), .A2(n29003), .Z(n35909) );
  XOR2_X1 U23280 ( .A1(n19047), .A2(n35910), .Z(n30221) );
  XOR2_X1 U23296 ( .A1(n17159), .A2(n28985), .Z(n35910) );
  XOR2_X1 U23297 ( .A1(n38171), .A2(n1553), .Z(n25141) );
  INV_X2 U23300 ( .I(n38629), .ZN(n35911) );
  NAND2_X2 U23305 ( .A1(n14910), .A2(n14908), .ZN(n20643) );
  NAND2_X1 U23308 ( .A1(n17538), .A2(n17617), .ZN(n17616) );
  XOR2_X1 U23332 ( .A1(n26393), .A2(n26466), .Z(n13244) );
  AOI21_X2 U23348 ( .A1(n33849), .A2(n4686), .B(n31678), .ZN(n27045) );
  XOR2_X1 U23354 ( .A1(n25268), .A2(n25162), .Z(n10407) );
  XOR2_X1 U23355 ( .A1(n13917), .A2(n25096), .Z(n25162) );
  INV_X2 U23361 ( .I(n31107), .ZN(n3662) );
  NAND2_X1 U23365 ( .A1(n5988), .A2(n31107), .ZN(n28235) );
  INV_X2 U23389 ( .I(n11970), .ZN(n32017) );
  AOI21_X2 U23404 ( .A1(n8328), .A2(n18150), .B(n8325), .ZN(n28398) );
  XOR2_X1 U23428 ( .A1(n35923), .A2(n17759), .Z(n26906) );
  NAND2_X2 U23435 ( .A1(n1039), .A2(n30574), .ZN(n23039) );
  OAI21_X2 U23436 ( .A1(n33240), .A2(n2192), .B(n35924), .ZN(n14896) );
  NAND2_X2 U23440 ( .A1(n2518), .A2(n576), .ZN(n27637) );
  AOI22_X2 U23459 ( .A1(n20827), .A2(n15031), .B1(n33285), .B2(n18005), .ZN(
        n35926) );
  NAND3_X2 U23479 ( .A1(n7483), .A2(n28154), .A3(n17818), .ZN(n11296) );
  NAND2_X2 U23490 ( .A1(n35928), .A2(n18378), .ZN(n496) );
  OAI21_X2 U23493 ( .A1(n18379), .A2(n18380), .B(n27571), .ZN(n35928) );
  NOR2_X1 U23495 ( .A1(n5537), .A2(n26852), .ZN(n19207) );
  NOR2_X1 U23500 ( .A1(n5537), .A2(n20660), .ZN(n11674) );
  XOR2_X1 U23519 ( .A1(n25242), .A2(n25229), .Z(n25313) );
  NAND3_X2 U23549 ( .A1(n32182), .A2(n9663), .A3(n18150), .ZN(n9575) );
  NAND2_X2 U23566 ( .A1(n16235), .A2(n16488), .ZN(n23939) );
  XOR2_X1 U23567 ( .A1(n35941), .A2(n20486), .Z(n15471) );
  XOR2_X1 U23569 ( .A1(n37701), .A2(n35942), .Z(n35941) );
  INV_X2 U23577 ( .I(n11937), .ZN(n35942) );
  OAI21_X1 U23591 ( .A1(n20623), .A2(n7357), .B(n35943), .ZN(n20148) );
  BUF_X2 U23600 ( .I(n26039), .Z(n35944) );
  XOR2_X1 U23623 ( .A1(n25841), .A2(n30469), .Z(n857) );
  NOR2_X1 U23624 ( .A1(n11678), .A2(n23391), .ZN(n4859) );
  NAND2_X2 U23627 ( .A1(n21634), .A2(n21633), .ZN(n36397) );
  XOR2_X1 U23659 ( .A1(n13550), .A2(n36390), .Z(n36150) );
  XOR2_X1 U23676 ( .A1(n20846), .A2(n20772), .Z(n6049) );
  NAND2_X2 U23697 ( .A1(n25659), .A2(n25658), .ZN(n32095) );
  OAI22_X2 U23698 ( .A1(n22314), .A2(n15004), .B1(n18675), .B2(n18674), .ZN(
        n18087) );
  XOR2_X1 U23699 ( .A1(n2042), .A2(n35957), .Z(n36357) );
  INV_X2 U23729 ( .I(n2880), .ZN(n15388) );
  XOR2_X1 U23739 ( .A1(n3023), .A2(n3022), .Z(n2880) );
  NAND2_X2 U23741 ( .A1(n8070), .A2(n2148), .ZN(n35962) );
  XOR2_X1 U23745 ( .A1(n35964), .A2(n28630), .Z(n28631) );
  XOR2_X1 U23748 ( .A1(n29052), .A2(n19825), .Z(n35964) );
  NOR3_X1 U23762 ( .A1(n35966), .A2(n35965), .A3(n1406), .ZN(n21196) );
  NOR2_X1 U23763 ( .A1(n29310), .A2(n29384), .ZN(n35965) );
  XOR2_X1 U23770 ( .A1(n32135), .A2(n34345), .Z(n22747) );
  NAND2_X2 U23781 ( .A1(n37098), .A2(n19179), .ZN(n26760) );
  NOR2_X1 U23786 ( .A1(n14235), .A2(n35915), .ZN(n10839) );
  NAND2_X2 U23790 ( .A1(n13641), .A2(n13640), .ZN(n14235) );
  XOR2_X1 U23798 ( .A1(n35970), .A2(n23649), .Z(n35969) );
  NOR2_X2 U23803 ( .A1(n23942), .A2(n23941), .ZN(n11081) );
  XOR2_X1 U23805 ( .A1(n5629), .A2(n35971), .Z(n734) );
  XOR2_X1 U23808 ( .A1(n36128), .A2(n25025), .Z(n35971) );
  AOI21_X2 U23814 ( .A1(n35976), .A2(n35975), .B(n7191), .ZN(n18240) );
  NAND2_X1 U23817 ( .A1(n7193), .A2(n7194), .ZN(n35976) );
  BUF_X2 U23818 ( .I(n21111), .Z(n35977) );
  NAND3_X1 U23833 ( .A1(n27411), .A2(n27311), .A3(n997), .ZN(n35978) );
  XOR2_X1 U23854 ( .A1(n4646), .A2(n35983), .Z(n12431) );
  XOR2_X1 U23859 ( .A1(n37129), .A2(n35984), .Z(n35983) );
  INV_X1 U23861 ( .I(n30122), .ZN(n35984) );
  NAND2_X2 U23879 ( .A1(n7805), .A2(n7808), .ZN(n8402) );
  XOR2_X1 U23925 ( .A1(n35993), .A2(n33357), .Z(n384) );
  XOR2_X1 U23927 ( .A1(n26545), .A2(n744), .Z(n35993) );
  NOR2_X2 U23930 ( .A1(n20670), .A2(n22153), .ZN(n20335) );
  INV_X2 U23931 ( .I(n37643), .ZN(n16686) );
  NAND2_X2 U23933 ( .A1(n15502), .A2(n11671), .ZN(n30881) );
  INV_X1 U23935 ( .I(n36815), .ZN(n30436) );
  AND2_X1 U23938 ( .A1(n36815), .A2(n36658), .Z(n19215) );
  XOR2_X1 U23950 ( .A1(n11215), .A2(n19991), .Z(n9221) );
  NAND2_X2 U23955 ( .A1(n22062), .A2(n32886), .ZN(n32885) );
  NOR2_X2 U23986 ( .A1(n9803), .A2(n10775), .ZN(n26001) );
  XOR2_X1 U23987 ( .A1(n26450), .A2(n26451), .Z(n6681) );
  OR2_X1 U23996 ( .A1(n28389), .A2(n18960), .Z(n11911) );
  AOI22_X2 U23999 ( .A1(n22083), .A2(n23114), .B1(n23115), .B2(n8569), .ZN(
        n36001) );
  NOR2_X2 U24015 ( .A1(n36004), .A2(n8265), .ZN(n32002) );
  NOR2_X1 U24020 ( .A1(n2969), .A2(n36801), .ZN(n2967) );
  XOR2_X1 U24029 ( .A1(n26448), .A2(n37380), .Z(n659) );
  NAND2_X2 U24040 ( .A1(n20551), .A2(n12568), .ZN(n22645) );
  XOR2_X1 U24041 ( .A1(n36013), .A2(n19937), .Z(Ciphertext[164]) );
  NOR3_X1 U24055 ( .A1(n21248), .A2(n27508), .A3(n31287), .ZN(n27187) );
  INV_X4 U24060 ( .I(n36532), .ZN(n15677) );
  NAND2_X2 U24062 ( .A1(n5454), .A2(n5452), .ZN(n36532) );
  XOR2_X1 U24067 ( .A1(n19096), .A2(n2318), .Z(n2317) );
  OAI21_X2 U24074 ( .A1(n36020), .A2(n20105), .B(n911), .ZN(n18349) );
  INV_X2 U24119 ( .I(n36024), .ZN(n11060) );
  XOR2_X1 U24120 ( .A1(n11061), .A2(n11062), .Z(n36024) );
  XOR2_X1 U24124 ( .A1(n22543), .A2(n18751), .Z(n1947) );
  NOR2_X1 U24140 ( .A1(n17931), .A2(n23354), .ZN(n36026) );
  NAND3_X1 U24145 ( .A1(n31192), .A2(n2888), .A3(n3575), .ZN(n2889) );
  NOR2_X1 U24149 ( .A1(n36794), .A2(n24896), .ZN(n25584) );
  XOR2_X1 U24158 ( .A1(n36030), .A2(n36205), .Z(n14481) );
  XOR2_X1 U24159 ( .A1(n25265), .A2(n14672), .Z(n36030) );
  INV_X2 U24172 ( .I(n25283), .ZN(n30318) );
  NAND2_X2 U24177 ( .A1(n24546), .A2(n4694), .ZN(n25283) );
  NAND2_X1 U24180 ( .A1(n24146), .A2(n1602), .ZN(n8501) );
  NAND3_X2 U24206 ( .A1(n29767), .A2(n31059), .A3(n31517), .ZN(n29792) );
  NAND2_X2 U24208 ( .A1(n20028), .A2(n24439), .ZN(n36075) );
  XOR2_X1 U24211 ( .A1(n11753), .A2(n29528), .Z(n11207) );
  XOR2_X1 U24213 ( .A1(n36034), .A2(n5103), .Z(n14411) );
  OAI21_X2 U24215 ( .A1(n33380), .A2(n20870), .B(n36036), .ZN(n27781) );
  NAND2_X1 U24223 ( .A1(n21461), .A2(n21868), .ZN(n3564) );
  XOR2_X1 U24229 ( .A1(n2068), .A2(n2067), .Z(n2066) );
  XOR2_X1 U24238 ( .A1(n22592), .A2(n36038), .Z(n22596) );
  NAND2_X2 U24260 ( .A1(n32337), .A2(n11683), .ZN(n15871) );
  XOR2_X1 U24274 ( .A1(n32646), .A2(n36040), .Z(n2352) );
  NAND2_X1 U24277 ( .A1(n28807), .A2(n19759), .ZN(n28289) );
  XOR2_X1 U24280 ( .A1(n27598), .A2(n32686), .Z(n36041) );
  NAND2_X2 U24282 ( .A1(n5777), .A2(n5776), .ZN(n9824) );
  INV_X2 U24301 ( .I(n36044), .ZN(n1589) );
  XNOR2_X1 U24304 ( .A1(n36646), .A2(n2398), .ZN(n36044) );
  NOR2_X2 U24309 ( .A1(n36046), .A2(n4775), .ZN(n9999) );
  XOR2_X1 U24313 ( .A1(n33645), .A2(n29649), .Z(n17798) );
  NOR2_X1 U24325 ( .A1(n38609), .A2(n12235), .ZN(n18752) );
  XOR2_X1 U24335 ( .A1(n26208), .A2(n659), .Z(n12412) );
  OAI21_X1 U24364 ( .A1(n38156), .A2(n16889), .B(n36051), .ZN(n9559) );
  OAI21_X1 U24367 ( .A1(n1208), .A2(n39235), .B(n17770), .ZN(n9684) );
  NAND2_X2 U24374 ( .A1(n36053), .A2(n25339), .ZN(n26063) );
  OAI21_X1 U24385 ( .A1(n566), .A2(n33968), .B(n29719), .ZN(n16630) );
  NAND2_X2 U24389 ( .A1(n7251), .A2(n36935), .ZN(n28525) );
  XOR2_X1 U24398 ( .A1(n3110), .A2(n25182), .Z(n25312) );
  NOR2_X2 U24411 ( .A1(n21709), .A2(n36055), .ZN(n22092) );
  AOI21_X1 U24413 ( .A1(n21706), .A2(n21707), .B(n2045), .ZN(n36055) );
  NOR2_X1 U24416 ( .A1(n5709), .A2(n11622), .ZN(n30377) );
  XOR2_X1 U24429 ( .A1(n2935), .A2(n22453), .Z(n36057) );
  OR2_X1 U24434 ( .A1(n29756), .A2(n29754), .Z(n33607) );
  XOR2_X1 U24443 ( .A1(Plaintext[145]), .A2(Key[145]), .Z(n36062) );
  NAND2_X2 U24445 ( .A1(n15868), .A2(n17869), .ZN(n17335) );
  INV_X2 U24449 ( .I(n36063), .ZN(n7240) );
  INV_X2 U24450 ( .I(n36064), .ZN(n32775) );
  XOR2_X1 U24466 ( .A1(n26279), .A2(n19808), .Z(n13931) );
  BUF_X2 U24467 ( .I(n23899), .Z(n36065) );
  XOR2_X1 U24470 ( .A1(n36066), .A2(n6764), .Z(n24285) );
  XOR2_X1 U24483 ( .A1(n22597), .A2(n33177), .Z(n12863) );
  XOR2_X1 U24486 ( .A1(n36068), .A2(n24016), .Z(n3454) );
  XOR2_X1 U24492 ( .A1(n23667), .A2(n11739), .Z(n24016) );
  AOI21_X1 U24499 ( .A1(n36069), .A2(n1335), .B(n17989), .ZN(n4126) );
  XOR2_X1 U24509 ( .A1(n22574), .A2(n6047), .Z(n30661) );
  AOI21_X2 U24552 ( .A1(n4384), .A2(n1547), .B(n36133), .ZN(n36071) );
  OAI21_X2 U24557 ( .A1(n4456), .A2(n27946), .B(n36072), .ZN(n28651) );
  XOR2_X1 U24564 ( .A1(n36074), .A2(n873), .Z(n9373) );
  XOR2_X1 U24566 ( .A1(n27605), .A2(n32021), .Z(n36074) );
  BUF_X2 U24584 ( .I(n10907), .Z(n36076) );
  XOR2_X1 U24586 ( .A1(n36077), .A2(n6963), .Z(n26177) );
  XOR2_X1 U24587 ( .A1(n26554), .A2(n26245), .Z(n26488) );
  NAND2_X2 U24591 ( .A1(n4431), .A2(n4430), .ZN(n26245) );
  XOR2_X1 U24599 ( .A1(n26161), .A2(n29269), .Z(n9932) );
  NAND2_X2 U24618 ( .A1(n3013), .A2(n25799), .ZN(n3434) );
  XOR2_X1 U24619 ( .A1(n23997), .A2(n36079), .Z(n19960) );
  OAI22_X2 U24624 ( .A1(n36080), .A2(n1220), .B1(n2998), .B2(n10946), .ZN(
        n12341) );
  XOR2_X1 U24625 ( .A1(n36970), .A2(n36081), .Z(n33479) );
  XOR2_X1 U24627 ( .A1(n17363), .A2(n8780), .Z(n36081) );
  XOR2_X1 U24634 ( .A1(n15592), .A2(n19797), .Z(n1886) );
  XOR2_X1 U24635 ( .A1(n22670), .A2(n36290), .Z(n20412) );
  NAND2_X2 U24640 ( .A1(n21263), .A2(n21260), .ZN(n36290) );
  INV_X2 U24646 ( .I(n6947), .ZN(n22326) );
  OAI22_X2 U24656 ( .A1(n439), .A2(n440), .B1(n13557), .B2(n13556), .ZN(n6947)
         );
  INV_X4 U24657 ( .I(n7221), .ZN(n8082) );
  NAND2_X2 U24663 ( .A1(n6243), .A2(n6244), .ZN(n7221) );
  XOR2_X1 U24669 ( .A1(n23804), .A2(n6289), .Z(n36087) );
  NAND2_X2 U24700 ( .A1(n22059), .A2(n22100), .ZN(n36092) );
  NAND2_X2 U24708 ( .A1(n12542), .A2(n28492), .ZN(n29252) );
  AOI22_X2 U24720 ( .A1(n9726), .A2(n6775), .B1(n1475), .B2(n27130), .ZN(
        n27632) );
  NAND2_X1 U24729 ( .A1(n2339), .A2(n8155), .ZN(n36097) );
  NAND2_X1 U24737 ( .A1(n19285), .A2(n4748), .ZN(n36098) );
  NAND2_X1 U24741 ( .A1(n36099), .A2(n2678), .ZN(n33517) );
  INV_X2 U24752 ( .I(n36104), .ZN(n30317) );
  XOR2_X1 U24764 ( .A1(n26279), .A2(n26404), .Z(n15530) );
  NAND2_X2 U24766 ( .A1(n15870), .A2(n15869), .ZN(n26404) );
  NOR2_X2 U24775 ( .A1(n6421), .A2(n6684), .ZN(n3309) );
  INV_X2 U24778 ( .I(n23310), .ZN(n6421) );
  NAND2_X2 U24786 ( .A1(n36444), .A2(n2088), .ZN(n7693) );
  NAND3_X2 U24802 ( .A1(n2587), .A2(n2586), .A3(n14597), .ZN(n15346) );
  NAND2_X2 U24803 ( .A1(n36109), .A2(n36108), .ZN(n17732) );
  INV_X1 U24806 ( .I(n36775), .ZN(n36108) );
  XOR2_X1 U24810 ( .A1(n9762), .A2(n36111), .Z(n10655) );
  XOR2_X1 U24811 ( .A1(n16082), .A2(n34161), .Z(n36111) );
  INV_X2 U24824 ( .I(n36113), .ZN(n2597) );
  XOR2_X1 U24833 ( .A1(n27837), .A2(n13878), .Z(n36114) );
  OAI22_X2 U24835 ( .A1(n33206), .A2(n33394), .B1(n37083), .B2(n30196), .ZN(
        n32925) );
  INV_X2 U24847 ( .I(n36117), .ZN(n37060) );
  XOR2_X1 U24848 ( .A1(n6852), .A2(n6855), .Z(n36117) );
  XOR2_X1 U24859 ( .A1(n38514), .A2(n18004), .Z(n5119) );
  XOR2_X1 U24871 ( .A1(n9390), .A2(n36119), .Z(n6593) );
  XOR2_X1 U24872 ( .A1(n31872), .A2(n7990), .Z(n36119) );
  AOI21_X2 U24874 ( .A1(n27232), .A2(n945), .B(n36120), .ZN(n20823) );
  XOR2_X1 U24882 ( .A1(n36123), .A2(n29017), .Z(Ciphertext[173]) );
  AOI22_X1 U24890 ( .A1(n29015), .A2(n30131), .B1(n29016), .B2(n3896), .ZN(
        n36123) );
  XOR2_X1 U24892 ( .A1(n27842), .A2(n7549), .Z(n21087) );
  NAND3_X2 U24900 ( .A1(n20434), .A2(n36126), .A3(n36125), .ZN(n20437) );
  XOR2_X1 U24912 ( .A1(n5750), .A2(n27855), .Z(n10782) );
  AND2_X2 U24926 ( .A1(n5899), .A2(n5966), .Z(n4915) );
  XOR2_X1 U24932 ( .A1(n13076), .A2(n18395), .Z(n36128) );
  OAI22_X2 U24944 ( .A1(n8968), .A2(n24866), .B1(n7970), .B2(n8314), .ZN(n7967) );
  OAI21_X1 U24947 ( .A1(n33976), .A2(n36135), .B(n25328), .ZN(n36134) );
  INV_X2 U24948 ( .I(n36136), .ZN(n4803) );
  NAND2_X2 U24955 ( .A1(n7781), .A2(n8248), .ZN(n16216) );
  NOR2_X2 U24961 ( .A1(n5734), .A2(n36139), .ZN(n4497) );
  XOR2_X1 U24964 ( .A1(n30913), .A2(n26499), .Z(n13673) );
  OAI21_X2 U24972 ( .A1(n5392), .A2(n5391), .B(n36140), .ZN(n5777) );
  INV_X2 U24973 ( .I(n36141), .ZN(n36140) );
  OAI21_X2 U24981 ( .A1(n19587), .A2(n5132), .B(n1155), .ZN(n36141) );
  OAI21_X1 U24984 ( .A1(n18910), .A2(n12543), .B(n36144), .ZN(n13028) );
  NOR3_X1 U25004 ( .A1(n1427), .A2(n28611), .A3(n8787), .ZN(n5927) );
  XOR2_X1 U25008 ( .A1(n6751), .A2(n6753), .Z(n28127) );
  BUF_X2 U25009 ( .I(n9616), .Z(n36151) );
  NAND2_X2 U25014 ( .A1(n20464), .A2(n20463), .ZN(n25345) );
  OAI21_X1 U25016 ( .A1(n19557), .A2(n27337), .B(n36152), .ZN(n27135) );
  XOR2_X1 U25043 ( .A1(n15844), .A2(n34162), .Z(n32842) );
  NAND2_X2 U25054 ( .A1(n29491), .A2(n1179), .ZN(n12428) );
  OR2_X1 U25061 ( .A1(n17072), .A2(n13699), .Z(n32962) );
  NOR2_X2 U25062 ( .A1(n33668), .A2(n16124), .ZN(n17072) );
  NAND2_X2 U25068 ( .A1(n28433), .A2(n39423), .ZN(n28460) );
  OAI21_X2 U25083 ( .A1(n36164), .A2(n26799), .B(n10203), .ZN(n7973) );
  OAI21_X2 U25094 ( .A1(n14409), .A2(n14439), .B(n22804), .ZN(n12960) );
  INV_X2 U25107 ( .I(n36160), .ZN(n37045) );
  XOR2_X1 U25108 ( .A1(n5937), .A2(n5936), .Z(n36160) );
  OAI21_X2 U25115 ( .A1(n36816), .A2(n13460), .B(n1113), .ZN(n13320) );
  NAND2_X2 U25116 ( .A1(n5896), .A2(n24492), .ZN(n24763) );
  NAND3_X2 U25118 ( .A1(n36163), .A2(n25070), .A3(n25067), .ZN(n31242) );
  XOR2_X1 U25121 ( .A1(n8972), .A2(n30126), .Z(n25809) );
  NAND2_X1 U25134 ( .A1(n36524), .A2(n11150), .ZN(n30381) );
  XOR2_X1 U25140 ( .A1(n36168), .A2(n34239), .Z(Ciphertext[88]) );
  INV_X2 U25147 ( .I(n18032), .ZN(n25965) );
  NAND2_X2 U25157 ( .A1(n30988), .A2(n36612), .ZN(n18032) );
  NAND2_X2 U25168 ( .A1(n36170), .A2(n29173), .ZN(n13559) );
  AND2_X2 U25178 ( .A1(n30597), .A2(n36931), .Z(n26727) );
  INV_X1 U25183 ( .I(n29206), .ZN(n36171) );
  NAND2_X2 U25189 ( .A1(n1782), .A2(n1785), .ZN(n4302) );
  NAND3_X1 U25207 ( .A1(n29922), .A2(n31570), .A3(n3860), .ZN(n8583) );
  NOR2_X2 U25230 ( .A1(n15644), .A2(n36172), .ZN(n33512) );
  INV_X2 U25233 ( .I(n36173), .ZN(n833) );
  XOR2_X1 U25234 ( .A1(n15938), .A2(n15937), .Z(n36173) );
  AOI21_X2 U25257 ( .A1(n26834), .A2(n26835), .B(n38852), .ZN(n36175) );
  BUF_X4 U25277 ( .I(n23354), .Z(n36564) );
  NOR2_X1 U25285 ( .A1(n22171), .A2(n36176), .ZN(n1840) );
  XOR2_X1 U25302 ( .A1(n13235), .A2(n22638), .Z(n4560) );
  XOR2_X1 U25304 ( .A1(n19725), .A2(n24982), .Z(n25245) );
  NAND2_X2 U25307 ( .A1(n11906), .A2(n24823), .ZN(n24982) );
  NAND2_X2 U25308 ( .A1(n9824), .A2(n4179), .ZN(n33581) );
  NAND2_X1 U25314 ( .A1(n36180), .A2(n24819), .ZN(n8648) );
  XOR2_X1 U25321 ( .A1(n23740), .A2(n36181), .Z(n6156) );
  XOR2_X1 U25323 ( .A1(n6227), .A2(n20317), .Z(n36181) );
  NAND2_X1 U25324 ( .A1(n2487), .A2(n36182), .ZN(n2485) );
  BUF_X2 U25330 ( .I(n32205), .Z(n36183) );
  NAND2_X1 U25331 ( .A1(n17691), .A2(n17692), .ZN(n36184) );
  XOR2_X1 U25346 ( .A1(n24436), .A2(n21174), .Z(n36205) );
  INV_X2 U25349 ( .I(n19979), .ZN(n5896) );
  INV_X2 U25350 ( .I(n24492), .ZN(n36186) );
  NAND2_X2 U25384 ( .A1(n16964), .A2(n385), .ZN(n18910) );
  NAND2_X2 U25387 ( .A1(n28290), .A2(n877), .ZN(n27896) );
  XOR2_X1 U25394 ( .A1(n22736), .A2(n22737), .Z(n36190) );
  NAND2_X2 U25405 ( .A1(n33844), .A2(n36193), .ZN(n29437) );
  NAND2_X2 U25413 ( .A1(n36194), .A2(n25508), .ZN(n20851) );
  OAI21_X2 U25415 ( .A1(n10850), .A2(n38825), .B(n33327), .ZN(n36194) );
  OAI21_X1 U25417 ( .A1(n28750), .A2(n28745), .B(n33283), .ZN(n28523) );
  AOI21_X2 U25451 ( .A1(n22945), .A2(n19488), .B(n17083), .ZN(n23390) );
  XOR2_X1 U25454 ( .A1(n36195), .A2(n1765), .Z(n13587) );
  NAND2_X2 U25474 ( .A1(n12466), .A2(n3097), .ZN(n36588) );
  NAND2_X1 U25475 ( .A1(n36199), .A2(n1598), .ZN(n23816) );
  OAI21_X1 U25481 ( .A1(n24294), .A2(n8824), .B(n33939), .ZN(n36199) );
  AOI22_X1 U25490 ( .A1(n36201), .A2(n626), .B1(n10342), .B2(n11673), .ZN(
        n31437) );
  OAI21_X1 U25514 ( .A1(n1606), .A2(n18329), .B(n3398), .ZN(n36201) );
  INV_X2 U25523 ( .I(n37014), .ZN(n1135) );
  XOR2_X1 U25531 ( .A1(n36204), .A2(n15932), .Z(n30839) );
  XOR2_X1 U25542 ( .A1(n386), .A2(n19774), .Z(n36204) );
  XOR2_X1 U25547 ( .A1(n16021), .A2(n23790), .Z(n36206) );
  XNOR2_X1 U25548 ( .A1(n4278), .A2(n4277), .ZN(n36698) );
  NAND2_X2 U25554 ( .A1(n11006), .A2(n11005), .ZN(n19631) );
  NAND2_X2 U25558 ( .A1(n25261), .A2(n37052), .ZN(n25725) );
  XOR2_X1 U25560 ( .A1(n1463), .A2(n12999), .Z(n36211) );
  NOR2_X2 U25565 ( .A1(n34121), .A2(n11108), .ZN(n36212) );
  XOR2_X1 U25566 ( .A1(n22490), .A2(n13478), .Z(n13477) );
  NOR2_X1 U25568 ( .A1(n35260), .A2(n9815), .ZN(n37049) );
  NAND2_X1 U25571 ( .A1(n31199), .A2(n23380), .ZN(n14974) );
  NAND2_X2 U25572 ( .A1(n454), .A2(n10670), .ZN(n30097) );
  NAND2_X2 U25583 ( .A1(n30350), .A2(n36936), .ZN(n5028) );
  XOR2_X1 U25588 ( .A1(n25173), .A2(n24921), .Z(n11061) );
  OR2_X1 U25596 ( .A1(n36471), .A2(n35901), .Z(n31625) );
  INV_X2 U25619 ( .I(n17353), .ZN(n36216) );
  BUF_X2 U25636 ( .I(n14231), .Z(n36218) );
  XNOR2_X1 U25649 ( .A1(n28896), .A2(n32608), .ZN(n32465) );
  XOR2_X1 U25676 ( .A1(n8904), .A2(n35970), .Z(n18404) );
  INV_X2 U25688 ( .I(n14015), .ZN(n6908) );
  NAND3_X2 U25690 ( .A1(n30715), .A2(n12565), .A3(n12566), .ZN(n14015) );
  NAND2_X2 U25691 ( .A1(n17107), .A2(n2114), .ZN(n27767) );
  XOR2_X1 U25701 ( .A1(n8605), .A2(n25040), .Z(n17623) );
  XOR2_X1 U25704 ( .A1(n28796), .A2(n28795), .Z(n19224) );
  XOR2_X1 U25707 ( .A1(n26513), .A2(n844), .Z(n5177) );
  INV_X2 U25709 ( .I(n14751), .ZN(n24963) );
  NOR2_X2 U25717 ( .A1(n32347), .A2(n32348), .ZN(n32205) );
  OR3_X2 U25731 ( .A1(n32775), .A2(n25487), .A3(n10938), .Z(n14656) );
  OR2_X1 U25732 ( .A1(n15865), .A2(n8193), .Z(n12564) );
  XOR2_X1 U25745 ( .A1(n26207), .A2(n1507), .Z(n26393) );
  BUF_X4 U25760 ( .I(n30504), .Z(n36340) );
  NOR2_X2 U25766 ( .A1(n21319), .A2(n9846), .ZN(n36229) );
  XOR2_X1 U25768 ( .A1(n36231), .A2(n2120), .Z(n2117) );
  XOR2_X1 U25771 ( .A1(n39209), .A2(n6561), .Z(n36233) );
  XOR2_X1 U25775 ( .A1(n29095), .A2(n29145), .Z(n29255) );
  XOR2_X1 U25782 ( .A1(n7337), .A2(n22714), .Z(n22719) );
  NAND2_X2 U25786 ( .A1(n28091), .A2(n36236), .ZN(n28463) );
  XOR2_X1 U25794 ( .A1(n7055), .A2(n36238), .Z(n33315) );
  INV_X1 U25799 ( .I(n22715), .ZN(n36238) );
  NAND2_X2 U25800 ( .A1(n22090), .A2(n7490), .ZN(n22715) );
  NOR2_X1 U25806 ( .A1(n14704), .A2(n30280), .ZN(n11760) );
  NAND2_X2 U25814 ( .A1(n16034), .A2(n20019), .ZN(n36320) );
  XOR2_X1 U25840 ( .A1(n36240), .A2(n36239), .Z(n15386) );
  XOR2_X1 U25844 ( .A1(n8586), .A2(n11050), .Z(n36240) );
  XOR2_X1 U25850 ( .A1(n22710), .A2(n22464), .Z(n22667) );
  XOR2_X1 U25855 ( .A1(n37957), .A2(n23710), .Z(n23662) );
  XOR2_X1 U25858 ( .A1(n31410), .A2(n30756), .Z(n31305) );
  NAND2_X2 U25860 ( .A1(n8305), .A2(n34150), .ZN(n260) );
  BUF_X2 U25864 ( .I(n9422), .Z(n36245) );
  NAND2_X1 U25865 ( .A1(n32695), .A2(n20133), .ZN(n36250) );
  INV_X2 U25870 ( .I(n36253), .ZN(n37057) );
  INV_X2 U25875 ( .I(n38165), .ZN(n36254) );
  INV_X2 U25883 ( .I(n36257), .ZN(n26763) );
  XOR2_X1 U25884 ( .A1(n32734), .A2(n36258), .Z(n2895) );
  XOR2_X1 U25889 ( .A1(n25103), .A2(n36259), .Z(n36258) );
  BUF_X4 U25896 ( .I(n34603), .Z(n36263) );
  NAND3_X2 U25897 ( .A1(n23069), .A2(n6000), .A3(n11366), .ZN(n19005) );
  XOR2_X1 U25901 ( .A1(n5721), .A2(n5722), .Z(n252) );
  INV_X2 U25948 ( .I(n8182), .ZN(n15164) );
  XOR2_X1 U25951 ( .A1(n27697), .A2(n36260), .Z(n8182) );
  XOR2_X1 U25952 ( .A1(n19717), .A2(n36265), .Z(n10239) );
  NAND2_X2 U25957 ( .A1(n22381), .A2(n22380), .ZN(n19717) );
  NAND2_X2 U25959 ( .A1(n30780), .A2(n36266), .ZN(n28677) );
  NAND2_X1 U25965 ( .A1(n1086), .A2(n27589), .ZN(n12263) );
  NAND2_X2 U25980 ( .A1(n3264), .A2(n9609), .ZN(n11937) );
  XOR2_X1 U25990 ( .A1(n25141), .A2(n15779), .Z(n21207) );
  XOR2_X1 U26016 ( .A1(n26169), .A2(n9776), .Z(n36270) );
  INV_X2 U26025 ( .I(n28514), .ZN(n1881) );
  NAND2_X2 U26034 ( .A1(n32759), .A2(n1882), .ZN(n28514) );
  OAI21_X2 U26035 ( .A1(n26), .A2(n12793), .B(n37011), .ZN(n36271) );
  NAND2_X2 U26053 ( .A1(n27192), .A2(n31421), .ZN(n19355) );
  AOI22_X2 U26056 ( .A1(n36273), .A2(n15319), .B1(n32297), .B2(n14558), .ZN(
        n13624) );
  INV_X4 U26078 ( .I(n17424), .ZN(n36275) );
  XOR2_X1 U26085 ( .A1(n3488), .A2(n11722), .Z(n16647) );
  OAI21_X2 U26102 ( .A1(n33926), .A2(n23328), .B(n36279), .ZN(n18279) );
  NAND2_X1 U26106 ( .A1(n1763), .A2(n531), .ZN(n16954) );
  NAND3_X1 U26112 ( .A1(n12564), .A2(n19426), .A3(n38839), .ZN(n11521) );
  INV_X2 U26117 ( .I(n36283), .ZN(n8413) );
  XOR2_X1 U26118 ( .A1(n2594), .A2(n33653), .Z(n36284) );
  AOI22_X2 U26120 ( .A1(n8686), .A2(n26179), .B1(n924), .B2(n5746), .ZN(n5745)
         );
  XOR2_X1 U26127 ( .A1(n36286), .A2(n20874), .Z(n23074) );
  XOR2_X1 U26132 ( .A1(n30444), .A2(n22387), .Z(n36286) );
  NAND2_X2 U26143 ( .A1(n37103), .A2(n1092), .ZN(n26817) );
  OR2_X2 U26152 ( .A1(n19250), .A2(n36655), .Z(n36523) );
  XOR2_X1 U26155 ( .A1(n36289), .A2(n27732), .Z(n10002) );
  XOR2_X1 U26159 ( .A1(n7651), .A2(n7549), .Z(n36289) );
  AOI22_X1 U26176 ( .A1(n12450), .A2(n38420), .B1(n1404), .B2(n31667), .ZN(
        n2410) );
  XOR2_X1 U26177 ( .A1(n36291), .A2(n20502), .Z(n4633) );
  NAND2_X1 U26185 ( .A1(n17261), .A2(n187), .ZN(n36446) );
  BUF_X2 U26199 ( .I(n33440), .Z(n36293) );
  XOR2_X1 U26212 ( .A1(n8554), .A2(n8553), .Z(n9775) );
  NAND2_X2 U26220 ( .A1(n10650), .A2(n10649), .ZN(n17074) );
  OAI22_X2 U26229 ( .A1(n18028), .A2(n20476), .B1(n32164), .B2(n14450), .ZN(
        n17923) );
  XOR2_X1 U26236 ( .A1(n26208), .A2(n32386), .Z(n26211) );
  NOR2_X2 U26237 ( .A1(n36297), .A2(n21614), .ZN(n9736) );
  INV_X2 U26238 ( .I(n15113), .ZN(n32759) );
  NAND2_X2 U26243 ( .A1(n13458), .A2(n13455), .ZN(n15113) );
  XOR2_X1 U26244 ( .A1(n1794), .A2(n1792), .Z(n20026) );
  NAND3_X2 U26246 ( .A1(n20999), .A2(n22284), .A3(n21000), .ZN(n22464) );
  XOR2_X1 U26248 ( .A1(n33179), .A2(n23732), .Z(n18922) );
  INV_X2 U26255 ( .I(n12633), .ZN(n1122) );
  NAND2_X2 U26256 ( .A1(n16446), .A2(n16450), .ZN(n12633) );
  XOR2_X1 U26277 ( .A1(n17137), .A2(n17136), .Z(n17984) );
  NAND3_X2 U26278 ( .A1(n14444), .A2(n31820), .A3(n14656), .ZN(n18176) );
  XOR2_X1 U26288 ( .A1(n22466), .A2(n18189), .Z(n10107) );
  NAND2_X2 U26298 ( .A1(n36300), .A2(n18426), .ZN(n26582) );
  NAND2_X2 U26299 ( .A1(n23242), .A2(n21130), .ZN(n36876) );
  XOR2_X1 U26301 ( .A1(n25312), .A2(n25074), .Z(n15937) );
  XOR2_X1 U26304 ( .A1(n37038), .A2(n24935), .Z(n25074) );
  XOR2_X1 U26316 ( .A1(n13634), .A2(n15625), .Z(n21259) );
  NAND2_X2 U26320 ( .A1(n14593), .A2(n12817), .ZN(n15625) );
  NAND3_X2 U26323 ( .A1(n10795), .A2(n10796), .A3(n21255), .ZN(n27252) );
  XOR2_X1 U26326 ( .A1(n7256), .A2(n4009), .Z(n882) );
  OAI22_X2 U26327 ( .A1(n14129), .A2(n36263), .B1(n6514), .B2(n23594), .ZN(
        n11098) );
  NOR2_X2 U26339 ( .A1(n37237), .A2(n611), .ZN(n36302) );
  XOR2_X1 U26359 ( .A1(n17344), .A2(n1971), .Z(n36305) );
  NAND2_X2 U26389 ( .A1(n30728), .A2(n4916), .ZN(n4377) );
  OAI21_X2 U26390 ( .A1(n8392), .A2(n930), .B(n36308), .ZN(n18631) );
  NAND3_X2 U26391 ( .A1(n7258), .A2(n2534), .A3(n9959), .ZN(n36308) );
  NOR2_X1 U26395 ( .A1(n36310), .A2(n36309), .ZN(n20187) );
  NOR2_X1 U26396 ( .A1(n19813), .A2(n6448), .ZN(n36310) );
  XOR2_X1 U26397 ( .A1(n25141), .A2(n20409), .Z(n15265) );
  XOR2_X1 U26412 ( .A1(n22604), .A2(n6893), .Z(n22755) );
  XOR2_X1 U26416 ( .A1(n10112), .A2(n36311), .Z(n10111) );
  XOR2_X1 U26418 ( .A1(n26468), .A2(n34157), .Z(n36311) );
  OAI21_X1 U26428 ( .A1(n36490), .A2(n13998), .B(n21555), .ZN(n7414) );
  INV_X1 U26447 ( .I(n5750), .ZN(n36317) );
  XOR2_X1 U26452 ( .A1(n26370), .A2(n26486), .Z(n12114) );
  OAI22_X1 U26461 ( .A1(n34156), .A2(n9529), .B1(n26063), .B2(n19793), .ZN(
        n9086) );
  NAND2_X2 U26473 ( .A1(n36322), .A2(n9209), .ZN(n19670) );
  OAI22_X1 U26479 ( .A1(n17985), .A2(n20671), .B1(n17422), .B2(n11910), .ZN(
        n17420) );
  XOR2_X1 U26489 ( .A1(n3956), .A2(n36326), .Z(n3134) );
  XOR2_X1 U26493 ( .A1(n26529), .A2(n745), .Z(n36326) );
  XOR2_X1 U26498 ( .A1(n12818), .A2(n36327), .Z(n3663) );
  XOR2_X1 U26506 ( .A1(n22772), .A2(n37042), .Z(n36327) );
  NOR2_X1 U26507 ( .A1(n14011), .A2(n35232), .ZN(n43) );
  XOR2_X1 U26513 ( .A1(n26279), .A2(n32003), .Z(n25735) );
  XOR2_X1 U26533 ( .A1(n15222), .A2(n27816), .Z(n36329) );
  OR2_X1 U26539 ( .A1(n19203), .A2(n27383), .Z(n33370) );
  NAND2_X2 U26553 ( .A1(n2657), .A2(n25532), .ZN(n11292) );
  NAND2_X2 U26569 ( .A1(n9175), .A2(n5356), .ZN(n26083) );
  OR2_X1 U26580 ( .A1(n28152), .A2(n32186), .Z(n36712) );
  XOR2_X1 U26601 ( .A1(n36334), .A2(n3331), .Z(n36447) );
  XOR2_X1 U26606 ( .A1(n36335), .A2(n11553), .Z(n17292) );
  XOR2_X1 U26607 ( .A1(n14385), .A2(n25155), .Z(n36335) );
  NOR2_X2 U26616 ( .A1(n36337), .A2(n36336), .ZN(n12567) );
  INV_X2 U26620 ( .I(n36338), .ZN(n11512) );
  NAND2_X2 U26669 ( .A1(n17810), .A2(n19070), .ZN(n36341) );
  OAI22_X1 U26681 ( .A1(n21678), .A2(n36455), .B1(n21825), .B2(n21861), .ZN(
        n21679) );
  OAI22_X2 U26682 ( .A1(n36346), .A2(n14549), .B1(n18712), .B2(n18710), .ZN(
        n18711) );
  XOR2_X1 U26694 ( .A1(n36349), .A2(n1169), .Z(n17812) );
  OAI21_X1 U26696 ( .A1(n39830), .A2(n21023), .B(n35252), .ZN(n18107) );
  BUF_X2 U26697 ( .I(n21858), .Z(n36351) );
  OR2_X1 U26707 ( .A1(n14139), .A2(n22262), .Z(n21990) );
  OR2_X1 U26714 ( .A1(n33644), .A2(n7512), .Z(n36352) );
  NOR2_X2 U26722 ( .A1(n36606), .A2(n36353), .ZN(n33140) );
  INV_X1 U26724 ( .I(n36354), .ZN(n21919) );
  AOI21_X2 U26727 ( .A1(n21921), .A2(n36354), .B(n8468), .ZN(n15441) );
  NAND2_X1 U26728 ( .A1(n670), .A2(n293), .ZN(n36354) );
  NAND2_X2 U26746 ( .A1(n423), .A2(n422), .ZN(n36471) );
  INV_X2 U26749 ( .I(n36357), .ZN(n12246) );
  OAI21_X2 U26756 ( .A1(n1351), .A2(n36887), .B(n21656), .ZN(n36358) );
  XOR2_X1 U26760 ( .A1(n36360), .A2(n37129), .Z(n27643) );
  XOR2_X1 U26769 ( .A1(n27523), .A2(n27852), .Z(n36360) );
  INV_X2 U26773 ( .I(n22215), .ZN(n6576) );
  OAI22_X2 U26775 ( .A1(n15274), .A2(n15292), .B1(n11172), .B2(n21629), .ZN(
        n22215) );
  XOR2_X1 U26781 ( .A1(n37101), .A2(n36364), .Z(n36363) );
  INV_X1 U26789 ( .I(n29983), .ZN(n36364) );
  XOR2_X1 U26796 ( .A1(n4039), .A2(n26500), .Z(n36366) );
  XNOR2_X1 U26811 ( .A1(n23904), .A2(n23681), .ZN(n36646) );
  INV_X2 U26816 ( .I(n11354), .ZN(n36369) );
  AOI22_X1 U26818 ( .A1(n18483), .A2(n30112), .B1(n32933), .B2(n30102), .ZN(
        n30105) );
  OAI22_X2 U26826 ( .A1(n28611), .A2(n35173), .B1(n1434), .B2(n28496), .ZN(
        n28539) );
  NAND2_X2 U26827 ( .A1(n33620), .A2(n15570), .ZN(n28356) );
  OR2_X1 U26831 ( .A1(n34019), .A2(n21001), .Z(n20999) );
  XOR2_X1 U26834 ( .A1(n36372), .A2(n36373), .Z(n33008) );
  NAND2_X1 U26846 ( .A1(n35895), .A2(n27320), .ZN(n18669) );
  XOR2_X1 U26858 ( .A1(n36377), .A2(n29162), .Z(n11384) );
  XOR2_X1 U26860 ( .A1(n9131), .A2(n1411), .Z(n36377) );
  NOR2_X2 U26861 ( .A1(n1603), .A2(n15320), .ZN(n32297) );
  XOR2_X1 U26864 ( .A1(n31563), .A2(n34135), .Z(n12830) );
  XOR2_X1 U26880 ( .A1(n24006), .A2(n24007), .Z(n36379) );
  XOR2_X1 U26888 ( .A1(n25155), .A2(n24922), .Z(n14214) );
  NAND2_X2 U26890 ( .A1(n685), .A2(n10652), .ZN(n15350) );
  XOR2_X1 U26897 ( .A1(n13504), .A2(n36388), .Z(n13503) );
  XOR2_X1 U26898 ( .A1(n8113), .A2(n8982), .Z(n36388) );
  XOR2_X1 U26903 ( .A1(n11372), .A2(n23898), .Z(n36389) );
  OR2_X1 U26904 ( .A1(n25808), .A2(n33997), .Z(n3806) );
  INV_X2 U26928 ( .I(n20573), .ZN(n36392) );
  XOR2_X1 U26932 ( .A1(n17039), .A2(n6433), .Z(n28946) );
  AOI21_X2 U26937 ( .A1(n28799), .A2(n28798), .B(n28670), .ZN(n17039) );
  INV_X2 U26947 ( .I(n19675), .ZN(n28669) );
  OAI22_X2 U26948 ( .A1(n15204), .A2(n31832), .B1(n15014), .B2(n17477), .ZN(
        n19675) );
  INV_X2 U26953 ( .I(n36396), .ZN(n37061) );
  NOR2_X2 U26968 ( .A1(n1119), .A2(n7810), .ZN(n548) );
  XOR2_X1 U26995 ( .A1(n7744), .A2(n30122), .Z(n9777) );
  NOR2_X2 U26998 ( .A1(n38302), .A2(n6849), .ZN(n6850) );
  XOR2_X1 U26999 ( .A1(n36400), .A2(n30682), .Z(Ciphertext[130]) );
  NOR2_X1 U27010 ( .A1(n31726), .A2(n31727), .ZN(n36400) );
  XOR2_X1 U27013 ( .A1(n11667), .A2(n38218), .Z(n25595) );
  XOR2_X1 U27016 ( .A1(n28984), .A2(n31398), .Z(n31377) );
  XOR2_X1 U27017 ( .A1(n10237), .A2(n36406), .Z(n10247) );
  NAND2_X2 U27027 ( .A1(n36408), .A2(n2635), .ZN(n25284) );
  AOI21_X1 U27047 ( .A1(n31231), .A2(n13986), .B(n15189), .ZN(n36410) );
  OAI21_X2 U27049 ( .A1(n36412), .A2(n36411), .B(n19813), .ZN(n20186) );
  NOR3_X1 U27080 ( .A1(n36415), .A2(n36413), .A3(n5152), .ZN(n5151) );
  NOR2_X1 U27083 ( .A1(n36671), .A2(n36414), .ZN(n36413) );
  AND2_X1 U27093 ( .A1(n36671), .A2(n31015), .Z(n36415) );
  NAND2_X2 U27097 ( .A1(n36416), .A2(n15017), .ZN(n12243) );
  NAND3_X1 U27099 ( .A1(n34019), .A2(n13980), .A3(n21001), .ZN(n36416) );
  XOR2_X1 U27100 ( .A1(n24838), .A2(n36418), .Z(n7377) );
  XOR2_X1 U27103 ( .A1(n34142), .A2(n24836), .Z(n36418) );
  OR2_X1 U27108 ( .A1(n11726), .A2(n8413), .Z(n3255) );
  XOR2_X1 U27112 ( .A1(n23782), .A2(n599), .Z(n3167) );
  XOR2_X1 U27116 ( .A1(n31563), .A2(n34032), .Z(n36423) );
  NAND2_X1 U27126 ( .A1(n16366), .A2(n18920), .ZN(n30368) );
  AOI21_X2 U27132 ( .A1(n4226), .A2(n4225), .B(n34123), .ZN(n4224) );
  OAI21_X2 U27143 ( .A1(n14065), .A2(n3449), .B(n20004), .ZN(n33001) );
  INV_X2 U27154 ( .I(n36435), .ZN(n12066) );
  NAND2_X2 U27157 ( .A1(n16237), .A2(n997), .ZN(n27011) );
  NOR2_X2 U27176 ( .A1(n9835), .A2(n23477), .ZN(n12008) );
  OAI21_X2 U27187 ( .A1(n36441), .A2(n20752), .B(n21939), .ZN(n20751) );
  OAI21_X2 U27194 ( .A1(n36621), .A2(n36622), .B(n24357), .ZN(n33224) );
  XOR2_X1 U27200 ( .A1(n12997), .A2(n9808), .Z(n13413) );
  NAND2_X2 U27206 ( .A1(n36446), .A2(n4372), .ZN(n5084) );
  INV_X2 U27209 ( .I(n36447), .ZN(n32623) );
  BUF_X2 U27217 ( .I(n32024), .Z(n36448) );
  NOR2_X1 U27218 ( .A1(n36450), .A2(n3509), .ZN(n36449) );
  INV_X1 U27220 ( .I(n16569), .ZN(n36451) );
  INV_X1 U27224 ( .I(n36452), .ZN(n28172) );
  NAND2_X1 U27227 ( .A1(n19467), .A2(n32474), .ZN(n36452) );
  NAND2_X2 U27234 ( .A1(n4), .A2(n3), .ZN(n1487) );
  INV_X2 U27241 ( .I(n36454), .ZN(n7160) );
  INV_X1 U27247 ( .I(n21858), .ZN(n36455) );
  XOR2_X1 U27249 ( .A1(Plaintext[46]), .A2(Key[46]), .Z(n21858) );
  XOR2_X1 U27262 ( .A1(n13673), .A2(n13674), .Z(n36456) );
  XOR2_X1 U27269 ( .A1(n3530), .A2(n3529), .Z(n20482) );
  NAND2_X1 U27276 ( .A1(n37776), .A2(n28458), .ZN(n28383) );
  BUF_X2 U27286 ( .I(n23873), .Z(n36461) );
  XOR2_X1 U27290 ( .A1(n29294), .A2(n5991), .Z(n36939) );
  AOI21_X1 U27301 ( .A1(n27311), .A2(n16243), .B(n27412), .ZN(n33261) );
  XOR2_X1 U27303 ( .A1(n8782), .A2(n9038), .Z(n8781) );
  OAI21_X2 U27306 ( .A1(n21940), .A2(n21941), .B(n21939), .ZN(n36464) );
  XOR2_X1 U27339 ( .A1(n22704), .A2(n22702), .Z(n36869) );
  XOR2_X1 U27344 ( .A1(n22464), .A2(n19931), .Z(n22702) );
  XOR2_X1 U27349 ( .A1(n7762), .A2(n5517), .Z(n5709) );
  INV_X1 U27357 ( .I(n4123), .ZN(n22483) );
  NAND2_X2 U27365 ( .A1(n4121), .A2(n4122), .ZN(n4123) );
  XOR2_X1 U27371 ( .A1(n36468), .A2(n14302), .Z(n14060) );
  AOI22_X2 U27372 ( .A1(n12079), .A2(n2186), .B1(n22030), .B2(n11508), .ZN(
        n11507) );
  NOR2_X2 U27374 ( .A1(n5075), .A2(n37217), .ZN(n12079) );
  XOR2_X1 U27398 ( .A1(n22543), .A2(n6711), .Z(n6710) );
  XOR2_X1 U27399 ( .A1(n23933), .A2(n23883), .Z(n23835) );
  NOR2_X2 U27410 ( .A1(n16758), .A2(n16757), .ZN(n23933) );
  NOR2_X2 U27423 ( .A1(n27053), .A2(n27337), .ZN(n27344) );
  INV_X2 U27425 ( .I(n36470), .ZN(n19426) );
  XNOR2_X1 U27426 ( .A1(n16942), .A2(n20767), .ZN(n36470) );
  XOR2_X1 U27433 ( .A1(n18359), .A2(n22603), .Z(n17284) );
  NAND2_X1 U27441 ( .A1(n3869), .A2(n24477), .ZN(n16159) );
  OAI21_X2 U27447 ( .A1(n20565), .A2(n25526), .B(n1539), .ZN(n36472) );
  OR2_X1 U27456 ( .A1(n20735), .A2(n21145), .Z(n36474) );
  NAND2_X2 U27462 ( .A1(n36476), .A2(n13698), .ZN(n27392) );
  OAI21_X2 U27485 ( .A1(n34040), .A2(n24514), .B(n31797), .ZN(n25104) );
  XOR2_X1 U27499 ( .A1(n26290), .A2(n26379), .Z(n26242) );
  AND2_X1 U27524 ( .A1(n18157), .A2(n33550), .Z(n33141) );
  BUF_X2 U27537 ( .I(n24411), .Z(n36485) );
  AOI21_X2 U27553 ( .A1(n36885), .A2(n32930), .B(n32024), .ZN(n17093) );
  INV_X2 U27561 ( .I(n39820), .ZN(n36486) );
  NOR2_X2 U27562 ( .A1(n36488), .A2(n36487), .ZN(n18838) );
  NAND2_X2 U27581 ( .A1(n18605), .A2(n30585), .ZN(n16835) );
  XNOR2_X1 U27584 ( .A1(n14902), .A2(n22787), .ZN(n16802) );
  XOR2_X1 U27590 ( .A1(n22671), .A2(n16798), .Z(n14902) );
  OAI22_X2 U27602 ( .A1(n34067), .A2(n36490), .B1(n19483), .B2(n10144), .ZN(
        n11173) );
  INV_X2 U27603 ( .I(n13959), .ZN(n36490) );
  XOR2_X1 U27610 ( .A1(n36491), .A2(n19879), .Z(Ciphertext[63]) );
  NAND3_X2 U27615 ( .A1(n7437), .A2(n7436), .A3(n7435), .ZN(n36491) );
  XOR2_X1 U27622 ( .A1(n2662), .A2(n36493), .Z(n33947) );
  XOR2_X1 U27636 ( .A1(n24981), .A2(n36494), .Z(n36493) );
  OAI22_X2 U27652 ( .A1(n20496), .A2(n20495), .B1(n28460), .B2(n28378), .ZN(
        n20492) );
  XOR2_X1 U27665 ( .A1(n28041), .A2(n36498), .Z(n19920) );
  XOR2_X1 U27666 ( .A1(n28040), .A2(n18159), .Z(n36498) );
  NAND2_X2 U27673 ( .A1(n3004), .A2(n36499), .ZN(n2349) );
  INV_X4 U27679 ( .I(n3455), .ZN(n16200) );
  NAND2_X2 U27681 ( .A1(n3175), .A2(n30813), .ZN(n3455) );
  NAND2_X2 U27682 ( .A1(n18718), .A2(n19504), .ZN(n36840) );
  NAND2_X2 U27687 ( .A1(n8990), .A2(n36501), .ZN(n8798) );
  NAND2_X2 U27696 ( .A1(n36502), .A2(n24856), .ZN(n18536) );
  OAI21_X2 U27703 ( .A1(n20690), .A2(n20689), .B(n24853), .ZN(n36502) );
  OR2_X1 U27726 ( .A1(n28205), .A2(n118), .Z(n14361) );
  XOR2_X1 U27732 ( .A1(n26181), .A2(n34165), .Z(n26368) );
  NOR3_X1 U27742 ( .A1(n10436), .A2(n8452), .A3(n23159), .ZN(n36506) );
  NOR2_X1 U27753 ( .A1(n16786), .A2(n14254), .ZN(n7194) );
  XOR2_X1 U27754 ( .A1(n33962), .A2(n16787), .Z(n16786) );
  NAND3_X2 U27760 ( .A1(n33675), .A2(n8914), .A3(n8913), .ZN(n29052) );
  XOR2_X1 U27767 ( .A1(n32766), .A2(n26542), .Z(n36508) );
  XOR2_X1 U27776 ( .A1(n26415), .A2(n36511), .Z(n36510) );
  XOR2_X1 U27791 ( .A1(n36758), .A2(n36513), .Z(n746) );
  INV_X2 U27813 ( .I(n36514), .ZN(n30186) );
  XOR2_X1 U27827 ( .A1(n7944), .A2(n36516), .Z(n36515) );
  INV_X2 U27830 ( .I(n3448), .ZN(n36516) );
  NAND2_X2 U27835 ( .A1(n25354), .A2(n25353), .ZN(n36922) );
  NAND2_X2 U27844 ( .A1(n35232), .A2(n31612), .ZN(n23636) );
  OAI21_X2 U27858 ( .A1(n18742), .A2(n15437), .B(n36518), .ZN(n9616) );
  XOR2_X1 U27862 ( .A1(n19862), .A2(n1553), .Z(n2184) );
  INV_X4 U27868 ( .I(n36523), .ZN(n5101) );
  NAND2_X1 U27880 ( .A1(n17710), .A2(n24145), .ZN(n14051) );
  INV_X2 U27899 ( .I(n28117), .ZN(n3159) );
  NOR2_X1 U27905 ( .A1(n36532), .A2(n1827), .ZN(n8156) );
  XOR2_X1 U27921 ( .A1(n21098), .A2(n20082), .Z(n14319) );
  NOR2_X1 U27934 ( .A1(n34279), .A2(n31433), .ZN(n30486) );
  OAI21_X2 U27937 ( .A1(n26353), .A2(n18606), .B(n14824), .ZN(n31433) );
  INV_X2 U27943 ( .I(n29113), .ZN(n5153) );
  NAND2_X2 U27944 ( .A1(n5154), .A2(n1741), .ZN(n29113) );
  XOR2_X1 U27945 ( .A1(n36537), .A2(n12179), .Z(n14401) );
  AND2_X1 U27954 ( .A1(n6592), .A2(n18545), .Z(n25676) );
  XOR2_X1 U27974 ( .A1(n23959), .A2(n36541), .Z(n36540) );
  INV_X2 U27976 ( .I(n23487), .ZN(n21247) );
  NAND2_X2 U27977 ( .A1(n22983), .A2(n22984), .ZN(n23487) );
  NAND2_X1 U28002 ( .A1(n5207), .A2(n5206), .ZN(n5205) );
  INV_X2 U28012 ( .I(n36543), .ZN(n668) );
  XOR2_X1 U28013 ( .A1(Plaintext[180]), .A2(Key[180]), .Z(n36543) );
  XOR2_X1 U28024 ( .A1(n6513), .A2(n6511), .Z(n18707) );
  INV_X1 U28035 ( .I(n26828), .ZN(n32892) );
  NAND2_X1 U28036 ( .A1(n15386), .A2(n32623), .ZN(n26828) );
  NOR2_X1 U28044 ( .A1(n29384), .A2(n31279), .ZN(n36550) );
  NAND2_X2 U28048 ( .A1(n21246), .A2(n36551), .ZN(n23600) );
  INV_X2 U28049 ( .I(n22973), .ZN(n36554) );
  NAND2_X1 U28064 ( .A1(n21052), .A2(n35809), .ZN(n30728) );
  NAND2_X1 U28069 ( .A1(n23034), .A2(n23035), .ZN(n23037) );
  NOR2_X1 U28078 ( .A1(n28048), .A2(n34410), .ZN(n36558) );
  INV_X1 U28081 ( .I(n4975), .ZN(n36559) );
  NOR2_X1 U28085 ( .A1(n30015), .A2(n30037), .ZN(n30031) );
  XOR2_X1 U28113 ( .A1(n23980), .A2(n32174), .Z(n21267) );
  NAND2_X2 U28116 ( .A1(n8138), .A2(n32506), .ZN(n23980) );
  OAI21_X2 U28121 ( .A1(n2574), .A2(n36568), .B(n2679), .ZN(n5031) );
  INV_X4 U28157 ( .I(n23426), .ZN(n2798) );
  XOR2_X1 U28195 ( .A1(n27756), .A2(n9184), .Z(n10818) );
  NOR2_X1 U28196 ( .A1(n29683), .A2(n31538), .ZN(n18794) );
  AND2_X1 U28235 ( .A1(n36571), .A2(n33440), .Z(n10889) );
  XOR2_X1 U28248 ( .A1(n23852), .A2(n36572), .Z(n16245) );
  XOR2_X1 U28249 ( .A1(n13978), .A2(n6561), .Z(n36572) );
  XOR2_X1 U28252 ( .A1(n36576), .A2(n24990), .Z(n25546) );
  XOR2_X1 U28255 ( .A1(n9389), .A2(n729), .Z(n36576) );
  NAND2_X2 U28267 ( .A1(n36577), .A2(n17441), .ZN(n23888) );
  OAI21_X2 U28295 ( .A1(n6514), .A2(n36263), .B(n19232), .ZN(n23416) );
  XOR2_X1 U28304 ( .A1(n26454), .A2(n26433), .Z(n11072) );
  NAND2_X2 U28311 ( .A1(n14988), .A2(n14990), .ZN(n27448) );
  NOR3_X1 U28324 ( .A1(n11226), .A2(n36480), .A3(n38377), .ZN(n3402) );
  NAND2_X1 U28338 ( .A1(n13226), .A2(n1143), .ZN(n22369) );
  NAND2_X1 U28345 ( .A1(n6543), .A2(n25860), .ZN(n36581) );
  NAND2_X2 U28365 ( .A1(n1587), .A2(n24398), .ZN(n9583) );
  NAND2_X2 U28366 ( .A1(n9783), .A2(n33574), .ZN(n10079) );
  INV_X1 U28373 ( .I(n998), .ZN(n27189) );
  NOR2_X2 U28384 ( .A1(n36584), .A2(n24163), .ZN(n7770) );
  NAND2_X1 U28420 ( .A1(n17677), .A2(n38656), .ZN(n36587) );
  OR2_X1 U28429 ( .A1(n7291), .A2(n9875), .Z(n36679) );
  NAND2_X2 U28457 ( .A1(n20604), .A2(n36589), .ZN(n21272) );
  NOR2_X2 U28480 ( .A1(n29779), .A2(n29776), .ZN(n36590) );
  AOI21_X2 U28506 ( .A1(n36593), .A2(n36592), .B(n35611), .ZN(n18565) );
  NAND2_X2 U28513 ( .A1(n36594), .A2(n3083), .ZN(n11922) );
  NOR2_X2 U28521 ( .A1(n12324), .A2(n12325), .ZN(n20353) );
  OAI21_X2 U28546 ( .A1(n21564), .A2(n19397), .B(n11433), .ZN(n22113) );
  NOR2_X2 U28547 ( .A1(n30835), .A2(n9190), .ZN(n16236) );
  NAND2_X2 U28548 ( .A1(n36598), .A2(n14762), .ZN(n18273) );
  OR2_X1 U28553 ( .A1(n12235), .A2(n8205), .Z(n16666) );
  XOR2_X1 U28557 ( .A1(n32219), .A2(n14978), .Z(n15037) );
  OAI21_X1 U28558 ( .A1(n4192), .A2(n32566), .B(n38187), .ZN(n2502) );
  AOI21_X2 U28559 ( .A1(n2428), .A2(n3088), .B(n32940), .ZN(n27845) );
  NOR2_X2 U28562 ( .A1(n33412), .A2(n24821), .ZN(n6770) );
  NAND2_X1 U28589 ( .A1(n29699), .A2(n29195), .ZN(n29633) );
  INV_X2 U28605 ( .I(n36601), .ZN(n858) );
  XOR2_X1 U28611 ( .A1(n15818), .A2(n15821), .Z(n36601) );
  NOR2_X1 U28614 ( .A1(n36981), .A2(n27240), .ZN(n17354) );
  XOR2_X1 U28618 ( .A1(n36603), .A2(n36602), .Z(n31272) );
  NOR2_X1 U28644 ( .A1(n28330), .A2(n17583), .ZN(n28738) );
  XOR2_X1 U28662 ( .A1(n14294), .A2(n36604), .Z(n550) );
  XOR2_X1 U28663 ( .A1(n9937), .A2(n36605), .Z(n36604) );
  NOR3_X1 U28669 ( .A1(n14600), .A2(n14158), .A3(n29815), .ZN(n17912) );
  AOI21_X2 U28670 ( .A1(n21558), .A2(n21559), .B(n21920), .ZN(n36606) );
  XOR2_X1 U28673 ( .A1(n36608), .A2(n8547), .Z(n8546) );
  XOR2_X1 U28674 ( .A1(n17812), .A2(n22444), .Z(n36608) );
  XOR2_X1 U28703 ( .A1(n31563), .A2(n3576), .Z(n3579) );
  NOR2_X2 U28737 ( .A1(n2759), .A2(n21672), .ZN(n31480) );
  NAND2_X1 U28755 ( .A1(n14877), .A2(n19724), .ZN(n14876) );
  AOI21_X2 U28759 ( .A1(n36611), .A2(n20515), .B(n3602), .ZN(n10775) );
  NAND2_X2 U28767 ( .A1(n7802), .A2(n19495), .ZN(n36611) );
  NAND2_X1 U28775 ( .A1(n29632), .A2(n29701), .ZN(n29197) );
  XOR2_X1 U28778 ( .A1(n36613), .A2(n33309), .Z(n21126) );
  XOR2_X1 U28789 ( .A1(n36223), .A2(n10673), .Z(n36613) );
  XOR2_X1 U28810 ( .A1(n32448), .A2(n11923), .Z(n11015) );
  AND3_X1 U28832 ( .A1(n16240), .A2(n31362), .A3(n33514), .Z(n7888) );
  NAND3_X2 U28837 ( .A1(n36615), .A2(n10676), .A3(n35777), .ZN(n9955) );
  OAI21_X1 U28854 ( .A1(n32651), .A2(n24565), .B(n36618), .ZN(n20301) );
  NAND2_X2 U28876 ( .A1(n17687), .A2(n18986), .ZN(n27466) );
  INV_X2 U28877 ( .I(n36620), .ZN(n10047) );
  XOR2_X1 U28880 ( .A1(n16563), .A2(n16560), .Z(n36620) );
  XOR2_X1 U28890 ( .A1(n5836), .A2(n3233), .Z(n3232) );
  NOR2_X2 U28892 ( .A1(n11173), .A2(n11174), .ZN(n11327) );
  NOR2_X1 U28918 ( .A1(n32099), .A2(n19499), .ZN(n7261) );
  NAND2_X2 U28921 ( .A1(n7263), .A2(n10791), .ZN(n9053) );
  XOR2_X1 U28934 ( .A1(n27840), .A2(n18650), .Z(n13791) );
  NAND2_X2 U29008 ( .A1(n19539), .A2(n19540), .ZN(n30096) );
  AOI21_X2 U29018 ( .A1(n18328), .A2(n30526), .B(n1606), .ZN(n36626) );
  XOR2_X1 U29024 ( .A1(n36627), .A2(n27881), .Z(n29483) );
  XOR2_X1 U29026 ( .A1(n13381), .A2(n27880), .Z(n36627) );
  OAI21_X2 U29029 ( .A1(n10564), .A2(n10565), .B(n32009), .ZN(n31048) );
  XOR2_X1 U29031 ( .A1(n38560), .A2(n30865), .Z(n16431) );
  OAI21_X1 U29033 ( .A1(n31859), .A2(n1331), .B(n31860), .ZN(n18729) );
  XOR2_X1 U29041 ( .A1(n31261), .A2(n19881), .Z(n32001) );
  XOR2_X1 U29051 ( .A1(n4612), .A2(n23717), .Z(n23722) );
  XOR2_X1 U29056 ( .A1(n25286), .A2(n25081), .Z(n5816) );
  XOR2_X1 U29063 ( .A1(n11321), .A2(n25014), .Z(n25081) );
  INV_X1 U29072 ( .I(n25355), .ZN(n25449) );
  XOR2_X1 U29073 ( .A1(n17108), .A2(n36799), .Z(n25355) );
  NAND2_X2 U29074 ( .A1(n36629), .A2(n12075), .ZN(n27697) );
  NOR2_X2 U29077 ( .A1(n12073), .A2(n12072), .ZN(n36629) );
  OAI21_X2 U29081 ( .A1(n36443), .A2(n32609), .B(n36631), .ZN(n9735) );
  NAND2_X2 U29086 ( .A1(n36632), .A2(n32609), .ZN(n36631) );
  XOR2_X1 U29122 ( .A1(n36637), .A2(n8401), .Z(n8301) );
  XOR2_X1 U29143 ( .A1(n9712), .A2(n32203), .Z(n17198) );
  INV_X2 U29148 ( .I(n2430), .ZN(n22899) );
  XOR2_X1 U29152 ( .A1(n2200), .A2(n2198), .Z(n2430) );
  NAND2_X1 U29171 ( .A1(n5966), .A2(n17405), .ZN(n28045) );
  XOR2_X1 U29180 ( .A1(n25809), .A2(n16294), .Z(n36644) );
  XOR2_X1 U29203 ( .A1(n12515), .A2(n16278), .Z(n36645) );
  XOR2_X1 U29204 ( .A1(n737), .A2(n26401), .Z(n6963) );
  NAND2_X1 U29209 ( .A1(n5174), .A2(n11616), .ZN(n36957) );
  BUF_X2 U29214 ( .I(n4342), .Z(n36649) );
  OR2_X1 U29219 ( .A1(n13998), .A2(n18959), .Z(n13956) );
  OAI21_X1 U29220 ( .A1(n34066), .A2(n21645), .B(n36651), .ZN(n21648) );
  NAND2_X1 U29223 ( .A1(n21642), .A2(n21645), .ZN(n36651) );
  NAND2_X2 U29226 ( .A1(n16732), .A2(n16731), .ZN(n32024) );
  NAND2_X1 U29228 ( .A1(n22822), .A2(n7387), .ZN(n36654) );
  XOR2_X1 U29240 ( .A1(n10399), .A2(n1457), .Z(n36656) );
  NAND2_X2 U29246 ( .A1(n2736), .A2(n2737), .ZN(n4108) );
  XOR2_X1 U29247 ( .A1(n5802), .A2(n12139), .Z(n13205) );
  AOI22_X2 U29259 ( .A1(n13009), .A2(n11044), .B1(n8792), .B2(n196), .ZN(
        n13008) );
  NAND2_X2 U29276 ( .A1(n32832), .A2(n8362), .ZN(n17454) );
  OAI21_X2 U29286 ( .A1(n7216), .A2(n1339), .B(n36661), .ZN(n36660) );
  XOR2_X1 U29287 ( .A1(n13977), .A2(n19344), .Z(n19343) );
  XOR2_X1 U29295 ( .A1(n25263), .A2(n18432), .Z(n17593) );
  BUF_X2 U29297 ( .I(n7063), .Z(n36663) );
  XOR2_X1 U29298 ( .A1(n31823), .A2(n26480), .Z(n26182) );
  XOR2_X1 U29306 ( .A1(n36727), .A2(n16753), .Z(n33182) );
  NAND2_X2 U29312 ( .A1(n32292), .A2(n18825), .ZN(n22240) );
  INV_X2 U29333 ( .I(n26128), .ZN(n36666) );
  XOR2_X1 U29371 ( .A1(n4875), .A2(n6523), .Z(n5534) );
  NAND2_X1 U29377 ( .A1(n36674), .A2(n8691), .ZN(n20074) );
  OAI21_X2 U29386 ( .A1(n29988), .A2(n30051), .B(n10943), .ZN(n30038) );
  OAI22_X2 U29392 ( .A1(n15936), .A2(n36673), .B1(n7267), .B2(n24799), .ZN(
        n14781) );
  NAND2_X2 U29400 ( .A1(n22828), .A2(n20907), .ZN(n5258) );
  XOR2_X1 U29445 ( .A1(n38816), .A2(n31218), .Z(n36687) );
  XOR2_X1 U29470 ( .A1(n6661), .A2(n30101), .Z(n28986) );
  NAND2_X1 U29483 ( .A1(n29207), .A2(n11973), .ZN(n9807) );
  NOR2_X1 U29494 ( .A1(n19610), .A2(n36691), .ZN(n19482) );
  NOR2_X1 U29498 ( .A1(n21141), .A2(n19893), .ZN(n36691) );
  XOR2_X1 U29516 ( .A1(n20554), .A2(n36692), .Z(n30562) );
  XOR2_X1 U29517 ( .A1(n25016), .A2(n25324), .Z(n36692) );
  XOR2_X1 U29518 ( .A1(n23725), .A2(n17563), .Z(n10941) );
  NAND3_X1 U29520 ( .A1(n15043), .A2(n15044), .A3(n29410), .ZN(n7733) );
  AND2_X1 U29528 ( .A1(n31287), .A2(n27424), .Z(n30475) );
  NAND2_X1 U29529 ( .A1(n33201), .A2(n33202), .ZN(n33200) );
  NAND2_X2 U29541 ( .A1(n22805), .A2(n36696), .ZN(n14856) );
  OAI22_X2 U29552 ( .A1(n12960), .A2(n32740), .B1(n22892), .B2(n33925), .ZN(
        n36696) );
  OAI22_X1 U29553 ( .A1(n3039), .A2(n5569), .B1(n38601), .B2(n3040), .ZN(
        n16197) );
  XOR2_X1 U29554 ( .A1(n4279), .A2(n36698), .Z(n31920) );
  NOR2_X1 U29557 ( .A1(n31271), .A2(n8193), .ZN(n5) );
  NOR2_X2 U29561 ( .A1(n29591), .A2(n28550), .ZN(n2296) );
  XOR2_X1 U29585 ( .A1(n29835), .A2(n36702), .Z(n12763) );
  XOR2_X1 U29587 ( .A1(n12765), .A2(n28819), .Z(n36702) );
  AOI21_X2 U29588 ( .A1(n9816), .A2(n13375), .B(n12417), .ZN(n12416) );
  NOR2_X2 U29594 ( .A1(n39671), .A2(n20740), .ZN(n27232) );
  NOR2_X1 U29607 ( .A1(n16154), .A2(n37671), .ZN(n36703) );
  XOR2_X1 U29615 ( .A1(n3521), .A2(n5185), .Z(n12973) );
  INV_X2 U29619 ( .I(n18994), .ZN(n1245) );
  NAND2_X1 U29635 ( .A1(n1046), .A2(n23140), .ZN(n21047) );
  AOI22_X2 U29667 ( .A1(n20411), .A2(n3120), .B1(n11710), .B2(n24847), .ZN(
        n24731) );
  OR2_X1 U29671 ( .A1(n21339), .A2(n21687), .Z(n4750) );
  AOI21_X2 U29682 ( .A1(n9721), .A2(n36712), .B(n33902), .ZN(n30837) );
  OAI22_X2 U29716 ( .A1(n1071), .A2(n20157), .B1(n28118), .B2(n19667), .ZN(
        n28140) );
  XOR2_X1 U29717 ( .A1(n22754), .A2(n18001), .Z(n5571) );
  INV_X2 U29737 ( .I(n36717), .ZN(n37051) );
  XOR2_X1 U29745 ( .A1(n36718), .A2(n13928), .Z(n17022) );
  XOR2_X1 U29749 ( .A1(n31790), .A2(n26408), .Z(n36718) );
  XOR2_X1 U29753 ( .A1(n3553), .A2(n36719), .Z(n5078) );
  XOR2_X1 U29760 ( .A1(n35065), .A2(n13193), .Z(n2739) );
  NOR2_X2 U29779 ( .A1(n15466), .A2(n12044), .ZN(n21929) );
  NAND2_X2 U29797 ( .A1(n32577), .A2(n26717), .ZN(n21101) );
  XOR2_X1 U29799 ( .A1(n22678), .A2(n36723), .Z(n23131) );
  XOR2_X1 U29801 ( .A1(n11985), .A2(n11984), .Z(n36723) );
  NAND2_X1 U29802 ( .A1(n22313), .A2(n36151), .ZN(n22314) );
  NOR2_X2 U29804 ( .A1(n18636), .A2(n32753), .ZN(n36726) );
  XOR2_X1 U29806 ( .A1(n10982), .A2(n10984), .Z(n27882) );
  XOR2_X1 U29816 ( .A1(n1658), .A2(n4819), .Z(n36727) );
  NOR2_X2 U29820 ( .A1(n22254), .A2(n32675), .ZN(n22126) );
  XOR2_X1 U29826 ( .A1(n10484), .A2(n10486), .Z(n19746) );
  OAI21_X1 U29833 ( .A1(n1787), .A2(n1095), .B(n14380), .ZN(n26954) );
  NAND2_X2 U29849 ( .A1(n13096), .A2(n26958), .ZN(n19529) );
  OAI21_X2 U29852 ( .A1(n12461), .A2(n12460), .B(n36729), .ZN(n25301) );
  XOR2_X1 U29861 ( .A1(n24974), .A2(n36730), .Z(n31410) );
  XOR2_X1 U29863 ( .A1(n26376), .A2(n26289), .Z(n8844) );
  XOR2_X1 U29882 ( .A1(n19384), .A2(n26582), .Z(n26286) );
  XOR2_X1 U29888 ( .A1(n36734), .A2(n25311), .Z(n15034) );
  XOR2_X1 U29891 ( .A1(n25031), .A2(n6066), .Z(n36734) );
  XOR2_X1 U29899 ( .A1(Plaintext[55]), .A2(Key[55]), .Z(n7703) );
  INV_X2 U29900 ( .I(n13359), .ZN(n36735) );
  NAND2_X1 U29918 ( .A1(n36738), .A2(n30217), .ZN(n36737) );
  NAND3_X1 U29941 ( .A1(n14869), .A2(n30211), .A3(n33437), .ZN(n31987) );
  NOR2_X1 U29945 ( .A1(n1068), .A2(n28591), .ZN(n4992) );
  OAI22_X2 U29948 ( .A1(n36944), .A2(n28176), .B1(n28265), .B2(n28175), .ZN(
        n28591) );
  OR2_X1 U29958 ( .A1(n26090), .A2(n35828), .Z(n25363) );
  NAND2_X1 U29961 ( .A1(n28267), .A2(n37079), .ZN(n31766) );
  NAND2_X2 U29963 ( .A1(n36741), .A2(n37279), .ZN(n2950) );
  NAND2_X2 U29966 ( .A1(n23340), .A2(n23341), .ZN(n36741) );
  NAND3_X2 U29973 ( .A1(n13282), .A2(n13281), .A3(n13280), .ZN(n6130) );
  NAND2_X1 U29979 ( .A1(n18412), .A2(n35977), .ZN(n8467) );
  AND2_X1 U29983 ( .A1(n38848), .A2(n33996), .Z(n18459) );
  NAND2_X1 U29992 ( .A1(n36745), .A2(n22317), .ZN(n36902) );
  NOR2_X1 U29994 ( .A1(n31766), .A2(n31765), .ZN(n36944) );
  OAI21_X2 U29998 ( .A1(n9735), .A2(n38746), .B(n9734), .ZN(n22657) );
  XOR2_X1 U29999 ( .A1(n35221), .A2(n22775), .Z(n22689) );
  NOR2_X2 U30000 ( .A1(n14800), .A2(n14801), .ZN(n11644) );
  AOI22_X1 U30008 ( .A1(n15230), .A2(n23042), .B1(n38329), .B2(n4714), .ZN(
        n11914) );
  INV_X2 U30020 ( .I(n24038), .ZN(n36748) );
  XOR2_X1 U30024 ( .A1(n36894), .A2(n19801), .Z(n16857) );
  XOR2_X1 U30025 ( .A1(n29245), .A2(n11127), .Z(n19727) );
  AOI21_X2 U30026 ( .A1(n21631), .A2(n36519), .B(n36751), .ZN(n21634) );
  OR2_X1 U30031 ( .A1(n10631), .A2(n20238), .Z(n36753) );
  XOR2_X1 U30032 ( .A1(n3823), .A2(n4118), .Z(n36992) );
  XNOR2_X1 U30033 ( .A1(n29300), .A2(n15617), .ZN(n28836) );
  NAND2_X2 U30036 ( .A1(n15514), .A2(n19726), .ZN(n29300) );
  OAI22_X2 U30040 ( .A1(n11213), .A2(n15237), .B1(n12090), .B2(n13186), .ZN(
        n31132) );
  XOR2_X1 U30057 ( .A1(n3616), .A2(n12664), .Z(n36759) );
  NAND2_X2 U30062 ( .A1(n7614), .A2(n36857), .ZN(n20159) );
  NAND2_X2 U30063 ( .A1(n33893), .A2(n5363), .ZN(n27452) );
  INV_X2 U30069 ( .I(n9917), .ZN(n28749) );
  NOR2_X2 U30076 ( .A1(n31934), .A2(n36761), .ZN(n17687) );
  BUF_X2 U30083 ( .I(n6205), .Z(n36764) );
  XOR2_X1 U30094 ( .A1(Plaintext[29]), .A2(Key[29]), .Z(n36772) );
  INV_X2 U30102 ( .I(n36772), .ZN(n21445) );
  NAND2_X1 U30124 ( .A1(n33765), .A2(n31664), .ZN(n36774) );
  NAND2_X2 U30125 ( .A1(n28700), .A2(n36777), .ZN(n36776) );
  NAND2_X2 U30128 ( .A1(n21956), .A2(n21957), .ZN(n22580) );
  NAND2_X2 U30133 ( .A1(n21486), .A2(n36779), .ZN(n22085) );
  AOI21_X2 U30136 ( .A1(n21120), .A2(n36782), .B(n21119), .ZN(n23473) );
  NAND2_X1 U30140 ( .A1(n13373), .A2(n36783), .ZN(n36782) );
  XOR2_X1 U30151 ( .A1(n30842), .A2(n9420), .Z(n18433) );
  XOR2_X1 U30157 ( .A1(n16492), .A2(n25269), .Z(n25161) );
  NAND3_X2 U30160 ( .A1(n16747), .A2(n2503), .A3(n16746), .ZN(n16492) );
  INV_X2 U30177 ( .I(n9339), .ZN(n10698) );
  NAND2_X1 U30180 ( .A1(n23152), .A2(n2572), .ZN(n9339) );
  XOR2_X1 U30206 ( .A1(n10039), .A2(n10248), .Z(n25581) );
  XOR2_X1 U30208 ( .A1(n24892), .A2(n24891), .Z(n36799) );
  XOR2_X1 U30209 ( .A1(n23736), .A2(n10771), .Z(n8016) );
  NOR3_X1 U30216 ( .A1(n14704), .A2(n4986), .A3(n12771), .ZN(n36800) );
  XOR2_X1 U30217 ( .A1(n19009), .A2(n11458), .Z(n11459) );
  XOR2_X1 U30221 ( .A1(n12588), .A2(n26285), .Z(n36803) );
  XOR2_X1 U30222 ( .A1(n479), .A2(n27648), .Z(n36804) );
  AOI21_X2 U30230 ( .A1(n25878), .A2(n25879), .B(n25877), .ZN(n6989) );
  NAND2_X2 U30232 ( .A1(n12889), .A2(n12888), .ZN(n28886) );
  OAI21_X2 U30233 ( .A1(n1521), .A2(n11036), .B(n36807), .ZN(n26403) );
  AOI21_X2 U30239 ( .A1(n37116), .A2(n1521), .B(n11032), .ZN(n36807) );
  AOI21_X1 U30244 ( .A1(n24228), .A2(n24328), .B(n1607), .ZN(n15496) );
  XOR2_X1 U30250 ( .A1(n36808), .A2(n1358), .Z(Ciphertext[107]) );
  XOR2_X1 U30257 ( .A1(n27673), .A2(n36809), .Z(n31043) );
  OAI21_X2 U30259 ( .A1(n18924), .A2(n13289), .B(n12240), .ZN(n27843) );
  NAND3_X2 U30260 ( .A1(n25405), .A2(n25406), .A3(n25404), .ZN(n3413) );
  AOI22_X1 U30261 ( .A1(n30185), .A2(n31846), .B1(n39122), .B2(n30182), .ZN(
        n4780) );
  XOR2_X1 U30270 ( .A1(n29246), .A2(n36837), .Z(n16787) );
  NAND2_X2 U30272 ( .A1(n33833), .A2(n13818), .ZN(n29246) );
  XOR2_X1 U30278 ( .A1(n36812), .A2(n19200), .Z(n15463) );
  INV_X2 U30288 ( .I(n30597), .ZN(n3449) );
  XOR2_X1 U30297 ( .A1(n38269), .A2(n38502), .Z(n26415) );
  NAND2_X2 U30303 ( .A1(n38874), .A2(n2716), .ZN(n36817) );
  NAND3_X2 U30305 ( .A1(n24511), .A2(n30414), .A3(n31986), .ZN(n24869) );
  XOR2_X1 U30306 ( .A1(n36822), .A2(n17406), .Z(n17405) );
  NAND2_X1 U30309 ( .A1(n30058), .A2(n37253), .ZN(n36824) );
  NAND2_X1 U30323 ( .A1(n37014), .A2(n36829), .ZN(n37010) );
  XOR2_X1 U30330 ( .A1(n36830), .A2(n16225), .Z(n16704) );
  XOR2_X1 U30337 ( .A1(n28979), .A2(n2914), .Z(n36830) );
  INV_X2 U30338 ( .I(n36831), .ZN(n30443) );
  XOR2_X1 U30340 ( .A1(n28983), .A2(n17880), .Z(n29026) );
  NAND2_X2 U30343 ( .A1(n15295), .A2(n7030), .ZN(n17880) );
  NAND2_X2 U30347 ( .A1(n15360), .A2(n3313), .ZN(n36833) );
  XOR2_X1 U30350 ( .A1(n31339), .A2(n39136), .Z(n12818) );
  NOR2_X2 U30352 ( .A1(n22376), .A2(n22375), .ZN(n31339) );
  AOI21_X2 U30364 ( .A1(n10618), .A2(n36835), .B(n888), .ZN(n3221) );
  XOR2_X1 U30372 ( .A1(n29289), .A2(n29081), .Z(n36837) );
  BUF_X2 U30374 ( .I(n4472), .Z(n36839) );
  XOR2_X1 U30376 ( .A1(n21267), .A2(n23784), .Z(n182) );
  XOR2_X1 U30377 ( .A1(n22542), .A2(n22656), .Z(n6709) );
  NAND2_X2 U30378 ( .A1(n36843), .A2(n8419), .ZN(n18081) );
  NOR2_X1 U30379 ( .A1(n6657), .A2(n32486), .ZN(n12131) );
  OAI22_X2 U30380 ( .A1(n11848), .A2(n33263), .B1(n8481), .B2(n834), .ZN(
        n25819) );
  XOR2_X1 U30392 ( .A1(n22771), .A2(n22393), .Z(n18914) );
  XOR2_X1 U30400 ( .A1(n36847), .A2(n13426), .Z(n13425) );
  XOR2_X1 U30403 ( .A1(n26258), .A2(n26257), .Z(n15453) );
  XOR2_X1 U30407 ( .A1(n35231), .A2(n19749), .Z(n16458) );
  XOR2_X1 U30421 ( .A1(n32309), .A2(n7481), .Z(n36851) );
  OAI21_X2 U30427 ( .A1(n26640), .A2(n26918), .B(n36853), .ZN(n5554) );
  NAND2_X1 U30428 ( .A1(n11700), .A2(n13786), .ZN(n13363) );
  NAND2_X2 U30438 ( .A1(n12379), .A2(n12378), .ZN(n12989) );
  OR2_X1 U30442 ( .A1(n25991), .A2(n25760), .Z(n33328) );
  INV_X2 U30446 ( .I(n36856), .ZN(n31557) );
  XOR2_X1 U30450 ( .A1(n4334), .A2(n4332), .Z(n36856) );
  XOR2_X1 U30457 ( .A1(n2739), .A2(n2738), .Z(n9022) );
  NAND2_X1 U30458 ( .A1(n550), .A2(n18415), .ZN(n6499) );
  NOR3_X1 U30459 ( .A1(n23042), .A2(n39096), .A3(n33431), .ZN(n14882) );
  XOR2_X1 U30462 ( .A1(n18051), .A2(n6523), .Z(n26500) );
  NAND2_X2 U30463 ( .A1(n5705), .A2(n16063), .ZN(n31015) );
  NAND2_X2 U30465 ( .A1(n21732), .A2(n11124), .ZN(n17126) );
  NAND2_X2 U30466 ( .A1(n33148), .A2(n21730), .ZN(n21732) );
  OAI22_X2 U30467 ( .A1(n20813), .A2(n1512), .B1(n10015), .B2(n26215), .ZN(
        n26038) );
  OAI22_X2 U30468 ( .A1(n12826), .A2(n17183), .B1(n31843), .B2(n31842), .ZN(
        n26215) );
  XOR2_X1 U30474 ( .A1(n27730), .A2(n9164), .Z(n36861) );
  XOR2_X1 U30487 ( .A1(n25080), .A2(n25196), .Z(n25286) );
  XOR2_X1 U30495 ( .A1(n33027), .A2(n26338), .Z(n26450) );
  AOI21_X2 U30497 ( .A1(n26053), .A2(n926), .B(n34153), .ZN(n2751) );
  INV_X2 U30498 ( .I(n36868), .ZN(n13686) );
  XOR2_X1 U30499 ( .A1(n10485), .A2(n25289), .Z(n10484) );
  INV_X4 U30512 ( .I(n36871), .ZN(n23531) );
  OAI22_X2 U30513 ( .A1(n23206), .A2(n36422), .B1(n23207), .B2(n14994), .ZN(
        n36871) );
  XOR2_X1 U30515 ( .A1(n26358), .A2(n32386), .Z(n33385) );
  INV_X1 U30522 ( .I(n21617), .ZN(n37033) );
  AOI22_X1 U30540 ( .A1(n122), .A2(n36910), .B1(n29218), .B2(n12691), .ZN(
        n33350) );
  NAND2_X2 U30549 ( .A1(n5258), .A2(n23523), .ZN(n23526) );
  XOR2_X1 U30552 ( .A1(n36880), .A2(n15398), .Z(n32154) );
  INV_X1 U30558 ( .I(n13374), .ZN(n1469) );
  XNOR2_X1 U30559 ( .A1(n13374), .A2(n27787), .ZN(n27748) );
  NAND2_X2 U30563 ( .A1(n18586), .A2(n15979), .ZN(n27358) );
  XOR2_X1 U30565 ( .A1(n5587), .A2(n36884), .Z(n29769) );
  XOR2_X1 U30566 ( .A1(n22758), .A2(n9205), .Z(n3529) );
  XOR2_X1 U30580 ( .A1(n10317), .A2(n10546), .Z(n10316) );
  INV_X4 U30581 ( .I(n36889), .ZN(n9231) );
  INV_X2 U30586 ( .I(n36890), .ZN(n30484) );
  XOR2_X1 U30587 ( .A1(n4967), .A2(n5743), .Z(n36890) );
  OAI21_X2 U30600 ( .A1(n24326), .A2(n13884), .B(n24390), .ZN(n36891) );
  OR2_X2 U30601 ( .A1(n21395), .A2(n21394), .Z(n17869) );
  OR2_X1 U30602 ( .A1(n25540), .A2(n30317), .Z(n16825) );
  NOR2_X2 U30603 ( .A1(n17800), .A2(n11614), .ZN(n36892) );
  NAND2_X1 U30604 ( .A1(n253), .A2(n30494), .ZN(n16884) );
  XOR2_X1 U30609 ( .A1(n17461), .A2(n36899), .Z(n22854) );
  XOR2_X1 U30610 ( .A1(n10939), .A2(n2234), .Z(n36899) );
  AOI22_X2 U30612 ( .A1(n23090), .A2(n19488), .B1(n15163), .B2(n23091), .ZN(
        n32025) );
  XOR2_X1 U30615 ( .A1(n8068), .A2(n8065), .Z(n8539) );
  OR2_X1 U30619 ( .A1(n24536), .A2(n33946), .Z(n25680) );
  XOR2_X1 U30620 ( .A1(n38905), .A2(n23914), .Z(n30502) );
  NAND3_X1 U30623 ( .A1(n37010), .A2(n39133), .A3(n15941), .ZN(n6521) );
  INV_X2 U30627 ( .I(n36909), .ZN(n18959) );
  XOR2_X1 U30628 ( .A1(Plaintext[175]), .A2(Key[175]), .Z(n36909) );
  INV_X2 U30629 ( .I(n33581), .ZN(n12435) );
  XOR2_X1 U30635 ( .A1(n37855), .A2(n10131), .Z(n36916) );
  NOR2_X1 U30636 ( .A1(n32696), .A2(n3605), .ZN(n32695) );
  XOR2_X1 U30640 ( .A1(n36919), .A2(n19799), .Z(Ciphertext[86]) );
  OR2_X1 U30641 ( .A1(n26058), .A2(n38416), .Z(n14573) );
  OAI21_X2 U30642 ( .A1(n34065), .A2(n12353), .B(n36923), .ZN(n21300) );
  NAND2_X2 U30643 ( .A1(n9394), .A2(n5414), .ZN(n36924) );
  INV_X2 U30645 ( .I(n28790), .ZN(n7288) );
  XOR2_X1 U30646 ( .A1(n6795), .A2(n36925), .Z(n6796) );
  XOR2_X1 U30647 ( .A1(n38816), .A2(n6847), .Z(n36925) );
  NAND3_X1 U30648 ( .A1(n30931), .A2(n18960), .A3(n28653), .ZN(n4523) );
  XOR2_X1 U30649 ( .A1(n22772), .A2(n11315), .Z(n11314) );
  XOR2_X1 U30650 ( .A1(n25313), .A2(n25312), .Z(n4273) );
  AOI22_X2 U30651 ( .A1(n7897), .A2(n36926), .B1(n8519), .B2(n7896), .ZN(n7895) );
  NAND2_X2 U30652 ( .A1(n1328), .A2(n22287), .ZN(n36926) );
  NOR2_X2 U30655 ( .A1(n36930), .A2(n17544), .ZN(n11568) );
  INV_X2 U30657 ( .I(n36932), .ZN(n6327) );
  XOR2_X1 U30661 ( .A1(n8400), .A2(n6360), .Z(n11451) );
  NAND2_X2 U30662 ( .A1(n3352), .A2(n2771), .ZN(n23069) );
  OAI21_X2 U30664 ( .A1(n36938), .A2(n31277), .B(n15251), .ZN(n27424) );
  OAI22_X2 U30666 ( .A1(n34077), .A2(n7440), .B1(n2439), .B2(n1031), .ZN(
        n23942) );
  NAND2_X1 U30669 ( .A1(n33894), .A2(n33609), .ZN(n23341) );
  AOI21_X2 U30671 ( .A1(n14203), .A2(n14205), .B(n24185), .ZN(n17351) );
  NAND2_X2 U30672 ( .A1(n6303), .A2(n23484), .ZN(n23306) );
  NOR2_X1 U30674 ( .A1(n9751), .A2(n19746), .ZN(n36940) );
  NOR2_X2 U30675 ( .A1(n26727), .A2(n13588), .ZN(n26774) );
  OAI21_X2 U30676 ( .A1(n14966), .A2(n1489), .B(n36942), .ZN(n14949) );
  INV_X1 U30678 ( .I(n28848), .ZN(n1178) );
  NOR2_X1 U30682 ( .A1(n4318), .A2(n22225), .ZN(n36946) );
  OAI22_X1 U30685 ( .A1(n21837), .A2(n8736), .B1(n690), .B2(n21435), .ZN(
        n14909) );
  NAND2_X1 U30689 ( .A1(n28562), .A2(n28563), .ZN(n28564) );
  NAND2_X2 U30690 ( .A1(n10640), .A2(n13484), .ZN(n6384) );
  XOR2_X1 U30693 ( .A1(n36959), .A2(n10748), .Z(n15883) );
  XOR2_X1 U30695 ( .A1(n29056), .A2(n29028), .Z(n12039) );
  NOR2_X2 U30696 ( .A1(n21370), .A2(n21369), .ZN(n31573) );
  XOR2_X1 U30697 ( .A1(n26473), .A2(n26472), .Z(n36961) );
  NOR2_X2 U30698 ( .A1(n4849), .A2(n344), .ZN(n20289) );
  XOR2_X1 U30699 ( .A1(n36962), .A2(n12228), .Z(n33144) );
  AND2_X1 U30703 ( .A1(n20660), .A2(n14453), .Z(n15668) );
  XOR2_X1 U30704 ( .A1(n27809), .A2(n10983), .Z(n10982) );
  OAI21_X2 U30709 ( .A1(n3012), .A2(n7075), .B(n36967), .ZN(n7901) );
  XOR2_X1 U30710 ( .A1(n31581), .A2(n23660), .Z(n8512) );
  OAI22_X1 U30713 ( .A1(n6851), .A2(n29421), .B1(n20018), .B2(n32946), .ZN(
        n36968) );
  XOR2_X1 U30715 ( .A1(n12411), .A2(n26145), .Z(n5737) );
  XNOR2_X1 U30718 ( .A1(n27855), .A2(n27607), .ZN(n27732) );
  NAND2_X2 U30719 ( .A1(n15772), .A2(n27453), .ZN(n27855) );
  NOR2_X1 U30720 ( .A1(n4116), .A2(n7935), .ZN(n21723) );
  NAND2_X2 U30723 ( .A1(n8595), .A2(n36974), .ZN(n3313) );
  NOR3_X1 U30724 ( .A1(n37378), .A2(n17791), .A3(n36798), .ZN(n15831) );
  NAND2_X2 U30727 ( .A1(n27068), .A2(n15120), .ZN(n27864) );
  XOR2_X1 U30730 ( .A1(n33132), .A2(n35900), .Z(n36980) );
  NAND2_X2 U30734 ( .A1(n36985), .A2(n18098), .ZN(n2) );
  NAND2_X2 U30735 ( .A1(n15015), .A2(n31194), .ZN(n36985) );
  NAND2_X2 U30736 ( .A1(n29270), .A2(n29271), .ZN(n19085) );
  NAND2_X1 U30738 ( .A1(n36216), .A2(n10104), .ZN(n13467) );
  XOR2_X1 U30744 ( .A1(n26393), .A2(n20212), .Z(n12622) );
  AOI22_X2 U30745 ( .A1(n29461), .A2(n29389), .B1(n17426), .B2(n19151), .ZN(
        n29402) );
  XOR2_X1 U30748 ( .A1(n17653), .A2(n31112), .Z(n24836) );
  INV_X2 U30749 ( .I(n24928), .ZN(n31112) );
  AOI22_X2 U30750 ( .A1(n24834), .A2(n1271), .B1(n24866), .B2(n13220), .ZN(
        n24928) );
  OAI21_X1 U30751 ( .A1(n3792), .A2(n3793), .B(n24733), .ZN(n4063) );
  NAND2_X2 U30755 ( .A1(n33929), .A2(n21424), .ZN(n4179) );
  OAI21_X2 U30757 ( .A1(n2668), .A2(n2671), .B(n9341), .ZN(n22443) );
  NAND3_X2 U30758 ( .A1(n32196), .A2(n1529), .A3(n35333), .ZN(n26218) );
  NAND3_X1 U30760 ( .A1(n29673), .A2(n19497), .A3(n20672), .ZN(n18944) );
  NAND2_X1 U30762 ( .A1(n16838), .A2(n1387), .ZN(n18431) );
  BUF_X2 U30766 ( .I(n22943), .Z(n36996) );
  NOR2_X1 U30767 ( .A1(n36998), .A2(n36997), .ZN(n16837) );
  INV_X1 U30768 ( .I(n8399), .ZN(n36998) );
  XOR2_X1 U30769 ( .A1(n33308), .A2(n31791), .Z(n36999) );
  NOR2_X1 U30773 ( .A1(n459), .A2(n1483), .ZN(n37002) );
  INV_X2 U30774 ( .I(n37003), .ZN(n6106) );
  XOR2_X1 U30775 ( .A1(n6109), .A2(n6107), .Z(n37003) );
  NAND2_X1 U30777 ( .A1(n2981), .A2(n2983), .ZN(n37006) );
  OR2_X2 U30778 ( .A1(n20897), .A2(n19167), .Z(n23121) );
  NAND2_X2 U30779 ( .A1(n37007), .A2(n25967), .ZN(n26516) );
  NOR2_X1 U30780 ( .A1(n25964), .A2(n25962), .ZN(n37008) );
  NAND2_X2 U30782 ( .A1(n528), .A2(n530), .ZN(n9611) );
  AOI22_X2 U30783 ( .A1(n27287), .A2(n27218), .B1(n31146), .B2(n30486), .ZN(
        n27564) );
  OAI21_X2 U30784 ( .A1(n34359), .A2(n1470), .B(n6013), .ZN(n27287) );
  NOR2_X1 U30787 ( .A1(n1297), .A2(n23468), .ZN(n37012) );
  INV_X2 U30788 ( .I(n37013), .ZN(n20616) );
  XNOR2_X1 U30789 ( .A1(n4140), .A2(n4141), .ZN(n37013) );
  NAND2_X2 U30791 ( .A1(n24571), .A2(n37017), .ZN(n13200) );
  AND2_X1 U30792 ( .A1(n3389), .A2(n37018), .Z(n5535) );
  XOR2_X1 U30793 ( .A1(n16833), .A2(n37019), .Z(n331) );
  XOR2_X1 U30794 ( .A1(n8704), .A2(n23980), .Z(n37019) );
  INV_X2 U30795 ( .I(n37020), .ZN(n37056) );
  XOR2_X1 U30796 ( .A1(n2757), .A2(n2758), .Z(n37020) );
  XOR2_X1 U30798 ( .A1(n30966), .A2(n14043), .Z(n14045) );
  AOI21_X2 U30804 ( .A1(n37026), .A2(n14082), .B(n7097), .ZN(n26086) );
  OR2_X1 U30805 ( .A1(n14257), .A2(n25642), .Z(n37026) );
  INV_X2 U30808 ( .I(n20616), .ZN(n32894) );
  NAND2_X2 U30809 ( .A1(n37027), .A2(n9313), .ZN(n9290) );
  OAI21_X2 U30810 ( .A1(n30369), .A2(n10236), .B(n18603), .ZN(n37027) );
  NAND3_X2 U30815 ( .A1(n13858), .A2(n13859), .A3(n13855), .ZN(n37030) );
  OR3_X1 U30816 ( .A1(n38159), .A2(n17751), .A3(n8944), .Z(n9745) );
  NAND3_X2 U30824 ( .A1(n14994), .A2(n14409), .A3(n31300), .ZN(n31918) );
  NAND2_X2 U30825 ( .A1(n20831), .A2(n21552), .ZN(n22349) );
  XOR2_X1 U30830 ( .A1(n37034), .A2(n12918), .Z(n9973) );
  NAND2_X2 U30833 ( .A1(n37036), .A2(n18822), .ZN(n18819) );
  OAI22_X2 U30834 ( .A1(n32740), .A2(n14994), .B1(n13946), .B2(n14439), .ZN(
        n37036) );
  XOR2_X1 U30838 ( .A1(n10837), .A2(n37038), .Z(n37037) );
  XOR2_X1 U30840 ( .A1(n5317), .A2(n5318), .Z(n12829) );
  OAI21_X2 U30842 ( .A1(n32837), .A2(n30288), .B(n27182), .ZN(n27746) );
  XOR2_X1 U30843 ( .A1(n11059), .A2(n10593), .Z(n10592) );
  NOR2_X1 U30845 ( .A1(n37039), .A2(n7175), .ZN(n19563) );
  BUF_X2 U30846 ( .I(n27417), .Z(n37040) );
  BUF_X2 U30847 ( .I(n7560), .Z(n37042) );
  XOR2_X1 U30848 ( .A1(n22517), .A2(n37660), .Z(n1868) );
  INV_X2 U30849 ( .I(n35469), .ZN(n274) );
  INV_X2 U30850 ( .I(n32191), .ZN(n1082) );
  INV_X2 U30853 ( .I(n32838), .ZN(n10659) );
  INV_X2 U30854 ( .I(n24316), .ZN(n24467) );
  XOR2_X1 U30855 ( .A1(n2107), .A2(n2104), .Z(n37047) );
  OAI21_X2 U30857 ( .A1(n13340), .A2(n32019), .B(n17453), .ZN(n31579) );
  OAI22_X2 U30858 ( .A1(n2746), .A2(n37202), .B1(n16541), .B2(n2745), .ZN(
        n31543) );
  XOR2_X1 U30859 ( .A1(n12830), .A2(n12833), .Z(n37048) );
  INV_X2 U30863 ( .I(n13877), .ZN(n12999) );
  INV_X1 U30867 ( .I(n29210), .ZN(n17121) );
  OAI21_X2 U30868 ( .A1(n15141), .A2(n15139), .B(n15138), .ZN(n29802) );
  NAND2_X2 U241 ( .A1(n2), .A2(n5543), .ZN(n6317) );
  INV_X2 U5878 ( .I(n8253), .ZN(n8385) );
  INV_X2 U1627 ( .I(n8173), .ZN(n32619) );
  INV_X2 U7284 ( .I(n668), .ZN(n21910) );
  NAND2_X2 U4261 ( .A1(n17118), .A2(n22177), .ZN(n22137) );
  INV_X2 U59 ( .I(n10118), .ZN(n1052) );
  NAND2_X2 U20202 ( .A1(n27266), .A2(n35990), .ZN(n20403) );
  OAI21_X2 U1704 ( .A1(n959), .A2(n33712), .B(n18238), .ZN(n33354) );
  NAND2_X2 U5464 ( .A1(n16579), .A2(n1843), .ZN(n1842) );
  NAND2_X2 U2347 ( .A1(n38629), .A2(n1419), .ZN(n28682) );
  INV_X2 U6509 ( .I(n22359), .ZN(n36337) );
  INV_X2 U10258 ( .I(n18429), .ZN(n4318) );
  INV_X2 U23027 ( .I(n20995), .ZN(n17047) );
  BUF_X4 U967 ( .I(n18983), .Z(n12159) );
  OAI22_X2 U17487 ( .A1(n2842), .A2(n2841), .B1(n1671), .B2(n22182), .ZN(n1745) );
  INV_X2 U5236 ( .I(n22897), .ZN(n1654) );
  NAND2_X2 U12157 ( .A1(n7724), .A2(n26134), .ZN(n3244) );
  NAND2_X2 U5990 ( .A1(n35779), .A2(n19053), .ZN(n12067) );
  INV_X2 U7621 ( .I(n30131), .ZN(n30144) );
  NAND2_X2 U2525 ( .A1(n36960), .A2(n35780), .ZN(n17813) );
  INV_X2 U6787 ( .I(n6291), .ZN(n5802) );
  BUF_X4 U6080 ( .I(n24140), .Z(n2439) );
  INV_X4 U1379 ( .I(n25867), .ZN(n5886) );
  NAND2_X2 U2394 ( .A1(n14130), .A2(n34013), .ZN(n22959) );
  INV_X2 U17116 ( .I(n24515), .ZN(n1270) );
  INV_X2 U22586 ( .I(n10679), .ZN(n29960) );
  OAI21_X2 U10169 ( .A1(n1778), .A2(n14028), .B(n14038), .ZN(n1777) );
  INV_X2 U1092 ( .I(n37593), .ZN(n34513) );
  INV_X4 U6911 ( .I(n14472), .ZN(n8070) );
  INV_X2 U4968 ( .I(n36913), .ZN(n7088) );
  INV_X2 U5911 ( .I(n26796), .ZN(n26734) );
  NAND3_X2 U28603 ( .A1(n978), .A2(n13508), .A3(n33100), .ZN(n12604) );
  OAI21_X2 U2367 ( .A1(n14130), .A2(n34013), .B(n17691), .ZN(n34715) );
  NAND2_X2 U8654 ( .A1(n20579), .A2(n20581), .ZN(n21980) );
  NOR2_X2 U1610 ( .A1(n12460), .A2(n31712), .ZN(n31711) );
  AOI21_X2 U3407 ( .A1(n27883), .A2(n28255), .B(n27885), .ZN(n10151) );
  INV_X2 U20427 ( .I(n7674), .ZN(n20372) );
  BUF_X4 U3791 ( .I(n6106), .Z(n32105) );
  NAND2_X2 U17987 ( .A1(n22402), .A2(n22183), .ZN(n22398) );
  NAND2_X2 U28416 ( .A1(n35429), .A2(n1047), .ZN(n22183) );
  INV_X2 U6937 ( .I(n20614), .ZN(n18831) );
  INV_X4 U16853 ( .I(n1276), .ZN(n24336) );
  INV_X2 U326 ( .I(n28250), .ZN(n13457) );
  NAND2_X2 U861 ( .A1(n20094), .A2(n26831), .ZN(n36507) );
  NOR2_X2 U4971 ( .A1(n13502), .A2(n19889), .ZN(n13501) );
  INV_X2 U23874 ( .I(n35901), .ZN(n15664) );
  INV_X2 U2138 ( .I(n23967), .ZN(n34451) );
  INV_X4 U7170 ( .I(n22935), .ZN(n1042) );
  BUF_X2 U4267 ( .I(n13989), .Z(n33516) );
  INV_X2 U15517 ( .I(n7810), .ZN(n8127) );
  NAND2_X2 U2172 ( .A1(n25337), .A2(n20052), .ZN(n25550) );
  INV_X2 U18960 ( .I(n6550), .ZN(n28159) );
  INV_X2 U1338 ( .I(n2047), .ZN(n1143) );
  INV_X2 U17145 ( .I(n29672), .ZN(n20672) );
  NAND2_X2 U3603 ( .A1(n1072), .A2(n34008), .ZN(n28108) );
  NOR2_X2 U1687 ( .A1(n3451), .A2(n25359), .ZN(n31900) );
  OAI21_X2 U7601 ( .A1(n29990), .A2(n3986), .B(n621), .ZN(n4011) );
  NAND2_X2 U1206 ( .A1(n19889), .A2(n11003), .ZN(n4852) );
  NAND2_X2 U7206 ( .A1(n26761), .A2(n26809), .ZN(n26653) );
  OAI21_X2 U22538 ( .A1(n19261), .A2(n22137), .B(n35802), .ZN(n5874) );
  INV_X4 U589 ( .I(n14408), .ZN(n1493) );
  INV_X2 U3542 ( .I(n23404), .ZN(n3366) );
  BUF_X2 U6276 ( .I(n13704), .Z(n35505) );
  INV_X2 U302 ( .I(n16108), .ZN(n15112) );
  NAND2_X2 U359 ( .A1(n28281), .A2(n37754), .ZN(n11280) );
  INV_X2 U20032 ( .I(n32010), .ZN(n33937) );
  INV_X2 U28095 ( .I(n27745), .ZN(n27535) );
  NAND2_X2 U7386 ( .A1(n9217), .A2(n13495), .ZN(n6409) );
  BUF_X4 U5213 ( .I(n2319), .Z(n35062) );
  INV_X2 U18781 ( .I(n5960), .ZN(n9147) );
  NAND2_X2 U729 ( .A1(n26870), .A2(n7973), .ZN(n27007) );
  OAI21_X2 U18464 ( .A1(n12146), .A2(n10008), .B(n33104), .ZN(n31759) );
  INV_X2 U141 ( .I(n34179), .ZN(n30052) );
  INV_X2 U653 ( .I(n4815), .ZN(n21149) );
  NAND2_X2 U29506 ( .A1(n7635), .A2(n28023), .ZN(n27918) );
  INV_X4 U5757 ( .I(n11003), .ZN(n927) );
  INV_X2 U3026 ( .I(n17529), .ZN(n1671) );
  INV_X4 U30812 ( .I(n31994), .ZN(n37028) );
  INV_X2 U3834 ( .I(n34526), .ZN(n24708) );
  INV_X2 U5877 ( .I(n16627), .ZN(n35722) );
  AOI22_X2 U18045 ( .A1(n17309), .A2(n32385), .B1(n11980), .B2(n38694), .ZN(
        n35212) );
  INV_X2 U3923 ( .I(n24317), .ZN(n17546) );
  INV_X2 U13744 ( .I(n692), .ZN(n25999) );
  NOR2_X1 U11009 ( .A1(n32497), .A2(n35720), .ZN(n18218) );
  INV_X2 U5270 ( .I(n24285), .ZN(n24119) );
  INV_X4 U6679 ( .I(n22682), .ZN(n22856) );
  BUF_X4 U1384 ( .I(n18987), .Z(n596) );
  NOR2_X2 U9089 ( .A1(n33669), .A2(n39132), .ZN(n2614) );
  NOR2_X2 U2391 ( .A1(n1045), .A2(n20173), .ZN(n35863) );
  BUF_X4 U5605 ( .I(n12667), .Z(n6131) );
  INV_X2 U4655 ( .I(n9165), .ZN(n10681) );
  NAND2_X2 U5742 ( .A1(n27011), .A2(n31875), .ZN(n10357) );
  NAND2_X1 U28849 ( .A1(n4239), .A2(n22390), .ZN(n36616) );
  INV_X2 U22096 ( .I(n9958), .ZN(n12302) );
  INV_X4 U2254 ( .I(n11033), .ZN(n930) );
  INV_X4 U3343 ( .I(n217), .ZN(n5702) );
  BUF_X2 U7714 ( .I(n3014), .Z(n33841) );
  NOR2_X2 U22616 ( .A1(n32542), .A2(n20732), .ZN(n8925) );
  NOR2_X2 U2242 ( .A1(n217), .A2(n7160), .ZN(n22932) );
  INV_X2 U19626 ( .I(n7133), .ZN(n26244) );
  INV_X2 U2369 ( .I(n25337), .ZN(n25460) );
  NOR2_X1 U10213 ( .A1(n16432), .A2(n34382), .ZN(n6104) );
  OAI21_X2 U6587 ( .A1(n38555), .A2(n31383), .B(n21995), .ZN(n20089) );
  NOR2_X2 U1721 ( .A1(n31698), .A2(n18148), .ZN(n20038) );
  NOR2_X2 U1080 ( .A1(n26056), .A2(n9743), .ZN(n15703) );
  OAI22_X2 U17473 ( .A1(n39576), .A2(n16468), .B1(n1057), .B2(n30051), .ZN(
        n7166) );
  NAND2_X2 U3191 ( .A1(n9363), .A2(n24707), .ZN(n34192) );
  NOR2_X2 U12702 ( .A1(n33986), .A2(n34526), .ZN(n9363) );
  NAND2_X2 U12056 ( .A1(n9326), .A2(n19241), .ZN(n1849) );
  NOR2_X2 U5051 ( .A1(n37072), .A2(n39454), .ZN(n9326) );
  INV_X2 U652 ( .I(n8402), .ZN(n8302) );
  INV_X4 U28451 ( .I(n34562), .ZN(n33369) );
  NOR2_X2 U12405 ( .A1(n6894), .A2(n560), .ZN(n21136) );
  INV_X2 U650 ( .I(n27825), .ZN(n1463) );
  NAND2_X2 U238 ( .A1(n10587), .A2(n9648), .ZN(n33724) );
  OAI21_X2 U5564 ( .A1(n20134), .A2(n20612), .B(n34417), .ZN(n16643) );
  NAND2_X2 U4895 ( .A1(n19546), .A2(n32138), .ZN(n12751) );
  INV_X2 U17390 ( .I(n5921), .ZN(n17708) );
  NOR2_X2 U5702 ( .A1(n39085), .A2(n1027), .ZN(n11199) );
  INV_X2 U2048 ( .I(n690), .ZN(n1158) );
  BUF_X4 U4150 ( .I(n8742), .Z(n557) );
  AOI22_X2 U17960 ( .A1(n21449), .A2(n1342), .B1(n32817), .B2(n22173), .ZN(
        n21453) );
  NOR2_X2 U2310 ( .A1(n12946), .A2(n20696), .ZN(n31123) );
  OR2_X1 U3897 ( .A1(n10896), .A2(n31596), .Z(n10870) );
  NAND2_X2 U16641 ( .A1(n28238), .A2(n1453), .ZN(n4150) );
  INV_X2 U17288 ( .I(n16054), .ZN(n3395) );
  NAND2_X2 U8624 ( .A1(n9242), .A2(n31971), .ZN(n2604) );
  NOR2_X2 U1120 ( .A1(n32157), .A2(n32156), .ZN(n34883) );
  NAND2_X2 U18281 ( .A1(n18062), .A2(n25801), .ZN(n25903) );
  INV_X2 U17589 ( .I(n30894), .ZN(n89) );
  NAND2_X2 U17232 ( .A1(n29986), .A2(n16468), .ZN(n6602) );
  NAND2_X2 U6855 ( .A1(n24337), .A2(n14558), .ZN(n7811) );
  INV_X2 U600 ( .I(n27730), .ZN(n27833) );
  AND2_X2 U17064 ( .A1(n889), .A2(n13492), .Z(n14642) );
  BUF_X2 U3387 ( .I(n17425), .Z(n15089) );
  INV_X2 U3233 ( .I(n19260), .ZN(n29525) );
  INV_X2 U2112 ( .I(n36272), .ZN(n14558) );
  AOI21_X2 U464 ( .A1(n35846), .A2(n16851), .B(n4152), .ZN(n12466) );
  NOR2_X2 U19587 ( .A1(n1650), .A2(n9472), .ZN(n5215) );
  NAND2_X2 U3424 ( .A1(n6161), .A2(n32617), .ZN(n6732) );
  INV_X4 U5846 ( .I(n25498), .ZN(n25379) );
  AOI21_X2 U18651 ( .A1(n21996), .A2(n3687), .B(n22071), .ZN(n16028) );
  INV_X4 U7232 ( .I(n11149), .ZN(n22267) );
  INV_X4 U1888 ( .I(n6944), .ZN(n24723) );
  INV_X2 U26225 ( .I(n32080), .ZN(n20572) );
  NAND2_X2 U1256 ( .A1(n37151), .A2(n26008), .ZN(n20049) );
  OAI21_X2 U9258 ( .A1(n3224), .A2(n11130), .B(n33858), .ZN(n3095) );
  INV_X4 U5583 ( .I(n29598), .ZN(n1404) );
  INV_X2 U7182 ( .I(n57), .ZN(n14304) );
  INV_X4 U5821 ( .I(n32617), .ZN(n21762) );
  NAND2_X2 U13678 ( .A1(n17635), .A2(n22107), .ZN(n17634) );
  AOI21_X2 U4236 ( .A1(n15715), .A2(n33061), .B(n38527), .ZN(n15713) );
  INV_X2 U13781 ( .I(n7768), .ZN(n8621) );
  INV_X4 U8954 ( .I(n33384), .ZN(n30694) );
  AND2_X1 U4001 ( .A1(n11562), .A2(n26269), .Z(n854) );
  OAI21_X2 U24461 ( .A1(n18734), .A2(n4664), .B(n32419), .ZN(n16809) );
  NOR2_X2 U6750 ( .A1(n23528), .A2(n36539), .ZN(n23529) );
  INV_X2 U4277 ( .I(n24337), .ZN(n8174) );
  INV_X2 U608 ( .I(n28219), .ZN(n36860) );
  INV_X2 U11367 ( .I(n28141), .ZN(n28142) );
  INV_X2 U4175 ( .I(n14463), .ZN(n10477) );
  INV_X2 U1717 ( .I(n25194), .ZN(n2318) );
  INV_X2 U3806 ( .I(n3313), .ZN(n992) );
  INV_X1 U9200 ( .I(n1472), .ZN(n3088) );
  AOI21_X2 U18104 ( .A1(n31680), .A2(n16480), .B(n16479), .ZN(n6110) );
  AOI22_X1 U10313 ( .A1(n21756), .A2(n11916), .B1(n11917), .B2(n11918), .ZN(
        n10324) );
  INV_X2 U9128 ( .I(n28153), .ZN(n1203) );
  INV_X2 U177 ( .I(n29642), .ZN(n35571) );
  INV_X1 U12780 ( .I(n16502), .ZN(n1581) );
  INV_X4 U2120 ( .I(n1589), .ZN(n2396) );
  NAND2_X2 U3264 ( .A1(n29981), .A2(n29968), .ZN(n29971) );
  INV_X2 U6363 ( .I(n20408), .ZN(n5907) );
  BUF_X4 U4208 ( .I(n28807), .Z(n33577) );
  INV_X2 U1099 ( .I(n801), .ZN(n24267) );
  AOI22_X2 U6925 ( .A1(n24084), .A2(n24853), .B1(n24855), .B2(n32064), .ZN(
        n24085) );
  INV_X2 U5747 ( .I(n23464), .ZN(n23238) );
  NAND2_X2 U17203 ( .A1(n35960), .A2(n24637), .ZN(n20414) );
  OAI22_X2 U13900 ( .A1(n21605), .A2(n16128), .B1(n21944), .B2(n19133), .ZN(
        n11302) );
  AOI22_X2 U2363 ( .A1(n22863), .A2(n1650), .B1(n1651), .B2(n6385), .ZN(n4160)
         );
  INV_X2 U79 ( .I(n31428), .ZN(n3693) );
  AOI21_X2 U857 ( .A1(n17785), .A2(n11513), .B(n35877), .ZN(n36520) );
  OAI21_X2 U1736 ( .A1(n11271), .A2(n37106), .B(n11082), .ZN(n13494) );
  NOR2_X2 U14416 ( .A1(n37137), .A2(n20625), .ZN(n31465) );
  NOR2_X2 U14439 ( .A1(n948), .A2(n26660), .ZN(n31264) );
  INV_X4 U3419 ( .I(n35377), .ZN(n21130) );
  INV_X2 U11532 ( .I(n30959), .ZN(n28168) );
  INV_X2 U6368 ( .I(n8765), .ZN(n962) );
  INV_X2 U2518 ( .I(n22335), .ZN(n36632) );
  INV_X2 U27619 ( .I(n19458), .ZN(n29998) );
  NOR2_X2 U21142 ( .A1(n8818), .A2(n18261), .ZN(n28111) );
  NAND2_X2 U9685 ( .A1(n9584), .A2(n34620), .ZN(n9580) );
  BUF_X4 U5741 ( .I(n5126), .Z(n31827) );
  OAI21_X2 U1604 ( .A1(n4625), .A2(n2149), .B(n34636), .ZN(n7695) );
  INV_X4 U3466 ( .I(n1275), .ZN(n9101) );
  OAI22_X1 U10220 ( .A1(n22889), .A2(n19469), .B1(n5656), .B2(n23125), .ZN(
        n34713) );
  INV_X2 U676 ( .I(n27595), .ZN(n31163) );
  NAND2_X2 U1432 ( .A1(n1048), .A2(n22108), .ZN(n22107) );
  INV_X2 U203 ( .I(n20006), .ZN(n11721) );
  NOR2_X2 U1615 ( .A1(n25327), .A2(n37237), .ZN(n18786) );
  NAND2_X2 U18361 ( .A1(n32902), .A2(n28377), .ZN(n9111) );
  CLKBUF_X4 U6087 ( .I(n23992), .Z(n24443) );
  INV_X2 U15189 ( .I(n13193), .ZN(n24018) );
  INV_X2 U5798 ( .I(n22122), .ZN(n22266) );
  AOI21_X2 U6996 ( .A1(n2057), .A2(n7210), .B(n20989), .ZN(n20988) );
  AOI22_X2 U2922 ( .A1(n38851), .A2(n19538), .B1(n1314), .B2(n14725), .ZN(
        n33706) );
  NAND2_X2 U1628 ( .A1(n37238), .A2(n5798), .ZN(n34636) );
  INV_X4 U7856 ( .I(n2532), .ZN(n21751) );
  INV_X2 U13217 ( .I(n23365), .ZN(n1953) );
  INV_X2 U11385 ( .I(n35895), .ZN(n32961) );
  INV_X2 U20655 ( .I(n32151), .ZN(n3969) );
  INV_X4 U8715 ( .I(n18205), .ZN(n21788) );
  NOR2_X2 U4466 ( .A1(n27326), .A2(n39216), .ZN(n8763) );
  INV_X4 U4911 ( .I(n12443), .ZN(n28103) );
  NAND2_X2 U4215 ( .A1(n7552), .A2(n39681), .ZN(n11126) );
  OR2_X1 U3875 ( .A1(n31558), .A2(n7584), .Z(n23161) );
  INV_X2 U3133 ( .I(n20372), .ZN(n23082) );
  OAI21_X2 U13650 ( .A1(n37189), .A2(n14823), .B(n9715), .ZN(n14822) );
  NOR2_X2 U13530 ( .A1(n35586), .A2(n19870), .ZN(n4099) );
  OAI21_X2 U27421 ( .A1(n1625), .A2(n6217), .B(n23528), .ZN(n23283) );
  INV_X4 U877 ( .I(n21254), .ZN(n954) );
  OAI21_X2 U2106 ( .A1(n4993), .A2(n19837), .B(n18163), .ZN(n33487) );
  NAND2_X2 U7027 ( .A1(n955), .A2(n15541), .ZN(n25452) );
  INV_X2 U15586 ( .I(n24427), .ZN(n19070) );
  OAI21_X2 U7035 ( .A1(n32085), .A2(n560), .B(n17353), .ZN(n5355) );
  AND2_X2 U1055 ( .A1(n36283), .A2(n12682), .Z(n26955) );
  INV_X2 U3812 ( .I(n20087), .ZN(n344) );
  INV_X2 U6938 ( .I(n6106), .ZN(n14708) );
  NAND2_X2 U2233 ( .A1(n35545), .A2(n39316), .ZN(n9011) );
  INV_X2 U6128 ( .I(n3779), .ZN(n4152) );
  OAI22_X2 U2968 ( .A1(n6181), .A2(n1390), .B1(n29662), .B2(n39689), .ZN(
        n29665) );
  OAI21_X2 U2523 ( .A1(n5945), .A2(n1989), .B(n5944), .ZN(n4328) );
  INV_X2 U6300 ( .I(n22038), .ZN(n34216) );
  INV_X2 U344 ( .I(n28717), .ZN(n35491) );
  INV_X2 U25211 ( .I(n25557), .ZN(n17281) );
  OAI21_X2 U7051 ( .A1(n38531), .A2(n31310), .B(n1524), .ZN(n35956) );
  NOR2_X2 U51 ( .A1(n3818), .A2(n30076), .ZN(n30066) );
  AOI22_X2 U29543 ( .A1(n6534), .A2(n36911), .B1(n39632), .B2(n7542), .ZN(
        n3920) );
  NOR2_X2 U3384 ( .A1(n20498), .A2(n17730), .ZN(n29717) );
  NOR2_X2 U1696 ( .A1(n9781), .A2(n18077), .ZN(n35748) );
  INV_X2 U3414 ( .I(n34120), .ZN(n17477) );
  AOI22_X2 U319 ( .A1(n18910), .A2(n6932), .B1(n28651), .B2(n11120), .ZN(
        n28389) );
  NAND2_X2 U5475 ( .A1(n22038), .A2(n21802), .ZN(n22076) );
  NAND2_X2 U4805 ( .A1(n13114), .A2(n1284), .ZN(n13113) );
  NAND2_X2 U4580 ( .A1(n39401), .A2(n23426), .ZN(n31787) );
  NOR2_X2 U1473 ( .A1(n1346), .A2(n11703), .ZN(n35) );
  INV_X2 U5994 ( .I(n4862), .ZN(n21143) );
  INV_X2 U7569 ( .I(n29761), .ZN(n30747) );
  INV_X2 U5472 ( .I(n28339), .ZN(n34007) );
  NAND2_X2 U7356 ( .A1(n1227), .A2(n3313), .ZN(n11140) );
  INV_X2 U428 ( .I(n19631), .ZN(n32338) );
  NAND2_X2 U430 ( .A1(n13601), .A2(n28728), .ZN(n15752) );
  INV_X4 U5724 ( .I(n13555), .ZN(n7086) );
  BUF_X4 U7444 ( .I(n28033), .Z(n37) );
  NAND2_X2 U2953 ( .A1(n5430), .A2(n28272), .ZN(n31027) );
  NOR2_X2 U19589 ( .A1(n32926), .A2(n33593), .ZN(n27245) );
  INV_X2 U2441 ( .I(n13352), .ZN(n23124) );
  INV_X2 U5809 ( .I(n11703), .ZN(n9288) );
  AOI21_X2 U3944 ( .A1(n25690), .A2(n14481), .B(n19963), .ZN(n25687) );
  NAND2_X2 U4159 ( .A1(n38610), .A2(n29040), .ZN(n15733) );
  AOI21_X2 U4253 ( .A1(n2927), .A2(n39266), .B(n12699), .ZN(n12698) );
  NOR2_X2 U626 ( .A1(n1070), .A2(n1448), .ZN(n4375) );
  BUF_X2 U3680 ( .I(n29456), .Z(n19065) );
  NAND3_X1 U19672 ( .A1(n1893), .A2(n1894), .A3(n17521), .ZN(n445) );
  NAND2_X2 U1312 ( .A1(n30443), .A2(n11658), .ZN(n23100) );
  OAI21_X2 U10327 ( .A1(n21810), .A2(n13472), .B(n2166), .ZN(n21566) );
  AOI21_X2 U2404 ( .A1(n22303), .A2(n22076), .B(n33886), .ZN(n14363) );
  INV_X2 U4953 ( .I(n14601), .ZN(n34004) );
  INV_X2 U1139 ( .I(n15679), .ZN(n20317) );
  NAND2_X2 U30862 ( .A1(n26863), .A2(n1230), .ZN(n37055) );
  INV_X2 U6872 ( .I(n5897), .ZN(n6273) );
  INV_X2 U14903 ( .I(n20416), .ZN(n25716) );
  NOR2_X2 U791 ( .A1(n27213), .A2(n16043), .ZN(n27214) );
  NAND2_X2 U1909 ( .A1(n24784), .A2(n32898), .ZN(n24875) );
  NAND2_X2 U5315 ( .A1(n37227), .A2(n17709), .ZN(n19028) );
  NAND2_X2 U16552 ( .A1(n3694), .A2(n15996), .ZN(n15822) );
  NOR2_X1 U14240 ( .A1(n34821), .A2(n15735), .ZN(n18715) );
  AND2_X2 U2027 ( .A1(n8151), .A2(n11643), .Z(n22870) );
  OR2_X2 U4819 ( .A1(n35252), .A2(n20087), .Z(n29581) );
  NOR2_X2 U2614 ( .A1(n21412), .A2(n21475), .ZN(n21564) );
  INV_X2 U7815 ( .I(n35287), .ZN(n27410) );
  AND2_X2 U13447 ( .A1(n32855), .A2(n21767), .Z(n21766) );
  AOI22_X2 U15198 ( .A1(n27990), .A2(n28103), .B1(n27991), .B2(n2740), .ZN(
        n27993) );
  NAND2_X2 U4152 ( .A1(n28394), .A2(n28395), .ZN(n33574) );
  NOR2_X2 U8429 ( .A1(n14088), .A2(n30659), .ZN(n9140) );
  INV_X4 U1334 ( .I(n21132), .ZN(n3803) );
  INV_X2 U24379 ( .I(n22796), .ZN(n18750) );
  INV_X2 U22261 ( .I(n10111), .ZN(n14394) );
  AOI21_X2 U1269 ( .A1(n26081), .A2(n13869), .B(n10724), .ZN(n30659) );
  NAND2_X2 U20968 ( .A1(n7494), .A2(n7612), .ZN(n27037) );
  NAND2_X2 U9845 ( .A1(n23331), .A2(n23636), .ZN(n3264) );
  INV_X4 U6085 ( .I(n17240), .ZN(n971) );
  INV_X2 U4590 ( .I(n24802), .ZN(n34354) );
  INV_X2 U9574 ( .I(n14045), .ZN(n1252) );
  INV_X1 U21057 ( .I(n8517), .ZN(n21839) );
  NAND2_X2 U2348 ( .A1(n12696), .A2(n10299), .ZN(n35441) );
  OAI22_X2 U18313 ( .A1(n3930), .A2(n11364), .B1(n31383), .B2(n22328), .ZN(
        n8503) );
  NOR2_X2 U10176 ( .A1(n13163), .A2(n22326), .ZN(n8504) );
  INV_X4 U30215 ( .I(n18619), .ZN(n24395) );
  NOR2_X2 U1826 ( .A1(n4225), .A2(n1566), .ZN(n18063) );
  AOI21_X2 U19371 ( .A1(n7535), .A2(n6969), .B(n5487), .ZN(n23244) );
  INV_X2 U16955 ( .I(n28159), .ZN(n19541) );
  INV_X4 U3078 ( .I(n15153), .ZN(n5669) );
  NOR2_X2 U8410 ( .A1(n31234), .A2(n34307), .ZN(n19119) );
  NAND2_X2 U555 ( .A1(n37056), .A2(n28153), .ZN(n28420) );
  NAND2_X2 U3431 ( .A1(n2639), .A2(n8476), .ZN(n28369) );
  NOR2_X1 U4825 ( .A1(n4126), .A2(n30878), .ZN(n30877) );
  INV_X2 U178 ( .I(n5977), .ZN(n29632) );
  INV_X2 U595 ( .I(n17934), .ZN(n26660) );
  NAND2_X2 U18103 ( .A1(n20039), .A2(n35813), .ZN(n24872) );
  INV_X2 U325 ( .I(n32682), .ZN(n34861) );
  INV_X4 U8003 ( .I(n9242), .ZN(n28278) );
  NAND3_X2 U2329 ( .A1(n35208), .A2(n13823), .A3(n37248), .ZN(n13818) );
  CLKBUF_X2 U6054 ( .I(Key[64]), .Z(n19583) );
  NAND2_X1 U27621 ( .A1(n9444), .A2(n28504), .ZN(n28507) );
  NAND2_X2 U17464 ( .A1(n6602), .A2(n39576), .ZN(n454) );
  OAI21_X2 U30129 ( .A1(n15568), .A2(n15569), .B(n28229), .ZN(n33620) );
  AOI21_X2 U5501 ( .A1(n35694), .A2(n16576), .B(n1203), .ZN(n10466) );
  INV_X2 U24952 ( .I(n4120), .ZN(n32902) );
  BUF_X2 U6367 ( .I(n22796), .Z(n23128) );
  INV_X1 U16980 ( .I(n38228), .ZN(n27576) );
  OAI21_X2 U17212 ( .A1(n6160), .A2(n31275), .B(n31785), .ZN(n31554) );
  INV_X2 U1389 ( .I(n36666), .ZN(n34745) );
  INV_X2 U17370 ( .I(n35151), .ZN(n26112) );
  NAND2_X1 U9383 ( .A1(n17213), .A2(n25939), .ZN(n13525) );
  NOR2_X2 U37 ( .A1(n18384), .A2(n29534), .ZN(n29519) );
  AOI22_X2 U3236 ( .A1(n26775), .A2(n26866), .B1(n20004), .B2(n26774), .ZN(
        n30617) );
  BUF_X4 U4350 ( .I(n14401), .Z(n1109) );
  INV_X2 U14216 ( .I(n19559), .ZN(n23602) );
  OAI21_X2 U3710 ( .A1(n20396), .A2(n21310), .B(n1126), .ZN(n24135) );
  OR2_X2 U5504 ( .A1(n16382), .A2(n13062), .Z(n14271) );
  NAND2_X2 U17520 ( .A1(n29341), .A2(n29336), .ZN(n29333) );
  INV_X4 U4290 ( .I(n34717), .ZN(n1217) );
  INV_X2 U30362 ( .I(n19515), .ZN(n33782) );
  INV_X2 U171 ( .I(n15270), .ZN(n15271) );
  NAND2_X2 U1565 ( .A1(n13516), .A2(n19886), .ZN(n12161) );
  NOR2_X2 U1025 ( .A1(n26920), .A2(n26922), .ZN(n35629) );
  INV_X2 U9803 ( .I(n9458), .ZN(n1275) );
  NAND2_X2 U25808 ( .A1(n9514), .A2(n759), .ZN(n15334) );
  NAND2_X2 U2943 ( .A1(n19728), .A2(n8527), .ZN(n2158) );
  INV_X2 U25872 ( .I(n39528), .ZN(n15448) );
  INV_X4 U2578 ( .I(n22294), .ZN(n22246) );
  NAND2_X2 U5807 ( .A1(n14083), .A2(n25642), .ZN(n34465) );
  NOR2_X2 U25074 ( .A1(n16140), .A2(n35290), .ZN(n15890) );
  INV_X4 U3851 ( .I(n22899), .ZN(n22849) );
  NAND2_X1 U25188 ( .A1(n14657), .A2(n24775), .ZN(n17971) );
  INV_X4 U598 ( .I(n15594), .ZN(n26354) );
  OAI21_X2 U16592 ( .A1(n36095), .A2(n22915), .B(n19293), .ZN(n4102) );
  NOR2_X2 U2296 ( .A1(n35377), .A2(n31944), .ZN(n2633) );
  BUF_X4 U17752 ( .I(n20156), .Z(n7251) );
  NAND2_X2 U11629 ( .A1(n26790), .A2(n4781), .ZN(n12352) );
  OAI21_X2 U9121 ( .A1(n13366), .A2(n14480), .B(n17447), .ZN(n11408) );
  NAND2_X2 U17830 ( .A1(n8735), .A2(n16366), .ZN(n35782) );
  NAND2_X1 U1516 ( .A1(n7696), .A2(n21868), .ZN(n12332) );
  NOR2_X2 U221 ( .A1(n35173), .A2(n28356), .ZN(n28535) );
  INV_X2 U2463 ( .I(n35859), .ZN(n11307) );
  AOI21_X2 U26558 ( .A1(n13339), .A2(n15272), .B(n20782), .ZN(n33135) );
  INV_X2 U2429 ( .I(n23085), .ZN(n20230) );
  INV_X2 U2414 ( .I(n29792), .ZN(n29782) );
  INV_X2 U6027 ( .I(n22197), .ZN(n1687) );
  AOI21_X2 U17715 ( .A1(n28649), .A2(n29494), .B(n29420), .ZN(n18725) );
  OAI21_X2 U25963 ( .A1(n5653), .A2(n5210), .B(n24909), .ZN(n5209) );
  INV_X2 U1381 ( .I(n11308), .ZN(n11315) );
  NOR2_X2 U26557 ( .A1(n14079), .A2(n17034), .ZN(n26662) );
  OAI21_X2 U7539 ( .A1(n8658), .A2(n8657), .B(n1066), .ZN(n8656) );
  OAI22_X2 U3591 ( .A1(n24136), .A2(n24086), .B1(n24309), .B2(n7730), .ZN(
        n11630) );
  NAND2_X2 U13880 ( .A1(n9539), .A2(n21854), .ZN(n6270) );
  OAI21_X2 U10197 ( .A1(n9546), .A2(n38246), .B(n7916), .ZN(n19011) );
  BUF_X2 U10892 ( .I(n16009), .Z(n4849) );
  INV_X2 U5955 ( .I(n524), .ZN(n35088) );
  AOI21_X2 U28586 ( .A1(n23010), .A2(n23009), .B(n23308), .ZN(n23016) );
  NAND2_X2 U165 ( .A1(n35571), .A2(n19962), .ZN(n7373) );
  NAND2_X2 U1910 ( .A1(n17087), .A2(n24623), .ZN(n35693) );
  NAND2_X2 U4585 ( .A1(n10143), .A2(n39401), .ZN(n31164) );
  INV_X4 U13563 ( .I(n17692), .ZN(n14130) );
  OAI21_X2 U627 ( .A1(n944), .A2(n1475), .B(n19662), .ZN(n31498) );
  OAI21_X2 U2212 ( .A1(n13489), .A2(n12236), .B(n37289), .ZN(n13488) );
  AOI21_X2 U4763 ( .A1(n38283), .A2(n19645), .B(n19469), .ZN(n15627) );
  INV_X4 U1070 ( .I(n1607), .ZN(n24330) );
  OAI22_X2 U10308 ( .A1(n21635), .A2(n32138), .B1(n12754), .B2(n21944), .ZN(
        n11303) );
  INV_X2 U1445 ( .I(n21802), .ZN(n22073) );
  NAND3_X2 U17386 ( .A1(n13294), .A2(n8262), .A3(n5101), .ZN(n27242) );
  NOR2_X2 U6392 ( .A1(n20034), .A2(n39284), .ZN(n9485) );
  NAND2_X2 U15413 ( .A1(n24076), .A2(n23911), .ZN(n7114) );
  INV_X2 U10141 ( .I(n33510), .ZN(n36517) );
  BUF_X4 U18633 ( .I(n11562), .Z(n948) );
  INV_X2 U761 ( .I(n16736), .ZN(n944) );
  OAI21_X2 U16132 ( .A1(n36461), .A2(n30775), .B(n6583), .ZN(n24056) );
  AOI21_X2 U2488 ( .A1(n22359), .A2(n22358), .B(n31939), .ZN(n14801) );
  INV_X2 U13069 ( .I(n19188), .ZN(n8884) );
  AOI21_X2 U16788 ( .A1(n7404), .A2(n36922), .B(n34402), .ZN(n14722) );
  OAI21_X2 U13846 ( .A1(n19553), .A2(n39672), .B(n19552), .ZN(n21686) );
  INV_X2 U6399 ( .I(n22041), .ZN(n17530) );
  AND2_X1 U18840 ( .A1(n16039), .A2(n15370), .Z(n11900) );
  NOR2_X2 U2586 ( .A1(n31480), .A2(n6102), .ZN(n6099) );
  INV_X2 U26196 ( .I(n14481), .ZN(n19813) );
  INV_X2 U27605 ( .I(n10231), .ZN(n26645) );
  INV_X4 U7712 ( .I(n33957), .ZN(n12784) );
  INV_X2 U6160 ( .I(n35191), .ZN(n1634) );
  NAND2_X2 U5901 ( .A1(n28698), .A2(n28696), .ZN(n28366) );
  BUF_X4 U16229 ( .I(n33736), .Z(n31504) );
  NOR2_X2 U12420 ( .A1(n23389), .A2(n38408), .ZN(n20450) );
  BUF_X2 U24220 ( .I(n15463), .Z(n32815) );
  CLKBUF_X4 U2294 ( .I(n39401), .Z(n36885) );
  INV_X2 U9933 ( .I(n18866), .ZN(n23404) );
  NAND3_X2 U282 ( .A1(n28213), .A2(n28212), .A3(n16869), .ZN(n28352) );
  INV_X2 U6782 ( .I(n10370), .ZN(n5699) );
  INV_X2 U14110 ( .I(n13966), .ZN(n31198) );
  INV_X2 U31 ( .I(n11067), .ZN(n13804) );
  NAND2_X2 U675 ( .A1(n17994), .A2(n25954), .ZN(n9589) );
  NOR2_X2 U7443 ( .A1(n1446), .A2(n8368), .ZN(n14585) );
  OAI21_X2 U11624 ( .A1(n27391), .A2(n27035), .B(n27200), .ZN(n27036) );
  NAND3_X2 U1420 ( .A1(n25697), .A2(n25698), .A3(n32654), .ZN(n32615) );
  NAND2_X2 U6608 ( .A1(n5616), .A2(n5618), .ZN(n34259) );
  NAND2_X2 U18277 ( .A1(n2340), .A2(n15136), .ZN(n31723) );
  INV_X4 U14576 ( .I(n2153), .ZN(n22262) );
  INV_X2 U26313 ( .I(n22247), .ZN(n16140) );
  BUF_X4 U8237 ( .I(n3441), .Z(n2747) );
  AOI21_X2 U1469 ( .A1(n10044), .A2(n21693), .B(n8971), .ZN(n21494) );
  NAND2_X2 U6672 ( .A1(n22129), .A2(n8245), .ZN(n16463) );
  OAI21_X2 U1137 ( .A1(n25764), .A2(n10724), .B(n25989), .ZN(n4801) );
  INV_X2 U7164 ( .I(n15290), .ZN(n6647) );
  INV_X2 U19558 ( .I(n13880), .ZN(n975) );
  NAND2_X2 U17979 ( .A1(n16115), .A2(n33845), .ZN(n18673) );
  NOR2_X2 U1647 ( .A1(n34689), .A2(n32131), .ZN(n18438) );
  AOI22_X2 U17873 ( .A1(n31326), .A2(n29990), .B1(n30045), .B2(n4011), .ZN(
        n35234) );
  NAND3_X2 U3278 ( .A1(n98), .A2(n9346), .A3(n23413), .ZN(n36927) );
  INV_X2 U21040 ( .I(n36075), .ZN(n10199) );
  NAND2_X2 U151 ( .A1(n37100), .A2(n14422), .ZN(n29449) );
  AOI22_X2 U3626 ( .A1(n14249), .A2(n33086), .B1(n14250), .B2(n14139), .ZN(
        n14248) );
  INV_X2 U18355 ( .I(n36623), .ZN(n17714) );
  OAI21_X2 U3241 ( .A1(n32802), .A2(n39537), .B(n17343), .ZN(n20959) );
  NAND2_X2 U13554 ( .A1(n23166), .A2(n22973), .ZN(n23088) );
  INV_X4 U5042 ( .I(n5541), .ZN(n12533) );
  INV_X4 U19815 ( .I(n20931), .ZN(n29990) );
  NOR2_X2 U2248 ( .A1(n23480), .A2(n9078), .ZN(n35013) );
  NAND2_X2 U18419 ( .A1(n3633), .A2(n11923), .ZN(n36594) );
  NAND2_X2 U28460 ( .A1(n20638), .A2(n20408), .ZN(n5464) );
  AOI21_X2 U7517 ( .A1(n28608), .A2(n11390), .B(n34737), .ZN(n6095) );
  OAI21_X2 U7151 ( .A1(n19944), .A2(n23171), .B(n23172), .ZN(n18331) );
  INV_X2 U2609 ( .I(n17923), .ZN(n16288) );
  INV_X2 U16342 ( .I(n26112), .ZN(n33753) );
  OAI21_X2 U2676 ( .A1(n17433), .A2(n33226), .B(n38878), .ZN(n17435) );
  NOR2_X2 U2789 ( .A1(n10931), .A2(n37355), .ZN(n32641) );
  INV_X2 U3467 ( .I(n14704), .ZN(n11265) );
  INV_X4 U833 ( .I(n12327), .ZN(n11910) );
  INV_X4 U1023 ( .I(n19886), .ZN(n1027) );
  NOR3_X2 U15338 ( .A1(n365), .A2(n33871), .A3(n13971), .ZN(n25759) );
  BUF_X2 U3448 ( .I(n7696), .Z(n19549) );
  INV_X2 U832 ( .I(n7676), .ZN(n35184) );
  NAND3_X1 U25604 ( .A1(n36217), .A2(n4976), .A3(n36216), .ZN(n11252) );
  INV_X4 U1655 ( .I(n4914), .ZN(n35449) );
  OAI21_X2 U1162 ( .A1(n33464), .A2(n33465), .B(n25345), .ZN(n26067) );
  INV_X2 U5159 ( .I(n5044), .ZN(n23572) );
  NAND2_X2 U18267 ( .A1(n4013), .A2(n18988), .ZN(n31114) );
  INV_X2 U894 ( .I(n5271), .ZN(n25154) );
  NAND2_X2 U18275 ( .A1(n18348), .A2(n37259), .ZN(n18347) );
  NAND2_X2 U5713 ( .A1(n37732), .A2(n20339), .ZN(n16881) );
  NAND2_X2 U3037 ( .A1(n9310), .A2(n32870), .ZN(n27270) );
  INV_X2 U18602 ( .I(n26063), .ZN(n25742) );
  OAI21_X2 U1135 ( .A1(n14793), .A2(n1106), .B(n3356), .ZN(n36574) );
  INV_X2 U3732 ( .I(n25943), .ZN(n6302) );
  OAI21_X2 U17046 ( .A1(n10055), .A2(n12629), .B(n34010), .ZN(n12601) );
  NAND2_X2 U3020 ( .A1(n30210), .A2(n30213), .ZN(n30212) );
  INV_X2 U351 ( .I(n37079), .ZN(n17032) );
  AND2_X1 U4773 ( .A1(n11044), .A2(n22222), .Z(n14474) );
  NAND2_X2 U1512 ( .A1(n18028), .A2(n20476), .ZN(n18954) );
  INV_X4 U8844 ( .I(n33514), .ZN(n13971) );
  NAND2_X2 U17449 ( .A1(n9265), .A2(n35290), .ZN(n164) );
  BUF_X2 U5070 ( .I(n23083), .Z(n19865) );
  OAI21_X2 U1855 ( .A1(n10840), .A2(n1301), .B(n32401), .ZN(n10842) );
  NAND2_X2 U467 ( .A1(n1074), .A2(n28180), .ZN(n27946) );
  OAI21_X2 U235 ( .A1(n35369), .A2(n35370), .B(n31269), .ZN(n34395) );
  INV_X2 U379 ( .I(n10883), .ZN(n33424) );
  NOR2_X2 U2931 ( .A1(n19728), .A2(n8527), .ZN(n8587) );
  NAND2_X2 U5903 ( .A1(n24558), .A2(n24757), .ZN(n31257) );
  INV_X4 U12427 ( .I(n25468), .ZN(n25409) );
  NAND3_X2 U10149 ( .A1(n12091), .A2(n937), .A3(n22252), .ZN(n22000) );
  INV_X2 U1713 ( .I(n24938), .ZN(n25031) );
  NAND2_X2 U9464 ( .A1(n14025), .A2(n1115), .ZN(n11954) );
  INV_X4 U2764 ( .I(n33933), .ZN(n20872) );
  AOI22_X2 U5800 ( .A1(n35157), .A2(n35156), .B1(n25592), .B2(n32105), .ZN(
        n19401) );
  OAI21_X2 U15187 ( .A1(n33094), .A2(n37936), .B(n33093), .ZN(n28960) );
  INV_X2 U245 ( .I(n28673), .ZN(n1068) );
  NOR2_X2 U5648 ( .A1(n26972), .A2(n5935), .ZN(n16000) );
  NOR2_X2 U2928 ( .A1(n30197), .A2(n30198), .ZN(n30199) );
  NOR2_X2 U858 ( .A1(n20052), .A2(n31809), .ZN(n8980) );
  NOR2_X2 U6404 ( .A1(n21879), .A2(n21878), .ZN(n22041) );
  NOR2_X2 U4271 ( .A1(n23550), .A2(n38614), .ZN(n23347) );
  AND2_X2 U143 ( .A1(n10422), .A2(n36426), .Z(n17444) );
  NAND2_X2 U22681 ( .A1(n4699), .A2(n3669), .ZN(n10321) );
  OAI22_X2 U12074 ( .A1(n25903), .A2(n33474), .B1(n26016), .B2(n38825), .ZN(
        n12458) );
  INV_X4 U7041 ( .I(n20517), .ZN(n1032) );
  NOR2_X2 U2355 ( .A1(n6005), .A2(n36230), .ZN(n32943) );
  NAND2_X2 U2214 ( .A1(n17816), .A2(n39371), .ZN(n32207) );
  NAND2_X1 U30050 ( .A1(n8580), .A2(n8579), .ZN(n7971) );
  INV_X2 U217 ( .I(n28791), .ZN(n248) );
  NAND2_X2 U7056 ( .A1(n25820), .A2(n36798), .ZN(n25931) );
  INV_X2 U14845 ( .I(n37954), .ZN(n24228) );
  NAND2_X2 U2500 ( .A1(n5876), .A2(n22236), .ZN(n35802) );
  NOR2_X2 U3497 ( .A1(n13038), .A2(n23349), .ZN(n16443) );
  NOR2_X2 U276 ( .A1(n14232), .A2(n28012), .ZN(n11876) );
  INV_X2 U3373 ( .I(n18545), .ZN(n1546) );
  INV_X1 U5707 ( .I(n37355), .ZN(n1578) );
  INV_X4 U6876 ( .I(n26086), .ZN(n25874) );
  INV_X2 U7479 ( .I(n1448), .ZN(n986) );
  INV_X2 U1970 ( .I(n9583), .ZN(n9579) );
  INV_X4 U11548 ( .I(n9893), .ZN(n955) );
  NAND2_X2 U8376 ( .A1(n23537), .A2(n23539), .ZN(n23225) );
  INV_X2 U7258 ( .I(n8413), .ZN(n8103) );
  INV_X2 U3909 ( .I(n38194), .ZN(n14064) );
  INV_X2 U12366 ( .I(n13988), .ZN(n9541) );
  AOI22_X2 U18050 ( .A1(n36092), .A2(n34128), .B1(n22060), .B2(n8618), .ZN(
        n22784) );
  NOR2_X2 U3868 ( .A1(n7387), .A2(n38724), .ZN(n36137) );
  OAI21_X2 U9750 ( .A1(n18141), .A2(n13710), .B(n1601), .ZN(n13709) );
  AND2_X2 U13820 ( .A1(n15697), .A2(n4342), .Z(n8618) );
  INV_X2 U7045 ( .I(n24095), .ZN(n24477) );
  INV_X2 U2142 ( .I(n23697), .ZN(n23779) );
  INV_X2 U26305 ( .I(n17605), .ZN(n22762) );
  NOR2_X2 U666 ( .A1(n16904), .A2(n16903), .ZN(n21265) );
  OAI21_X2 U27173 ( .A1(n28226), .A2(n35659), .B(n19921), .ZN(n20226) );
  AOI21_X2 U2178 ( .A1(n13691), .A2(n23645), .B(n35312), .ZN(n35285) );
  INV_X4 U20709 ( .I(n39678), .ZN(n8014) );
  NAND2_X2 U9861 ( .A1(n23462), .A2(n18090), .ZN(n18155) );
  NOR2_X1 U21571 ( .A1(n1275), .A2(n1131), .ZN(n9459) );
  OAI21_X2 U7796 ( .A1(n3515), .A2(n3514), .B(n27072), .ZN(n4492) );
  NAND2_X2 U6867 ( .A1(n7198), .A2(n24795), .ZN(n9614) );
  AOI22_X2 U465 ( .A1(n8880), .A2(n28194), .B1(n9897), .B2(n37251), .ZN(n3846)
         );
  NOR2_X2 U6314 ( .A1(n14392), .A2(n24300), .ZN(n13112) );
  AOI21_X2 U21139 ( .A1(n23452), .A2(n10480), .B(n8668), .ZN(n16713) );
  NOR2_X2 U14727 ( .A1(n34399), .A2(n11003), .ZN(n31299) );
  NAND2_X2 U4925 ( .A1(n8971), .A2(n21804), .ZN(n4298) );
  NAND2_X2 U12575 ( .A1(n24736), .A2(n37687), .ZN(n2850) );
  NAND3_X2 U2684 ( .A1(n19123), .A2(n19124), .A3(n19125), .ZN(n36072) );
  NAND2_X2 U16810 ( .A1(n32974), .A2(n25874), .ZN(n26088) );
  INV_X2 U2570 ( .I(n31573), .ZN(n36960) );
  INV_X2 U5030 ( .I(n35244), .ZN(n1288) );
  NAND2_X2 U6950 ( .A1(n14999), .A2(n13966), .ZN(n24757) );
  AOI21_X2 U3557 ( .A1(n25840), .A2(n11807), .B(n8233), .ZN(n8234) );
  AOI22_X2 U450 ( .A1(n37136), .A2(n28283), .B1(n13993), .B2(n16544), .ZN(
        n28170) );
  NAND2_X1 U14100 ( .A1(n34805), .A2(n29587), .ZN(n34804) );
  INV_X2 U27288 ( .I(n22349), .ZN(n1332) );
  BUF_X4 U30631 ( .I(n21912), .Z(n36912) );
  OAI22_X2 U3571 ( .A1(n14495), .A2(n15651), .B1(n16171), .B2(n30238), .ZN(
        n5632) );
  BUF_X2 U2491 ( .I(n32932), .Z(n31607) );
  OAI21_X1 U16049 ( .A1(n980), .A2(n28690), .B(n2639), .ZN(n31461) );
  INV_X2 U6695 ( .I(n9845), .ZN(n14451) );
  NOR2_X2 U13752 ( .A1(n14251), .A2(n22259), .ZN(n17001) );
  INV_X4 U8351 ( .I(n15461), .ZN(n1128) );
  INV_X4 U4436 ( .I(n31679), .ZN(n1265) );
  NAND3_X2 U13118 ( .A1(n17959), .A2(n17958), .A3(n38055), .ZN(n16031) );
  NOR2_X2 U9114 ( .A1(n18277), .A2(n18276), .ZN(n7034) );
  AND2_X1 U17676 ( .A1(n31917), .A2(n26090), .Z(n5682) );
  INV_X2 U8835 ( .I(n3257), .ZN(n27624) );
  INV_X2 U1392 ( .I(n260), .ZN(n16073) );
  BUF_X2 U10933 ( .I(n29296), .Z(n4816) );
  OR2_X1 U4450 ( .A1(n36827), .A2(n7023), .Z(n28606) );
  NOR2_X2 U571 ( .A1(n12260), .A2(n876), .ZN(n13984) );
  NAND2_X1 U4244 ( .A1(n5034), .A2(n9503), .ZN(n31640) );
  NAND3_X2 U1790 ( .A1(n13896), .A2(n30412), .A3(n27259), .ZN(n5374) );
  NOR2_X2 U7096 ( .A1(n603), .A2(n25797), .ZN(n25855) );
  NAND3_X2 U18732 ( .A1(n30470), .A2(n25519), .A3(n20924), .ZN(n5902) );
  OAI22_X2 U454 ( .A1(n33481), .A2(n28152), .B1(n16412), .B2(n8960), .ZN(
        n28402) );
  NAND2_X2 U1649 ( .A1(n31509), .A2(n5541), .ZN(n25416) );
  INV_X4 U16912 ( .I(n9733), .ZN(n32671) );
  INV_X4 U22334 ( .I(n28771), .ZN(n35777) );
  INV_X4 U190 ( .I(n28768), .ZN(n28771) );
  NAND2_X2 U213 ( .A1(n11488), .A2(n11490), .ZN(n28529) );
  NAND2_X2 U668 ( .A1(n10946), .A2(n36865), .ZN(n1835) );
  INV_X4 U994 ( .I(n17993), .ZN(n32745) );
  OAI21_X2 U60 ( .A1(n16988), .A2(n6863), .B(n39392), .ZN(n29273) );
  INV_X2 U6141 ( .I(n27777), .ZN(n1460) );
  NAND2_X2 U1085 ( .A1(n14378), .A2(n17709), .ZN(n14123) );
  NAND2_X2 U15923 ( .A1(n30290), .A2(n27282), .ZN(n26264) );
  INV_X2 U39 ( .I(n29568), .ZN(n29567) );
  INV_X2 U6211 ( .I(n23214), .ZN(n17568) );
  NAND2_X2 U6165 ( .A1(n36035), .A2(n35536), .ZN(n31475) );
  OR2_X1 U4426 ( .A1(n19658), .A2(n33937), .Z(n24225) );
  NOR2_X2 U25352 ( .A1(n20585), .A2(n21328), .ZN(n22306) );
  INV_X2 U936 ( .I(n26743), .ZN(n35877) );
  INV_X2 U7482 ( .I(n31279), .ZN(n1406) );
  INV_X2 U6045 ( .I(n21577), .ZN(n21593) );
  INV_X2 U1695 ( .I(n37050), .ZN(n17246) );
  NAND2_X2 U7050 ( .A1(n39301), .A2(n8212), .ZN(n8211) );
  NAND2_X2 U8924 ( .A1(n25604), .A2(n9029), .ZN(n34261) );
  INV_X2 U7617 ( .I(n29517), .ZN(n33427) );
  OAI21_X2 U929 ( .A1(n19886), .A2(n36296), .B(n12159), .ZN(n11198) );
  BUF_X2 U4755 ( .I(n12396), .Z(n33538) );
  BUF_X2 U10452 ( .I(Key[6]), .Z(n29649) );
  INV_X4 U7502 ( .I(n28396), .ZN(n32791) );
  INV_X2 U4845 ( .I(n1154), .ZN(n31649) );
  NOR2_X2 U9957 ( .A1(n10297), .A2(n10296), .ZN(n10295) );
  OAI21_X2 U8476 ( .A1(n8707), .A2(n1313), .B(n23142), .ZN(n10297) );
  INV_X1 U25462 ( .I(n36196), .ZN(n6898) );
  OAI22_X2 U30103 ( .A1(n25991), .A2(n11807), .B1(n18289), .B2(n9883), .ZN(
        n4854) );
  INV_X2 U1949 ( .I(n23619), .ZN(n20835) );
  NAND2_X2 U2353 ( .A1(n34185), .A2(n34184), .ZN(n22907) );
  NOR2_X2 U12977 ( .A1(n32683), .A2(n37107), .ZN(n4244) );
  NAND2_X2 U3798 ( .A1(n22055), .A2(n22132), .ZN(n22056) );
  AND2_X1 U4186 ( .A1(n25782), .A2(n8407), .Z(n13119) );
  AOI21_X2 U826 ( .A1(n25562), .A2(n25637), .B(n25436), .ZN(n25439) );
  NOR2_X2 U9703 ( .A1(n9634), .A2(n13809), .ZN(n21211) );
  BUF_X2 U17990 ( .I(n27211), .Z(n36203) );
  INV_X2 U30119 ( .I(n28109), .ZN(n33612) );
  NAND2_X2 U4628 ( .A1(n3013), .A2(n38168), .ZN(n9962) );
  INV_X4 U9353 ( .I(n19332), .ZN(n1235) );
  INV_X4 U11454 ( .I(n27478), .ZN(n27815) );
  NAND2_X2 U13732 ( .A1(n22107), .A2(n7613), .ZN(n17898) );
  INV_X2 U13611 ( .I(n22573), .ZN(n13768) );
  BUF_X4 U14090 ( .I(n3713), .Z(n32260) );
  NAND2_X2 U11321 ( .A1(n15389), .A2(n42), .ZN(n27936) );
  INV_X2 U5951 ( .I(n24794), .ZN(n1563) );
  NOR2_X2 U166 ( .A1(n1175), .A2(n35210), .ZN(n34619) );
  INV_X2 U6772 ( .I(n5323), .ZN(n23831) );
  OAI21_X2 U14696 ( .A1(n20395), .A2(n12286), .B(n24156), .ZN(n34895) );
  INV_X2 U13555 ( .I(n23189), .ZN(n1647) );
  NAND2_X2 U23637 ( .A1(n935), .A2(n35684), .ZN(n8869) );
  OAI21_X2 U808 ( .A1(n36262), .A2(n33026), .B(n33025), .ZN(n26153) );
  INV_X2 U438 ( .I(n27506), .ZN(n601) );
  OAI21_X2 U17190 ( .A1(n35897), .A2(n21248), .B(n30544), .ZN(n27506) );
  INV_X2 U4167 ( .I(n24308), .ZN(n24446) );
  INV_X2 U7300 ( .I(n1217), .ZN(n34943) );
  NOR2_X2 U23074 ( .A1(n1094), .A2(n1786), .ZN(n26957) );
  OAI21_X2 U3411 ( .A1(n13053), .A2(n27955), .B(n17477), .ZN(n385) );
  NOR2_X2 U1698 ( .A1(n25725), .A2(n38661), .ZN(n36686) );
  OAI21_X2 U5411 ( .A1(n14712), .A2(n14713), .B(n28627), .ZN(n36255) );
  NOR2_X2 U8929 ( .A1(n13714), .A2(n20896), .ZN(n27955) );
  AOI22_X2 U9604 ( .A1(n34666), .A2(n1121), .B1(n24782), .B2(n24658), .ZN(
        n4694) );
  NAND2_X2 U9478 ( .A1(n4217), .A2(n4216), .ZN(n4215) );
  AOI21_X2 U1164 ( .A1(n10290), .A2(n35109), .B(n20769), .ZN(n20768) );
  NAND2_X2 U2385 ( .A1(n18365), .A2(n17578), .ZN(n7012) );
  OAI21_X2 U695 ( .A1(n37191), .A2(n3998), .B(n3996), .ZN(n35037) );
  INV_X4 U7833 ( .I(n35919), .ZN(n1081) );
  INV_X4 U604 ( .I(n26695), .ZN(n1495) );
  NAND2_X2 U4602 ( .A1(n24693), .A2(n24721), .ZN(n30862) );
  INV_X4 U18359 ( .I(n30161), .ZN(n33277) );
  INV_X4 U5689 ( .I(n25434), .ZN(n25674) );
  INV_X2 U3970 ( .I(n6686), .ZN(n27416) );
  OAI21_X2 U960 ( .A1(n14921), .A2(n14922), .B(n1490), .ZN(n12684) );
  BUF_X2 U7912 ( .I(n20394), .Z(n17076) );
  NAND2_X2 U24130 ( .A1(n25622), .A2(n33785), .ZN(n2417) );
  INV_X2 U16 ( .I(n19297), .ZN(n29658) );
  NOR2_X2 U1205 ( .A1(n39061), .A2(n39160), .ZN(n4455) );
  OAI22_X2 U4058 ( .A1(n11009), .A2(n31321), .B1(n28716), .B2(n33591), .ZN(
        n16503) );
  AOI21_X1 U25465 ( .A1(n26606), .A2(n13219), .B(n26986), .ZN(n36196) );
  INV_X2 U24725 ( .I(n15004), .ZN(n16935) );
  INV_X2 U5876 ( .I(n4192), .ZN(n991) );
  OAI21_X2 U12916 ( .A1(n24142), .A2(n18302), .B(n14123), .ZN(n14780) );
  OAI21_X1 U1567 ( .A1(n18218), .A2(n34156), .B(n18217), .ZN(n25655) );
  NAND2_X2 U22515 ( .A1(n32526), .A2(n15324), .ZN(n16055) );
  NAND2_X2 U3436 ( .A1(n1783), .A2(n24700), .ZN(n1782) );
  NOR2_X2 U12045 ( .A1(n25781), .A2(n25774), .ZN(n15870) );
  INV_X4 U2323 ( .I(n21068), .ZN(n23518) );
  NAND3_X2 U1231 ( .A1(n25409), .A2(n14635), .A3(n25467), .ZN(n25339) );
  AOI21_X2 U14496 ( .A1(n24426), .A2(n3142), .B(n8041), .ZN(n2089) );
  NAND2_X2 U4515 ( .A1(n33392), .A2(n19507), .ZN(n12517) );
  NAND2_X2 U13240 ( .A1(n23362), .A2(n23480), .ZN(n15681) );
  AOI22_X2 U1905 ( .A1(n8916), .A2(n20863), .B1(n20864), .B2(n38302), .ZN(
        n11577) );
  BUF_X4 U16866 ( .I(n24745), .Z(n35137) );
  INV_X2 U10799 ( .I(n17978), .ZN(n30858) );
  INV_X2 U5928 ( .I(n17458), .ZN(n1243) );
  INV_X2 U7235 ( .I(n11327), .ZN(n22360) );
  INV_X2 U7082 ( .I(n17269), .ZN(n9227) );
  NAND2_X2 U2078 ( .A1(n253), .A2(n24443), .ZN(n24310) );
  AOI22_X2 U18655 ( .A1(n22072), .A2(n3687), .B1(n22071), .B2(n33623), .ZN(
        n22380) );
  AOI22_X2 U13831 ( .A1(n17264), .A2(n18417), .B1(n14542), .B2(n21712), .ZN(
        n12024) );
  INV_X4 U17461 ( .I(n19410), .ZN(n20157) );
  INV_X2 U6740 ( .I(n6176), .ZN(n20972) );
  NOR2_X2 U968 ( .A1(n36262), .A2(n36261), .ZN(n7859) );
  INV_X2 U1858 ( .I(n24707), .ZN(n24700) );
  AOI22_X2 U12911 ( .A1(n1274), .A2(n232), .B1(n1123), .B2(n24116), .ZN(n11133) );
  NOR2_X2 U5343 ( .A1(n1602), .A2(n23819), .ZN(n8690) );
  INV_X2 U1585 ( .I(n12836), .ZN(n26876) );
  NAND2_X2 U8683 ( .A1(n21727), .A2(n18293), .ZN(n11172) );
  INV_X4 U20951 ( .I(n1029), .ZN(n35578) );
  AOI21_X2 U9958 ( .A1(n11301), .A2(n33361), .B(n11299), .ZN(n18034) );
  NOR2_X2 U10200 ( .A1(n1675), .A2(n18656), .ZN(n17156) );
  OAI21_X1 U13890 ( .A1(n21715), .A2(n21714), .B(n21713), .ZN(n21716) );
  NAND2_X2 U813 ( .A1(n26148), .A2(n36262), .ZN(n33025) );
  NAND2_X2 U706 ( .A1(n5297), .A2(n1217), .ZN(n35144) );
  BUF_X2 U4544 ( .I(n10665), .Z(n33785) );
  NOR2_X2 U678 ( .A1(n15245), .A2(n35604), .ZN(n35603) );
  NOR2_X2 U22843 ( .A1(n17691), .A2(n17692), .ZN(n11159) );
  NOR2_X2 U30570 ( .A1(n12814), .A2(n22270), .ZN(n5147) );
  BUF_X4 U17894 ( .I(n26893), .Z(n33396) );
  NAND3_X2 U8952 ( .A1(n35392), .A2(n29520), .A3(n29521), .ZN(n29523) );
  NAND2_X2 U2374 ( .A1(n8707), .A2(n35591), .ZN(n8706) );
  AOI21_X2 U16487 ( .A1(n14229), .A2(n13712), .B(n1019), .ZN(n14224) );
  NAND2_X2 U9520 ( .A1(n25665), .A2(n4001), .ZN(n20442) );
  NAND2_X2 U118 ( .A1(n19896), .A2(n17295), .ZN(n17294) );
  INV_X2 U1631 ( .I(n20153), .ZN(n25327) );
  AOI21_X2 U19123 ( .A1(n6375), .A2(n6374), .B(n28287), .ZN(n6587) );
  INV_X2 U6749 ( .I(n20418), .ZN(n12638) );
  OAI21_X2 U502 ( .A1(n20941), .A2(n18013), .B(n14152), .ZN(n34965) );
  NOR2_X2 U1880 ( .A1(n2553), .A2(n23456), .ZN(n18763) );
  INV_X4 U26905 ( .I(n14501), .ZN(n21656) );
  AOI21_X2 U4572 ( .A1(n35023), .A2(n37081), .B(n38529), .ZN(n16255) );
  INV_X4 U946 ( .I(n5935), .ZN(n3694) );
  INV_X2 U8047 ( .I(n29794), .ZN(n16682) );
  NAND2_X2 U911 ( .A1(n26840), .A2(n32345), .ZN(n18095) );
  BUF_X4 U11048 ( .I(n19771), .Z(n7486) );
  NAND3_X2 U19876 ( .A1(n14437), .A2(n16060), .A3(n36850), .ZN(n31980) );
  NAND2_X1 U2923 ( .A1(n35787), .A2(n14664), .ZN(n16075) );
  INV_X2 U9029 ( .I(n8944), .ZN(n1433) );
  NAND2_X2 U6630 ( .A1(n20372), .A2(n34419), .ZN(n22843) );
  INV_X2 U6459 ( .I(n21982), .ZN(n1686) );
  AOI21_X2 U1154 ( .A1(n26107), .A2(n25825), .B(n16200), .ZN(n15551) );
  NOR2_X2 U5905 ( .A1(n18541), .A2(n16908), .ZN(n24716) );
  INV_X2 U30576 ( .I(n39067), .ZN(n24464) );
  INV_X2 U8360 ( .I(n23590), .ZN(n23874) );
  INV_X4 U3855 ( .I(n23053), .ZN(n1043) );
  NAND2_X2 U8427 ( .A1(n31644), .A2(n32260), .ZN(n3714) );
  BUF_X2 U7546 ( .I(n29042), .Z(n31782) );
  INV_X2 U17525 ( .I(n16539), .ZN(n31891) );
  NOR2_X1 U15894 ( .A1(n936), .A2(n14089), .ZN(n2272) );
  OAI21_X2 U947 ( .A1(n2929), .A2(n20578), .B(n38238), .ZN(n17416) );
  OR2_X1 U4700 ( .A1(n17594), .A2(n37085), .Z(n25615) );
  NAND2_X2 U2621 ( .A1(n5075), .A2(n9252), .ZN(n29) );
  INV_X4 U2129 ( .I(n23819), .ZN(n1123) );
  NAND2_X2 U28774 ( .A1(n33648), .A2(n18031), .ZN(n36612) );
  INV_X2 U6157 ( .I(n21808), .ZN(n1345) );
  NOR2_X2 U6869 ( .A1(n19484), .A2(n38884), .ZN(n24518) );
  NAND2_X2 U24437 ( .A1(n16729), .A2(n7379), .ZN(n16728) );
  AOI22_X2 U6213 ( .A1(n37073), .A2(n11858), .B1(n25888), .B2(n928), .ZN(
        n12941) );
  NAND2_X2 U2284 ( .A1(n36263), .A2(n17887), .ZN(n36131) );
  AOI21_X2 U7531 ( .A1(n33229), .A2(n28478), .B(n2191), .ZN(n16036) );
  AOI21_X2 U2859 ( .A1(n18999), .A2(n5821), .B(n31649), .ZN(n31953) );
  NAND2_X1 U17703 ( .A1(n21220), .A2(n20885), .ZN(n4901) );
  NAND2_X2 U1356 ( .A1(n34898), .A2(n26075), .ZN(n26079) );
  INV_X2 U1707 ( .I(n25392), .ZN(n25587) );
  INV_X4 U8256 ( .I(n32091), .ZN(n19484) );
  INV_X4 U4265 ( .I(n17118), .ZN(n22236) );
  NAND2_X2 U5715 ( .A1(n20545), .A2(n38899), .ZN(n36458) );
  AOI22_X2 U2447 ( .A1(n20590), .A2(n20344), .B1(n22793), .B2(n20174), .ZN(
        n34664) );
  NOR2_X2 U8480 ( .A1(n23121), .A2(n19440), .ZN(n30663) );
  INV_X2 U1407 ( .I(n31809), .ZN(n1537) );
  INV_X2 U12649 ( .I(n24770), .ZN(n12460) );
  INV_X2 U6643 ( .I(n20638), .ZN(n14524) );
  INV_X4 U413 ( .I(n36320), .ZN(n2191) );
  AOI21_X2 U2366 ( .A1(n36234), .A2(n27149), .B(n27235), .ZN(n5997) );
  INV_X2 U8553 ( .I(n17021), .ZN(n22921) );
  NAND2_X2 U11612 ( .A1(n5082), .A2(n37076), .ZN(n5297) );
  NAND2_X2 U704 ( .A1(n31150), .A2(n31298), .ZN(n34579) );
  AOI21_X2 U288 ( .A1(n33436), .A2(n1194), .B(n1431), .ZN(n19688) );
  INV_X4 U1361 ( .I(n35059), .ZN(n20813) );
  NAND2_X1 U9851 ( .A1(n9862), .A2(n23555), .ZN(n15325) );
  NAND2_X2 U2736 ( .A1(n27149), .A2(n27436), .ZN(n15983) );
  OAI21_X2 U14432 ( .A1(n11042), .A2(n11041), .B(n2035), .ZN(n11040) );
  INV_X2 U338 ( .I(n28570), .ZN(n37018) );
  OAI21_X2 U19003 ( .A1(n18617), .A2(n34121), .B(n34245), .ZN(n6463) );
  NOR2_X2 U20220 ( .A1(n11547), .A2(n1532), .ZN(n7513) );
  INV_X2 U2058 ( .I(n30000), .ZN(n21167) );
  OAI22_X2 U10718 ( .A1(n6862), .A2(n11056), .B1(n29421), .B2(n13153), .ZN(
        n6866) );
  NOR2_X2 U2493 ( .A1(n36085), .A2(n36084), .ZN(n4111) );
  NAND2_X2 U262 ( .A1(n12543), .A2(n28651), .ZN(n36144) );
  NOR2_X2 U3128 ( .A1(n19865), .A2(n20372), .ZN(n10470) );
  AOI21_X2 U845 ( .A1(n39117), .A2(n14079), .B(n1008), .ZN(n12405) );
  OAI21_X2 U23083 ( .A1(n365), .A2(n34154), .B(n2942), .ZN(n2941) );
  NOR2_X2 U12117 ( .A1(n39824), .A2(n11616), .ZN(n31018) );
  INV_X2 U399 ( .I(n32002), .ZN(n36775) );
  INV_X2 U6627 ( .I(n13686), .ZN(n925) );
  INV_X2 U22234 ( .I(n21721), .ZN(n21645) );
  AOI21_X2 U24714 ( .A1(n21573), .A2(n15839), .B(n20580), .ZN(n20579) );
  NOR2_X2 U13703 ( .A1(n18129), .A2(n1148), .ZN(n7868) );
  OAI21_X2 U9921 ( .A1(n17556), .A2(n23569), .B(n23543), .ZN(n23546) );
  INV_X2 U17034 ( .I(n25602), .ZN(n35157) );
  NAND2_X2 U4232 ( .A1(n1029), .A2(n9825), .ZN(n24752) );
  OAI22_X2 U19849 ( .A1(n31975), .A2(n17266), .B1(n21745), .B2(n19542), .ZN(
        n19906) );
  NAND2_X2 U19188 ( .A1(n1148), .A2(n584), .ZN(n6450) );
  INV_X4 U11103 ( .I(n865), .ZN(n6615) );
  NAND2_X2 U6579 ( .A1(n22133), .A2(n22132), .ZN(n4121) );
  NAND2_X2 U154 ( .A1(n36924), .A2(n12353), .ZN(n36923) );
  INV_X2 U5748 ( .I(n14477), .ZN(n1136) );
  INV_X2 U1063 ( .I(n36858), .ZN(n865) );
  INV_X4 U6959 ( .I(n17658), .ZN(n1118) );
  NAND2_X1 U8298 ( .A1(n30651), .A2(n2889), .ZN(n4460) );
  INV_X4 U1156 ( .I(n18142), .ZN(n31133) );
  NAND2_X2 U2555 ( .A1(n33571), .A2(n35290), .ZN(n22141) );
  OAI21_X2 U14770 ( .A1(n4367), .A2(n30175), .B(n39122), .ZN(n34903) );
  NAND2_X2 U15651 ( .A1(n39501), .A2(n17658), .ZN(n24161) );
  OAI21_X2 U1479 ( .A1(n14666), .A2(n9602), .B(n1249), .ZN(n35492) );
  NAND2_X2 U30066 ( .A1(n1432), .A2(n4232), .ZN(n28605) );
  NAND2_X1 U20475 ( .A1(n16868), .A2(n12192), .ZN(n18019) );
  NOR3_X2 U28376 ( .A1(n39284), .A2(n32039), .A3(n196), .ZN(n21965) );
  OAI21_X2 U6028 ( .A1(n18752), .A2(n30378), .B(n16081), .ZN(n36725) );
  NOR2_X2 U10271 ( .A1(n34025), .A2(n34393), .ZN(n34392) );
  NOR2_X2 U11881 ( .A1(n26982), .A2(n26979), .ZN(n4982) );
  NOR3_X2 U2182 ( .A1(n32858), .A2(n1297), .A3(n6969), .ZN(n18680) );
  NAND3_X2 U1200 ( .A1(n17003), .A2(n26133), .A3(n25936), .ZN(n21306) );
  NAND2_X2 U11593 ( .A1(n37201), .A2(n27284), .ZN(n9493) );
  AND3_X1 U13792 ( .A1(n22315), .A2(n15004), .A3(n22277), .Z(n14508) );
  INV_X2 U24678 ( .I(n35832), .ZN(n20692) );
  NOR2_X1 U12796 ( .A1(n19453), .A2(n12040), .ZN(n33468) );
  NOR2_X2 U9714 ( .A1(n5714), .A2(n20653), .ZN(n5713) );
  OAI21_X2 U22491 ( .A1(n23060), .A2(n36724), .B(n19535), .ZN(n22705) );
  BUF_X4 U5216 ( .I(n23592), .Z(n4147) );
  INV_X2 U2161 ( .I(n23976), .ZN(n1616) );
  AOI21_X2 U9243 ( .A1(n26667), .A2(n17237), .B(n1002), .ZN(n14280) );
  AOI21_X2 U442 ( .A1(n6714), .A2(n879), .B(n38365), .ZN(n6713) );
  INV_X4 U17069 ( .I(n33453), .ZN(n6217) );
  NOR2_X2 U19489 ( .A1(n6770), .A2(n37210), .ZN(n14168) );
  OR2_X2 U6947 ( .A1(n1118), .A2(n24226), .Z(n24964) );
  INV_X2 U9365 ( .I(n26463), .ZN(n1238) );
  INV_X2 U747 ( .I(n27404), .ZN(n1079) );
  NAND2_X1 U24476 ( .A1(n2726), .A2(n17319), .ZN(n2725) );
  OAI21_X2 U1552 ( .A1(n13949), .A2(n13948), .B(n26986), .ZN(n13947) );
  INV_X4 U6723 ( .I(n34962), .ZN(n1642) );
  OAI21_X2 U6488 ( .A1(n22265), .A2(n19515), .B(n22267), .ZN(n33781) );
  BUF_X4 U1906 ( .I(n22234), .Z(n19261) );
  NOR2_X1 U6331 ( .A1(n23529), .A2(n18236), .ZN(n8928) );
  NOR2_X1 U13093 ( .A1(n36248), .A2(n36247), .ZN(n36246) );
  OAI21_X2 U2530 ( .A1(n1327), .A2(n11329), .B(n22287), .ZN(n34822) );
  INV_X1 U1539 ( .I(n21722), .ZN(n21640) );
  OAI21_X2 U15423 ( .A1(n10473), .A2(n32782), .B(n25748), .ZN(n26478) );
  OAI21_X2 U7851 ( .A1(n3417), .A2(n1500), .B(n33689), .ZN(n2238) );
  BUF_X4 U1781 ( .I(n7923), .Z(n2576) );
  INV_X1 U3927 ( .I(n25490), .ZN(n25517) );
  AOI22_X2 U13238 ( .A1(n23556), .A2(n31234), .B1(n16443), .B2(n32616), .ZN(
        n23558) );
  AOI21_X2 U8589 ( .A1(n916), .A2(n22349), .B(n2910), .ZN(n7814) );
  OAI21_X2 U11772 ( .A1(n10678), .A2(n10187), .B(n26354), .ZN(n10186) );
  OAI21_X2 U12438 ( .A1(n9526), .A2(n18837), .B(n38685), .ZN(n12599) );
  BUF_X4 U7247 ( .I(n22113), .Z(n1049) );
  NOR2_X1 U13230 ( .A1(n596), .A2(n3926), .ZN(n32721) );
  NAND2_X2 U2420 ( .A1(n10345), .A2(n21402), .ZN(n14846) );
  INV_X4 U8518 ( .I(n33745), .ZN(n11328) );
  AOI21_X2 U17009 ( .A1(n683), .A2(n123), .B(n35153), .ZN(n10128) );
  NAND2_X1 U17565 ( .A1(n9278), .A2(n17456), .ZN(n5015) );
  OR3_X1 U4658 ( .A1(n15414), .A2(n20128), .A3(n14064), .Z(n13664) );
  NAND2_X2 U7848 ( .A1(n13156), .A2(n14757), .ZN(n27390) );
  OAI21_X2 U532 ( .A1(n1494), .A2(n20211), .B(n13757), .ZN(n20636) );
  INV_X4 U14844 ( .I(n2395), .ZN(n12733) );
  OAI21_X2 U5615 ( .A1(n4776), .A2(n25897), .B(n37582), .ZN(n6397) );
  INV_X4 U4467 ( .I(n1302), .ZN(n17167) );
  INV_X4 U27294 ( .I(n18585), .ZN(n19262) );
  CLKBUF_X4 U5845 ( .I(n25157), .Z(n25754) );
  NOR2_X2 U7360 ( .A1(n13266), .A2(n1079), .ZN(n36080) );
  NOR2_X2 U17528 ( .A1(n12955), .A2(n10569), .ZN(n12954) );
  OAI21_X2 U8412 ( .A1(n23588), .A2(n19686), .B(n37757), .ZN(n8046) );
  NOR2_X2 U9898 ( .A1(n23620), .A2(n33080), .ZN(n9587) );
  BUF_X2 U6873 ( .I(n13779), .Z(n31385) );
  INV_X2 U24081 ( .I(n13635), .ZN(n17691) );
  NAND2_X2 U247 ( .A1(n35479), .A2(n35478), .ZN(n30786) );
  CLKBUF_X4 U2312 ( .I(n18525), .Z(n20525) );
  INV_X4 U25847 ( .I(n1257), .ZN(n25467) );
  NOR2_X2 U167 ( .A1(n14437), .A2(n29937), .ZN(n12275) );
  INV_X4 U2213 ( .I(n1109), .ZN(n25661) );
  INV_X2 U21661 ( .I(n9539), .ZN(n11598) );
  NAND2_X2 U17981 ( .A1(n24244), .A2(n11673), .ZN(n30526) );
  INV_X4 U14842 ( .I(n2393), .ZN(n24327) );
  NAND2_X2 U10361 ( .A1(n36728), .A2(n35116), .ZN(n21945) );
  NAND2_X2 U24378 ( .A1(n18524), .A2(n4664), .ZN(n17232) );
  OAI22_X2 U24896 ( .A1(n18734), .A2(n19637), .B1(n25386), .B2(n4048), .ZN(
        n18524) );
  NOR2_X2 U30001 ( .A1(n13491), .A2(n37671), .ZN(n3234) );
  BUF_X4 U10331 ( .I(n35828), .Z(n34399) );
  INV_X4 U22940 ( .I(n8042), .ZN(n33104) );
  OAI22_X2 U4657 ( .A1(n10160), .A2(n37525), .B1(n35901), .B2(n10161), .ZN(
        n10159) );
  OAI21_X2 U7969 ( .A1(n17179), .A2(n10807), .B(n17178), .ZN(n25441) );
  AOI21_X2 U5721 ( .A1(n26805), .A2(n26804), .B(n13713), .ZN(n20245) );
  BUF_X4 U5393 ( .I(n28550), .Z(n29596) );
  OAI21_X2 U10376 ( .A1(n21751), .A2(n17102), .B(n21889), .ZN(n5979) );
  OAI21_X2 U17679 ( .A1(n38100), .A2(n15555), .B(n7024), .ZN(n35191) );
  OAI21_X2 U1265 ( .A1(n20105), .A2(n31131), .B(n32722), .ZN(n31634) );
  INV_X2 U13030 ( .I(n39815), .ZN(n8581) );
  NOR2_X2 U16389 ( .A1(n28051), .A2(n19750), .ZN(n10516) );
  INV_X2 U24736 ( .I(n35116), .ZN(n20242) );
  INV_X4 U6633 ( .I(n28238), .ZN(n2740) );
  OAI21_X1 U21976 ( .A1(n15967), .A2(n13411), .B(n22258), .ZN(n22767) );
  NAND2_X2 U6032 ( .A1(n7608), .A2(n5305), .ZN(n22197) );
  NOR2_X2 U9334 ( .A1(n39117), .A2(n1008), .ZN(n12173) );
  NAND2_X2 U20405 ( .A1(n14085), .A2(n37075), .ZN(n14084) );
  INV_X2 U5172 ( .I(n15423), .ZN(n23380) );
  AOI21_X2 U7407 ( .A1(n32961), .A2(n27391), .B(n13699), .ZN(n14797) );
  NAND3_X2 U835 ( .A1(n33333), .A2(n4007), .A3(n26933), .ZN(n26644) );
  NOR2_X2 U13686 ( .A1(n5932), .A2(n34776), .ZN(n17221) );
  NAND2_X2 U11810 ( .A1(n20562), .A2(n26610), .ZN(n7855) );
  NAND2_X1 U16642 ( .A1(n17811), .A2(n35122), .ZN(n24380) );
  INV_X2 U12311 ( .I(n25470), .ZN(n2962) );
  NAND2_X2 U7028 ( .A1(n1257), .A2(n10004), .ZN(n25470) );
  BUF_X2 U13024 ( .I(n18269), .Z(n10008) );
  NOR2_X1 U24401 ( .A1(n15206), .A2(n15205), .ZN(n15223) );
  NOR2_X2 U3969 ( .A1(n32488), .A2(n36634), .ZN(n10374) );
  BUF_X4 U3952 ( .I(n16174), .Z(n2771) );
  NOR2_X2 U18553 ( .A1(n5707), .A2(n5706), .ZN(n28713) );
  INV_X1 U25670 ( .I(n17197), .ZN(n28192) );
  NOR2_X2 U18765 ( .A1(n32944), .A2(n12056), .ZN(n31810) );
  CLKBUF_X4 U3548 ( .I(n3903), .Z(n32012) );
  CLKBUF_X4 U3312 ( .I(n21567), .Z(n3293) );
  INV_X4 U30070 ( .I(n37107), .ZN(n33580) );
  NOR2_X2 U12637 ( .A1(n10606), .A2(n10605), .ZN(n31060) );
  INV_X2 U886 ( .I(n7377), .ZN(n24896) );
  NAND3_X2 U1270 ( .A1(n7026), .A2(n7025), .A3(n6366), .ZN(n6860) );
  AOI21_X2 U18192 ( .A1(n1404), .A2(n29486), .B(n31667), .ZN(n33425) );
  BUF_X2 U11967 ( .I(n26512), .Z(n26934) );
  INV_X2 U1349 ( .I(n16678), .ZN(n23011) );
  BUF_X2 U11965 ( .I(n26779), .Z(n5537) );
  OAI22_X2 U3713 ( .A1(n27300), .A2(n36989), .B1(n27171), .B2(n27170), .ZN(
        n27172) );
  INV_X4 U8197 ( .I(n9526), .ZN(n1115) );
  BUF_X2 U25231 ( .I(n17915), .Z(n32924) );
  INV_X2 U2388 ( .I(n18204), .ZN(n1630) );
  NAND2_X1 U7272 ( .A1(n9614), .A2(n36321), .ZN(n9612) );
  NOR2_X2 U12025 ( .A1(n4794), .A2(n6062), .ZN(n8135) );
  OR3_X1 U4681 ( .A1(n33333), .A2(n26932), .A3(n37235), .Z(n32072) );
  NAND2_X2 U2996 ( .A1(n6366), .A2(n8245), .ZN(n8594) );
  NAND2_X2 U161 ( .A1(n14178), .A2(n14179), .ZN(n8726) );
  INV_X4 U17632 ( .I(n19544), .ZN(n31603) );
  NAND2_X2 U976 ( .A1(n30348), .A2(n38238), .ZN(n17739) );
  NAND3_X2 U7986 ( .A1(n26076), .A2(n11807), .A3(n26077), .ZN(n7171) );
  BUF_X4 U3363 ( .I(n17810), .Z(n33101) );
  INV_X2 U21858 ( .I(n37498), .ZN(n25316) );
  AOI21_X2 U1140 ( .A1(n25996), .A2(n25995), .B(n37211), .ZN(n36949) );
  BUF_X2 U1225 ( .I(n2349), .Z(n586) );
  INV_X2 U618 ( .I(n37104), .ZN(n7195) );
  OAI21_X2 U919 ( .A1(n26805), .A2(n13713), .B(n1091), .ZN(n31447) );
  INV_X4 U15833 ( .I(n34813), .ZN(n916) );
  INV_X2 U5644 ( .I(n4458), .ZN(n13713) );
  NAND2_X2 U1614 ( .A1(n6696), .A2(n591), .ZN(n14443) );
  BUF_X4 U4909 ( .I(n13973), .Z(n1890) );
  INV_X2 U18222 ( .I(n10143), .ZN(n35313) );
  AOI21_X2 U2761 ( .A1(n15084), .A2(n33745), .B(n35564), .ZN(n15082) );
  NAND2_X2 U2448 ( .A1(n18244), .A2(n23101), .ZN(n35528) );
  NOR2_X2 U883 ( .A1(n4748), .A2(n18870), .ZN(n2339) );
  INV_X2 U2023 ( .I(n27385), .ZN(n19132) );
  NOR2_X2 U796 ( .A1(n31710), .A2(n31708), .ZN(n34776) );
  NOR2_X1 U12396 ( .A1(n7583), .A2(n35271), .ZN(n1873) );
  NOR2_X2 U7234 ( .A1(n26794), .A2(n925), .ZN(n12172) );
  BUF_X4 U6161 ( .I(n3092), .Z(n2035) );
  NOR2_X1 U3982 ( .A1(n20363), .A2(n20362), .ZN(n14351) );
  INV_X2 U6503 ( .I(n17127), .ZN(n18867) );
  NAND2_X2 U17097 ( .A1(n17693), .A2(n16271), .ZN(n17711) );
  INV_X4 U26779 ( .I(n36361), .ZN(n14501) );
  NAND2_X2 U1575 ( .A1(n24612), .A2(n6977), .ZN(n32367) );
  NOR2_X1 U1258 ( .A1(n32510), .A2(n26134), .ZN(n6749) );
  AOI21_X2 U5423 ( .A1(n30740), .A2(n28480), .B(n3532), .ZN(n34266) );
  BUF_X2 U4817 ( .I(n8365), .Z(n591) );
  OAI22_X2 U9387 ( .A1(n1242), .A2(n5883), .B1(n1523), .B2(n5882), .ZN(n5881)
         );
  NAND2_X2 U9279 ( .A1(n16267), .A2(n22352), .ZN(n3972) );
  OAI22_X2 U9999 ( .A1(n18072), .A2(n22799), .B1(n22800), .B2(n23209), .ZN(
        n22801) );
  INV_X2 U7267 ( .I(n21912), .ZN(n1155) );
  INV_X2 U18123 ( .I(n5131), .ZN(n19587) );
  AOI22_X2 U18540 ( .A1(n39365), .A2(n37880), .B1(n37981), .B2(n28302), .ZN(
        n28304) );
  INV_X1 U10893 ( .I(n29900), .ZN(n6204) );
  INV_X1 U6353 ( .I(n21687), .ZN(n6234) );
  INV_X2 U554 ( .I(n26802), .ZN(n26804) );
  NAND2_X1 U23858 ( .A1(n32743), .A2(n39595), .ZN(n33302) );
  NOR2_X2 U12245 ( .A1(n12096), .A2(n12097), .ZN(n31028) );
  NOR2_X2 U9095 ( .A1(n30952), .A2(n30951), .ZN(n18891) );
  INV_X2 U17524 ( .I(n31584), .ZN(n31585) );
  AOI21_X1 U11503 ( .A1(n36969), .A2(n27214), .B(n2922), .ZN(n8645) );
  NOR2_X2 U7446 ( .A1(n1200), .A2(n4457), .ZN(n32585) );
  NOR2_X1 U10975 ( .A1(n14787), .A2(n14773), .ZN(n31717) );
  NAND2_X2 U12131 ( .A1(n491), .A2(n18420), .ZN(n31795) );
  NAND2_X2 U6656 ( .A1(n8197), .A2(n1831), .ZN(n7025) );
  AOI21_X2 U10316 ( .A1(n21909), .A2(n21462), .B(n668), .ZN(n7526) );
  BUF_X2 U16553 ( .I(n38901), .Z(n15996) );
  INV_X2 U1100 ( .I(n8193), .ZN(n20537) );
  AOI21_X2 U8671 ( .A1(n6349), .A2(n6350), .B(n21561), .ZN(n6348) );
  OAI21_X1 U9244 ( .A1(n30942), .A2(n1493), .B(n4651), .ZN(n11306) );
  INV_X2 U724 ( .I(n13712), .ZN(n14228) );
  NOR2_X2 U27468 ( .A1(n35839), .A2(n19084), .ZN(n21943) );
  INV_X2 U18100 ( .I(n24419), .ZN(n16917) );
  INV_X2 U28291 ( .I(n21602), .ZN(n21662) );
  NAND2_X2 U4607 ( .A1(n5662), .A2(n38566), .ZN(n36615) );
  NOR2_X2 U26165 ( .A1(n21987), .A2(n22342), .ZN(n22345) );
  NOR2_X2 U3256 ( .A1(n24694), .A2(n24590), .ZN(n24576) );
  INV_X1 U17051 ( .I(n9828), .ZN(n35175) );
  NAND2_X2 U13887 ( .A1(n21580), .A2(n1847), .ZN(n10652) );
  AOI21_X2 U7129 ( .A1(n25979), .A2(n34265), .B(n37175), .ZN(n25984) );
  OR2_X1 U17137 ( .A1(n33561), .A2(n17022), .Z(n20666) );
  CLKBUF_X4 U20873 ( .I(n19713), .Z(n35560) );
  OR3_X2 U12626 ( .A1(n19586), .A2(n31093), .A3(n33745), .Z(n22820) );
  BUF_X4 U9570 ( .I(n13410), .Z(n9526) );
  NAND2_X1 U10499 ( .A1(n37228), .A2(n13817), .ZN(n20969) );
  INV_X4 U3291 ( .I(n5089), .ZN(n30851) );
  INV_X2 U27549 ( .I(n19298), .ZN(n26932) );
  INV_X4 U4697 ( .I(n22307), .ZN(n4200) );
  OAI22_X2 U13183 ( .A1(n20278), .A2(n37014), .B1(n20620), .B2(n22987), .ZN(
        n7041) );
  NOR2_X2 U4932 ( .A1(n19549), .A2(n16305), .ZN(n21336) );
  NAND2_X2 U797 ( .A1(n27347), .A2(n19477), .ZN(n8165) );
  INV_X1 U25461 ( .I(n25412), .ZN(n17020) );
  INV_X2 U27706 ( .I(n21869), .ZN(n21570) );
  NAND3_X2 U12063 ( .A1(n34116), .A2(n1781), .A3(n1777), .ZN(n22742) );
  INV_X2 U17311 ( .I(n197), .ZN(n35176) );
  INV_X2 U4992 ( .I(n4210), .ZN(n15513) );
  NAND2_X2 U12867 ( .A1(n18256), .A2(n15143), .ZN(n16744) );
  NAND2_X2 U24787 ( .A1(n19697), .A2(n12392), .ZN(n19530) );
  INV_X2 U6048 ( .I(n20778), .ZN(n14499) );
  OAI21_X2 U2173 ( .A1(n9669), .A2(n9670), .B(n20588), .ZN(n17819) );
  INV_X2 U1527 ( .I(n21484), .ZN(n9670) );
  INV_X2 U12501 ( .I(n20333), .ZN(n16673) );
  INV_X2 U4309 ( .I(n24817), .ZN(n24828) );
  NOR2_X2 U15603 ( .A1(n35019), .A2(n22030), .ZN(n35818) );
  NAND2_X2 U2948 ( .A1(n8734), .A2(n28725), .ZN(n8733) );
  OAI21_X2 U5573 ( .A1(n30696), .A2(n30695), .B(n26004), .ZN(n16118) );
  INV_X2 U1474 ( .I(n19543), .ZN(n6504) );
  AOI21_X2 U242 ( .A1(n37018), .A2(n28448), .B(n979), .ZN(n13806) );
  NAND2_X1 U5543 ( .A1(n33887), .A2(n34037), .ZN(n10949) );
  NOR2_X2 U18695 ( .A1(n15155), .A2(n32114), .ZN(n32113) );
  NAND3_X2 U829 ( .A1(n10567), .A2(n10098), .A3(n17047), .ZN(n18605) );
  NAND2_X2 U30485 ( .A1(n6615), .A2(n16834), .ZN(n10098) );
  OAI21_X2 U5298 ( .A1(n21661), .A2(n21946), .B(n32664), .ZN(n15805) );
  NAND2_X1 U22541 ( .A1(n28770), .A2(n28769), .ZN(n10596) );
  AOI22_X2 U7487 ( .A1(n32324), .A2(n2876), .B1(n32705), .B2(n39132), .ZN(
        n2873) );
  OR2_X1 U17811 ( .A1(n3827), .A2(n3826), .Z(n3825) );
  NAND2_X2 U426 ( .A1(n17735), .A2(n33765), .ZN(n14737) );
  CLKBUF_X4 U2642 ( .I(n7062), .Z(n35071) );
  INV_X2 U20317 ( .I(n26512), .ZN(n26937) );
  NAND2_X2 U825 ( .A1(n26774), .A2(n3919), .ZN(n3918) );
  INV_X1 U18052 ( .I(n11297), .ZN(n17535) );
  BUF_X4 U1014 ( .I(n26485), .Z(n33194) );
  NAND2_X2 U29427 ( .A1(n30629), .A2(n17458), .ZN(n25889) );
  INV_X1 U7957 ( .I(n25261), .ZN(n3568) );
  NAND2_X2 U2773 ( .A1(n28544), .A2(n13372), .ZN(n34870) );
  NOR2_X2 U24516 ( .A1(n15314), .A2(n32849), .ZN(n8595) );
  INV_X2 U7722 ( .I(n28205), .ZN(n1438) );
  NOR2_X2 U2189 ( .A1(n39666), .A2(n12144), .ZN(n33226) );
  INV_X2 U16786 ( .I(n6548), .ZN(n11375) );
  INV_X2 U6281 ( .I(n2186), .ZN(n35019) );
  INV_X4 U11781 ( .I(n27184), .ZN(n30986) );
  AOI21_X2 U9382 ( .A1(n26083), .A2(n4163), .B(n3277), .ZN(n9174) );
  INV_X2 U18471 ( .I(n37094), .ZN(n17117) );
  NAND3_X2 U811 ( .A1(n30851), .A2(n35904), .A3(n27081), .ZN(n30556) );
  CLKBUF_X4 U2287 ( .I(n23523), .Z(n30835) );
  OR2_X2 U23582 ( .A1(n10379), .A2(n37043), .Z(n10378) );
  CLKBUF_X4 U8168 ( .I(n38197), .Z(n10055) );
  BUF_X4 U13618 ( .I(n22573), .Z(n9874) );
  NOR2_X2 U9497 ( .A1(n13218), .A2(n19367), .ZN(n13197) );
  NAND2_X2 U23019 ( .A1(n11484), .A2(n12446), .ZN(n15287) );
  INV_X4 U3003 ( .I(n23108), .ZN(n1142) );
  INV_X2 U10229 ( .I(n20397), .ZN(n19778) );
  BUF_X4 U27068 ( .I(n23108), .Z(n33196) );
  NAND2_X2 U14277 ( .A1(n19028), .A2(n1597), .ZN(n13026) );
  INV_X2 U22577 ( .I(n10655), .ZN(n17237) );
  INV_X2 U23963 ( .I(n13417), .ZN(n20018) );
  INV_X4 U1592 ( .I(n24694), .ZN(n9656) );
  BUF_X2 U4652 ( .I(n30447), .Z(n545) );
  NAND3_X2 U1739 ( .A1(n7847), .A2(n18509), .A3(n37389), .ZN(n13629) );
  NOR2_X2 U22895 ( .A1(n37033), .A2(n37032), .ZN(n14813) );
  OAI21_X2 U3135 ( .A1(n12983), .A2(n3101), .B(n1116), .ZN(n17173) );
  NAND2_X2 U2767 ( .A1(n31283), .A2(n5570), .ZN(n29188) );
  BUF_X2 U11952 ( .I(n26919), .Z(n13392) );
  INV_X2 U1087 ( .I(n6130), .ZN(n26573) );
  INV_X2 U6374 ( .I(n2147), .ZN(n28750) );
  INV_X2 U6761 ( .I(n9518), .ZN(n9154) );
  NAND2_X2 U8315 ( .A1(n34216), .A2(n38687), .ZN(n22303) );
  OAI21_X2 U1688 ( .A1(n38702), .A2(n15049), .B(n17163), .ZN(n33187) );
  NAND2_X2 U2229 ( .A1(n23039), .A2(n17995), .ZN(n15799) );
  NAND2_X2 U924 ( .A1(n26810), .A2(n14377), .ZN(n26812) );
  NOR2_X2 U16861 ( .A1(n35135), .A2(n30384), .ZN(n33755) );
  NAND2_X2 U16864 ( .A1(n4321), .A2(n18744), .ZN(n35135) );
  NOR2_X2 U8716 ( .A1(n14499), .A2(n21521), .ZN(n21412) );
  NAND2_X2 U17723 ( .A1(n2878), .A2(n11283), .ZN(n2874) );
  NOR2_X2 U287 ( .A1(n17532), .A2(n32705), .ZN(n2878) );
  INV_X2 U13281 ( .I(n23039), .ZN(n11797) );
  INV_X2 U9 ( .I(n20437), .ZN(n29570) );
  INV_X2 U5489 ( .I(n25509), .ZN(n33834) );
  INV_X4 U27814 ( .I(n15102), .ZN(n16460) );
  INV_X1 U4483 ( .I(n20566), .ZN(n5384) );
  OAI21_X2 U19771 ( .A1(n27278), .A2(n9875), .B(n38305), .ZN(n7694) );
  INV_X2 U1531 ( .I(n21857), .ZN(n21860) );
  NAND2_X2 U12137 ( .A1(n1012), .A2(n6506), .ZN(n8236) );
  NAND2_X2 U23407 ( .A1(n18188), .A2(n19410), .ZN(n28119) );
  NAND2_X2 U11905 ( .A1(n5997), .A2(n5998), .ZN(n34836) );
  NAND3_X2 U9841 ( .A1(n18155), .A2(n23459), .A3(n35808), .ZN(n23241) );
  BUF_X4 U5687 ( .I(n25720), .Z(n18519) );
  AOI21_X1 U18131 ( .A1(n5145), .A2(n29813), .B(n5144), .ZN(n5143) );
  NOR2_X2 U15731 ( .A1(n33270), .A2(n831), .ZN(n4952) );
  OAI21_X2 U622 ( .A1(n31000), .A2(n11088), .B(n35114), .ZN(n11087) );
  AOI22_X2 U10036 ( .A1(n19054), .A2(n33969), .B1(n38752), .B2(n1653), .ZN(
        n18748) );
  OR2_X2 U1566 ( .A1(n15159), .A2(n30844), .Z(n12705) );
  NAND2_X1 U12252 ( .A1(n12780), .A2(n12779), .ZN(n12778) );
  INV_X4 U7202 ( .I(n10440), .ZN(n30795) );
  INV_X2 U18567 ( .I(n19473), .ZN(n24309) );
  NOR2_X2 U24402 ( .A1(n277), .A2(n24168), .ZN(n24182) );
  INV_X4 U14366 ( .I(n2416), .ZN(n25622) );
  INV_X1 U199 ( .I(n11348), .ZN(n35870) );
  OAI21_X2 U24756 ( .A1(n18408), .A2(n1676), .B(n17869), .ZN(n17557) );
  NOR2_X2 U2671 ( .A1(n10441), .A2(n10442), .ZN(n35038) );
  INV_X2 U22419 ( .I(n39096), .ZN(n22937) );
  OAI21_X2 U17684 ( .A1(n38100), .A2(n15555), .B(n7024), .ZN(n35192) );
  INV_X2 U3356 ( .I(n12856), .ZN(n17810) );
  OAI21_X2 U8687 ( .A1(n21551), .A2(n21763), .B(n33771), .ZN(n6670) );
  BUF_X4 U17635 ( .I(n21608), .Z(n12144) );
  AOI21_X2 U1925 ( .A1(n34046), .A2(n33513), .B(n35086), .ZN(n5330) );
  NAND2_X2 U12417 ( .A1(n19767), .A2(n32722), .ZN(n4454) );
  BUF_X4 U2823 ( .I(n33417), .Z(n32131) );
  INV_X2 U17634 ( .I(n21608), .ZN(n17233) );
  NOR2_X2 U4245 ( .A1(n12144), .A2(n21779), .ZN(n21535) );
  NOR2_X2 U11213 ( .A1(n17615), .A2(n32352), .ZN(n17085) );
  AOI21_X2 U9411 ( .A1(n12457), .A2(n25751), .B(n1522), .ZN(n12456) );
  NAND3_X2 U4919 ( .A1(n21788), .A2(n32456), .A3(n21787), .ZN(n16951) );
  NOR2_X2 U11913 ( .A1(n7978), .A2(n26703), .ZN(n13644) );
  INV_X2 U8907 ( .I(n29777), .ZN(n1402) );
  NAND2_X1 U13724 ( .A1(n1838), .A2(n554), .ZN(n1837) );
  BUF_X2 U10418 ( .I(n15354), .Z(n11274) );
  OAI21_X2 U2257 ( .A1(n21208), .A2(n37012), .B(n17167), .ZN(n12268) );
  AOI21_X2 U9858 ( .A1(n23462), .A2(n1140), .B(n5083), .ZN(n23299) );
  OR2_X2 U1377 ( .A1(n25351), .A2(n18121), .Z(n19264) );
  INV_X4 U15862 ( .I(n1606), .ZN(n9547) );
  INV_X2 U3705 ( .I(n33997), .ZN(n1107) );
  AOI21_X2 U4444 ( .A1(n14810), .A2(n26110), .B(n33753), .ZN(n33752) );
  BUF_X2 U4243 ( .I(n21857), .Z(n455) );
  INV_X2 U5548 ( .I(n26018), .ZN(n1239) );
  INV_X2 U1911 ( .I(n24732), .ZN(n24839) );
  INV_X2 U17362 ( .I(n20208), .ZN(n35180) );
  OAI21_X2 U15281 ( .A1(n2812), .A2(n38748), .B(n36210), .ZN(n2813) );
  OAI21_X2 U27275 ( .A1(n21588), .A2(n19397), .B(n17792), .ZN(n18560) );
  BUF_X2 U10447 ( .I(Key[143]), .Z(n29647) );
  BUF_X2 U3165 ( .I(n21270), .Z(n32720) );
  BUF_X4 U4868 ( .I(n5988), .Z(n36854) );
  NAND2_X2 U20147 ( .A1(n32041), .A2(n32040), .ZN(n23065) );
  INV_X2 U13343 ( .I(n4847), .ZN(n33893) );
  INV_X4 U6306 ( .I(n19915), .ZN(n1127) );
  NAND2_X2 U17411 ( .A1(n22342), .A2(n17074), .ZN(n21966) );
  INV_X2 U6507 ( .I(n17074), .ZN(n22171) );
  AOI21_X2 U6718 ( .A1(n22803), .A2(n5657), .B(n8461), .ZN(n8460) );
  INV_X4 U20454 ( .I(n16200), .ZN(n10807) );
  INV_X4 U15541 ( .I(n585), .ZN(n5572) );
  AOI22_X2 U2249 ( .A1(n18606), .A2(n26740), .B1(n6615), .B2(n18706), .ZN(
        n30585) );
  NOR3_X2 U2754 ( .A1(n1417), .A2(n209), .A3(n1192), .ZN(n5156) );
  NOR2_X2 U8956 ( .A1(n27653), .A2(n11412), .ZN(n14237) );
  NAND2_X2 U5954 ( .A1(n978), .A2(n13508), .ZN(n32004) );
  AOI21_X2 U4693 ( .A1(n37737), .A2(n24746), .B(n32882), .ZN(n2549) );
  BUF_X2 U7489 ( .I(n8944), .Z(n36796) );
  AOI22_X2 U4614 ( .A1(n9352), .A2(n38566), .B1(n9353), .B2(n10618), .ZN(
        n33686) );
  BUF_X4 U2533 ( .I(n19712), .Z(n31157) );
  INV_X2 U30561 ( .I(n8556), .ZN(n2292) );
  NOR2_X2 U2712 ( .A1(n12702), .A2(n12703), .ZN(n56) );
  INV_X2 U19298 ( .I(n6591), .ZN(n19589) );
  INV_X4 U4899 ( .I(n14378), .ZN(n1597) );
  BUF_X4 U1065 ( .I(n18500), .Z(n17194) );
  NOR2_X1 U7256 ( .A1(n17617), .A2(n5405), .ZN(n36307) );
  INV_X2 U395 ( .I(n36791), .ZN(n13133) );
  NAND2_X2 U1267 ( .A1(n26119), .A2(n7423), .ZN(n35401) );
  NOR2_X2 U13658 ( .A1(n11012), .A2(n21965), .ZN(n9343) );
  NAND2_X2 U9987 ( .A1(n22959), .A2(n11157), .ZN(n11156) );
  NAND2_X1 U9197 ( .A1(n18730), .A2(n1331), .ZN(n31860) );
  OAI22_X1 U10552 ( .A1(n25363), .A2(n424), .B1(n9568), .B2(n26090), .ZN(
        n34413) );
  CLKBUF_X8 U12706 ( .I(n2634), .Z(n2340) );
  OAI21_X2 U25964 ( .A1(n12477), .A2(n13081), .B(n37057), .ZN(n36266) );
  OAI21_X2 U12801 ( .A1(n28590), .A2(n3598), .B(n14701), .ZN(n35961) );
  NAND2_X2 U8847 ( .A1(n31583), .A2(n37061), .ZN(n20371) );
  NAND3_X2 U3650 ( .A1(n32712), .A2(n27146), .A3(n27354), .ZN(n36492) );
  NOR2_X1 U30348 ( .A1(n9056), .A2(n154), .ZN(n36834) );
  OR3_X2 U13033 ( .A1(n18342), .A2(n12951), .A3(n11795), .Z(n7279) );
  BUF_X2 U1794 ( .I(n30454), .Z(n33240) );
  AOI22_X2 U2217 ( .A1(n23253), .A2(n23610), .B1(n9639), .B2(n1132), .ZN(
        n33702) );
  NOR2_X1 U18766 ( .A1(n32619), .A2(n32618), .ZN(n3761) );
  NAND2_X1 U8616 ( .A1(n23548), .A2(n23472), .ZN(n2688) );
  NOR2_X2 U1112 ( .A1(n6104), .A2(n6103), .ZN(n6154) );
  OAI21_X1 U8261 ( .A1(n4531), .A2(n32703), .B(n32702), .ZN(n10640) );
  NAND2_X2 U19812 ( .A1(n15121), .A2(n1101), .ZN(n7135) );
  INV_X2 U179 ( .I(n36595), .ZN(n3633) );
  INV_X4 U128 ( .I(n37100), .ZN(n29446) );
  NOR3_X2 U2343 ( .A1(n14396), .A2(n19538), .A3(n31093), .ZN(n35564) );
  BUF_X2 U3860 ( .I(n29307), .Z(n29498) );
  OR2_X2 U689 ( .A1(n27108), .A2(n6686), .Z(n30434) );
  OR2_X2 U13020 ( .A1(n10733), .A2(n14290), .Z(n15775) );
  NAND2_X2 U1290 ( .A1(n32436), .A2(n260), .ZN(n31964) );
  NAND2_X2 U21579 ( .A1(n35665), .A2(n34087), .ZN(n32436) );
  INV_X4 U23324 ( .I(n12066), .ZN(n12065) );
  NAND2_X1 U26021 ( .A1(n33054), .A2(n33052), .ZN(n33051) );
  INV_X2 U6860 ( .I(n17915), .ZN(n1528) );
  NAND2_X2 U28144 ( .A1(n19238), .A2(n17112), .ZN(n21511) );
  INV_X2 U7081 ( .I(n32377), .ZN(n23579) );
  INV_X2 U908 ( .I(n10987), .ZN(n3426) );
  INV_X2 U27577 ( .I(n16835), .ZN(n19334) );
  NAND2_X2 U1664 ( .A1(n32831), .A2(n24878), .ZN(n8125) );
  OAI21_X2 U12267 ( .A1(n25687), .A2(n25686), .B(n25685), .ZN(n20008) );
  NOR2_X2 U7494 ( .A1(n11412), .A2(n11164), .ZN(n11163) );
  NOR2_X1 U20357 ( .A1(n32950), .A2(n6534), .ZN(n35466) );
  CLKBUF_X4 U3496 ( .I(n9847), .Z(n2018) );
  INV_X1 U17621 ( .I(n38199), .ZN(n26754) );
  BUF_X4 U3984 ( .I(n33987), .Z(n33986) );
  OAI21_X2 U9688 ( .A1(n19027), .A2(n13026), .B(n19026), .ZN(n23754) );
  NAND2_X2 U5631 ( .A1(n26696), .A2(n923), .ZN(n4583) );
  NOR2_X2 U21152 ( .A1(n17040), .A2(n7730), .ZN(n8682) );
  NAND2_X2 U1128 ( .A1(n20088), .A2(n26021), .ZN(n33423) );
  NAND2_X2 U3975 ( .A1(n34969), .A2(n8537), .ZN(n13364) );
  NOR2_X2 U1347 ( .A1(n37238), .A2(n5798), .ZN(n13034) );
  INV_X2 U2416 ( .I(n12909), .ZN(n14461) );
  NAND2_X1 U3919 ( .A1(n27114), .A2(n33088), .ZN(n32757) );
  NAND2_X2 U1313 ( .A1(n8006), .A2(n17008), .ZN(n7941) );
  INV_X2 U9327 ( .I(n1091), .ZN(n10890) );
  INV_X2 U7490 ( .I(n15187), .ZN(n18667) );
  CLKBUF_X4 U2709 ( .I(n22854), .Z(n22993) );
  BUF_X2 U7310 ( .I(Key[51]), .Z(n29223) );
  INV_X1 U5332 ( .I(n37916), .ZN(n1279) );
  OAI21_X2 U313 ( .A1(n20188), .A2(n33842), .B(n21239), .ZN(n14330) );
  OAI21_X2 U4042 ( .A1(n1112), .A2(n7866), .B(n33950), .ZN(n11332) );
  INV_X4 U8188 ( .I(n25692), .ZN(n1112) );
  NAND2_X2 U5006 ( .A1(n21806), .A2(n36735), .ZN(n21274) );
  AOI21_X2 U11830 ( .A1(n3125), .A2(n35960), .B(n3124), .ZN(n35022) );
  NOR2_X2 U2610 ( .A1(n123), .A2(n19545), .ZN(n9041) );
  NAND2_X2 U3623 ( .A1(n22080), .A2(n38337), .ZN(n4337) );
  INV_X2 U10888 ( .I(n11573), .ZN(n30220) );
  INV_X2 U13567 ( .I(n20077), .ZN(n1653) );
  NAND3_X1 U7002 ( .A1(n24269), .A2(n24444), .A3(n24311), .ZN(n11104) );
  AOI21_X2 U272 ( .A1(n27996), .A2(n16461), .B(n27995), .ZN(n28002) );
  NOR2_X2 U4425 ( .A1(n2078), .A2(n3541), .ZN(n2077) );
  INV_X1 U8187 ( .I(n37604), .ZN(n32634) );
  NAND2_X2 U22313 ( .A1(n17501), .A2(n32747), .ZN(n10224) );
  AND3_X1 U4090 ( .A1(n24812), .A2(n24565), .A3(n19294), .Z(n14532) );
  INV_X4 U840 ( .I(n25487), .ZN(n1535) );
  INV_X2 U2320 ( .I(n23296), .ZN(n35808) );
  AOI21_X1 U5454 ( .A1(n15372), .A2(n28220), .B(n11650), .ZN(n11649) );
  CLKBUF_X2 U14028 ( .I(Key[44]), .Z(n30090) );
  INV_X2 U14385 ( .I(n2000), .ZN(n13758) );
  NOR2_X2 U12324 ( .A1(n8222), .A2(n7866), .ZN(n8221) );
  NAND2_X2 U25311 ( .A1(n28361), .A2(n28362), .ZN(n18836) );
  NOR2_X2 U8719 ( .A1(n14499), .A2(n8597), .ZN(n8599) );
  INV_X4 U6769 ( .I(n14488), .ZN(n26823) );
  NAND2_X1 U16404 ( .A1(n35447), .A2(n20306), .ZN(n36972) );
  NOR2_X2 U1918 ( .A1(n17120), .A2(n9996), .ZN(n12669) );
  AOI21_X2 U6267 ( .A1(n1267), .A2(n2341), .B(n1576), .ZN(n6636) );
  OAI21_X2 U11337 ( .A1(n15313), .A2(n28720), .B(n37311), .ZN(n15312) );
  NOR2_X2 U4439 ( .A1(n25586), .A2(n10062), .ZN(n32157) );
  INV_X2 U12668 ( .I(n18110), .ZN(n16211) );
  NAND2_X2 U16802 ( .A1(n4345), .A2(n9201), .ZN(n3998) );
  NAND2_X2 U3892 ( .A1(n16922), .A2(n16921), .ZN(n16920) );
  AOI22_X2 U9048 ( .A1(n19139), .A2(n1446), .B1(n20577), .B2(n28111), .ZN(
        n18309) );
  INV_X2 U13295 ( .I(n23347), .ZN(n10048) );
  CLKBUF_X4 U8382 ( .I(n10162), .Z(n36422) );
  CLKBUF_X4 U2872 ( .I(n28704), .Z(n18281) );
  BUF_X2 U2457 ( .I(n22887), .Z(n31300) );
  BUF_X4 U6118 ( .I(n9878), .Z(n2937) );
  NOR2_X2 U4395 ( .A1(n19777), .A2(n5698), .ZN(n17841) );
  INV_X2 U5785 ( .I(n18246), .ZN(n19564) );
  AOI22_X2 U20025 ( .A1(n16105), .A2(n16104), .B1(n1316), .B2(n20173), .ZN(
        n7366) );
  NOR2_X2 U4360 ( .A1(n7320), .A2(n26304), .ZN(n31274) );
  NAND2_X2 U15070 ( .A1(n6446), .A2(n27070), .ZN(n34944) );
  INV_X1 U11969 ( .I(n26358), .ZN(n4591) );
  CLKBUF_X2 U7592 ( .I(n14422), .Z(n357) );
  NOR2_X2 U8865 ( .A1(n9394), .A2(n5669), .ZN(n30190) );
  INV_X2 U6442 ( .I(n3443), .ZN(n9316) );
  NAND3_X1 U2967 ( .A1(n4919), .A2(n16985), .A3(n20480), .ZN(n32188) );
  INV_X2 U9530 ( .I(n12394), .ZN(n1536) );
  NAND2_X2 U12314 ( .A1(n25444), .A2(n38338), .ZN(n9503) );
  NAND2_X2 U9962 ( .A1(n2049), .A2(n1989), .ZN(n5944) );
  INV_X2 U13802 ( .I(n17869), .ZN(n17207) );
  INV_X2 U16333 ( .I(n5080), .ZN(n25328) );
  INV_X2 U6419 ( .I(n21923), .ZN(n1689) );
  NOR2_X2 U5402 ( .A1(n37852), .A2(n8954), .ZN(n8968) );
  BUF_X4 U28226 ( .I(n16760), .Z(n33359) );
  NOR2_X2 U2625 ( .A1(n4759), .A2(n21888), .ZN(n21601) );
  NAND2_X2 U2505 ( .A1(n22342), .A2(n22341), .ZN(n10487) );
  NOR3_X2 U2009 ( .A1(n17127), .A2(n1989), .A3(n37791), .ZN(n33034) );
  NOR2_X2 U7099 ( .A1(n26135), .A2(n31626), .ZN(n15449) );
  NAND2_X2 U5287 ( .A1(n15240), .A2(n1608), .ZN(n20083) );
  INV_X2 U565 ( .I(n33960), .ZN(n32977) );
  OR2_X2 U1185 ( .A1(n34609), .A2(n4553), .Z(n25916) );
  INV_X4 U1936 ( .I(n1140), .ZN(n32061) );
  AOI22_X2 U11230 ( .A1(n28759), .A2(n18701), .B1(n1416), .B2(n30917), .ZN(
        n28761) );
  OAI21_X1 U21369 ( .A1(n29741), .A2(n29754), .B(n29737), .ZN(n29726) );
  INV_X2 U18388 ( .I(n17567), .ZN(n17784) );
  INV_X4 U6545 ( .I(n11329), .ZN(n8520) );
  NAND2_X2 U20121 ( .A1(n7062), .A2(n32456), .ZN(n21794) );
  OAI21_X2 U3701 ( .A1(n923), .A2(n37102), .B(n26695), .ZN(n16707) );
  NOR2_X2 U12116 ( .A1(n25758), .A2(n33514), .ZN(n2498) );
  INV_X2 U17498 ( .I(n27786), .ZN(n18733) );
  NOR2_X2 U7434 ( .A1(n36197), .A2(n28278), .ZN(n7840) );
  BUF_X4 U27642 ( .I(n18342), .Z(n33289) );
  NAND2_X2 U7461 ( .A1(n18461), .A2(n38262), .ZN(n18457) );
  NAND2_X2 U24181 ( .A1(n19043), .A2(n17714), .ZN(n13890) );
  INV_X1 U15745 ( .I(n14130), .ZN(n23178) );
  INV_X1 U30764 ( .I(n36995), .ZN(n30338) );
  AOI21_X2 U6813 ( .A1(n9892), .A2(n931), .B(n7460), .ZN(n24968) );
  NAND3_X1 U12532 ( .A1(n18264), .A2(n24413), .A3(n18263), .ZN(n24415) );
  NOR2_X2 U1208 ( .A1(n32044), .A2(n2957), .ZN(n2955) );
  NAND2_X2 U8260 ( .A1(n1028), .A2(n24782), .ZN(n13415) );
  INV_X2 U16321 ( .I(n9385), .ZN(n14211) );
  INV_X2 U1072 ( .I(n18238), .ZN(n1591) );
  OAI21_X2 U13291 ( .A1(n8459), .A2(n8458), .B(n19469), .ZN(n4698) );
  AOI21_X2 U28818 ( .A1(n34906), .A2(n24732), .B(n4973), .ZN(n24254) );
  BUF_X2 U11861 ( .I(n27141), .Z(n9593) );
  NOR2_X2 U1975 ( .A1(n5942), .A2(n5943), .ZN(n5946) );
  NAND2_X2 U12443 ( .A1(n25467), .A2(n38210), .ZN(n14679) );
  NAND2_X1 U8096 ( .A1(n17038), .A2(n17020), .ZN(n17037) );
  OAI21_X2 U16531 ( .A1(n1689), .A2(n9316), .B(n37612), .ZN(n4057) );
  NAND2_X2 U7438 ( .A1(n28214), .A2(n11512), .ZN(n18020) );
  NAND2_X2 U22803 ( .A1(n8385), .A2(n11083), .ZN(n13178) );
  AOI21_X2 U17154 ( .A1(n7767), .A2(n17212), .B(n834), .ZN(n25772) );
  NAND3_X2 U4221 ( .A1(n36638), .A2(n33247), .A3(n3683), .ZN(n31343) );
  INV_X2 U8352 ( .I(n14491), .ZN(n24453) );
  NOR2_X2 U2174 ( .A1(n37190), .A2(n34981), .ZN(n4538) );
  NOR2_X2 U24744 ( .A1(n33709), .A2(n15879), .ZN(n7625) );
  OAI21_X2 U8959 ( .A1(n33424), .A2(n18035), .B(n11030), .ZN(n4926) );
  NAND2_X1 U495 ( .A1(n27981), .A2(n28047), .ZN(n36914) );
  INV_X1 U27151 ( .I(n36755), .ZN(n36433) );
  INV_X2 U27903 ( .I(n20958), .ZN(n23076) );
  NOR2_X1 U3087 ( .A1(n18884), .A2(n8480), .ZN(n16642) );
  INV_X2 U4737 ( .I(n23198), .ZN(n1044) );
  OR2_X1 U12043 ( .A1(n19137), .A2(n16510), .Z(n10148) );
  NOR2_X2 U11727 ( .A1(n4927), .A2(n34569), .ZN(n32206) );
  AOI22_X2 U21872 ( .A1(n18822), .A2(n22892), .B1(n13946), .B2(n22804), .ZN(
        n32397) );
  NOR2_X2 U13287 ( .A1(n30386), .A2(n3761), .ZN(n36729) );
  NAND2_X2 U6369 ( .A1(n19375), .A2(n34923), .ZN(n21778) );
  NAND2_X2 U5621 ( .A1(n34658), .A2(n26316), .ZN(n31253) );
  NOR2_X2 U12843 ( .A1(n6914), .A2(n6170), .ZN(n6913) );
  INV_X4 U347 ( .I(n20860), .ZN(n7872) );
  NOR2_X2 U10032 ( .A1(n31005), .A2(n20872), .ZN(n16892) );
  INV_X1 U17394 ( .I(n26905), .ZN(n15485) );
  AOI21_X2 U19238 ( .A1(n23174), .A2(n3803), .B(n20840), .ZN(n11157) );
  AOI21_X1 U11937 ( .A1(n38548), .A2(n14212), .B(n25951), .ZN(n12869) );
  INV_X1 U7198 ( .I(n735), .ZN(n26470) );
  BUF_X2 U4473 ( .I(n18062), .Z(n31719) );
  INV_X2 U1738 ( .I(n37395), .ZN(n34746) );
  NAND2_X2 U7826 ( .A1(n7612), .A2(n5035), .ZN(n5366) );
  INV_X1 U15781 ( .I(n33995), .ZN(n31513) );
  NAND2_X2 U26689 ( .A1(n5366), .A2(n5367), .ZN(n5361) );
  NOR2_X2 U14613 ( .A1(n9587), .A2(n9588), .ZN(n34884) );
  AOI21_X1 U18928 ( .A1(n2681), .A2(n38248), .B(n31836), .ZN(n2684) );
  AOI21_X2 U6010 ( .A1(n17793), .A2(n22108), .B(n1684), .ZN(n12155) );
  INV_X2 U24726 ( .I(n22272), .ZN(n15029) );
  NAND2_X2 U23396 ( .A1(n17167), .A2(n12191), .ZN(n23334) );
  OAI21_X2 U22203 ( .A1(n14392), .A2(n24184), .B(n35690), .ZN(n10046) );
  NAND3_X2 U2221 ( .A1(n23494), .A2(n33638), .A3(n36630), .ZN(n23500) );
  INV_X2 U575 ( .I(n38002), .ZN(n26840) );
  NAND2_X2 U2063 ( .A1(n37216), .A2(n36227), .ZN(n31168) );
  INV_X4 U1261 ( .I(n23399), .ZN(n961) );
  NAND3_X1 U9189 ( .A1(n28042), .A2(n28043), .A3(n1073), .ZN(n36832) );
  NOR2_X1 U1310 ( .A1(n832), .A2(n14778), .ZN(n30945) );
  NAND2_X2 U11875 ( .A1(n6909), .A2(n35537), .ZN(n12566) );
  NOR3_X2 U29184 ( .A1(n26240), .A2(n26239), .A3(n26238), .ZN(n26439) );
  NAND2_X2 U6654 ( .A1(n18948), .A2(n15925), .ZN(n18696) );
  OAI21_X2 U29248 ( .A1(n33689), .A2(n37585), .B(n26444), .ZN(n26445) );
  AOI21_X2 U2930 ( .A1(n14382), .A2(n19728), .B(n1500), .ZN(n26444) );
  NOR2_X2 U6647 ( .A1(n16638), .A2(n22993), .ZN(n34643) );
  OR2_X2 U2116 ( .A1(n30280), .A2(n31278), .Z(n15018) );
  OAI21_X2 U506 ( .A1(n7934), .A2(n8498), .B(n28045), .ZN(n27988) );
  NOR2_X2 U21197 ( .A1(n27507), .A2(n35265), .ZN(n35604) );
  NAND2_X2 U11492 ( .A1(n8092), .A2(n8093), .ZN(n34525) );
  OAI22_X2 U29054 ( .A1(n33428), .A2(n33427), .B1(n29536), .B2(n29519), .ZN(
        n29510) );
  NAND3_X2 U24877 ( .A1(n24118), .A2(n24372), .A3(n38609), .ZN(n14895) );
  INV_X2 U5915 ( .I(n26541), .ZN(n16169) );
  BUF_X4 U18303 ( .I(n38669), .Z(n31088) );
  INV_X2 U17576 ( .I(n4841), .ZN(n28238) );
  NOR2_X2 U9581 ( .A1(n35000), .A2(n33640), .ZN(n2328) );
  NOR2_X2 U8854 ( .A1(n17374), .A2(n19120), .ZN(n13388) );
  NOR2_X2 U20065 ( .A1(n5415), .A2(n8112), .ZN(n33281) );
  AOI21_X2 U6554 ( .A1(n12353), .A2(n5669), .B(n30155), .ZN(n8112) );
  OAI21_X2 U15056 ( .A1(n32802), .A2(n37097), .B(n2608), .ZN(n2607) );
  NAND2_X2 U13252 ( .A1(n14739), .A2(n8146), .ZN(n8145) );
  INV_X2 U2413 ( .I(n30304), .ZN(n8093) );
  AOI21_X1 U12285 ( .A1(n33826), .A2(n19237), .B(n19236), .ZN(n17868) );
  NAND2_X2 U2201 ( .A1(n3497), .A2(n15787), .ZN(n36394) );
  OAI21_X2 U8423 ( .A1(n23624), .A2(n35938), .B(n3498), .ZN(n3497) );
  OAI22_X2 U3992 ( .A1(n10906), .A2(n36663), .B1(n18871), .B2(n10883), .ZN(
        n28314) );
  AOI22_X2 U3396 ( .A1(n14484), .A2(n19366), .B1(n28148), .B2(n18392), .ZN(
        n30608) );
  NOR2_X2 U8398 ( .A1(n1298), .A2(n32351), .ZN(n5790) );
  AOI22_X2 U16680 ( .A1(n12544), .A2(n12543), .B1(n36145), .B2(n18961), .ZN(
        n12542) );
  BUF_X4 U20222 ( .I(n30504), .Z(n35443) );
  AOI22_X2 U13147 ( .A1(n8390), .A2(n32858), .B1(n23421), .B2(n1302), .ZN(
        n7482) );
  BUF_X2 U17287 ( .I(n36397), .Z(n35754) );
  OAI21_X1 U4688 ( .A1(n24626), .A2(n24627), .B(n9847), .ZN(n13747) );
  INV_X2 U28297 ( .I(n9736), .ZN(n22334) );
  INV_X2 U15163 ( .I(n7324), .ZN(n31353) );
  NAND2_X2 U26622 ( .A1(n26964), .A2(n26963), .ZN(n17602) );
  NAND3_X2 U1073 ( .A1(n30665), .A2(n35537), .A3(n1231), .ZN(n26963) );
  INV_X4 U27859 ( .I(n21939), .ZN(n36519) );
  NAND2_X1 U4458 ( .A1(n27011), .A2(n16263), .ZN(n8196) );
  OAI21_X2 U12784 ( .A1(n6175), .A2(n10690), .B(n9844), .ZN(n16406) );
  NAND2_X2 U26478 ( .A1(n5351), .A2(n36325), .ZN(n7325) );
  INV_X1 U1344 ( .I(n23102), .ZN(n23103) );
  INV_X2 U17540 ( .I(n29555), .ZN(n29541) );
  OAI22_X2 U6705 ( .A1(n22809), .A2(n36554), .B1(n531), .B2(n23169), .ZN(
        n22812) );
  NOR2_X2 U23409 ( .A1(n16081), .A2(n24373), .ZN(n24191) );
  NAND2_X2 U671 ( .A1(n26084), .A2(n26114), .ZN(n4372) );
  INV_X4 U3287 ( .I(n14729), .ZN(n1577) );
  INV_X2 U29245 ( .I(n26439), .ZN(n26440) );
  BUF_X4 U1801 ( .I(n39816), .Z(n250) );
  INV_X1 U30574 ( .I(n23654), .ZN(n238) );
  INV_X2 U7060 ( .I(n23599), .ZN(n23601) );
  INV_X2 U5864 ( .I(n20896), .ZN(n941) );
  AOI22_X2 U2590 ( .A1(n8434), .A2(n21834), .B1(n8436), .B2(n21436), .ZN(
        n34220) );
  INV_X2 U25457 ( .I(n25716), .ZN(n25562) );
  NAND2_X2 U2977 ( .A1(n23308), .A2(n38704), .ZN(n23311) );
  AOI21_X2 U5697 ( .A1(n24708), .A2(n24529), .B(n33986), .ZN(n8389) );
  NOR2_X2 U12187 ( .A1(n26079), .A2(n15283), .ZN(n7170) );
  AOI21_X2 U19536 ( .A1(n30702), .A2(n28133), .B(n2870), .ZN(n3070) );
  NAND2_X1 U5437 ( .A1(n4874), .A2(n13837), .ZN(n6556) );
  OR2_X1 U10037 ( .A1(n1484), .A2(n32870), .Z(n16480) );
  INV_X2 U9587 ( .I(n24944), .ZN(n13259) );
  INV_X4 U1339 ( .I(n34014), .ZN(n9050) );
  INV_X4 U105 ( .I(n8805), .ZN(n3986) );
  NOR2_X1 U19058 ( .A1(n20915), .A2(n14692), .ZN(n20914) );
  NOR2_X1 U860 ( .A1(n20815), .A2(n35271), .ZN(n219) );
  BUF_X4 U12684 ( .I(n8805), .Z(n34652) );
  NOR2_X1 U14559 ( .A1(n4459), .A2(n2140), .ZN(n10903) );
  NOR2_X2 U19714 ( .A1(n32543), .A2(n28486), .ZN(n8657) );
  NAND2_X2 U1916 ( .A1(n31945), .A2(n30506), .ZN(n32598) );
  NOR2_X2 U866 ( .A1(n13427), .A2(n4686), .ZN(n27044) );
  BUF_X2 U1558 ( .I(n24819), .Z(n31714) );
  AOI22_X2 U541 ( .A1(n13984), .A2(n27969), .B1(n12257), .B2(n13983), .ZN(
        n14277) );
  NAND3_X2 U27587 ( .A1(n24906), .A2(n32802), .A3(n24905), .ZN(n24907) );
  INV_X2 U4035 ( .I(n18302), .ZN(n20058) );
  NAND2_X2 U4111 ( .A1(n21117), .A2(n38448), .ZN(n2128) );
  INV_X2 U1726 ( .I(n20774), .ZN(n1209) );
  NAND2_X2 U183 ( .A1(n6163), .A2(n8805), .ZN(n29992) );
  BUF_X2 U18027 ( .I(Key[99]), .Z(n30094) );
  CLKBUF_X4 U17379 ( .I(n14462), .Z(n12443) );
  CLKBUF_X4 U4082 ( .I(n9383), .Z(n1606) );
  INV_X2 U1064 ( .I(n39648), .ZN(n7658) );
  INV_X2 U17193 ( .I(n33316), .ZN(n36965) );
  INV_X2 U6800 ( .I(n9214), .ZN(n26901) );
  NOR2_X2 U780 ( .A1(n27273), .A2(n27274), .ZN(n8382) );
  INV_X1 U10909 ( .I(n7766), .ZN(n28947) );
  BUF_X2 U6603 ( .I(n15871), .Z(n35532) );
  NOR2_X1 U11801 ( .A1(n7393), .A2(n7392), .ZN(n14966) );
  NOR2_X2 U23787 ( .A1(n10806), .A2(n39571), .ZN(n32727) );
  NAND2_X2 U17347 ( .A1(n33116), .A2(n8272), .ZN(n35529) );
  OAI21_X2 U226 ( .A1(n18096), .A2(n37295), .B(n5662), .ZN(n19726) );
  INV_X2 U10110 ( .I(n23140), .ZN(n22949) );
  AOI21_X2 U2766 ( .A1(n25365), .A2(n25623), .B(n1532), .ZN(n3012) );
  INV_X2 U7106 ( .I(n25856), .ZN(n26008) );
  NAND2_X1 U20992 ( .A1(n32215), .A2(n15411), .ZN(n11222) );
  NOR2_X2 U6973 ( .A1(n24824), .A2(n24819), .ZN(n24629) );
  OAI21_X2 U26800 ( .A1(n32425), .A2(n38292), .B(n38042), .ZN(n23328) );
  NAND3_X2 U15239 ( .A1(n16520), .A2(n27406), .A3(n2947), .ZN(n16516) );
  INV_X2 U13676 ( .I(n22352), .ZN(n4993) );
  OAI21_X2 U29724 ( .A1(n24509), .A2(n14213), .B(n24799), .ZN(n7396) );
  OAI21_X2 U24157 ( .A1(n1038), .A2(n32424), .B(n1635), .ZN(n15702) );
  INV_X2 U28768 ( .I(n25797), .ZN(n25912) );
  OR3_X1 U4633 ( .A1(n38168), .A2(n35855), .A3(n14375), .Z(n13282) );
  NAND3_X2 U28682 ( .A1(n34494), .A2(n37279), .A3(n17927), .ZN(n23627) );
  INV_X2 U6053 ( .I(n24257), .ZN(n36342) );
  NOR2_X2 U9069 ( .A1(n30431), .A2(n30714), .ZN(n11026) );
  NOR2_X2 U4789 ( .A1(n20968), .A2(n20967), .ZN(n20966) );
  INV_X2 U3773 ( .I(n32601), .ZN(n23477) );
  OAI21_X1 U1481 ( .A1(n18593), .A2(n18592), .B(n21431), .ZN(n18591) );
  NAND2_X1 U14791 ( .A1(n26945), .A2(n34908), .ZN(n35613) );
  NAND3_X2 U80 ( .A1(n481), .A2(n29776), .A3(n34914), .ZN(n9063) );
  NAND3_X2 U10253 ( .A1(n8869), .A2(n8491), .A3(n18865), .ZN(n30815) );
  NOR3_X2 U2098 ( .A1(n6849), .A2(n20537), .A3(n24469), .ZN(n34366) );
  OAI21_X1 U20236 ( .A1(n20305), .A2(n28064), .B(n21239), .ZN(n35447) );
  OAI21_X2 U2177 ( .A1(n34996), .A2(n7333), .B(n38292), .ZN(n14012) );
  NAND3_X1 U21960 ( .A1(n37210), .A2(n24387), .A3(n31714), .ZN(n4938) );
  NOR2_X2 U21714 ( .A1(n32359), .A2(n972), .ZN(n6649) );
  OAI21_X2 U14587 ( .A1(n22843), .A2(n19865), .B(n2163), .ZN(n22456) );
  AOI22_X2 U6014 ( .A1(n28425), .A2(n39724), .B1(n9935), .B2(n10906), .ZN(
        n30748) );
  INV_X2 U7830 ( .I(n27399), .ZN(n1473) );
  BUF_X2 U3516 ( .I(n22802), .Z(n272) );
  INV_X2 U6318 ( .I(n12612), .ZN(n24116) );
  NOR2_X1 U21797 ( .A1(n24822), .A2(n13214), .ZN(n24823) );
  NAND2_X1 U5709 ( .A1(n25854), .A2(n36048), .ZN(n15919) );
  NOR2_X2 U5016 ( .A1(n1686), .A2(n3644), .ZN(n21421) );
  NOR2_X2 U9890 ( .A1(n10174), .A2(n13150), .ZN(n15624) );
  INV_X2 U5467 ( .I(n7324), .ZN(n1197) );
  NAND2_X2 U18205 ( .A1(n28418), .A2(n9169), .ZN(n18378) );
  NOR2_X2 U1466 ( .A1(n11851), .A2(n543), .ZN(n6671) );
  NAND2_X2 U24299 ( .A1(n17577), .A2(n14196), .ZN(n17576) );
  OAI21_X2 U13758 ( .A1(n2458), .A2(n18408), .B(n16511), .ZN(n17577) );
  NOR2_X2 U14811 ( .A1(n35782), .A2(n24406), .ZN(n35781) );
  INV_X4 U22230 ( .I(n6684), .ZN(n19869) );
  NAND2_X1 U1921 ( .A1(n31267), .A2(n36157), .ZN(n34438) );
  INV_X4 U6240 ( .I(n16043), .ZN(n15276) );
  NOR2_X1 U871 ( .A1(n14989), .A2(n3402), .ZN(n14988) );
  NAND3_X1 U8387 ( .A1(n3048), .A2(n15123), .A3(n9924), .ZN(n15324) );
  NAND2_X2 U1037 ( .A1(n24118), .A2(n24372), .ZN(n24430) );
  INV_X4 U5143 ( .I(n22709), .ZN(n1650) );
  NAND2_X2 U30763 ( .A1(n31574), .A2(n39389), .ZN(n13537) );
  INV_X2 U3625 ( .I(n293), .ZN(n21917) );
  NOR2_X2 U15421 ( .A1(n2439), .A2(n2975), .ZN(n2974) );
  NOR2_X2 U7204 ( .A1(n22287), .A2(n22197), .ZN(n22134) );
  NAND2_X1 U8827 ( .A1(n9046), .A2(n35405), .ZN(n9045) );
  NAND2_X2 U2245 ( .A1(n8964), .A2(n35536), .ZN(n8138) );
  AOI22_X2 U2512 ( .A1(n23215), .A2(n23413), .B1(n23412), .B2(n6421), .ZN(
        n18381) );
  NAND3_X1 U7610 ( .A1(n30136), .A2(n34177), .A3(n18588), .ZN(n31258) );
  NAND3_X2 U13474 ( .A1(n23068), .A2(n3906), .A3(n37984), .ZN(n11366) );
  OAI22_X2 U1192 ( .A1(n25916), .A2(n34265), .B1(n26034), .B2(n37300), .ZN(
        n12708) );
  OAI21_X2 U24789 ( .A1(n22962), .A2(n39303), .B(n22816), .ZN(n19528) );
  NAND2_X2 U29311 ( .A1(n26777), .A2(n32256), .ZN(n26778) );
  NOR2_X2 U8390 ( .A1(n32858), .A2(n5487), .ZN(n21208) );
  OAI22_X2 U12561 ( .A1(n7938), .A2(n31055), .B1(n30345), .B2(n33864), .ZN(
        n3348) );
  AOI21_X2 U3652 ( .A1(n13150), .A2(n32377), .B(n1626), .ZN(n10613) );
  INV_X2 U15442 ( .I(n23226), .ZN(n31332) );
  OAI21_X2 U3132 ( .A1(n32425), .A2(n6637), .B(n6639), .ZN(n6994) );
  AOI21_X2 U6726 ( .A1(n6638), .A2(n6637), .B(n30881), .ZN(n6639) );
  NAND2_X2 U253 ( .A1(n36814), .A2(n27907), .ZN(n12312) );
  NAND2_X2 U2134 ( .A1(n22150), .A2(n33678), .ZN(n16511) );
  INV_X2 U17799 ( .I(n33937), .ZN(n18455) );
  INV_X2 U4824 ( .I(n22465), .ZN(n30322) );
  INV_X4 U6218 ( .I(n25962), .ZN(n25803) );
  NAND2_X1 U2340 ( .A1(n27374), .A2(n27373), .ZN(n27375) );
  INV_X1 U23915 ( .I(n11636), .ZN(n1095) );
  INV_X1 U2805 ( .I(n29087), .ZN(n6675) );
  NAND3_X1 U8640 ( .A1(n3333), .A2(n39507), .A3(n13065), .ZN(n3332) );
  INV_X2 U2049 ( .I(n22528), .ZN(n22454) );
  INV_X2 U23222 ( .I(n26249), .ZN(n36801) );
  AOI21_X2 U17959 ( .A1(n10857), .A2(n38275), .B(n32075), .ZN(n10856) );
  INV_X1 U23093 ( .I(n686), .ZN(n35881) );
  OAI21_X2 U10687 ( .A1(n8717), .A2(n8716), .B(n29183), .ZN(n20219) );
  NAND2_X2 U7123 ( .A1(n22803), .A2(n37883), .ZN(n4439) );
  NOR2_X2 U12807 ( .A1(n24293), .A2(n24295), .ZN(n13809) );
  OAI21_X2 U3725 ( .A1(n25401), .A2(n37926), .B(n16234), .ZN(n24937) );
  INV_X2 U18040 ( .I(n22263), .ZN(n19471) );
  NAND2_X1 U21490 ( .A1(n841), .A2(n25495), .ZN(n19311) );
  NAND2_X2 U16658 ( .A1(n38483), .A2(n26970), .ZN(n4171) );
  BUF_X4 U5655 ( .I(n37054), .Z(n1786) );
  NOR2_X2 U8583 ( .A1(n37217), .A2(n2186), .ZN(n11508) );
  NOR2_X1 U3883 ( .A1(n27420), .A2(n31287), .ZN(n13793) );
  NAND2_X2 U13722 ( .A1(n10433), .A2(n35019), .ZN(n4122) );
  NOR3_X2 U13184 ( .A1(n5380), .A2(n34014), .A3(n22958), .ZN(n34716) );
  INV_X2 U21107 ( .I(n14383), .ZN(n14382) );
  NAND2_X2 U10184 ( .A1(n22132), .A2(n37217), .ZN(n22029) );
  NAND2_X1 U26315 ( .A1(n16146), .A2(n34720), .ZN(n16147) );
  NAND2_X2 U6563 ( .A1(n14037), .A2(n14038), .ZN(n14036) );
  OAI21_X2 U3351 ( .A1(n29760), .A2(n29764), .B(n29762), .ZN(n17540) );
  INV_X2 U1232 ( .I(n25702), .ZN(n16072) );
  NAND2_X2 U4185 ( .A1(n38408), .A2(n1627), .ZN(n8146) );
  NOR2_X1 U12242 ( .A1(n8689), .A2(n25723), .ZN(n7239) );
  NAND2_X2 U7052 ( .A1(n20450), .A2(n1627), .ZN(n5839) );
  BUF_X4 U9237 ( .I(n14015), .Z(n2761) );
  OR2_X2 U3942 ( .A1(n14481), .A2(n19963), .Z(n25685) );
  AOI21_X2 U26215 ( .A1(n24472), .A2(n19818), .B(n33085), .ZN(n20378) );
  NAND2_X1 U11896 ( .A1(n18946), .A2(n6606), .ZN(n8019) );
  AOI21_X2 U27342 ( .A1(n20150), .A2(n18743), .B(n38079), .ZN(n20149) );
  NAND2_X2 U15367 ( .A1(n31390), .A2(n31389), .ZN(n28435) );
  NAND2_X2 U1287 ( .A1(n1044), .A2(n38282), .ZN(n5658) );
  NOR2_X2 U3646 ( .A1(n2451), .A2(n33396), .ZN(n6313) );
  AND2_X1 U27520 ( .A1(n14583), .A2(n11227), .Z(n36483) );
  NAND2_X2 U3353 ( .A1(n17105), .A2(n29764), .ZN(n28962) );
  OAI21_X2 U5792 ( .A1(n27319), .A2(n2304), .B(n1081), .ZN(n2303) );
  INV_X4 U3039 ( .I(n17105), .ZN(n29762) );
  NOR2_X2 U1403 ( .A1(n22115), .A2(n22114), .ZN(n22375) );
  OAI21_X2 U12854 ( .A1(n32590), .A2(n1312), .B(n31081), .ZN(n31080) );
  NOR2_X1 U8286 ( .A1(n7085), .A2(n7084), .ZN(n7083) );
  AOI21_X2 U11571 ( .A1(n27295), .A2(n39531), .B(n35485), .ZN(n27296) );
  NAND2_X1 U10518 ( .A1(n12321), .A2(n15840), .ZN(n12320) );
  NOR2_X2 U2246 ( .A1(n36430), .A2(n36431), .ZN(n36429) );
  NAND2_X2 U30203 ( .A1(n2127), .A2(n2128), .ZN(n36795) );
  NOR2_X1 U2076 ( .A1(n7504), .A2(n20109), .ZN(n20108) );
  OAI21_X2 U3381 ( .A1(n11095), .A2(n11468), .B(n38055), .ZN(n2933) );
  NAND2_X2 U17348 ( .A1(n33116), .A2(n8272), .ZN(n35255) );
  NAND3_X2 U28550 ( .A1(n23213), .A2(n14561), .A3(n4472), .ZN(n23510) );
  NAND2_X1 U23721 ( .A1(n35959), .A2(n35958), .ZN(n32394) );
  INV_X1 U7280 ( .I(n686), .ZN(n1352) );
  INV_X4 U6923 ( .I(n13300), .ZN(n19507) );
  NAND2_X2 U6154 ( .A1(n32740), .A2(n36422), .ZN(n30326) );
  BUF_X4 U7470 ( .I(n20453), .Z(n1399) );
  NOR2_X2 U16080 ( .A1(n24333), .A2(n14581), .ZN(n31484) );
  NAND2_X2 U333 ( .A1(n28221), .A2(n18841), .ZN(n19852) );
  NAND2_X2 U11741 ( .A1(n14135), .A2(n33689), .ZN(n14134) );
  NOR2_X1 U15969 ( .A1(n32808), .A2(n18274), .ZN(n19907) );
  NOR2_X2 U2346 ( .A1(n37984), .A2(n23143), .ZN(n23156) );
  NOR2_X2 U15653 ( .A1(n1118), .A2(n38794), .ZN(n12407) );
  OAI21_X1 U696 ( .A1(n35768), .A2(n35767), .B(n35766), .ZN(n27052) );
  NAND2_X1 U23016 ( .A1(n3430), .A2(n19765), .ZN(n10209) );
  INV_X2 U4293 ( .I(n14450), .ZN(n21498) );
  NOR2_X2 U8128 ( .A1(n25583), .A2(n1253), .ZN(n17815) );
  OAI22_X1 U4935 ( .A1(n7302), .A2(n7303), .B1(n29464), .B2(n9105), .ZN(n616)
         );
  OAI21_X2 U11900 ( .A1(n27226), .A2(n35427), .B(n11256), .ZN(n27228) );
  NAND2_X2 U11091 ( .A1(n28705), .A2(n31088), .ZN(n8272) );
  NOR3_X2 U1994 ( .A1(n18867), .A2(n35442), .A3(n1989), .ZN(n5943) );
  INV_X2 U12436 ( .I(n25625), .ZN(n1532) );
  NAND2_X2 U17686 ( .A1(n15803), .A2(n15802), .ZN(n15801) );
  INV_X2 U8358 ( .I(n6402), .ZN(n1131) );
  INV_X2 U23194 ( .I(n16039), .ZN(n20277) );
  NAND3_X2 U25228 ( .A1(n8674), .A2(n8673), .A3(n20872), .ZN(n33138) );
  NAND3_X2 U12360 ( .A1(n24943), .A2(n1112), .A3(n1531), .ZN(n12391) );
  NAND2_X2 U2104 ( .A1(n15175), .A2(n16635), .ZN(n17943) );
  NAND2_X1 U23638 ( .A1(n16982), .A2(n24214), .ZN(n35948) );
  NAND2_X2 U23102 ( .A1(n7861), .A2(n36262), .ZN(n32607) );
  NAND2_X1 U1985 ( .A1(n18402), .A2(n24383), .ZN(n35985) );
  INV_X2 U30527 ( .I(n33895), .ZN(n20423) );
  NAND2_X2 U10822 ( .A1(n15424), .A2(n29776), .ZN(n5923) );
  NAND2_X1 U20997 ( .A1(n18534), .A2(n33726), .ZN(n32215) );
  NAND2_X2 U21785 ( .A1(n28475), .A2(n31088), .ZN(n9673) );
  NOR2_X1 U24674 ( .A1(n4800), .A2(n36188), .ZN(n13480) );
  INV_X2 U15371 ( .I(n34987), .ZN(n20407) );
  NOR3_X1 U13393 ( .A1(n18506), .A2(n17578), .A3(n18462), .ZN(n18505) );
  NAND3_X2 U17057 ( .A1(n26645), .A2(n26751), .A3(n26754), .ZN(n26352) );
  NAND3_X2 U232 ( .A1(n31347), .A2(n2469), .A3(n1195), .ZN(n6370) );
  INV_X1 U816 ( .I(n25481), .ZN(n1534) );
  NOR2_X2 U28387 ( .A1(n1152), .A2(n22092), .ZN(n22091) );
  INV_X2 U9110 ( .I(n10255), .ZN(n19750) );
  OAI21_X2 U6598 ( .A1(n22093), .A2(n22094), .B(n35060), .ZN(n22095) );
  NAND3_X1 U10599 ( .A1(n16126), .A2(n31662), .A3(n31661), .ZN(n34416) );
  NAND2_X2 U3320 ( .A1(n8131), .A2(n28807), .ZN(n2469) );
  INV_X4 U8333 ( .I(n24266), .ZN(n1601) );
  NOR2_X2 U13275 ( .A1(n7939), .A2(n38119), .ZN(n7938) );
  NAND2_X2 U29242 ( .A1(n34892), .A2(n1089), .ZN(n26422) );
  AOI21_X2 U2637 ( .A1(n36912), .A2(n6604), .B(n5392), .ZN(n35699) );
  NAND2_X1 U17385 ( .A1(n15719), .A2(n36649), .ZN(n4745) );
  NAND2_X2 U7417 ( .A1(n11574), .A2(n1177), .ZN(n10408) );
  AND2_X1 U3936 ( .A1(n14450), .A2(n19313), .Z(n32410) );
  NAND2_X1 U11545 ( .A1(n16919), .A2(n1000), .ZN(n27024) );
  INV_X1 U21539 ( .I(n32310), .ZN(n33450) );
  NOR2_X1 U10216 ( .A1(n3435), .A2(n1687), .ZN(n4902) );
  INV_X4 U7858 ( .I(n27306), .ZN(n1086) );
  NOR2_X1 U8078 ( .A1(n5664), .A2(n33662), .ZN(n33908) );
  INV_X2 U12076 ( .I(n26021), .ZN(n10474) );
  NAND2_X2 U13773 ( .A1(n31940), .A2(n35754), .ZN(n22212) );
  AOI22_X2 U1427 ( .A1(n2246), .A2(n36083), .B1(n2247), .B2(n517), .ZN(n35371)
         );
  INV_X2 U605 ( .I(n26974), .ZN(n1497) );
  INV_X4 U7329 ( .I(n1746), .ZN(n2840) );
  BUF_X2 U6912 ( .I(n25106), .Z(n25448) );
  NAND2_X1 U10096 ( .A1(n35440), .A2(n4647), .ZN(n36053) );
  NAND2_X2 U10003 ( .A1(n22886), .A2(n20638), .ZN(n18365) );
  AOI21_X2 U7896 ( .A1(n1231), .A2(n35537), .B(n8651), .ZN(n12694) );
  INV_X2 U12282 ( .I(n11332), .ZN(n11331) );
  NAND2_X2 U329 ( .A1(n36414), .A2(n36671), .ZN(n35478) );
  NAND2_X1 U20217 ( .A1(n32063), .A2(n32062), .ZN(n24624) );
  NAND2_X2 U4288 ( .A1(n13542), .A2(n935), .ZN(n465) );
  BUF_X4 U29360 ( .I(n31132), .Z(n36673) );
  INV_X1 U130 ( .I(n19783), .ZN(n30232) );
  BUF_X4 U2751 ( .I(n36791), .Z(n209) );
  INV_X2 U28975 ( .I(n25469), .ZN(n25609) );
  NOR2_X1 U16916 ( .A1(n5682), .A2(n4677), .ZN(n5679) );
  INV_X4 U13025 ( .I(n19990), .ZN(n21310) );
  NOR2_X1 U770 ( .A1(n34660), .A2(n37241), .ZN(n35768) );
  NOR2_X2 U2335 ( .A1(n33737), .A2(n36506), .ZN(n35361) );
  AOI22_X2 U954 ( .A1(n26994), .A2(n1229), .B1(n26996), .B2(n19364), .ZN(
        n34257) );
  OAI21_X1 U15884 ( .A1(n7418), .A2(n27180), .B(n31459), .ZN(n27004) );
  AOI21_X2 U7415 ( .A1(n29420), .A2(n505), .B(n12262), .ZN(n12261) );
  NOR3_X2 U95 ( .A1(n505), .A2(n9993), .A3(n29494), .ZN(n12262) );
  BUF_X2 U3064 ( .I(n18866), .Z(n9190) );
  NOR2_X1 U19330 ( .A1(n18628), .A2(n1073), .ZN(n36060) );
  INV_X2 U1114 ( .I(n39055), .ZN(n13446) );
  INV_X2 U11169 ( .I(n24661), .ZN(n1028) );
  OAI21_X2 U6885 ( .A1(n16779), .A2(n9922), .B(n7949), .ZN(n32250) );
  NOR2_X2 U13344 ( .A1(n11583), .A2(n4963), .ZN(n12254) );
  NAND2_X2 U10343 ( .A1(n21413), .A2(n19543), .ZN(n11433) );
  BUF_X4 U8037 ( .I(n20406), .Z(n1755) );
  NOR2_X2 U24051 ( .A1(n19488), .A2(n1763), .ZN(n23091) );
  INV_X1 U10593 ( .I(n12369), .ZN(n7302) );
  OAI21_X2 U2979 ( .A1(n35830), .A2(n12543), .B(n34702), .ZN(n18259) );
  BUF_X4 U8776 ( .I(Key[102]), .Z(n30170) );
  NAND2_X1 U24360 ( .A1(n372), .A2(n20921), .ZN(n32884) );
  NAND2_X2 U5368 ( .A1(n35330), .A2(n35329), .ZN(n139) );
  NOR2_X2 U18416 ( .A1(n31994), .A2(n34265), .ZN(n25981) );
  NAND3_X1 U6379 ( .A1(n17998), .A2(n1049), .A3(n21117), .ZN(n10744) );
  BUF_X4 U5974 ( .I(n24276), .Z(n14378) );
  INV_X2 U14792 ( .I(n26019), .ZN(n31310) );
  AOI21_X2 U22277 ( .A1(n38673), .A2(n10154), .B(n22114), .ZN(n11439) );
  NAND2_X2 U5355 ( .A1(n33855), .A2(n9799), .ZN(n34688) );
  AND2_X2 U3274 ( .A1(n15461), .A2(n7240), .Z(n24472) );
  NAND2_X2 U7615 ( .A1(n28069), .A2(n5020), .ZN(n10826) );
  OAI21_X2 U7016 ( .A1(n24314), .A2(n33077), .B(n5572), .ZN(n1877) );
  INV_X2 U1115 ( .I(n16590), .ZN(n20791) );
  NOR2_X1 U20266 ( .A1(n28270), .A2(n1198), .ZN(n12497) );
  NOR2_X1 U21317 ( .A1(n34063), .A2(n35629), .ZN(n36853) );
  INV_X4 U18431 ( .I(n5558), .ZN(n5935) );
  INV_X4 U17458 ( .I(n11092), .ZN(n20924) );
  INV_X1 U1095 ( .I(n18790), .ZN(n24372) );
  NAND3_X2 U9707 ( .A1(n17592), .A2(n24242), .A3(n1593), .ZN(n17591) );
  NAND2_X1 U6770 ( .A1(n30507), .A2(n16079), .ZN(n16078) );
  OAI21_X2 U3112 ( .A1(n17900), .A2(n30851), .B(n30556), .ZN(n16953) );
  INV_X4 U9591 ( .I(n24925), .ZN(n1259) );
  OAI21_X2 U20051 ( .A1(n16841), .A2(n37355), .B(n17350), .ZN(n24509) );
  NOR2_X1 U5516 ( .A1(n7840), .A2(n7839), .ZN(n35523) );
  BUF_X2 U26685 ( .I(n10054), .Z(n33151) );
  NOR2_X1 U6820 ( .A1(n4821), .A2(n24395), .ZN(n12803) );
  OAI22_X2 U18877 ( .A1(n36244), .A2(n7978), .B1(n26702), .B2(n30795), .ZN(
        n26707) );
  NAND2_X2 U2072 ( .A1(n2192), .A2(n36500), .ZN(n4183) );
  INV_X4 U22999 ( .I(n3644), .ZN(n22114) );
  INV_X2 U4408 ( .I(n18722), .ZN(n21478) );
  INV_X2 U1107 ( .I(n13584), .ZN(n10747) );
  NAND2_X2 U23700 ( .A1(n17294), .A2(n17296), .ZN(n32714) );
  AOI21_X2 U25012 ( .A1(n29481), .A2(n29454), .B(n29426), .ZN(n17296) );
  BUF_X2 U5125 ( .I(n8646), .Z(n33412) );
  AOI21_X1 U20574 ( .A1(n3067), .A2(n3066), .B(n3065), .ZN(n32132) );
  NAND2_X2 U12665 ( .A1(n12517), .A2(n37421), .ZN(n9826) );
  NAND2_X1 U13734 ( .A1(n28507), .A2(n34794), .ZN(n34781) );
  NAND2_X1 U12873 ( .A1(n12803), .A2(n24397), .ZN(n12802) );
  OAI21_X2 U23107 ( .A1(n28342), .A2(n28401), .B(n28341), .ZN(n11665) );
  NAND2_X1 U4651 ( .A1(n18384), .A2(n29531), .ZN(n17103) );
  INV_X4 U13533 ( .I(n6885), .ZN(n17286) );
  INV_X2 U9129 ( .I(n31494), .ZN(n1204) );
  BUF_X4 U3879 ( .I(n3213), .Z(n362) );
  OAI21_X2 U12858 ( .A1(n7730), .A2(n19745), .B(n13707), .ZN(n13706) );
  NAND2_X2 U6352 ( .A1(n5907), .A2(n20638), .ZN(n20637) );
  NAND2_X1 U5784 ( .A1(n32266), .A2(n31359), .ZN(n35440) );
  OAI21_X1 U28397 ( .A1(n25469), .A2(n32556), .B(n19968), .ZN(n32266) );
  OAI21_X2 U13453 ( .A1(n22512), .A2(n23213), .B(n1312), .ZN(n2253) );
  OAI21_X2 U2102 ( .A1(n8682), .A2(n8681), .B(n24448), .ZN(n11631) );
  INV_X1 U13149 ( .I(n26497), .ZN(n34712) );
  AOI22_X2 U2790 ( .A1(n29482), .A2(n19896), .B1(n29378), .B2(n31521), .ZN(
        n6734) );
  INV_X1 U7994 ( .I(n27969), .ZN(n28233) );
  NOR2_X2 U4692 ( .A1(n5392), .A2(n37351), .ZN(n5451) );
  OAI21_X2 U24613 ( .A1(n7284), .A2(n1255), .B(n1256), .ZN(n16411) );
  BUF_X2 U7412 ( .I(n11083), .Z(n34360) );
  OAI22_X2 U4694 ( .A1(n27207), .A2(n27325), .B1(n27326), .B2(n1473), .ZN(n556) );
  INV_X4 U5415 ( .I(n19499), .ZN(n6337) );
  NAND2_X2 U5352 ( .A1(n30746), .A2(n30745), .ZN(n36947) );
  CLKBUF_X4 U5523 ( .I(n28174), .Z(n3989) );
  CLKBUF_X4 U20441 ( .I(n24195), .Z(n6515) );
  NAND3_X2 U21584 ( .A1(n24710), .A2(n6491), .A3(n33986), .ZN(n9364) );
  BUF_X2 U5637 ( .I(n13770), .Z(n36424) );
  OR2_X2 U14370 ( .A1(n32986), .A2(n31254), .Z(n18575) );
  NAND3_X1 U1 ( .A1(n32452), .A2(n18795), .A3(n20862), .ZN(n36919) );
  INV_X2 U9583 ( .I(n19572), .ZN(n19941) );
  NOR3_X2 U4603 ( .A1(n11271), .A2(n11081), .A3(n9218), .ZN(n9474) );
  NAND2_X2 U11324 ( .A1(n8351), .A2(n11407), .ZN(n8350) );
  BUF_X2 U2576 ( .I(n28157), .Z(n28269) );
  NAND2_X2 U17629 ( .A1(n13593), .A2(n18187), .ZN(n19305) );
  INV_X1 U25549 ( .I(n19631), .ZN(n976) );
  INV_X2 U7159 ( .I(n962), .ZN(n1313) );
  AOI22_X2 U8105 ( .A1(n2799), .A2(n954), .B1(n728), .B2(n21254), .ZN(n4132)
         );
  INV_X2 U7176 ( .I(n23162), .ZN(n22996) );
  BUF_X4 U4910 ( .I(n17650), .Z(n9776) );
  OAI22_X2 U1924 ( .A1(n15828), .A2(n24433), .B1(n1608), .B2(n30897), .ZN(
        n15826) );
  INV_X2 U29080 ( .I(n36263), .ZN(n36630) );
  NAND2_X2 U9286 ( .A1(n26996), .A2(n17655), .ZN(n20562) );
  NOR3_X2 U2974 ( .A1(n19412), .A2(n19411), .A3(n29656), .ZN(n18243) );
  INV_X4 U1900 ( .I(n3708), .ZN(n23521) );
  BUF_X2 U7092 ( .I(n25798), .Z(n34961) );
  INV_X1 U612 ( .I(n875), .ZN(n11337) );
  INV_X2 U6652 ( .I(n19823), .ZN(n23070) );
  OAI21_X2 U4129 ( .A1(n13111), .A2(n19364), .B(n26692), .ZN(n17826) );
  NAND2_X2 U2241 ( .A1(n23413), .A2(n5591), .ZN(n34635) );
  BUF_X2 U9127 ( .I(n27481), .Z(n28123) );
  BUF_X2 U5330 ( .I(n24369), .Z(n19942) );
  INV_X2 U1175 ( .I(n25820), .ZN(n1511) );
  NOR2_X1 U11215 ( .A1(n3055), .A2(n3056), .ZN(n36709) );
  INV_X1 U1053 ( .I(n24296), .ZN(n1598) );
  NAND2_X2 U2034 ( .A1(n20783), .A2(n1142), .ZN(n15272) );
  NAND2_X1 U5245 ( .A1(n15940), .A2(n17470), .ZN(n21128) );
  INV_X4 U4974 ( .I(n22132), .ZN(n22030) );
  INV_X4 U21390 ( .I(n11653), .ZN(n19544) );
  BUF_X2 U3088 ( .I(n12673), .Z(n30995) );
  BUF_X2 U7265 ( .I(n26665), .Z(n12290) );
  CLKBUF_X2 U8761 ( .I(Key[139]), .Z(n19839) );
  NOR2_X2 U20443 ( .A1(n12705), .A2(n38685), .ZN(n12702) );
  NAND2_X2 U29406 ( .A1(n22302), .A2(n22303), .ZN(n22305) );
  AOI21_X2 U7335 ( .A1(n26980), .A2(n26687), .B(n12290), .ZN(n12590) );
  NOR2_X2 U8224 ( .A1(n2697), .A2(n1996), .ZN(n1995) );
  AOI21_X2 U12115 ( .A1(n13168), .A2(n9605), .B(n32109), .ZN(n11764) );
  OAI21_X2 U14296 ( .A1(n27956), .A2(n16325), .B(n34832), .ZN(n11208) );
  NAND2_X1 U1234 ( .A1(n31432), .A2(n17952), .ZN(n35353) );
  NAND2_X2 U13138 ( .A1(n3383), .A2(n23117), .ZN(n3382) );
  BUF_X2 U16707 ( .I(n19467), .Z(n28048) );
  NAND2_X1 U25124 ( .A1(n23271), .A2(n23355), .ZN(n18197) );
  BUF_X4 U2065 ( .I(n7536), .Z(n123) );
  NAND2_X1 U26094 ( .A1(n28479), .A2(n1419), .ZN(n21190) );
  AOI21_X1 U11778 ( .A1(n21171), .A2(n26219), .B(n16298), .ZN(n5560) );
  OAI21_X1 U11596 ( .A1(n20709), .A2(n7499), .B(n20708), .ZN(n8208) );
  NOR2_X2 U7905 ( .A1(n21099), .A2(n26970), .ZN(n3541) );
  NAND2_X2 U8936 ( .A1(n1416), .A2(n2022), .ZN(n8849) );
  INV_X4 U6984 ( .I(n9276), .ZN(n10116) );
  INV_X2 U5027 ( .I(n22711), .ZN(n1322) );
  BUF_X4 U1393 ( .I(n25718), .Z(n19400) );
  NOR2_X2 U18172 ( .A1(n38609), .A2(n31697), .ZN(n13) );
  BUF_X4 U6688 ( .I(n18229), .Z(n12392) );
  INV_X2 U7731 ( .I(n1445), .ZN(n1207) );
  NAND2_X1 U25190 ( .A1(n33109), .A2(n14839), .ZN(n12105) );
  OAI22_X1 U17941 ( .A1(n23309), .A2(n39626), .B1(n23607), .B2(n23311), .ZN(
        n5592) );
  AOI22_X2 U9789 ( .A1(n863), .A2(n1093), .B1(n36477), .B2(n34163), .ZN(n34335) );
  INV_X2 U4442 ( .I(n19465), .ZN(n10902) );
  BUF_X4 U2137 ( .I(n27249), .Z(n7676) );
  NAND2_X1 U28428 ( .A1(n33370), .A2(n33369), .ZN(n7806) );
  NOR2_X2 U17638 ( .A1(n38914), .A2(n25849), .ZN(n2424) );
  NAND3_X1 U4949 ( .A1(n4750), .A2(n7367), .A3(n21808), .ZN(n7999) );
  NOR2_X2 U12040 ( .A1(n11858), .A2(n26068), .ZN(n2541) );
  BUF_X2 U25423 ( .I(n22674), .Z(n18072) );
  BUF_X2 U8009 ( .I(n3158), .Z(n3032) );
  CLKBUF_X4 U2959 ( .I(n13545), .Z(n611) );
  CLKBUF_X2 U10467 ( .I(Key[80]), .Z(n29282) );
  BUF_X2 U4333 ( .I(n20591), .Z(n20173) );
  INV_X1 U8395 ( .I(n10174), .ZN(n1626) );
  NAND2_X1 U12653 ( .A1(n34646), .A2(n34645), .ZN(n25972) );
  NAND3_X1 U13547 ( .A1(n10146), .A2(n10147), .A3(n971), .ZN(n34763) );
  INV_X4 U5793 ( .I(n7357), .ZN(n18429) );
  NAND2_X2 U315 ( .A1(n7325), .A2(n8056), .ZN(n7946) );
  NOR2_X1 U6658 ( .A1(n10353), .A2(n36090), .ZN(n10354) );
  INV_X4 U19807 ( .I(n28560), .ZN(n28654) );
  OAI21_X2 U5780 ( .A1(n22301), .A2(n22075), .B(n22076), .ZN(n20356) );
  NAND2_X1 U4449 ( .A1(n24917), .A2(n18876), .ZN(n33209) );
  NAND2_X1 U12201 ( .A1(n17037), .A2(n39821), .ZN(n36693) );
  NAND3_X1 U2539 ( .A1(n13723), .A2(n13441), .A3(n18997), .ZN(n2555) );
  NOR2_X1 U5363 ( .A1(n29425), .A2(n20830), .ZN(n35296) );
  OR2_X1 U10323 ( .A1(n34483), .A2(n34597), .Z(n34613) );
  INV_X2 U1105 ( .I(n12235), .ZN(n24118) );
  NAND2_X1 U14436 ( .A1(n34855), .A2(n31430), .ZN(n18554) );
  AOI21_X1 U312 ( .A1(n36742), .A2(n35804), .B(n32800), .ZN(n6371) );
  INV_X4 U10105 ( .I(n37589), .ZN(n23213) );
  NOR2_X2 U6924 ( .A1(n9703), .A2(n24853), .ZN(n14934) );
  OAI22_X2 U22350 ( .A1(n10116), .A2(n17087), .B1(n9277), .B2(n32064), .ZN(
        n9703) );
  NAND2_X1 U5629 ( .A1(n5070), .A2(n33708), .ZN(n14201) );
  NAND3_X1 U11229 ( .A1(n27986), .A2(n38874), .A3(n20053), .ZN(n27987) );
  AOI21_X2 U5496 ( .A1(n13826), .A2(n11806), .B(n1117), .ZN(n32365) );
  NAND2_X1 U18278 ( .A1(n18346), .A2(n13653), .ZN(n9280) );
  INV_X2 U4568 ( .I(n9861), .ZN(n31139) );
  NOR2_X1 U13757 ( .A1(n14777), .A2(n22245), .ZN(n20731) );
  NOR2_X2 U3473 ( .A1(n24698), .A2(n37097), .ZN(n1909) );
  NAND2_X1 U11832 ( .A1(n31238), .A2(n31237), .ZN(n31236) );
  INV_X2 U5969 ( .I(n24408), .ZN(n24406) );
  INV_X2 U30367 ( .I(n14234), .ZN(n23115) );
  INV_X2 U12136 ( .I(n25889), .ZN(n7293) );
  NAND2_X2 U12184 ( .A1(n26079), .A2(n1012), .ZN(n18876) );
  BUF_X4 U30742 ( .I(n5831), .Z(n36989) );
  NAND2_X1 U21912 ( .A1(n30393), .A2(n21533), .ZN(n16930) );
  NAND3_X2 U7792 ( .A1(n27072), .A2(n34943), .A3(n39338), .ZN(n5294) );
  INV_X2 U23072 ( .I(n12141), .ZN(n14933) );
  INV_X2 U1045 ( .I(n20936), .ZN(n35764) );
  BUF_X4 U3434 ( .I(n29897), .Z(n30059) );
  INV_X2 U27300 ( .I(n33244), .ZN(n33935) );
  INV_X1 U5591 ( .I(n16520), .ZN(n27310) );
  AOI21_X1 U4781 ( .A1(n3637), .A2(n12527), .B(n33647), .ZN(n31036) );
  INV_X2 U9968 ( .I(n6355), .ZN(n27412) );
  AOI21_X2 U7402 ( .A1(n29378), .A2(n31521), .B(n16877), .ZN(n16876) );
  INV_X1 U21016 ( .I(n23202), .ZN(n35576) );
  INV_X2 U17427 ( .I(n13414), .ZN(n1036) );
  NAND2_X1 U11732 ( .A1(n11222), .A2(n11220), .ZN(n11225) );
  INV_X2 U1424 ( .I(n20351), .ZN(n1329) );
  NAND2_X2 U8178 ( .A1(n32223), .A2(n32221), .ZN(n24365) );
  NAND2_X2 U13405 ( .A1(n3683), .A2(n22902), .ZN(n14331) );
  BUF_X4 U5278 ( .I(n35614), .Z(n34014) );
  OR2_X2 U4671 ( .A1(n24483), .A2(n32360), .Z(n30373) );
  NAND2_X1 U24465 ( .A1(n25708), .A2(n33218), .ZN(n18215) );
  NAND2_X2 U1579 ( .A1(n39258), .A2(n1909), .ZN(n3399) );
  NAND3_X2 U7845 ( .A1(n4583), .A2(n946), .A3(n4582), .ZN(n4581) );
  AOI21_X2 U8368 ( .A1(n20036), .A2(n23559), .B(n23560), .ZN(n20035) );
  NAND2_X2 U3546 ( .A1(n23430), .A2(n34494), .ZN(n20036) );
  NOR2_X2 U3524 ( .A1(n26980), .A2(n26687), .ZN(n14830) );
  INV_X2 U9322 ( .I(n26655), .ZN(n13645) );
  OAI22_X2 U200 ( .A1(n9692), .A2(n7063), .B1(n18035), .B2(n39724), .ZN(n14091) );
  OR2_X2 U21510 ( .A1(n35748), .A2(n25606), .Z(n25608) );
  NAND2_X2 U1285 ( .A1(n7941), .A2(n31523), .ZN(n35499) );
  OAI21_X1 U12537 ( .A1(n2704), .A2(n2703), .B(n33195), .ZN(n2701) );
  BUF_X2 U30108 ( .I(n15922), .Z(n33603) );
  INV_X1 U4782 ( .I(n12527), .ZN(n1430) );
  NAND2_X2 U909 ( .A1(n34538), .A2(n37585), .ZN(n9535) );
  INV_X4 U21060 ( .I(n8526), .ZN(n19728) );
  NOR2_X1 U5801 ( .A1(n9926), .A2(n27187), .ZN(n27192) );
  BUF_X4 U5949 ( .I(n28660), .Z(n33436) );
  NAND3_X2 U1174 ( .A1(n8860), .A2(n8858), .A3(n34482), .ZN(n34481) );
  NOR2_X2 U10226 ( .A1(n34085), .A2(n25435), .ZN(n11442) );
  INV_X4 U6978 ( .I(n19507), .ZN(n20696) );
  NOR2_X1 U2040 ( .A1(n8979), .A2(n8978), .ZN(n8977) );
  NAND2_X2 U657 ( .A1(n2518), .A2(n576), .ZN(n35218) );
  OAI21_X1 U8287 ( .A1(n12975), .A2(n24433), .B(n10023), .ZN(n13072) );
  INV_X2 U7495 ( .I(n6317), .ZN(n5542) );
  INV_X4 U3998 ( .I(n28669), .ZN(n14209) );
  NAND2_X2 U10148 ( .A1(n36008), .A2(n36007), .ZN(n25845) );
  AOI21_X2 U12251 ( .A1(n11268), .A2(n953), .B(n11944), .ZN(n16737) );
  OAI21_X2 U1524 ( .A1(n2288), .A2(n33480), .B(n30941), .ZN(n171) );
  INV_X4 U26698 ( .I(n18077), .ZN(n25468) );
  NAND2_X2 U9815 ( .A1(n33804), .A2(n33805), .ZN(n34342) );
  NOR3_X2 U26201 ( .A1(n17346), .A2(n26564), .A3(n17194), .ZN(n15879) );
  NOR2_X1 U10247 ( .A1(n6822), .A2(n24527), .ZN(n15168) );
  NAND3_X1 U21967 ( .A1(n32485), .A2(n21224), .A3(n36844), .ZN(n32411) );
  INV_X2 U27278 ( .I(n33242), .ZN(n728) );
  OAI21_X1 U1056 ( .A1(n33539), .A2(n1239), .B(n7415), .ZN(n20802) );
  INV_X1 U26367 ( .I(n26643), .ZN(n36306) );
  NOR2_X2 U1679 ( .A1(n33532), .A2(n33530), .ZN(n33529) );
  INV_X1 U12423 ( .I(n25483), .ZN(n6248) );
  OAI21_X1 U11821 ( .A1(n14427), .A2(n21091), .B(n18469), .ZN(n17144) );
  AOI21_X2 U24050 ( .A1(n23169), .A2(n1763), .B(n22810), .ZN(n22811) );
  OAI21_X1 U7008 ( .A1(n25614), .A2(n25613), .B(n25612), .ZN(n25618) );
  NAND2_X1 U11560 ( .A1(n26622), .A2(n1500), .ZN(n34538) );
  NOR2_X2 U6073 ( .A1(n21236), .A2(n9048), .ZN(n9047) );
  OR2_X2 U24577 ( .A1(n6163), .A2(n7140), .Z(n7141) );
  NAND4_X2 U8953 ( .A1(n29847), .A2(n5108), .A3(n5107), .A4(n34267), .ZN(
        n34552) );
  INV_X4 U1355 ( .I(n9854), .ZN(n23160) );
  INV_X2 U2468 ( .I(n12393), .ZN(n34789) );
  INV_X4 U14922 ( .I(n35883), .ZN(n34923) );
  INV_X2 U4815 ( .I(n20321), .ZN(n26841) );
  NAND2_X1 U13190 ( .A1(n23249), .A2(n6637), .ZN(n11528) );
  CLKBUF_X2 U2008 ( .I(n22993), .Z(n32084) );
  BUF_X2 U10473 ( .I(Key[11]), .Z(n29849) );
  BUF_X2 U4871 ( .I(n34122), .Z(n33899) );
  INV_X2 U14314 ( .I(n9266), .ZN(n17447) );
  BUF_X2 U6468 ( .I(Key[49]), .Z(n17428) );
  BUF_X2 U10482 ( .I(Key[21]), .Z(n19755) );
  BUF_X2 U14049 ( .I(Key[148]), .Z(n19534) );
  BUF_X2 U10445 ( .I(Key[12]), .Z(n19722) );
  BUF_X2 U7313 ( .I(Key[126]), .Z(n19815) );
  BUF_X2 U14053 ( .I(Key[86]), .Z(n19879) );
  CLKBUF_X2 U10448 ( .I(Key[155]), .Z(n30122) );
  INV_X1 U28501 ( .I(Key[3]), .ZN(n29528) );
  BUF_X2 U8760 ( .I(Key[22]), .Z(n19730) );
  BUF_X2 U6466 ( .I(Key[187]), .Z(n19761) );
  INV_X1 U20774 ( .I(n29887), .ZN(n32174) );
  CLKBUF_X4 U10437 ( .I(n21790), .Z(n18205) );
  INV_X1 U8863 ( .I(n28821), .ZN(n30682) );
  INV_X2 U10411 ( .I(n8936), .ZN(n21833) );
  INV_X1 U25516 ( .I(n19763), .ZN(n14820) );
  INV_X1 U26977 ( .I(n29463), .ZN(n33184) );
  INV_X2 U8722 ( .I(n34122), .ZN(n21923) );
  CLKBUF_X2 U30573 ( .I(n32370), .Z(n36887) );
  INV_X1 U27790 ( .I(n30016), .ZN(n33311) );
  CLKBUF_X4 U7296 ( .I(n11576), .Z(n10120) );
  CLKBUF_X2 U14006 ( .I(n21752), .Z(n19416) );
  BUF_X2 U4969 ( .I(n21496), .Z(n16128) );
  INV_X1 U14007 ( .I(n29141), .ZN(n18700) );
  CLKBUF_X2 U26650 ( .I(n695), .Z(n33148) );
  INV_X2 U1518 ( .I(n17209), .ZN(n21894) );
  CLKBUF_X2 U4879 ( .I(n12670), .Z(n33885) );
  CLKBUF_X2 U14002 ( .I(n21841), .Z(n18152) );
  INV_X1 U25500 ( .I(n29337), .ZN(n20479) );
  CLKBUF_X2 U6436 ( .I(n20810), .Z(n10044) );
  INV_X2 U8662 ( .I(n34247), .ZN(n20923) );
  INV_X2 U23225 ( .I(n21761), .ZN(n11851) );
  INV_X2 U7866 ( .I(n17799), .ZN(n18028) );
  CLKBUF_X2 U27618 ( .I(n21840), .Z(n33285) );
  INV_X1 U27516 ( .I(n21789), .ZN(n21527) );
  OR2_X1 U23244 ( .A1(n11900), .A2(n18293), .Z(n15274) );
  NAND2_X1 U22005 ( .A1(n21728), .A2(n36721), .ZN(n35723) );
  NAND2_X1 U17056 ( .A1(n21867), .A2(n15359), .ZN(n12333) );
  AOI21_X1 U13825 ( .A1(n21059), .A2(n21058), .B(n7640), .ZN(n21057) );
  OAI21_X1 U20143 ( .A1(n17866), .A2(n21859), .B(n36351), .ZN(n35437) );
  BUF_X2 U7728 ( .I(n8040), .Z(n3676) );
  CLKBUF_X4 U3304 ( .I(n22354), .Z(n9685) );
  NAND2_X1 U16900 ( .A1(n4424), .A2(n20679), .ZN(n5796) );
  CLKBUF_X2 U21260 ( .I(n22122), .Z(n32259) );
  BUF_X2 U4045 ( .I(n2696), .Z(n32434) );
  CLKBUF_X4 U5791 ( .I(n11327), .Z(n11171) );
  INV_X2 U15527 ( .I(n22292), .ZN(n33713) );
  CLKBUF_X2 U27270 ( .I(n8882), .Z(n36457) );
  BUF_X2 U30132 ( .I(n19773), .Z(n33623) );
  INV_X2 U1426 ( .I(n22281), .ZN(n19486) );
  CLKBUF_X4 U25788 ( .I(n19655), .Z(n36237) );
  AOI21_X1 U6495 ( .A1(n1686), .A2(n13191), .B(n38375), .ZN(n11234) );
  INV_X1 U6021 ( .I(n22045), .ZN(n10924) );
  INV_X1 U17744 ( .I(n12964), .ZN(n20773) );
  NOR2_X1 U10144 ( .A1(n22199), .A2(n8518), .ZN(n14270) );
  CLKBUF_X4 U14112 ( .I(n1326), .Z(n34808) );
  NAND2_X1 U28422 ( .A1(n22353), .A2(n21288), .ZN(n22208) );
  NAND2_X1 U17545 ( .A1(n22009), .A2(n22214), .ZN(n21105) );
  OAI21_X1 U28413 ( .A1(n22204), .A2(n19837), .B(n22207), .ZN(n22163) );
  CLKBUF_X4 U2531 ( .I(n22334), .Z(n36443) );
  OAI21_X1 U24186 ( .A1(n15294), .A2(n13910), .B(n22156), .ZN(n13909) );
  NAND2_X1 U20007 ( .A1(n12433), .A2(n7093), .ZN(n36436) );
  NOR2_X1 U6564 ( .A1(n8701), .A2(n22172), .ZN(n33228) );
  NAND2_X1 U27606 ( .A1(n22144), .A2(n33438), .ZN(n19430) );
  INV_X1 U27748 ( .I(n21298), .ZN(n20239) );
  AOI21_X1 U25088 ( .A1(n21337), .A2(n14024), .B(n33359), .ZN(n19216) );
  NAND2_X1 U2208 ( .A1(n21335), .A2(n21334), .ZN(n21338) );
  NAND2_X1 U13690 ( .A1(n11142), .A2(n1149), .ZN(n11141) );
  INV_X1 U4162 ( .I(n34345), .ZN(n36778) );
  CLKBUF_X4 U2938 ( .I(n6014), .Z(n5284) );
  INV_X1 U24425 ( .I(n16798), .ZN(n22174) );
  NAND2_X1 U20955 ( .A1(n22026), .A2(n22027), .ZN(n4630) );
  BUF_X2 U8053 ( .I(n3528), .Z(n34188) );
  CLKBUF_X2 U6266 ( .I(n33227), .Z(n36362) );
  BUF_X1 U13602 ( .I(n22773), .Z(n19848) );
  NAND2_X1 U15263 ( .A1(n33072), .A2(n33780), .ZN(n34972) );
  CLKBUF_X2 U20866 ( .I(n15346), .Z(n35559) );
  INV_X2 U25494 ( .I(n22430), .ZN(n21215) );
  INV_X1 U6258 ( .I(n7560), .ZN(n34691) );
  CLKBUF_X2 U11465 ( .I(n22711), .Z(n30950) );
  CLKBUF_X2 U6239 ( .I(n23140), .Z(n36763) );
  CLKBUF_X2 U23928 ( .I(n5337), .Z(n35994) );
  CLKBUF_X4 U10088 ( .I(n23152), .Z(n8569) );
  CLKBUF_X1 U4008 ( .I(n12631), .Z(n31183) );
  CLKBUF_X2 U6231 ( .I(n13668), .Z(n34419) );
  BUF_X2 U2006 ( .I(n22709), .Z(n383) );
  INV_X2 U2462 ( .I(n8539), .ZN(n33925) );
  CLKBUF_X2 U2458 ( .I(n407), .Z(n32515) );
  BUF_X2 U6224 ( .I(n23164), .Z(n36095) );
  CLKBUF_X4 U6235 ( .I(n22946), .Z(n34013) );
  CLKBUF_X4 U13568 ( .I(n23102), .Z(n18244) );
  INV_X2 U8550 ( .I(n14442), .ZN(n1147) );
  INV_X2 U1368 ( .I(n7160), .ZN(n16678) );
  BUF_X2 U6655 ( .I(n21291), .Z(n11582) );
  BUF_X2 U4784 ( .I(n39811), .Z(n33082) );
  INV_X1 U6617 ( .I(n12029), .ZN(n35667) );
  INV_X1 U23236 ( .I(n32636), .ZN(n23052) );
  INV_X1 U1359 ( .I(n22864), .ZN(n22994) );
  NAND2_X1 U13469 ( .A1(n9255), .A2(n23123), .ZN(n3046) );
  INV_X1 U6226 ( .I(n11913), .ZN(n35851) );
  INV_X2 U2432 ( .I(n23020), .ZN(n23138) );
  INV_X2 U14767 ( .I(n22833), .ZN(n1141) );
  NAND2_X1 U10563 ( .A1(n32084), .A2(n15239), .ZN(n15238) );
  INV_X2 U1326 ( .I(n781), .ZN(n1045) );
  NOR2_X1 U8481 ( .A1(n17124), .A2(n35442), .ZN(n5810) );
  NAND2_X1 U25339 ( .A1(n23177), .A2(n23174), .ZN(n36185) );
  OR2_X1 U4031 ( .A1(n23066), .A2(n22994), .Z(n14747) );
  NAND2_X1 U27440 ( .A1(n19013), .A2(n14390), .ZN(n22918) );
  NOR2_X1 U5264 ( .A1(n33763), .A2(n19697), .ZN(n36043) );
  NOR2_X1 U2349 ( .A1(n14879), .A2(n30394), .ZN(n35347) );
  NAND2_X1 U19635 ( .A1(n22997), .A2(n35586), .ZN(n9330) );
  NAND2_X1 U6192 ( .A1(n3811), .A2(n10828), .ZN(n36094) );
  INV_X1 U19030 ( .I(n13719), .ZN(n23184) );
  INV_X1 U19691 ( .I(n19528), .ZN(n7010) );
  NAND2_X1 U6182 ( .A1(n36043), .A2(n18386), .ZN(n35092) );
  OAI21_X1 U23540 ( .A1(n23020), .A2(n36763), .B(n35939), .ZN(n4690) );
  NAND2_X1 U22717 ( .A1(n22280), .A2(n22833), .ZN(n32552) );
  OAI21_X1 U28599 ( .A1(n23063), .A2(n23062), .B(n23061), .ZN(n23064) );
  OAI21_X1 U3226 ( .A1(n37062), .A2(n22999), .B(n23000), .ZN(n8058) );
  CLKBUF_X4 U3391 ( .I(n38704), .Z(n5591) );
  BUF_X2 U13332 ( .I(n23464), .Z(n5083) );
  INV_X1 U13475 ( .I(n17968), .ZN(n23185) );
  CLKBUF_X4 U5231 ( .I(n33453), .Z(n31685) );
  CLKBUF_X2 U2302 ( .I(n12028), .Z(n35525) );
  CLKBUF_X4 U7100 ( .I(n11669), .Z(n6637) );
  INV_X2 U14384 ( .I(n4644), .ZN(n35545) );
  CLKBUF_X2 U9956 ( .I(n31908), .Z(n34357) );
  INV_X2 U14940 ( .I(n15953), .ZN(n23539) );
  BUF_X4 U23171 ( .I(n23631), .Z(n32616) );
  CLKBUF_X4 U2215 ( .I(n23251), .Z(n23493) );
  INV_X2 U7097 ( .I(n16013), .ZN(n16774) );
  BUF_X2 U4270 ( .I(n38614), .Z(n36210) );
  NAND2_X1 U13178 ( .A1(n3174), .A2(n20322), .ZN(n3031) );
  CLKBUF_X2 U13341 ( .I(n23530), .Z(n18086) );
  BUF_X2 U28117 ( .I(n13038), .Z(n33349) );
  INV_X2 U18884 ( .I(n9395), .ZN(n23452) );
  INV_X1 U23135 ( .I(n23622), .ZN(n23621) );
  CLKBUF_X4 U20806 ( .I(n9395), .Z(n33080) );
  INV_X2 U9936 ( .I(n15122), .ZN(n17960) );
  INV_X1 U13330 ( .I(n23586), .ZN(n13897) );
  INV_X1 U6127 ( .I(n19389), .ZN(n35344) );
  INV_X1 U9971 ( .I(n38881), .ZN(n1307) );
  NOR2_X1 U13288 ( .A1(n13897), .A2(n39261), .ZN(n7629) );
  INV_X1 U7868 ( .I(n31164), .ZN(n23469) );
  NAND2_X1 U1915 ( .A1(n30789), .A2(n23321), .ZN(n30788) );
  NAND2_X1 U1940 ( .A1(n7387), .A2(n19686), .ZN(n23324) );
  NAND2_X1 U3447 ( .A1(n23216), .A2(n23606), .ZN(n18382) );
  INV_X1 U13206 ( .I(n23397), .ZN(n20066) );
  CLKBUF_X4 U24028 ( .I(n9968), .Z(n36011) );
  INV_X1 U13191 ( .I(n7224), .ZN(n11097) );
  INV_X1 U2153 ( .I(n9347), .ZN(n35279) );
  NAND2_X1 U27764 ( .A1(n19923), .A2(n19922), .ZN(n23633) );
  NAND2_X1 U13198 ( .A1(n16863), .A2(n15842), .ZN(n7487) );
  INV_X1 U16327 ( .I(n37957), .ZN(n2512) );
  INV_X1 U25120 ( .I(n20509), .ZN(n24059) );
  INV_X1 U5277 ( .I(n23777), .ZN(n12857) );
  NOR2_X1 U2159 ( .A1(n1616), .A2(n10110), .ZN(n10109) );
  INV_X1 U13065 ( .I(n23663), .ZN(n7360) );
  INV_X1 U13075 ( .I(n14220), .ZN(n23716) );
  INV_X1 U1808 ( .I(n18602), .ZN(n24203) );
  INV_X1 U2371 ( .I(n19949), .ZN(n20457) );
  CLKBUF_X2 U3544 ( .I(n19949), .Z(n277) );
  CLKBUF_X2 U9823 ( .I(n14471), .Z(n10152) );
  CLKBUF_X2 U9819 ( .I(n24095), .Z(n23694) );
  BUF_X2 U3822 ( .I(n8250), .Z(n30311) );
  CLKBUF_X2 U3316 ( .I(n19295), .Z(n10073) );
  CLKBUF_X2 U4702 ( .I(n16816), .Z(n32069) );
  INV_X2 U9808 ( .I(n23827), .ZN(n1276) );
  NOR2_X1 U24838 ( .A1(n24133), .A2(n19864), .ZN(n18277) );
  BUF_X2 U9820 ( .I(n16179), .Z(n9066) );
  INV_X1 U5302 ( .I(n24271), .ZN(n1124) );
  INV_X2 U1763 ( .I(n9371), .ZN(n33513) );
  CLKBUF_X4 U1797 ( .I(n15754), .Z(n3869) );
  CLKBUF_X4 U27662 ( .I(n24420), .Z(n19584) );
  CLKBUF_X4 U1132 ( .I(n18790), .Z(n16081) );
  BUF_X1 U13745 ( .I(n94), .Z(n34783) );
  INV_X2 U2028 ( .I(n15385), .ZN(n19382) );
  INV_X1 U5967 ( .I(n24370), .ZN(n12580) );
  INV_X2 U8582 ( .I(n24381), .ZN(n24214) );
  CLKBUF_X1 U19754 ( .I(n24169), .Z(n35384) );
  INV_X1 U28796 ( .I(n24412), .ZN(n24112) );
  BUF_X2 U5319 ( .I(n24427), .Z(n3142) );
  INV_X2 U12971 ( .I(n800), .ZN(n18466) );
  NOR2_X1 U9786 ( .A1(n24168), .A2(n24169), .ZN(n4821) );
  INV_X1 U14752 ( .I(n32250), .ZN(n3190) );
  NAND2_X1 U1982 ( .A1(n23845), .A2(n34620), .ZN(n17584) );
  INV_X2 U22797 ( .I(n3142), .ZN(n32937) );
  NAND2_X1 U28804 ( .A1(n24137), .A2(n17040), .ZN(n24138) );
  NOR2_X1 U12861 ( .A1(n24398), .A2(n12801), .ZN(n12800) );
  NOR2_X1 U25570 ( .A1(n24081), .A2(n1126), .ZN(n24082) );
  AOI21_X1 U12938 ( .A1(n1034), .A2(n305), .B(n4286), .ZN(n5014) );
  BUF_X2 U26853 ( .I(n19499), .Z(n36376) );
  NAND2_X1 U12602 ( .A1(n34637), .A2(n4051), .ZN(n4050) );
  NOR2_X1 U5337 ( .A1(n10783), .A2(n31003), .ZN(n10777) );
  INV_X2 U6932 ( .I(n24903), .ZN(n20155) );
  INV_X2 U18783 ( .I(n24799), .ZN(n24655) );
  CLKBUF_X4 U5074 ( .I(n14283), .Z(n19) );
  INV_X2 U12728 ( .I(n17087), .ZN(n19868) );
  CLKBUF_X4 U1945 ( .I(n9385), .Z(n4973) );
  CLKBUF_X4 U3976 ( .I(n32831), .Z(n30843) );
  CLKBUF_X4 U30856 ( .I(n7810), .Z(n3076) );
  INV_X2 U23317 ( .I(n24668), .ZN(n24750) );
  NOR2_X1 U1675 ( .A1(n24735), .A2(n24814), .ZN(n33818) );
  CLKBUF_X4 U3785 ( .I(n12686), .Z(n8314) );
  INV_X1 U12648 ( .I(n36955), .ZN(n3122) );
  INV_X2 U6909 ( .I(n6357), .ZN(n24686) );
  BUF_X2 U17781 ( .I(n24877), .Z(n33705) );
  INV_X1 U19777 ( .I(n24566), .ZN(n3624) );
  CLKBUF_X4 U27110 ( .I(n24883), .Z(n18114) );
  NAND2_X1 U6968 ( .A1(n14338), .A2(n24762), .ZN(n12632) );
  NAND2_X1 U27670 ( .A1(n24840), .A2(n24843), .ZN(n19597) );
  INV_X2 U22944 ( .I(n24250), .ZN(n24733) );
  INV_X1 U17383 ( .I(n24763), .ZN(n6023) );
  NAND2_X1 U9666 ( .A1(n31722), .A2(n1582), .ZN(n16669) );
  NAND2_X1 U24858 ( .A1(n4601), .A2(n20926), .ZN(n20925) );
  NAND2_X1 U3490 ( .A1(n15688), .A2(n2018), .ZN(n14782) );
  NAND2_X1 U1785 ( .A1(n17495), .A2(n34947), .ZN(n36672) );
  NAND2_X1 U12550 ( .A1(n10115), .A2(n4688), .ZN(n7321) );
  AOI22_X1 U21908 ( .A1(n32400), .A2(n13901), .B1(n38973), .B2(n13903), .ZN(
        n12817) );
  OAI21_X1 U26868 ( .A1(n34115), .A2(n9277), .B(n14936), .ZN(n14935) );
  NOR2_X1 U11218 ( .A1(n1119), .A2(n30915), .ZN(n31144) );
  NAND2_X1 U1573 ( .A1(n13746), .A2(n24832), .ZN(n30930) );
  NAND2_X1 U29350 ( .A1(n25052), .A2(n1273), .ZN(n36669) );
  NAND2_X1 U12539 ( .A1(n18844), .A2(n6336), .ZN(n24580) );
  NAND2_X1 U5931 ( .A1(n2076), .A2(n2075), .ZN(n36295) );
  OAI21_X1 U20341 ( .A1(n15849), .A2(n24648), .B(n15848), .ZN(n32087) );
  NAND2_X1 U27669 ( .A1(n19597), .A2(n24841), .ZN(n19596) );
  NAND2_X1 U2216 ( .A1(n31520), .A2(n31891), .ZN(n33043) );
  CLKBUF_X4 U9600 ( .I(n8542), .Z(n30761) );
  INV_X1 U1709 ( .I(n25016), .ZN(n34653) );
  INV_X1 U5853 ( .I(n39600), .ZN(n34856) );
  CLKBUF_X4 U9596 ( .I(n7328), .Z(n5208) );
  CLKBUF_X2 U11907 ( .I(n25569), .Z(n31004) );
  CLKBUF_X4 U12482 ( .I(n25309), .Z(n25469) );
  CLKBUF_X4 U4547 ( .I(n10584), .Z(n31780) );
  BUF_X2 U4527 ( .I(n835), .Z(n32580) );
  BUF_X2 U2640 ( .I(n25421), .Z(n12309) );
  CLKBUF_X2 U12477 ( .I(n25598), .Z(n9815) );
  CLKBUF_X2 U6252 ( .I(n5709), .Z(n5519) );
  CLKBUF_X4 U8181 ( .I(n13018), .Z(n12500) );
  BUF_X2 U9569 ( .I(n25694), .Z(n19767) );
  CLKBUF_X4 U17341 ( .I(n25613), .Z(n18031) );
  INV_X1 U17603 ( .I(n25158), .ZN(n13811) );
  CLKBUF_X4 U9571 ( .I(n25552), .Z(n12825) );
  CLKBUF_X2 U4353 ( .I(n16203), .Z(n3985) );
  CLKBUF_X4 U8183 ( .I(n25722), .Z(n19367) );
  CLKBUF_X2 U4522 ( .I(n252), .Z(n32868) );
  CLKBUF_X2 U1665 ( .I(n33948), .Z(n19548) );
  NOR2_X1 U3375 ( .A1(n18545), .A2(n19589), .ZN(n14257) );
  CLKBUF_X2 U5325 ( .I(n25355), .Z(n25583) );
  CLKBUF_X2 U30302 ( .I(n34576), .Z(n36816) );
  CLKBUF_X4 U9535 ( .I(n730), .Z(n7986) );
  NAND2_X1 U7460 ( .A1(n15541), .A2(n1552), .ZN(n25349) );
  NOR2_X1 U1676 ( .A1(n35508), .A2(n36162), .ZN(n36142) );
  AOI21_X1 U15988 ( .A1(n18545), .A2(n19589), .B(n25502), .ZN(n15254) );
  CLKBUF_X4 U23740 ( .I(n25696), .Z(n32722) );
  INV_X2 U26410 ( .I(n7075), .ZN(n33115) );
  CLKBUF_X1 U5039 ( .I(n31010), .Z(n35696) );
  CLKBUF_X2 U10742 ( .I(n14805), .Z(n34436) );
  NOR2_X1 U15948 ( .A1(n31619), .A2(n33115), .ZN(n7924) );
  NAND2_X1 U5480 ( .A1(n17815), .A2(n36792), .ZN(n4216) );
  NOR2_X1 U819 ( .A1(n4469), .A2(n1545), .ZN(n4465) );
  NAND2_X1 U9448 ( .A1(n10788), .A2(n1534), .ZN(n10787) );
  NOR2_X1 U12333 ( .A1(n6748), .A2(n25666), .ZN(n25667) );
  NAND2_X1 U12320 ( .A1(n12462), .A2(n12463), .ZN(n12996) );
  AOI22_X1 U29082 ( .A1(n25633), .A2(n25728), .B1(n16168), .B2(n18294), .ZN(
        n25634) );
  OAI21_X1 U29061 ( .A1(n1022), .A2(n14413), .B(n36019), .ZN(n25515) );
  NAND2_X1 U27461 ( .A1(n36475), .A2(n36793), .ZN(n20626) );
  OAI21_X1 U9467 ( .A1(n25528), .A2(n517), .B(n25333), .ZN(n1992) );
  NOR2_X1 U19228 ( .A1(n25478), .A2(n8980), .ZN(n8979) );
  INV_X1 U11749 ( .I(n34572), .ZN(n34571) );
  NAND2_X1 U17665 ( .A1(n15404), .A2(n14679), .ZN(n4888) );
  NAND2_X1 U27104 ( .A1(n33204), .A2(n30381), .ZN(n15445) );
  AOI21_X1 U18322 ( .A1(n30633), .A2(n32279), .B(n19398), .ZN(n32278) );
  OAI21_X1 U12241 ( .A1(n17868), .A2(n19235), .B(n19234), .ZN(n25573) );
  NAND2_X1 U3364 ( .A1(n11549), .A2(n25621), .ZN(n10041) );
  NAND2_X1 U14629 ( .A1(n4756), .A2(n4754), .ZN(n34886) );
  NAND2_X1 U12294 ( .A1(n6173), .A2(n6172), .ZN(n6171) );
  INV_X2 U7920 ( .I(n26106), .ZN(n1017) );
  BUF_X1 U4994 ( .I(n37393), .Z(n34417) );
  INV_X2 U12206 ( .I(n37393), .ZN(n11848) );
  CLKBUF_X4 U3679 ( .I(n26115), .Z(n30302) );
  INV_X2 U725 ( .I(n33293), .ZN(n1106) );
  NAND2_X1 U4050 ( .A1(n26093), .A2(n26329), .ZN(n15003) );
  CLKBUF_X4 U2706 ( .I(n33909), .Z(n31205) );
  INV_X2 U16974 ( .I(n26124), .ZN(n5098) );
  INV_X2 U18849 ( .I(n32691), .ZN(n26003) );
  CLKBUF_X4 U4302 ( .I(n7901), .Z(n3013) );
  BUF_X2 U7103 ( .I(n33644), .Z(n31263) );
  CLKBUF_X4 U6848 ( .I(n18032), .Z(n16407) );
  CLKBUF_X4 U4470 ( .I(n34609), .Z(n30883) );
  INV_X2 U775 ( .I(n37730), .ZN(n1524) );
  CLKBUF_X4 U3090 ( .I(n18994), .Z(n7767) );
  INV_X2 U3259 ( .I(n17400), .ZN(n1011) );
  CLKBUF_X4 U1923 ( .I(n26070), .Z(n11858) );
  AOI21_X1 U27612 ( .A1(n39729), .A2(n33237), .B(n35744), .ZN(n19439) );
  AOI21_X1 U12096 ( .A1(n949), .A2(n18003), .B(n18002), .ZN(n11010) );
  NOR2_X1 U26145 ( .A1(n25459), .A2(n33348), .ZN(n18314) );
  OAI21_X1 U12122 ( .A1(n931), .A2(n7460), .B(n13067), .ZN(n13066) );
  NAND2_X1 U1255 ( .A1(n34647), .A2(n39676), .ZN(n34646) );
  NAND2_X1 U29110 ( .A1(n25959), .A2(n25793), .ZN(n25794) );
  OAI21_X1 U23049 ( .A1(n25957), .A2(n11552), .B(n11551), .ZN(n18745) );
  AOI21_X1 U8004 ( .A1(n12569), .A2(n26012), .B(n39661), .ZN(n4401) );
  INV_X1 U6826 ( .I(n26072), .ZN(n11859) );
  NAND2_X1 U5698 ( .A1(n36766), .A2(n26214), .ZN(n25833) );
  NOR2_X1 U4355 ( .A1(n195), .A2(n30436), .ZN(n36300) );
  INV_X1 U11799 ( .I(n8858), .ZN(n9378) );
  NAND2_X1 U9039 ( .A1(n25857), .A2(n26072), .ZN(n34275) );
  AOI21_X1 U672 ( .A1(n10889), .A2(n7110), .B(n7111), .ZN(n9983) );
  NAND2_X1 U3345 ( .A1(n12105), .A2(n34685), .ZN(n10016) );
  NAND2_X1 U7119 ( .A1(n25651), .A2(n39015), .ZN(n3914) );
  OAI21_X1 U1893 ( .A1(n11859), .A2(n26071), .B(n15796), .ZN(n17187) );
  INV_X1 U6577 ( .I(n26565), .ZN(n1507) );
  CLKBUF_X4 U1138 ( .I(n14393), .Z(n37024) );
  INV_X1 U7101 ( .I(n9174), .ZN(n10269) );
  NAND2_X1 U12021 ( .A1(n34595), .A2(n36293), .ZN(n9077) );
  CLKBUF_X2 U4427 ( .I(n18490), .Z(n31941) );
  BUF_X2 U11997 ( .I(n26565), .Z(n19289) );
  CLKBUF_X4 U8798 ( .I(n2055), .Z(n33812) );
  CLKBUF_X4 U4430 ( .I(n14346), .Z(n33308) );
  CLKBUF_X1 U5682 ( .I(n17455), .Z(n36765) );
  INV_X2 U8831 ( .I(n26234), .ZN(n7603) );
  CLKBUF_X4 U4424 ( .I(n26559), .Z(n32464) );
  CLKBUF_X2 U15549 ( .I(n20613), .Z(n19700) );
  CLKBUF_X2 U17950 ( .I(n3827), .Z(n36480) );
  CLKBUF_X2 U4390 ( .I(n36355), .Z(n31502) );
  CLKBUF_X4 U5662 ( .I(n26809), .Z(n14377) );
  CLKBUF_X2 U11963 ( .I(n26796), .Z(n7725) );
  CLKBUF_X2 U2698 ( .I(n14440), .Z(n7516) );
  CLKBUF_X2 U11075 ( .I(n14488), .Z(n34484) );
  OR2_X1 U21952 ( .A1(n35197), .A2(n19442), .Z(n14659) );
  CLKBUF_X2 U27962 ( .I(n384), .Z(n33333) );
  CLKBUF_X2 U9357 ( .I(n14080), .Z(n14079) );
  CLKBUF_X4 U21256 ( .I(n8413), .Z(n32256) );
  CLKBUF_X2 U3996 ( .I(n26885), .Z(n7305) );
  CLKBUF_X4 U7181 ( .I(n14962), .Z(n34892) );
  INV_X2 U21017 ( .I(n8479), .ZN(n10187) );
  NAND2_X1 U11834 ( .A1(n18575), .A2(n106), .ZN(n20790) );
  INV_X1 U15099 ( .I(n11224), .ZN(n11226) );
  BUF_X2 U3939 ( .I(n17252), .Z(n33301) );
  INV_X1 U11892 ( .I(n26652), .ZN(n26738) );
  NAND2_X1 U27513 ( .A1(n26798), .A2(n26797), .ZN(n19210) );
  NAND2_X1 U11803 ( .A1(n16049), .A2(n26721), .ZN(n27124) );
  INV_X2 U530 ( .I(n26751), .ZN(n26898) );
  NOR2_X1 U3933 ( .A1(n26987), .A2(n26986), .ZN(n5480) );
  NAND2_X1 U9315 ( .A1(n26907), .A2(n26926), .ZN(n26912) );
  NAND2_X1 U11524 ( .A1(n26912), .A2(n9166), .ZN(n30958) );
  OAI21_X1 U15275 ( .A1(n11616), .A2(n26751), .B(n26738), .ZN(n34974) );
  NOR2_X1 U12023 ( .A1(n15594), .A2(n20797), .ZN(n9015) );
  NAND2_X1 U19272 ( .A1(n17514), .A2(n6555), .ZN(n6554) );
  OAI21_X1 U16934 ( .A1(n4459), .A2(n12549), .B(n33952), .ZN(n4580) );
  NOR2_X1 U30395 ( .A1(n26843), .A2(n1002), .ZN(n36846) );
  NAND2_X1 U11867 ( .A1(n26911), .A2(n26910), .ZN(n12659) );
  NAND2_X1 U14290 ( .A1(n16939), .A2(n14659), .ZN(n34830) );
  NAND2_X1 U5625 ( .A1(n31226), .A2(n31225), .ZN(n36938) );
  OR2_X1 U11811 ( .A1(n26898), .A2(n15317), .Z(n5172) );
  NAND2_X1 U7328 ( .A1(n26352), .A2(n34843), .ZN(n5590) );
  OAI21_X1 U3050 ( .A1(n17279), .A2(n17278), .B(n1236), .ZN(n15550) );
  NAND2_X1 U25286 ( .A1(n9619), .A2(n17786), .ZN(n36521) );
  NAND2_X1 U523 ( .A1(n4689), .A2(n9075), .ZN(n26733) );
  INV_X2 U14128 ( .I(n1788), .ZN(n8137) );
  INV_X1 U5627 ( .I(n26760), .ZN(n11517) );
  NOR2_X1 U12726 ( .A1(n9015), .A2(n9014), .ZN(n36501) );
  INV_X1 U11789 ( .I(n14280), .ZN(n3136) );
  CLKBUF_X2 U11747 ( .I(n5831), .Z(n3513) );
  NAND2_X1 U11774 ( .A1(n26138), .A2(n11522), .ZN(n15685) );
  CLKBUF_X2 U15140 ( .I(n27358), .Z(n34952) );
  CLKBUF_X4 U5767 ( .I(n21272), .Z(n2760) );
  CLKBUF_X2 U13593 ( .I(n19135), .Z(n34769) );
  CLKBUF_X2 U5888 ( .I(n27399), .Z(n18228) );
  CLKBUF_X1 U7361 ( .I(n27131), .Z(n7620) );
  INV_X2 U755 ( .I(n33662), .ZN(n14261) );
  BUF_X2 U4915 ( .I(n9267), .Z(n31672) );
  CLKBUF_X4 U7391 ( .I(n9037), .Z(n2522) );
  INV_X2 U8573 ( .I(n27288), .ZN(n1470) );
  NAND2_X1 U7819 ( .A1(n19334), .A2(n18195), .ZN(n9488) );
  INV_X2 U23329 ( .I(n17166), .ZN(n12074) );
  CLKBUF_X4 U7821 ( .I(n27275), .Z(n10677) );
  CLKBUF_X4 U5745 ( .I(n27435), .Z(n17754) );
  OAI21_X1 U18229 ( .A1(n18232), .A2(n19619), .B(n27271), .ZN(n19329) );
  AOI21_X1 U11644 ( .A1(n27273), .A2(n20244), .B(n38900), .ZN(n20243) );
  NOR2_X1 U406 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  NAND2_X1 U18566 ( .A1(n34520), .A2(n33803), .ZN(n7403) );
  NOR2_X1 U25327 ( .A1(n2208), .A2(n32557), .ZN(n33376) );
  NAND2_X1 U13598 ( .A1(n34770), .A2(n27388), .ZN(n36036) );
  NOR2_X1 U7414 ( .A1(n17354), .A2(n7894), .ZN(n18861) );
  NAND2_X1 U11582 ( .A1(n16360), .A2(n27273), .ZN(n14057) );
  CLKBUF_X1 U12138 ( .I(n27738), .Z(n31020) );
  INV_X1 U23651 ( .I(n27528), .ZN(n35986) );
  CLKBUF_X2 U3906 ( .I(n14456), .Z(n32783) );
  INV_X1 U30258 ( .I(n27843), .ZN(n36809) );
  CLKBUF_X4 U7704 ( .I(n18688), .Z(n1454) );
  CLKBUF_X2 U30386 ( .I(n28117), .Z(n36844) );
  CLKBUF_X4 U559 ( .I(n20531), .Z(n7635) );
  INV_X1 U371 ( .I(n21159), .ZN(n19417) );
  CLKBUF_X2 U7725 ( .I(n9775), .Z(n7591) );
  CLKBUF_X4 U5403 ( .I(n28093), .Z(n28214) );
  CLKBUF_X2 U17906 ( .I(n17533), .Z(n32324) );
  CLKBUF_X4 U3318 ( .I(n28125), .Z(n10254) );
  INV_X2 U7719 ( .I(n19435), .ZN(n1071) );
  CLKBUF_X4 U7720 ( .I(n28186), .Z(n15357) );
  CLKBUF_X2 U2421 ( .I(n8148), .Z(n288) );
  CLKBUF_X2 U22708 ( .I(n6990), .Z(n35827) );
  CLKBUF_X2 U19801 ( .I(n33955), .Z(n31966) );
  OR2_X1 U17964 ( .A1(n20531), .A2(n6640), .Z(n14618) );
  CLKBUF_X4 U4098 ( .I(n28188), .Z(n9969) );
  INV_X1 U4266 ( .I(n27989), .ZN(n33020) );
  OR3_X1 U4132 ( .A1(n9688), .A2(n17314), .A3(n32352), .Z(n27994) );
  NAND2_X1 U299 ( .A1(n13714), .A2(n1212), .ZN(n13663) );
  AOI21_X1 U22782 ( .A1(n15597), .A2(n20896), .B(n18603), .ZN(n11055) );
  INV_X1 U11340 ( .I(n28108), .ZN(n6789) );
  INV_X2 U3358 ( .I(n36838), .ZN(n28194) );
  OAI21_X1 U9047 ( .A1(n35607), .A2(n19280), .B(n13251), .ZN(n13250) );
  OAI21_X1 U7670 ( .A1(n35607), .A2(n1205), .B(n11147), .ZN(n6790) );
  AOI21_X1 U5490 ( .A1(n20993), .A2(n28045), .B(n4915), .ZN(n32869) );
  INV_X1 U5483 ( .I(n28420), .ZN(n18380) );
  NAND2_X1 U14234 ( .A1(n13250), .A2(n13249), .ZN(n5237) );
  NAND2_X1 U11329 ( .A1(n19324), .A2(n19325), .ZN(n5906) );
  NAND2_X1 U11189 ( .A1(n35657), .A2(n19946), .ZN(n4724) );
  NAND2_X1 U21877 ( .A1(n27891), .A2(n34447), .ZN(n14736) );
  CLKBUF_X4 U3675 ( .I(n28578), .Z(n34667) );
  CLKBUF_X4 U3619 ( .I(n9290), .Z(n5662) );
  BUF_X2 U3899 ( .I(n28595), .Z(n16295) );
  BUF_X2 U4421 ( .I(n1882), .Z(n31321) );
  CLKBUF_X2 U30153 ( .I(n20445), .Z(n36788) );
  NAND2_X1 U11179 ( .A1(n12487), .A2(n12486), .ZN(n7745) );
  CLKBUF_X4 U3900 ( .I(n6932), .Z(n30931) );
  BUF_X2 U9019 ( .I(n9575), .Z(n7555) );
  CLKBUF_X4 U7505 ( .I(n28396), .Z(n36814) );
  INV_X2 U260 ( .I(n28433), .ZN(n28458) );
  OAI22_X1 U29584 ( .A1(n7454), .A2(n36788), .B1(n28354), .B2(n28353), .ZN(
        n28355) );
  NAND2_X1 U18088 ( .A1(n28533), .A2(n8743), .ZN(n28504) );
  CLKBUF_X4 U3999 ( .I(n13880), .Z(n33843) );
  INV_X2 U9757 ( .I(n8743), .ZN(n17800) );
  INV_X2 U5477 ( .I(n28356), .ZN(n28611) );
  CLKBUF_X4 U28689 ( .I(n28494), .Z(n36609) );
  INV_X2 U7526 ( .I(n17800), .ZN(n5890) );
  NAND2_X1 U14818 ( .A1(n1430), .A2(n28726), .ZN(n12610) );
  CLKBUF_X4 U11167 ( .I(n28696), .Z(n9648) );
  NAND2_X1 U18299 ( .A1(n12610), .A2(n32178), .ZN(n12607) );
  NAND2_X1 U5420 ( .A1(n10361), .A2(n36567), .ZN(n31404) );
  NAND2_X1 U20539 ( .A1(n21188), .A2(n21190), .ZN(n18103) );
  NAND2_X1 U19562 ( .A1(n28366), .A2(n37081), .ZN(n16343) );
  NAND2_X1 U10992 ( .A1(n13060), .A2(n17045), .ZN(n7647) );
  OAI21_X1 U10947 ( .A1(n4025), .A2(n28746), .B(n4023), .ZN(n28752) );
  NAND2_X1 U3271 ( .A1(n35030), .A2(n15964), .ZN(n4878) );
  NOR2_X1 U19561 ( .A1(n17322), .A2(n37081), .ZN(n17321) );
  NAND2_X1 U229 ( .A1(n7478), .A2(n34305), .ZN(n2900) );
  AOI22_X1 U205 ( .A1(n9598), .A2(n17320), .B1(n17321), .B2(n10587), .ZN(
        n17338) );
  INV_X2 U16698 ( .I(n7710), .ZN(n29832) );
  BUF_X2 U6574 ( .I(n29249), .Z(n18242) );
  INV_X1 U4121 ( .I(n28869), .ZN(n31841) );
  OAI21_X1 U6808 ( .A1(n16656), .A2(n16655), .B(n5645), .ZN(n33375) );
  CLKBUF_X4 U4298 ( .I(n18305), .Z(n467) );
  CLKBUF_X2 U17403 ( .I(n29903), .Z(n18222) );
  BUF_X2 U8046 ( .I(n11415), .Z(n482) );
  CLKBUF_X1 U18373 ( .I(n38186), .Z(n33404) );
  CLKBUF_X2 U2781 ( .I(n15853), .Z(n105) );
  CLKBUF_X4 U1671 ( .I(n28899), .Z(n29491) );
  OAI21_X1 U19034 ( .A1(n30229), .A2(n19765), .B(n10590), .ZN(n14281) );
  INV_X2 U97 ( .I(n17238), .ZN(n1175) );
  NAND2_X1 U2444 ( .A1(n8726), .A2(n29286), .ZN(n32648) );
  NAND2_X1 U109 ( .A1(n20405), .A2(n35695), .ZN(n35057) );
  INV_X1 U4094 ( .I(n21290), .ZN(n32499) );
  AOI21_X1 U7398 ( .A1(n29629), .A2(n31511), .B(n13722), .ZN(n2554) );
  BUF_X1 U4101 ( .I(n30049), .Z(n32628) );
  NOR2_X1 U24292 ( .A1(n30165), .A2(n14184), .ZN(n14183) );
  NAND2_X1 U30605 ( .A1(n36893), .A2(n29389), .ZN(n8147) );
  NAND2_X1 U21880 ( .A1(n29861), .A2(n17779), .ZN(n17302) );
  NAND2_X1 U23989 ( .A1(n32762), .A2(n30001), .ZN(n15644) );
  NAND2_X1 U10651 ( .A1(n29953), .A2(n19196), .ZN(n19195) );
  BUF_X2 U10594 ( .I(n29930), .Z(n9591) );
  CLKBUF_X4 U17354 ( .I(n19260), .Z(n18384) );
  BUF_X2 U10618 ( .I(n29530), .Z(n19362) );
  CLKBUF_X2 U5340 ( .I(n30178), .Z(n35899) );
  INV_X4 U27 ( .I(n9231), .ZN(n30024) );
  AOI21_X1 U29181 ( .A1(n35175), .A2(n30093), .B(n1382), .ZN(n30083) );
  NAND3_X1 U24024 ( .A1(n9263), .A2(n9264), .A3(n32508), .ZN(n36005) );
  OR2_X1 U4291 ( .A1(n30180), .A2(n17997), .Z(n896) );
  AOI22_X1 U9638 ( .A1(n29669), .A2(n29668), .B1(n29676), .B2(n29670), .ZN(
        n34323) );
  NOR2_X1 U4 ( .A1(n13606), .A2(n29811), .ZN(n36365) );
  CLKBUF_X2 U8792 ( .I(Key[112]), .Z(n19735) );
  CLKBUF_X2 U6461 ( .I(Key[100]), .Z(n19674) );
  CLKBUF_X2 U10457 ( .I(Key[123]), .Z(n28821) );
  CLKBUF_X2 U8754 ( .I(Key[114]), .Z(n19943) );
  CLKBUF_X2 U8758 ( .I(Key[34]), .Z(n29666) );
  CLKBUF_X2 U10475 ( .I(Key[72]), .Z(n30104) );
  CLKBUF_X2 U10483 ( .I(Key[115]), .Z(n19729) );
  BUF_X2 U8784 ( .I(Key[159]), .Z(n19835) );
  INV_X1 U4064 ( .I(n19786), .ZN(n33866) );
  INV_X1 U30194 ( .I(n19943), .ZN(n33661) );
  INV_X1 U27794 ( .I(n19883), .ZN(n36513) );
  AOI22_X1 U16870 ( .A1(n21902), .A2(n526), .B1(n35921), .B2(n7304), .ZN(
        n21904) );
  NOR2_X1 U25073 ( .A1(n21748), .A2(n21713), .ZN(n21649) );
  CLKBUF_X2 U6313 ( .I(n22042), .Z(n36428) );
  INV_X2 U1444 ( .I(n22306), .ZN(n1335) );
  BUF_X2 U4848 ( .I(n8431), .Z(n32817) );
  OR2_X1 U25402 ( .A1(n22293), .A2(n9265), .Z(n14498) );
  CLKBUF_X2 U29160 ( .I(n22348), .Z(n36641) );
  CLKBUF_X4 U2096 ( .I(n22549), .Z(n7055) );
  NAND2_X2 U1376 ( .A1(n17339), .A2(n17340), .ZN(n22700) );
  CLKBUF_X4 U21821 ( .I(n2126), .Z(n36596) );
  CLKBUF_X2 U4801 ( .I(n23214), .Z(n32590) );
  INV_X2 U23587 ( .I(n9797), .ZN(n23061) );
  INV_X2 U6685 ( .I(n22895), .ZN(n20174) );
  OAI21_X1 U8464 ( .A1(n9770), .A2(n9769), .B(n22964), .ZN(n12816) );
  INV_X2 U17624 ( .I(n388), .ZN(n1635) );
  CLKBUF_X4 U2289 ( .I(n14235), .Z(n35963) );
  CLKBUF_X2 U6152 ( .I(n5357), .Z(n35130) );
  CLKBUF_X4 U6756 ( .I(n17508), .Z(n15176) );
  CLKBUF_X1 U27904 ( .I(n23337), .Z(n36530) );
  AOI21_X1 U1163 ( .A1(n35664), .A2(n12597), .B(n11969), .ZN(n20222) );
  NOR2_X1 U13315 ( .A1(n16774), .A2(n37431), .ZN(n16863) );
  CLKBUF_X1 U14360 ( .I(n3609), .Z(n34844) );
  CLKBUF_X2 U3979 ( .I(n18602), .Z(n33314) );
  CLKBUF_X2 U8354 ( .I(n8193), .Z(n5599) );
  CLKBUF_X2 U4171 ( .I(n14463), .Z(n370) );
  INV_X2 U17265 ( .I(n24203), .ZN(n7210) );
  CLKBUF_X1 U4537 ( .I(n24202), .Z(n18304) );
  BUF_X2 U5204 ( .I(n35134), .Z(n35690) );
  NAND2_X1 U9726 ( .A1(n24294), .A2(n8463), .ZN(n9083) );
  AOI21_X1 U2030 ( .A1(n24214), .A2(n6567), .B(n34673), .ZN(n34252) );
  NOR2_X1 U12603 ( .A1(n4053), .A2(n1031), .ZN(n34637) );
  INV_X1 U8282 ( .I(n24737), .ZN(n1582) );
  INV_X2 U5072 ( .I(n31986), .ZN(n24648) );
  NAND2_X1 U27711 ( .A1(n39196), .A2(n19565), .ZN(n6169) );
  NAND2_X1 U26565 ( .A1(n24839), .A2(n34906), .ZN(n24840) );
  NAND2_X1 U17737 ( .A1(n6187), .A2(n24806), .ZN(n6183) );
  CLKBUF_X2 U17983 ( .I(n31181), .Z(n35972) );
  CLKBUF_X4 U4539 ( .I(n15030), .Z(n518) );
  CLKBUF_X4 U4222 ( .I(n24924), .Z(n449) );
  CLKBUF_X2 U5866 ( .I(n25266), .Z(n35953) );
  BUF_X2 U3920 ( .I(n15907), .Z(n371) );
  CLKBUF_X2 U17442 ( .I(n20416), .Z(n31574) );
  CLKBUF_X2 U5827 ( .I(n20838), .Z(n36019) );
  CLKBUF_X2 U12757 ( .I(n25158), .Z(n25756) );
  INV_X1 U23936 ( .I(n25727), .ZN(n16168) );
  CLKBUF_X2 U5471 ( .I(n17594), .Z(n13460) );
  NAND2_X1 U27987 ( .A1(n15329), .A2(n15172), .ZN(n33204) );
  AOI21_X1 U2648 ( .A1(n32172), .A2(n16677), .B(n25449), .ZN(n4620) );
  AOI21_X1 U11751 ( .A1(n20888), .A2(n19463), .B(n25616), .ZN(n34572) );
  NOR2_X1 U9409 ( .A1(n12768), .A2(n9944), .ZN(n34309) );
  NOR2_X1 U12292 ( .A1(n8123), .A2(n8122), .ZN(n8121) );
  INV_X1 U754 ( .I(n9833), .ZN(n19121) );
  BUF_X2 U6868 ( .I(n26106), .Z(n18162) );
  BUF_X2 U4489 ( .I(n26215), .Z(n9868) );
  INV_X1 U17021 ( .I(n15992), .ZN(n35155) );
  INV_X2 U8039 ( .I(n14890), .ZN(n25928) );
  BUF_X2 U25607 ( .I(n10834), .Z(n32979) );
  BUF_X2 U4475 ( .I(n21204), .Z(n31340) );
  BUF_X2 U5540 ( .I(n19240), .Z(n33474) );
  CLKBUF_X2 U4977 ( .I(n26131), .Z(n35109) );
  BUF_X2 U3950 ( .I(n25900), .Z(n33327) );
  NAND2_X1 U1342 ( .A1(n1019), .A2(n35151), .ZN(n34647) );
  OAI21_X1 U5442 ( .A1(n11835), .A2(n11833), .B(n19740), .ZN(n12523) );
  NAND2_X1 U11715 ( .A1(n34573), .A2(n34574), .ZN(n34565) );
  NAND2_X1 U21264 ( .A1(n25110), .A2(n25510), .ZN(n18864) );
  CLKBUF_X2 U1598 ( .I(n26968), .Z(n13181) );
  AND2_X1 U10521 ( .A1(n34160), .A2(n26968), .Z(n2969) );
  CLKBUF_X2 U11966 ( .I(n20891), .Z(n19972) );
  CLKBUF_X2 U3941 ( .I(n866), .Z(n31701) );
  BUF_X2 U7229 ( .I(n20704), .Z(n9178) );
  CLKBUF_X2 U11951 ( .I(n26630), .Z(n26811) );
  CLKBUF_X2 U4398 ( .I(n11224), .Z(n33726) );
  NAND2_X1 U2564 ( .A1(n26860), .A2(n12682), .ZN(n11652) );
  INV_X1 U21897 ( .I(n35732), .ZN(n30347) );
  NOR2_X1 U20632 ( .A1(n26812), .A2(n33849), .ZN(n12795) );
  BUF_X2 U2735 ( .I(n27436), .Z(n30671) );
  CLKBUF_X2 U11707 ( .I(n27252), .Z(n9756) );
  BUF_X2 U5599 ( .I(n35051), .Z(n34689) );
  CLKBUF_X4 U760 ( .I(n8537), .Z(n31875) );
  AND2_X2 U720 ( .A1(n8798), .A2(n27349), .Z(n27351) );
  CLKBUF_X2 U23578 ( .I(n27253), .Z(n32697) );
  CLKBUF_X2 U4342 ( .I(n30358), .Z(n31683) );
  INV_X1 U3610 ( .I(n27492), .ZN(n4885) );
  BUF_X2 U5401 ( .I(n36838), .Z(n19657) );
  CLKBUF_X4 U5474 ( .I(n28651), .Z(n35830) );
  CLKBUF_X2 U11115 ( .I(n28596), .Z(n9598) );
  CLKBUF_X2 U4852 ( .I(n33100), .Z(n34915) );
  CLKBUF_X2 U17300 ( .I(n5028), .Z(n32595) );
  BUF_X2 U17206 ( .I(n12168), .Z(n33647) );
  NAND2_X1 U23047 ( .A1(n10618), .A2(n32286), .ZN(n35875) );
  BUF_X2 U25962 ( .I(n29052), .Z(n33041) );
  CLKBUF_X2 U6102 ( .I(n29120), .Z(n29286) );
  BUF_X2 U24059 ( .I(n21299), .Z(n32777) );
  NAND2_X1 U19231 ( .A1(n8445), .A2(n6496), .ZN(n30001) );
  BUF_X2 U2847 ( .I(n18896), .Z(n13705) );
  CLKBUF_X4 U16847 ( .I(n17347), .Z(n6252) );
  INV_X2 U6505 ( .I(n13559), .ZN(n1382) );
  INV_X1 U8839 ( .I(n3896), .ZN(n3897) );
  BUF_X4 U5675 ( .I(n7959), .Z(n36244) );
  BUF_X4 U6382 ( .I(n21387), .Z(n18417) );
  NAND2_X1 U9503 ( .A1(n32053), .A2(n7915), .ZN(n30808) );
  NAND2_X2 U405 ( .A1(n30370), .A2(n28118), .ZN(n20410) );
  BUF_X2 U11968 ( .I(n26770), .Z(n19442) );
  OAI21_X2 U27212 ( .A1(n19660), .A2(n19659), .B(n23070), .ZN(n19360) );
  NAND2_X1 U4311 ( .A1(n19596), .A2(n19595), .ZN(n14826) );
  OR2_X1 U2885 ( .A1(n37079), .A2(n8604), .Z(n27989) );
  NOR2_X2 U27188 ( .A1(n34923), .A2(n19350), .ZN(n36441) );
  OAI21_X2 U5038 ( .A1(n24685), .A2(n12460), .B(n7930), .ZN(n8107) );
  NAND2_X2 U30500 ( .A1(n33284), .A2(n15876), .ZN(n29401) );
  NOR2_X2 U1215 ( .A1(n30936), .A2(n25467), .ZN(n33270) );
  INV_X4 U25361 ( .I(n12049), .ZN(n32946) );
  BUF_X4 U2149 ( .I(n23963), .Z(n30612) );
  NOR2_X2 U12851 ( .A1(n24336), .A2(n24332), .ZN(n24333) );
  BUF_X4 U6777 ( .I(n855), .Z(n12373) );
  INV_X4 U5280 ( .I(n12953), .ZN(n1603) );
  INV_X4 U6425 ( .I(n21692), .ZN(n1355) );
  NOR2_X2 U8062 ( .A1(n1018), .A2(n31626), .ZN(n1852) );
  BUF_X2 U3978 ( .I(n205), .Z(n33379) );
  BUF_X4 U15539 ( .I(n4322), .Z(n32974) );
  NAND2_X1 U13480 ( .A1(n16955), .A2(n16954), .ZN(n22945) );
  NOR2_X2 U13923 ( .A1(n14577), .A2(n21932), .ZN(n18025) );
  NOR2_X2 U12758 ( .A1(n10691), .A2(n10690), .ZN(n10689) );
  NAND3_X2 U20527 ( .A1(n13738), .A2(n13739), .A3(n29286), .ZN(n35502) );
  OAI21_X2 U19520 ( .A1(n23596), .A2(n36720), .B(n23595), .ZN(n14993) );
  OR2_X1 U4154 ( .A1(n2572), .A2(n18433), .Z(n32636) );
  INV_X4 U21069 ( .I(n36214), .ZN(n14196) );
  NAND2_X2 U17660 ( .A1(n4948), .A2(n17465), .ZN(n12415) );
  NOR2_X2 U17271 ( .A1(n7631), .A2(n8757), .ZN(n6519) );
  NAND2_X2 U18926 ( .A1(n9700), .A2(n9698), .ZN(n31835) );
  NAND2_X2 U360 ( .A1(n36478), .A2(n28537), .ZN(n4228) );
  INV_X2 U7154 ( .I(n26009), .ZN(n26158) );
  BUF_X2 U4112 ( .I(n30154), .Z(n33081) );
  NAND2_X2 U14850 ( .A1(n7941), .A2(n31318), .ZN(n31654) );
  NOR2_X2 U3491 ( .A1(n26140), .A2(n11485), .ZN(n11484) );
  NAND2_X2 U18774 ( .A1(n24770), .A2(n5957), .ZN(n24351) );
  INV_X4 U12968 ( .I(n921), .ZN(n9508) );
  NOR2_X1 U12925 ( .A1(n10695), .A2(n1283), .ZN(n10694) );
  INV_X2 U2140 ( .I(n8113), .ZN(n1993) );
  INV_X2 U2951 ( .I(n29166), .ZN(n36928) );
  BUF_X4 U800 ( .I(n39583), .Z(n33088) );
  NAND2_X2 U2615 ( .A1(n19075), .A2(n21778), .ZN(n36346) );
  NOR2_X2 U11756 ( .A1(n16401), .A2(n12177), .ZN(n8332) );
  INV_X2 U5781 ( .I(n22075), .ZN(n22039) );
  NAND3_X2 U27543 ( .A1(n1299), .A2(n33538), .A3(n19283), .ZN(n23266) );
  NOR2_X2 U144 ( .A1(n29286), .A2(n1062), .ZN(n11409) );
  AND2_X2 U11724 ( .A1(n27583), .A2(n27304), .Z(n8696) );
  OAI21_X1 U13414 ( .A1(n23050), .A2(n9854), .B(n4566), .ZN(n4565) );
  NAND2_X2 U12781 ( .A1(n24135), .A2(n24464), .ZN(n7033) );
  NOR2_X2 U29924 ( .A1(n4182), .A2(n33531), .ZN(n33530) );
  BUF_X4 U18667 ( .I(n26553), .Z(n31791) );
  OAI21_X2 U16476 ( .A1(n11709), .A2(n11708), .B(n11707), .ZN(n17415) );
  NOR2_X1 U22564 ( .A1(n13547), .A2(n24029), .ZN(n35803) );
  BUF_X4 U2686 ( .I(n17220), .Z(n36384) );
  NAND2_X2 U3695 ( .A1(n26802), .A2(n26747), .ZN(n4458) );
  INV_X4 U19982 ( .I(n35422), .ZN(n15102) );
  INV_X4 U14442 ( .I(n27275), .ZN(n4434) );
  BUF_X4 U16578 ( .I(n24104), .Z(n24328) );
  NAND2_X2 U2858 ( .A1(n29483), .A2(n29643), .ZN(n29443) );
  INV_X1 U14919 ( .I(n21776), .ZN(n34922) );
  INV_X1 U22578 ( .I(n10656), .ZN(n21868) );
  INV_X1 U2288 ( .I(n7062), .ZN(n2990) );
  INV_X1 U5009 ( .I(n12670), .ZN(n21895) );
  INV_X1 U22214 ( .I(n18027), .ZN(n14769) );
  BUF_X2 U3520 ( .I(n7304), .Z(n275) );
  INV_X2 U10419 ( .I(n19262), .ZN(n1350) );
  NOR2_X1 U5816 ( .A1(n35883), .A2(n21465), .ZN(n4084) );
  INV_X2 U22693 ( .I(n13998), .ZN(n19483) );
  INV_X1 U2199 ( .I(n21713), .ZN(n30731) );
  INV_X2 U23516 ( .I(n15359), .ZN(n16305) );
  INV_X2 U19590 ( .I(n35359), .ZN(n5392) );
  INV_X1 U1538 ( .I(n13996), .ZN(n13959) );
  INV_X1 U24311 ( .I(n14245), .ZN(n14373) );
  INV_X1 U15320 ( .I(n31381), .ZN(n17242) );
  INV_X1 U7304 ( .I(n20810), .ZN(n21492) );
  INV_X1 U10426 ( .I(n694), .ZN(n1353) );
  NAND2_X1 U28217 ( .A1(n19822), .A2(n1372), .ZN(n21393) );
  AOI21_X1 U30656 ( .A1(n17847), .A2(n21839), .B(n452), .ZN(n36930) );
  NOR2_X1 U25067 ( .A1(n21893), .A2(n21568), .ZN(n21569) );
  NAND2_X1 U8658 ( .A1(n19036), .A2(n21702), .ZN(n9425) );
  NOR2_X1 U1477 ( .A1(n19479), .A2(n21775), .ZN(n18742) );
  NOR2_X1 U4639 ( .A1(n21762), .A2(n9642), .ZN(n538) );
  NOR2_X1 U13955 ( .A1(n21894), .A2(n21893), .ZN(n21896) );
  INV_X2 U8686 ( .I(n21840), .ZN(n15031) );
  INV_X2 U6427 ( .I(n19434), .ZN(n21592) );
  INV_X1 U10338 ( .I(n19483), .ZN(n6654) );
  BUF_X2 U4917 ( .I(n21517), .Z(n587) );
  NOR2_X1 U30029 ( .A1(n19375), .A2(n8700), .ZN(n36751) );
  INV_X2 U7855 ( .I(n21751), .ZN(n15910) );
  NAND2_X1 U4933 ( .A1(n21897), .A2(n17242), .ZN(n21838) );
  NAND2_X1 U6413 ( .A1(n21507), .A2(n9670), .ZN(n21591) );
  NAND2_X1 U19081 ( .A1(n19016), .A2(n21432), .ZN(n21825) );
  NOR2_X1 U2655 ( .A1(n21684), .A2(n19262), .ZN(n19403) );
  INV_X1 U1525 ( .I(n9316), .ZN(n21724) );
  NAND2_X1 U8690 ( .A1(n21429), .A2(n14373), .ZN(n13805) );
  INV_X1 U1520 ( .I(n21823), .ZN(n21861) );
  NAND2_X1 U20008 ( .A1(n37111), .A2(n32123), .ZN(n10345) );
  INV_X1 U27635 ( .I(n21655), .ZN(n21779) );
  INV_X2 U1495 ( .I(n10120), .ZN(n1159) );
  NOR2_X1 U21870 ( .A1(n19768), .A2(n21682), .ZN(n21812) );
  INV_X1 U28187 ( .I(n21835), .ZN(n21837) );
  INV_X1 U4918 ( .I(n21849), .ZN(n21667) );
  NOR2_X1 U2814 ( .A1(n21659), .A2(n21660), .ZN(n13257) );
  OAI21_X1 U28206 ( .A1(n21660), .A2(n21767), .B(n21788), .ZN(n21384) );
  NAND2_X1 U19315 ( .A1(n6604), .A2(n33154), .ZN(n21718) );
  INV_X1 U6433 ( .I(n21767), .ZN(n21528) );
  INV_X2 U18302 ( .I(n5392), .ZN(n21914) );
  AND2_X1 U5140 ( .A1(n21492), .A2(n21805), .Z(n683) );
  NAND2_X1 U17280 ( .A1(n20266), .A2(n21478), .ZN(n14946) );
  NOR2_X1 U24732 ( .A1(n19434), .A2(n19238), .ZN(n20587) );
  NAND2_X1 U13950 ( .A1(n21787), .A2(n21528), .ZN(n4829) );
  AOI21_X1 U3245 ( .A1(n14783), .A2(n20277), .B(n15466), .ZN(n14811) );
  NAND2_X1 U29319 ( .A1(n6198), .A2(n31604), .ZN(n21448) );
  NAND2_X1 U16014 ( .A1(n2533), .A2(n21751), .ZN(n15928) );
  INV_X1 U13925 ( .I(n21850), .ZN(n21423) );
  INV_X1 U19078 ( .I(n21825), .ZN(n17866) );
  NAND3_X1 U10283 ( .A1(n15115), .A2(n21727), .A3(n917), .ZN(n14848) );
  NAND2_X1 U17891 ( .A1(n8441), .A2(n21899), .ZN(n8440) );
  NAND2_X1 U8691 ( .A1(n21817), .A2(n2155), .ZN(n2154) );
  NAND2_X1 U28145 ( .A1(n21327), .A2(n21511), .ZN(n21328) );
  AOI21_X1 U13853 ( .A1(n20762), .A2(n19756), .B(n35977), .ZN(n20761) );
  NAND2_X1 U6412 ( .A1(n19470), .A2(n6241), .ZN(n21483) );
  INV_X1 U6411 ( .I(n21924), .ZN(n21469) );
  INV_X1 U7301 ( .I(n20923), .ZN(n21636) );
  INV_X2 U3721 ( .I(n21339), .ZN(n1156) );
  OAI21_X1 U22705 ( .A1(n10915), .A2(n10918), .B(n21804), .ZN(n10914) );
  NOR3_X1 U17011 ( .A1(n19545), .A2(n21806), .A3(n21410), .ZN(n35153) );
  INV_X1 U28971 ( .I(n1847), .ZN(n33413) );
  AOI21_X1 U6037 ( .A1(n4373), .A2(n19133), .B(n16130), .ZN(n16129) );
  NOR2_X1 U10298 ( .A1(n11378), .A2(n21414), .ZN(n21415) );
  NAND2_X1 U26061 ( .A1(n17966), .A2(n39627), .ZN(n15802) );
  CLKBUF_X2 U4649 ( .I(n32617), .Z(n543) );
  NOR2_X1 U28312 ( .A1(n21433), .A2(n18174), .ZN(n36578) );
  NAND2_X1 U4662 ( .A1(n15761), .A2(n13855), .ZN(n17763) );
  NAND2_X1 U27980 ( .A1(n21775), .A2(n19479), .ZN(n21612) );
  NOR2_X1 U28302 ( .A1(n21942), .A2(n21770), .ZN(n21637) );
  NAND2_X1 U28746 ( .A1(n19517), .A2(n21445), .ZN(n2759) );
  INV_X1 U1475 ( .I(n21810), .ZN(n1346) );
  NAND2_X1 U2193 ( .A1(n18174), .A2(n36351), .ZN(n30874) );
  NOR2_X1 U17279 ( .A1(n21478), .A2(n19388), .ZN(n533) );
  INV_X1 U1465 ( .I(n9616), .ZN(n14928) );
  OAI22_X1 U10299 ( .A1(n5047), .A2(n6234), .B1(n21854), .B2(n1156), .ZN(
        n21855) );
  AOI21_X1 U10907 ( .A1(n30874), .A2(n455), .B(n33053), .ZN(n21419) );
  OAI21_X1 U2620 ( .A1(n12927), .A2(n21498), .B(n32164), .ZN(n15125) );
  NAND3_X1 U17562 ( .A1(n35071), .A2(n21789), .A3(n4829), .ZN(n21529) );
  NAND2_X1 U24512 ( .A1(n21779), .A2(n21656), .ZN(n17161) );
  NAND2_X1 U24526 ( .A1(n39426), .A2(n5132), .ZN(n19856) );
  NAND2_X1 U3063 ( .A1(n21644), .A2(n19647), .ZN(n7954) );
  OAI21_X1 U16182 ( .A1(n37155), .A2(n21515), .B(n3670), .ZN(n21516) );
  NOR2_X1 U28165 ( .A1(n18174), .A2(n19609), .ZN(n21342) );
  NOR2_X1 U18894 ( .A1(n14868), .A2(n19392), .ZN(n6102) );
  AOI21_X1 U10326 ( .A1(n21582), .A2(n19699), .B(n21581), .ZN(n21586) );
  NAND2_X1 U10320 ( .A1(n5505), .A2(n5391), .ZN(n5504) );
  AOI21_X1 U10286 ( .A1(n10127), .A2(n8971), .B(n10125), .ZN(n10126) );
  AOI21_X1 U2606 ( .A1(n21448), .A2(n31292), .B(n21672), .ZN(n35737) );
  NAND2_X1 U1486 ( .A1(n9041), .A2(n21492), .ZN(n4296) );
  NOR2_X1 U21448 ( .A1(n12927), .A2(n35651), .ZN(n21797) );
  AOI21_X1 U28277 ( .A1(n32544), .A2(n21509), .B(n33852), .ZN(n21510) );
  NAND2_X1 U10304 ( .A1(n12852), .A2(n15369), .ZN(n2481) );
  AND2_X1 U5141 ( .A1(n16165), .A2(n1766), .Z(n685) );
  NAND2_X1 U16180 ( .A1(n21583), .A2(n3670), .ZN(n21584) );
  AOI21_X1 U3881 ( .A1(n17112), .A2(n38480), .B(n21592), .ZN(n21597) );
  NOR2_X1 U26124 ( .A1(n21497), .A2(n21656), .ZN(n17482) );
  NOR2_X1 U7251 ( .A1(n21836), .A2(n1158), .ZN(n15952) );
  INV_X2 U18740 ( .I(n36425), .ZN(n1680) );
  NAND2_X1 U28278 ( .A1(n21511), .A2(n21510), .ZN(n21512) );
  NOR2_X1 U1478 ( .A1(n4373), .A2(n2645), .ZN(n2644) );
  OAI21_X1 U13936 ( .A1(n21457), .A2(n21456), .B(n19337), .ZN(n13789) );
  INV_X1 U19124 ( .I(n6381), .ZN(n21501) );
  NAND2_X1 U23732 ( .A1(n21648), .A2(n21647), .ZN(n22008) );
  INV_X1 U20711 ( .I(n10820), .ZN(n22221) );
  INV_X1 U5806 ( .I(n22047), .ZN(n22108) );
  NOR2_X1 U17771 ( .A1(n8493), .A2(n22155), .ZN(n4935) );
  INV_X1 U8603 ( .I(n31202), .ZN(n7046) );
  INV_X2 U4647 ( .I(n22100), .ZN(n20391) );
  NOR2_X1 U21068 ( .A1(n33678), .A2(n14196), .ZN(n4765) );
  NAND2_X1 U6540 ( .A1(n22362), .A2(n36397), .ZN(n22358) );
  INV_X1 U13754 ( .I(n2840), .ZN(n14038) );
  INV_X2 U9374 ( .I(n5061), .ZN(n1149) );
  INV_X2 U27208 ( .I(n14423), .ZN(n12230) );
  INV_X1 U30354 ( .I(n38375), .ZN(n10930) );
  BUF_X2 U6292 ( .I(n22243), .Z(n35429) );
  NAND2_X1 U7219 ( .A1(n22040), .A2(n2839), .ZN(n22181) );
  INV_X1 U6020 ( .I(n16880), .ZN(n11091) );
  INV_X1 U13816 ( .I(n22277), .ZN(n22313) );
  NAND2_X1 U10205 ( .A1(n1680), .A2(n16880), .ZN(n7578) );
  INV_X2 U8628 ( .I(n19737), .ZN(n22229) );
  INV_X1 U26324 ( .I(n22130), .ZN(n22189) );
  INV_X1 U10270 ( .I(n17861), .ZN(n17897) );
  INV_X1 U8631 ( .I(n22177), .ZN(n20943) );
  NOR2_X1 U13736 ( .A1(n11044), .A2(n196), .ZN(n8948) );
  INV_X2 U3402 ( .I(n21864), .ZN(n1047) );
  BUF_X2 U4961 ( .I(n8493), .Z(n396) );
  NAND2_X1 U4957 ( .A1(n19471), .A2(n33738), .ZN(n22079) );
  NOR2_X1 U26617 ( .A1(n22358), .A2(n5077), .ZN(n36336) );
  INV_X1 U7224 ( .I(n22353), .ZN(n1678) );
  NOR2_X1 U6533 ( .A1(n1328), .A2(n22196), .ZN(n20758) );
  OAI21_X1 U15455 ( .A1(n31407), .A2(n19655), .B(n17359), .ZN(n22026) );
  NAND3_X1 U26109 ( .A1(n8749), .A2(n21864), .A3(n8439), .ZN(n36680) );
  INV_X1 U1429 ( .I(n2257), .ZN(n6297) );
  CLKBUF_X2 U29244 ( .I(n21864), .Z(n33438) );
  INV_X2 U6435 ( .I(n39075), .ZN(n5232) );
  INV_X1 U2118 ( .I(n22296), .ZN(n13626) );
  INV_X1 U2566 ( .I(n34379), .ZN(n34407) );
  BUF_X2 U26262 ( .I(n474), .Z(n33091) );
  NAND2_X1 U3025 ( .A1(n2840), .A2(n17530), .ZN(n17529) );
  NAND2_X1 U8606 ( .A1(n22267), .A2(n22122), .ZN(n17308) );
  NOR2_X1 U8588 ( .A1(n22190), .A2(n5819), .ZN(n21002) );
  BUF_X2 U22300 ( .I(n22306), .Z(n32478) );
  BUF_X2 U3768 ( .I(n22332), .Z(n30306) );
  INV_X2 U16390 ( .I(n22322), .ZN(n11276) );
  INV_X1 U18729 ( .I(n22222), .ZN(n22017) );
  INV_X1 U1428 ( .I(n22295), .ZN(n22248) );
  NAND2_X1 U5778 ( .A1(n4388), .A2(n22038), .ZN(n3266) );
  INV_X1 U5796 ( .I(n133), .ZN(n1684) );
  NOR2_X1 U17680 ( .A1(n22151), .A2(n35771), .ZN(n15175) );
  INV_X1 U9113 ( .I(n22310), .ZN(n34282) );
  INV_X1 U4443 ( .I(n22058), .ZN(n20234) );
  NAND2_X1 U2619 ( .A1(n10154), .A2(n10930), .ZN(n2127) );
  NOR2_X1 U6530 ( .A1(n19471), .A2(n33086), .ZN(n35014) );
  INV_X1 U2549 ( .I(n22080), .ZN(n35514) );
  NAND2_X1 U25635 ( .A1(n22176), .A2(n20234), .ZN(n4746) );
  NAND2_X1 U13707 ( .A1(n4932), .A2(n17793), .ZN(n8348) );
  NAND2_X1 U21476 ( .A1(n17897), .A2(n20996), .ZN(n35652) );
  NAND2_X1 U13710 ( .A1(n16888), .A2(n22238), .ZN(n21826) );
  NOR2_X1 U19515 ( .A1(n32313), .A2(n35526), .ZN(n6807) );
  OAI21_X1 U17507 ( .A1(n39075), .A2(n6128), .B(n1680), .ZN(n14823) );
  NOR2_X1 U19291 ( .A1(n35618), .A2(n22364), .ZN(n22157) );
  OAI21_X1 U4108 ( .A1(n22313), .A2(n15493), .B(n14925), .ZN(n14924) );
  OAI22_X1 U8587 ( .A1(n1684), .A2(n21972), .B1(n21971), .B2(n1048), .ZN(
        n17027) );
  NAND3_X1 U16812 ( .A1(n8520), .A2(n22197), .A3(n22196), .ZN(n22198) );
  NOR2_X1 U10203 ( .A1(n39075), .A2(n16880), .ZN(n18271) );
  NAND2_X1 U8594 ( .A1(n22323), .A2(n22324), .ZN(n1866) );
  INV_X1 U15126 ( .I(n7355), .ZN(n14181) );
  OAI21_X1 U26683 ( .A1(n19253), .A2(n15499), .B(n11044), .ZN(n9342) );
  AOI21_X1 U13716 ( .A1(n7294), .A2(n16936), .B(n16935), .ZN(n16934) );
  NOR2_X1 U10245 ( .A1(n35429), .A2(n1047), .ZN(n2434) );
  NOR2_X1 U20719 ( .A1(n22143), .A2(n8679), .ZN(n8029) );
  NOR2_X1 U25089 ( .A1(n22236), .A2(n33860), .ZN(n16227) );
  NAND3_X1 U29791 ( .A1(n3266), .A2(n22073), .A3(n3269), .ZN(n3265) );
  NOR2_X1 U16722 ( .A1(n12230), .A2(n4240), .ZN(n22172) );
  NOR2_X1 U13133 ( .A1(n14035), .A2(n14034), .ZN(n22043) );
  NAND2_X1 U7203 ( .A1(n8949), .A2(n22224), .ZN(n8745) );
  INV_X2 U6589 ( .I(n36006), .ZN(n1344) );
  NOR2_X1 U24769 ( .A1(n22017), .A2(n32039), .ZN(n18803) );
  NAND2_X1 U4775 ( .A1(n32408), .A2(n22222), .ZN(n22015) );
  NAND2_X1 U24264 ( .A1(n6127), .A2(n1149), .ZN(n18928) );
  NOR2_X1 U16829 ( .A1(n22101), .A2(n22335), .ZN(n22103) );
  NOR2_X1 U13811 ( .A1(n1342), .A2(n20679), .ZN(n22173) );
  INV_X1 U4032 ( .I(n22194), .ZN(n30996) );
  INV_X1 U1419 ( .I(n20643), .ZN(n22225) );
  NAND2_X1 U2509 ( .A1(n36649), .A2(n36731), .ZN(n502) );
  NOR2_X1 U18038 ( .A1(n22261), .A2(n19471), .ZN(n19975) );
  INV_X1 U24424 ( .I(n22059), .ZN(n15347) );
  BUF_X2 U6556 ( .I(n22058), .Z(n32609) );
  NAND2_X1 U6504 ( .A1(n1047), .A2(n37089), .ZN(n8751) );
  OAI22_X1 U20876 ( .A1(n22006), .A2(n8275), .B1(n22007), .B2(n22225), .ZN(
        n21103) );
  AOI21_X1 U5002 ( .A1(n22065), .A2(n22066), .B(n39151), .ZN(n4479) );
  NOR2_X1 U5000 ( .A1(n22034), .A2(n18854), .ZN(n22037) );
  AOI21_X1 U10175 ( .A1(n11276), .A2(n33091), .B(n31092), .ZN(n17537) );
  OAI21_X1 U17071 ( .A1(n12814), .A2(n36683), .B(n22154), .ZN(n12813) );
  OAI21_X1 U16674 ( .A1(n35755), .A2(n33359), .B(n32478), .ZN(n4198) );
  NOR3_X1 U24545 ( .A1(n22328), .A2(n36303), .A3(n38555), .ZN(n22329) );
  OAI21_X1 U27009 ( .A1(n11276), .A2(n18253), .B(n22324), .ZN(n17782) );
  NAND2_X1 U4406 ( .A1(n13632), .A2(n22146), .ZN(n7911) );
  NOR2_X1 U6381 ( .A1(n14269), .A2(n22134), .ZN(n9391) );
  OAI21_X1 U2083 ( .A1(n22236), .A2(n19261), .B(n33859), .ZN(n20386) );
  AOI21_X1 U10191 ( .A1(n8751), .A2(n8749), .B(n35429), .ZN(n8750) );
  INV_X1 U1443 ( .I(n22254), .ZN(n20308) );
  OAI21_X1 U3515 ( .A1(n8687), .A2(n33438), .B(n19430), .ZN(n13614) );
  OAI21_X1 U2081 ( .A1(n1048), .A2(n32640), .B(n20254), .ZN(n33655) );
  OAI21_X1 U25383 ( .A1(n6724), .A2(n12255), .B(n22281), .ZN(n6723) );
  NAND2_X1 U13695 ( .A1(n15029), .A2(n31649), .ZN(n19654) );
  NOR2_X1 U19954 ( .A1(n584), .A2(n19261), .ZN(n15837) );
  NAND2_X1 U8072 ( .A1(n35754), .A2(n22360), .ZN(n34189) );
  NAND2_X1 U28839 ( .A1(n36616), .A2(n916), .ZN(n2883) );
  NOR2_X1 U23468 ( .A1(n18928), .A2(n22248), .ZN(n12325) );
  OAI21_X1 U19836 ( .A1(n18803), .A2(n18804), .B(n35400), .ZN(n19819) );
  NAND2_X1 U1394 ( .A1(n18429), .A2(n22227), .ZN(n22367) );
  INV_X1 U5586 ( .I(n19815), .ZN(n31771) );
  NAND2_X1 U30434 ( .A1(n15852), .A2(n22272), .ZN(n22499) );
  INV_X1 U30329 ( .I(n22740), .ZN(n33756) );
  NAND2_X1 U26083 ( .A1(n15837), .A2(n20351), .ZN(n15836) );
  OAI21_X1 U10180 ( .A1(n18999), .A2(n36661), .B(n7131), .ZN(n7132) );
  NAND2_X1 U4022 ( .A1(n17782), .A2(n32803), .ZN(n21832) );
  INV_X1 U13606 ( .I(n22651), .ZN(n7530) );
  NOR3_X1 U6373 ( .A1(n3109), .A2(n9485), .A3(n8947), .ZN(n3106) );
  AOI21_X1 U8071 ( .A1(n34189), .A2(n34246), .B(n22361), .ZN(n14800) );
  INV_X1 U28502 ( .I(n29528), .ZN(n27739) );
  INV_X1 U16661 ( .I(n22648), .ZN(n20608) );
  INV_X1 U13614 ( .I(n22542), .ZN(n13236) );
  BUF_X2 U2292 ( .I(n3610), .Z(n2585) );
  INV_X1 U6437 ( .I(n30085), .ZN(n1713) );
  INV_X1 U8738 ( .I(n19407), .ZN(n1375) );
  INV_X1 U1380 ( .I(n29325), .ZN(n1718) );
  INV_X2 U2054 ( .I(n12195), .ZN(n22670) );
  INV_X1 U6441 ( .I(Key[97]), .ZN(n1697) );
  INV_X1 U13639 ( .I(n17756), .ZN(n1664) );
  INV_X1 U8557 ( .I(n22371), .ZN(n22732) );
  INV_X1 U5823 ( .I(n19835), .ZN(n965) );
  INV_X1 U8745 ( .I(n19940), .ZN(n1369) );
  INV_X1 U16168 ( .I(n12818), .ZN(n22482) );
  INV_X1 U14160 ( .I(n1805), .ZN(n7584) );
  INV_X1 U1365 ( .I(n23074), .ZN(n20873) );
  INV_X1 U8537 ( .I(n7584), .ZN(n1320) );
  INV_X2 U18789 ( .I(n5976), .ZN(n14390) );
  INV_X2 U26964 ( .I(n906), .ZN(n23077) );
  INV_X1 U26497 ( .I(n16593), .ZN(n23164) );
  INV_X1 U2401 ( .I(n15289), .ZN(n19307) );
  INV_X1 U26695 ( .I(n33152), .ZN(n14560) );
  AND2_X1 U30835 ( .A1(n407), .A2(n10162), .Z(n22892) );
  BUF_X4 U3735 ( .I(n19680), .Z(n6366) );
  NAND2_X1 U27875 ( .A1(n23188), .A2(n23190), .ZN(n20364) );
  NAND3_X1 U5046 ( .A1(n23078), .A2(n23077), .A3(n33933), .ZN(n23079) );
  NAND2_X1 U24561 ( .A1(n33925), .A2(n22892), .ZN(n20264) );
  NAND2_X1 U25859 ( .A1(n33817), .A2(n22935), .ZN(n17205) );
  INV_X1 U2822 ( .I(n7518), .ZN(n12630) );
  INV_X1 U4281 ( .I(n18220), .ZN(n7960) );
  INV_X1 U13496 ( .I(n20782), .ZN(n13336) );
  CLKBUF_X2 U6626 ( .I(n2047), .Z(n35442) );
  INV_X2 U10056 ( .I(n23060), .ZN(n14765) );
  NOR2_X1 U23680 ( .A1(n301), .A2(n12729), .ZN(n33544) );
  NAND2_X1 U1305 ( .A1(n7266), .A2(n14442), .ZN(n22979) );
  INV_X2 U5997 ( .I(n10436), .ZN(n935) );
  BUF_X2 U4007 ( .I(n22798), .Z(n3273) );
  INV_X2 U1367 ( .I(n20267), .ZN(n936) );
  INV_X1 U6629 ( .I(n36554), .ZN(n34467) );
  INV_X2 U5020 ( .I(n640), .ZN(n23013) );
  INV_X2 U13328 ( .I(n33925), .ZN(n32740) );
  INV_X2 U10061 ( .I(n3452), .ZN(n22919) );
  INV_X1 U7167 ( .I(n22368), .ZN(n20439) );
  INV_X1 U10094 ( .I(n20407), .ZN(n18071) );
  CLKBUF_X2 U29917 ( .I(n10334), .Z(n36736) );
  INV_X2 U1323 ( .I(n23149), .ZN(n9699) );
  INV_X1 U7171 ( .I(n23165), .ZN(n22975) );
  INV_X2 U3183 ( .I(n22795), .ZN(n5380) );
  INV_X1 U28543 ( .I(n23129), .ZN(n22958) );
  INV_X1 U8554 ( .I(n12631), .ZN(n23095) );
  INV_X1 U8497 ( .I(n39527), .ZN(n1318) );
  INV_X1 U7175 ( .I(n550), .ZN(n22859) );
  INV_X1 U23017 ( .I(n11481), .ZN(n20840) );
  AND2_X1 U27279 ( .A1(n217), .A2(n32981), .Z(n23012) );
  INV_X1 U1325 ( .I(n19697), .ZN(n23110) );
  INV_X1 U7169 ( .I(n16174), .ZN(n3906) );
  INV_X2 U2995 ( .I(n8245), .ZN(n1831) );
  NOR2_X1 U5085 ( .A1(n32815), .A2(n22915), .ZN(n22997) );
  NOR2_X1 U2433 ( .A1(n23169), .A2(n23167), .ZN(n17498) );
  NOR3_X1 U15618 ( .A1(n9797), .A2(n23058), .A3(n23060), .ZN(n284) );
  NOR2_X1 U16549 ( .A1(n22804), .A2(n301), .ZN(n14880) );
  NAND2_X1 U20148 ( .A1(n14765), .A2(n23058), .ZN(n32040) );
  OAI21_X1 U21147 ( .A1(n20872), .A2(n23077), .B(n23182), .ZN(n8676) );
  INV_X1 U10065 ( .I(n23047), .ZN(n8720) );
  NOR2_X1 U6616 ( .A1(n2350), .A2(n22900), .ZN(n15199) );
  NAND2_X1 U27432 ( .A1(n19082), .A2(n17131), .ZN(n20373) );
  NOR2_X1 U3302 ( .A1(n2771), .A2(n8942), .ZN(n10296) );
  NOR2_X1 U16752 ( .A1(n35684), .A2(n17205), .ZN(n35791) );
  NAND2_X1 U16335 ( .A1(n14130), .A2(n3803), .ZN(n15741) );
  INV_X1 U13503 ( .I(n9080), .ZN(n11160) );
  INV_X1 U6661 ( .I(n37922), .ZN(n22926) );
  NAND2_X1 U13485 ( .A1(n20590), .A2(n1316), .ZN(n15678) );
  NAND2_X1 U13521 ( .A1(n1315), .A2(n15290), .ZN(n5309) );
  NOR2_X1 U28578 ( .A1(n19697), .A2(n20782), .ZN(n22982) );
  INV_X1 U13463 ( .I(n14804), .ZN(n15041) );
  INV_X1 U1297 ( .I(n15388), .ZN(n5569) );
  BUF_X2 U27230 ( .I(n18415), .Z(n36453) );
  NOR2_X1 U7150 ( .A1(n7960), .A2(n19293), .ZN(n18572) );
  INV_X2 U2297 ( .I(n22920), .ZN(n18518) );
  BUF_X2 U7177 ( .I(n19167), .Z(n19134) );
  INV_X2 U16736 ( .I(n33431), .ZN(n22833) );
  INV_X1 U1330 ( .I(n17691), .ZN(n23177) );
  INV_X1 U7160 ( .I(n33935), .ZN(n19614) );
  CLKBUF_X2 U29294 ( .I(n23101), .Z(n36662) );
  NOR2_X1 U10100 ( .A1(n23095), .A2(n6466), .ZN(n22985) );
  INV_X1 U5770 ( .I(n19840), .ZN(n19440) );
  NAND2_X1 U7136 ( .A1(n1313), .A2(n5581), .ZN(n8705) );
  NOR2_X1 U18429 ( .A1(n4713), .A2(n15045), .ZN(n5555) );
  INV_X1 U10109 ( .I(n39155), .ZN(n1319) );
  OR2_X1 U2406 ( .A1(n4472), .A2(n2880), .Z(n9155) );
  INV_X1 U5531 ( .I(n14395), .ZN(n14725) );
  INV_X1 U5019 ( .I(n9472), .ZN(n1651) );
  INV_X1 U5054 ( .I(n39811), .ZN(n23098) );
  NAND2_X1 U2024 ( .A1(n33972), .A2(n217), .ZN(n5038) );
  NAND2_X1 U10073 ( .A1(n1652), .A2(n17226), .ZN(n10299) );
  NOR2_X1 U13520 ( .A1(n1316), .A2(n22895), .ZN(n16105) );
  AOI21_X1 U21527 ( .A1(n19134), .A2(n19351), .B(n32228), .ZN(n9255) );
  NAND3_X1 U17651 ( .A1(n23028), .A2(n20077), .A3(n15290), .ZN(n17009) );
  AOI22_X1 U18735 ( .A1(n17578), .A2(n23211), .B1(n23209), .B2(n5907), .ZN(
        n18065) );
  AOI21_X1 U14555 ( .A1(n23020), .A2(n22949), .B(n37108), .ZN(n35880) );
  NAND3_X1 U2854 ( .A1(n5380), .A2(n19621), .A3(n59), .ZN(n3628) );
  AOI22_X1 U24269 ( .A1(n18572), .A2(n22915), .B1(n32815), .B2(n22870), .ZN(
        n8013) );
  NAND2_X1 U1990 ( .A1(n35040), .A2(n22880), .ZN(n30599) );
  NOR2_X1 U8488 ( .A1(n1648), .A2(n1316), .ZN(n2795) );
  NAND3_X1 U15062 ( .A1(n6366), .A2(n19614), .A3(n1831), .ZN(n18660) );
  OAI22_X1 U16505 ( .A1(n36736), .A2(n8730), .B1(n4714), .B2(n1144), .ZN(
        n22280) );
  NOR2_X1 U3647 ( .A1(n36453), .A2(n10074), .ZN(n5413) );
  NOR3_X1 U2557 ( .A1(n34014), .A2(n19621), .A3(n34457), .ZN(n11240) );
  AOI21_X1 U7135 ( .A1(n37589), .A2(n36839), .B(n38601), .ZN(n13275) );
  NAND3_X1 U3858 ( .A1(n1146), .A2(n23053), .A3(n14556), .ZN(n13077) );
  NOR2_X1 U15310 ( .A1(n34979), .A2(n22985), .ZN(n10876) );
  NOR2_X1 U30740 ( .A1(n2771), .A2(n15911), .ZN(n2772) );
  NOR2_X1 U6356 ( .A1(n15330), .A2(n23098), .ZN(n7590) );
  NOR3_X1 U28443 ( .A1(n13734), .A2(n18244), .A3(n19788), .ZN(n22397) );
  NAND2_X1 U10101 ( .A1(n23138), .A2(n34368), .ZN(n12618) );
  OAI22_X1 U22906 ( .A1(n18518), .A2(n9725), .B1(n22682), .B2(n22920), .ZN(
        n11301) );
  OAI21_X1 U13514 ( .A1(n1824), .A2(n13734), .B(n36662), .ZN(n23081) );
  AOI22_X1 U26175 ( .A1(n33075), .A2(n33074), .B1(n1824), .B2(n18244), .ZN(
        n3145) );
  NAND3_X1 U2762 ( .A1(n14396), .A2(n19586), .A3(n33745), .ZN(n31748) );
  NAND2_X1 U15585 ( .A1(n35016), .A2(n35918), .ZN(n4611) );
  OAI21_X1 U13298 ( .A1(n34727), .A2(n34726), .B(n39356), .ZN(n7722) );
  NAND2_X1 U20637 ( .A1(n6466), .A2(n6366), .ZN(n7902) );
  NOR2_X1 U2000 ( .A1(n1044), .A2(n19469), .ZN(n32873) );
  NOR2_X1 U8504 ( .A1(n13650), .A2(n39811), .ZN(n2658) );
  NAND3_X1 U22032 ( .A1(n23045), .A2(n15330), .A3(n13650), .ZN(n36903) );
  NAND3_X1 U24034 ( .A1(n18867), .A2(n19181), .A3(n1989), .ZN(n32918) );
  NAND2_X1 U13371 ( .A1(n15041), .A2(n32270), .ZN(n3535) );
  NOR2_X1 U28570 ( .A1(n22949), .A2(n1046), .ZN(n22951) );
  NOR2_X1 U13534 ( .A1(n19966), .A2(n16104), .ZN(n2794) );
  NAND3_X1 U5754 ( .A1(n20637), .A2(n18072), .A3(n22886), .ZN(n18066) );
  NOR2_X1 U4366 ( .A1(n5702), .A2(n39350), .ZN(n6901) );
  NOR2_X1 U24734 ( .A1(n6646), .A2(n20077), .ZN(n19944) );
  INV_X1 U28446 ( .I(n22838), .ZN(n22396) );
  INV_X1 U5089 ( .I(n16967), .ZN(n23031) );
  NOR2_X1 U2395 ( .A1(n23209), .A2(n23135), .ZN(n35806) );
  NOR2_X1 U24549 ( .A1(n15289), .A2(n23028), .ZN(n23171) );
  INV_X2 U30324 ( .I(n2553), .ZN(n36829) );
  NAND2_X1 U26757 ( .A1(n19083), .A2(n20373), .ZN(n23145) );
  NAND2_X1 U5165 ( .A1(n22923), .A2(n5838), .ZN(n5837) );
  OAI21_X1 U13426 ( .A1(n13311), .A2(n23028), .B(n6646), .ZN(n18330) );
  OAI22_X1 U1276 ( .A1(n23197), .A2(n31049), .B1(n23199), .B2(n23198), .ZN(
        n15589) );
  AOI22_X1 U13483 ( .A1(n17226), .A2(n23142), .B1(n5581), .B2(n8508), .ZN(
        n8507) );
  NAND2_X1 U8460 ( .A1(n23012), .A2(n23011), .ZN(n6903) );
  OAI22_X1 U6701 ( .A1(n1045), .A2(n22884), .B1(n20590), .B2(n4340), .ZN(n4704) );
  AOI22_X1 U2356 ( .A1(n2795), .A2(n22895), .B1(n2794), .B2(n20173), .ZN(
        n31657) );
  NAND2_X1 U13461 ( .A1(n23155), .A2(n37674), .ZN(n9700) );
  NOR2_X1 U1282 ( .A1(n23123), .A2(n22876), .ZN(n22878) );
  NAND2_X1 U6692 ( .A1(n5582), .A2(n1652), .ZN(n36527) );
  NAND3_X1 U18811 ( .A1(n8706), .A2(n8705), .A3(n1652), .ZN(n6000) );
  OAI21_X1 U21412 ( .A1(n35851), .A2(n9322), .B(n1141), .ZN(n35644) );
  OAI21_X1 U15119 ( .A1(n23031), .A2(n22954), .B(n18750), .ZN(n6087) );
  OAI21_X1 U16650 ( .A1(n5413), .A2(n4162), .B(n383), .ZN(n4161) );
  NAND2_X1 U17375 ( .A1(n4143), .A2(n9080), .ZN(n7639) );
  INV_X1 U24441 ( .I(n22937), .ZN(n23096) );
  INV_X1 U13524 ( .I(n23156), .ZN(n3561) );
  NAND2_X1 U6349 ( .A1(n16617), .A2(n7130), .ZN(n23432) );
  OAI21_X1 U6348 ( .A1(n10698), .A2(n23114), .B(n1043), .ZN(n10697) );
  NOR2_X1 U1268 ( .A1(n15740), .A2(n15742), .ZN(n6088) );
  NAND2_X1 U7140 ( .A1(n9339), .A2(n9699), .ZN(n9698) );
  NOR2_X1 U13465 ( .A1(n23187), .A2(n14724), .ZN(n4936) );
  OAI21_X1 U5752 ( .A1(n18072), .A2(n18065), .B(n18066), .ZN(n23464) );
  OR2_X1 U6690 ( .A1(n9155), .A2(n17568), .Z(n23511) );
  INV_X1 U6336 ( .I(n17931), .ZN(n12093) );
  INV_X1 U1237 ( .I(n35534), .ZN(n1306) );
  CLKBUF_X2 U2508 ( .I(n23352), .Z(n32158) );
  BUF_X2 U5247 ( .I(n23587), .Z(n19686) );
  BUF_X2 U2293 ( .I(n4644), .Z(n36859) );
  NAND2_X1 U1264 ( .A1(n8569), .A2(n23151), .ZN(n23158) );
  INV_X1 U8435 ( .I(n23303), .ZN(n23488) );
  INV_X1 U5744 ( .I(n7712), .ZN(n12083) );
  INV_X1 U1955 ( .I(n23349), .ZN(n13305) );
  INV_X1 U11695 ( .I(n17508), .ZN(n34558) );
  INV_X1 U5169 ( .I(n23613), .ZN(n14739) );
  INV_X2 U8475 ( .I(n23237), .ZN(n1140) );
  INV_X1 U5261 ( .I(n31908), .ZN(n1290) );
  INV_X2 U6722 ( .I(n35915), .ZN(n4207) );
  NOR2_X1 U2332 ( .A1(n16013), .A2(n23390), .ZN(n23622) );
  NAND2_X1 U9901 ( .A1(n14011), .A2(n23637), .ZN(n7009) );
  INV_X1 U4255 ( .I(n7577), .ZN(n32425) );
  INV_X1 U1239 ( .I(n23461), .ZN(n23370) );
  INV_X1 U6732 ( .I(n35664), .ZN(n1632) );
  INV_X2 U12178 ( .I(n4147), .ZN(n36130) );
  NOR2_X1 U1914 ( .A1(n10839), .A2(n35545), .ZN(n32401) );
  INV_X1 U17322 ( .I(n22493), .ZN(n4542) );
  INV_X1 U8330 ( .I(n18682), .ZN(n1297) );
  INV_X1 U8407 ( .I(n23535), .ZN(n23537) );
  INV_X2 U9963 ( .I(n36539), .ZN(n1300) );
  INV_X1 U1954 ( .I(n10480), .ZN(n52) );
  INV_X2 U13218 ( .I(n7379), .ZN(n23645) );
  NAND2_X1 U6727 ( .A1(n23325), .A2(n35534), .ZN(n23586) );
  NOR2_X1 U2602 ( .A1(n23639), .A2(n7712), .ZN(n10633) );
  NAND2_X1 U3361 ( .A1(n34506), .A2(n23548), .ZN(n13752) );
  INV_X1 U9954 ( .I(n18425), .ZN(n1295) );
  INV_X2 U8453 ( .I(n12028), .ZN(n1310) );
  INV_X1 U5022 ( .I(n23532), .ZN(n1625) );
  INV_X1 U1242 ( .I(n23473), .ZN(n1139) );
  INV_X2 U7197 ( .I(n8668), .ZN(n33496) );
  INV_X2 U4922 ( .I(n36810), .ZN(n23401) );
  INV_X1 U18705 ( .I(n23478), .ZN(n23483) );
  INV_X1 U2319 ( .I(n6159), .ZN(n35367) );
  AND2_X1 U7835 ( .A1(n23423), .A2(n17094), .Z(n34121) );
  AND2_X1 U19428 ( .A1(n39194), .A2(n7225), .Z(n20031) );
  INV_X1 U17353 ( .I(n33840), .ZN(n960) );
  OAI22_X1 U25144 ( .A1(n23483), .A2(n9078), .B1(n23361), .B2(n6176), .ZN(
        n23363) );
  NAND2_X1 U25639 ( .A1(n23526), .A2(n23404), .ZN(n36219) );
  INV_X2 U10227 ( .I(n36564), .ZN(n23270) );
  INV_X1 U13169 ( .I(n23227), .ZN(n23277) );
  NOR2_X1 U8433 ( .A1(n23325), .A2(n19481), .ZN(n23264) );
  NOR2_X1 U9896 ( .A1(n23306), .A2(n23483), .ZN(n8784) );
  NOR2_X1 U28637 ( .A1(n18284), .A2(n35808), .ZN(n23298) );
  NAND2_X1 U13299 ( .A1(n23347), .A2(n14845), .ZN(n5253) );
  NAND2_X1 U8619 ( .A1(n7335), .A2(n3496), .ZN(n23343) );
  AOI22_X1 U6771 ( .A1(n7598), .A2(n4600), .B1(n32226), .B2(n23425), .ZN(
        n18370) );
  NAND2_X1 U20764 ( .A1(n23302), .A2(n37774), .ZN(n32407) );
  NAND2_X1 U13273 ( .A1(n23533), .A2(n23534), .ZN(n16369) );
  NAND2_X1 U7078 ( .A1(n15642), .A2(n35377), .ZN(n2632) );
  CLKBUF_X2 U6345 ( .I(n23461), .Z(n18090) );
  NAND2_X1 U24169 ( .A1(n5591), .A2(n32246), .ZN(n23010) );
  NOR2_X1 U21138 ( .A1(n23453), .A2(n605), .ZN(n9588) );
  INV_X1 U1210 ( .I(n23358), .ZN(n8965) );
  NOR2_X1 U15352 ( .A1(n23306), .A2(n8692), .ZN(n34981) );
  NAND2_X1 U6138 ( .A1(n36027), .A2(n36026), .ZN(n23275) );
  NOR2_X1 U6728 ( .A1(n32425), .A2(n6638), .ZN(n22989) );
  NAND2_X1 U18763 ( .A1(n1644), .A2(n37923), .ZN(n23286) );
  INV_X1 U13266 ( .I(n23534), .ZN(n16086) );
  INV_X1 U13246 ( .I(n23620), .ZN(n13603) );
  NAND2_X1 U9879 ( .A1(n8239), .A2(n10763), .ZN(n10207) );
  BUF_X2 U18870 ( .I(n23567), .Z(n31829) );
  NOR2_X1 U2316 ( .A1(n23251), .A2(n5357), .ZN(n36888) );
  INV_X1 U4740 ( .I(n23572), .ZN(n33721) );
  INV_X2 U5237 ( .I(n2798), .ZN(n31661) );
  NOR2_X1 U15472 ( .A1(n31787), .A2(n35313), .ZN(n35312) );
  INV_X2 U7091 ( .I(n23577), .ZN(n1134) );
  BUF_X2 U2290 ( .I(n36442), .Z(n9835) );
  INV_X1 U11244 ( .I(n23441), .ZN(n11095) );
  INV_X2 U1209 ( .I(n23531), .ZN(n18236) );
  NOR2_X1 U24170 ( .A1(n1631), .A2(n5591), .ZN(n23215) );
  NAND2_X1 U9869 ( .A1(n36564), .A2(n23350), .ZN(n30974) );
  NAND2_X1 U5180 ( .A1(n23572), .A2(n1134), .ZN(n33719) );
  AOI21_X1 U8369 ( .A1(n35039), .A2(n39812), .B(n4396), .ZN(n4251) );
  AOI21_X1 U6763 ( .A1(n23444), .A2(n4207), .B(n36859), .ZN(n23447) );
  NAND3_X1 U8372 ( .A1(n23599), .A2(n23489), .A3(n12597), .ZN(n7825) );
  AOI22_X1 U30624 ( .A1(n8680), .A2(n36885), .B1(n18391), .B2(n33287), .ZN(
        n36945) );
  OAI21_X1 U13193 ( .A1(n22989), .A2(n23256), .B(n1293), .ZN(n17441) );
  NAND3_X1 U22903 ( .A1(n23553), .A2(n14623), .A3(n18236), .ZN(n35864) );
  NOR2_X1 U9855 ( .A1(n23397), .A2(n23264), .ZN(n7630) );
  NOR3_X1 U5255 ( .A1(n30440), .A2(n35001), .A3(n18763), .ZN(n7042) );
  INV_X1 U2258 ( .I(n23526), .ZN(n36878) );
  OAI21_X1 U28271 ( .A1(n2853), .A2(n6637), .B(n6638), .ZN(n36577) );
  OAI21_X1 U24384 ( .A1(n23493), .A2(n23315), .B(n19358), .ZN(n23418) );
  NOR2_X1 U20402 ( .A1(n9192), .A2(n7426), .ZN(n35477) );
  INV_X1 U5217 ( .I(n23476), .ZN(n12009) );
  OAI21_X1 U15286 ( .A1(n20991), .A2(n20992), .B(n16182), .ZN(n31376) );
  INV_X1 U1228 ( .I(n23400), .ZN(n19146) );
  OAI21_X1 U1193 ( .A1(n16086), .A2(n23533), .B(n5184), .ZN(n5183) );
  NAND2_X1 U19184 ( .A1(n39012), .A2(n6217), .ZN(n18237) );
  AOI21_X1 U1835 ( .A1(n23286), .A2(n31091), .B(n33080), .ZN(n31037) );
  OAI21_X1 U19736 ( .A1(n31949), .A2(n16456), .B(n36564), .ZN(n15604) );
  INV_X1 U25123 ( .I(n23581), .ZN(n21297) );
  NAND2_X1 U6764 ( .A1(n23275), .A2(n23274), .ZN(n9889) );
  NAND2_X1 U2665 ( .A1(n5371), .A2(n16370), .ZN(n31074) );
  NAND2_X1 U25848 ( .A1(n12642), .A2(n12641), .ZN(n36241) );
  INV_X1 U9918 ( .I(n23560), .ZN(n17927) );
  NAND2_X1 U15823 ( .A1(n23525), .A2(n3365), .ZN(n3364) );
  NAND2_X1 U13234 ( .A1(n12638), .A2(n1304), .ZN(n23262) );
  NAND2_X1 U5021 ( .A1(n31829), .A2(n32260), .ZN(n4417) );
  INV_X1 U1179 ( .I(n23554), .ZN(n6286) );
  INV_X1 U2151 ( .I(n24012), .ZN(n23659) );
  OAI21_X1 U25150 ( .A1(n18762), .A2(n39133), .B(n18763), .ZN(n16056) );
  OAI22_X1 U8377 ( .A1(n23365), .A2(n3715), .B1(n32260), .B2(n2921), .ZN(n2920) );
  AOI21_X1 U25152 ( .A1(n23278), .A2(n31332), .B(n23277), .ZN(n15562) );
  NAND2_X1 U28591 ( .A1(n39214), .A2(n30524), .ZN(n23038) );
  NAND3_X1 U13215 ( .A1(n18237), .A2(n18235), .A3(n18086), .ZN(n23224) );
  NAND2_X1 U3861 ( .A1(n37279), .A2(n23560), .ZN(n8238) );
  OAI21_X1 U26540 ( .A1(n37923), .A2(n23452), .B(n16713), .ZN(n16712) );
  NAND3_X1 U28594 ( .A1(n23040), .A2(n34386), .A3(n18090), .ZN(n23041) );
  NAND2_X1 U13095 ( .A1(n30364), .A2(n5999), .ZN(n7149) );
  NAND2_X1 U2255 ( .A1(n37005), .A2(n23458), .ZN(n23239) );
  AOI22_X1 U26162 ( .A1(n23640), .A2(n32226), .B1(n1310), .B2(n43), .ZN(n3275)
         );
  INV_X1 U5212 ( .I(n2319), .ZN(n34315) );
  NAND2_X1 U20242 ( .A1(n18680), .A2(n23468), .ZN(n12413) );
  NAND2_X1 U13179 ( .A1(n23579), .A2(n15624), .ZN(n23329) );
  NAND2_X1 U13194 ( .A1(n7425), .A2(n7427), .ZN(n3795) );
  NOR2_X1 U5978 ( .A1(n23054), .A2(n23048), .ZN(n23597) );
  BUF_X2 U6776 ( .I(n9611), .Z(n36895) );
  INV_X1 U1155 ( .I(n23873), .ZN(n2390) );
  INV_X1 U13089 ( .I(n23695), .ZN(n14345) );
  INV_X1 U7811 ( .I(n23900), .ZN(n1620) );
  AOI22_X1 U14958 ( .A1(n18918), .A2(n18917), .B1(n16047), .B2(n23403), .ZN(
        n23712) );
  INV_X1 U1145 ( .I(n23667), .ZN(n1617) );
  INV_X1 U2141 ( .I(n18301), .ZN(n34498) );
  INV_X1 U28056 ( .I(n23655), .ZN(n24005) );
  INV_X1 U1144 ( .I(n17925), .ZN(n23930) );
  INV_X1 U13088 ( .I(n16055), .ZN(n23661) );
  INV_X1 U1829 ( .I(n23778), .ZN(n31227) );
  INV_X1 U3007 ( .I(n9979), .ZN(n12174) );
  INV_X1 U9003 ( .I(n34269), .ZN(n15532) );
  INV_X1 U6324 ( .I(n23671), .ZN(n24024) );
  INV_X1 U6786 ( .I(n24015), .ZN(n3571) );
  BUF_X2 U1131 ( .I(n24463), .Z(n19864) );
  INV_X2 U27146 ( .I(n18178), .ZN(n18402) );
  NAND2_X1 U28803 ( .A1(n17076), .A2(n19864), .ZN(n24134) );
  BUF_X2 U6822 ( .I(n4243), .Z(n33061) );
  NOR2_X1 U12973 ( .A1(n9371), .A2(n17911), .ZN(n9370) );
  BUF_X2 U13052 ( .I(n24164), .Z(n24346) );
  INV_X1 U1077 ( .I(n1609), .ZN(n24478) );
  INV_X1 U1791 ( .I(n24196), .ZN(n31452) );
  NAND2_X1 U6805 ( .A1(n12733), .A2(n24327), .ZN(n24329) );
  CLKBUF_X2 U22682 ( .I(n9520), .Z(n33712) );
  INV_X1 U5033 ( .I(n24169), .ZN(n24398) );
  NAND2_X1 U7039 ( .A1(n24087), .A2(n802), .ZN(n24223) );
  BUF_X2 U12996 ( .I(n24404), .Z(n12360) );
  BUF_X2 U3377 ( .I(n24287), .Z(n232) );
  INV_X2 U5300 ( .I(n6515), .ZN(n24282) );
  BUF_X2 U2206 ( .I(n31403), .Z(n8735) );
  INV_X2 U15201 ( .I(n2741), .ZN(n14392) );
  INV_X1 U6536 ( .I(n16832), .ZN(n1285) );
  INV_X1 U9829 ( .I(n13144), .ZN(n1283) );
  INV_X2 U7941 ( .I(n18402), .ZN(n17066) );
  INV_X1 U15863 ( .I(n15892), .ZN(n18238) );
  INV_X1 U7897 ( .I(n7240), .ZN(n16377) );
  INV_X1 U8342 ( .I(n17709), .ZN(n24143) );
  INV_X1 U23367 ( .I(n12138), .ZN(n19880) );
  INV_X1 U8348 ( .I(n37230), .ZN(n1282) );
  NAND2_X1 U13043 ( .A1(n2192), .A2(n24366), .ZN(n4182) );
  INV_X2 U1767 ( .I(n38886), .ZN(n2336) );
  INV_X1 U18971 ( .I(n6226), .ZN(n21043) );
  INV_X1 U7014 ( .I(n24360), .ZN(n24458) );
  INV_X2 U15853 ( .I(n1129), .ZN(n1031) );
  NOR2_X1 U24247 ( .A1(n1131), .A2(n1275), .ZN(n17163) );
  NOR2_X1 U6830 ( .A1(n37134), .A2(n3226), .ZN(n3228) );
  NAND3_X1 U3711 ( .A1(n21310), .A2(n24461), .A3(n19864), .ZN(n24305) );
  NOR2_X1 U8296 ( .A1(n1595), .A2(n5985), .ZN(n4359) );
  NAND2_X1 U8320 ( .A1(n37045), .A2(n39815), .ZN(n24400) );
  NAND3_X1 U1770 ( .A1(n24390), .A2(n9963), .A3(n13584), .ZN(n30580) );
  NAND2_X1 U4312 ( .A1(n13884), .A2(n10747), .ZN(n12481) );
  INV_X1 U4155 ( .I(n807), .ZN(n17040) );
  INV_X1 U19458 ( .I(n39699), .ZN(n1035) );
  INV_X1 U9811 ( .I(n33599), .ZN(n24283) );
  INV_X2 U5972 ( .I(n19426), .ZN(n20863) );
  NOR2_X1 U4679 ( .A1(n9370), .A2(n24282), .ZN(n32322) );
  INV_X1 U2094 ( .I(n13412), .ZN(n14004) );
  BUF_X2 U4699 ( .I(n24241), .Z(n32360) );
  INV_X1 U8149 ( .I(n39415), .ZN(n34210) );
  INV_X1 U5732 ( .I(n9066), .ZN(n1599) );
  AOI21_X1 U6288 ( .A1(n1586), .A2(n17709), .B(n36757), .ZN(n6215) );
  INV_X1 U12797 ( .I(n24466), .ZN(n12288) );
  NAND2_X1 U12875 ( .A1(n24312), .A2(n24313), .ZN(n12329) );
  CLKBUF_X2 U5193 ( .I(n1609), .Z(n36740) );
  BUF_X2 U9825 ( .I(n18721), .Z(n12146) );
  NOR2_X1 U1044 ( .A1(n914), .A2(n14558), .ZN(n24338) );
  INV_X1 U9788 ( .I(n16366), .ZN(n1594) );
  INV_X1 U19565 ( .I(n18721), .ZN(n24258) );
  INV_X1 U20142 ( .I(n24279), .ZN(n32891) );
  NAND2_X1 U1086 ( .A1(n1032), .A2(n13555), .ZN(n7082) );
  NOR2_X1 U18848 ( .A1(n1129), .A2(n24140), .ZN(n24141) );
  NOR2_X1 U26437 ( .A1(n12733), .A2(n2396), .ZN(n24166) );
  INV_X1 U8347 ( .I(n24287), .ZN(n1602) );
  INV_X1 U8353 ( .I(n35134), .ZN(n1284) );
  OR2_X1 U17515 ( .A1(n10073), .A2(n5211), .Z(n17456) );
  INV_X1 U6312 ( .I(n24116), .ZN(n1274) );
  INV_X1 U2082 ( .I(n16459), .ZN(n33077) );
  INV_X1 U18559 ( .I(n18342), .ZN(n20027) );
  INV_X1 U5973 ( .I(n33939), .ZN(n24295) );
  INV_X1 U20627 ( .I(n17871), .ZN(n7883) );
  AOI21_X1 U9738 ( .A1(n1033), .A2(n24346), .B(n34330), .ZN(n23702) );
  NOR2_X1 U3716 ( .A1(n24134), .A2(n21310), .ZN(n18276) );
  NAND2_X1 U2021 ( .A1(n5953), .A2(n24346), .ZN(n35916) );
  NAND2_X1 U5733 ( .A1(n34547), .A2(n9066), .ZN(n24293) );
  AOI22_X1 U2689 ( .A1(n24231), .A2(n15385), .B1(n1595), .B2(n24335), .ZN(
        n4360) );
  OAI21_X1 U5147 ( .A1(n38302), .A2(n24469), .B(n5599), .ZN(n35504) );
  NOR3_X1 U7023 ( .A1(n1609), .A2(n3869), .A3(n94), .ZN(n15755) );
  NOR2_X1 U26670 ( .A1(n23702), .A2(n23704), .ZN(n36343) );
  NOR2_X1 U1753 ( .A1(n24412), .A2(n24411), .ZN(n4308) );
  INV_X1 U19628 ( .I(n36852), .ZN(n13167) );
  NOR2_X1 U12998 ( .A1(n18116), .A2(n2192), .ZN(n3620) );
  OAI21_X1 U1061 ( .A1(n23820), .A2(n14704), .B(n15018), .ZN(n9846) );
  NOR2_X1 U6847 ( .A1(n8735), .A2(n18920), .ZN(n15872) );
  NOR2_X1 U1036 ( .A1(n19426), .A2(n8193), .ZN(n13350) );
  NAND2_X1 U1066 ( .A1(n17711), .A2(n14378), .ZN(n19026) );
  NOR2_X1 U9787 ( .A1(n35314), .A2(n33061), .ZN(n14899) );
  OAI21_X1 U6286 ( .A1(n24136), .A2(n24267), .B(n19745), .ZN(n24139) );
  NOR2_X1 U15329 ( .A1(n24233), .A2(n23694), .ZN(n15206) );
  NOR2_X1 U3712 ( .A1(n19864), .A2(n21310), .ZN(n12286) );
  OAI21_X1 U25044 ( .A1(n2336), .A2(n7440), .B(n2439), .ZN(n36154) );
  INV_X1 U1742 ( .I(n4475), .ZN(n9909) );
  OAI21_X1 U21215 ( .A1(n11169), .A2(n19864), .B(n19466), .ZN(n32247) );
  OAI21_X1 U21728 ( .A1(n24166), .A2(n24327), .B(n1607), .ZN(n24167) );
  NAND3_X1 U1048 ( .A1(n12367), .A2(n19007), .A3(n7082), .ZN(n7081) );
  OAI21_X1 U10659 ( .A1(n24214), .A2(n18402), .B(n7210), .ZN(n7209) );
  NAND2_X1 U12887 ( .A1(n23844), .A2(n24395), .ZN(n18101) );
  NOR2_X1 U9816 ( .A1(n12771), .A2(n9844), .ZN(n10695) );
  NAND2_X1 U28844 ( .A1(n19415), .A2(n18455), .ZN(n24429) );
  NAND3_X1 U2041 ( .A1(n15145), .A2(n15146), .A3(n24330), .ZN(n36209) );
  NOR2_X1 U9752 ( .A1(n13708), .A2(n1601), .ZN(n13707) );
  AOI22_X1 U15930 ( .A1(n11132), .A2(n24119), .B1(n14684), .B2(n23819), .ZN(
        n11131) );
  NAND2_X1 U9760 ( .A1(n24114), .A2(n12771), .ZN(n7344) );
  NAND2_X1 U23110 ( .A1(n11673), .A2(n24245), .ZN(n21081) );
  INV_X1 U7902 ( .I(n24140), .ZN(n24459) );
  BUF_X2 U4617 ( .I(n16445), .Z(n14705) );
  NOR2_X1 U3392 ( .A1(n1593), .A2(n35244), .ZN(n24165) );
  INV_X1 U7017 ( .I(n1128), .ZN(n1588) );
  INV_X1 U9804 ( .I(n19857), .ZN(n1604) );
  AND2_X1 U7746 ( .A1(n32518), .A2(n9520), .Z(n34080) );
  AOI21_X1 U2969 ( .A1(n13446), .A2(n1032), .B(n13444), .ZN(n13445) );
  AND2_X1 U6062 ( .A1(n18721), .A2(n18269), .Z(n34044) );
  NOR2_X1 U9692 ( .A1(n11317), .A2(n34074), .ZN(n9805) );
  OAI22_X1 U5719 ( .A1(n24293), .A2(n326), .B1(n1599), .B2(n24295), .ZN(n8840)
         );
  NAND2_X1 U24077 ( .A1(n24353), .A2(n24233), .ZN(n13625) );
  AOI21_X1 U19593 ( .A1(n37134), .A2(n24298), .B(n17081), .ZN(n13308) );
  AOI22_X1 U6857 ( .A1(n24149), .A2(n12248), .B1(n20839), .B2(n24207), .ZN(
        n7179) );
  OAI21_X1 U6293 ( .A1(n18698), .A2(n18697), .B(n24274), .ZN(n19537) );
  NAND3_X1 U17821 ( .A1(n37651), .A2(n24407), .A3(n39504), .ZN(n20583) );
  NAND2_X1 U30294 ( .A1(n33727), .A2(n12360), .ZN(n17299) );
  AOI21_X1 U9705 ( .A1(n10220), .A2(n9101), .B(n15049), .ZN(n9888) );
  OAI21_X1 U1969 ( .A1(n2348), .A2(n39478), .B(n36561), .ZN(n16069) );
  OAI21_X1 U1928 ( .A1(n35873), .A2(n35872), .B(n18348), .ZN(n30914) );
  OAI21_X1 U6865 ( .A1(n16829), .A2(n14630), .B(n36378), .ZN(n6953) );
  NAND2_X1 U18916 ( .A1(n39478), .A2(n9963), .ZN(n24391) );
  AOI21_X1 U6850 ( .A1(n19382), .A2(n1127), .B(n24102), .ZN(n30652) );
  NAND2_X1 U1986 ( .A1(n13386), .A2(n36852), .ZN(n9840) );
  NAND2_X1 U28822 ( .A1(n807), .A2(n1601), .ZN(n24265) );
  NOR2_X1 U22345 ( .A1(n24402), .A2(n32484), .ZN(n13741) );
  INV_X1 U6829 ( .I(n24129), .ZN(n3949) );
  AOI21_X1 U23985 ( .A1(n19426), .A2(n38302), .B(n20537), .ZN(n13481) );
  NOR2_X1 U12943 ( .A1(n11758), .A2(n24173), .ZN(n9842) );
  OAI22_X1 U12852 ( .A1(n19381), .A2(n24176), .B1(n24336), .B2(n18295), .ZN(
        n6956) );
  NAND2_X1 U21430 ( .A1(n31270), .A2(n37803), .ZN(n19052) );
  NOR2_X1 U22627 ( .A1(n35815), .A2(n35814), .ZN(n1949) );
  NOR2_X1 U12963 ( .A1(n585), .A2(n32507), .ZN(n34690) );
  NAND2_X1 U19100 ( .A1(n7083), .A2(n7081), .ZN(n6357) );
  NOR2_X1 U14702 ( .A1(n17509), .A2(n24459), .ZN(n34899) );
  AOI21_X1 U21103 ( .A1(n24401), .A2(n8581), .B(n39703), .ZN(n24301) );
  NOR2_X1 U12903 ( .A1(n19682), .A2(n36378), .ZN(n9931) );
  INV_X1 U26358 ( .I(n33108), .ZN(n23765) );
  OAI21_X1 U1759 ( .A1(n24441), .A2(n20903), .B(n19584), .ZN(n33616) );
  OAI22_X1 U20590 ( .A1(n7800), .A2(n24346), .B1(n39156), .B2(n24348), .ZN(
        n12050) );
  NAND2_X1 U19505 ( .A1(n13481), .A2(n19052), .ZN(n35348) );
  OAI21_X1 U10751 ( .A1(n34899), .A2(n35854), .B(n19895), .ZN(n34437) );
  INV_X1 U1672 ( .I(n24746), .ZN(n16196) );
  CLKBUF_X2 U3973 ( .I(n24864), .Z(n32093) );
  CLKBUF_X2 U1643 ( .I(n24661), .Z(n16210) );
  CLKBUF_X2 U1669 ( .I(n3760), .Z(n3487) );
  OAI21_X1 U13510 ( .A1(n13351), .A2(n13350), .B(n5613), .ZN(n31519) );
  INV_X2 U23619 ( .I(n24634), .ZN(n12672) );
  INV_X2 U5704 ( .I(n17986), .ZN(n24630) );
  INV_X2 U6890 ( .I(n15281), .ZN(n934) );
  INV_X2 U4249 ( .I(n9197), .ZN(n457) );
  NAND2_X1 U1844 ( .A1(n12672), .A2(n36634), .ZN(n36690) );
  INV_X1 U4048 ( .I(n19713), .ZN(n24876) );
  INV_X2 U20221 ( .I(n10116), .ZN(n32064) );
  INV_X2 U1886 ( .I(n11081), .ZN(n13495) );
  INV_X1 U14275 ( .I(n13221), .ZN(n24833) );
  INV_X1 U8250 ( .I(n24589), .ZN(n1263) );
  BUF_X2 U21709 ( .I(n17986), .Z(n33012) );
  NAND2_X1 U8144 ( .A1(n37389), .A2(n24589), .ZN(n34199) );
  NAND2_X1 U25924 ( .A1(n24226), .A2(n2747), .ZN(n25018) );
  CLKBUF_X2 U1815 ( .I(n24683), .Z(n33392) );
  NOR2_X1 U15871 ( .A1(n15332), .A2(n24847), .ZN(n36955) );
  INV_X1 U1673 ( .I(n16238), .ZN(n7198) );
  INV_X1 U1897 ( .I(n1265), .ZN(n34198) );
  INV_X2 U6994 ( .I(n5056), .ZN(n24692) );
  NAND2_X1 U12679 ( .A1(n9581), .A2(n9580), .ZN(n9578) );
  INV_X1 U5952 ( .I(n17101), .ZN(n1267) );
  INV_X1 U993 ( .I(n24814), .ZN(n24853) );
  INV_X1 U1629 ( .I(n24686), .ZN(n31712) );
  INV_X1 U8247 ( .I(n7770), .ZN(n36716) );
  INV_X1 U17043 ( .I(n20326), .ZN(n24826) );
  NAND2_X1 U1834 ( .A1(n37983), .A2(n24746), .ZN(n2906) );
  NAND2_X1 U9623 ( .A1(n24572), .A2(n24832), .ZN(n4188) );
  NOR2_X1 U15182 ( .A1(n13045), .A2(n5897), .ZN(n6492) );
  NAND2_X1 U15510 ( .A1(n13966), .A2(n24864), .ZN(n21018) );
  INV_X2 U27302 ( .I(n24883), .ZN(n18845) );
  NOR2_X1 U27540 ( .A1(n16990), .A2(n24737), .ZN(n19278) );
  NOR2_X1 U21937 ( .A1(n24828), .A2(n11081), .ZN(n32403) );
  NOR3_X1 U1583 ( .A1(n1271), .A2(n933), .A3(n7286), .ZN(n32504) );
  NAND3_X1 U5413 ( .A1(n16097), .A2(n32045), .A3(n37411), .ZN(n9209) );
  NAND2_X1 U30055 ( .A1(n24699), .A2(n37097), .ZN(n2608) );
  NAND2_X1 U21025 ( .A1(n24663), .A2(n1029), .ZN(n35579) );
  NOR2_X1 U17431 ( .A1(n19484), .A2(n36376), .ZN(n443) );
  INV_X2 U6878 ( .I(n2340), .ZN(n15137) );
  NAND2_X1 U5944 ( .A1(n36988), .A2(n36340), .ZN(n15427) );
  INV_X1 U28903 ( .I(n37067), .ZN(n24743) );
  NOR2_X1 U28878 ( .A1(n11271), .A2(n24630), .ZN(n24569) );
  NAND3_X1 U3492 ( .A1(n31625), .A2(n23705), .A3(n2018), .ZN(n20975) );
  NAND2_X1 U21043 ( .A1(n30282), .A2(n24691), .ZN(n32223) );
  INV_X2 U977 ( .I(n24877), .ZN(n1119) );
  BUF_X2 U6883 ( .I(n24545), .Z(n34666) );
  INV_X1 U25713 ( .I(n15136), .ZN(n20930) );
  NOR2_X1 U8142 ( .A1(n34199), .A2(n34198), .ZN(n34197) );
  BUF_X4 U1650 ( .I(n33919), .Z(n31161) );
  BUF_X2 U23783 ( .I(n24863), .Z(n35968) );
  BUF_X2 U5375 ( .I(n7506), .Z(n33317) );
  INV_X2 U6282 ( .I(n6977), .ZN(n9212) );
  INV_X1 U1806 ( .I(n36321), .ZN(n35521) );
  CLKBUF_X2 U17710 ( .I(n8966), .Z(n30554) );
  INV_X1 U14264 ( .I(n24698), .ZN(n24900) );
  NAND3_X1 U6908 ( .A1(n24824), .A2(n24821), .A3(n24819), .ZN(n4351) );
  INV_X1 U6893 ( .I(n30534), .ZN(n36920) );
  AND2_X1 U7690 ( .A1(n24250), .A2(n9385), .Z(n34055) );
  INV_X1 U5037 ( .I(n9825), .ZN(n4601) );
  NOR2_X1 U15985 ( .A1(n3510), .A2(n24912), .ZN(n5210) );
  OAI21_X1 U5372 ( .A1(n24789), .A2(n24788), .B(n20039), .ZN(n24510) );
  NAND2_X1 U9654 ( .A1(n957), .A2(n1026), .ZN(n13581) );
  AOI21_X1 U3005 ( .A1(n36988), .A2(n19901), .B(n37477), .ZN(n24651) );
  INV_X1 U12577 ( .I(n12643), .ZN(n1560) );
  AOI22_X1 U1824 ( .A1(n17496), .A2(n24799), .B1(n19679), .B2(n37355), .ZN(
        n34947) );
  NOR2_X1 U9669 ( .A1(n31698), .A2(n31161), .ZN(n4909) );
  NAND3_X1 U22559 ( .A1(n6822), .A2(n5431), .A3(n24828), .ZN(n24571) );
  AOI21_X1 U10989 ( .A1(n2904), .A2(n30699), .B(n37983), .ZN(n2903) );
  NAND2_X1 U3218 ( .A1(n1030), .A2(n35952), .ZN(n24558) );
  NAND2_X1 U3142 ( .A1(n14241), .A2(n36340), .ZN(n33666) );
  OAI21_X1 U12306 ( .A1(n14523), .A2(n18504), .B(n1263), .ZN(n11907) );
  NAND2_X1 U12620 ( .A1(n457), .A2(n9198), .ZN(n11751) );
  NOR2_X1 U24018 ( .A1(n24659), .A2(n19), .ZN(n36046) );
  NAND2_X1 U1756 ( .A1(n16815), .A2(n34906), .ZN(n34747) );
  NAND2_X1 U2626 ( .A1(n6838), .A2(n4323), .ZN(n6574) );
  AOI21_X1 U9617 ( .A1(n6337), .A2(n19484), .B(n9997), .ZN(n10793) );
  AOI21_X1 U24239 ( .A1(n2340), .A2(n24664), .B(n1029), .ZN(n20927) );
  NAND2_X1 U1811 ( .A1(n35579), .A2(n35577), .ZN(n24666) );
  NAND2_X1 U5916 ( .A1(n24177), .A2(n19), .ZN(n35697) );
  NAND2_X1 U2729 ( .A1(n3122), .A2(n24593), .ZN(n62) );
  AOI21_X1 U14779 ( .A1(n32403), .A2(n6822), .B(n9474), .ZN(n34905) );
  NAND2_X1 U12660 ( .A1(n24569), .A2(n37106), .ZN(n13202) );
  INV_X1 U1734 ( .I(n31161), .ZN(n5224) );
  NOR2_X1 U8273 ( .A1(n35968), .A2(n32093), .ZN(n4226) );
  OAI21_X1 U4203 ( .A1(n2731), .A2(n934), .B(n38794), .ZN(n2746) );
  NOR2_X1 U9595 ( .A1(n24965), .A2(n38631), .ZN(n9177) );
  INV_X1 U6261 ( .I(n9021), .ZN(n11642) );
  AND2_X1 U7928 ( .A1(n36321), .A2(n16238), .Z(n34138) );
  NOR2_X1 U23260 ( .A1(n19679), .A2(n31213), .ZN(n11943) );
  AOI21_X1 U19939 ( .A1(n934), .A2(n15282), .B(n12409), .ZN(n12408) );
  AOI21_X1 U15787 ( .A1(n24752), .A2(n1576), .B(n24664), .ZN(n5245) );
  OAI21_X1 U28773 ( .A1(n17658), .A2(n18115), .B(n2731), .ZN(n11769) );
  AOI21_X1 U8229 ( .A1(n24639), .A2(n34906), .B(n14211), .ZN(n2505) );
  AOI22_X1 U1837 ( .A1(n3487), .A2(n11846), .B1(n9921), .B2(n5957), .ZN(n12461) );
  NAND3_X1 U3585 ( .A1(n14241), .A2(n19901), .A3(n38848), .ZN(n15846) );
  NAND3_X1 U25192 ( .A1(n9656), .A2(n958), .A3(n24692), .ZN(n24210) );
  OAI22_X1 U30027 ( .A1(n24728), .A2(n25048), .B1(n12672), .B2(n25053), .ZN(
        n14827) );
  NAND2_X1 U12583 ( .A1(n24629), .A2(n24821), .ZN(n24389) );
  AOI21_X1 U1535 ( .A1(n6957), .A2(n24696), .B(n957), .ZN(n12503) );
  AOI22_X1 U1962 ( .A1(n24644), .A2(n6977), .B1(n32045), .B2(n24643), .ZN(
        n9683) );
  OAI22_X1 U14889 ( .A1(n5653), .A2(n24909), .B1(n25053), .B2(n37105), .ZN(
        n13030) );
  NAND2_X1 U5424 ( .A1(n16841), .A2(n24799), .ZN(n32643) );
  NAND2_X1 U12556 ( .A1(n37210), .A2(n24629), .ZN(n14165) );
  NOR2_X1 U15132 ( .A1(n34138), .A2(n1563), .ZN(n13340) );
  NAND2_X1 U3672 ( .A1(n24736), .A2(n7846), .ZN(n7845) );
  AOI21_X1 U25652 ( .A1(n20158), .A2(n38285), .B(n33317), .ZN(n17343) );
  NAND2_X1 U4581 ( .A1(n8317), .A2(n8318), .ZN(n8316) );
  NAND2_X1 U12590 ( .A1(n24709), .A2(n13050), .ZN(n13049) );
  AOI21_X1 U950 ( .A1(n24556), .A2(n19886), .B(n14532), .ZN(n15586) );
  NAND2_X1 U1775 ( .A1(n6023), .A2(n24691), .ZN(n36918) );
  AOI21_X1 U12991 ( .A1(n6707), .A2(n19484), .B(n6706), .ZN(n4840) );
  NAND2_X1 U28881 ( .A1(n24579), .A2(n24578), .ZN(n24885) );
  NAND2_X1 U1784 ( .A1(n36280), .A2(n7831), .ZN(n10467) );
  AOI21_X1 U2547 ( .A1(n14523), .A2(n37687), .B(n13628), .ZN(n4703) );
  NOR2_X1 U9609 ( .A1(n11943), .A2(n36673), .ZN(n3879) );
  OAI22_X1 U22571 ( .A1(n2340), .A2(n35578), .B1(n38523), .B2(n2341), .ZN(
        n20438) );
  INV_X1 U24255 ( .I(n33271), .ZN(n33197) );
  INV_X1 U12517 ( .I(n24991), .ZN(n5845) );
  INV_X1 U3635 ( .I(n12534), .ZN(n10837) );
  NOR3_X1 U1768 ( .A1(n20411), .A2(n24847), .A3(n11710), .ZN(n12388) );
  NAND2_X1 U6941 ( .A1(n20806), .A2(n19507), .ZN(n20697) );
  OAI22_X1 U18491 ( .A1(n24730), .A2(n39157), .B1(n24731), .B2(n11712), .ZN(
        n35245) );
  BUF_X2 U4561 ( .I(n19725), .Z(n32195) );
  AOI21_X1 U15170 ( .A1(n24531), .A2(n8389), .B(n8388), .ZN(n25229) );
  AOI21_X1 U5693 ( .A1(n24499), .A2(n38369), .B(n12207), .ZN(n12206) );
  INV_X1 U5427 ( .I(n24959), .ZN(n25225) );
  INV_X1 U21794 ( .I(n3015), .ZN(n11756) );
  INV_X1 U896 ( .I(n24994), .ZN(n25083) );
  INV_X1 U8202 ( .I(n25263), .ZN(n5308) );
  INV_X1 U4579 ( .I(n2653), .ZN(n31628) );
  INV_X1 U25184 ( .I(n25160), .ZN(n24676) );
  INV_X1 U9836 ( .I(n16526), .ZN(n7352) );
  NAND2_X1 U15344 ( .A1(n16542), .A2(n9528), .ZN(n25238) );
  INV_X1 U5691 ( .I(n15030), .ZN(n1558) );
  NOR2_X1 U26312 ( .A1(n25022), .A2(n25021), .ZN(n25165) );
  INV_X1 U12586 ( .I(n24985), .ZN(n1561) );
  INV_X1 U6945 ( .I(n24922), .ZN(n25192) );
  INV_X1 U25179 ( .I(n4302), .ZN(n25076) );
  INV_X1 U6943 ( .I(n25247), .ZN(n3647) );
  INV_X1 U22530 ( .I(n24927), .ZN(n16674) );
  NAND2_X1 U16155 ( .A1(n817), .A2(n9181), .ZN(n25202) );
  INV_X1 U6987 ( .I(n24931), .ZN(n4348) );
  INV_X1 U30582 ( .I(n15907), .ZN(n8304) );
  NOR2_X1 U13535 ( .A1(n5100), .A2(n32989), .ZN(n31156) );
  INV_X2 U3139 ( .I(n841), .ZN(n1116) );
  BUF_X2 U9580 ( .I(n14751), .Z(n5798) );
  INV_X1 U5041 ( .I(n34483), .ZN(n9740) );
  INV_X1 U10664 ( .I(n34427), .ZN(n319) );
  INV_X1 U1683 ( .I(n25421), .ZN(n34576) );
  INV_X1 U26453 ( .I(n18121), .ZN(n25574) );
  INV_X1 U876 ( .I(n25581), .ZN(n1253) );
  INV_X1 U8167 ( .I(n18831), .ZN(n19235) );
  NAND2_X1 U25214 ( .A1(n25558), .A2(n25557), .ZN(n17450) );
  INV_X1 U3193 ( .I(n31557), .ZN(n36593) );
  NOR2_X1 U9528 ( .A1(n33826), .A2(n25721), .ZN(n10532) );
  INV_X2 U1613 ( .I(n25540), .ZN(n36991) );
  NAND2_X1 U1639 ( .A1(n12309), .A2(n17594), .ZN(n20888) );
  INV_X1 U3719 ( .I(n33130), .ZN(n9481) );
  INV_X1 U24174 ( .I(n13873), .ZN(n16264) );
  INV_X2 U11620 ( .I(n25606), .ZN(n31359) );
  NAND2_X1 U1748 ( .A1(n8771), .A2(n24963), .ZN(n4625) );
  INV_X1 U19881 ( .I(n12162), .ZN(n7236) );
  CLKBUF_X2 U3788 ( .I(n8069), .Z(n2148) );
  INV_X1 U5458 ( .I(n25647), .ZN(n32279) );
  CLKBUF_X2 U21244 ( .I(n733), .Z(n35611) );
  CLKBUF_X2 U4530 ( .I(n25543), .Z(n517) );
  INV_X2 U27493 ( .I(n19153), .ZN(n25577) );
  INV_X2 U30851 ( .I(n36105), .ZN(n1249) );
  NAND2_X1 U5522 ( .A1(n25665), .A2(n25361), .ZN(n4469) );
  INV_X1 U30171 ( .I(n19941), .ZN(n36792) );
  INV_X2 U9562 ( .I(n24536), .ZN(n19398) );
  INV_X1 U1387 ( .I(n25600), .ZN(n32101) );
  INV_X1 U9568 ( .I(n14473), .ZN(n25401) );
  AND2_X1 U25594 ( .A1(n11060), .A2(n16186), .Z(n16316) );
  INV_X1 U12480 ( .I(n31305), .ZN(n1551) );
  INV_X1 U5942 ( .I(n21042), .ZN(n25670) );
  INV_X1 U9529 ( .I(n33947), .ZN(n7802) );
  INV_X1 U10529 ( .I(n39061), .ZN(n1022) );
  INV_X1 U5683 ( .I(n25696), .ZN(n911) );
  AND2_X1 U23534 ( .A1(n36105), .A2(n25619), .Z(n25142) );
  NAND2_X1 U28861 ( .A1(n25682), .A2(n30633), .ZN(n24535) );
  NAND2_X1 U5843 ( .A1(n32580), .A2(n30377), .ZN(n16372) );
  NAND3_X1 U1363 ( .A1(n25399), .A2(n25400), .A3(n25401), .ZN(n32789) );
  NAND2_X1 U15349 ( .A1(n9526), .A2(n25307), .ZN(n13849) );
  NOR2_X1 U6906 ( .A1(n25487), .A2(n35216), .ZN(n7052) );
  NAND2_X1 U12388 ( .A1(n25603), .A2(n14708), .ZN(n5857) );
  INV_X2 U7926 ( .I(n25513), .ZN(n13461) );
  NOR2_X1 U9488 ( .A1(n9893), .A2(n826), .ZN(n8739) );
  INV_X1 U2037 ( .I(n25484), .ZN(n1547) );
  NAND2_X1 U12402 ( .A1(n12616), .A2(n826), .ZN(n9029) );
  NAND2_X1 U1657 ( .A1(n7705), .A2(n33946), .ZN(n25679) );
  NAND2_X1 U823 ( .A1(n25545), .A2(n1539), .ZN(n13375) );
  AOI21_X1 U27888 ( .A1(n10674), .A2(n19863), .B(n25379), .ZN(n12462) );
  INV_X1 U12428 ( .I(n1252), .ZN(n6064) );
  INV_X2 U870 ( .I(n14081), .ZN(n25642) );
  NOR2_X1 U18245 ( .A1(n4914), .A2(n11060), .ZN(n13468) );
  NAND2_X1 U12316 ( .A1(n25435), .A2(n25248), .ZN(n11441) );
  NAND2_X1 U6249 ( .A1(n16246), .A2(n19696), .ZN(n25698) );
  AOI21_X1 U1286 ( .A1(n15443), .A2(n19095), .B(n31984), .ZN(n31158) );
  OAI21_X1 U9465 ( .A1(n5011), .A2(n5010), .B(n8014), .ZN(n5277) );
  AOI21_X1 U12355 ( .A1(n20440), .A2(n20442), .B(n25361), .ZN(n7339) );
  NOR2_X1 U1275 ( .A1(n14619), .A2(n10530), .ZN(n31159) );
  AOI21_X1 U9517 ( .A1(n7075), .A2(n30694), .B(n37905), .ZN(n7926) );
  INV_X1 U17465 ( .I(n15443), .ZN(n15329) );
  INV_X1 U29571 ( .I(n6592), .ZN(n20855) );
  NAND2_X1 U1581 ( .A1(n19400), .A2(n14410), .ZN(n36907) );
  INV_X1 U4428 ( .I(n138), .ZN(n15406) );
  NAND2_X1 U8112 ( .A1(n12825), .A2(n19581), .ZN(n11278) );
  OR2_X1 U1632 ( .A1(n16203), .A2(n33949), .Z(n4384) );
  AND2_X1 U18573 ( .A1(n25498), .A2(n25380), .Z(n12404) );
  AND2_X1 U3479 ( .A1(n25695), .A2(n25694), .Z(n20105) );
  AND2_X1 U3254 ( .A1(n31669), .A2(n20838), .Z(n25514) );
  INV_X1 U814 ( .I(n34150), .ZN(n19296) );
  INV_X1 U2146 ( .I(n541), .ZN(n15215) );
  INV_X1 U6898 ( .I(n25660), .ZN(n25381) );
  AOI21_X1 U1277 ( .A1(n12394), .A2(n20648), .B(n8014), .ZN(n32255) );
  NAND2_X1 U9451 ( .A1(n4048), .A2(n4664), .ZN(n8907) );
  OAI21_X1 U6899 ( .A1(n10563), .A2(n9915), .B(n9441), .ZN(n9440) );
  NOR2_X1 U1546 ( .A1(n15406), .A2(n36708), .ZN(n36941) );
  NAND2_X1 U1463 ( .A1(n36907), .A2(n1024), .ZN(n21220) );
  OAI21_X1 U19435 ( .A1(n25637), .A2(n6731), .B(n37993), .ZN(n20885) );
  NAND2_X1 U12370 ( .A1(n952), .A2(n15406), .ZN(n8568) );
  NAND2_X1 U6954 ( .A1(n24937), .A2(n14805), .ZN(n31165) );
  INV_X1 U10963 ( .I(n20855), .ZN(n34464) );
  NAND2_X1 U9555 ( .A1(n10882), .A2(n16836), .ZN(n11641) );
  NAND2_X1 U17261 ( .A1(n35449), .A2(n18909), .ZN(n36217) );
  NAND2_X1 U1522 ( .A1(n25625), .A2(n25365), .ZN(n34719) );
  AOI21_X1 U4049 ( .A1(n12382), .A2(n33950), .B(n12500), .ZN(n35117) );
  NAND2_X1 U4496 ( .A1(n31984), .A2(n30705), .ZN(n9427) );
  NAND2_X1 U12335 ( .A1(n1112), .A2(n12500), .ZN(n4642) );
  AOI21_X1 U14381 ( .A1(n36345), .A2(n1984), .B(n7924), .ZN(n34846) );
  OAI21_X1 U30037 ( .A1(n25422), .A2(n18031), .B(n12309), .ZN(n36755) );
  OAI21_X1 U9456 ( .A1(n2416), .A2(n2576), .B(n33785), .ZN(n11547) );
  NOR2_X1 U23541 ( .A1(n12675), .A2(n25754), .ZN(n32684) );
  INV_X1 U30529 ( .I(n25566), .ZN(n33897) );
  NOR2_X1 U24913 ( .A1(n25474), .A2(n36486), .ZN(n16026) );
  INV_X1 U2999 ( .I(n25577), .ZN(n25662) );
  NAND2_X1 U12412 ( .A1(n13016), .A2(n12500), .ZN(n13015) );
  AOI21_X1 U12271 ( .A1(n20746), .A2(n17613), .B(n7802), .ZN(n9803) );
  NOR2_X1 U9495 ( .A1(n11278), .A2(n20052), .ZN(n10719) );
  NOR2_X1 U12415 ( .A1(n25756), .A2(n38338), .ZN(n25627) );
  NOR2_X1 U9772 ( .A1(n31745), .A2(n10034), .ZN(n14794) );
  NAND2_X1 U8944 ( .A1(n32207), .A2(n4214), .ZN(n34264) );
  NOR2_X1 U1254 ( .A1(n10674), .A2(n25660), .ZN(n229) );
  NAND2_X1 U1662 ( .A1(n35882), .A2(n11647), .ZN(n30813) );
  INV_X1 U12411 ( .I(n11363), .ZN(n14316) );
  NOR2_X1 U9501 ( .A1(n15172), .A2(n1108), .ZN(n15924) );
  OAI21_X1 U3093 ( .A1(n36486), .A2(n13461), .B(n13744), .ZN(n25476) );
  NOR2_X1 U3286 ( .A1(n25608), .A2(n25472), .ZN(n17013) );
  INV_X1 U8154 ( .I(n25545), .ZN(n25480) );
  NAND2_X1 U1217 ( .A1(n25195), .A2(n32722), .ZN(n2496) );
  NOR2_X1 U1471 ( .A1(n25682), .A2(n25681), .ZN(n34393) );
  NAND3_X1 U29092 ( .A1(n20856), .A2(n25677), .A3(n14081), .ZN(n25678) );
  NAND2_X1 U12336 ( .A1(n25448), .A2(n39371), .ZN(n14486) );
  OAI21_X1 U15458 ( .A1(n3005), .A2(n591), .B(n38245), .ZN(n3004) );
  OAI21_X1 U22205 ( .A1(n14472), .A2(n32450), .B(n32449), .ZN(n15881) );
  NOR2_X1 U776 ( .A1(n32101), .A2(n3058), .ZN(n3057) );
  INV_X2 U4627 ( .I(n25887), .ZN(n928) );
  NAND3_X1 U18221 ( .A1(n31707), .A2(n12675), .A3(n9441), .ZN(n25755) );
  NOR2_X1 U27394 ( .A1(n33251), .A2(n33250), .ZN(n2248) );
  NAND3_X1 U1405 ( .A1(n34078), .A2(n25562), .A3(n35349), .ZN(n1855) );
  INV_X2 U3802 ( .I(n25345), .ZN(n9530) );
  OAI21_X1 U18873 ( .A1(n10973), .A2(n7987), .B(n6065), .ZN(n10972) );
  NAND2_X1 U8103 ( .A1(n4792), .A2(n4791), .ZN(n25775) );
  AOI21_X1 U1401 ( .A1(n2576), .A2(n25623), .B(n34719), .ZN(n11548) );
  NOR2_X1 U16146 ( .A1(n14613), .A2(n16428), .ZN(n36897) );
  INV_X2 U7069 ( .I(n18062), .ZN(n26016) );
  NAND2_X1 U12228 ( .A1(n11734), .A2(n26128), .ZN(n1827) );
  INV_X2 U16489 ( .I(n25971), .ZN(n1019) );
  INV_X2 U6859 ( .I(n8683), .ZN(n1012) );
  INV_X2 U17864 ( .I(n9412), .ZN(n18406) );
  NOR2_X1 U1314 ( .A1(n26016), .A2(n26015), .ZN(n10850) );
  NAND2_X1 U12234 ( .A1(n15991), .A2(n37184), .ZN(n11952) );
  NAND2_X1 U3948 ( .A1(n31375), .A2(n26020), .ZN(n31312) );
  OAI21_X1 U1396 ( .A1(n954), .A2(n4914), .B(n17353), .ZN(n36624) );
  INV_X2 U7058 ( .I(n17791), .ZN(n26135) );
  BUF_X2 U7741 ( .I(n10223), .Z(n30595) );
  NAND2_X1 U1399 ( .A1(n26019), .A2(n26020), .ZN(n26045) );
  INV_X1 U8051 ( .I(n18176), .ZN(n19793) );
  INV_X1 U764 ( .I(n25993), .ZN(n25957) );
  BUF_X2 U1371 ( .I(n35903), .Z(n31994) );
  INV_X1 U3803 ( .I(n38416), .ZN(n20456) );
  INV_X1 U15898 ( .I(n33879), .ZN(n26185) );
  INV_X1 U6823 ( .I(n25941), .ZN(n26061) );
  INV_X2 U735 ( .I(n10015), .ZN(n5908) );
  INV_X2 U28208 ( .I(n15085), .ZN(n36571) );
  INV_X1 U1333 ( .I(n31362), .ZN(n25998) );
  INV_X2 U7076 ( .I(n37613), .ZN(n11552) );
  NAND2_X1 U1336 ( .A1(n18176), .A2(n25345), .ZN(n25769) );
  NOR2_X1 U1332 ( .A1(n596), .A2(n25941), .ZN(n35720) );
  NOR2_X1 U7077 ( .A1(n3356), .A2(n36226), .ZN(n34382) );
  NAND2_X1 U17766 ( .A1(n26045), .A2(n5886), .ZN(n20088) );
  NOR2_X1 U22033 ( .A1(n25822), .A2(n18142), .ZN(n15832) );
  INV_X1 U722 ( .I(n25798), .ZN(n26004) );
  CLKBUF_X2 U12194 ( .I(n8683), .Z(n9883) );
  NAND2_X1 U24604 ( .A1(n25971), .A2(n18661), .ZN(n26110) );
  CLKBUF_X2 U3068 ( .I(n6830), .Z(n2888) );
  NAND2_X1 U14591 ( .A1(n1017), .A2(n17180), .ZN(n26042) );
  NAND2_X1 U18601 ( .A1(n25770), .A2(n26063), .ZN(n26060) );
  INV_X1 U1978 ( .I(n26001), .ZN(n9379) );
  INV_X1 U17783 ( .I(n26116), .ZN(n31624) );
  INV_X1 U12195 ( .I(n7136), .ZN(n15121) );
  INV_X1 U1186 ( .I(n18827), .ZN(n19259) );
  INV_X2 U5562 ( .I(n39030), .ZN(n26005) );
  INV_X1 U4250 ( .I(n17180), .ZN(n1518) );
  INV_X1 U20294 ( .I(n10834), .ZN(n929) );
  INV_X2 U16575 ( .I(n8375), .ZN(n6056) );
  INV_X1 U17697 ( .I(n13717), .ZN(n9380) );
  INV_X1 U16033 ( .I(n9413), .ZN(n12234) );
  INV_X1 U1303 ( .I(n26329), .ZN(n1240) );
  INV_X1 U730 ( .I(n2349), .ZN(n926) );
  AOI21_X1 U12210 ( .A1(n25975), .A2(n17458), .B(n6056), .ZN(n25793) );
  INV_X2 U1089 ( .I(n6222), .ZN(n33365) );
  NAND3_X1 U1130 ( .A1(n13869), .A2(n38548), .A3(n10724), .ZN(n2418) );
  NOR2_X1 U29127 ( .A1(n25876), .A2(n25875), .ZN(n25877) );
  NAND3_X1 U8718 ( .A1(n38548), .A2(n35003), .A3(n14212), .ZN(n30674) );
  AOI21_X1 U25248 ( .A1(n33263), .A2(n15178), .B(n18884), .ZN(n15177) );
  NAND2_X1 U9378 ( .A1(n14375), .A2(n31263), .ZN(n4293) );
  NOR2_X1 U14581 ( .A1(n8156), .A2(n25738), .ZN(n10510) );
  NOR2_X1 U8041 ( .A1(n6506), .A2(n8683), .ZN(n25760) );
  NOR2_X1 U1248 ( .A1(n32196), .A2(n31340), .ZN(n35046) );
  NOR2_X1 U18574 ( .A1(n25874), .A2(n4322), .ZN(n2891) );
  OAI21_X1 U28982 ( .A1(n25995), .A2(n318), .B(n25111), .ZN(n25110) );
  NAND2_X1 U7086 ( .A1(n11807), .A2(n9883), .ZN(n24917) );
  NAND2_X1 U12102 ( .A1(n10062), .A2(n1102), .ZN(n8710) );
  NAND2_X1 U25238 ( .A1(n25657), .A2(n34402), .ZN(n19214) );
  INV_X1 U12012 ( .I(n26083), .ZN(n11773) );
  INV_X1 U16125 ( .I(n7961), .ZN(n33366) );
  INV_X1 U12244 ( .I(n9694), .ZN(n26032) );
  NOR2_X1 U17284 ( .A1(n30302), .A2(n4163), .ZN(n25788) );
  INV_X1 U4409 ( .I(n35855), .ZN(n1527) );
  BUF_X2 U14965 ( .I(n26054), .Z(n32109) );
  BUF_X2 U18025 ( .I(n1011), .Z(n36722) );
  INV_X1 U12205 ( .I(n19259), .ZN(n2835) );
  INV_X1 U8077 ( .I(n11734), .ZN(n26126) );
  CLKBUF_X2 U4465 ( .I(n6180), .Z(n33795) );
  CLKBUF_X2 U12204 ( .I(n26329), .Z(n7460) );
  NAND2_X1 U1271 ( .A1(n26016), .A2(n26015), .ZN(n26123) );
  NAND2_X1 U14780 ( .A1(n1239), .A2(n586), .ZN(n25745) );
  INV_X1 U4135 ( .I(n26031), .ZN(n1016) );
  INV_X1 U8060 ( .I(n6506), .ZN(n15283) );
  INV_X1 U12243 ( .I(n1107), .ZN(n12711) );
  INV_X1 U10608 ( .I(n26070), .ZN(n15796) );
  INV_X1 U6879 ( .I(n26054), .ZN(n1020) );
  AND2_X1 U5740 ( .A1(n26054), .A2(n2349), .Z(n34153) );
  OAI21_X1 U12106 ( .A1(n25886), .A2(n15796), .B(n928), .ZN(n25858) );
  AOI22_X1 U684 ( .A1(n25862), .A2(n33218), .B1(n38982), .B2(n25861), .ZN(
        n15946) );
  BUF_X2 U7109 ( .I(n25836), .Z(n31954) );
  AOI22_X1 U12162 ( .A1(n33348), .A2(n26050), .B1(n31311), .B2(n1523), .ZN(
        n26051) );
  OAI22_X1 U2568 ( .A1(n32056), .A2(n32690), .B1(n26005), .B2(n26006), .ZN(
        n25531) );
  NAND2_X1 U24608 ( .A1(n20813), .A2(n31340), .ZN(n26213) );
  NAND3_X1 U6201 ( .A1(n10724), .A2(n30937), .A3(n12199), .ZN(n12152) );
  NOR2_X1 U8867 ( .A1(n16200), .A2(n38760), .ZN(n19218) );
  AOI21_X1 U12049 ( .A1(n5326), .A2(n25870), .B(n17501), .ZN(n5325) );
  NAND3_X1 U659 ( .A1(n30900), .A2(n425), .A3(n32052), .ZN(n25406) );
  NAND2_X1 U12145 ( .A1(n25855), .A2(n26004), .ZN(n16612) );
  AOI21_X1 U11034 ( .A1(n25768), .A2(n4832), .B(n1097), .ZN(n21307) );
  AOI22_X1 U14726 ( .A1(n31299), .A2(n9743), .B1(n927), .B2(n949), .ZN(n19368)
         );
  NOR2_X1 U1054 ( .A1(n9568), .A2(n15703), .ZN(n31470) );
  OAI21_X1 U7105 ( .A1(n17502), .A2(n950), .B(n10765), .ZN(n26099) );
  NOR2_X1 U19147 ( .A1(n25771), .A2(n35109), .ZN(n6401) );
  OAI21_X1 U23128 ( .A1(n6578), .A2(n34018), .B(n35891), .ZN(n9087) );
  OAI21_X1 U1190 ( .A1(n34519), .A2(n25996), .B(n11834), .ZN(n11625) );
  NAND3_X1 U18417 ( .A1(n16478), .A2(n16477), .A3(n34265), .ZN(n20507) );
  OAI21_X1 U7934 ( .A1(n32109), .A2(n25745), .B(n30611), .ZN(n25746) );
  NOR2_X1 U7063 ( .A1(n17951), .A2(n14375), .ZN(n26186) );
  NOR3_X1 U17921 ( .A1(n14564), .A2(n31994), .A3(n19898), .ZN(n12709) );
  NAND2_X1 U8717 ( .A1(n30425), .A2(n30674), .ZN(n30934) );
  NAND3_X1 U9375 ( .A1(n25922), .A2(n18038), .A3(n25803), .ZN(n13165) );
  BUF_X2 U5674 ( .I(n26113), .Z(n1521) );
  NAND3_X1 U29111 ( .A1(n26030), .A2(n10062), .A3(n25965), .ZN(n25796) );
  NOR2_X1 U26997 ( .A1(n362), .A2(n25835), .ZN(n18376) );
  NAND2_X1 U18290 ( .A1(n5886), .A2(n38531), .ZN(n5882) );
  OR2_X1 U20853 ( .A1(n14854), .A2(n32185), .Z(n3361) );
  INV_X1 U6158 ( .I(n26215), .ZN(n1529) );
  INV_X1 U6214 ( .I(n8120), .ZN(n26078) );
  INV_X1 U12082 ( .I(n26214), .ZN(n26212) );
  NAND2_X1 U23358 ( .A1(n12721), .A2(n32243), .ZN(n13281) );
  NOR2_X1 U30826 ( .A1(n362), .A2(n18375), .ZN(n5283) );
  OAI21_X1 U18642 ( .A1(n26078), .A2(n26075), .B(n11762), .ZN(n12151) );
  AOI22_X1 U7980 ( .A1(n14685), .A2(n6578), .B1(n6302), .B2(n26061), .ZN(n4430) );
  NAND2_X1 U16375 ( .A1(n35099), .A2(n25977), .ZN(n2574) );
  NAND2_X1 U12120 ( .A1(n25898), .A2(n36293), .ZN(n6396) );
  OAI21_X1 U26613 ( .A1(n36819), .A2(n1015), .B(n36581), .ZN(n25838) );
  AOI22_X1 U1136 ( .A1(n5283), .A2(n1015), .B1(n14694), .B2(n362), .ZN(n34499)
         );
  INV_X1 U27382 ( .I(n25919), .ZN(n18863) );
  INV_X1 U7116 ( .I(n10225), .ZN(n31073) );
  NAND2_X1 U4319 ( .A1(n25831), .A2(n25921), .ZN(n25834) );
  BUF_X2 U640 ( .I(n9858), .Z(n343) );
  OAI21_X1 U5666 ( .A1(n14984), .A2(n25749), .B(n14983), .ZN(n26165) );
  OAI21_X1 U21416 ( .A1(n3361), .A2(n3360), .B(n35646), .ZN(n3781) );
  NAND2_X1 U14570 ( .A1(n9077), .A2(n20116), .ZN(n26530) );
  BUF_X2 U3621 ( .I(n11752), .Z(n291) );
  INV_X1 U6811 ( .I(n6154), .ZN(n16294) );
  NOR2_X1 U17617 ( .A1(n26078), .A2(n9855), .ZN(n2421) );
  NAND2_X1 U1016 ( .A1(n34148), .A2(n18273), .ZN(n7862) );
  INV_X1 U26588 ( .I(n26585), .ZN(n36333) );
  INV_X1 U12005 ( .I(n32095), .ZN(n9870) );
  INV_X1 U1599 ( .I(n17263), .ZN(n8110) );
  INV_X1 U7963 ( .I(n1009), .ZN(n11298) );
  NAND2_X1 U2131 ( .A1(n7603), .A2(n7602), .ZN(n7781) );
  AOI22_X1 U14386 ( .A1(n32747), .A2(n32748), .B1(n26097), .B2(n39351), .ZN(
        n35239) );
  BUF_X2 U15111 ( .I(n4828), .Z(n36958) );
  INV_X1 U20345 ( .I(n34768), .ZN(n35463) );
  INV_X1 U12001 ( .I(n26436), .ZN(n16830) );
  NAND2_X1 U9360 ( .A1(n3100), .A2(n1504), .ZN(n3099) );
  INV_X1 U11976 ( .I(n32464), .ZN(n20843) );
  INV_X1 U623 ( .I(n13062), .ZN(n26729) );
  BUF_X2 U6778 ( .I(n26861), .Z(n8817) );
  BUF_X2 U1082 ( .I(n19423), .Z(n34005) );
  INV_X2 U17785 ( .I(n12682), .ZN(n14380) );
  INV_X2 U16889 ( .I(n13605), .ZN(n26933) );
  INV_X1 U7915 ( .I(n26861), .ZN(n20223) );
  INV_X1 U26192 ( .I(n36292), .ZN(n14453) );
  INV_X1 U1081 ( .I(n740), .ZN(n33858) );
  INV_X1 U11972 ( .I(n37054), .ZN(n1787) );
  INV_X1 U5362 ( .I(n30284), .ZN(n20004) );
  BUF_X2 U962 ( .I(n10355), .Z(n33689) );
  INV_X2 U1034 ( .I(n167), .ZN(n26944) );
  BUF_X2 U7909 ( .I(n11335), .Z(n11334) );
  NAND2_X1 U13250 ( .A1(n19353), .A2(n33561), .ZN(n26987) );
  BUF_X2 U4410 ( .I(n13528), .Z(n33849) );
  CLKBUF_X2 U16312 ( .I(n19615), .Z(n36882) );
  INV_X2 U10744 ( .I(n30853), .ZN(n14355) );
  BUF_X2 U4196 ( .I(n6454), .Z(n441) );
  INV_X2 U5656 ( .I(n26992), .ZN(n26692) );
  INV_X1 U987 ( .I(n39825), .ZN(n17655) );
  INV_X1 U7958 ( .I(n9118), .ZN(n9117) );
  INV_X1 U23229 ( .I(n17252), .ZN(n11864) );
  INV_X1 U18917 ( .I(n26746), .ZN(n20120) );
  INV_X2 U16503 ( .I(n36392), .ZN(n1002) );
  INV_X1 U2899 ( .I(n18210), .ZN(n1008) );
  INV_X1 U30829 ( .I(n17022), .ZN(n26986) );
  INV_X1 U592 ( .I(n34005), .ZN(n26903) );
  INV_X1 U550 ( .I(n10355), .ZN(n1491) );
  INV_X2 U585 ( .I(n8527), .ZN(n26857) );
  NOR3_X1 U3924 ( .A1(n15411), .A2(n17217), .A3(n33726), .ZN(n32849) );
  INV_X1 U22931 ( .I(n34160), .ZN(n14455) );
  INV_X2 U6754 ( .I(n17047), .ZN(n11679) );
  NAND2_X1 U21409 ( .A1(n11138), .A2(n14412), .ZN(n9062) );
  NAND2_X1 U2279 ( .A1(n26920), .A2(n38188), .ZN(n33063) );
  NOR2_X1 U13588 ( .A1(n1497), .A2(n15996), .ZN(n34767) );
  NOR2_X1 U29322 ( .A1(n20399), .A2(n26863), .ZN(n26864) );
  NOR2_X1 U15288 ( .A1(n26943), .A2(n15670), .ZN(n33548) );
  INV_X1 U19191 ( .I(n6454), .ZN(n10479) );
  INV_X1 U7937 ( .I(n35197), .ZN(n26825) );
  INV_X1 U5641 ( .I(n13056), .ZN(n8816) );
  NOR2_X1 U11863 ( .A1(n14488), .A2(n36882), .ZN(n21192) );
  INV_X1 U11807 ( .I(n26950), .ZN(n8815) );
  INV_X1 U934 ( .I(n1003), .ZN(n32344) );
  INV_X1 U887 ( .I(n14065), .ZN(n31225) );
  NOR2_X1 U24812 ( .A1(n1092), .A2(n13757), .ZN(n3961) );
  INV_X2 U6779 ( .I(n14636), .ZN(n26701) );
  INV_X2 U11946 ( .I(n4411), .ZN(n4007) );
  NOR2_X1 U7895 ( .A1(n8814), .A2(n8817), .ZN(n26731) );
  INV_X1 U907 ( .I(n26860), .ZN(n8415) );
  NAND2_X1 U881 ( .A1(n33849), .A2(n37098), .ZN(n31670) );
  INV_X1 U5218 ( .I(n37103), .ZN(n1090) );
  NAND2_X1 U21108 ( .A1(n10355), .A2(n14383), .ZN(n15371) );
  INV_X1 U15211 ( .I(n2752), .ZN(n26800) );
  INV_X2 U1018 ( .I(n858), .ZN(n1490) );
  INV_X1 U24471 ( .I(n26763), .ZN(n26923) );
  INV_X1 U9300 ( .I(n14459), .ZN(n1229) );
  INV_X1 U25629 ( .I(n32986), .ZN(n849) );
  INV_X1 U9341 ( .I(n26770), .ZN(n18903) );
  AOI21_X1 U4546 ( .A1(n5935), .A2(n858), .B(n20423), .ZN(n15998) );
  INV_X1 U553 ( .I(n9618), .ZN(n26740) );
  INV_X1 U23261 ( .I(n11948), .ZN(n17034) );
  INV_X1 U5657 ( .I(n30859), .ZN(n13088) );
  INV_X1 U26505 ( .I(n26795), .ZN(n20699) );
  NAND2_X1 U9336 ( .A1(n3449), .A2(n20399), .ZN(n3919) );
  NOR2_X1 U9301 ( .A1(n31982), .A2(n12682), .ZN(n3742) );
  NAND2_X1 U5690 ( .A1(n11696), .A2(n17515), .ZN(n15650) );
  OAI22_X1 U25401 ( .A1(n31670), .A2(n6891), .B1(n26653), .B2(n37856), .ZN(
        n36655) );
  NAND3_X1 U952 ( .A1(n26828), .A2(n11138), .A3(n17260), .ZN(n36974) );
  NOR3_X1 U4018 ( .A1(n30665), .A2(n26961), .A3(n2292), .ZN(n35403) );
  OAI21_X1 U11850 ( .A1(n14732), .A2(n2491), .B(n13588), .ZN(n12887) );
  NOR2_X1 U7281 ( .A1(n2226), .A2(n32168), .ZN(n4172) );
  NOR2_X1 U11760 ( .A1(n13427), .A2(n37856), .ZN(n7627) );
  OAI21_X1 U6760 ( .A1(n26720), .A2(n1234), .B(n735), .ZN(n13454) );
  OAI21_X1 U16918 ( .A1(n26996), .A2(n14459), .B(n26692), .ZN(n13036) );
  OAI21_X1 U996 ( .A1(n26951), .A2(n31701), .B(n35409), .ZN(n31638) );
  NOR2_X1 U24048 ( .A1(n8478), .A2(n2752), .ZN(n10678) );
  NAND2_X1 U999 ( .A1(n10314), .A2(n5537), .ZN(n36147) );
  NAND2_X1 U19273 ( .A1(n441), .A2(n26639), .ZN(n6555) );
  NAND2_X1 U3006 ( .A1(n8817), .A2(n26780), .ZN(n34426) );
  NAND2_X1 U11964 ( .A1(n26876), .A2(n14455), .ZN(n12328) );
  NAND2_X1 U3054 ( .A1(n26833), .A2(n26724), .ZN(n2882) );
  NAND2_X1 U29193 ( .A1(n26992), .A2(n19364), .ZN(n26284) );
  INV_X2 U2985 ( .I(n862), .ZN(n18809) );
  NAND2_X1 U24637 ( .A1(n33279), .A2(n26970), .ZN(n15196) );
  NOR2_X1 U30654 ( .A1(n36929), .A2(n37055), .ZN(n31277) );
  NAND3_X1 U930 ( .A1(n19939), .A2(n37154), .A3(n11334), .ZN(n32036) );
  NAND2_X1 U7223 ( .A1(n1490), .A2(n5935), .ZN(n15823) );
  AOI21_X1 U19266 ( .A1(n34061), .A2(n11707), .B(n36647), .ZN(n35321) );
  NOR2_X1 U2944 ( .A1(n26857), .A2(n19728), .ZN(n35028) );
  OAI21_X1 U30089 ( .A1(n34108), .A2(n13487), .B(n33396), .ZN(n36769) );
  AOI21_X1 U6691 ( .A1(n32941), .A2(n26679), .B(n36078), .ZN(n30500) );
  NOR2_X1 U17539 ( .A1(n167), .A2(n26614), .ZN(n19206) );
  NAND2_X1 U28379 ( .A1(n14134), .A2(n12220), .ZN(n36582) );
  NAND2_X1 U3357 ( .A1(n1492), .A2(n2140), .ZN(n26976) );
  NOR2_X1 U11884 ( .A1(n852), .A2(n26979), .ZN(n14831) );
  OAI21_X1 U1995 ( .A1(n1088), .A2(n14636), .B(n26700), .ZN(n10441) );
  INV_X2 U15302 ( .I(n38519), .ZN(n8154) );
  NAND2_X1 U21532 ( .A1(n9269), .A2(n19225), .ZN(n26834) );
  OAI21_X1 U23033 ( .A1(n26700), .A2(n14636), .B(n36244), .ZN(n32602) );
  INV_X1 U30553 ( .I(n3574), .ZN(n26663) );
  INV_X1 U7210 ( .I(n7596), .ZN(n26710) );
  INV_X1 U6796 ( .I(n13393), .ZN(n1232) );
  OAI22_X1 U17248 ( .A1(n15650), .A2(n18809), .B1(n10479), .B2(n11696), .ZN(
        n18776) );
  NAND3_X1 U21427 ( .A1(n13801), .A2(n14807), .A3(n1493), .ZN(n9098) );
  OAI21_X1 U9292 ( .A1(n13758), .A2(n26220), .B(n1092), .ZN(n7691) );
  OAI21_X1 U20661 ( .A1(n38852), .A2(n38928), .B(n26772), .ZN(n19172) );
  NAND3_X1 U943 ( .A1(n16686), .A2(n14488), .A3(n36882), .ZN(n26427) );
  AOI21_X1 U24941 ( .A1(n18587), .A2(n19331), .B(n14921), .ZN(n18586) );
  AOI21_X1 U19227 ( .A1(n39824), .A2(n26899), .B(n26898), .ZN(n35311) );
  NOR2_X1 U519 ( .A1(n17574), .A2(n17573), .ZN(n19687) );
  NAND2_X1 U8926 ( .A1(n17097), .A2(n33301), .ZN(n34262) );
  OAI21_X1 U29316 ( .A1(n1091), .A2(n26802), .B(n26801), .ZN(n26806) );
  NAND2_X1 U931 ( .A1(n26877), .A2(n17655), .ZN(n13870) );
  NOR2_X1 U948 ( .A1(n26909), .A2(n9117), .ZN(n26787) );
  NAND2_X1 U9230 ( .A1(n27141), .A2(n946), .ZN(n17916) );
  NAND2_X1 U899 ( .A1(n26653), .A2(n36424), .ZN(n31678) );
  NOR2_X1 U9330 ( .A1(n8155), .A2(n38519), .ZN(n7511) );
  NOR2_X1 U15394 ( .A1(n30347), .A2(n10202), .ZN(n36164) );
  NAND2_X1 U959 ( .A1(n1494), .A2(n37103), .ZN(n26838) );
  NAND3_X1 U22316 ( .A1(n15341), .A2(n14097), .A3(n39117), .ZN(n35772) );
  NAND2_X1 U11809 ( .A1(n8652), .A2(n35537), .ZN(n2129) );
  OAI21_X1 U10293 ( .A1(n36146), .A2(n36147), .B(n34396), .ZN(n32577) );
  NAND3_X1 U26179 ( .A1(n16686), .A2(n26826), .A3(n18903), .ZN(n26425) );
  NOR2_X1 U20765 ( .A1(n33633), .A2(n34034), .ZN(n33631) );
  NAND2_X1 U889 ( .A1(n30665), .A2(n35764), .ZN(n27129) );
  INV_X1 U26321 ( .I(n12756), .ZN(n33097) );
  INV_X1 U7903 ( .I(n26709), .ZN(n18606) );
  INV_X1 U11889 ( .I(n2158), .ZN(n3417) );
  OAI21_X1 U9302 ( .A1(n12373), .A2(n11696), .B(n441), .ZN(n6078) );
  NAND2_X1 U9287 ( .A1(n948), .A2(n26696), .ZN(n10340) );
  OAI21_X1 U5898 ( .A1(n9147), .A2(n4946), .B(n36873), .ZN(n12936) );
  AOI21_X1 U9239 ( .A1(n32633), .A2(n32634), .B(n1492), .ZN(n17143) );
  AOI21_X1 U15746 ( .A1(n3283), .A2(n19449), .B(n3282), .ZN(n27283) );
  NAND2_X1 U17875 ( .A1(n26650), .A2(n18719), .ZN(n18718) );
  NAND2_X1 U7269 ( .A1(n20636), .A2(n1090), .ZN(n14757) );
  NOR2_X1 U1762 ( .A1(n1232), .A2(n3606), .ZN(n12714) );
  OAI21_X1 U23458 ( .A1(n30363), .A2(n32669), .B(n13392), .ZN(n20792) );
  INV_X1 U7288 ( .I(n32926), .ZN(n2660) );
  OAI22_X1 U862 ( .A1(n32693), .A2(n34004), .B1(n8465), .B2(n1002), .ZN(n35573) );
  NAND3_X1 U2039 ( .A1(n26564), .A2(n17194), .A3(n26636), .ZN(n26637) );
  NAND3_X1 U4073 ( .A1(n26750), .A2(n17194), .A3(n15897), .ZN(n15896) );
  NAND2_X1 U890 ( .A1(n21182), .A2(n36445), .ZN(n21050) );
  NOR2_X1 U29844 ( .A1(n19529), .A2(n27508), .ZN(n27420) );
  INV_X1 U750 ( .I(n27361), .ZN(n27282) );
  INV_X1 U4680 ( .I(n17132), .ZN(n13333) );
  INV_X1 U21544 ( .I(n36833), .ZN(n30290) );
  INV_X2 U484 ( .I(n12485), .ZN(n17142) );
  BUF_X2 U806 ( .I(n27361), .Z(n32557) );
  INV_X1 U19721 ( .I(n39424), .ZN(n35381) );
  INV_X2 U17978 ( .I(n11910), .ZN(n20671) );
  INV_X1 U4474 ( .I(n7973), .ZN(n1480) );
  INV_X2 U24262 ( .I(n34644), .ZN(n27081) );
  INV_X1 U3188 ( .I(n35051), .ZN(n11736) );
  INV_X2 U793 ( .I(n15360), .ZN(n31298) );
  INV_X2 U5880 ( .I(n35500), .ZN(n12326) );
  INV_X2 U15027 ( .I(n39826), .ZN(n14327) );
  CLKBUF_X2 U4153 ( .I(n5363), .Z(n11765) );
  INV_X1 U5700 ( .I(n3540), .ZN(n995) );
  INV_X2 U28310 ( .I(n27448), .ZN(n16043) );
  INV_X2 U8081 ( .I(n11729), .ZN(n27180) );
  INV_X2 U5891 ( .I(n7632), .ZN(n1000) );
  INV_X1 U30562 ( .I(n27358), .ZN(n1227) );
  INV_X1 U19112 ( .I(n19135), .ZN(n35299) );
  INV_X1 U5381 ( .I(n27365), .ZN(n5772) );
  INV_X2 U5581 ( .I(n30358), .ZN(n10946) );
  NAND2_X1 U2881 ( .A1(n27415), .A2(n30434), .ZN(n33234) );
  OAI21_X1 U23988 ( .A1(n27372), .A2(n38578), .B(n16042), .ZN(n16041) );
  NAND3_X1 U9157 ( .A1(n13294), .A2(n6534), .A3(n27240), .ZN(n8263) );
  NOR2_X1 U17558 ( .A1(n27341), .A2(n7096), .ZN(n27342) );
  NAND2_X1 U7782 ( .A1(n36528), .A2(n4192), .ZN(n16849) );
  NAND2_X1 U18665 ( .A1(n36989), .A2(n27379), .ZN(n6446) );
  INV_X1 U27384 ( .I(n20740), .ZN(n27147) );
  BUF_X2 U9706 ( .I(n19529), .Z(n30768) );
  INV_X1 U3576 ( .I(n8537), .ZN(n16263) );
  NAND2_X1 U29390 ( .A1(n39414), .A2(n27240), .ZN(n27238) );
  INV_X2 U19794 ( .I(n27269), .ZN(n19662) );
  NAND2_X1 U29382 ( .A1(n12326), .A2(n38060), .ZN(n27206) );
  NAND2_X1 U17192 ( .A1(n1225), .A2(n7096), .ZN(n4037) );
  NOR3_X1 U21123 ( .A1(n17467), .A2(n20574), .A3(n8627), .ZN(n27092) );
  NAND2_X1 U16275 ( .A1(n13526), .A2(n20377), .ZN(n12375) );
  NAND2_X1 U4654 ( .A1(n27108), .A2(n6686), .ZN(n27181) );
  INV_X2 U18865 ( .I(n993), .ZN(n33146) );
  NAND3_X1 U18483 ( .A1(n1000), .A2(n31298), .A3(n27357), .ZN(n15429) );
  INV_X1 U6588 ( .I(n20133), .ZN(n9512) );
  INV_X1 U479 ( .I(n27424), .ZN(n3059) );
  INV_X1 U16313 ( .I(n7975), .ZN(n27247) );
  NAND2_X1 U7344 ( .A1(n27275), .A2(n27314), .ZN(n6648) );
  INV_X1 U788 ( .I(n18743), .ZN(n7706) );
  INV_X1 U507 ( .I(n15616), .ZN(n1080) );
  INV_X1 U746 ( .I(n4034), .ZN(n1224) );
  INV_X1 U18683 ( .I(n39583), .ZN(n1481) );
  NAND2_X1 U18369 ( .A1(n6191), .A2(n27292), .ZN(n27295) );
  NOR2_X1 U728 ( .A1(n38578), .A2(n19662), .ZN(n3470) );
  NAND2_X1 U3486 ( .A1(n27251), .A2(n35184), .ZN(n2377) );
  AOI21_X1 U6143 ( .A1(n16170), .A2(n19997), .B(n1477), .ZN(n8640) );
  OAI21_X1 U9182 ( .A1(n38630), .A2(n27409), .B(n10677), .ZN(n4570) );
  AOI21_X1 U30226 ( .A1(n27250), .A2(n27007), .B(n27027), .ZN(n36806) );
  NOR3_X1 U30081 ( .A1(n11765), .A2(n15276), .A3(n33893), .ZN(n36761) );
  NAND3_X1 U6155 ( .A1(n37653), .A2(n13278), .A3(n35485), .ZN(n17500) );
  NOR2_X1 U9191 ( .A1(n2761), .A2(n39826), .ZN(n2580) );
  NAND2_X1 U22453 ( .A1(n2035), .A2(n27402), .ZN(n3978) );
  NOR2_X1 U18444 ( .A1(n38926), .A2(n2923), .ZN(n14634) );
  INV_X1 U11604 ( .I(n27299), .ZN(n27377) );
  NAND2_X1 U656 ( .A1(n27297), .A2(n27225), .ZN(n31273) );
  NOR2_X1 U686 ( .A1(n1475), .A2(n27269), .ZN(n34990) );
  INV_X1 U5743 ( .I(n10032), .ZN(n17903) );
  INV_X1 U663 ( .I(n27245), .ZN(n33619) );
  NAND2_X1 U24248 ( .A1(n14086), .A2(n8385), .ZN(n14085) );
  NAND2_X1 U799 ( .A1(n27398), .A2(n17142), .ZN(n32631) );
  NAND3_X1 U13451 ( .A1(n31150), .A2(n11140), .A3(n15360), .ZN(n15120) );
  NAND2_X1 U28843 ( .A1(n13178), .A2(n33403), .ZN(n11591) );
  NOR2_X1 U9148 ( .A1(n12074), .A2(n27090), .ZN(n12073) );
  CLKBUF_X2 U18648 ( .I(n27407), .Z(n7606) );
  NAND2_X1 U2378 ( .A1(n31298), .A2(n34952), .ZN(n27360) );
  NAND2_X1 U14328 ( .A1(n16849), .A2(n16847), .ZN(n16848) );
  NOR2_X1 U29275 ( .A1(n37598), .A2(n36203), .ZN(n26623) );
  BUF_X2 U30772 ( .I(n495), .Z(n37001) );
  NOR2_X1 U11529 ( .A1(n1220), .A2(n1797), .ZN(n1796) );
  NOR2_X1 U687 ( .A1(n17754), .A2(n945), .ZN(n36120) );
  INV_X1 U14209 ( .I(n27408), .ZN(n27155) );
  INV_X1 U19128 ( .I(n27347), .ZN(n11682) );
  INV_X1 U7347 ( .I(n36989), .ZN(n27072) );
  OAI22_X1 U705 ( .A1(n4037), .A2(n8486), .B1(n27133), .B2(n1225), .ZN(n36467)
         );
  NAND2_X1 U14448 ( .A1(n15360), .A2(n27357), .ZN(n2207) );
  INV_X1 U721 ( .I(n495), .ZN(n27154) );
  AOI22_X1 U9144 ( .A1(n30429), .A2(n11682), .B1(n993), .B2(n27348), .ZN(
        n18075) );
  NAND3_X1 U29365 ( .A1(n1486), .A2(n27196), .A3(n27364), .ZN(n27122) );
  NAND3_X1 U29405 ( .A1(n27371), .A2(n1475), .A3(n944), .ZN(n27376) );
  AOI21_X1 U2446 ( .A1(n1472), .A2(n27447), .B(n32926), .ZN(n1940) );
  AOI21_X1 U6148 ( .A1(n8453), .A2(n27403), .B(n35258), .ZN(n15464) );
  NAND3_X1 U434 ( .A1(n1217), .A2(n1224), .A3(n3513), .ZN(n27382) );
  NAND3_X1 U29375 ( .A1(n18246), .A2(n1085), .A3(n27416), .ZN(n27182) );
  AOI21_X1 U3111 ( .A1(n30851), .A2(n33254), .B(n27081), .ZN(n10337) );
  AOI22_X1 U5773 ( .A1(n38146), .A2(n27403), .B1(n33803), .B2(n994), .ZN(
        n32184) );
  AOI22_X1 U24245 ( .A1(n36865), .A2(n27404), .B1(n27390), .B2(n13730), .ZN(
        n2998) );
  OAI21_X1 U6703 ( .A1(n27560), .A2(n1082), .B(n10508), .ZN(n27078) );
  NAND2_X1 U16550 ( .A1(n35115), .A2(n35114), .ZN(n35113) );
  NAND3_X1 U1653 ( .A1(n37198), .A2(n39203), .A3(n27154), .ZN(n27083) );
  NAND2_X1 U21956 ( .A1(n10359), .A2(n13364), .ZN(n10358) );
  NAND2_X1 U11551 ( .A1(n27329), .A2(n27328), .ZN(n21164) );
  AOI21_X1 U628 ( .A1(n27245), .A2(n4192), .B(n2006), .ZN(n2114) );
  NOR2_X1 U4898 ( .A1(n34606), .A2(n4782), .ZN(n8933) );
  NAND2_X1 U18422 ( .A1(n17903), .A2(n27284), .ZN(n17902) );
  NAND2_X1 U22390 ( .A1(n16248), .A2(n4743), .ZN(n35790) );
  NAND2_X1 U21642 ( .A1(n27319), .A2(n37508), .ZN(n9491) );
  OAI21_X1 U9174 ( .A1(n18768), .A2(n2580), .B(n27291), .ZN(n18767) );
  NAND2_X1 U1988 ( .A1(n10066), .A2(n18268), .ZN(n19803) );
  NOR2_X1 U25260 ( .A1(n1217), .A2(n27072), .ZN(n19062) );
  NAND2_X1 U11577 ( .A1(n37162), .A2(n7291), .ZN(n20561) );
  OAI21_X1 U14203 ( .A1(n27155), .A2(n5311), .B(n37001), .ZN(n3674) );
  AOI21_X1 U4479 ( .A1(n27006), .A2(n7973), .B(n32976), .ZN(n5769) );
  NAND2_X1 U15066 ( .A1(n34944), .A2(n34943), .ZN(n35293) );
  NAND2_X1 U4307 ( .A1(n33088), .A2(n31668), .ZN(n27258) );
  NOR2_X1 U20969 ( .A1(n7494), .A2(n39448), .ZN(n13895) );
  NAND2_X1 U2810 ( .A1(n36797), .A2(n19203), .ZN(n35423) );
  INV_X1 U392 ( .I(n27852), .ZN(n1458) );
  OAI21_X1 U11506 ( .A1(n27065), .A2(n26273), .B(n1221), .ZN(n6027) );
  NAND3_X1 U19471 ( .A1(n20740), .A2(n36234), .A3(n945), .ZN(n27148) );
  NAND2_X1 U11543 ( .A1(n7694), .A2(n17058), .ZN(n10953) );
  NAND2_X1 U22752 ( .A1(n37162), .A2(n38305), .ZN(n10999) );
  INV_X1 U3053 ( .I(n37881), .ZN(n4709) );
  INV_X1 U3535 ( .I(n27834), .ZN(n32160) );
  OAI21_X1 U25272 ( .A1(n14482), .A2(n15986), .B(n17754), .ZN(n15985) );
  INV_X1 U381 ( .I(n27554), .ZN(n27853) );
  INV_X1 U17733 ( .I(n8894), .ZN(n33595) );
  OAI21_X1 U18800 ( .A1(n11486), .A2(n14667), .B(n26196), .ZN(n27794) );
  BUF_X2 U16663 ( .I(n19606), .Z(n32931) );
  BUF_X2 U19263 ( .I(n10301), .Z(n35318) );
  INV_X1 U10104 ( .I(n27464), .ZN(n27669) );
  INV_X1 U5835 ( .I(n27672), .ZN(n27849) );
  INV_X1 U11447 ( .I(n27756), .ZN(n16972) );
  INV_X1 U5810 ( .I(n27760), .ZN(n9162) );
  INV_X1 U6697 ( .I(n14260), .ZN(n27676) );
  NAND2_X1 U17329 ( .A1(n36639), .A2(n35603), .ZN(n35178) );
  INV_X1 U6696 ( .I(n27607), .ZN(n27460) );
  INV_X1 U7750 ( .I(n17417), .ZN(n17418) );
  INV_X1 U5829 ( .I(n27830), .ZN(n1456) );
  BUF_X2 U5524 ( .I(n28204), .Z(n9514) );
  INV_X2 U557 ( .I(n10817), .ZN(n7528) );
  INV_X1 U12018 ( .I(n34594), .ZN(n12218) );
  INV_X1 U5860 ( .I(n759), .ZN(n1441) );
  INV_X2 U3907 ( .I(n5352), .ZN(n1442) );
  AOI21_X1 U13947 ( .A1(n1212), .A2(n15357), .B(n32783), .ZN(n15204) );
  INV_X2 U497 ( .I(n19750), .ZN(n1451) );
  INV_X1 U24082 ( .I(n13989), .ZN(n15038) );
  INV_X1 U343 ( .I(n8148), .ZN(n8149) );
  INV_X1 U27296 ( .I(n36463), .ZN(n879) );
  NOR2_X1 U340 ( .A1(n1202), .A2(n15704), .ZN(n10779) );
  NOR2_X1 U19758 ( .A1(n1209), .A2(n8078), .ZN(n11737) );
  NAND2_X1 U2914 ( .A1(n1439), .A2(n28205), .ZN(n16261) );
  INV_X1 U4134 ( .I(n17314), .ZN(n28102) );
  BUF_X2 U21722 ( .I(n28237), .Z(n32352) );
  INV_X1 U6648 ( .I(n877), .ZN(n28156) );
  INV_X2 U26373 ( .I(n28279), .ZN(n1076) );
  INV_X1 U543 ( .I(n12673), .ZN(n5020) );
  AND2_X1 U9665 ( .A1(n34166), .A2(n35225), .Z(n28064) );
  INV_X1 U29356 ( .I(n27481), .ZN(n28050) );
  INV_X1 U6650 ( .I(n7528), .ZN(n27980) );
  INV_X1 U23243 ( .I(n32638), .ZN(n13081) );
  INV_X1 U593 ( .I(n28133), .ZN(n28015) );
  NOR2_X1 U28028 ( .A1(n33603), .A2(n879), .ZN(n20941) );
  NAND3_X1 U6644 ( .A1(n18673), .A2(n13769), .A3(n15704), .ZN(n7717) );
  NAND2_X1 U584 ( .A1(n19410), .A2(n19667), .ZN(n345) );
  NAND2_X1 U461 ( .A1(n20053), .A2(n15925), .ZN(n27940) );
  NOR2_X1 U514 ( .A1(n4915), .A2(n2717), .ZN(n36818) );
  INV_X1 U334 ( .I(n878), .ZN(n28001) );
  INV_X1 U515 ( .I(n12038), .ZN(n32728) );
  AOI21_X1 U7467 ( .A1(n12784), .A2(n28283), .B(n16544), .ZN(n30565) );
  BUF_X2 U2678 ( .I(n18261), .Z(n42) );
  NOR2_X1 U522 ( .A1(n983), .A2(n10836), .ZN(n10519) );
  CLKBUF_X2 U572 ( .I(n5352), .Z(n35607) );
  BUF_X2 U2333 ( .I(n15692), .Z(n9897) );
  NOR2_X1 U6677 ( .A1(n883), .A2(n20860), .ZN(n20977) );
  INV_X2 U510 ( .I(n28024), .ZN(n33331) );
  INV_X2 U17028 ( .I(n8818), .ZN(n28109) );
  INV_X2 U20871 ( .I(n27894), .ZN(n28165) );
  INV_X1 U2501 ( .I(n9534), .ZN(n11754) );
  OR2_X1 U15417 ( .A1(n15922), .A2(n28159), .Z(n11501) );
  AND2_X1 U8017 ( .A1(n19891), .A2(n19605), .Z(n34170) );
  AND2_X1 U11342 ( .A1(n20010), .A2(n19995), .Z(n15623) );
  INV_X1 U549 ( .I(n37056), .ZN(n28151) );
  INV_X1 U9111 ( .I(n28157), .ZN(n28012) );
  INV_X1 U322 ( .I(n886), .ZN(n1205) );
  INV_X2 U7713 ( .I(n18261), .ZN(n1444) );
  INV_X1 U6684 ( .I(n14451), .ZN(n28230) );
  INV_X2 U15061 ( .I(n5988), .ZN(n7690) );
  INV_X2 U18125 ( .I(n2716), .ZN(n1440) );
  OAI21_X1 U3455 ( .A1(n1070), .A2(n28215), .B(n1448), .ZN(n28081) );
  NAND3_X1 U20416 ( .A1(n8232), .A2(n28229), .A3(n28228), .ZN(n19921) );
  NAND2_X1 U9755 ( .A1(n3983), .A2(n30773), .ZN(n15622) );
  NAND2_X1 U20545 ( .A1(n3032), .A2(n3159), .ZN(n35507) );
  AOI21_X1 U16253 ( .A1(n11375), .A2(n32080), .B(n28159), .ZN(n5671) );
  NOR2_X1 U3665 ( .A1(n37057), .A2(n988), .ZN(n13469) );
  INV_X1 U13223 ( .I(n889), .ZN(n7310) );
  AOI21_X1 U27952 ( .A1(n11754), .A2(n27948), .B(n33331), .ZN(n10352) );
  INV_X1 U30038 ( .I(n28043), .ZN(n2664) );
  NAND2_X1 U26487 ( .A1(n18603), .A2(n15357), .ZN(n15518) );
  NOR2_X1 U3216 ( .A1(n11628), .A2(n28272), .ZN(n13776) );
  NAND2_X1 U11331 ( .A1(n18392), .A2(n12260), .ZN(n12258) );
  NAND2_X1 U25824 ( .A1(n36818), .A2(n36817), .ZN(n16034) );
  INV_X2 U11360 ( .I(n1074), .ZN(n19124) );
  NAND2_X1 U3931 ( .A1(n19366), .A2(n99), .ZN(n28053) );
  NOR2_X1 U27193 ( .A1(n1207), .A2(n28290), .ZN(n28291) );
  INV_X1 U7729 ( .I(n9089), .ZN(n21020) );
  OAI21_X1 U9058 ( .A1(n6050), .A2(n5239), .B(n35607), .ZN(n13695) );
  INV_X1 U7702 ( .I(n30484), .ZN(n1435) );
  INV_X1 U30818 ( .I(n8604), .ZN(n28266) );
  INV_X1 U6135 ( .I(n38579), .ZN(n28217) );
  INV_X1 U501 ( .I(n1454), .ZN(n1073) );
  NOR2_X1 U14558 ( .A1(n9969), .A2(n28189), .ZN(n28190) );
  NAND2_X1 U482 ( .A1(n28215), .A2(n987), .ZN(n16971) );
  NOR2_X1 U4338 ( .A1(n38996), .A2(n14562), .ZN(n31765) );
  NOR2_X1 U11271 ( .A1(n28032), .A2(n4347), .ZN(n6114) );
  NAND3_X1 U7622 ( .A1(n9534), .A2(n27948), .A3(n28024), .ZN(n18149) );
  NAND2_X1 U463 ( .A1(n21239), .A2(n27896), .ZN(n31848) );
  INV_X1 U6131 ( .I(n20977), .ZN(n28216) );
  AOI21_X1 U9027 ( .A1(n9702), .A2(n18841), .B(n1069), .ZN(n27711) );
  NOR2_X1 U7394 ( .A1(n15014), .A2(n27955), .ZN(n10052) );
  NAND2_X1 U29492 ( .A1(n1200), .A2(n19124), .ZN(n27872) );
  NOR2_X1 U16785 ( .A1(n1446), .A2(n4306), .ZN(n28242) );
  NAND2_X1 U3376 ( .A1(n14397), .A2(n28181), .ZN(n19123) );
  NAND3_X1 U29560 ( .A1(n28171), .A2(n19601), .A3(n28260), .ZN(n28173) );
  OAI21_X1 U400 ( .A1(n14562), .A2(n1454), .B(n1206), .ZN(n3230) );
  OAI21_X1 U6660 ( .A1(n1202), .A2(n38666), .B(n11737), .ZN(n9237) );
  OAI21_X1 U19708 ( .A1(n31616), .A2(n33292), .B(n31607), .ZN(n13455) );
  NOR2_X1 U11206 ( .A1(n28227), .A2(n19891), .ZN(n20225) );
  NAND2_X1 U2376 ( .A1(n27900), .A2(n11461), .ZN(n28203) );
  NAND2_X1 U14904 ( .A1(n7635), .A2(n31022), .ZN(n28085) );
  NAND2_X1 U5895 ( .A1(n17770), .A2(n7851), .ZN(n16994) );
  NOR2_X1 U11170 ( .A1(n4415), .A2(n3832), .ZN(n2667) );
  OAI21_X1 U9036 ( .A1(n6245), .A2(n7223), .B(n38762), .ZN(n6244) );
  NOR2_X1 U29476 ( .A1(n36689), .A2(n6693), .ZN(n6243) );
  NAND2_X1 U24491 ( .A1(n15572), .A2(n15571), .ZN(n15570) );
  NOR2_X1 U26253 ( .A1(n31607), .A2(n28114), .ZN(n15993) );
  NAND2_X1 U2683 ( .A1(n28274), .A2(n37057), .ZN(n33867) );
  INV_X2 U339 ( .I(n37671), .ZN(n3235) );
  AND2_X1 U17395 ( .A1(n11368), .A2(n28286), .Z(n31871) );
  NAND2_X1 U18268 ( .A1(n28661), .A2(n28660), .ZN(n6041) );
  NAND3_X1 U296 ( .A1(n1451), .A2(n27962), .A3(n10254), .ZN(n11893) );
  AOI21_X1 U7668 ( .A1(n15249), .A2(n42), .B(n28111), .ZN(n11518) );
  OAI22_X1 U19497 ( .A1(n27918), .A2(n200), .B1(n7635), .B2(n6777), .ZN(n20533) );
  INV_X1 U6129 ( .I(n16261), .ZN(n7541) );
  NAND2_X1 U5923 ( .A1(n28284), .A2(n28283), .ZN(n11323) );
  NAND2_X1 U29384 ( .A1(n38579), .A2(n28079), .ZN(n28351) );
  NAND2_X1 U18987 ( .A1(n7555), .A2(n28458), .ZN(n31854) );
  NOR2_X1 U28497 ( .A1(n14615), .A2(n36591), .ZN(n16964) );
  OAI21_X1 U353 ( .A1(n28168), .A2(n20398), .B(n30995), .ZN(n11322) );
  AOI21_X1 U1992 ( .A1(n27920), .A2(n1070), .B(n987), .ZN(n27921) );
  AOI21_X1 U22881 ( .A1(n33669), .A2(n32705), .B(n35862), .ZN(n17476) );
  AOI21_X1 U9023 ( .A1(n28243), .A2(n1444), .B(n28242), .ZN(n28244) );
  NAND2_X1 U3197 ( .A1(n6117), .A2(n8149), .ZN(n6116) );
  OAI21_X1 U28075 ( .A1(n36559), .A2(n36558), .B(n3990), .ZN(n28263) );
  NAND2_X1 U17455 ( .A1(n7719), .A2(n1072), .ZN(n7718) );
  NAND2_X1 U29512 ( .A1(n27935), .A2(n28142), .ZN(n28346) );
  NAND2_X1 U3059 ( .A1(n12227), .A2(n33048), .ZN(n28087) );
  BUF_X2 U17250 ( .I(n19675), .Z(n16777) );
  INV_X1 U4600 ( .I(n3664), .ZN(n28657) );
  INV_X1 U10584 ( .I(n1823), .ZN(n31855) );
  OAI21_X1 U328 ( .A1(n28660), .A2(n1431), .B(n6041), .ZN(n6040) );
  INV_X2 U22893 ( .I(n1195), .ZN(n28812) );
  NOR2_X1 U7492 ( .A1(n3252), .A2(n28369), .ZN(n13820) );
  INV_X1 U23003 ( .I(n28661), .ZN(n28553) );
  NAND2_X1 U387 ( .A1(n2822), .A2(n89), .ZN(n36986) );
  NAND2_X1 U29630 ( .A1(n16778), .A2(n16777), .ZN(n12653) );
  NAND2_X1 U14405 ( .A1(n31597), .A2(n14760), .ZN(n15024) );
  NAND2_X1 U17068 ( .A1(n11005), .A2(n11006), .ZN(n31542) );
  INV_X2 U1605 ( .I(n2191), .ZN(n1419) );
  INV_X2 U424 ( .I(n37758), .ZN(n28554) );
  CLKBUF_X2 U16637 ( .I(n16067), .Z(n32543) );
  INV_X1 U6124 ( .I(n8476), .ZN(n28690) );
  OR2_X1 U11158 ( .A1(n496), .A2(n14193), .Z(n16398) );
  INV_X1 U12547 ( .I(n20445), .ZN(n1434) );
  INV_X2 U23536 ( .I(n28677), .ZN(n18883) );
  INV_X1 U3620 ( .I(n9290), .ZN(n9329) );
  INV_X1 U6611 ( .I(n28728), .ZN(n28323) );
  INV_X1 U15324 ( .I(n3538), .ZN(n14987) );
  INV_X2 U5123 ( .I(n6405), .ZN(n28378) );
  NOR2_X1 U2443 ( .A1(n28724), .A2(n37311), .ZN(n20736) );
  INV_X1 U11085 ( .I(n15024), .ZN(n12715) );
  NOR2_X1 U10699 ( .A1(n28727), .A2(n15752), .ZN(n34433) );
  NAND2_X1 U11001 ( .A1(n3252), .A2(n38556), .ZN(n3250) );
  NAND2_X1 U7577 ( .A1(n974), .A2(n28339), .ZN(n12539) );
  NAND3_X1 U18307 ( .A1(n36775), .A2(n38669), .A3(n36774), .ZN(n36773) );
  NAND2_X1 U19673 ( .A1(n32791), .A2(n28753), .ZN(n12313) );
  OAI21_X1 U194 ( .A1(n28697), .A2(n9648), .B(n10587), .ZN(n16495) );
  NOR2_X1 U11011 ( .A1(n14605), .A2(n28654), .ZN(n11800) );
  NOR2_X1 U16960 ( .A1(n2330), .A2(n33436), .ZN(n33640) );
  INV_X1 U309 ( .I(n6067), .ZN(n33046) );
  INV_X2 U420 ( .I(n33047), .ZN(n28639) );
  INV_X2 U1817 ( .I(n11164), .ZN(n9444) );
  NAND2_X1 U224 ( .A1(n14621), .A2(n11697), .ZN(n28444) );
  INV_X2 U6609 ( .I(n6892), .ZN(n28530) );
  INV_X1 U6623 ( .I(n15224), .ZN(n1192) );
  INV_X1 U24550 ( .I(n28434), .ZN(n28380) );
  INV_X2 U211 ( .I(n13690), .ZN(n18871) );
  INV_X1 U23547 ( .I(n9575), .ZN(n20494) );
  INV_X1 U5598 ( .I(n19759), .ZN(n28808) );
  INV_X1 U6112 ( .I(n11831), .ZN(n1066) );
  INV_X1 U7572 ( .I(n31015), .ZN(n28312) );
  NAND2_X1 U16872 ( .A1(n1194), .A2(n28659), .ZN(n28555) );
  OAI21_X1 U7522 ( .A1(n28732), .A2(n17073), .B(n32595), .ZN(n13784) );
  NAND3_X1 U26291 ( .A1(n15112), .A2(n31321), .A3(n28717), .ZN(n28709) );
  NAND2_X1 U19535 ( .A1(n35777), .A2(n902), .ZN(n18088) );
  NAND2_X1 U11089 ( .A1(n13061), .A2(n8349), .ZN(n13060) );
  NOR2_X1 U9101 ( .A1(n36892), .A2(n13891), .ZN(n31206) );
  NOR2_X1 U2375 ( .A1(n28765), .A2(n28812), .ZN(n13964) );
  NAND2_X1 U27381 ( .A1(n1426), .A2(n39363), .ZN(n18859) );
  NOR2_X1 U27004 ( .A1(n10618), .A2(n17771), .ZN(n18096) );
  NAND3_X1 U17230 ( .A1(n18281), .A2(n36775), .A3(n37863), .ZN(n8320) );
  OAI22_X1 U16199 ( .A1(n28554), .A2(n28551), .B1(n28427), .B2(n1431), .ZN(
        n28428) );
  INV_X1 U15567 ( .I(n36685), .ZN(n28415) );
  INV_X1 U2583 ( .I(n18960), .ZN(n28450) );
  NOR2_X1 U8947 ( .A1(n12539), .A2(n11488), .ZN(n12538) );
  INV_X1 U22568 ( .I(n32338), .ZN(n35804) );
  INV_X1 U13367 ( .I(n39435), .ZN(n34737) );
  NAND2_X1 U7519 ( .A1(n16255), .A2(n16295), .ZN(n16256) );
  AOI21_X1 U12528 ( .A1(n8637), .A2(n12336), .B(n34559), .ZN(n34627) );
  INV_X1 U5444 ( .I(n18972), .ZN(n36145) );
  NAND2_X1 U8841 ( .A1(n32376), .A2(n14222), .ZN(n16657) );
  NAND2_X1 U7508 ( .A1(n33100), .A2(n978), .ZN(n15457) );
  NAND2_X1 U6575 ( .A1(n14816), .A2(n14604), .ZN(n21145) );
  INV_X2 U185 ( .I(n28530), .ZN(n11390) );
  BUF_X2 U284 ( .I(n28638), .Z(n4369) );
  NAND2_X1 U305 ( .A1(n33436), .A2(n1431), .ZN(n28439) );
  NOR2_X1 U2817 ( .A1(n3598), .A2(n18883), .ZN(n32952) );
  AND2_X1 U18767 ( .A1(n28478), .A2(n1414), .Z(n28309) );
  NAND2_X1 U5417 ( .A1(n7486), .A2(n38231), .ZN(n34958) );
  NOR2_X1 U30542 ( .A1(n11438), .A2(n11490), .ZN(n33910) );
  NAND2_X1 U17096 ( .A1(n28494), .A2(n1434), .ZN(n12890) );
  NOR2_X1 U7528 ( .A1(n28530), .A2(n12237), .ZN(n10910) );
  NAND2_X1 U19623 ( .A1(n18972), .A2(n30931), .ZN(n28489) );
  NAND2_X1 U23221 ( .A1(n32703), .A2(n15580), .ZN(n14506) );
  OAI21_X1 U3465 ( .A1(n4969), .A2(n28510), .B(n28715), .ZN(n7799) );
  OAI21_X1 U13605 ( .A1(n888), .A2(n28293), .B(n32286), .ZN(n15514) );
  NAND3_X1 U19563 ( .A1(n10587), .A2(n9598), .A3(n37081), .ZN(n28520) );
  NAND2_X1 U27412 ( .A1(n34244), .A2(n9917), .ZN(n28522) );
  OAI21_X1 U1705 ( .A1(n28386), .A2(n4950), .B(n4949), .ZN(n27958) );
  NAND2_X1 U1812 ( .A1(n28754), .A2(n28755), .ZN(n16922) );
  OAI21_X1 U1700 ( .A1(n28368), .A2(n18972), .B(n28490), .ZN(n9625) );
  NAND2_X1 U11043 ( .A1(n28293), .A2(n28771), .ZN(n11465) );
  OAI21_X1 U2832 ( .A1(n27457), .A2(n28535), .B(n28537), .ZN(n3129) );
  NAND2_X1 U5991 ( .A1(n28756), .A2(n21027), .ZN(n21026) );
  OAI21_X1 U25310 ( .A1(n37758), .A2(n33436), .B(n19688), .ZN(n28558) );
  NAND2_X1 U10926 ( .A1(n28343), .A2(n34007), .ZN(n11664) );
  AOI21_X1 U9282 ( .A1(n38556), .A2(n28604), .B(n34298), .ZN(n35621) );
  AOI21_X1 U258 ( .A1(n28617), .A2(n3664), .B(n28654), .ZN(n28618) );
  OAI21_X1 U11039 ( .A1(n9638), .A2(n28348), .B(n9141), .ZN(n16932) );
  OAI22_X1 U16555 ( .A1(n5399), .A2(n5396), .B1(n9586), .B2(n38203), .ZN(n5398) );
  OAI21_X1 U7504 ( .A1(n11438), .A2(n7913), .B(n11490), .ZN(n8854) );
  NOR2_X1 U6591 ( .A1(n20497), .A2(n1823), .ZN(n20493) );
  NAND3_X1 U6105 ( .A1(n12990), .A2(n28453), .A3(n37204), .ZN(n12378) );
  CLKBUF_X2 U4056 ( .I(n11695), .Z(n3703) );
  OR2_X1 U8935 ( .A1(n28529), .A2(n37619), .Z(n11491) );
  NOR2_X1 U29616 ( .A1(n36777), .A2(n28516), .ZN(n28518) );
  AOI22_X1 U8940 ( .A1(n12605), .A2(n28608), .B1(n11390), .B2(n33647), .ZN(
        n6094) );
  OAI21_X1 U4645 ( .A1(n8323), .A2(n8322), .B(n7555), .ZN(n8321) );
  CLKBUF_X2 U5406 ( .I(n7744), .Z(n32448) );
  CLKBUF_X2 U20153 ( .I(n29160), .Z(n33511) );
  INV_X1 U12735 ( .I(n10079), .ZN(n29127) );
  AOI21_X1 U16185 ( .A1(n28808), .A2(n33577), .B(n35083), .ZN(n35082) );
  INV_X1 U24689 ( .I(n28874), .ZN(n16310) );
  INV_X1 U16688 ( .I(n9787), .ZN(n21007) );
  BUF_X2 U16761 ( .I(n20465), .Z(n2392) );
  BUF_X2 U12189 ( .I(n9036), .Z(n3665) );
  INV_X1 U10970 ( .I(n10080), .ZN(n28927) );
  INV_X1 U15141 ( .I(n14941), .ZN(n28977) );
  INV_X1 U209 ( .I(n28827), .ZN(n28978) );
  INV_X2 U14654 ( .I(n20686), .ZN(n29862) );
  INV_X2 U3894 ( .I(n10896), .ZN(n19962) );
  INV_X1 U15637 ( .I(n6163), .ZN(n31428) );
  INV_X2 U3162 ( .I(n21270), .ZN(n13441) );
  CLKBUF_X2 U10903 ( .I(n29424), .Z(n19896) );
  BUF_X2 U15438 ( .I(n28436), .Z(n29700) );
  INV_X2 U27831 ( .I(n19424), .ZN(n1407) );
  INV_X1 U15667 ( .I(n32251), .ZN(n29195) );
  INV_X2 U138 ( .I(n18315), .ZN(n29595) );
  INV_X1 U30866 ( .I(n12829), .ZN(n31279) );
  INV_X1 U189 ( .I(n20026), .ZN(n29310) );
  INV_X1 U14084 ( .I(n18288), .ZN(n30195) );
  INV_X1 U18048 ( .I(n14254), .ZN(n17238) );
  NAND2_X1 U7442 ( .A1(n1179), .A2(n18720), .ZN(n4655) );
  INV_X1 U30865 ( .I(n18667), .ZN(n33928) );
  INV_X1 U3505 ( .I(n29701), .ZN(n8941) );
  INV_X2 U5081 ( .I(n30043), .ZN(n1056) );
  OR2_X1 U4102 ( .A1(n30049), .A2(n33256), .Z(n4255) );
  INV_X1 U19400 ( .I(n16217), .ZN(n29935) );
  INV_X2 U8853 ( .I(n20979), .ZN(n30680) );
  INV_X1 U4963 ( .I(n15854), .ZN(n29996) );
  NAND2_X1 U30098 ( .A1(n6019), .A2(n1057), .ZN(n29986) );
  INV_X2 U6555 ( .I(n30220), .ZN(n1177) );
  INV_X1 U18092 ( .I(n16599), .ZN(n20982) );
  INV_X2 U8079 ( .I(n34000), .ZN(n29779) );
  OR2_X1 U180 ( .A1(n33256), .A2(n11896), .Z(n30048) );
  INV_X1 U1576 ( .I(n20687), .ZN(n29863) );
  INV_X1 U127 ( .I(n11428), .ZN(n30162) );
  INV_X1 U156 ( .I(n33967), .ZN(n29445) );
  INV_X1 U94 ( .I(n21023), .ZN(n17644) );
  NOR2_X1 U10035 ( .A1(n20525), .A2(n30153), .ZN(n30796) );
  INV_X1 U23169 ( .I(n11783), .ZN(n30241) );
  INV_X2 U74 ( .I(n29596), .ZN(n12450) );
  NAND2_X1 U16855 ( .A1(n3700), .A2(n3631), .ZN(n3698) );
  NOR2_X1 U27617 ( .A1(n30048), .A2(n32628), .ZN(n19454) );
  INV_X1 U9831 ( .I(n34344), .ZN(n18007) );
  NOR2_X1 U4808 ( .A1(n32945), .A2(n13153), .ZN(n32944) );
  INV_X1 U25496 ( .I(n29586), .ZN(n21264) );
  NAND2_X1 U2753 ( .A1(n9394), .A2(n15153), .ZN(n14495) );
  NAND2_X1 U23797 ( .A1(n16510), .A2(n971), .ZN(n13085) );
  INV_X1 U3284 ( .I(n20982), .ZN(n1398) );
  NOR2_X1 U10835 ( .A1(n30187), .A2(n39280), .ZN(n29061) );
  NAND2_X1 U7483 ( .A1(n29777), .A2(n33964), .ZN(n29780) );
  INV_X2 U87 ( .I(n6019), .ZN(n29987) );
  AOI21_X1 U8856 ( .A1(n771), .A2(n29446), .B(n1401), .ZN(n16508) );
  AOI21_X1 U2816 ( .A1(n29378), .A2(n29458), .B(n29377), .ZN(n29345) );
  AOI21_X1 U7413 ( .A1(n5570), .A2(n921), .B(n3700), .ZN(n9799) );
  INV_X1 U8875 ( .I(n1399), .ZN(n11574) );
  INV_X1 U120 ( .I(n21285), .ZN(n21287) );
  NOR2_X1 U7399 ( .A1(n28864), .A2(n29587), .ZN(n13670) );
  INV_X1 U29771 ( .I(n32906), .ZN(n29266) );
  NOR2_X1 U15054 ( .A1(n29348), .A2(n29286), .ZN(n29211) );
  INV_X1 U116 ( .I(n20018), .ZN(n11056) );
  NAND2_X1 U4964 ( .A1(n29946), .A2(n32571), .ZN(n19137) );
  OR2_X1 U5374 ( .A1(n29701), .A2(n16599), .Z(n34180) );
  AND2_X1 U10861 ( .A1(n21023), .A2(n28843), .Z(n29634) );
  INV_X1 U142 ( .I(n29941), .ZN(n30051) );
  INV_X1 U5584 ( .I(n344), .ZN(n16209) );
  INV_X2 U5587 ( .I(n32946), .ZN(n907) );
  NOR2_X1 U111 ( .A1(n1181), .A2(n30160), .ZN(n35849) );
  NOR2_X1 U6526 ( .A1(n2456), .A2(n19992), .ZN(n2016) );
  NOR2_X1 U3536 ( .A1(n29449), .A2(n771), .ZN(n29350) );
  NAND2_X1 U7400 ( .A1(n16074), .A2(n14151), .ZN(n2132) );
  NOR2_X1 U7388 ( .A1(n13670), .A2(n13672), .ZN(n13669) );
  NOR2_X1 U2459 ( .A1(n1404), .A2(n29595), .ZN(n2378) );
  NAND2_X1 U29679 ( .A1(n30159), .A2(n1399), .ZN(n33488) );
  OAI21_X1 U10754 ( .A1(n14755), .A2(n12054), .B(n38262), .ZN(n12060) );
  INV_X1 U16558 ( .I(n32894), .ZN(n30045) );
  AOI21_X1 U30336 ( .A1(n29694), .A2(n21037), .B(n2559), .ZN(n33760) );
  NAND2_X1 U14473 ( .A1(n33094), .A2(n34858), .ZN(n30396) );
  NAND2_X1 U3084 ( .A1(n33277), .A2(n1400), .ZN(n7908) );
  OAI21_X1 U2418 ( .A1(n29634), .A2(n29704), .B(n16209), .ZN(n17348) );
  NAND2_X1 U93 ( .A1(n36207), .A2(n1755), .ZN(n33393) );
  NOR2_X1 U3540 ( .A1(n29449), .A2(n1176), .ZN(n19791) );
  OAI21_X1 U10808 ( .A1(n2121), .A2(n18815), .B(n19508), .ZN(n3245) );
  OAI21_X1 U27258 ( .A1(n29843), .A2(n773), .B(n18477), .ZN(n29873) );
  NOR2_X1 U67 ( .A1(n33394), .A2(n33393), .ZN(n18590) );
  NOR2_X1 U77 ( .A1(n34973), .A2(n29378), .ZN(n35295) );
  NAND2_X1 U75 ( .A1(n36023), .A2(n36022), .ZN(n4799) );
  INV_X1 U18838 ( .I(n6332), .ZN(n10869) );
  AOI21_X1 U16296 ( .A1(n17842), .A2(n39416), .B(n14183), .ZN(n35096) );
  INV_X1 U17289 ( .I(n9828), .ZN(n14126) );
  INV_X1 U72 ( .I(n20208), .ZN(n29534) );
  INV_X2 U26258 ( .I(n18081), .ZN(n1174) );
  INV_X1 U4068 ( .I(n29277), .ZN(n1379) );
  INV_X2 U46 ( .I(n9105), .ZN(n969) );
  INV_X1 U26874 ( .I(n29659), .ZN(n17382) );
  INV_X1 U9482 ( .I(n29930), .ZN(n29922) );
  CLKBUF_X2 U5567 ( .I(n29475), .Z(n18873) );
  CLKBUF_X2 U2906 ( .I(n30079), .Z(n31120) );
  INV_X1 U2890 ( .I(n17469), .ZN(n30129) );
  INV_X1 U3016 ( .I(n29979), .ZN(n29975) );
  INV_X1 U23831 ( .I(n29208), .ZN(n13142) );
  INV_X1 U61 ( .I(n29367), .ZN(n16683) );
  INV_X1 U6126 ( .I(n30262), .ZN(n1172) );
  NOR2_X1 U49 ( .A1(n28585), .A2(n28584), .ZN(n17262) );
  INV_X1 U4040 ( .I(n29684), .ZN(n29675) );
  NAND2_X1 U18806 ( .A1(n31821), .A2(n10978), .ZN(n30134) );
  INV_X1 U41 ( .I(n20078), .ZN(n30069) );
  INV_X1 U6066 ( .I(n20307), .ZN(n30132) );
  AND2_X1 U55 ( .A1(n31821), .A2(n10978), .Z(n34177) );
  INV_X1 U29921 ( .I(n33437), .ZN(n36738) );
  INV_X1 U5831 ( .I(n29929), .ZN(n3860) );
  INV_X1 U23 ( .I(n30022), .ZN(n30035) );
  NAND2_X1 U17382 ( .A1(n38164), .A2(n17192), .ZN(n33207) );
  NAND2_X1 U2186 ( .A1(n29478), .A2(n29468), .ZN(n29464) );
  INV_X1 U7363 ( .I(n29981), .ZN(n29977) );
  INV_X1 U30801 ( .I(n30107), .ZN(n30119) );
  INV_X1 U14 ( .I(n13192), .ZN(n29811) );
  INV_X1 U3836 ( .I(n15509), .ZN(n29209) );
  NAND2_X1 U3577 ( .A1(n30038), .A2(n9231), .ZN(n30014) );
  INV_X2 U47 ( .I(n29859), .ZN(n29851) );
  NOR2_X1 U17211 ( .A1(n1385), .A2(n32508), .ZN(n8286) );
  NAND2_X1 U2919 ( .A1(n29567), .A2(n31899), .ZN(n29565) );
  INV_X1 U7371 ( .I(n29530), .ZN(n29527) );
  INV_X1 U17564 ( .I(n29740), .ZN(n19348) );
  INV_X1 U7370 ( .I(n30093), .ZN(n30098) );
  INV_X1 U19739 ( .I(n37096), .ZN(n29369) );
  INV_X1 U18 ( .I(n17192), .ZN(n17193) );
  NAND2_X1 U20893 ( .A1(n10813), .A2(n8286), .ZN(n9261) );
  NAND3_X1 U2 ( .A1(n29368), .A2(n13839), .A3(n13804), .ZN(n39677) );
  AOI22_X1 U6 ( .A1(n19090), .A2(n5530), .B1(n29277), .B2(n37157), .ZN(n17773)
         );
  AND2_X1 U7 ( .A1(n4368), .A2(n12198), .Z(n4367) );
  NOR2_X1 U8 ( .A1(n20538), .A2(n4368), .ZN(n30171) );
  INV_X1 U10 ( .I(n29336), .ZN(n29335) );
  NAND2_X1 U11 ( .A1(n2792), .A2(n29802), .ZN(n29806) );
  NAND2_X1 U15 ( .A1(n10118), .A2(n30117), .ZN(n30106) );
  BUF_X2 U20 ( .I(n3096), .Z(n36096) );
  INV_X1 U21 ( .I(n29231), .ZN(n1387) );
  INV_X1 U22 ( .I(n29802), .ZN(n29813) );
  AND2_X1 U24 ( .A1(n30097), .A2(n31601), .Z(n16471) );
  NAND2_X1 U26 ( .A1(n35272), .A2(n16260), .ZN(n15044) );
  INV_X1 U30 ( .I(n85), .ZN(n9913) );
  INV_X1 U33 ( .I(n29678), .ZN(n1173) );
  INV_X2 U34 ( .I(n12198), .ZN(n20538) );
  INV_X2 U36 ( .I(n20274), .ZN(n10813) );
  INV_X1 U38 ( .I(n30213), .ZN(n33521) );
  INV_X1 U45 ( .I(n31899), .ZN(n1053) );
  NOR2_X1 U48 ( .A1(n38164), .A2(n1385), .ZN(n37724) );
  NAND2_X1 U52 ( .A1(n29810), .A2(n13192), .ZN(n5970) );
  OR2_X1 U54 ( .A1(n19475), .A2(n20160), .Z(n37157) );
  NAND2_X1 U56 ( .A1(n4072), .A2(n33071), .ZN(n33070) );
  INV_X2 U57 ( .I(n8039), .ZN(n30034) );
  AOI22_X1 U58 ( .A1(n29595), .A2(n2296), .B1(n31667), .B2(n14417), .ZN(n36193) );
  NAND2_X1 U62 ( .A1(n29427), .A2(n29449), .ZN(n38805) );
  AOI21_X1 U66 ( .A1(n30165), .A2(n30046), .B(n39416), .ZN(n36023) );
  OAI21_X1 U69 ( .A1(n7207), .A2(n39322), .B(n19162), .ZN(n20160) );
  AND2_X1 U70 ( .A1(n29942), .A2(n30059), .Z(n37177) );
  OAI21_X1 U71 ( .A1(n29485), .A2(n19962), .B(n32197), .ZN(n29489) );
  NAND2_X1 U76 ( .A1(n37752), .A2(n20673), .ZN(n5924) );
  NAND2_X1 U83 ( .A1(n37376), .A2(n37614), .ZN(n37375) );
  NAND2_X1 U84 ( .A1(n16508), .A2(n32671), .ZN(n37797) );
  OAI21_X1 U85 ( .A1(n38919), .A2(n6938), .B(n29202), .ZN(n38773) );
  OAI21_X1 U86 ( .A1(n20289), .A2(n29635), .B(n18107), .ZN(n35762) );
  NAND2_X1 U89 ( .A1(n2954), .A2(n29459), .ZN(n34194) );
  OAI22_X1 U99 ( .A1(n29457), .A2(n31521), .B1(n13261), .B2(n29458), .ZN(n8924) );
  AOI22_X1 U102 ( .A1(n29939), .A2(n6019), .B1(n29987), .B2(n30051), .ZN(
        n34681) );
  AND2_X1 U103 ( .A1(n5348), .A2(n20080), .Z(n29899) );
  INV_X1 U107 ( .I(n773), .ZN(n29867) );
  INV_X1 U110 ( .I(n28882), .ZN(n8762) );
  NAND2_X1 U113 ( .A1(n16672), .A2(n1755), .ZN(n31065) );
  CLKBUF_X2 U122 ( .I(n29454), .Z(n39647) );
  OR2_X1 U123 ( .A1(n1056), .A2(n4220), .Z(n37082) );
  CLKBUF_X4 U124 ( .I(n4879), .Z(n37936) );
  OAI21_X1 U125 ( .A1(n37729), .A2(n37728), .B(n37727), .ZN(n29011) );
  NOR2_X1 U129 ( .A1(n36102), .A2(n30680), .ZN(n36101) );
  NAND2_X1 U133 ( .A1(n11634), .A2(n29263), .ZN(n11595) );
  NAND2_X1 U136 ( .A1(n773), .A2(n4879), .ZN(n33093) );
  NAND2_X1 U140 ( .A1(n36481), .A2(n30160), .ZN(n38883) );
  NAND2_X1 U145 ( .A1(n29781), .A2(n34000), .ZN(n10746) );
  INV_X1 U146 ( .I(n15089), .ZN(n37858) );
  OAI21_X1 U148 ( .A1(n37368), .A2(n29942), .B(n30059), .ZN(n29171) );
  BUF_X4 U149 ( .I(n29500), .Z(n38051) );
  INV_X1 U152 ( .I(n29642), .ZN(n37879) );
  BUF_X2 U155 ( .I(n30195), .Z(n36225) );
  INV_X1 U159 ( .I(n28843), .ZN(n28882) );
  INV_X1 U164 ( .I(n29346), .ZN(n38822) );
  CLKBUF_X2 U168 ( .I(n777), .Z(n39322) );
  INV_X1 U170 ( .I(n3631), .ZN(n38709) );
  NAND2_X1 U172 ( .A1(n29642), .A2(n29643), .ZN(n38129) );
  INV_X1 U173 ( .I(n30156), .ZN(n29210) );
  BUF_X2 U174 ( .I(n4671), .Z(n31511) );
  INV_X2 U175 ( .I(n30057), .ZN(n37021) );
  INV_X1 U176 ( .I(n19428), .ZN(n31689) );
  NOR2_X1 U184 ( .A1(n35823), .A2(n16036), .ZN(n38161) );
  NAND2_X1 U186 ( .A1(n28636), .A2(n10061), .ZN(n29025) );
  INV_X1 U187 ( .I(n19571), .ZN(n37726) );
  INV_X1 U188 ( .I(n28830), .ZN(n1410) );
  NAND2_X1 U192 ( .A1(n5342), .A2(n8048), .ZN(n37637) );
  NOR2_X1 U195 ( .A1(n38855), .A2(n39473), .ZN(n38463) );
  NOR2_X1 U196 ( .A1(n34173), .A2(n35997), .ZN(n37555) );
  NAND2_X1 U197 ( .A1(n34958), .A2(n39555), .ZN(n28331) );
  NAND2_X1 U198 ( .A1(n39000), .A2(n38997), .ZN(n28648) );
  OAI21_X1 U202 ( .A1(n3018), .A2(n3019), .B(n28390), .ZN(n37990) );
  NAND2_X1 U206 ( .A1(n38399), .A2(n37285), .ZN(n31393) );
  NOR2_X1 U207 ( .A1(n9444), .A2(n11614), .ZN(n37558) );
  NAND2_X1 U208 ( .A1(n28268), .A2(n16691), .ZN(n15109) );
  NAND2_X1 U210 ( .A1(n28439), .A2(n34176), .ZN(n37577) );
  NAND2_X1 U214 ( .A1(n28336), .A2(n32178), .ZN(n38062) );
  OAI22_X1 U215 ( .A1(n28525), .A2(n28735), .B1(n28736), .B2(n38172), .ZN(
        n38017) );
  AND2_X1 U216 ( .A1(n18871), .A2(n28686), .Z(n18996) );
  OAI21_X1 U218 ( .A1(n28726), .A2(n12237), .B(n38500), .ZN(n3634) );
  AND2_X1 U220 ( .A1(n9878), .A2(n28620), .Z(n28401) );
  NOR2_X1 U223 ( .A1(n28386), .A2(n28653), .ZN(n28368) );
  NOR2_X1 U225 ( .A1(n2937), .A2(n1189), .ZN(n7913) );
  NAND2_X1 U227 ( .A1(n39664), .A2(n28755), .ZN(n21027) );
  NOR2_X1 U228 ( .A1(n28485), .A2(n28390), .ZN(n28178) );
  NAND2_X1 U230 ( .A1(n36776), .A2(n36773), .ZN(n38469) );
  AND2_X1 U233 ( .A1(n1186), .A2(n14987), .Z(n37128) );
  OAI21_X1 U236 ( .A1(n16307), .A2(n17596), .B(n5396), .ZN(n9585) );
  NAND3_X1 U237 ( .A1(n28721), .A2(n28362), .A3(n28361), .ZN(n38399) );
  BUF_X2 U250 ( .I(n28464), .Z(n19827) );
  OAI21_X1 U251 ( .A1(n37561), .A2(n37560), .B(n28724), .ZN(n36585) );
  NOR2_X1 U255 ( .A1(n15235), .A2(n15737), .ZN(n38861) );
  NAND3_X1 U257 ( .A1(n15709), .A2(n37981), .A3(n28639), .ZN(n35351) );
  AND2_X1 U263 ( .A1(n16559), .A2(n16067), .Z(n34173) );
  INV_X1 U266 ( .I(n28730), .ZN(n50) );
  NOR2_X1 U267 ( .A1(n37080), .A2(n33283), .ZN(n32781) );
  NAND2_X1 U271 ( .A1(n31888), .A2(n28473), .ZN(n8094) );
  NAND2_X1 U275 ( .A1(n28580), .A2(n1196), .ZN(n3052) );
  NOR2_X1 U277 ( .A1(n28485), .A2(n16559), .ZN(n3018) );
  NOR2_X1 U278 ( .A1(n16067), .A2(n28484), .ZN(n6629) );
  NOR2_X1 U281 ( .A1(n28699), .A2(n28698), .ZN(n38503) );
  INV_X1 U285 ( .I(n1823), .ZN(n37777) );
  OR2_X1 U286 ( .A1(n38159), .A2(n17751), .Z(n28725) );
  NAND2_X1 U290 ( .A1(n28716), .A2(n1882), .ZN(n28515) );
  NAND2_X1 U291 ( .A1(n31663), .A2(n37758), .ZN(n28440) );
  INV_X2 U294 ( .I(n33283), .ZN(n28746) );
  OR2_X1 U297 ( .A1(n38203), .A2(n39227), .Z(n8158) );
  OR2_X1 U303 ( .A1(n28720), .A2(n28723), .Z(n14604) );
  INV_X2 U304 ( .I(n5418), .ZN(n36414) );
  BUF_X2 U306 ( .I(n28503), .Z(n13891) );
  BUF_X2 U314 ( .I(n28676), .Z(n9599) );
  NAND2_X1 U316 ( .A1(n34861), .A2(n7251), .ZN(n38065) );
  AND2_X1 U317 ( .A1(n28686), .A2(n39724), .Z(n10038) );
  AND2_X1 U318 ( .A1(n10883), .A2(n7063), .Z(n5641) );
  NAND2_X1 U321 ( .A1(n8082), .A2(n11831), .ZN(n21141) );
  OR2_X1 U330 ( .A1(n39227), .A2(n37484), .Z(n34510) );
  NOR2_X1 U331 ( .A1(n28700), .A2(n19349), .ZN(n33793) );
  NOR2_X1 U332 ( .A1(n976), .A2(n13170), .ZN(n38657) );
  NAND2_X1 U345 ( .A1(n38231), .A2(n7429), .ZN(n28073) );
  NAND3_X1 U348 ( .A1(n11330), .A2(n12527), .A3(n36588), .ZN(n38500) );
  NAND2_X1 U352 ( .A1(n28643), .A2(n14448), .ZN(n38999) );
  INV_X1 U354 ( .I(n7905), .ZN(n36110) );
  INV_X2 U365 ( .I(n36588), .ZN(n39435) );
  AND2_X1 U366 ( .A1(n31027), .A2(n30668), .Z(n38231) );
  NOR2_X1 U368 ( .A1(n35203), .A2(n34559), .ZN(n36742) );
  INV_X2 U369 ( .I(n31663), .ZN(n1194) );
  BUF_X2 U370 ( .I(n31378), .Z(n902) );
  BUF_X1 U373 ( .I(n31663), .Z(n39147) );
  INV_X1 U374 ( .I(n28503), .ZN(n28533) );
  CLKBUF_X2 U383 ( .I(n33765), .Z(n33629) );
  INV_X2 U386 ( .I(n17234), .ZN(n32682) );
  INV_X2 U390 ( .I(n34695), .ZN(n1196) );
  OAI21_X1 U396 ( .A1(n15389), .A2(n1444), .B(n8368), .ZN(n20584) );
  NAND2_X1 U401 ( .A1(n11512), .A2(n36643), .ZN(n28349) );
  NAND2_X1 U404 ( .A1(n37785), .A2(n37782), .ZN(n27925) );
  BUF_X4 U411 ( .I(n8366), .Z(n37758) );
  OAI21_X1 U412 ( .A1(n39795), .A2(n39794), .B(n898), .ZN(n27938) );
  NAND2_X1 U416 ( .A1(n38490), .A2(n14461), .ZN(n28038) );
  NAND3_X1 U417 ( .A1(n13491), .A2(n37671), .A3(n19525), .ZN(n28144) );
  OAI21_X1 U418 ( .A1(n30623), .A2(n28028), .B(n27948), .ZN(n38288) );
  OAI21_X1 U421 ( .A1(n12784), .A2(n30995), .B(n16544), .ZN(n28284) );
  OAI22_X1 U427 ( .A1(n36979), .A2(n9969), .B1(n13851), .B2(n16325), .ZN(
        n38490) );
  NAND3_X1 U432 ( .A1(n35507), .A2(n21238), .A3(n28249), .ZN(n38923) );
  NOR2_X1 U433 ( .A1(n37642), .A2(n17057), .ZN(n17055) );
  NAND2_X1 U436 ( .A1(n13409), .A2(n27969), .ZN(n35005) );
  NAND3_X1 U437 ( .A1(n37322), .A2(n28199), .A3(n16461), .ZN(n28202) );
  INV_X1 U439 ( .I(n3990), .ZN(n39188) );
  NAND2_X1 U440 ( .A1(n37784), .A2(n1204), .ZN(n37782) );
  NOR2_X1 U443 ( .A1(n28024), .A2(n14829), .ZN(n30623) );
  OR2_X1 U445 ( .A1(n8207), .A2(n288), .Z(n37126) );
  NAND2_X1 U446 ( .A1(n4347), .A2(n1435), .ZN(n38308) );
  OAI22_X1 U453 ( .A1(n37057), .A2(n988), .B1(n13081), .B2(n14399), .ZN(n8946)
         );
  NOR3_X1 U456 ( .A1(n7872), .A2(n1448), .A3(n38579), .ZN(n38868) );
  INV_X1 U457 ( .I(n38419), .ZN(n20577) );
  NAND2_X1 U460 ( .A1(n14562), .A2(n18689), .ZN(n27887) );
  NAND2_X1 U468 ( .A1(n10466), .A2(n10465), .ZN(n37334) );
  AOI21_X1 U469 ( .A1(n37159), .A2(n27896), .B(n27973), .ZN(n16706) );
  BUF_X2 U470 ( .I(n27964), .Z(n28118) );
  NAND2_X1 U473 ( .A1(n35061), .A2(n28274), .ZN(n32374) );
  NAND2_X1 U474 ( .A1(n3990), .A2(n3989), .ZN(n27981) );
  NAND3_X1 U476 ( .A1(n28165), .A2(n10642), .A3(n988), .ZN(n37035) );
  NAND3_X1 U477 ( .A1(n11375), .A2(n11501), .A3(n37078), .ZN(n406) );
  OR2_X1 U485 ( .A1(n28152), .A2(n16576), .Z(n10465) );
  AND2_X1 U490 ( .A1(n28152), .A2(n16576), .Z(n18770) );
  INV_X1 U492 ( .I(n31494), .ZN(n37783) );
  OR2_X1 U498 ( .A1(n9242), .A2(n36197), .Z(n2603) );
  NAND2_X1 U503 ( .A1(n28282), .A2(n33957), .ZN(n28067) );
  CLKBUF_X2 U504 ( .I(n18689), .Z(n38996) );
  NOR2_X1 U505 ( .A1(n31942), .A2(n28214), .ZN(n34817) );
  NOR2_X1 U508 ( .A1(n14397), .A2(n36573), .ZN(n4767) );
  NAND3_X1 U511 ( .A1(n37), .A2(n1448), .A3(n38579), .ZN(n28325) );
  OAI21_X1 U512 ( .A1(n38307), .A2(n30995), .B(n7528), .ZN(n12809) );
  AOI21_X1 U513 ( .A1(n37754), .A2(n37753), .B(n30773), .ZN(n38327) );
  INV_X1 U525 ( .I(n16576), .ZN(n10420) );
  NAND3_X1 U526 ( .A1(n18777), .A2(n16261), .A3(n34447), .ZN(n12420) );
  NAND2_X1 U535 ( .A1(n39126), .A2(n39127), .ZN(n38678) );
  NAND2_X1 U536 ( .A1(n28238), .A2(n28236), .ZN(n17615) );
  INV_X1 U537 ( .I(n18853), .ZN(n39112) );
  BUF_X2 U544 ( .I(n7741), .Z(n38579) );
  BUF_X2 U545 ( .I(n33957), .Z(n38307) );
  NOR2_X1 U547 ( .A1(n14397), .A2(n28181), .ZN(n39696) );
  INV_X1 U548 ( .I(n11676), .ZN(n1436) );
  INV_X1 U551 ( .I(n38453), .ZN(n34166) );
  BUF_X2 U561 ( .I(n17405), .Z(n2717) );
  INV_X1 U562 ( .I(n2281), .ZN(n38620) );
  INV_X1 U566 ( .I(n13877), .ZN(n37307) );
  INV_X1 U568 ( .I(n21093), .ZN(n38648) );
  INV_X1 U569 ( .I(n31355), .ZN(n8364) );
  AOI21_X1 U573 ( .A1(n27287), .A2(n1080), .B(n6010), .ZN(n16162) );
  NAND3_X1 U576 ( .A1(n10998), .A2(n27059), .A3(n10999), .ZN(n10997) );
  BUF_X2 U577 ( .I(n31767), .Z(n37812) );
  NOR2_X1 U579 ( .A1(n27172), .A2(n19062), .ZN(n27549) );
  AND2_X1 U587 ( .A1(n8253), .A2(n1082), .Z(n8252) );
  NAND3_X1 U590 ( .A1(n37552), .A2(n16514), .A3(n16516), .ZN(n35718) );
  NAND2_X1 U594 ( .A1(n3672), .A2(n3674), .ZN(n38078) );
  OAI22_X1 U596 ( .A1(n5059), .A2(n27310), .B1(n37001), .B2(n27155), .ZN(
        n35123) );
  OR2_X1 U599 ( .A1(n16520), .A2(n27153), .Z(n37552) );
  OAI21_X1 U601 ( .A1(n30871), .A2(n2035), .B(n33335), .ZN(n30584) );
  AOI21_X1 U603 ( .A1(n27250), .A2(n27007), .B(n27251), .ZN(n5770) );
  NAND2_X1 U607 ( .A1(n30582), .A2(n37170), .ZN(n17107) );
  NAND2_X1 U609 ( .A1(n10032), .A2(n35905), .ZN(n38047) );
  OAI21_X1 U610 ( .A1(n37704), .A2(n37703), .B(n37040), .ZN(n35914) );
  NAND2_X1 U611 ( .A1(n36744), .A2(n33619), .ZN(n16306) );
  NAND2_X1 U613 ( .A1(n37512), .A2(n27398), .ZN(n27073) );
  INV_X1 U614 ( .I(n35243), .ZN(n31584) );
  OAI22_X1 U620 ( .A1(n14327), .A2(n6908), .B1(n2761), .B2(n27165), .ZN(n14326) );
  NOR2_X1 U621 ( .A1(n2207), .A2(n32020), .ZN(n39236) );
  NAND2_X1 U624 ( .A1(n5059), .A2(n39206), .ZN(n38481) );
  OAI21_X1 U631 ( .A1(n39632), .A2(n6534), .B(n38690), .ZN(n34570) );
  AND2_X1 U634 ( .A1(n17095), .A2(n3977), .Z(n11038) );
  NAND3_X1 U636 ( .A1(n7588), .A2(n33088), .A3(n18717), .ZN(n10578) );
  INV_X1 U639 ( .I(n26749), .ZN(n491) );
  INV_X1 U645 ( .I(n27393), .ZN(n31400) );
  NAND2_X1 U646 ( .A1(n39632), .A2(n6534), .ZN(n37854) );
  NAND2_X1 U648 ( .A1(n37655), .A2(n37652), .ZN(n32545) );
  NOR2_X1 U649 ( .A1(n32555), .A2(n34167), .ZN(n39230) );
  NOR2_X1 U655 ( .A1(n32566), .A2(n38187), .ZN(n3531) );
  NAND2_X1 U658 ( .A1(n12020), .A2(n35826), .ZN(n39565) );
  NOR2_X1 U660 ( .A1(n161), .A2(n160), .ZN(n30667) );
  CLKBUF_X2 U664 ( .I(n1226), .Z(n34520) );
  OR2_X1 U665 ( .A1(n32926), .A2(n36496), .Z(n37170) );
  INV_X1 U667 ( .I(n37603), .ZN(n30732) );
  NAND2_X1 U674 ( .A1(n27021), .A2(n15360), .ZN(n38276) );
  NAND2_X1 U677 ( .A1(n38489), .A2(n38488), .ZN(n6195) );
  NAND2_X1 U679 ( .A1(n13294), .A2(n36911), .ZN(n38565) );
  OR2_X1 U680 ( .A1(n14881), .A2(n35895), .Z(n32960) );
  NAND2_X1 U682 ( .A1(n14327), .A2(n27389), .ZN(n34733) );
  NAND2_X1 U691 ( .A1(n20133), .A2(n10051), .ZN(n37465) );
  NAND2_X1 U693 ( .A1(n35332), .A2(n27304), .ZN(n39283) );
  NOR2_X1 U694 ( .A1(n27230), .A2(n1085), .ZN(n37704) );
  NAND3_X1 U698 ( .A1(n4782), .A2(n16782), .A3(n33593), .ZN(n36744) );
  OAI21_X1 U700 ( .A1(n27270), .A2(n27196), .B(n27272), .ZN(n38739) );
  OAI21_X1 U701 ( .A1(n19557), .A2(n7096), .B(n1225), .ZN(n39573) );
  NAND2_X1 U707 ( .A1(n27357), .A2(n27358), .ZN(n2208) );
  NAND2_X1 U708 ( .A1(n5101), .A2(n39414), .ZN(n27456) );
  OR2_X1 U709 ( .A1(n10171), .A2(n2722), .Z(n27090) );
  OR2_X1 U711 ( .A1(n1788), .A2(n7757), .Z(n37076) );
  AND2_X1 U712 ( .A1(n31006), .A2(n7424), .Z(n37246) );
  INV_X2 U713 ( .I(n27164), .ZN(n20981) );
  OR2_X1 U714 ( .A1(n27248), .A2(n7975), .Z(n35730) );
  BUF_X2 U716 ( .I(n3540), .Z(n36865) );
  NAND2_X1 U717 ( .A1(n27378), .A2(n1788), .ZN(n27071) );
  NAND2_X1 U718 ( .A1(n11083), .A2(n14153), .ZN(n14086) );
  OAI22_X1 U727 ( .A1(n998), .A2(n35265), .B1(n32829), .B2(n27424), .ZN(n9268)
         );
  AND2_X1 U731 ( .A1(n19455), .A2(n27197), .Z(n14695) );
  INV_X1 U733 ( .I(n31014), .ZN(n30758) );
  NAND2_X1 U734 ( .A1(n36200), .A2(n34969), .ZN(n16170) );
  INV_X1 U736 ( .I(n27452), .ZN(n5932) );
  INV_X1 U737 ( .I(n36969), .ZN(n2923) );
  INV_X1 U738 ( .I(n27095), .ZN(n33593) );
  INV_X1 U743 ( .I(n5588), .ZN(n39546) );
  INV_X2 U748 ( .I(n9875), .ZN(n21144) );
  NAND2_X1 U752 ( .A1(n27211), .A2(n34977), .ZN(n27441) );
  INV_X2 U762 ( .I(n11820), .ZN(n10051) );
  INV_X1 U765 ( .I(n27434), .ZN(n39150) );
  CLKBUF_X4 U766 ( .I(n32566), .Z(n36528) );
  NAND3_X1 U768 ( .A1(n4782), .A2(n2660), .A3(n36496), .ZN(n38618) );
  NAND2_X1 U769 ( .A1(n4272), .A2(n6191), .ZN(n15641) );
  INV_X2 U771 ( .I(n39050), .ZN(n39826) );
  BUF_X2 U772 ( .I(n27446), .Z(n4782) );
  OAI21_X1 U773 ( .A1(n30365), .A2(n32958), .B(n36477), .ZN(n36476) );
  BUF_X2 U774 ( .I(n998), .Z(n30544) );
  NAND3_X1 U777 ( .A1(n26892), .A2(n4325), .A3(n33396), .ZN(n4324) );
  NOR3_X1 U778 ( .A1(n26663), .A2(n32009), .A3(n26662), .ZN(n39754) );
  NOR2_X1 U782 ( .A1(n38234), .A2(n38233), .ZN(n38232) );
  NOR2_X1 U784 ( .A1(n35403), .A2(n37373), .ZN(n37694) );
  NAND2_X1 U787 ( .A1(n37133), .A2(n38393), .ZN(n5264) );
  NOR2_X1 U789 ( .A1(n9058), .A2(n15352), .ZN(n37735) );
  NAND2_X1 U792 ( .A1(n26755), .A2(n38268), .ZN(n32917) );
  NAND2_X1 U798 ( .A1(n38955), .A2(n6261), .ZN(n31406) );
  NAND2_X1 U802 ( .A1(n38498), .A2(n4489), .ZN(n30689) );
  OAI21_X1 U803 ( .A1(n14458), .A2(n39342), .B(n7596), .ZN(n3283) );
  NAND2_X1 U804 ( .A1(n10736), .A2(n26695), .ZN(n32928) );
  OAI21_X1 U805 ( .A1(n26661), .A2(n19449), .B(n16773), .ZN(n3282) );
  AOI21_X1 U807 ( .A1(n26799), .A2(n39514), .B(n18773), .ZN(n9240) );
  NAND2_X1 U809 ( .A1(n7619), .A2(n1235), .ZN(n10567) );
  NAND2_X1 U815 ( .A1(n4007), .A2(n33352), .ZN(n30643) );
  NAND2_X1 U817 ( .A1(n26618), .A2(n31701), .ZN(n20604) );
  AOI21_X1 U818 ( .A1(n875), .A2(n26937), .B(n11334), .ZN(n37549) );
  NAND2_X1 U824 ( .A1(n26459), .A2(n735), .ZN(n9166) );
  NOR2_X1 U828 ( .A1(n1231), .A2(n30665), .ZN(n26624) );
  AND2_X1 U838 ( .A1(n849), .A2(n9178), .Z(n37074) );
  NAND2_X1 U844 ( .A1(n33063), .A2(n33062), .ZN(n37766) );
  NAND2_X1 U847 ( .A1(n38715), .A2(n16941), .ZN(n39222) );
  OAI21_X1 U848 ( .A1(n11325), .A2(n4970), .B(n1093), .ZN(n38498) );
  INV_X1 U850 ( .I(n11334), .ZN(n38824) );
  NAND2_X1 U851 ( .A1(n26944), .A2(n26849), .ZN(n38393) );
  INV_X1 U853 ( .I(n26943), .ZN(n36146) );
  OAI21_X1 U864 ( .A1(n278), .A2(n1786), .B(n8917), .ZN(n37562) );
  NOR2_X1 U867 ( .A1(n26639), .A2(n862), .ZN(n37286) );
  INV_X1 U872 ( .I(n37288), .ZN(n37287) );
  NAND2_X1 U873 ( .A1(n17047), .A2(n6615), .ZN(n38684) );
  NAND2_X1 U875 ( .A1(n11248), .A2(n26910), .ZN(n38549) );
  OAI21_X1 U878 ( .A1(n5935), .A2(n19331), .B(n15998), .ZN(n39646) );
  NOR3_X1 U879 ( .A1(n13686), .A2(n5960), .A3(n14080), .ZN(n5963) );
  AOI22_X1 U880 ( .A1(n21192), .A2(n26826), .B1(n26769), .B2(n14488), .ZN(
        n39557) );
  NAND2_X1 U882 ( .A1(n39758), .A2(n26923), .ZN(n39508) );
  NOR2_X1 U884 ( .A1(n13854), .A2(n13088), .ZN(n38233) );
  AOI21_X1 U885 ( .A1(n278), .A2(n1786), .B(n8415), .ZN(n34601) );
  NAND3_X1 U888 ( .A1(n26991), .A2(n26989), .A3(n26990), .ZN(n5477) );
  NAND3_X1 U891 ( .A1(n11616), .A2(n38644), .A3(n10231), .ZN(n38268) );
  AND2_X1 U895 ( .A1(n20321), .A2(n37084), .Z(n2929) );
  AND2_X1 U901 ( .A1(n11636), .A2(n38280), .Z(n26777) );
  AND2_X1 U910 ( .A1(n15037), .A2(n35256), .Z(n2491) );
  INV_X1 U918 ( .I(n860), .ZN(n37955) );
  NOR2_X1 U926 ( .A1(n32345), .A2(n20211), .ZN(n3935) );
  NOR2_X1 U927 ( .A1(n33279), .A2(n32168), .ZN(n37281) );
  BUF_X2 U928 ( .I(n26704), .Z(n7978) );
  NOR2_X1 U932 ( .A1(n441), .A2(n26639), .ZN(n34108) );
  OR2_X1 U937 ( .A1(n875), .A2(n17993), .Z(n37154) );
  NOR2_X1 U941 ( .A1(n2451), .A2(n26639), .ZN(n12236) );
  OR2_X1 U953 ( .A1(n26932), .A2(n37235), .Z(n17617) );
  AOI21_X1 U955 ( .A1(n862), .A2(n9690), .B(n37289), .ZN(n37288) );
  INV_X1 U956 ( .I(n33455), .ZN(n9081) );
  INV_X1 U958 ( .I(n9801), .ZN(n38591) );
  INV_X1 U969 ( .I(n19728), .ZN(n38592) );
  INV_X1 U971 ( .I(n859), .ZN(n36477) );
  INV_X1 U973 ( .I(n13528), .ZN(n37856) );
  INV_X1 U974 ( .I(n26704), .ZN(n6190) );
  OR2_X1 U980 ( .A1(n18390), .A2(n31897), .Z(n35622) );
  INV_X1 U984 ( .I(n26988), .ZN(n26819) );
  CLKBUF_X2 U986 ( .I(n5274), .Z(n33352) );
  OR2_X1 U988 ( .A1(n20321), .A2(n37084), .Z(n26667) );
  NAND2_X1 U989 ( .A1(n30859), .A2(n26988), .ZN(n26606) );
  INV_X1 U990 ( .I(n36355), .ZN(n36873) );
  INV_X1 U992 ( .I(n36931), .ZN(n30284) );
  INV_X1 U997 ( .I(n39353), .ZN(n36355) );
  INV_X1 U998 ( .I(n39207), .ZN(n39825) );
  INV_X1 U1001 ( .I(n37588), .ZN(n6454) );
  INV_X1 U1003 ( .I(n26511), .ZN(n39561) );
  BUF_X2 U1006 ( .I(n32253), .Z(n38844) );
  CLKBUF_X2 U1007 ( .I(n31965), .Z(n36758) );
  INV_X1 U1008 ( .I(n26420), .ZN(n3330) );
  INV_X1 U1011 ( .I(n13853), .ZN(n26451) );
  INV_X1 U1015 ( .I(n26356), .ZN(n33504) );
  BUF_X2 U1017 ( .I(n10076), .Z(n39129) );
  INV_X2 U1021 ( .I(n26517), .ZN(n39662) );
  AOI21_X1 U1024 ( .A1(n26236), .A2(n26237), .B(n30883), .ZN(n26240) );
  NOR2_X1 U1030 ( .A1(n25785), .A2(n30595), .ZN(n10457) );
  AOI21_X1 U1033 ( .A1(n38953), .A2(n10724), .B(n13869), .ZN(n11424) );
  INV_X1 U1035 ( .I(n6989), .ZN(n39135) );
  NOR2_X1 U1039 ( .A1(n38437), .A2(n8407), .ZN(n13121) );
  NAND2_X1 U1042 ( .A1(n37745), .A2(n38501), .ZN(n32380) );
  OAI21_X1 U1047 ( .A1(n20235), .A2(n25800), .B(n17951), .ZN(n37618) );
  NOR2_X1 U1050 ( .A1(n34339), .A2(n12910), .ZN(n38386) );
  NOR2_X1 U1051 ( .A1(n16867), .A2(n25965), .ZN(n2837) );
  NAND2_X1 U1057 ( .A1(n16977), .A2(n37996), .ZN(n25918) );
  NAND3_X1 U1060 ( .A1(n1098), .A2(n38409), .A3(n26119), .ZN(n20062) );
  NAND2_X1 U1071 ( .A1(n3518), .A2(n26084), .ZN(n10270) );
  NAND2_X1 U1076 ( .A1(n32243), .A2(n18354), .ZN(n18353) );
  OAI21_X1 U1078 ( .A1(n14650), .A2(n25978), .B(n31496), .ZN(n37365) );
  NAND3_X1 U1079 ( .A1(n25764), .A2(n13869), .A3(n34217), .ZN(n30571) );
  AOI22_X1 U1088 ( .A1(n1515), .A2(n7460), .B1(n8005), .B2(n1240), .ZN(n34554)
         );
  AOI22_X1 U1090 ( .A1(n25788), .A2(n1514), .B1(n17371), .B2(n17372), .ZN(
        n13389) );
  INV_X1 U1111 ( .I(n9859), .ZN(n25886) );
  INV_X1 U1116 ( .I(n34399), .ZN(n37416) );
  INV_X1 U1118 ( .I(n37462), .ZN(n34117) );
  NOR2_X1 U1122 ( .A1(n25836), .A2(n3213), .ZN(n25861) );
  NAND2_X1 U1125 ( .A1(n35151), .A2(n18661), .ZN(n26111) );
  BUF_X2 U1129 ( .I(n7512), .Z(n32243) );
  NOR2_X1 U1146 ( .A1(n15832), .A2(n15831), .ZN(n39509) );
  AOI22_X1 U1147 ( .A1(n11552), .A2(n25993), .B1(n25956), .B2(n9413), .ZN(
        n25510) );
  INV_X1 U1148 ( .I(n31624), .ZN(n3518) );
  CLKBUF_X2 U1149 ( .I(n9802), .Z(n33218) );
  NAND2_X1 U1151 ( .A1(n32924), .A2(n38432), .ZN(n33764) );
  AND2_X1 U1158 ( .A1(n26125), .A2(n39454), .Z(n4191) );
  NAND2_X1 U1159 ( .A1(n38437), .A2(n26041), .ZN(n34254) );
  NAND2_X1 U1165 ( .A1(n39030), .A2(n32690), .ZN(n25910) );
  NAND2_X1 U1166 ( .A1(n10223), .A2(n10764), .ZN(n7915) );
  OR2_X1 U1172 ( .A1(n26015), .A2(n25801), .Z(n26121) );
  NOR2_X1 U1176 ( .A1(n26120), .A2(n25903), .ZN(n39143) );
  OAI21_X1 U1184 ( .A1(n25978), .A2(n1100), .B(n34265), .ZN(n37930) );
  OAI22_X1 U1191 ( .A1(n1523), .A2(n25868), .B1(n26021), .B2(n1524), .ZN(
        n13440) );
  AND2_X1 U1195 ( .A1(n6904), .A2(n26124), .Z(n37072) );
  BUF_X2 U1196 ( .I(n26048), .Z(n1523) );
  INV_X2 U1197 ( .I(n35003), .ZN(n13869) );
  INV_X2 U1212 ( .I(n3575), .ZN(n6222) );
  NOR3_X1 U1214 ( .A1(n37683), .A2(n1012), .A3(n25992), .ZN(n8233) );
  BUF_X2 U1216 ( .I(n14890), .Z(n4163) );
  CLKBUF_X4 U1219 ( .I(n10986), .Z(n446) );
  NAND2_X1 U1220 ( .A1(n25989), .A2(n34217), .ZN(n38550) );
  INV_X1 U1224 ( .I(n598), .ZN(n1018) );
  CLKBUF_X4 U1226 ( .I(n6904), .Z(n4602) );
  NAND2_X1 U1227 ( .A1(n32196), .A2(n20813), .ZN(n38509) );
  NAND2_X1 U1229 ( .A1(n951), .A2(n13712), .ZN(n32558) );
  INV_X2 U1236 ( .I(n26134), .ZN(n1105) );
  NAND2_X1 U1238 ( .A1(n37393), .A2(n17212), .ZN(n17211) );
  INV_X1 U1241 ( .I(n34350), .ZN(n10404) );
  NAND2_X1 U1243 ( .A1(n38663), .A2(n39782), .ZN(n38185) );
  NAND2_X1 U1247 ( .A1(n12548), .A2(n25798), .ZN(n25856) );
  BUF_X2 U1249 ( .I(n10015), .Z(n32196) );
  CLKBUF_X2 U1251 ( .I(n598), .Z(n38247) );
  INV_X2 U1252 ( .I(n6830), .ZN(n6390) );
  CLKBUF_X2 U1253 ( .I(n25801), .Z(n7423) );
  AOI22_X1 U1257 ( .A1(n25541), .A2(n36486), .B1(n5042), .B2(n25542), .ZN(
        n39782) );
  NOR2_X1 U1260 ( .A1(n38675), .A2(n13301), .ZN(n37596) );
  OAI21_X1 U1272 ( .A1(n39390), .A2(n37174), .B(n11951), .ZN(n32827) );
  OAI21_X1 U1274 ( .A1(n33597), .A2(n25364), .B(n37905), .ZN(n38662) );
  NOR2_X1 U1279 ( .A1(n25697), .A2(n37119), .ZN(n16230) );
  OAI21_X1 U1283 ( .A1(n25622), .A2(n25365), .B(n33114), .ZN(n7890) );
  NAND2_X1 U1289 ( .A1(n33268), .A2(n25248), .ZN(n9146) );
  AND2_X1 U1291 ( .A1(n25699), .A2(n31721), .Z(n37181) );
  NOR2_X1 U1292 ( .A1(n39327), .A2(n30317), .ZN(n38675) );
  AND2_X1 U1293 ( .A1(n14401), .A2(n19863), .Z(n34099) );
  OAI21_X1 U1295 ( .A1(n32076), .A2(n2149), .B(n1530), .ZN(n39144) );
  AND2_X1 U1296 ( .A1(n25577), .A2(n1109), .Z(n37174) );
  NOR2_X1 U1301 ( .A1(n37336), .A2(n19767), .ZN(n36020) );
  OAI21_X1 U1302 ( .A1(n25448), .A2(n25583), .B(n38782), .ZN(n38004) );
  AND2_X1 U1316 ( .A1(n15515), .A2(n32026), .Z(n25525) );
  NAND2_X1 U1317 ( .A1(n7926), .A2(n36345), .ZN(n39352) );
  NOR2_X1 U1320 ( .A1(n10158), .A2(n7284), .ZN(n16410) );
  OAI21_X1 U1321 ( .A1(n31721), .A2(n25699), .B(n12931), .ZN(n5034) );
  NOR2_X1 U1324 ( .A1(n25381), .A2(n1109), .ZN(n39390) );
  NOR3_X1 U1327 ( .A1(n15443), .A2(n11150), .A3(n14553), .ZN(n15422) );
  OAI21_X1 U1328 ( .A1(n19336), .A2(n25248), .B(n12896), .ZN(n37647) );
  OAI21_X1 U1337 ( .A1(n6747), .A2(n20441), .B(n38223), .ZN(n9336) );
  NAND2_X1 U1340 ( .A1(n25682), .A2(n25681), .ZN(n19490) );
  INV_X1 U1343 ( .I(n25489), .ZN(n38364) );
  OR2_X1 U1345 ( .A1(n13413), .A2(n11060), .Z(n16315) );
  OR2_X1 U1353 ( .A1(n19941), .A2(n24896), .Z(n20296) );
  BUF_X2 U1354 ( .I(n25513), .Z(n39327) );
  NAND2_X1 U1358 ( .A1(n1551), .A2(n371), .ZN(n14805) );
  CLKBUF_X2 U1360 ( .I(n25359), .Z(n39321) );
  CLKBUF_X2 U1366 ( .I(n25619), .Z(n9594) );
  CLKBUF_X1 U1370 ( .I(n24741), .Z(n36249) );
  NOR2_X1 U1372 ( .A1(n10055), .A2(n6300), .ZN(n4824) );
  NOR2_X1 U1374 ( .A1(n33114), .A2(n33384), .ZN(n33113) );
  OAI21_X1 U1375 ( .A1(n25142), .A2(n20924), .B(n37844), .ZN(n39568) );
  NAND2_X1 U1397 ( .A1(n37845), .A2(n38782), .ZN(n4217) );
  NOR2_X1 U1400 ( .A1(n20924), .A2(n11874), .ZN(n11873) );
  NAND2_X1 U1404 ( .A1(n9132), .A2(n37051), .ZN(n2462) );
  NAND2_X1 U1410 ( .A1(n25674), .A2(n25677), .ZN(n39700) );
  NAND3_X1 U1415 ( .A1(n6065), .A2(n32450), .A3(n1252), .ZN(n35710) );
  AOI21_X1 U1416 ( .A1(n25600), .A2(n33491), .B(n25601), .ZN(n37348) );
  INV_X1 U1417 ( .I(n32989), .ZN(n19678) );
  INV_X1 U1418 ( .I(n33491), .ZN(n34755) );
  INV_X1 U1421 ( .I(n38849), .ZN(n18545) );
  INV_X1 U1422 ( .I(n32775), .ZN(n20815) );
  CLKBUF_X2 U1423 ( .I(n31669), .Z(n39160) );
  CLKBUF_X2 U1425 ( .I(n19941), .Z(n39371) );
  AND2_X1 U1433 ( .A1(n20595), .A2(n19696), .Z(n34060) );
  NAND2_X1 U1434 ( .A1(n12944), .A2(n20924), .ZN(n37844) );
  BUF_X2 U1435 ( .I(n32989), .Z(n5166) );
  INV_X1 U1439 ( .I(n25619), .ZN(n11874) );
  NOR2_X1 U1447 ( .A1(n25449), .A2(n25582), .ZN(n37845) );
  NOR2_X1 U1448 ( .A1(n1548), .A2(n17774), .ZN(n15620) );
  INV_X1 U1449 ( .I(n39778), .ZN(n34150) );
  INV_X1 U1450 ( .I(n25072), .ZN(n5800) );
  INV_X1 U1451 ( .I(n25254), .ZN(n20347) );
  INV_X1 U1452 ( .I(n15930), .ZN(n25250) );
  CLKBUF_X2 U1457 ( .I(n25136), .Z(n39756) );
  INV_X1 U1460 ( .I(n13935), .ZN(n6984) );
  INV_X1 U1480 ( .I(n25237), .ZN(n39582) );
  INV_X2 U1482 ( .I(n25259), .ZN(n1260) );
  INV_X1 U1483 ( .I(n9701), .ZN(n38336) );
  NAND2_X1 U1487 ( .A1(n38242), .A2(n2505), .ZN(n2503) );
  INV_X1 U1488 ( .I(n25079), .ZN(n25258) );
  OAI21_X1 U1502 ( .A1(n33317), .A2(n37115), .B(n38521), .ZN(n20665) );
  NAND2_X1 U1509 ( .A1(n39469), .A2(n33666), .ZN(n38083) );
  CLKBUF_X2 U1511 ( .I(n36908), .Z(n36228) );
  CLKBUF_X2 U1513 ( .I(n20411), .Z(n39157) );
  NOR2_X1 U1514 ( .A1(n31698), .A2(n39704), .ZN(n33449) );
  AOI21_X1 U1521 ( .A1(n31213), .A2(n37355), .B(n24655), .ZN(n24657) );
  NOR2_X1 U1526 ( .A1(n24789), .A2(n20039), .ZN(n37830) );
  NAND2_X1 U1542 ( .A1(n33317), .A2(n24899), .ZN(n38521) );
  NAND2_X1 U1544 ( .A1(n957), .A2(n31845), .ZN(n15585) );
  AND2_X1 U1547 ( .A1(n2731), .A2(n24674), .Z(n37202) );
  NOR2_X1 U1548 ( .A1(n19886), .A2(n24565), .ZN(n39712) );
  NAND2_X1 U1549 ( .A1(n6791), .A2(n1784), .ZN(n1783) );
  AND2_X1 U1550 ( .A1(n24715), .A2(n39268), .Z(n16908) );
  AOI21_X1 U1555 ( .A1(n24909), .A2(n36634), .B(n36752), .ZN(n6229) );
  NOR2_X1 U1562 ( .A1(n31198), .A2(n3697), .ZN(n37684) );
  NOR2_X1 U1564 ( .A1(n1120), .A2(n36082), .ZN(n24765) );
  NAND2_X1 U1568 ( .A1(n38978), .A2(n8264), .ZN(n33401) );
  NAND2_X1 U1570 ( .A1(n39817), .A2(n5888), .ZN(n9071) );
  INV_X1 U1574 ( .I(n34141), .ZN(n38293) );
  NOR2_X1 U1580 ( .A1(n31861), .A2(n38182), .ZN(n20944) );
  NOR3_X1 U1582 ( .A1(n24775), .A2(n24292), .A3(n35801), .ZN(n4578) );
  NAND2_X1 U1586 ( .A1(n5063), .A2(n37474), .ZN(n38286) );
  NOR2_X1 U1591 ( .A1(n39085), .A2(n37276), .ZN(n37275) );
  NOR2_X1 U1597 ( .A1(n9197), .A2(n9198), .ZN(n30384) );
  NAND2_X1 U1600 ( .A1(n2731), .A2(n15282), .ZN(n38795) );
  OAI21_X1 U1606 ( .A1(n36988), .A2(n24648), .B(n37477), .ZN(n24514) );
  AOI21_X1 U1612 ( .A1(n31385), .A2(n24866), .B(n30554), .ZN(n7970) );
  NOR2_X1 U1618 ( .A1(n16210), .A2(n18110), .ZN(n16949) );
  NOR2_X1 U1619 ( .A1(n24899), .A2(n1268), .ZN(n35170) );
  NOR3_X1 U1620 ( .A1(n9921), .A2(n24685), .A3(n24686), .ZN(n815) );
  INV_X1 U1623 ( .I(n24572), .ZN(n16208) );
  NAND2_X1 U1625 ( .A1(n24529), .A2(n5897), .ZN(n13050) );
  NAND3_X1 U1633 ( .A1(n34662), .A2(n16815), .A3(n37395), .ZN(n38389) );
  CLKBUF_X2 U1637 ( .I(n39098), .Z(n38984) );
  INV_X1 U1641 ( .I(n24712), .ZN(n24899) );
  INV_X1 U1642 ( .I(n39279), .ZN(n30699) );
  INV_X1 U1644 ( .I(n10054), .ZN(n14857) );
  INV_X2 U1652 ( .I(n14283), .ZN(n1121) );
  INV_X1 U1654 ( .I(n35250), .ZN(n16815) );
  NAND2_X1 U1656 ( .A1(n35443), .A2(n24650), .ZN(n24868) );
  INV_X2 U1660 ( .I(n37477), .ZN(n14241) );
  BUF_X2 U1667 ( .I(n5634), .Z(n37737) );
  BUF_X2 U1668 ( .I(n2616), .Z(n31213) );
  NAND2_X1 U1677 ( .A1(n24811), .A2(n37277), .ZN(n37276) );
  INV_X1 U1678 ( .I(n24227), .ZN(n38744) );
  CLKBUF_X2 U1680 ( .I(n32637), .Z(n39085) );
  NOR2_X1 U1681 ( .A1(n7871), .A2(n1577), .ZN(n37318) );
  INV_X2 U1686 ( .I(n3510), .ZN(n36752) );
  NOR2_X1 U1690 ( .A1(n36716), .A2(n5768), .ZN(n6744) );
  NOR2_X1 U1691 ( .A1(n24875), .A2(n24876), .ZN(n36017) );
  AOI21_X1 U1694 ( .A1(n24829), .A2(n14064), .B(n13665), .ZN(n13666) );
  NOR2_X1 U1703 ( .A1(n24565), .A2(n32637), .ZN(n24528) );
  AOI21_X1 U1708 ( .A1(n24592), .A2(n24847), .B(n35960), .ZN(n24593) );
  NAND2_X1 U1710 ( .A1(n23857), .A2(n31845), .ZN(n37537) );
  NAND2_X1 U1714 ( .A1(n24855), .A2(n35373), .ZN(n24856) );
  INV_X2 U1716 ( .I(n39406), .ZN(n9198) );
  NAND2_X1 U1718 ( .A1(n39523), .A2(n36395), .ZN(n24897) );
  NOR2_X1 U1720 ( .A1(n38658), .A2(n24783), .ZN(n24177) );
  NOR2_X1 U1724 ( .A1(n8317), .A2(n31385), .ZN(n31483) );
  OR2_X1 U1725 ( .A1(n5282), .A2(n38749), .Z(n32390) );
  INV_X1 U1727 ( .I(n39098), .ZN(n18324) );
  NOR2_X1 U1731 ( .A1(n31796), .A2(n38848), .ZN(n39265) );
  AOI21_X1 U1733 ( .A1(n31845), .A2(n1574), .B(n1026), .ZN(n10403) );
  NAND2_X1 U1740 ( .A1(n7810), .A2(n32831), .ZN(n38978) );
  INV_X1 U1746 ( .I(n32651), .ZN(n37277) );
  INV_X1 U1747 ( .I(n30845), .ZN(n24820) );
  INV_X1 U1750 ( .I(n15414), .ZN(n13665) );
  INV_X1 U1751 ( .I(n36908), .ZN(n38973) );
  BUF_X2 U1758 ( .I(n14729), .Z(n7286) );
  BUF_X2 U1760 ( .I(n24827), .Z(n5431) );
  BUF_X4 U1765 ( .I(n24817), .Z(n37106) );
  NAND2_X1 U1766 ( .A1(n19420), .A2(n36385), .ZN(n7871) );
  NOR2_X1 U1773 ( .A1(n1120), .A2(n39098), .ZN(n18168) );
  BUF_X2 U1779 ( .I(n18788), .Z(n9997) );
  NAND2_X1 U1780 ( .A1(n24674), .A2(n15281), .ZN(n24226) );
  NAND2_X1 U1782 ( .A1(n24746), .A2(n39279), .ZN(n24602) );
  OAI21_X1 U1786 ( .A1(n12250), .A2(n12277), .B(n19915), .ZN(n12249) );
  BUF_X4 U1789 ( .I(n32136), .Z(n37097) );
  NOR2_X1 U1799 ( .A1(n5957), .A2(n3760), .ZN(n5495) );
  OR2_X1 U1800 ( .A1(n1125), .A2(n9371), .Z(n37065) );
  OR2_X1 U1802 ( .A1(n24098), .A2(n24403), .Z(n2342) );
  NOR2_X1 U1803 ( .A1(n39398), .A2(n39397), .ZN(n39244) );
  AOI22_X1 U1805 ( .A1(n37068), .A2(n1128), .B1(n1588), .B2(n2579), .ZN(n38036) );
  NAND2_X1 U1810 ( .A1(n24140), .A2(n2336), .ZN(n31267) );
  NOR2_X1 U1816 ( .A1(n4308), .A2(n32818), .ZN(n37977) );
  NAND2_X1 U1818 ( .A1(n36740), .A2(n24234), .ZN(n38821) );
  NAND2_X1 U1819 ( .A1(n39381), .A2(n33531), .ZN(n39243) );
  AOI21_X1 U1820 ( .A1(n24395), .A2(n24182), .B(n19739), .ZN(n38526) );
  NOR2_X1 U1821 ( .A1(n250), .A2(n24443), .ZN(n24441) );
  INV_X1 U1822 ( .I(n35314), .ZN(n39397) );
  OAI21_X1 U1832 ( .A1(n8987), .A2(n24219), .B(n1124), .ZN(n37388) );
  NOR2_X1 U1839 ( .A1(n5853), .A2(n31464), .ZN(n37672) );
  NOR2_X1 U1840 ( .A1(n9101), .A2(n1131), .ZN(n38405) );
  NAND2_X1 U1841 ( .A1(n34422), .A2(n33531), .ZN(n15365) );
  INV_X1 U1845 ( .I(n32683), .ZN(n39398) );
  OR2_X1 U1848 ( .A1(n1130), .A2(n7240), .Z(n37068) );
  INV_X1 U1849 ( .I(n35954), .ZN(n35958) );
  OR2_X1 U1850 ( .A1(n1276), .A2(n15385), .Z(n19381) );
  INV_X1 U1851 ( .I(n6715), .ZN(n38422) );
  NOR2_X1 U1852 ( .A1(n24401), .A2(n14392), .ZN(n24402) );
  NAND2_X1 U1854 ( .A1(n33104), .A2(n24258), .ZN(n24378) );
  AOI22_X1 U1859 ( .A1(n10220), .A2(n15049), .B1(n1131), .B2(n19140), .ZN(
        n38446) );
  NOR2_X1 U1862 ( .A1(n24382), .A2(n24381), .ZN(n17067) );
  OAI22_X1 U1863 ( .A1(n39156), .A2(n35916), .B1(n24345), .B2(n20404), .ZN(
        n24350) );
  NOR2_X1 U1864 ( .A1(n11361), .A2(n24141), .ZN(n2989) );
  NAND2_X1 U1865 ( .A1(n24225), .A2(n16081), .ZN(n37958) );
  AOI22_X1 U1866 ( .A1(n24331), .A2(n24327), .B1(n24174), .B2(n39057), .ZN(
        n36640) );
  NAND2_X1 U1868 ( .A1(n24484), .A2(n24241), .ZN(n24345) );
  NAND2_X1 U1879 ( .A1(n1131), .A2(n2597), .ZN(n4702) );
  INV_X1 U1881 ( .I(n24433), .ZN(n15240) );
  AND2_X1 U1885 ( .A1(n35233), .A2(n15903), .Z(n24207) );
  AND2_X1 U1889 ( .A1(n12759), .A2(n12758), .Z(n24231) );
  INV_X1 U1890 ( .I(n24216), .ZN(n38527) );
  NOR2_X1 U1891 ( .A1(n14655), .A2(n15751), .ZN(n12926) );
  NAND2_X1 U1892 ( .A1(n32683), .A2(n33580), .ZN(n24261) );
  CLKBUF_X2 U1894 ( .I(n17693), .Z(n37377) );
  INV_X2 U1896 ( .I(n2192), .ZN(n39373) );
  NAND2_X1 U1907 ( .A1(n24328), .A2(n1589), .ZN(n15146) );
  NAND3_X1 U1917 ( .A1(n2439), .A2(n24458), .A3(n38431), .ZN(n32881) );
  NAND2_X1 U1930 ( .A1(n24169), .A2(n20457), .ZN(n24397) );
  NOR2_X1 U1931 ( .A1(n33314), .A2(n20196), .ZN(n20989) );
  OR2_X1 U1932 ( .A1(n20619), .A2(n24470), .Z(n24132) );
  NAND2_X1 U1934 ( .A1(n16449), .A2(n1283), .ZN(n23820) );
  NAND2_X1 U1939 ( .A1(n35450), .A2(n37267), .ZN(n24133) );
  INV_X1 U1941 ( .I(n30494), .ZN(n1289) );
  NAND2_X1 U1943 ( .A1(n1129), .A2(n24360), .ZN(n24457) );
  CLKBUF_X1 U1944 ( .I(n6226), .Z(n34786) );
  NOR2_X1 U1948 ( .A1(n2395), .A2(n1589), .ZN(n38948) );
  BUF_X2 U1951 ( .I(n33599), .Z(n39605) );
  INV_X1 U1952 ( .I(n35242), .ZN(n39055) );
  INV_X1 U1959 ( .I(n23598), .ZN(n36067) );
  INV_X1 U1960 ( .I(n23775), .ZN(n38022) );
  INV_X1 U1961 ( .I(n20205), .ZN(n39314) );
  CLKBUF_X4 U1965 ( .I(n39161), .Z(n38021) );
  INV_X1 U1968 ( .I(n24034), .ZN(n37861) );
  OAI21_X1 U1972 ( .A1(n23600), .A2(n12597), .B(n37649), .ZN(n14107) );
  BUF_X2 U1980 ( .I(n23419), .Z(n39408) );
  NAND2_X1 U1981 ( .A1(n3506), .A2(n23561), .ZN(n1830) );
  AOI21_X1 U1996 ( .A1(n37278), .A2(n17927), .B(n23625), .ZN(n17926) );
  OAI21_X1 U1998 ( .A1(n16715), .A2(n23455), .B(n605), .ZN(n33155) );
  INV_X1 U1999 ( .I(n23939), .ZN(n39412) );
  INV_X1 U2003 ( .I(n23636), .ZN(n23640) );
  INV_X1 U2005 ( .I(n23460), .ZN(n37005) );
  NOR2_X1 U2011 ( .A1(n23521), .A2(n2273), .ZN(n9672) );
  INV_X2 U2019 ( .I(n23430), .ZN(n37279) );
  NAND2_X1 U2020 ( .A1(n33869), .A2(n38806), .ZN(n18538) );
  NAND2_X1 U2022 ( .A1(n37528), .A2(n30506), .ZN(n32596) );
  NOR2_X1 U2026 ( .A1(n38335), .A2(n38334), .ZN(n35398) );
  NOR2_X1 U2029 ( .A1(n23522), .A2(n2273), .ZN(n23405) );
  NOR2_X1 U2031 ( .A1(n16728), .A2(n2798), .ZN(n39281) );
  OR2_X1 U2033 ( .A1(n23272), .A2(n36564), .Z(n15603) );
  AND2_X1 U2043 ( .A1(n33786), .A2(n10216), .Z(n7886) );
  NAND2_X1 U2046 ( .A1(n23401), .A2(n32471), .ZN(n20867) );
  NOR2_X1 U2052 ( .A1(n39805), .A2(n17768), .ZN(n37482) );
  NAND2_X1 U2055 ( .A1(n39012), .A2(n23283), .ZN(n33911) );
  OAI21_X1 U2056 ( .A1(n37207), .A2(n36448), .B(n37802), .ZN(n23648) );
  NOR2_X1 U2059 ( .A1(n37839), .A2(n16726), .ZN(n34942) );
  NOR2_X1 U2061 ( .A1(n21130), .A2(n38380), .ZN(n23393) );
  NAND2_X1 U2062 ( .A1(n15458), .A2(n1644), .ZN(n37320) );
  NAND2_X1 U2067 ( .A1(n23302), .A2(n12597), .ZN(n37649) );
  NOR2_X1 U2070 ( .A1(n17995), .A2(n39133), .ZN(n37976) );
  INV_X1 U2074 ( .I(n23453), .ZN(n16715) );
  AND2_X1 U2075 ( .A1(n35938), .A2(n23430), .Z(n37278) );
  NOR2_X1 U2077 ( .A1(n3174), .A2(n32061), .ZN(n32060) );
  NAND2_X1 U2080 ( .A1(n23116), .A2(n23117), .ZN(n23335) );
  OAI21_X1 U2085 ( .A1(n11097), .A2(n20031), .B(n1036), .ZN(n39276) );
  NOR2_X1 U2086 ( .A1(n1136), .A2(n38248), .ZN(n37569) );
  OAI21_X1 U2087 ( .A1(n4859), .A2(n1642), .B(n23392), .ZN(n6052) );
  AND2_X1 U2090 ( .A1(n23531), .A2(n33453), .Z(n39812) );
  INV_X1 U2092 ( .I(n23505), .ZN(n39301) );
  INV_X1 U2105 ( .I(n23568), .ZN(n1298) );
  AND2_X1 U2107 ( .A1(n23440), .A2(n9862), .Z(n2454) );
  NOR2_X1 U2109 ( .A1(n23459), .A2(n35808), .ZN(n36431) );
  NOR3_X1 U2114 ( .A1(n31685), .A2(n18086), .A3(n36539), .ZN(n4396) );
  CLKBUF_X2 U2115 ( .I(n4618), .Z(n32351) );
  NOR2_X1 U2122 ( .A1(n7379), .A2(n10143), .ZN(n18391) );
  NAND2_X1 U2133 ( .A1(n5044), .A2(n6159), .ZN(n23574) );
  NAND2_X1 U2135 ( .A1(n23401), .A2(n33703), .ZN(n22872) );
  NOR2_X1 U2136 ( .A1(n39803), .A2(n9772), .ZN(n39428) );
  CLKBUF_X2 U2143 ( .I(n23577), .Z(n39214) );
  BUF_X2 U2144 ( .I(n3708), .Z(n36103) );
  CLKBUF_X2 U2145 ( .I(n23518), .Z(n38252) );
  NOR2_X1 U2148 ( .A1(n23645), .A2(n37839), .ZN(n30417) );
  NOR2_X1 U2150 ( .A1(n23460), .A2(n23458), .ZN(n36430) );
  NAND2_X1 U2156 ( .A1(n23360), .A2(n14974), .ZN(n37779) );
  NAND2_X1 U2157 ( .A1(n22680), .A2(n22681), .ZN(n37514) );
  NAND2_X1 U2163 ( .A1(n23611), .A2(n4525), .ZN(n38651) );
  NAND2_X1 U2165 ( .A1(n1634), .A2(n38614), .ZN(n11436) );
  INV_X2 U2169 ( .I(n23580), .ZN(n1138) );
  NAND2_X1 U2170 ( .A1(n23620), .A2(n16774), .ZN(n38971) );
  NOR2_X1 U2180 ( .A1(n1299), .A2(n39001), .ZN(n7048) );
  INV_X1 U2184 ( .I(n38792), .ZN(n20278) );
  AND2_X1 U2185 ( .A1(n12966), .A2(n9862), .Z(n23282) );
  NOR2_X1 U2187 ( .A1(n15353), .A2(n8692), .ZN(n32111) );
  NAND2_X1 U2192 ( .A1(n23637), .A2(n12028), .ZN(n23247) );
  BUF_X2 U2195 ( .I(n7644), .Z(n32930) );
  AND2_X1 U2196 ( .A1(n8660), .A2(n38704), .Z(n23412) );
  CLKBUF_X2 U2198 ( .I(n35331), .Z(n39316) );
  INV_X1 U2204 ( .I(n38614), .ZN(n23346) );
  NOR2_X1 U2209 ( .A1(n38441), .A2(n39070), .ZN(n23556) );
  INV_X2 U2219 ( .I(n33747), .ZN(n23571) );
  INV_X2 U2224 ( .I(n23337), .ZN(n31331) );
  NAND2_X1 U2226 ( .A1(n17931), .A2(n13029), .ZN(n23272) );
  NAND2_X1 U2227 ( .A1(n23456), .A2(n2553), .ZN(n15941) );
  NOR2_X1 U2231 ( .A1(n30574), .A2(n2553), .ZN(n38792) );
  CLKBUF_X2 U2234 ( .I(n10216), .Z(n8190) );
  NAND2_X1 U2235 ( .A1(n19559), .A2(n23487), .ZN(n36551) );
  INV_X2 U2237 ( .I(n39001), .ZN(n7049) );
  INV_X1 U2238 ( .I(n23296), .ZN(n37308) );
  CLKBUF_X2 U2240 ( .I(n33840), .Z(n39805) );
  AOI21_X1 U2244 ( .A1(n33082), .A2(n22907), .B(n22906), .ZN(n38173) );
  INV_X2 U2250 ( .I(n13733), .ZN(n37774) );
  INV_X2 U2251 ( .I(n37088), .ZN(n23389) );
  CLKBUF_X2 U2252 ( .I(n30299), .Z(n38119) );
  BUF_X4 U2253 ( .I(n20346), .Z(n39401) );
  NOR2_X1 U2256 ( .A1(n35950), .A2(n37063), .ZN(n34615) );
  NAND2_X1 U2259 ( .A1(n19481), .A2(n35534), .ZN(n9856) );
  INV_X1 U2264 ( .I(n16094), .ZN(n21293) );
  NAND2_X1 U2268 ( .A1(n23160), .A2(n38074), .ZN(n32909) );
  NAND2_X1 U2269 ( .A1(n22830), .A2(n22831), .ZN(n37980) );
  OAI21_X1 U2272 ( .A1(n23162), .A2(n22871), .B(n22915), .ZN(n37548) );
  OAI22_X1 U2273 ( .A1(n4714), .A2(n36736), .B1(n1144), .B2(n8730), .ZN(n2102)
         );
  NOR2_X1 U2275 ( .A1(n35684), .A2(n10436), .ZN(n38074) );
  NOR2_X1 U2276 ( .A1(n18415), .A2(n22859), .ZN(n22863) );
  NAND2_X1 U2277 ( .A1(n11295), .A2(n22802), .ZN(n23123) );
  NOR2_X1 U2278 ( .A1(n37500), .A2(n284), .ZN(n37749) );
  NAND2_X1 U2280 ( .A1(n18147), .A2(n38789), .ZN(n36374) );
  OAI21_X1 U2282 ( .A1(n1146), .A2(n23053), .B(n23114), .ZN(n19229) );
  NOR2_X1 U2283 ( .A1(n6691), .A2(n37629), .ZN(n36167) );
  INV_X1 U2285 ( .I(n11476), .ZN(n10507) );
  NAND3_X1 U2286 ( .A1(n15330), .A2(n13650), .A3(n38986), .ZN(n39819) );
  NAND2_X1 U2298 ( .A1(n9854), .A2(n35684), .ZN(n39526) );
  AOI21_X1 U2300 ( .A1(n22558), .A2(n39518), .B(n6674), .ZN(n38559) );
  NOR2_X1 U2303 ( .A1(n37589), .A2(n23212), .ZN(n38492) );
  NOR2_X1 U2306 ( .A1(n7071), .A2(n1042), .ZN(n38541) );
  NAND2_X1 U2311 ( .A1(n22836), .A2(n23047), .ZN(n38800) );
  CLKBUF_X4 U2313 ( .I(n23125), .Z(n37883) );
  NAND2_X1 U2314 ( .A1(n3862), .A2(n23066), .ZN(n35310) );
  AOI21_X1 U2315 ( .A1(n20872), .A2(n23078), .B(n23077), .ZN(n15040) );
  INV_X1 U2318 ( .I(n22800), .ZN(n23210) );
  NAND2_X1 U2322 ( .A1(n5515), .A2(n20372), .ZN(n12163) );
  NAND2_X1 U2324 ( .A1(n14765), .A2(n19535), .ZN(n39046) );
  NAND2_X1 U2325 ( .A1(n17128), .A2(n9651), .ZN(n17319) );
  INV_X1 U2326 ( .I(n15330), .ZN(n11584) );
  OAI21_X1 U2331 ( .A1(n936), .A2(n10047), .B(n14089), .ZN(n34368) );
  NOR2_X1 U2339 ( .A1(n15163), .A2(n22944), .ZN(n17497) );
  NAND2_X1 U2345 ( .A1(n12729), .A2(n36422), .ZN(n14877) );
  INV_X1 U2351 ( .I(n38790), .ZN(n38789) );
  OAI21_X1 U2354 ( .A1(n10047), .A2(n39303), .B(n22816), .ZN(n12621) );
  NOR2_X1 U2361 ( .A1(n23188), .A2(n22979), .ZN(n39205) );
  NAND2_X1 U2362 ( .A1(n7160), .A2(n33972), .ZN(n22473) );
  INV_X1 U2365 ( .I(n4573), .ZN(n4931) );
  OR2_X1 U2368 ( .A1(n7518), .A2(n39446), .Z(n23047) );
  INV_X2 U2370 ( .I(n783), .ZN(n37922) );
  BUF_X2 U2373 ( .I(n37218), .Z(n4713) );
  CLKBUF_X2 U2379 ( .I(n15388), .Z(n38601) );
  OAI21_X1 U2383 ( .A1(n23169), .A2(n36554), .B(n23167), .ZN(n38790) );
  NAND2_X1 U2386 ( .A1(n39811), .A2(n19938), .ZN(n23099) );
  INV_X1 U2389 ( .I(n780), .ZN(n8730) );
  NAND2_X1 U2390 ( .A1(n13995), .A2(n17127), .ZN(n17124) );
  BUF_X2 U2392 ( .I(n14494), .Z(n6646) );
  INV_X1 U2397 ( .I(n11307), .ZN(n20783) );
  INV_X1 U2398 ( .I(n22678), .ZN(n37764) );
  BUF_X2 U2399 ( .I(n22740), .Z(n31863) );
  CLKBUF_X2 U2407 ( .I(n19931), .Z(n39682) );
  INV_X1 U2409 ( .I(n19814), .ZN(n39559) );
  OAI21_X1 U2411 ( .A1(n35014), .A2(n34090), .B(n22125), .ZN(n36849) );
  NAND2_X1 U2419 ( .A1(n37454), .A2(n37302), .ZN(n17536) );
  NOR2_X1 U2425 ( .A1(n16403), .A2(n8618), .ZN(n38747) );
  NAND2_X1 U2430 ( .A1(n7355), .A2(n1344), .ZN(n38479) );
  NOR2_X1 U2436 ( .A1(n20299), .A2(n1673), .ZN(n20298) );
  OAI21_X1 U2437 ( .A1(n38287), .A2(n2816), .B(n36006), .ZN(n6808) );
  NAND3_X1 U2438 ( .A1(n554), .A2(n22171), .A3(n18766), .ZN(n16435) );
  NAND3_X1 U2439 ( .A1(n5345), .A2(n18360), .A3(n5894), .ZN(n39111) );
  NAND2_X1 U2449 ( .A1(n22152), .A2(n17335), .ZN(n22153) );
  AND2_X1 U2450 ( .A1(n21968), .A2(n35780), .Z(n8574) );
  AND2_X1 U2451 ( .A1(n22349), .A2(n34813), .Z(n2909) );
  AOI21_X1 U2452 ( .A1(n21974), .A2(n21975), .B(n32640), .ZN(n21976) );
  NAND2_X1 U2454 ( .A1(n37794), .A2(n37793), .ZN(n22062) );
  OAI21_X1 U2461 ( .A1(n20758), .A2(n20759), .B(n37911), .ZN(n38869) );
  NOR2_X1 U2465 ( .A1(n33713), .A2(n22294), .ZN(n39237) );
  NOR2_X1 U2470 ( .A1(n7768), .A2(n1332), .ZN(n38911) );
  OAI22_X1 U2475 ( .A1(n37838), .A2(n22360), .B1(n11171), .B2(n31940), .ZN(
        n11379) );
  NAND2_X1 U2477 ( .A1(n33489), .A2(n22365), .ZN(n22006) );
  NAND2_X1 U2479 ( .A1(n11276), .A2(n22324), .ZN(n37454) );
  NAND2_X1 U2480 ( .A1(n5894), .A2(n5693), .ZN(n4874) );
  AOI21_X1 U2482 ( .A1(n4108), .A2(n6361), .B(n22327), .ZN(n34790) );
  OR2_X1 U2484 ( .A1(n915), .A2(n3863), .Z(n38917) );
  OAI21_X1 U2486 ( .A1(n6485), .A2(n21002), .B(n9987), .ZN(n15017) );
  NAND3_X1 U2492 ( .A1(n39010), .A2(n1337), .A3(n6297), .ZN(n22020) );
  NOR2_X1 U2494 ( .A1(n1049), .A2(n3907), .ZN(n22045) );
  OR2_X1 U2496 ( .A1(n22277), .A2(n8493), .Z(n37199) );
  BUF_X2 U2497 ( .I(n15697), .Z(n38830) );
  NAND2_X1 U2498 ( .A1(n14423), .A2(n32107), .ZN(n22390) );
  INV_X1 U2503 ( .I(n9938), .ZN(n37838) );
  NOR2_X1 U2507 ( .A1(n19873), .A2(n22349), .ZN(n38007) );
  NAND3_X1 U2513 ( .A1(n30893), .A2(n14020), .A3(n38448), .ZN(n37709) );
  BUF_X2 U2514 ( .I(n22240), .Z(n16888) );
  NAND2_X1 U2520 ( .A1(n22073), .A2(n38687), .ZN(n39377) );
  INV_X1 U2526 ( .I(n584), .ZN(n37794) );
  NOR2_X1 U2527 ( .A1(n22324), .A2(n22322), .ZN(n7636) );
  INV_X2 U2529 ( .I(n33086), .ZN(n22261) );
  NOR2_X1 U2532 ( .A1(n22282), .A2(n22281), .ZN(n38700) );
  BUF_X2 U2534 ( .I(n11568), .Z(n2910) );
  BUF_X2 U2538 ( .I(n7497), .Z(n584) );
  BUF_X2 U2540 ( .I(n20397), .Z(n33886) );
  NAND2_X1 U2541 ( .A1(n32313), .A2(n22263), .ZN(n39357) );
  INV_X2 U2550 ( .I(n35780), .ZN(n2186) );
  BUF_X2 U2553 ( .I(n18929), .Z(n6127) );
  OR2_X1 U2554 ( .A1(n21345), .A2(n21433), .Z(n37180) );
  BUF_X4 U2556 ( .I(n22400), .Z(n37089) );
  AOI21_X1 U2558 ( .A1(n39620), .A2(n21713), .B(n39619), .ZN(n39618) );
  NAND2_X1 U2561 ( .A1(n38546), .A2(n39192), .ZN(n38545) );
  NOR2_X1 U2567 ( .A1(n19650), .A2(n21876), .ZN(n21455) );
  INV_X1 U2569 ( .I(n38546), .ZN(n39620) );
  NAND2_X1 U2571 ( .A1(n1372), .A2(n21702), .ZN(n38340) );
  OR2_X1 U2573 ( .A1(n18968), .A2(n917), .Z(n37142) );
  AOI21_X1 U2577 ( .A1(n21784), .A2(n21405), .B(n21783), .ZN(n38938) );
  NOR3_X1 U2580 ( .A1(n21869), .A2(n21870), .A3(n15359), .ZN(n684) );
  NOR2_X1 U2584 ( .A1(n21808), .A2(n39639), .ZN(n21690) );
  NOR2_X1 U2585 ( .A1(n21914), .A2(n1352), .ZN(n5505) );
  OR2_X1 U2589 ( .A1(n37939), .A2(n39411), .Z(n21789) );
  CLKBUF_X2 U2591 ( .I(n33154), .Z(n39426) );
  BUF_X2 U2598 ( .I(n21848), .Z(n19517) );
  OR2_X1 U2600 ( .A1(n21669), .A2(n21848), .Z(n21850) );
  NAND2_X1 U2603 ( .A1(n21902), .A2(n35921), .ZN(n21422) );
  NOR2_X1 U2604 ( .A1(n21577), .A2(n21594), .ZN(n18784) );
  AND2_X1 U2617 ( .A1(n20476), .A2(n14769), .Z(n14577) );
  NAND2_X1 U2618 ( .A1(n4094), .A2(n19262), .ZN(n39368) );
  NAND2_X1 U2628 ( .A1(n19084), .A2(n21944), .ZN(n12752) );
  NAND3_X1 U2630 ( .A1(n20277), .A2(n21928), .A3(n12044), .ZN(n21728) );
  INV_X2 U2631 ( .I(n1157), .ZN(n38546) );
  CLKBUF_X2 U2633 ( .I(n18467), .Z(n5132) );
  AOI21_X2 U2638 ( .A1(n35302), .A2(n31739), .B(n23610), .ZN(n31816) );
  NAND3_X2 U2650 ( .A1(n30680), .A2(n19147), .A3(n19962), .ZN(n32197) );
  NAND2_X2 U2651 ( .A1(n30881), .A2(n388), .ZN(n8362) );
  NAND2_X2 U2654 ( .A1(n39305), .A2(n27449), .ZN(n31708) );
  NAND2_X2 U2656 ( .A1(n33091), .A2(n11344), .ZN(n11277) );
  INV_X2 U2658 ( .I(n25691), .ZN(n17271) );
  AOI22_X2 U2663 ( .A1(n18562), .A2(n5220), .B1(n5219), .B2(n1221), .ZN(n7680)
         );
  INV_X2 U2664 ( .I(n25351), .ZN(n25614) );
  INV_X4 U2667 ( .I(n29241), .ZN(n1062) );
  AND2_X1 U2668 ( .A1(n16933), .A2(n15515), .Z(n2246) );
  BUF_X4 U2670 ( .I(n32304), .Z(n10702) );
  AND2_X1 U2677 ( .A1(n15330), .A2(n20570), .Z(n37124) );
  NOR2_X2 U2679 ( .A1(n6443), .A2(n30153), .ZN(n14520) );
  BUF_X4 U2680 ( .I(n30249), .Z(n19663) );
  BUF_X4 U2682 ( .I(n20987), .Z(n39320) );
  BUF_X2 U2690 ( .I(n29166), .Z(n39798) );
  NOR2_X2 U2692 ( .A1(n24526), .A2(n37106), .ZN(n15169) );
  NAND2_X2 U2693 ( .A1(n9265), .A2(n38719), .ZN(n38718) );
  NAND2_X1 U2694 ( .A1(n31652), .A2(n18231), .ZN(n39234) );
  BUF_X2 U2695 ( .I(n8116), .Z(n124) );
  BUF_X4 U2697 ( .I(n16080), .Z(n36678) );
  BUF_X2 U2699 ( .I(n29174), .Z(n30160) );
  NOR2_X2 U2700 ( .A1(n28171), .A2(n28257), .ZN(n27885) );
  INV_X4 U2702 ( .I(n25801), .ZN(n1098) );
  OAI21_X2 U2710 ( .A1(n854), .A2(n26697), .B(n10736), .ZN(n26698) );
  NAND2_X2 U2714 ( .A1(n30587), .A2(n37432), .ZN(n5459) );
  NOR2_X2 U2715 ( .A1(n9310), .A2(n32870), .ZN(n27368) );
  BUF_X2 U2716 ( .I(n30454), .Z(n37319) );
  NAND3_X2 U2717 ( .A1(n17176), .A2(n37298), .A3(n9957), .ZN(n38697) );
  INV_X2 U2718 ( .I(n15368), .ZN(n15421) );
  NAND2_X1 U2719 ( .A1(n36485), .A2(n12425), .ZN(n12424) );
  BUF_X2 U2725 ( .I(n11297), .Z(n38491) );
  BUF_X2 U2728 ( .I(n6327), .Z(n37629) );
  AOI21_X2 U2731 ( .A1(n29182), .A2(n3986), .B(n32894), .ZN(n4072) );
  BUF_X4 U2732 ( .I(n32854), .Z(n34307) );
  INV_X2 U2733 ( .I(n18785), .ZN(n3965) );
  NAND2_X2 U2738 ( .A1(n4525), .A2(n23610), .ZN(n4527) );
  AOI21_X2 U2739 ( .A1(n39159), .A2(n27288), .B(n27069), .ZN(n6010) );
  INV_X4 U2740 ( .I(n22324), .ZN(n1683) );
  NOR2_X2 U2742 ( .A1(n14705), .A2(n16449), .ZN(n12772) );
  NAND2_X2 U2743 ( .A1(n39065), .A2(n31433), .ZN(n17661) );
  AOI22_X2 U2744 ( .A1(n21359), .A2(n1158), .B1(n21666), .B2(n19620), .ZN(
        n21362) );
  NAND2_X2 U2745 ( .A1(n23056), .A2(n23160), .ZN(n8758) );
  INV_X4 U2746 ( .I(n11150), .ZN(n952) );
  INV_X2 U2747 ( .I(n33347), .ZN(n28049) );
  OAI22_X2 U2748 ( .A1(n29335), .A2(n29341), .B1(n18601), .B2(n16889), .ZN(
        n29340) );
  NAND2_X2 U2749 ( .A1(n37859), .A2(n37858), .ZN(n37857) );
  INV_X2 U2750 ( .I(n33956), .ZN(n27996) );
  AOI21_X2 U2755 ( .A1(n9082), .A2(n18749), .B(n27318), .ZN(n3849) );
  BUF_X4 U2756 ( .I(n24034), .Z(n1614) );
  BUF_X2 U2759 ( .I(n39443), .Z(n37614) );
  INV_X2 U2765 ( .I(n197), .ZN(n691) );
  INV_X4 U2768 ( .I(n23889), .ZN(n17850) );
  INV_X2 U2769 ( .I(n4493), .ZN(n39176) );
  BUF_X4 U2775 ( .I(n26031), .Z(n37300) );
  INV_X2 U2776 ( .I(n13587), .ZN(n22944) );
  NOR2_X2 U2778 ( .A1(n13471), .A2(n35919), .ZN(n16101) );
  OAI22_X2 U2780 ( .A1(n26103), .A2(n18827), .B1(n1021), .B2(n17624), .ZN(
        n5327) );
  BUF_X4 U2782 ( .I(n7106), .Z(n269) );
  INV_X2 U2784 ( .I(n19318), .ZN(n29664) );
  INV_X4 U2786 ( .I(n12478), .ZN(n1531) );
  NOR2_X2 U2787 ( .A1(n24788), .A2(n19255), .ZN(n24609) );
  INV_X2 U2791 ( .I(n31433), .ZN(n34359) );
  INV_X2 U2792 ( .I(n18433), .ZN(n38604) );
  OR2_X2 U2796 ( .A1(n4899), .A2(n34987), .Z(n22886) );
  INV_X2 U2797 ( .I(n27564), .ZN(n990) );
  NAND2_X2 U2798 ( .A1(n4457), .A2(n36573), .ZN(n19125) );
  NAND2_X2 U2800 ( .A1(n12793), .A2(n4179), .ZN(n22154) );
  INV_X2 U2801 ( .I(n35705), .ZN(n38367) );
  NOR2_X2 U2806 ( .A1(n36371), .A2(n21982), .ZN(n21618) );
  AOI22_X2 U2807 ( .A1(n22176), .A2(n32609), .B1(n20234), .B2(n21616), .ZN(
        n2586) );
  INV_X2 U2809 ( .I(n17425), .ZN(n19151) );
  OAI21_X2 U2813 ( .A1(n1515), .A2(n37150), .B(n17008), .ZN(n39773) );
  NOR2_X2 U2820 ( .A1(n24753), .A2(n6756), .ZN(n24600) );
  INV_X1 U2824 ( .I(n37023), .ZN(n3734) );
  NAND2_X2 U2825 ( .A1(n13981), .A2(n29367), .ZN(n15958) );
  NAND2_X2 U2826 ( .A1(n11734), .A2(n5126), .ZN(n2139) );
  AOI21_X2 U2827 ( .A1(n23544), .A2(n17017), .B(n32351), .ZN(n23545) );
  NAND3_X2 U2829 ( .A1(n35193), .A2(n4497), .A3(n4493), .ZN(n4494) );
  INV_X2 U2830 ( .I(n2150), .ZN(n39386) );
  INV_X2 U2834 ( .I(n21687), .ZN(n38439) );
  NAND2_X2 U2835 ( .A1(n23468), .A2(n3256), .ZN(n7535) );
  BUF_X4 U2836 ( .I(n16631), .Z(n1448) );
  NAND2_X2 U2838 ( .A1(n5953), .A2(n1033), .ZN(n17592) );
  NAND2_X2 U2839 ( .A1(n26178), .A2(n26655), .ZN(n32482) );
  INV_X2 U2842 ( .I(n22475), .ZN(n22570) );
  NAND2_X1 U2844 ( .A1(n18070), .A2(n15259), .ZN(n15483) );
  NAND2_X1 U2845 ( .A1(n29236), .A2(n29231), .ZN(n15259) );
  OR2_X1 U2846 ( .A1(n28715), .A2(n19844), .Z(n28712) );
  BUF_X2 U2851 ( .I(n19844), .Z(n33460) );
  NOR2_X1 U2852 ( .A1(n33384), .A2(n25622), .ZN(n33597) );
  CLKBUF_X4 U2853 ( .I(n11657), .Z(n33384) );
  NOR2_X1 U2855 ( .A1(n759), .A2(n28205), .ZN(n7851) );
  NOR2_X1 U2862 ( .A1(n1439), .A2(n28205), .ZN(n39702) );
  INV_X1 U2864 ( .I(n30041), .ZN(n1405) );
  NAND2_X1 U2866 ( .A1(n16328), .A2(n30041), .ZN(n4220) );
  CLKBUF_X4 U2867 ( .I(n29149), .Z(n30041) );
  NAND2_X1 U2871 ( .A1(n39686), .A2(n39420), .ZN(n39567) );
  NAND2_X1 U2873 ( .A1(n4387), .A2(n3820), .ZN(n39420) );
  INV_X1 U2875 ( .I(n24040), .ZN(n30321) );
  NAND2_X1 U2876 ( .A1(n36824), .A2(n29171), .ZN(n36170) );
  NAND2_X1 U2878 ( .A1(n23392), .A2(n15642), .ZN(n23242) );
  INV_X1 U2880 ( .I(n23392), .ZN(n37528) );
  INV_X1 U2883 ( .I(n21813), .ZN(n35026) );
  OAI22_X1 U2884 ( .A1(n21813), .A2(n21682), .B1(n1350), .B2(n21684), .ZN(
        n21375) );
  NOR2_X1 U2888 ( .A1(n30196), .A2(n19693), .ZN(n38255) );
  NOR3_X1 U2889 ( .A1(n18261), .A2(n15248), .A3(n28109), .ZN(n38374) );
  CLKBUF_X2 U2891 ( .I(n22968), .Z(n45) );
  AOI22_X1 U2894 ( .A1(n35250), .A2(n34055), .B1(n12782), .B2(n14211), .ZN(
        n30960) );
  NOR2_X1 U2901 ( .A1(n9385), .A2(n35250), .ZN(n21049) );
  NAND2_X1 U2904 ( .A1(n5077), .A2(n22008), .ZN(n22214) );
  NOR2_X1 U2908 ( .A1(n25616), .A2(n25574), .ZN(n25420) );
  NAND2_X1 U2909 ( .A1(n25574), .A2(n38625), .ZN(n35419) );
  INV_X1 U2911 ( .I(n27470), .ZN(n27761) );
  INV_X2 U2912 ( .I(n14858), .ZN(n29338) );
  INV_X1 U2915 ( .I(n29501), .ZN(n37374) );
  OAI21_X1 U2916 ( .A1(n18374), .A2(n18743), .B(n10677), .ZN(n12108) );
  NAND2_X1 U2917 ( .A1(n18374), .A2(n35051), .ZN(n20150) );
  INV_X1 U2920 ( .I(n871), .ZN(n36223) );
  AOI22_X1 U2924 ( .A1(n18388), .A2(n33538), .B1(n18475), .B2(n7049), .ZN(
        n36091) );
  AOI22_X1 U2925 ( .A1(n1382), .A2(n30096), .B1(n14126), .B2(n30097), .ZN(
        n30099) );
  CLKBUF_X2 U2927 ( .I(n9267), .Z(n37890) );
  AOI22_X1 U2933 ( .A1(n3470), .A2(n9295), .B1(n3469), .B2(n16042), .ZN(n3468)
         );
  NAND2_X1 U2939 ( .A1(n8372), .A2(n19352), .ZN(n35424) );
  CLKBUF_X2 U2950 ( .I(n27095), .Z(n32046) );
  NAND2_X1 U2952 ( .A1(n14362), .A2(n3252), .ZN(n37809) );
  NOR2_X1 U2954 ( .A1(n6892), .A2(n12527), .ZN(n10908) );
  NAND2_X1 U2955 ( .A1(n11330), .A2(n6892), .ZN(n28726) );
  INV_X1 U2956 ( .I(n13223), .ZN(n27065) );
  NAND2_X1 U2960 ( .A1(n13223), .A2(n34562), .ZN(n12020) );
  BUF_X2 U2961 ( .I(n889), .Z(n13851) );
  NAND3_X1 U2965 ( .A1(n28189), .A2(n889), .A3(n16325), .ZN(n13322) );
  OAI21_X1 U2966 ( .A1(n39202), .A2(n32343), .B(n11513), .ZN(n31130) );
  NOR2_X1 U2970 ( .A1(n26748), .A2(n26800), .ZN(n2802) );
  INV_X1 U2983 ( .I(n31538), .ZN(n31539) );
  AOI21_X1 U2987 ( .A1(n28192), .A2(n9897), .B(n9553), .ZN(n15691) );
  NOR2_X1 U2988 ( .A1(n9897), .A2(n17598), .ZN(n33598) );
  INV_X2 U2989 ( .I(n20056), .ZN(n17598) );
  NAND2_X1 U2990 ( .A1(n27387), .A2(n2761), .ZN(n27289) );
  NAND2_X1 U2991 ( .A1(n11111), .A2(n4255), .ZN(n35787) );
  NAND2_X1 U2992 ( .A1(n30092), .A2(n30086), .ZN(n29175) );
  INV_X1 U2997 ( .I(n30096), .ZN(n30092) );
  NAND2_X1 U3000 ( .A1(n18562), .A2(n19203), .ZN(n13223) );
  INV_X2 U3004 ( .I(n27383), .ZN(n18562) );
  AND2_X1 U3008 ( .A1(n2522), .A2(n1891), .Z(n37191) );
  OAI21_X1 U3012 ( .A1(n35903), .A2(n9694), .B(n25978), .ZN(n31496) );
  NOR2_X1 U3013 ( .A1(n1221), .A2(n27385), .ZN(n13222) );
  CLKBUF_X1 U3014 ( .I(n15854), .Z(n32571) );
  NAND2_X1 U3015 ( .A1(n28657), .A2(n1197), .ZN(n14605) );
  NOR2_X1 U3018 ( .A1(n1197), .A2(n28560), .ZN(n38681) );
  NAND2_X1 U3019 ( .A1(n37592), .A2(n33383), .ZN(n37591) );
  INV_X1 U3021 ( .I(n29067), .ZN(n38087) );
  OR2_X1 U3022 ( .A1(n13587), .A2(n20555), .Z(n22974) );
  NAND2_X1 U3024 ( .A1(n7096), .A2(n27131), .ZN(n26889) );
  NAND2_X1 U3031 ( .A1(n12689), .A2(n2150), .ZN(n2152) );
  NAND2_X1 U3032 ( .A1(n29212), .A2(n13762), .ZN(n32267) );
  INV_X1 U3034 ( .I(n2139), .ZN(n4868) );
  AOI21_X1 U3036 ( .A1(n2139), .A2(n34745), .B(n1103), .ZN(n36387) );
  AOI22_X1 U3038 ( .A1(n2760), .A2(n2761), .B1(n34769), .B2(n20871), .ZN(
        n38873) );
  NOR2_X1 U3040 ( .A1(n30484), .A2(n1211), .ZN(n6733) );
  NAND2_X1 U3041 ( .A1(n1211), .A2(n30484), .ZN(n28032) );
  AOI21_X1 U3042 ( .A1(n8206), .A2(n1211), .B(n31808), .ZN(n30962) );
  INV_X1 U3043 ( .I(n14980), .ZN(n19765) );
  CLKBUF_X2 U3045 ( .I(n14980), .Z(n9872) );
  NAND3_X1 U3047 ( .A1(n34733), .A2(n35617), .A3(n2760), .ZN(n35616) );
  OAI22_X1 U3048 ( .A1(n9541), .A2(n18519), .B1(n18520), .B2(n19980), .ZN(
        n9540) );
  NAND2_X1 U3049 ( .A1(n19367), .A2(n18519), .ZN(n18520) );
  NAND2_X1 U3051 ( .A1(n38716), .A2(n18519), .ZN(n4792) );
  NAND3_X1 U3052 ( .A1(n3662), .A2(n36854), .A3(n32324), .ZN(n32752) );
  NOR2_X1 U3055 ( .A1(n7690), .A2(n3662), .ZN(n6058) );
  NAND2_X1 U3056 ( .A1(n38767), .A2(n4232), .ZN(n4005) );
  NAND2_X1 U3060 ( .A1(n34819), .A2(n28369), .ZN(n38767) );
  INV_X2 U3062 ( .I(n2269), .ZN(n29131) );
  AOI21_X1 U3066 ( .A1(n37858), .A2(n37375), .B(n37374), .ZN(n30353) );
  INV_X2 U3067 ( .I(n17017), .ZN(n1137) );
  NAND2_X1 U3069 ( .A1(n17017), .A2(n23566), .ZN(n23543) );
  NAND2_X1 U3070 ( .A1(n6040), .A2(n39147), .ZN(n6039) );
  NOR2_X1 U3072 ( .A1(n12218), .A2(n14426), .ZN(n5427) );
  CLKBUF_X1 U3073 ( .I(n30038), .Z(n35103) );
  NAND3_X1 U3075 ( .A1(n13006), .A2(n14997), .A3(n39603), .ZN(n38371) );
  OAI21_X1 U3076 ( .A1(n4882), .A2(n15615), .B(n30177), .ZN(n39603) );
  BUF_X1 U3077 ( .I(n35465), .Z(n37095) );
  AOI21_X1 U3081 ( .A1(n30255), .A2(n31529), .B(n39234), .ZN(n30256) );
  CLKBUF_X2 U3082 ( .I(n30262), .Z(n31529) );
  AOI22_X1 U3086 ( .A1(n19909), .A2(n29987), .B1(n29989), .B2(n31629), .ZN(
        n16589) );
  AOI22_X1 U3091 ( .A1(n907), .A2(n20018), .B1(n10451), .B2(n8918), .ZN(n35541) );
  OAI22_X1 U3095 ( .A1(n29176), .A2(n29175), .B1(n30099), .B2(n30087), .ZN(
        n37935) );
  NAND3_X1 U3096 ( .A1(n34621), .A2(n18431), .A3(n18070), .ZN(n20559) );
  NAND2_X1 U3097 ( .A1(n29351), .A2(n29385), .ZN(n29080) );
  INV_X1 U3098 ( .I(n29384), .ZN(n29351) );
  NAND2_X1 U3101 ( .A1(n16663), .A2(n13605), .ZN(n26643) );
  OAI21_X1 U3103 ( .A1(n26933), .A2(n4411), .B(n16663), .ZN(n18946) );
  BUF_X2 U3104 ( .I(n15855), .Z(n10587) );
  INV_X1 U3106 ( .I(n15855), .ZN(n28699) );
  CLKBUF_X2 U3110 ( .I(n15855), .Z(n38529) );
  NAND2_X1 U3113 ( .A1(n33784), .A2(n30241), .ZN(n7749) );
  NOR2_X1 U3114 ( .A1(n17501), .A2(n26098), .ZN(n25872) );
  INV_X1 U3117 ( .I(n26098), .ZN(n25447) );
  OR2_X1 U3120 ( .A1(n26098), .A2(n3874), .Z(n25445) );
  NAND3_X1 U3121 ( .A1(n33815), .A2(n26098), .A3(n31367), .ZN(n32053) );
  NAND2_X1 U3122 ( .A1(n26098), .A2(n10223), .ZN(n39250) );
  OAI21_X1 U3124 ( .A1(n26903), .A2(n26901), .B(n26652), .ZN(n17228) );
  INV_X1 U3125 ( .I(n26901), .ZN(n39287) );
  NAND3_X1 U3126 ( .A1(n34005), .A2(n26754), .A3(n26901), .ZN(n26755) );
  CLKBUF_X4 U3127 ( .I(n29347), .Z(n17225) );
  NOR2_X1 U3134 ( .A1(n2059), .A2(n36788), .ZN(n28538) );
  NOR2_X1 U3136 ( .A1(n2059), .A2(n1434), .ZN(n27457) );
  BUF_X1 U3145 ( .I(n8787), .Z(n2059) );
  NOR3_X1 U3146 ( .A1(n24266), .A2(n19745), .A3(n24267), .ZN(n24029) );
  OR2_X1 U3147 ( .A1(n39277), .A2(n14709), .Z(n9020) );
  NAND2_X1 U3148 ( .A1(n18398), .A2(n37809), .ZN(n12046) );
  NOR2_X1 U3149 ( .A1(n10346), .A2(n29586), .ZN(n29629) );
  NAND2_X1 U3154 ( .A1(n39018), .A2(n29810), .ZN(n29799) );
  NAND2_X1 U3156 ( .A1(n25924), .A2(n26027), .ZN(n15377) );
  AOI22_X1 U3157 ( .A1(n28657), .A2(n38681), .B1(n28442), .B2(n28559), .ZN(
        n3050) );
  OAI22_X1 U3158 ( .A1(n29904), .A2(n14600), .B1(n18222), .B2(n1407), .ZN(
        n31356) );
  INV_X1 U3159 ( .I(n12940), .ZN(n37914) );
  NAND2_X1 U3166 ( .A1(n12940), .A2(n18667), .ZN(n11597) );
  NOR2_X1 U3169 ( .A1(n12940), .A2(n19783), .ZN(n17794) );
  BUF_X2 U3170 ( .I(n33368), .Z(n38580) );
  NOR2_X1 U3172 ( .A1(n29630), .A2(n21269), .ZN(n10081) );
  NOR2_X1 U3174 ( .A1(n33784), .A2(n30796), .ZN(n31238) );
  AND2_X1 U3175 ( .A1(n30178), .A2(n12198), .Z(n4882) );
  NAND2_X1 U3178 ( .A1(n38407), .A2(n13757), .ZN(n20635) );
  NAND3_X1 U3180 ( .A1(n13757), .A2(n38407), .A3(n32345), .ZN(n26626) );
  AOI22_X1 U3181 ( .A1(n8761), .A2(n28882), .B1(n20085), .B2(n8762), .ZN(
        n38698) );
  NOR2_X1 U3182 ( .A1(n33482), .A2(n14417), .ZN(n2294) );
  BUF_X1 U3187 ( .I(n29591), .Z(n33482) );
  NAND2_X1 U3190 ( .A1(n105), .A2(n29996), .ZN(n21290) );
  NAND3_X1 U3192 ( .A1(n33130), .A2(n841), .A3(n21042), .ZN(n33304) );
  OAI21_X1 U3195 ( .A1(n841), .A2(n12131), .B(n25359), .ZN(n10935) );
  NOR2_X1 U3198 ( .A1(n5963), .A2(n3573), .ZN(n6012) );
  INV_X2 U3205 ( .I(n15189), .ZN(n38141) );
  NAND2_X1 U3207 ( .A1(n29732), .A2(n29755), .ZN(n29750) );
  NAND2_X1 U3208 ( .A1(n4368), .A2(n20342), .ZN(n30180) );
  NAND2_X1 U3210 ( .A1(n39274), .A2(n29459), .ZN(n37859) );
  AND2_X1 U3212 ( .A1(n25867), .A2(n5859), .Z(n25747) );
  NAND2_X1 U3217 ( .A1(n25367), .A2(n25513), .ZN(n15788) );
  NOR3_X1 U3222 ( .A1(n25367), .A2(n25540), .A3(n30317), .ZN(n16428) );
  INV_X2 U3223 ( .I(n25539), .ZN(n25367) );
  AOI21_X1 U3227 ( .A1(n29642), .A2(n30680), .B(n37303), .ZN(n29488) );
  NAND2_X1 U3230 ( .A1(n7373), .A2(n37304), .ZN(n37303) );
  INV_X1 U3232 ( .I(n28714), .ZN(n17077) );
  NAND2_X1 U3234 ( .A1(n1425), .A2(n31015), .ZN(n28714) );
  NAND3_X1 U3238 ( .A1(n35731), .A2(n15307), .A3(n15310), .ZN(n17366) );
  NAND2_X1 U3243 ( .A1(n14158), .A2(n19424), .ZN(n29904) );
  NOR2_X1 U3246 ( .A1(n8677), .A2(n14158), .ZN(n10610) );
  INV_X1 U3247 ( .I(n9106), .ZN(n34740) );
  INV_X1 U3249 ( .I(n26441), .ZN(n38530) );
  NAND3_X1 U3251 ( .A1(n28051), .A2(n11891), .A3(n28123), .ZN(n17236) );
  OAI22_X1 U3252 ( .A1(n29787), .A2(n15867), .B1(n29788), .B2(n29789), .ZN(
        n37781) );
  NAND2_X1 U3257 ( .A1(n30665), .A2(n34075), .ZN(n12565) );
  CLKBUF_X2 U3262 ( .I(n30043), .Z(n35809) );
  NOR2_X1 U3265 ( .A1(n30042), .A2(n16328), .ZN(n29898) );
  INV_X1 U3267 ( .I(n36827), .ZN(n980) );
  NOR2_X1 U3270 ( .A1(n8476), .A2(n36827), .ZN(n28604) );
  NAND2_X1 U3275 ( .A1(n8476), .A2(n36827), .ZN(n10542) );
  NAND2_X1 U3276 ( .A1(n27452), .A2(n15276), .ZN(n40) );
  INV_X1 U3277 ( .I(n12350), .ZN(n30139) );
  NAND3_X1 U3279 ( .A1(n34180), .A2(n37565), .A3(n35858), .ZN(n8996) );
  AOI21_X1 U3289 ( .A1(n27822), .A2(n28257), .B(n9880), .ZN(n12529) );
  NAND2_X1 U3290 ( .A1(n33928), .A2(n14940), .ZN(n37545) );
  CLKBUF_X2 U3292 ( .I(n30233), .Z(n14940) );
  OAI21_X1 U3293 ( .A1(n36481), .A2(n30046), .B(n29185), .ZN(n36328) );
  BUF_X2 U3296 ( .I(n14559), .Z(n36481) );
  OAI21_X1 U3297 ( .A1(n30162), .A2(n29185), .B(n36481), .ZN(n28822) );
  NAND2_X1 U3299 ( .A1(n30034), .A2(n30033), .ZN(n30017) );
  NAND2_X1 U3301 ( .A1(n30033), .A2(n30022), .ZN(n30032) );
  NAND2_X1 U3307 ( .A1(n30033), .A2(n8039), .ZN(n30026) );
  INV_X1 U3309 ( .I(n38196), .ZN(n37813) );
  CLKBUF_X2 U3310 ( .I(n19050), .Z(n38196) );
  BUF_X2 U3311 ( .I(n19226), .Z(n26764) );
  NOR2_X1 U3313 ( .A1(n19349), .A2(n32002), .ZN(n30334) );
  OAI21_X1 U3315 ( .A1(n19497), .A2(n5067), .B(n20672), .ZN(n29668) );
  NAND2_X1 U3317 ( .A1(n36471), .A2(n24802), .ZN(n13748) );
  INV_X1 U3319 ( .I(n36471), .ZN(n24804) );
  NAND2_X1 U3321 ( .A1(n26097), .A2(n17700), .ZN(n15618) );
  NOR2_X1 U3322 ( .A1(n39305), .A2(n36969), .ZN(n36762) );
  NOR2_X1 U3324 ( .A1(n27265), .A2(n39305), .ZN(n31934) );
  OAI21_X1 U3325 ( .A1(n29597), .A2(n29595), .B(n29596), .ZN(n39006) );
  NAND2_X1 U3327 ( .A1(n2292), .A2(n26959), .ZN(n2100) );
  INV_X2 U3328 ( .I(n26959), .ZN(n8651) );
  CLKBUF_X4 U3329 ( .I(n26959), .Z(n30665) );
  AOI21_X1 U3333 ( .A1(n29960), .A2(n29955), .B(n29862), .ZN(n17148) );
  NAND3_X1 U3337 ( .A1(n29960), .A2(n19878), .A3(n29862), .ZN(n29845) );
  INV_X1 U3338 ( .I(n5344), .ZN(n37638) );
  NOR2_X1 U3342 ( .A1(n865), .A2(n17535), .ZN(n39202) );
  OAI22_X1 U3344 ( .A1(n28714), .A2(n28715), .B1(n28712), .B2(n1193), .ZN(
        n37862) );
  AOI21_X1 U3347 ( .A1(n31015), .A2(n33460), .B(n1193), .ZN(n8216) );
  OAI22_X1 U3349 ( .A1(n29533), .A2(n35180), .B1(n37605), .B2(n29536), .ZN(
        n30645) );
  CLKBUF_X4 U3350 ( .I(n17730), .Z(n5921) );
  AND2_X1 U3352 ( .A1(n8293), .A2(n20361), .Z(n7962) );
  OAI21_X1 U3354 ( .A1(n38658), .A2(n34666), .B(n30421), .ZN(n24546) );
  INV_X1 U3355 ( .I(n34609), .ZN(n1100) );
  INV_X1 U3359 ( .I(n13365), .ZN(n7790) );
  NAND2_X1 U3362 ( .A1(n32791), .A2(n9848), .ZN(n17191) );
  INV_X1 U3366 ( .I(n9848), .ZN(n27907) );
  BUF_X2 U3367 ( .I(n9848), .Z(n39664) );
  NAND2_X1 U3368 ( .A1(n26687), .A2(n17097), .ZN(n11866) );
  NOR2_X1 U3370 ( .A1(n28723), .A2(n28722), .ZN(n15313) );
  NAND2_X1 U3374 ( .A1(n38145), .A2(n28722), .ZN(n28679) );
  CLKBUF_X2 U3378 ( .I(n29696), .Z(n29763) );
  NAND2_X1 U3380 ( .A1(n37349), .A2(n28637), .ZN(n38818) );
  NAND2_X1 U3385 ( .A1(n19115), .A2(n5009), .ZN(n37349) );
  AOI22_X1 U3388 ( .A1(n7048), .A2(n38535), .B1(n2175), .B2(n37463), .ZN(
        n38025) );
  INV_X1 U3389 ( .I(n28262), .ZN(n28257) );
  CLKBUF_X2 U3393 ( .I(n28262), .Z(n3990) );
  BUF_X1 U3394 ( .I(n33967), .Z(n31095) );
  CLKBUF_X4 U3395 ( .I(n15573), .Z(n15447) );
  NAND2_X1 U3400 ( .A1(n33972), .A2(n15033), .ZN(n39153) );
  NAND2_X1 U3403 ( .A1(n30056), .A2(n3818), .ZN(n35095) );
  AND2_X1 U3405 ( .A1(n29220), .A2(n18240), .Z(n14421) );
  AOI21_X1 U3408 ( .A1(n29870), .A2(n28), .B(n29692), .ZN(n29693) );
  INV_X2 U3409 ( .I(n29870), .ZN(n33094) );
  NOR2_X1 U3410 ( .A1(n10096), .A2(n29870), .ZN(n32359) );
  OR2_X1 U3416 ( .A1(n9214), .A2(n9235), .Z(n26652) );
  AOI22_X1 U3417 ( .A1(n38829), .A2(n33437), .B1(n30216), .B2(n38227), .ZN(
        n38267) );
  OR2_X1 U3418 ( .A1(n37013), .A2(n29005), .Z(n5736) );
  INV_X1 U3422 ( .I(n25252), .ZN(n38958) );
  CLKBUF_X4 U3426 ( .I(n30242), .Z(n32415) );
  NAND2_X1 U3427 ( .A1(n1068), .A2(n28676), .ZN(n28576) );
  AOI21_X1 U3428 ( .A1(n35199), .A2(n28591), .B(n28676), .ZN(n14701) );
  NOR2_X1 U3429 ( .A1(n39126), .A2(n28141), .ZN(n10756) );
  NOR2_X1 U3432 ( .A1(n33405), .A2(n28141), .ZN(n9655) );
  CLKBUF_X2 U3440 ( .I(n28141), .Z(n39298) );
  NAND3_X1 U3441 ( .A1(n30506), .A2(n35377), .A3(n36191), .ZN(n23290) );
  BUF_X2 U3442 ( .I(n6640), .Z(n200) );
  CLKBUF_X2 U3444 ( .I(n21792), .Z(n16945) );
  NOR2_X1 U3454 ( .A1(n2802), .A2(n2801), .ZN(n8990) );
  NAND2_X1 U3458 ( .A1(n29209), .A2(n11567), .ZN(n9806) );
  NAND2_X1 U3459 ( .A1(n37544), .A2(n14940), .ZN(n14892) );
  NAND2_X1 U3460 ( .A1(n1595), .A2(n19915), .ZN(n15143) );
  OAI22_X1 U3462 ( .A1(n26865), .A2(n39737), .B1(n39598), .B2(n36549), .ZN(
        n16124) );
  NOR2_X1 U3463 ( .A1(n39449), .A2(n36549), .ZN(n10974) );
  NAND2_X1 U3464 ( .A1(n17831), .A2(n18785), .ZN(n3966) );
  CLKBUF_X4 U3468 ( .I(n28692), .Z(n8349) );
  AOI21_X1 U3469 ( .A1(n29185), .A2(n482), .B(n1181), .ZN(n11803) );
  INV_X2 U3470 ( .I(n7907), .ZN(n30128) );
  CLKBUF_X2 U3471 ( .I(n7907), .Z(n32508) );
  AND2_X1 U3476 ( .A1(n39583), .A2(n27252), .Z(n10581) );
  OR2_X1 U3482 ( .A1(n27252), .A2(n39583), .Z(n4105) );
  AND2_X1 U3483 ( .A1(n5410), .A2(n8116), .Z(n3133) );
  CLKBUF_X4 U3484 ( .I(n29568), .Z(n29571) );
  NAND2_X1 U3485 ( .A1(n9200), .A2(n33521), .ZN(n30201) );
  NAND2_X1 U3487 ( .A1(n28722), .A2(n28680), .ZN(n2790) );
  NOR2_X1 U3488 ( .A1(n13594), .A2(n28680), .ZN(n28360) );
  CLKBUF_X4 U3489 ( .I(n15113), .Z(n5093) );
  AOI21_X1 U3494 ( .A1(n26847), .A2(n26614), .B(n26849), .ZN(n16941) );
  OAI21_X1 U3495 ( .A1(n26847), .A2(n167), .B(n26945), .ZN(n34396) );
  INV_X2 U3499 ( .I(n14453), .ZN(n26847) );
  INV_X2 U3500 ( .I(n15473), .ZN(n28724) );
  NAND2_X1 U3502 ( .A1(n37311), .A2(n15473), .ZN(n28501) );
  NAND2_X1 U3506 ( .A1(n4369), .A2(n28463), .ZN(n28095) );
  NAND2_X1 U3507 ( .A1(n19113), .A2(n28463), .ZN(n19115) );
  AOI21_X1 U3508 ( .A1(n30077), .A2(n3818), .B(n31120), .ZN(n6488) );
  NAND2_X1 U3511 ( .A1(n31120), .A2(n30077), .ZN(n39022) );
  INV_X2 U3512 ( .I(n28313), .ZN(n1193) );
  NOR2_X1 U3513 ( .A1(n28313), .A2(n19844), .ZN(n28510) );
  NAND2_X1 U3519 ( .A1(n22795), .A2(n35213), .ZN(n16967) );
  CLKBUF_X2 U3523 ( .I(n22795), .Z(n34457) );
  NAND2_X1 U3525 ( .A1(n34014), .A2(n22795), .ZN(n13688) );
  INV_X1 U3526 ( .I(n19384), .ZN(n37882) );
  NOR2_X1 U3527 ( .A1(n457), .A2(n39406), .ZN(n34277) );
  NAND2_X1 U3530 ( .A1(n39406), .A2(n9197), .ZN(n33541) );
  AOI21_X1 U3537 ( .A1(n9197), .A2(n39406), .B(n39405), .ZN(n37515) );
  NAND2_X1 U3538 ( .A1(n31095), .A2(n14400), .ZN(n29375) );
  NAND2_X1 U3541 ( .A1(n14400), .A2(n9333), .ZN(n38461) );
  INV_X2 U3547 ( .I(n4947), .ZN(n6065) );
  NOR2_X1 U3549 ( .A1(n4947), .A2(n1530), .ZN(n7467) );
  NAND2_X1 U3550 ( .A1(n2148), .A2(n4947), .ZN(n4755) );
  NAND2_X1 U3553 ( .A1(n3053), .A2(n3052), .ZN(n34291) );
  OAI21_X1 U3554 ( .A1(n4284), .A2(n1419), .B(n34695), .ZN(n3053) );
  CLKBUF_X2 U3558 ( .I(n5638), .Z(n5471) );
  INV_X1 U3559 ( .I(n28465), .ZN(n39365) );
  OAI21_X1 U3560 ( .A1(n28639), .A2(n33046), .B(n28465), .ZN(n31030) );
  NAND2_X1 U3562 ( .A1(n11389), .A2(n9955), .ZN(n5645) );
  INV_X1 U3563 ( .I(n18004), .ZN(n15591) );
  OR2_X1 U3564 ( .A1(n14000), .A2(n18903), .Z(n18904) );
  NAND2_X1 U3566 ( .A1(n20429), .A2(n13261), .ZN(n32987) );
  INV_X1 U3567 ( .I(n28638), .ZN(n19113) );
  NAND2_X1 U3578 ( .A1(n28638), .A2(n28464), .ZN(n28465) );
  NAND2_X1 U3579 ( .A1(n15573), .A2(n28638), .ZN(n5009) );
  NAND2_X1 U3580 ( .A1(n20453), .A2(n30186), .ZN(n34344) );
  OAI21_X1 U3583 ( .A1(n23469), .A2(n32930), .B(n36448), .ZN(n39670) );
  AOI22_X1 U3584 ( .A1(n30417), .A2(n36448), .B1(n8680), .B2(n37839), .ZN(
        n39333) );
  NOR2_X1 U3586 ( .A1(n23645), .A2(n36448), .ZN(n4634) );
  CLKBUF_X2 U3587 ( .I(n8026), .Z(n35590) );
  OAI21_X1 U3589 ( .A1(n29309), .A2(n31279), .B(n6262), .ZN(n39134) );
  AOI21_X1 U3592 ( .A1(n18031), .A2(n25614), .B(n2721), .ZN(n36434) );
  CLKBUF_X4 U3595 ( .I(n26249), .Z(n26970) );
  NAND2_X1 U3596 ( .A1(n26876), .A2(n26249), .ZN(n15124) );
  CLKBUF_X1 U3598 ( .I(n18186), .Z(n5062) );
  NAND2_X1 U3600 ( .A1(n23181), .A2(n22903), .ZN(n20957) );
  AOI22_X1 U3601 ( .A1(n15040), .A2(n15039), .B1(n18851), .B2(n23181), .ZN(
        n31319) );
  NAND2_X1 U3604 ( .A1(n28659), .A2(n31663), .ZN(n28437) );
  INV_X1 U3605 ( .I(n28437), .ZN(n28438) );
  NOR2_X1 U3607 ( .A1(n28437), .A2(n28554), .ZN(n35000) );
  AOI21_X1 U3608 ( .A1(n17031), .A2(n3538), .B(n28742), .ZN(n11474) );
  NAND2_X1 U3609 ( .A1(n11506), .A2(n29437), .ZN(n12321) );
  NOR2_X1 U3612 ( .A1(n1392), .A2(n29437), .ZN(n14414) );
  OR2_X1 U3616 ( .A1(n1812), .A2(n34475), .Z(n15229) );
  INV_X1 U3618 ( .I(n7506), .ZN(n1268) );
  NOR2_X1 U3622 ( .A1(n7506), .A2(n24903), .ZN(n24904) );
  NAND2_X1 U3628 ( .A1(n19050), .A2(n33963), .ZN(n4805) );
  NOR2_X1 U3629 ( .A1(n33288), .A2(n20889), .ZN(n20355) );
  NAND2_X1 U3631 ( .A1(n16398), .A2(n209), .ZN(n31643) );
  OAI21_X1 U3632 ( .A1(n36465), .A2(n13404), .B(n37898), .ZN(n32524) );
  NAND2_X1 U3633 ( .A1(n37898), .A2(n974), .ZN(n28340) );
  AOI21_X1 U3634 ( .A1(n19005), .A2(n33864), .B(n23380), .ZN(n6518) );
  INV_X1 U3636 ( .I(n11125), .ZN(n33278) );
  NOR2_X1 U3640 ( .A1(n34652), .A2(n7141), .ZN(n37274) );
  AOI21_X1 U3641 ( .A1(n28050), .A2(n28124), .B(n14404), .ZN(n27152) );
  INV_X2 U3649 ( .I(n14404), .ZN(n983) );
  AOI22_X1 U3651 ( .A1(n9660), .A2(n33697), .B1(n22902), .B2(n36369), .ZN(
        n12130) );
  AOI22_X1 U3654 ( .A1(n5982), .A2(n30883), .B1(n5981), .B2(n3345), .ZN(n31630) );
  NAND2_X1 U3655 ( .A1(n3345), .A2(n37997), .ZN(n26237) );
  NAND2_X1 U3656 ( .A1(n9694), .A2(n3345), .ZN(n35947) );
  NAND2_X1 U3657 ( .A1(n37997), .A2(n3345), .ZN(n37996) );
  INV_X2 U3658 ( .I(n34265), .ZN(n3345) );
  AOI21_X1 U3659 ( .A1(n17857), .A2(n2906), .B(n7044), .ZN(n2905) );
  NAND2_X1 U3662 ( .A1(n7044), .A2(n34011), .ZN(n2904) );
  NOR2_X1 U3668 ( .A1(n34011), .A2(n7044), .ZN(n24601) );
  NAND2_X1 U3669 ( .A1(n7044), .A2(n32882), .ZN(n3044) );
  OAI21_X1 U3670 ( .A1(n27377), .A2(n8137), .B(n6445), .ZN(n27381) );
  NAND2_X1 U3671 ( .A1(n39153), .A2(n34131), .ZN(n15452) );
  OAI21_X1 U3678 ( .A1(n27998), .A2(n18061), .B(n11461), .ZN(n8524) );
  NAND2_X1 U3681 ( .A1(n28200), .A2(n18061), .ZN(n37322) );
  NOR2_X1 U3682 ( .A1(n1022), .A2(n25695), .ZN(n31131) );
  NAND2_X1 U3684 ( .A1(n34424), .A2(n33579), .ZN(n34422) );
  NOR3_X1 U3685 ( .A1(n33579), .A2(n2192), .A3(n37107), .ZN(n37439) );
  CLKBUF_X2 U3686 ( .I(n11753), .Z(n37951) );
  OAI21_X1 U3687 ( .A1(n6902), .A2(n6901), .B(n4573), .ZN(n6900) );
  AOI21_X1 U3688 ( .A1(n4573), .A2(n640), .B(n33554), .ZN(n37750) );
  OAI21_X1 U3691 ( .A1(n4573), .A2(n640), .B(n1318), .ZN(n39297) );
  NAND2_X1 U3694 ( .A1(n25829), .A2(n2830), .ZN(n6097) );
  INV_X2 U3696 ( .I(n18017), .ZN(n25692) );
  NOR2_X1 U3697 ( .A1(n19914), .A2(n1006), .ZN(n11305) );
  OAI21_X1 U3698 ( .A1(n1493), .A2(n14458), .B(n19914), .ZN(n5746) );
  NAND2_X1 U3699 ( .A1(n13491), .A2(n281), .ZN(n27935) );
  NOR2_X1 U3702 ( .A1(n281), .A2(n12663), .ZN(n13059) );
  NAND3_X1 U3704 ( .A1(n32354), .A2(n8380), .A3(n8381), .ZN(n5622) );
  INV_X1 U3706 ( .I(n32354), .ZN(n37270) );
  NOR2_X1 U3707 ( .A1(n19782), .A2(n24465), .ZN(n24251) );
  OAI21_X1 U3708 ( .A1(n24465), .A2(n24467), .B(n18347), .ZN(n24158) );
  NOR2_X1 U3717 ( .A1(n18348), .A2(n24465), .ZN(n7361) );
  NAND2_X1 U3718 ( .A1(n35903), .A2(n4553), .ZN(n26034) );
  NOR2_X1 U3720 ( .A1(n26838), .A2(n1092), .ZN(n3093) );
  OAI22_X1 U3723 ( .A1(n24351), .A2(n9921), .B1(n3487), .B2(n18653), .ZN(
        n12643) );
  AOI21_X1 U3724 ( .A1(n5957), .A2(n18653), .B(n24770), .ZN(n13428) );
  NAND2_X1 U3726 ( .A1(n18653), .A2(n3487), .ZN(n39182) );
  NAND2_X1 U3727 ( .A1(n26219), .A2(n1494), .ZN(n20547) );
  NAND2_X1 U3728 ( .A1(n9268), .A2(n11162), .ZN(n8601) );
  AOI21_X1 U3729 ( .A1(n26953), .A2(n11162), .B(n30768), .ZN(n11463) );
  NAND2_X1 U3737 ( .A1(n27508), .A2(n998), .ZN(n11162) );
  AOI21_X1 U3741 ( .A1(n33935), .A2(n22129), .B(n8245), .ZN(n17778) );
  OAI21_X1 U3743 ( .A1(n12630), .A2(n33935), .B(n7496), .ZN(n7495) );
  AOI21_X1 U3745 ( .A1(n6366), .A2(n33935), .B(n1831), .ZN(n7496) );
  NAND2_X1 U3746 ( .A1(n1831), .A2(n33935), .ZN(n22909) );
  NOR2_X1 U3748 ( .A1(n16463), .A2(n33935), .ZN(n37517) );
  NOR3_X1 U3751 ( .A1(n28023), .A2(n6643), .A3(n16065), .ZN(n32150) );
  INV_X2 U3752 ( .I(n16065), .ZN(n989) );
  AOI22_X1 U3753 ( .A1(n15669), .A2(n26852), .B1(n15668), .B2(n167), .ZN(
        n15667) );
  NOR2_X1 U3754 ( .A1(n26852), .A2(n38797), .ZN(n39257) );
  BUF_X2 U3755 ( .I(n26852), .Z(n15670) );
  OAI21_X1 U3756 ( .A1(n11432), .A2(n27337), .B(n11431), .ZN(n26890) );
  NAND2_X1 U3757 ( .A1(n39417), .A2(n4886), .ZN(n27218) );
  INV_X1 U3759 ( .I(n39417), .ZN(n35745) );
  NAND2_X1 U3761 ( .A1(n27069), .A2(n39417), .ZN(n6013) );
  NAND2_X1 U3764 ( .A1(n38097), .A2(n2741), .ZN(n14203) );
  CLKBUF_X4 U3765 ( .I(n4378), .Z(n3818) );
  INV_X1 U3766 ( .I(n17184), .ZN(n17395) );
  CLKBUF_X2 U3767 ( .I(n17184), .Z(n38714) );
  NAND2_X1 U3769 ( .A1(n35523), .A2(n38327), .ZN(n38056) );
  AND2_X1 U3770 ( .A1(n5530), .A2(n29284), .Z(n6843) );
  NAND3_X1 U3774 ( .A1(n30258), .A2(n11700), .A3(n19663), .ZN(n31652) );
  INV_X1 U3775 ( .I(n26660), .ZN(n26697) );
  CLKBUF_X4 U3777 ( .I(n15423), .Z(n8757) );
  NAND2_X1 U3779 ( .A1(n6357), .A2(n30464), .ZN(n18653) );
  OAI21_X1 U3780 ( .A1(n13170), .A2(n35357), .B(n5465), .ZN(n8635) );
  NAND2_X1 U3782 ( .A1(n35357), .A2(n19759), .ZN(n31347) );
  AOI22_X1 U3783 ( .A1(n33577), .A2(n28812), .B1(n28764), .B2(n35357), .ZN(
        n32376) );
  OAI21_X1 U3786 ( .A1(n28808), .A2(n35357), .B(n31542), .ZN(n35083) );
  NAND3_X1 U3787 ( .A1(n30292), .A2(n35357), .A3(n28764), .ZN(n33675) );
  OAI21_X1 U3790 ( .A1(n30161), .A2(n30162), .B(n1400), .ZN(n11429) );
  NAND2_X1 U3793 ( .A1(n11125), .A2(n30161), .ZN(n39686) );
  OAI21_X1 U3796 ( .A1(n2522), .A2(n35919), .B(n38414), .ZN(n3996) );
  CLKBUF_X2 U3799 ( .I(n4771), .Z(n39448) );
  AND2_X1 U3800 ( .A1(n8412), .A2(n4771), .Z(n16144) );
  AND3_X1 U3801 ( .A1(n27440), .A2(n27438), .A3(n4771), .Z(n161) );
  INV_X1 U3804 ( .I(n4771), .ZN(n13992) );
  OR2_X1 U3811 ( .A1(n4771), .A2(n27438), .Z(n11638) );
  INV_X2 U3815 ( .I(n13650), .ZN(n34184) );
  AOI21_X1 U3817 ( .A1(n603), .A2(n32691), .B(n25912), .ZN(n32056) );
  AOI21_X1 U3819 ( .A1(n32691), .A2(n25912), .B(n32690), .ZN(n32689) );
  CLKBUF_X2 U3820 ( .I(n12572), .Z(n7892) );
  NOR2_X1 U3821 ( .A1(n9444), .A2(n28533), .ZN(n9443) );
  NOR2_X1 U3824 ( .A1(n8727), .A2(n29851), .ZN(n37390) );
  OAI21_X1 U3828 ( .A1(n2969), .A2(n32168), .B(n32559), .ZN(n2968) );
  NAND2_X1 U3830 ( .A1(n31716), .A2(n27049), .ZN(n12745) );
  INV_X1 U3837 ( .I(n27049), .ZN(n54) );
  OAI22_X1 U3841 ( .A1(n38611), .A2(n14739), .B1(n20788), .B2(n23610), .ZN(
        n4528) );
  INV_X1 U3842 ( .I(n856), .ZN(n17158) );
  BUF_X2 U3843 ( .I(n856), .Z(n11138) );
  NOR2_X1 U3845 ( .A1(n27405), .A2(n27155), .ZN(n32853) );
  OAI21_X1 U3846 ( .A1(n29310), .A2(n12880), .B(n10422), .ZN(n12879) );
  AND2_X1 U3847 ( .A1(n29384), .A2(n10422), .Z(n35966) );
  OR3_X1 U3849 ( .A1(n11084), .A2(n36426), .A3(n10422), .Z(n1822) );
  INV_X1 U3850 ( .I(n11383), .ZN(n37721) );
  NOR3_X1 U3852 ( .A1(n24473), .A2(n15461), .A3(n39309), .ZN(n33085) );
  CLKBUF_X1 U3862 ( .I(n24473), .Z(n37916) );
  BUF_X2 U3866 ( .I(n36894), .Z(n34829) );
  BUF_X2 U3869 ( .I(n9918), .Z(n39576) );
  NOR2_X1 U3873 ( .A1(n29940), .A2(n9918), .ZN(n29939) );
  NAND2_X1 U3874 ( .A1(n29940), .A2(n9918), .ZN(n9143) );
  NOR2_X1 U3877 ( .A1(n32854), .A2(n13305), .ZN(n16367) );
  NAND2_X1 U3878 ( .A1(n4805), .A2(n6938), .ZN(n31025) );
  INV_X1 U3885 ( .I(n10739), .ZN(n13691) );
  NAND2_X1 U3887 ( .A1(n10739), .A2(n19389), .ZN(n7820) );
  NAND2_X1 U3888 ( .A1(n23506), .A2(n23580), .ZN(n13833) );
  NAND2_X1 U3890 ( .A1(n18453), .A2(n7023), .ZN(n34819) );
  CLKBUF_X2 U3898 ( .I(n7023), .Z(n1432) );
  NAND2_X1 U3908 ( .A1(n13424), .A2(n209), .ZN(n7849) );
  NAND2_X1 U3913 ( .A1(n14752), .A2(n38491), .ZN(n27013) );
  CLKBUF_X2 U3914 ( .I(n14752), .Z(n7619) );
  BUF_X2 U3915 ( .I(Key[47]), .Z(n30169) );
  INV_X1 U3917 ( .I(n16989), .ZN(n3733) );
  INV_X2 U3918 ( .I(n3840), .ZN(n14027) );
  NAND2_X1 U3922 ( .A1(n3840), .A2(n18303), .ZN(n16989) );
  AND2_X1 U3929 ( .A1(n3840), .A2(n1338), .Z(n1778) );
  OR2_X1 U3930 ( .A1(n5028), .A2(n28729), .Z(n14497) );
  INV_X1 U3934 ( .I(n28729), .ZN(n15649) );
  INV_X1 U3935 ( .I(n28729), .ZN(n38998) );
  NAND2_X1 U3940 ( .A1(n21770), .A2(n21768), .ZN(n21605) );
  CLKBUF_X4 U3946 ( .I(n21768), .Z(n19546) );
  NOR2_X1 U3947 ( .A1(n21768), .A2(n21770), .ZN(n16052) );
  INV_X2 U3953 ( .I(n21768), .ZN(n19084) );
  CLKBUF_X2 U3954 ( .I(n9501), .Z(n31721) );
  INV_X1 U3955 ( .I(n9501), .ZN(n10563) );
  NAND2_X1 U3956 ( .A1(n425), .A2(n25894), .ZN(n5276) );
  BUF_X2 U3957 ( .I(n25894), .Z(n30900) );
  INV_X2 U3962 ( .I(n25894), .ZN(n1103) );
  NOR2_X1 U3964 ( .A1(n15677), .A2(n25894), .ZN(n25738) );
  NAND3_X1 U3971 ( .A1(n28383), .A2(n20494), .A3(n31855), .ZN(n28384) );
  NAND2_X1 U3972 ( .A1(n31854), .A2(n31855), .ZN(n30636) );
  NAND2_X1 U3977 ( .A1(n29675), .A2(n29683), .ZN(n29682) );
  INV_X1 U3980 ( .I(n29683), .ZN(n29677) );
  OR2_X1 U3983 ( .A1(n21885), .A2(n15839), .Z(n13858) );
  NOR2_X1 U3986 ( .A1(n18246), .A2(n11729), .ZN(n37703) );
  NAND3_X1 U3987 ( .A1(n9699), .A2(n8569), .A3(n20309), .ZN(n22830) );
  NAND2_X1 U3989 ( .A1(n20309), .A2(n19000), .ZN(n22934) );
  INV_X2 U3990 ( .I(n20313), .ZN(n24172) );
  NAND2_X1 U3993 ( .A1(n20312), .A2(n20313), .ZN(n263) );
  INV_X2 U3995 ( .I(n36840), .ZN(n7588) );
  AOI22_X1 U4005 ( .A1(n27255), .A2(n36840), .B1(n18716), .B2(n18195), .ZN(
        n27256) );
  NAND2_X1 U4014 ( .A1(n36840), .A2(n39583), .ZN(n27049) );
  NAND2_X1 U4017 ( .A1(n15911), .A2(n962), .ZN(n38001) );
  OAI21_X1 U4024 ( .A1(n8942), .A2(n962), .B(n5581), .ZN(n5582) );
  INV_X2 U4026 ( .I(n14415), .ZN(n1094) );
  NOR2_X1 U4027 ( .A1(n14415), .A2(n14380), .ZN(n34249) );
  AOI21_X1 U4034 ( .A1(n11636), .A2(n14415), .B(n8413), .ZN(n8917) );
  OAI21_X1 U4036 ( .A1(n39415), .A2(n21043), .B(n7658), .ZN(n4128) );
  OAI22_X1 U4037 ( .A1(n1034), .A2(n24425), .B1(n17456), .B2(n21043), .ZN(n298) );
  OAI21_X1 U4053 ( .A1(n21043), .A2(n38561), .B(n17456), .ZN(n31252) );
  NAND2_X1 U4057 ( .A1(n21043), .A2(n37580), .ZN(n17062) );
  NAND2_X1 U4061 ( .A1(n20643), .A2(n19518), .ZN(n33015) );
  INV_X1 U4063 ( .I(n35376), .ZN(n23730) );
  AOI21_X1 U4065 ( .A1(n24738), .A2(n31722), .B(n24737), .ZN(n35128) );
  NAND2_X1 U4069 ( .A1(n31722), .A2(n31679), .ZN(n16671) );
  NAND2_X1 U4071 ( .A1(n23535), .A2(n14759), .ZN(n23227) );
  NOR2_X1 U4072 ( .A1(n14759), .A2(n23535), .ZN(n20100) );
  INV_X1 U4074 ( .I(n14759), .ZN(n23538) );
  NAND2_X1 U4075 ( .A1(n3907), .A2(n22113), .ZN(n10154) );
  NAND3_X1 U4077 ( .A1(n1049), .A2(n3907), .A3(n38448), .ZN(n11456) );
  NAND3_X1 U4078 ( .A1(n10930), .A2(n13191), .A3(n3907), .ZN(n38484) );
  CLKBUF_X2 U4080 ( .I(n6285), .Z(n33656) );
  INV_X1 U4081 ( .I(n18160), .ZN(n5564) );
  AND2_X2 U4083 ( .A1(n37922), .A2(n38229), .Z(n37062) );
  INV_X1 U4088 ( .I(n10482), .ZN(n14089) );
  INV_X2 U4091 ( .I(n4574), .ZN(n39527) );
  AND3_X1 U4096 ( .A1(n15455), .A2(n1046), .A3(n20267), .Z(n37063) );
  CLKBUF_X4 U4097 ( .I(n4524), .Z(n38408) );
  INV_X2 U4099 ( .I(n4524), .ZN(n38611) );
  INV_X2 U4104 ( .I(n15299), .ZN(n32424) );
  OR2_X2 U4105 ( .A1(n7577), .A2(n15299), .Z(n37064) );
  INV_X2 U4114 ( .I(n15933), .ZN(n24394) );
  AND2_X1 U4115 ( .A1(n24090), .A2(n24442), .Z(n37066) );
  AND2_X2 U4116 ( .A1(n33616), .A2(n39191), .Z(n37067) );
  NAND2_X2 U4119 ( .A1(n31143), .A2(n39731), .ZN(n25085) );
  OR2_X1 U4120 ( .A1(n25513), .A2(n25540), .Z(n37069) );
  INV_X2 U4122 ( .I(n17624), .ZN(n32193) );
  AND3_X1 U4124 ( .A1(n178), .A2(n25359), .A3(n33130), .Z(n37070) );
  AND2_X1 U4125 ( .A1(n25367), .A2(n25540), .Z(n37071) );
  INV_X2 U4126 ( .I(n25288), .ZN(n25989) );
  CLKBUF_X4 U4130 ( .I(n25288), .Z(n38548) );
  INV_X1 U4131 ( .I(n17803), .ZN(n17951) );
  BUF_X4 U4133 ( .I(n17803), .Z(n38168) );
  AND2_X1 U4136 ( .A1(n9859), .A2(n25887), .Z(n37073) );
  OR2_X2 U4137 ( .A1(n38939), .A2(n38755), .Z(n37075) );
  INV_X4 U4140 ( .I(n13973), .ZN(n1891) );
  INV_X2 U4141 ( .I(n36050), .ZN(n38690) );
  OR2_X1 U4142 ( .A1(n27292), .A2(n6191), .Z(n37077) );
  INV_X2 U4143 ( .I(n19995), .ZN(n37754) );
  BUF_X2 U4144 ( .I(n27910), .Z(n580) );
  OR2_X1 U4146 ( .A1(n19541), .A2(n5525), .Z(n37078) );
  XOR2_X1 U4151 ( .A1(n3206), .A2(n35438), .Z(n37079) );
  INV_X4 U4160 ( .I(n7063), .ZN(n39724) );
  INV_X2 U4161 ( .I(n5028), .ZN(n30805) );
  INV_X1 U4168 ( .I(n14448), .ZN(n154) );
  OR2_X2 U4170 ( .A1(n28748), .A2(n28622), .Z(n37080) );
  AND2_X2 U4173 ( .A1(n32077), .A2(n6264), .Z(n37081) );
  NAND2_X2 U4177 ( .A1(n2868), .A2(n39112), .ZN(n35657) );
  INV_X2 U4178 ( .I(n20673), .ZN(n19992) );
  CLKBUF_X4 U4181 ( .I(n20673), .Z(n481) );
  NAND2_X2 U4188 ( .A1(n2784), .A2(n2789), .ZN(n38147) );
  OR2_X2 U4189 ( .A1(n35551), .A2(n18288), .Z(n37083) );
  NAND2_X1 U4190 ( .A1(n17861), .A2(n20255), .ZN(n21972) );
  INV_X2 U4195 ( .I(n20255), .ZN(n20996) );
  BUF_X2 U4199 ( .I(n20255), .Z(n7613) );
  AND2_X2 U4201 ( .A1(n11573), .A2(n30221), .Z(n9708) );
  OR2_X2 U4204 ( .A1(n20541), .A2(n30221), .Z(n30225) );
  OR2_X2 U4206 ( .A1(n14833), .A2(n5796), .Z(n5795) );
  CLKBUF_X4 U4211 ( .I(n9387), .Z(n32039) );
  AOI21_X1 U4212 ( .A1(n21726), .A2(n21727), .B(n18293), .ZN(n18979) );
  INV_X2 U4218 ( .I(n15868), .ZN(n18408) );
  NOR2_X1 U4223 ( .A1(n22274), .A2(n15868), .ZN(n15280) );
  NAND2_X1 U4224 ( .A1(n39059), .A2(n36908), .ZN(n24687) );
  OAI22_X1 U4227 ( .A1(n33151), .A2(n14265), .B1(n39059), .B2(n36908), .ZN(
        n8296) );
  OR2_X2 U4233 ( .A1(n33230), .A2(n36908), .Z(n37999) );
  OR2_X2 U4237 ( .A1(n7067), .A2(n7066), .Z(n31290) );
  NOR2_X2 U4240 ( .A1(n22146), .A2(n22240), .ZN(n22145) );
  CLKBUF_X12 U4241 ( .I(n734), .Z(n35216) );
  CLKBUF_X12 U4247 ( .I(n734), .Z(n7583) );
  INV_X2 U4251 ( .I(n29497), .ZN(n2954) );
  NAND2_X1 U4252 ( .A1(n29389), .A2(n29497), .ZN(n39274) );
  OAI21_X1 U4256 ( .A1(n29389), .A2(n19151), .B(n29497), .ZN(n15876) );
  NAND2_X1 U4257 ( .A1(n29459), .A2(n29497), .ZN(n29501) );
  NOR2_X1 U4258 ( .A1(n5127), .A2(n18929), .ZN(n10092) );
  INV_X2 U4264 ( .I(n18929), .ZN(n6128) );
  INV_X2 U4275 ( .I(n10047), .ZN(n15455) );
  INV_X1 U4276 ( .I(n35431), .ZN(n22299) );
  OAI21_X1 U4279 ( .A1(n2341), .A2(n19422), .B(n1029), .ZN(n20929) );
  INV_X1 U4282 ( .I(n19422), .ZN(n1576) );
  INV_X1 U4283 ( .I(n31367), .ZN(n950) );
  NAND3_X1 U4286 ( .A1(n24416), .A2(n37355), .A3(n31213), .ZN(n17979) );
  INV_X2 U4287 ( .I(n24416), .ZN(n19679) );
  CLKBUF_X4 U4296 ( .I(n24366), .Z(n32683) );
  INV_X2 U4297 ( .I(n24366), .ZN(n9135) );
  NAND2_X1 U4299 ( .A1(n24366), .A2(n37107), .ZN(n34424) );
  NOR2_X1 U4303 ( .A1(n2084), .A2(n2085), .ZN(n33775) );
  BUF_X2 U4305 ( .I(n37047), .Z(n36556) );
  INV_X1 U4310 ( .I(n37047), .ZN(n24426) );
  AND2_X2 U4315 ( .A1(n29377), .A2(n20726), .Z(n34973) );
  OR2_X2 U4316 ( .A1(n36357), .A2(n39456), .Z(n39535) );
  AND2_X2 U4317 ( .A1(n33510), .A2(n36357), .Z(n10288) );
  AND2_X2 U4318 ( .A1(n20669), .A2(n12012), .Z(n33633) );
  INV_X1 U4321 ( .I(n21848), .ZN(n6198) );
  OAI22_X1 U4322 ( .A1(n2643), .A2(n19133), .B1(n21944), .B2(n21605), .ZN(
        n38836) );
  OR2_X2 U4323 ( .A1(n5656), .A2(n10455), .Z(n12245) );
  NAND2_X1 U4325 ( .A1(n18850), .A2(n38704), .ZN(n32013) );
  NAND2_X1 U4326 ( .A1(n18850), .A2(n23310), .ZN(n23606) );
  INV_X1 U4327 ( .I(n18850), .ZN(n1636) );
  NAND2_X1 U4329 ( .A1(n33168), .A2(n18998), .ZN(n15852) );
  INV_X1 U4330 ( .I(n33168), .ZN(n32457) );
  AOI21_X1 U4331 ( .A1(n20376), .A2(n33168), .B(n7131), .ZN(n21977) );
  NOR2_X1 U4332 ( .A1(n9422), .A2(n33168), .ZN(n7216) );
  INV_X1 U4336 ( .I(n20662), .ZN(n28532) );
  NAND2_X1 U4339 ( .A1(n24565), .A2(n32637), .ZN(n24566) );
  AND3_X2 U4341 ( .A1(n24557), .A2(n24812), .A3(n32637), .Z(n39713) );
  NAND2_X1 U4344 ( .A1(n32637), .A2(n24565), .ZN(n36618) );
  OAI22_X1 U4345 ( .A1(n7878), .A2(n10158), .B1(n19637), .B2(n19636), .ZN(
        n7877) );
  OAI21_X1 U4346 ( .A1(n19637), .A2(n4048), .B(n25387), .ZN(n17231) );
  INV_X1 U4347 ( .I(n19637), .ZN(n1255) );
  CLKBUF_X12 U4352 ( .I(n9824), .Z(n36683) );
  AND2_X2 U4354 ( .A1(n20194), .A2(n25694), .Z(n25195) );
  CLKBUF_X4 U4356 ( .I(n6355), .Z(n4743) );
  OAI21_X1 U4357 ( .A1(n21923), .A2(n9316), .B(n21924), .ZN(n38898) );
  CLKBUF_X12 U4358 ( .I(n13039), .Z(n37084) );
  INV_X1 U4359 ( .I(n32230), .ZN(n4956) );
  BUF_X2 U4367 ( .I(n32230), .Z(n32122) );
  OAI22_X1 U4368 ( .A1(n19382), .A2(n1595), .B1(n545), .B2(n1276), .ZN(n37967)
         );
  NAND2_X1 U4369 ( .A1(n1276), .A2(n5985), .ZN(n24102) );
  INV_X1 U4370 ( .I(n19112), .ZN(n21257) );
  CLKBUF_X12 U4373 ( .I(n2145), .Z(n38468) );
  INV_X1 U4375 ( .I(n3213), .ZN(n6543) );
  INV_X2 U4378 ( .I(n22484), .ZN(n33415) );
  CLKBUF_X4 U4379 ( .I(n21214), .Z(n7916) );
  OR2_X1 U4380 ( .A1(n24600), .A2(n18788), .Z(n9073) );
  BUF_X2 U4381 ( .I(n16489), .Z(n11696) );
  INV_X1 U4383 ( .I(n26435), .ZN(n10878) );
  INV_X1 U4386 ( .I(n20423), .ZN(n32427) );
  AND2_X1 U4387 ( .A1(n20423), .A2(n19867), .Z(n18587) );
  NOR2_X1 U4392 ( .A1(n26972), .A2(n20423), .ZN(n26815) );
  NAND2_X1 U4393 ( .A1(n20423), .A2(n858), .ZN(n15980) );
  INV_X1 U4399 ( .I(n18549), .ZN(n37487) );
  NAND2_X1 U4400 ( .A1(n19203), .A2(n18549), .ZN(n19352) );
  NAND2_X1 U4401 ( .A1(n27383), .A2(n18549), .ZN(n36797) );
  NOR2_X1 U4403 ( .A1(n1221), .A2(n18549), .ZN(n27026) );
  CLKBUF_X12 U4405 ( .I(n18507), .Z(n37085) );
  CLKBUF_X12 U4407 ( .I(n6347), .Z(n39010) );
  INV_X1 U4411 ( .I(n6347), .ZN(n2818) );
  NAND2_X1 U4414 ( .A1(n7644), .A2(n4576), .ZN(n19389) );
  NAND2_X1 U4416 ( .A1(n7379), .A2(n7644), .ZN(n31662) );
  NAND2_X1 U4420 ( .A1(n33287), .A2(n7644), .ZN(n16126) );
  NAND2_X2 U4422 ( .A1(n21479), .A2(n2157), .ZN(n2156) );
  CLKBUF_X12 U4432 ( .I(n38839), .Z(n37803) );
  INV_X2 U4435 ( .I(n38839), .ZN(n38302) );
  BUF_X2 U4437 ( .I(n15299), .Z(n6638) );
  INV_X1 U4438 ( .I(n3003), .ZN(n20799) );
  BUF_X2 U4446 ( .I(n3003), .Z(n31407) );
  NAND2_X1 U4453 ( .A1(n36058), .A2(n13300), .ZN(n24605) );
  INV_X2 U4454 ( .I(n26229), .ZN(n34495) );
  NAND2_X1 U4455 ( .A1(n4149), .A2(n17887), .ZN(n5371) );
  OR2_X2 U4460 ( .A1(n19594), .A2(n35246), .Z(n4340) );
  NOR2_X1 U4461 ( .A1(n19966), .A2(n19594), .ZN(n22793) );
  INV_X1 U4463 ( .I(n26048), .ZN(n1242) );
  NOR2_X1 U4468 ( .A1(n26048), .A2(n1524), .ZN(n5475) );
  BUF_X2 U4469 ( .I(n37232), .Z(n37086) );
  OAI21_X1 U4471 ( .A1(n4147), .A2(n12790), .B(n36263), .ZN(n31951) );
  NAND2_X1 U4476 ( .A1(n27133), .A2(n1225), .ZN(n31734) );
  NAND2_X1 U4478 ( .A1(n5027), .A2(n27133), .ZN(n10066) );
  INV_X1 U4480 ( .I(n36750), .ZN(n15909) );
  CLKBUF_X12 U4485 ( .I(n36750), .Z(n39116) );
  AOI22_X1 U4488 ( .A1(n37985), .A2(n30764), .B1(n9656), .B2(n24591), .ZN(n819) );
  INV_X2 U4490 ( .I(n30764), .ZN(n958) );
  NAND2_X1 U4493 ( .A1(n878), .A2(n33956), .ZN(n27900) );
  CLKBUF_X12 U4499 ( .I(n33956), .Z(n310) );
  INV_X1 U4500 ( .I(n5274), .ZN(n16663) );
  INV_X2 U4502 ( .I(n9802), .ZN(n1015) );
  NAND2_X1 U4504 ( .A1(n9802), .A2(n33997), .ZN(n32035) );
  AOI22_X1 U4508 ( .A1(n1015), .A2(n25860), .B1(n362), .B2(n9802), .ZN(n12712)
         );
  NOR2_X1 U4509 ( .A1(n1520), .A2(n9802), .ZN(n37309) );
  OAI21_X1 U4510 ( .A1(n14881), .A2(n31006), .B(n35895), .ZN(n14795) );
  OR2_X2 U4512 ( .A1(n37662), .A2(n25636), .Z(n25717) );
  CLKBUF_X2 U4516 ( .I(n25636), .Z(n9132) );
  CLKBUF_X12 U4517 ( .I(n33847), .Z(n37087) );
  BUF_X4 U4518 ( .I(n33847), .Z(n37088) );
  INV_X1 U4523 ( .I(n10782), .ZN(n20820) );
  OAI22_X1 U4532 ( .A1(n38211), .A2(n8251), .B1(n8253), .B2(n1082), .ZN(n2380)
         );
  AND2_X2 U4534 ( .A1(n25481), .A2(n19928), .Z(n20565) );
  INV_X1 U4536 ( .I(n7497), .ZN(n6451) );
  NOR2_X1 U4541 ( .A1(n1151), .A2(n7497), .ZN(n5876) );
  INV_X1 U4542 ( .I(n8972), .ZN(n37995) );
  AOI22_X1 U4543 ( .A1(n2837), .A2(n26030), .B1(n25923), .B2(n25962), .ZN(
        n38102) );
  OR2_X2 U4545 ( .A1(n19478), .A2(n25553), .Z(n25477) );
  OR2_X1 U4548 ( .A1(n19992), .A2(n29781), .Z(n19993) );
  INV_X1 U4552 ( .I(n25163), .ZN(n10273) );
  NOR2_X1 U4554 ( .A1(n1097), .A2(n4604), .ZN(n3359) );
  NAND2_X1 U4556 ( .A1(n4604), .A2(n38416), .ZN(n25768) );
  BUF_X2 U4557 ( .I(n4604), .Z(n34402) );
  CLKBUF_X12 U4559 ( .I(n24403), .Z(n37904) );
  OAI22_X1 U4560 ( .A1(n1032), .A2(n39055), .B1(n13555), .B2(n24403), .ZN(
        n33727) );
  NAND2_X1 U4563 ( .A1(n24403), .A2(n13443), .ZN(n12366) );
  AND3_X2 U4564 ( .A1(n20517), .A2(n24403), .A3(n13555), .Z(n33500) );
  NAND2_X1 U4566 ( .A1(n22240), .A2(n21214), .ZN(n22147) );
  INV_X1 U4567 ( .I(n22240), .ZN(n21821) );
  NAND2_X1 U4571 ( .A1(n9387), .A2(n10820), .ZN(n20034) );
  INV_X2 U4576 ( .I(n30210), .ZN(n30214) );
  NAND2_X1 U4577 ( .A1(n21802), .A2(n8899), .ZN(n22075) );
  OR2_X2 U4588 ( .A1(n20397), .A2(n8899), .Z(n3269) );
  INV_X2 U4589 ( .I(n15515), .ZN(n25527) );
  NOR2_X1 U4593 ( .A1(n39415), .A2(n9193), .ZN(n38349) );
  NAND3_X2 U4594 ( .A1(n7472), .A2(n7471), .A3(n27149), .ZN(n38277) );
  AOI22_X1 U4598 ( .A1(n50), .A2(n14448), .B1(n28732), .B2(n36623), .ZN(n15321) );
  NOR2_X1 U4599 ( .A1(n7712), .A2(n31612), .ZN(n23425) );
  INV_X1 U4605 ( .I(n31612), .ZN(n7008) );
  BUF_X2 U4608 ( .I(n31612), .Z(n4600) );
  NOR2_X1 U4610 ( .A1(n12331), .A2(n14817), .ZN(n22992) );
  INV_X2 U4611 ( .I(n12331), .ZN(n6674) );
  NAND2_X1 U4613 ( .A1(n22865), .A2(n12331), .ZN(n16638) );
  NAND2_X1 U4626 ( .A1(n31744), .A2(n21248), .ZN(n32546) );
  INV_X2 U4629 ( .I(n13029), .ZN(n23350) );
  NAND2_X1 U4634 ( .A1(n6590), .A2(n26109), .ZN(n14229) );
  INV_X2 U4635 ( .I(n6590), .ZN(n951) );
  NOR2_X1 U4636 ( .A1(n6590), .A2(n26109), .ZN(n37462) );
  NOR2_X1 U4642 ( .A1(n23303), .A2(n11970), .ZN(n23420) );
  OR2_X1 U4646 ( .A1(n29939), .A2(n1057), .Z(n34086) );
  CLKBUF_X12 U4648 ( .I(n28179), .Z(n18832) );
  INV_X1 U4661 ( .I(n28873), .ZN(n33715) );
  INV_X1 U4663 ( .I(n8003), .ZN(n39725) );
  OAI22_X1 U4664 ( .A1(n29571), .A2(n31899), .B1(n1393), .B2(n17262), .ZN(
        n29577) );
  OAI21_X1 U4666 ( .A1(n30629), .A2(n17400), .B(n25975), .ZN(n17002) );
  AOI22_X1 U4667 ( .A1(n5311), .A2(n27407), .B1(n27153), .B2(n27406), .ZN(
        n5085) );
  AOI22_X1 U4669 ( .A1(n27153), .A2(n27407), .B1(n2947), .B2(n1487), .ZN(
        n27405) );
  NAND2_X1 U4674 ( .A1(n17714), .A2(n28729), .ZN(n38123) );
  NAND2_X1 U4683 ( .A1(n36623), .A2(n28729), .ZN(n36633) );
  OAI21_X1 U4689 ( .A1(n28178), .A2(n28031), .B(n16559), .ZN(n20084) );
  OR2_X2 U4696 ( .A1(n27964), .A2(n33960), .Z(n21322) );
  AND2_X2 U4698 ( .A1(n33960), .A2(n27964), .Z(n4640) );
  NAND2_X1 U4701 ( .A1(n13995), .A2(n2047), .ZN(n23146) );
  NOR2_X1 U4703 ( .A1(n13995), .A2(n2047), .ZN(n23044) );
  INV_X2 U4705 ( .I(n13995), .ZN(n37791) );
  NOR2_X1 U4708 ( .A1(n23145), .A2(n13995), .ZN(n23148) );
  NOR2_X1 U4710 ( .A1(n27325), .A2(n35500), .ZN(n17985) );
  NAND2_X1 U4712 ( .A1(n17142), .A2(n27325), .ZN(n37512) );
  NAND3_X1 U4718 ( .A1(n11910), .A2(n17142), .A3(n27325), .ZN(n38734) );
  AOI21_X1 U4719 ( .A1(n12326), .A2(n27325), .B(n11910), .ZN(n27329) );
  NOR2_X1 U4720 ( .A1(n12326), .A2(n27325), .ZN(n4253) );
  INV_X1 U4721 ( .I(n29041), .ZN(n5992) );
  INV_X1 U4722 ( .I(n26125), .ZN(n39661) );
  NOR2_X1 U4723 ( .A1(n14126), .A2(n30097), .ZN(n2489) );
  OAI21_X1 U4724 ( .A1(n32682), .A2(n38172), .B(n9686), .ZN(n4871) );
  INV_X2 U4726 ( .I(n9686), .ZN(n28736) );
  NAND2_X1 U4730 ( .A1(n9686), .A2(n17234), .ZN(n28547) );
  INV_X1 U4731 ( .I(n21754), .ZN(n21699) );
  NAND2_X1 U4732 ( .A1(n14493), .A2(n21754), .ZN(n21542) );
  BUF_X2 U4733 ( .I(n21754), .Z(n1372) );
  NAND2_X1 U4734 ( .A1(n26063), .A2(n25943), .ZN(n35679) );
  INV_X2 U4735 ( .I(n3874), .ZN(n4699) );
  NAND2_X1 U4738 ( .A1(n31367), .A2(n3874), .ZN(n25870) );
  NAND2_X1 U4739 ( .A1(n3669), .A2(n3874), .ZN(n17700) );
  NAND3_X1 U4745 ( .A1(n15577), .A2(n27305), .A3(n27304), .ZN(n10735) );
  OAI21_X1 U4747 ( .A1(n27305), .A2(n17166), .B(n35906), .ZN(n12072) );
  INV_X1 U4748 ( .I(n22669), .ZN(n35810) );
  OR2_X2 U4749 ( .A1(n20896), .A2(n34120), .Z(n12323) );
  INV_X2 U4750 ( .I(n27438), .ZN(n19719) );
  INV_X1 U4754 ( .I(n38981), .ZN(n23321) );
  CLKBUF_X4 U4757 ( .I(n38981), .Z(n16047) );
  AOI21_X1 U4758 ( .A1(n7424), .A2(n17072), .B(n14881), .ZN(n14796) );
  AOI21_X1 U4760 ( .A1(n7426), .A2(n34959), .B(n3708), .ZN(n7425) );
  NOR2_X2 U4761 ( .A1(n37070), .A2(n9482), .ZN(n9479) );
  INV_X1 U4762 ( .I(n26364), .ZN(n26366) );
  BUF_X2 U4764 ( .I(n26765), .Z(n26922) );
  OAI22_X1 U4765 ( .A1(n26765), .A2(n13543), .B1(n19371), .B2(n3606), .ZN(
        n39758) );
  INV_X2 U4766 ( .I(n180), .ZN(n1420) );
  NAND2_X1 U4767 ( .A1(n28616), .A2(n180), .ZN(n28615) );
  NOR2_X1 U4769 ( .A1(n6147), .A2(n14126), .ZN(n20099) );
  NOR2_X1 U4771 ( .A1(n30092), .A2(n6147), .ZN(n37356) );
  NAND2_X1 U4772 ( .A1(n6147), .A2(n31601), .ZN(n7600) );
  INV_X1 U4776 ( .I(n28972), .ZN(n4314) );
  NOR2_X1 U4777 ( .A1(n3434), .A2(n25800), .ZN(n32233) );
  NOR2_X1 U4779 ( .A1(n20031), .A2(n9862), .ZN(n2453) );
  NAND2_X1 U4787 ( .A1(n12952), .A2(n1145), .ZN(n38513) );
  NAND3_X1 U4791 ( .A1(n8260), .A2(n8261), .A3(n7542), .ZN(n37696) );
  NAND2_X1 U4798 ( .A1(n15135), .A2(n10171), .ZN(n27305) );
  INV_X2 U4799 ( .I(n10171), .ZN(n35332) );
  INV_X1 U4802 ( .I(n10611), .ZN(n25037) );
  AND3_X1 U4804 ( .A1(n1021), .A2(n17624), .A3(n11148), .Z(n25781) );
  OR2_X1 U4807 ( .A1(n11148), .A2(n15575), .Z(n37213) );
  OAI22_X1 U4813 ( .A1(n29723), .A2(n29717), .B1(n29710), .B2(n29709), .ZN(
        n32519) );
  NOR2_X1 U4814 ( .A1(n29723), .A2(n5951), .ZN(n39101) );
  AND2_X2 U4816 ( .A1(n22879), .A2(n5891), .Z(n6009) );
  OR2_X2 U4820 ( .A1(n22879), .A2(n5891), .Z(n12032) );
  CLKBUF_X12 U4821 ( .I(n3116), .Z(n37092) );
  BUF_X2 U4822 ( .I(n3116), .Z(n37093) );
  AOI21_X1 U4827 ( .A1(n38068), .A2(n4192), .B(n27446), .ZN(n32940) );
  NAND2_X1 U4833 ( .A1(n27446), .A2(n38187), .ZN(n5630) );
  INV_X1 U4836 ( .I(n17351), .ZN(n17350) );
  CLKBUF_X12 U4839 ( .I(n11627), .Z(n531) );
  NAND2_X1 U4843 ( .A1(n23566), .A2(n3713), .ZN(n5792) );
  CLKBUF_X4 U4849 ( .I(n33734), .Z(n2192) );
  INV_X1 U4857 ( .I(n33734), .ZN(n4243) );
  INV_X1 U4858 ( .I(n21488), .ZN(n19699) );
  NAND2_X1 U4860 ( .A1(n2765), .A2(n8679), .ZN(n22144) );
  INV_X4 U4866 ( .I(n1812), .ZN(n18253) );
  OAI21_X1 U4872 ( .A1(n38973), .A2(n39059), .B(n33230), .ZN(n8355) );
  NAND2_X1 U4875 ( .A1(n36908), .A2(n33230), .ZN(n13554) );
  NAND2_X1 U4876 ( .A1(n33230), .A2(n24761), .ZN(n14338) );
  INV_X2 U4881 ( .I(n23482), .ZN(n6303) );
  CLKBUF_X4 U4891 ( .I(n23482), .Z(n9078) );
  OAI21_X1 U4893 ( .A1(n1630), .A2(n38244), .B(n23586), .ZN(n34585) );
  INV_X2 U4897 ( .I(n12617), .ZN(n38244) );
  AND3_X2 U4900 ( .A1(n38976), .A2(n22196), .A3(n30800), .Z(n14269) );
  OAI22_X1 U4901 ( .A1(n38976), .A2(n1327), .B1(n8520), .B2(n22287), .ZN(n5557) );
  INV_X2 U4902 ( .I(n38976), .ZN(n1328) );
  OAI21_X1 U4904 ( .A1(n5396), .A2(n39227), .B(n13598), .ZN(n5397) );
  INV_X1 U4906 ( .I(n19370), .ZN(n21517) );
  CLKBUF_X12 U4920 ( .I(n19370), .Z(n17534) );
  OR3_X2 U4923 ( .A1(n20207), .A2(n9945), .A3(n24116), .Z(n4687) );
  AND2_X2 U4924 ( .A1(n24287), .A2(n20207), .Z(n11132) );
  AOI21_X1 U4926 ( .A1(n14423), .A2(n4239), .B(n34813), .ZN(n2907) );
  OR2_X2 U4936 ( .A1(n20449), .A2(n12100), .Z(n22990) );
  AND2_X2 U4940 ( .A1(n3861), .A2(n2858), .Z(n29852) );
  INV_X1 U4944 ( .I(n17758), .ZN(n26319) );
  NOR2_X1 U4946 ( .A1(n18502), .A2(n29438), .ZN(n17293) );
  NOR2_X1 U4948 ( .A1(n29439), .A2(n29438), .ZN(n29433) );
  INV_X1 U4952 ( .I(n31944), .ZN(n23450) );
  NAND2_X1 U4954 ( .A1(n31944), .A2(n11678), .ZN(n23394) );
  AND2_X2 U4956 ( .A1(n11585), .A2(n11586), .Z(n18193) );
  NAND3_X1 U4958 ( .A1(n21847), .A2(n19392), .A3(n21668), .ZN(n16653) );
  AOI21_X1 U4959 ( .A1(n19517), .A2(n18219), .B(n21847), .ZN(n6101) );
  NOR2_X1 U4966 ( .A1(n20538), .A2(n20342), .ZN(n2466) );
  NAND2_X1 U4970 ( .A1(n5450), .A2(n4424), .ZN(n3681) );
  AOI21_X1 U4972 ( .A1(n2480), .A2(n5450), .B(n18567), .ZN(n4045) );
  NAND2_X1 U4975 ( .A1(n5450), .A2(n14833), .ZN(n22256) );
  INV_X1 U4976 ( .I(n5450), .ZN(n22063) );
  NOR3_X1 U4981 ( .A1(n16094), .A2(n23477), .A3(n23473), .ZN(n17388) );
  NAND2_X1 U4986 ( .A1(n16094), .A2(n1139), .ZN(n12870) );
  NAND2_X1 U4990 ( .A1(n34558), .A2(n16094), .ZN(n23475) );
  OR2_X2 U4991 ( .A1(n36442), .A2(n16094), .Z(n8432) );
  NAND2_X1 U5004 ( .A1(n25583), .A2(n24896), .ZN(n20295) );
  INV_X1 U5007 ( .I(n25191), .ZN(n34788) );
  NAND3_X1 U5023 ( .A1(n28812), .A2(n33577), .A3(n19759), .ZN(n8913) );
  OR2_X2 U5025 ( .A1(n9845), .A2(n28231), .Z(n27970) );
  OR2_X2 U5029 ( .A1(n10216), .A2(n33786), .Z(n8027) );
  INV_X2 U5031 ( .I(n37016), .ZN(n32045) );
  INV_X1 U5032 ( .I(n9916), .ZN(n14132) );
  CLKBUF_X12 U5036 ( .I(n22223), .Z(n39284) );
  BUF_X4 U5040 ( .I(n21814), .Z(n19768) );
  CLKBUF_X12 U5047 ( .I(n29005), .Z(n621) );
  INV_X1 U5052 ( .I(n18399), .ZN(n33243) );
  CLKBUF_X12 U5053 ( .I(n13794), .Z(n36426) );
  OAI21_X1 U5059 ( .A1(n31845), .A2(n39268), .B(n24618), .ZN(n39562) );
  NAND2_X1 U5060 ( .A1(n37624), .A2(n39268), .ZN(n24534) );
  AOI21_X1 U5063 ( .A1(n31845), .A2(n39268), .B(n1026), .ZN(n6187) );
  NAND2_X1 U5076 ( .A1(n25813), .A2(n33909), .ZN(n35671) );
  INV_X1 U5080 ( .I(n25813), .ZN(n32510) );
  BUF_X4 U5083 ( .I(n22623), .Z(n37094) );
  CLKBUF_X4 U5084 ( .I(n24053), .Z(n38813) );
  NAND2_X1 U5087 ( .A1(n28463), .A2(n28464), .ZN(n1815) );
  INV_X2 U5093 ( .I(n28464), .ZN(n28637) );
  NAND3_X1 U5099 ( .A1(n38600), .A2(n34558), .A3(n36442), .ZN(n22681) );
  INV_X1 U5101 ( .I(n36442), .ZN(n20343) );
  NAND2_X1 U5102 ( .A1(n36442), .A2(n23473), .ZN(n11186) );
  CLKBUF_X4 U5103 ( .I(n26272), .Z(n26979) );
  NAND2_X1 U5106 ( .A1(n37341), .A2(n12633), .ZN(n39343) );
  OAI22_X1 U5107 ( .A1(n33151), .A2(n12633), .B1(n14857), .B2(n36908), .ZN(
        n13002) );
  INV_X1 U5117 ( .I(n17583), .ZN(n14968) );
  NAND2_X1 U5127 ( .A1(n17583), .A2(n28330), .ZN(n17031) );
  OR2_X2 U5128 ( .A1(n5732), .A2(n962), .Z(n8769) );
  AND2_X2 U5133 ( .A1(n8628), .A2(n5732), .Z(n8508) );
  BUF_X1 U5136 ( .I(n21885), .Z(n36754) );
  NOR3_X1 U5146 ( .A1(n34977), .A2(n27211), .A3(n8412), .ZN(n36407) );
  NAND2_X1 U5149 ( .A1(n19719), .A2(n8412), .ZN(n27097) );
  CLKBUF_X4 U5150 ( .I(n8412), .Z(n7494) );
  NAND2_X1 U5168 ( .A1(n7852), .A2(n36082), .ZN(n24768) );
  AND2_X1 U5175 ( .A1(n7852), .A2(n24764), .Z(n39099) );
  OAI22_X1 U5183 ( .A1(n21591), .A2(n21592), .B1(n38480), .B2(n21576), .ZN(
        n20585) );
  NOR3_X1 U5184 ( .A1(n8735), .A2(n37934), .A3(n24406), .ZN(n37551) );
  INV_X1 U5186 ( .I(n6756), .ZN(n30534) );
  AOI21_X1 U5191 ( .A1(n24126), .A2(n19484), .B(n6756), .ZN(n24127) );
  NOR2_X1 U5192 ( .A1(n23516), .A2(n23517), .ZN(n2175) );
  OAI22_X1 U5198 ( .A1(n7049), .A2(n18475), .B1(n23516), .B2(n39001), .ZN(
        n38024) );
  OR2_X2 U5202 ( .A1(n12950), .A2(n35954), .Z(n24206) );
  CLKBUF_X12 U5209 ( .I(n17397), .Z(n33646) );
  NAND2_X1 U5210 ( .A1(n17397), .A2(n28207), .ZN(n28361) );
  INV_X2 U5224 ( .I(n17397), .ZN(n28723) );
  BUF_X4 U5225 ( .I(n35465), .Z(n37096) );
  INV_X1 U5228 ( .I(n34685), .ZN(n25857) );
  NOR2_X1 U5232 ( .A1(n34685), .A2(n10404), .ZN(n34206) );
  AND3_X2 U5234 ( .A1(n15796), .A2(n25849), .A3(n34685), .Z(n12063) );
  CLKBUF_X12 U5240 ( .I(n18211), .Z(n5021) );
  NAND2_X1 U5241 ( .A1(n24765), .A2(n24764), .ZN(n24766) );
  AND2_X2 U5242 ( .A1(n26195), .A2(n35750), .Z(n14667) );
  NAND2_X1 U5244 ( .A1(n35750), .A2(n5089), .ZN(n34842) );
  OR2_X2 U5248 ( .A1(n26643), .A2(n26932), .Z(n26547) );
  NAND3_X1 U5251 ( .A1(n33352), .A2(n26933), .A3(n26932), .ZN(n33383) );
  INV_X1 U5254 ( .I(n26932), .ZN(n35912) );
  AND2_X2 U5258 ( .A1(n26932), .A2(n37235), .Z(n14485) );
  BUF_X1 U5260 ( .I(n26818), .Z(n19353) );
  NAND2_X1 U5266 ( .A1(n10404), .A2(n25887), .ZN(n26072) );
  NOR2_X1 U5273 ( .A1(n9859), .A2(n25887), .ZN(n26071) );
  OAI22_X1 U5274 ( .A1(n23342), .A2(n23430), .B1(n15787), .B2(n23343), .ZN(
        n1829) );
  NAND2_X1 U5281 ( .A1(n1628), .A2(n23430), .ZN(n3506) );
  NOR2_X1 U5288 ( .A1(n9685), .A2(n22092), .ZN(n22094) );
  NAND2_X1 U5289 ( .A1(n1152), .A2(n22092), .ZN(n22205) );
  NOR2_X1 U5292 ( .A1(n4190), .A2(n6904), .ZN(n17645) );
  OAI21_X1 U5293 ( .A1(n6904), .A2(n26125), .B(n5098), .ZN(n38783) );
  NAND3_X1 U5294 ( .A1(n39454), .A2(n6904), .A3(n4516), .ZN(n26010) );
  NAND2_X1 U5296 ( .A1(n39826), .A2(n27389), .ZN(n27167) );
  CLKBUF_X12 U5309 ( .I(n19478), .Z(n31580) );
  BUF_X2 U5311 ( .I(n25418), .Z(n19495) );
  NOR2_X1 U5314 ( .A1(n35260), .A2(n25418), .ZN(n25597) );
  AOI21_X1 U5317 ( .A1(n10623), .A2(n3840), .B(n3086), .ZN(n3085) );
  INV_X2 U5318 ( .I(n23076), .ZN(n23181) );
  CLKBUF_X12 U5322 ( .I(n26668), .Z(n19331) );
  INV_X1 U5323 ( .I(n26668), .ZN(n26973) );
  AND2_X2 U5324 ( .A1(n38901), .A2(n26668), .Z(n33006) );
  NAND2_X1 U5327 ( .A1(n26178), .A2(n26701), .ZN(n4641) );
  NOR2_X1 U5329 ( .A1(n23076), .A2(n23077), .ZN(n787) );
  NOR2_X1 U5331 ( .A1(n33933), .A2(n23076), .ZN(n9841) );
  NOR2_X1 U5336 ( .A1(n15641), .A2(n39424), .ZN(n21109) );
  NOR2_X1 U5339 ( .A1(n27221), .A2(n39424), .ZN(n4627) );
  INV_X1 U5341 ( .I(n39424), .ZN(n39531) );
  AOI21_X1 U5346 ( .A1(n27292), .A2(n39424), .B(n5588), .ZN(n4700) );
  NAND2_X1 U5347 ( .A1(n28748), .A2(n28622), .ZN(n28747) );
  INV_X2 U5348 ( .I(n28622), .ZN(n34244) );
  NAND2_X1 U5349 ( .A1(n24829), .A2(n24802), .ZN(n10161) );
  NOR2_X1 U5350 ( .A1(n24829), .A2(n38194), .ZN(n24572) );
  NAND2_X1 U5358 ( .A1(n2018), .A2(n24829), .ZN(n10160) );
  INV_X1 U5360 ( .I(n17405), .ZN(n5266) );
  INV_X4 U5369 ( .I(n29617), .ZN(n35405) );
  NAND2_X1 U5370 ( .A1(n28681), .A2(n28720), .ZN(n2788) );
  NOR2_X1 U5378 ( .A1(n28720), .A2(n28722), .ZN(n37560) );
  INV_X1 U5382 ( .I(n28720), .ZN(n28721) );
  AND2_X2 U5383 ( .A1(n862), .A2(n867), .Z(n13489) );
  CLKBUF_X4 U5387 ( .I(n867), .Z(n2451) );
  NAND2_X1 U5388 ( .A1(n32046), .A2(n32566), .ZN(n38068) );
  INV_X1 U5391 ( .I(n32566), .ZN(n16782) );
  INV_X1 U5398 ( .I(n15135), .ZN(n27586) );
  BUF_X2 U5400 ( .I(n15135), .Z(n4781) );
  NAND3_X1 U5405 ( .A1(n16181), .A2(n16071), .A3(n17624), .ZN(n16070) );
  INV_X1 U5407 ( .I(n15754), .ZN(n15751) );
  OAI21_X1 U5412 ( .A1(n30024), .A2(n30022), .B(n8039), .ZN(n30011) );
  NAND2_X1 U5414 ( .A1(n31371), .A2(n13151), .ZN(n15602) );
  NAND2_X1 U5416 ( .A1(n2534), .A2(n11034), .ZN(n35099) );
  INV_X2 U5418 ( .I(n11034), .ZN(n36099) );
  OR3_X2 U5426 ( .A1(n24883), .A2(n19499), .A3(n18788), .Z(n24681) );
  NOR2_X1 U5428 ( .A1(n24753), .A2(n18788), .ZN(n32099) );
  INV_X1 U5429 ( .I(n18788), .ZN(n24680) );
  NAND2_X1 U5432 ( .A1(n18788), .A2(n6756), .ZN(n5137) );
  OAI22_X1 U5435 ( .A1(n9066), .A2(n15903), .B1(n20839), .B2(n24296), .ZN(
        n37634) );
  INV_X1 U5436 ( .I(n16864), .ZN(n39468) );
  INV_X1 U5438 ( .I(n25303), .ZN(n12441) );
  INV_X1 U5439 ( .I(n24741), .ZN(n25386) );
  OR2_X2 U5440 ( .A1(n18722), .A2(n32820), .Z(n3215) );
  INV_X2 U5441 ( .I(n29284), .ZN(n19090) );
  OR2_X2 U5447 ( .A1(n11699), .A2(n10534), .Z(n15968) );
  NAND2_X1 U5451 ( .A1(n21882), .A2(n21883), .ZN(n21576) );
  NAND3_X1 U5455 ( .A1(n896), .A2(n2465), .A3(n11968), .ZN(n37644) );
  AOI21_X1 U5457 ( .A1(n30177), .A2(n20342), .B(n30183), .ZN(n7318) );
  CLKBUF_X2 U5459 ( .I(n16309), .Z(n39025) );
  INV_X1 U5465 ( .I(n28365), .ZN(n5738) );
  CLKBUF_X1 U5466 ( .I(n20597), .Z(n39363) );
  INV_X1 U5468 ( .I(n28615), .ZN(n32703) );
  CLKBUF_X1 U5473 ( .I(n5383), .Z(n32178) );
  NAND2_X1 U5478 ( .A1(n310), .A2(n16461), .ZN(n4503) );
  CLKBUF_X8 U5479 ( .I(n39126), .Z(n37671) );
  CLKBUF_X1 U5481 ( .I(n36463), .Z(n39786) );
  CLKBUF_X2 U5486 ( .I(n8078), .Z(n38762) );
  CLKBUF_X2 U5488 ( .I(n18860), .Z(n38419) );
  INV_X2 U5492 ( .I(n31683), .ZN(n38877) );
  NAND2_X1 U5494 ( .A1(n37654), .A2(n37653), .ZN(n37652) );
  NOR2_X1 U5497 ( .A1(n2923), .A2(n11765), .ZN(n37801) );
  INV_X2 U5498 ( .I(n18195), .ZN(n9633) );
  NOR2_X1 U5499 ( .A1(n27071), .A2(n36989), .ZN(n37384) );
  INV_X2 U5502 ( .I(n27292), .ZN(n38488) );
  NAND2_X1 U5503 ( .A1(n26762), .A2(n26761), .ZN(n37826) );
  CLKBUF_X1 U5510 ( .I(n5218), .Z(n39262) );
  NAND2_X1 U5512 ( .A1(n15196), .A2(n2081), .ZN(n32799) );
  OR3_X1 U5513 ( .A1(n38002), .A2(n1092), .A3(n37103), .Z(n36112) );
  BUF_X2 U5514 ( .I(n26724), .Z(n38928) );
  NOR2_X1 U5521 ( .A1(n7725), .A2(n7516), .ZN(n26798) );
  INV_X4 U5526 ( .I(n13770), .ZN(n37098) );
  CLKBUF_X2 U5529 ( .I(n26185), .Z(n39507) );
  AND2_X1 U5533 ( .A1(n1518), .A2(n1017), .Z(n37172) );
  AOI21_X1 U5534 ( .A1(n11552), .A2(n18406), .B(n9413), .ZN(n11551) );
  BUF_X2 U5538 ( .I(n25860), .Z(n36819) );
  BUF_X2 U5541 ( .I(n25971), .Z(n39248) );
  CLKBUF_X1 U5546 ( .I(n9833), .Z(n39165) );
  INV_X1 U5547 ( .I(n38004), .ZN(n20628) );
  NAND2_X1 U5550 ( .A1(n12748), .A2(n25517), .ZN(n37339) );
  NOR2_X1 U5551 ( .A1(n18294), .A2(n16264), .ZN(n39251) );
  INV_X2 U5552 ( .I(n5042), .ZN(n38728) );
  CLKBUF_X2 U5553 ( .I(n13811), .Z(n38300) );
  NAND2_X1 U5554 ( .A1(n32775), .A2(n10938), .ZN(n25486) );
  CLKBUF_X2 U5556 ( .I(n25140), .Z(n39295) );
  INV_X2 U5560 ( .I(n20128), .ZN(n24832) );
  OAI21_X1 U5568 ( .A1(n32785), .A2(n24478), .B(n32784), .ZN(n37504) );
  NOR2_X1 U5576 ( .A1(n38349), .A2(n38561), .ZN(n38652) );
  INV_X1 U5580 ( .I(n20119), .ZN(n9723) );
  NAND2_X1 U5590 ( .A1(n24397), .A2(n24396), .ZN(n37710) );
  NOR2_X1 U5592 ( .A1(n38812), .A2(n24123), .ZN(n37891) );
  NAND2_X1 U5594 ( .A1(n39415), .A2(n38251), .ZN(n38250) );
  CLKBUF_X2 U5602 ( .I(n16366), .Z(n39504) );
  NAND2_X1 U5603 ( .A1(n39067), .A2(n17076), .ZN(n24081) );
  INV_X2 U5604 ( .I(n30311), .ZN(n39706) );
  BUF_X4 U5606 ( .I(n4880), .Z(n39415) );
  CLKBUF_X2 U5607 ( .I(n20384), .Z(n37896) );
  CLKBUF_X2 U5608 ( .I(n13395), .Z(n39636) );
  CLKBUF_X2 U5610 ( .I(n18301), .Z(n37842) );
  NAND2_X1 U5616 ( .A1(n38894), .A2(n38893), .ZN(n35753) );
  NAND2_X1 U5617 ( .A1(n38792), .A2(n38299), .ZN(n6520) );
  CLKBUF_X2 U5620 ( .I(n16013), .Z(n37923) );
  OAI21_X1 U5624 ( .A1(n10867), .A2(n2116), .B(n19319), .ZN(n13641) );
  CLKBUF_X2 U5626 ( .I(n17511), .Z(n34823) );
  NAND2_X1 U5628 ( .A1(n39601), .A2(n17009), .ZN(n7491) );
  CLKBUF_X2 U5630 ( .I(n23162), .Z(n19870) );
  NAND2_X1 U5634 ( .A1(n23082), .A2(n14442), .ZN(n38903) );
  INV_X1 U5642 ( .I(n14494), .ZN(n23173) );
  OR2_X1 U5649 ( .A1(n23189), .A2(n34200), .Z(n23192) );
  AND2_X1 U5651 ( .A1(n39075), .A2(n1149), .Z(n37189) );
  AOI21_X1 U5652 ( .A1(n20756), .A2(n33549), .B(n37911), .ZN(n38522) );
  BUF_X2 U5658 ( .I(n31202), .Z(n37938) );
  CLKBUF_X2 U5661 ( .I(n36281), .Z(n37775) );
  INV_X2 U5667 ( .I(n10463), .ZN(n22143) );
  CLKBUF_X2 U5668 ( .I(n33993), .Z(n38375) );
  OAI21_X1 U5671 ( .A1(n21942), .A2(n16128), .B(n19133), .ZN(n37399) );
  INV_X1 U5677 ( .I(n21422), .ZN(n20827) );
  INV_X1 U5678 ( .I(n19831), .ZN(n37112) );
  BUF_X2 U5681 ( .I(n14245), .Z(n39716) );
  INV_X1 U5686 ( .I(n19629), .ZN(n37109) );
  INV_X1 U5688 ( .I(n29879), .ZN(n37110) );
  NOR3_X1 U5696 ( .A1(n30147), .A2(n30146), .A3(n3896), .ZN(n39510) );
  NAND2_X1 U5701 ( .A1(n29547), .A2(n6252), .ZN(n9837) );
  NAND3_X1 U5703 ( .A1(n29505), .A2(n29504), .A3(n16083), .ZN(n38802) );
  NAND3_X1 U5705 ( .A1(n10409), .A2(n10410), .A3(n10513), .ZN(n37825) );
  OAI22_X1 U5708 ( .A1(n29608), .A2(n29607), .B1(n37258), .B2(n37430), .ZN(
        n29610) );
  NOR3_X1 U5710 ( .A1(n2205), .A2(n2507), .A3(n1054), .ZN(n39079) );
  INV_X1 U5714 ( .I(n30026), .ZN(n30025) );
  CLKBUF_X2 U5716 ( .I(n85), .Z(n34534) );
  INV_X2 U5722 ( .I(n29612), .ZN(n29627) );
  CLKBUF_X4 U5726 ( .I(n17996), .Z(n17997) );
  NAND2_X1 U5727 ( .A1(n37531), .A2(n30432), .ZN(n31499) );
  INV_X1 U5728 ( .I(n39006), .ZN(n39005) );
  NAND2_X1 U5738 ( .A1(n36994), .A2(n31279), .ZN(n37359) );
  INV_X4 U5753 ( .I(n18815), .ZN(n3700) );
  CLKBUF_X4 U5758 ( .I(n35551), .Z(n36207) );
  CLKBUF_X2 U5759 ( .I(n29598), .Z(n38420) );
  BUF_X2 U5763 ( .I(n10006), .Z(n31583) );
  INV_X1 U5764 ( .I(n29498), .ZN(n37376) );
  INV_X1 U5765 ( .I(n29694), .ZN(n37752) );
  CLKBUF_X2 U5768 ( .I(n11783), .Z(n39187) );
  INV_X4 U5769 ( .I(n18720), .ZN(n37099) );
  INV_X2 U5771 ( .I(n29863), .ZN(n29957) );
  BUF_X2 U5782 ( .I(n30221), .Z(n6938) );
  BUF_X4 U5783 ( .I(n6449), .Z(n6019) );
  BUF_X4 U5787 ( .I(n29312), .Z(n37100) );
  INV_X1 U5790 ( .I(n18623), .ZN(n39634) );
  BUF_X2 U5795 ( .I(n29054), .Z(n6661) );
  INV_X1 U5799 ( .I(n39391), .ZN(n37059) );
  CLKBUF_X2 U5802 ( .I(n6930), .Z(n38703) );
  CLKBUF_X2 U5808 ( .I(n28610), .Z(n38290) );
  CLKBUF_X2 U5811 ( .I(n12244), .Z(n39536) );
  NAND2_X1 U5812 ( .A1(n35875), .A2(n37615), .ZN(n32758) );
  CLKBUF_X2 U5814 ( .I(n18453), .Z(n38556) );
  NAND2_X1 U5815 ( .A1(n28561), .A2(n38858), .ZN(n38857) );
  NAND2_X1 U5818 ( .A1(n28335), .A2(n33647), .ZN(n38061) );
  NOR2_X1 U5819 ( .A1(n6017), .A2(n28473), .ZN(n39332) );
  OAI21_X1 U5830 ( .A1(n33100), .A2(n28758), .B(n13508), .ZN(n32273) );
  INV_X1 U5833 ( .I(n28061), .ZN(n37414) );
  NAND2_X1 U5837 ( .A1(n28430), .A2(n9586), .ZN(n37413) );
  NAND2_X1 U5842 ( .A1(n28553), .A2(n1431), .ZN(n28556) );
  INV_X1 U5844 ( .I(n28440), .ZN(n37579) );
  INV_X1 U5854 ( .I(n28360), .ZN(n20879) );
  INV_X1 U5861 ( .I(n34176), .ZN(n28395) );
  BUF_X4 U5867 ( .I(n28621), .Z(n11490) );
  CLKBUF_X2 U5868 ( .I(n15540), .Z(n38566) );
  CLKBUF_X4 U5872 ( .I(n20662), .Z(n11614) );
  AND2_X1 U5873 ( .A1(n11831), .A2(n7221), .Z(n35172) );
  CLKBUF_X2 U5879 ( .I(n33707), .Z(n39425) );
  CLKBUF_X2 U5881 ( .I(n18480), .Z(n37804) );
  CLKBUF_X2 U5883 ( .I(n38854), .Z(n38075) );
  CLKBUF_X2 U5885 ( .I(n28753), .Z(n37460) );
  INV_X1 U5887 ( .I(n38203), .ZN(n37484) );
  NAND2_X1 U5889 ( .A1(n37895), .A2(n11754), .ZN(n38391) );
  NAND2_X1 U5893 ( .A1(n37445), .A2(n13366), .ZN(n18224) );
  NAND2_X1 U5894 ( .A1(n8525), .A2(n8524), .ZN(n39180) );
  NAND2_X1 U5897 ( .A1(n15364), .A2(n16869), .ZN(n37445) );
  OR2_X1 U5907 ( .A1(n28205), .A2(n438), .Z(n27891) );
  NAND2_X1 U5908 ( .A1(n27940), .A2(n39193), .ZN(n20019) );
  NAND2_X1 U5912 ( .A1(n4502), .A2(n4503), .ZN(n4508) );
  NOR2_X1 U5914 ( .A1(n28101), .A2(n5266), .ZN(n39193) );
  NAND2_X1 U5917 ( .A1(n28180), .A2(n14389), .ZN(n4766) );
  INV_X1 U5918 ( .I(n36643), .ZN(n2467) );
  BUF_X1 U5922 ( .I(n17197), .Z(n34668) );
  CLKBUF_X2 U5924 ( .I(n4945), .Z(n39132) );
  AND2_X1 U5925 ( .A1(n7528), .A2(n28282), .Z(n37136) );
  CLKBUF_X2 U5930 ( .I(n18628), .Z(n39789) );
  CLKBUF_X4 U5934 ( .I(n27624), .Z(n28419) );
  BUF_X4 U5935 ( .I(n28182), .Z(n14397) );
  BUF_X1 U5936 ( .I(n3159), .Z(n38010) );
  BUF_X2 U5937 ( .I(n14411), .Z(n16325) );
  BUF_X4 U5945 ( .I(n27604), .Z(n28272) );
  AND2_X1 U5953 ( .A1(n2868), .A2(n28224), .Z(n37186) );
  CLKBUF_X2 U5956 ( .I(n18451), .Z(n39574) );
  INV_X1 U5957 ( .I(n13883), .ZN(n37540) );
  INV_X1 U5960 ( .I(n27723), .ZN(n37427) );
  BUF_X2 U5970 ( .I(n13703), .Z(n386) );
  CLKBUF_X2 U5971 ( .I(n27647), .Z(n18577) );
  BUF_X2 U5977 ( .I(n4127), .Z(n35350) );
  CLKBUF_X4 U5979 ( .I(n12551), .Z(n37101) );
  NAND2_X1 U5982 ( .A1(n35681), .A2(n39572), .ZN(n32245) );
  NAND2_X1 U5985 ( .A1(n20203), .A2(n27312), .ZN(n38635) );
  INV_X1 U5986 ( .I(n38152), .ZN(n38515) );
  INV_X1 U5989 ( .I(n37433), .ZN(n37432) );
  NAND2_X1 U6002 ( .A1(n6508), .A2(n6507), .ZN(n38587) );
  NAND2_X1 U6013 ( .A1(n26647), .A2(n38690), .ZN(n38688) );
  NAND2_X1 U6015 ( .A1(n35978), .A2(n38637), .ZN(n38636) );
  INV_X1 U6024 ( .I(n27354), .ZN(n39485) );
  INV_X1 U6029 ( .I(n39573), .ZN(n39572) );
  NAND2_X1 U6033 ( .A1(n27289), .A2(n37130), .ZN(n18769) );
  INV_X1 U6041 ( .I(n15641), .ZN(n38489) );
  NOR2_X1 U6063 ( .A1(n37771), .A2(n37770), .ZN(n8535) );
  OR2_X1 U6064 ( .A1(n5101), .A2(n27240), .Z(n37158) );
  NOR2_X1 U6067 ( .A1(n37385), .A2(n37384), .ZN(n35294) );
  OAI21_X1 U6069 ( .A1(n27096), .A2(n13992), .B(n27441), .ZN(n37903) );
  NAND2_X1 U6072 ( .A1(n38306), .A2(n38305), .ZN(n31926) );
  NOR2_X1 U6074 ( .A1(n4627), .A2(n6191), .ZN(n37655) );
  OAI21_X1 U6075 ( .A1(n19326), .A2(n27131), .B(n27338), .ZN(n39336) );
  OR2_X1 U6079 ( .A1(n18195), .A2(n38193), .Z(n9632) );
  NOR2_X1 U6081 ( .A1(n38983), .A2(n27253), .ZN(n27255) );
  INV_X2 U6089 ( .I(n27435), .ZN(n27149) );
  INV_X1 U6092 ( .I(n12766), .ZN(n37827) );
  INV_X2 U6096 ( .I(n27379), .ZN(n27298) );
  CLKBUF_X2 U6097 ( .I(n39484), .Z(n38571) );
  CLKBUF_X2 U6100 ( .I(n9144), .Z(n33503) );
  INV_X2 U6104 ( .I(n15284), .ZN(n27278) );
  AND2_X1 U6110 ( .A1(n6908), .A2(n21272), .Z(n37192) );
  CLKBUF_X4 U6119 ( .I(n36200), .Z(n34387) );
  CLKBUF_X2 U6125 ( .I(n35500), .Z(n39216) );
  CLKBUF_X4 U6132 ( .I(n27438), .Z(n7612) );
  INV_X1 U6139 ( .I(n16835), .ZN(n38983) );
  CLKBUF_X4 U6142 ( .I(n6533), .Z(n39414) );
  CLKBUF_X2 U6144 ( .I(n4886), .Z(n39628) );
  CLKBUF_X2 U6145 ( .I(n16736), .Z(n38578) );
  NAND2_X1 U6147 ( .A1(n38363), .A2(n38362), .ZN(n26446) );
  NOR2_X1 U6159 ( .A1(n12795), .A2(n37161), .ZN(n33098) );
  AND3_X1 U6167 ( .A1(n33849), .A2(n19179), .A3(n37098), .Z(n37161) );
  AOI21_X1 U6168 ( .A1(n26618), .A2(n34003), .B(n26621), .ZN(n9658) );
  NAND2_X1 U6170 ( .A1(n26785), .A2(n26862), .ZN(n4) );
  NAND2_X1 U6172 ( .A1(n1491), .A2(n8746), .ZN(n38362) );
  AND2_X1 U6174 ( .A1(n26847), .A2(n26945), .Z(n37133) );
  NAND2_X1 U6175 ( .A1(n26443), .A2(n33689), .ZN(n38363) );
  AND2_X1 U6176 ( .A1(n32344), .A2(n7619), .Z(n37131) );
  OR2_X1 U6177 ( .A1(n10187), .A2(n8478), .Z(n37188) );
  INV_X1 U6178 ( .I(n32072), .ZN(n37590) );
  INV_X4 U6181 ( .I(n10338), .ZN(n37102) );
  INV_X1 U6184 ( .I(n27013), .ZN(n39064) );
  NAND2_X1 U6187 ( .A1(n26769), .A2(n19442), .ZN(n16939) );
  NOR2_X1 U6188 ( .A1(n20666), .A2(n26990), .ZN(n19191) );
  OR2_X1 U6189 ( .A1(n16160), .A2(n20858), .Z(n34003) );
  CLKBUF_X2 U6190 ( .I(n26837), .Z(n38407) );
  OR2_X1 U6195 ( .A1(n26876), .A2(n21099), .Z(n37140) );
  CLKBUF_X2 U6197 ( .I(n34160), .Z(n38483) );
  BUF_X4 U6199 ( .I(n11617), .Z(n11616) );
  OR2_X1 U6200 ( .A1(n20171), .A2(n26770), .Z(n4808) );
  CLKBUF_X2 U6204 ( .I(n11948), .Z(n39564) );
  BUF_X4 U6205 ( .I(n26836), .Z(n37103) );
  CLKBUF_X4 U6208 ( .I(n26808), .Z(n19179) );
  INV_X1 U6209 ( .I(n31546), .ZN(n39602) );
  CLKBUF_X4 U6210 ( .I(n12788), .Z(n37104) );
  INV_X1 U6212 ( .I(n39611), .ZN(n26475) );
  CLKBUF_X2 U6216 ( .I(n26361), .Z(n38896) );
  BUF_X2 U6219 ( .I(n4875), .Z(n39637) );
  CLKBUF_X2 U6220 ( .I(n30913), .Z(n39093) );
  NAND2_X1 U6221 ( .A1(n37930), .A2(n35947), .ZN(n30967) );
  NOR2_X1 U6222 ( .A1(n37372), .A2(n18801), .ZN(n6478) );
  NAND2_X1 U6223 ( .A1(n14985), .A2(n38783), .ZN(n14984) );
  NAND2_X2 U6225 ( .A1(n9868), .A2(n25920), .ZN(n25596) );
  INV_X1 U6228 ( .I(n38930), .ZN(n34512) );
  AND2_X1 U6229 ( .A1(n7258), .A2(n11033), .Z(n37116) );
  INV_X1 U6230 ( .I(n30957), .ZN(n37310) );
  BUF_X1 U6232 ( .I(n1015), .Z(n37837) );
  INV_X2 U6233 ( .I(n5753), .ZN(n34577) );
  CLKBUF_X1 U6237 ( .I(n9412), .Z(n37819) );
  CLKBUF_X2 U6241 ( .I(n9694), .Z(n39375) );
  CLKBUF_X2 U6242 ( .I(n33879), .Z(n37502) );
  INV_X1 U6246 ( .I(n31367), .ZN(n37746) );
  BUF_X1 U6250 ( .I(n26108), .Z(n38501) );
  CLKBUF_X2 U6253 ( .I(n17696), .Z(n38507) );
  CLKBUF_X2 U6254 ( .I(n17180), .Z(n38760) );
  CLKBUF_X4 U6255 ( .I(n25899), .Z(n38825) );
  NAND2_X1 U6256 ( .A1(n1932), .A2(n1933), .ZN(n21204) );
  CLKBUF_X2 U6257 ( .I(n26093), .Z(n39729) );
  NAND2_X1 U6259 ( .A1(n37713), .A2(n37712), .ZN(n37711) );
  OAI21_X1 U6262 ( .A1(n19829), .A2(n10444), .B(n38013), .ZN(n38132) );
  NAND2_X1 U6268 ( .A1(n25645), .A2(n4467), .ZN(n37616) );
  OAI21_X1 U6270 ( .A1(n39252), .A2(n39251), .B(n5051), .ZN(n25635) );
  NAND2_X1 U6271 ( .A1(n9429), .A2(n15329), .ZN(n38301) );
  OR2_X1 U6272 ( .A1(n219), .A2(n32879), .Z(n38933) );
  INV_X1 U6273 ( .I(n38050), .ZN(n6173) );
  OR2_X1 U6275 ( .A1(n39328), .A2(n17029), .Z(n37182) );
  AND2_X1 U6277 ( .A1(n14436), .A2(n12533), .Z(n6472) );
  CLKBUF_X2 U6291 ( .I(n31895), .Z(n37748) );
  BUF_X2 U6296 ( .I(n32775), .Z(n38245) );
  NAND2_X1 U6299 ( .A1(n38863), .A2(n38862), .ZN(n38113) );
  CLKBUF_X4 U6304 ( .I(n10414), .Z(n39599) );
  CLKBUF_X2 U6311 ( .I(n11622), .Z(n38178) );
  CLKBUF_X2 U6328 ( .I(n19582), .Z(n39389) );
  CLKBUF_X4 U6332 ( .I(n25700), .Z(n12675) );
  BUF_X2 U6334 ( .I(n32165), .Z(n15172) );
  CLKBUF_X2 U6335 ( .I(n13873), .Z(n38661) );
  CLKBUF_X2 U6341 ( .I(n32433), .Z(n38560) );
  CLKBUF_X2 U6343 ( .I(n25186), .Z(n39146) );
  CLKBUF_X2 U6344 ( .I(n33132), .Z(n37312) );
  CLKBUF_X4 U6346 ( .I(n25269), .Z(n39765) );
  CLKBUF_X2 U6350 ( .I(n25118), .Z(n38665) );
  CLKBUF_X2 U6360 ( .I(n24999), .Z(n38950) );
  NAND2_X1 U6362 ( .A1(n17106), .A2(n9612), .ZN(n39496) );
  NAND2_X1 U6365 ( .A1(n11367), .A2(n38389), .ZN(n4427) );
  INV_X1 U6366 ( .I(n39256), .ZN(n39255) );
  NAND2_X1 U6377 ( .A1(n10793), .A2(n37193), .ZN(n24884) );
  BUF_X2 U6385 ( .I(n8605), .Z(n507) );
  NAND2_X1 U6387 ( .A1(n30700), .A2(n30698), .ZN(n37664) );
  NOR2_X1 U6388 ( .A1(n37233), .A2(n6357), .ZN(n30386) );
  OR2_X1 U6397 ( .A1(n24898), .A2(n38317), .Z(n31455) );
  INV_X1 U6405 ( .I(n24776), .ZN(n39540) );
  CLKBUF_X2 U6409 ( .I(n1118), .Z(n38631) );
  NOR2_X1 U6420 ( .A1(n1263), .A2(n16671), .ZN(n37688) );
  NAND2_X1 U6426 ( .A1(n38347), .A2(n24696), .ZN(n23857) );
  CLKBUF_X8 U6467 ( .I(n33996), .Z(n37477) );
  BUF_X4 U6475 ( .I(n39681), .Z(n31845) );
  CLKBUF_X2 U6476 ( .I(n7769), .Z(n37640) );
  BUF_X1 U6477 ( .I(n7770), .Z(n39513) );
  BUF_X4 U6481 ( .I(n17607), .Z(n37355) );
  CLKBUF_X8 U6482 ( .I(n32825), .Z(n37105) );
  BUF_X2 U6485 ( .I(n24779), .Z(n38658) );
  NAND2_X1 U6489 ( .A1(n37891), .A2(n18647), .ZN(n18608) );
  CLKBUF_X1 U6491 ( .I(n24753), .Z(n38884) );
  INV_X2 U6492 ( .I(n24650), .ZN(n36988) );
  NAND2_X1 U6493 ( .A1(n38652), .A2(n38250), .ZN(n37472) );
  NAND2_X1 U6497 ( .A1(n39660), .A2(n39659), .ZN(n18647) );
  NAND2_X1 U6500 ( .A1(n34938), .A2(n24069), .ZN(n39092) );
  NAND2_X1 U6515 ( .A1(n37710), .A2(n24170), .ZN(n38925) );
  NAND2_X1 U6516 ( .A1(n24305), .A2(n39796), .ZN(n8319) );
  NAND2_X1 U6517 ( .A1(n24253), .A2(n19782), .ZN(n39587) );
  NAND2_X1 U6518 ( .A1(n37959), .A2(n37958), .ZN(n5716) );
  NAND2_X1 U6520 ( .A1(n18759), .A2(n7000), .ZN(n6999) );
  INV_X1 U6524 ( .I(n16377), .ZN(n38473) );
  NOR2_X1 U6525 ( .A1(n6933), .A2(n24453), .ZN(n37392) );
  NAND2_X1 U6546 ( .A1(n4359), .A2(n24336), .ZN(n37635) );
  NAND2_X1 U6558 ( .A1(n9083), .A2(n9084), .ZN(n39738) );
  AND2_X1 U6561 ( .A1(n24396), .A2(n24169), .Z(n37187) );
  NAND2_X1 U6567 ( .A1(n38948), .A2(n11477), .ZN(n12176) );
  NAND2_X1 U6570 ( .A1(n16666), .A2(n24372), .ZN(n37959) );
  CLKBUF_X2 U6571 ( .I(n24381), .Z(n38812) );
  CLKBUF_X4 U6582 ( .I(n1129), .Z(n38431) );
  INV_X1 U6583 ( .I(n24470), .ZN(n38032) );
  INV_X2 U6585 ( .I(n13099), .ZN(n24169) );
  CLKBUF_X2 U6590 ( .I(n18830), .Z(n38487) );
  CLKBUF_X2 U6593 ( .I(n17871), .Z(n37733) );
  INV_X1 U6594 ( .I(n32899), .ZN(n38251) );
  BUF_X1 U6595 ( .I(n12235), .Z(n37994) );
  BUF_X4 U6596 ( .I(n37267), .Z(n39067) );
  CLKBUF_X2 U6618 ( .I(n11795), .Z(n37480) );
  BUF_X2 U6619 ( .I(n24106), .Z(n24396) );
  INV_X1 U6620 ( .I(n23565), .ZN(n37352) );
  BUF_X4 U6622 ( .I(n2297), .Z(n37107) );
  INV_X1 U6625 ( .I(n20384), .ZN(n35134) );
  INV_X1 U6634 ( .I(n7558), .ZN(n17288) );
  INV_X1 U6637 ( .I(n16833), .ZN(n5667) );
  CLKBUF_X2 U6645 ( .I(n39163), .Z(n37899) );
  CLKBUF_X2 U6646 ( .I(n3601), .Z(n39014) );
  NAND2_X1 U6651 ( .A1(n2960), .A2(n7389), .ZN(n39506) );
  INV_X1 U6653 ( .I(n12362), .ZN(n32562) );
  CLKBUF_X2 U6657 ( .I(n39038), .Z(n38370) );
  NAND2_X1 U6668 ( .A1(n32407), .A2(n32406), .ZN(n37705) );
  NAND2_X1 U6678 ( .A1(n30788), .A2(n37924), .ZN(n39218) );
  CLKBUF_X2 U6680 ( .I(n23619), .Z(n37431) );
  NAND2_X1 U6682 ( .A1(n4534), .A2(n37266), .ZN(n36966) );
  INV_X2 U6687 ( .I(n36859), .ZN(n38894) );
  NAND2_X1 U6689 ( .A1(n30524), .A2(n38726), .ZN(n23385) );
  BUF_X2 U6704 ( .I(n18204), .Z(n7387) );
  AND3_X1 U6710 ( .A1(n23477), .A2(n1139), .A3(n15176), .Z(n37135) );
  CLKBUF_X2 U6712 ( .I(n23355), .Z(n39534) );
  CLKBUF_X4 U6714 ( .I(n13217), .Z(n37523) );
  INV_X2 U6715 ( .I(n18199), .ZN(n23355) );
  BUF_X1 U6719 ( .I(n23310), .Z(n39626) );
  BUF_X1 U6721 ( .I(n23548), .Z(n38656) );
  CLKBUF_X2 U6725 ( .I(n1635), .Z(n37622) );
  INV_X2 U6729 ( .I(n32471), .ZN(n1304) );
  CLKBUF_X2 U6730 ( .I(n23423), .Z(n37814) );
  CLKBUF_X2 U6731 ( .I(n19671), .Z(n37463) );
  INV_X2 U6735 ( .I(n11342), .ZN(n31234) );
  CLKBUF_X2 U6736 ( .I(n30881), .Z(n38042) );
  NOR2_X1 U6738 ( .A1(n783), .A2(n37127), .ZN(n37500) );
  AOI22_X1 U6741 ( .A1(n17498), .A2(n23165), .B1(n17497), .B2(n23169), .ZN(
        n37901) );
  NOR2_X1 U6744 ( .A1(n37840), .A2(n14851), .ZN(n20910) );
  CLKBUF_X2 U6752 ( .I(n38653), .Z(n38100) );
  OAI21_X1 U6755 ( .A1(n23061), .A2(n23000), .B(n36167), .ZN(n38967) );
  NAND2_X1 U6762 ( .A1(n39297), .A2(n15032), .ZN(n35067) );
  OAI21_X1 U6765 ( .A1(n23082), .A2(n5515), .B(n38903), .ZN(n22910) );
  NOR2_X1 U6767 ( .A1(n7626), .A2(n12630), .ZN(n37518) );
  CLKBUF_X2 U6774 ( .I(n23173), .Z(n38752) );
  NAND3_X1 U6775 ( .A1(n23209), .A2(n23135), .A3(n19859), .ZN(n23134) );
  BUF_X2 U6783 ( .I(n19731), .Z(n121) );
  CLKBUF_X2 U6784 ( .I(n780), .Z(n38329) );
  BUF_X2 U6788 ( .I(n22864), .Z(n19288) );
  CLKBUF_X2 U6792 ( .I(n7584), .Z(n38542) );
  BUF_X2 U6795 ( .I(n34200), .Z(n5515) );
  CLKBUF_X2 U6803 ( .I(n1319), .Z(n39034) );
  CLKBUF_X2 U6806 ( .I(n23074), .Z(n31005) );
  CLKBUF_X4 U6807 ( .I(n7518), .Z(n6466) );
  BUF_X2 U6818 ( .I(n22879), .Z(n4682) );
  INV_X4 U6819 ( .I(n1046), .ZN(n37108) );
  BUF_X4 U6821 ( .I(n22942), .Z(n19586) );
  CLKBUF_X1 U6825 ( .I(n10382), .Z(n38216) );
  CLKBUF_X4 U6828 ( .I(n4624), .Z(n39787) );
  CLKBUF_X2 U6835 ( .I(n16798), .Z(n39548) );
  CLKBUF_X2 U6842 ( .I(n9982), .Z(n38330) );
  NAND2_X1 U6844 ( .A1(n22141), .A2(n20731), .ZN(n37708) );
  INV_X1 U6845 ( .I(n38522), .ZN(n10996) );
  NAND2_X1 U6849 ( .A1(n22319), .A2(n38917), .ZN(n12815) );
  OAI21_X1 U6853 ( .A1(n21963), .A2(n9987), .B(n38699), .ZN(n20042) );
  INV_X1 U6854 ( .I(n21972), .ZN(n17636) );
  INV_X1 U6862 ( .I(n37491), .ZN(n37490) );
  INV_X1 U6863 ( .I(n22282), .ZN(n38105) );
  CLKBUF_X2 U6864 ( .I(n11329), .Z(n37911) );
  AND3_X1 U6866 ( .A1(n32107), .A2(n22349), .A3(n22389), .Z(n2886) );
  CLKBUF_X2 U6870 ( .I(n22254), .Z(n39151) );
  NAND2_X1 U6871 ( .A1(n22205), .A2(n21288), .ZN(n38931) );
  BUF_X2 U6877 ( .I(n22362), .Z(n34246) );
  BUF_X2 U6882 ( .I(n22170), .Z(n554) );
  BUF_X2 U6889 ( .I(n6947), .Z(n6361) );
  CLKBUF_X2 U6891 ( .I(n38395), .Z(n38246) );
  NAND2_X1 U6892 ( .A1(n13239), .A2(n13240), .ZN(n39746) );
  INV_X1 U6897 ( .I(n37789), .ZN(n17436) );
  NAND2_X1 U6900 ( .A1(n13345), .A2(n17161), .ZN(n34683) );
  AOI22_X1 U6902 ( .A1(n21343), .A2(n21861), .B1(n21342), .B2(n36351), .ZN(
        n39771) );
  NAND2_X1 U6907 ( .A1(n21649), .A2(n1157), .ZN(n38547) );
  NAND2_X1 U6910 ( .A1(n20367), .A2(n21950), .ZN(n39658) );
  INV_X1 U6915 ( .I(n37399), .ZN(n37398) );
  NAND2_X1 U6917 ( .A1(n21695), .A2(n21876), .ZN(n39732) );
  BUF_X2 U6918 ( .I(n21905), .Z(n19647) );
  CLKBUF_X2 U6920 ( .I(n21593), .Z(n38480) );
  BUF_X2 U6926 ( .I(n12754), .Z(n35839) );
  NAND2_X1 U6927 ( .A1(n19650), .A2(n21876), .ZN(n21873) );
  CLKBUF_X4 U6929 ( .I(n21883), .Z(n19434) );
  INV_X1 U6935 ( .I(n30170), .ZN(n38261) );
  CLKBUF_X2 U6936 ( .I(n21628), .Z(n32412) );
  CLKBUF_X2 U6942 ( .I(n10656), .Z(n39656) );
  CLKBUF_X2 U6944 ( .I(n21641), .Z(n39650) );
  INV_X1 U6948 ( .I(n19919), .ZN(n38962) );
  INV_X1 U6949 ( .I(n29805), .ZN(n37261) );
  BUF_X2 U6962 ( .I(n15009), .Z(n37111) );
  INV_X1 U6965 ( .I(Plaintext[151]), .ZN(n38991) );
  INV_X1 U6966 ( .I(n4759), .ZN(n37659) );
  INV_X1 U6971 ( .I(n9759), .ZN(n38273) );
  NOR2_X1 U6972 ( .A1(n20003), .A2(n18028), .ZN(n16537) );
  INV_X1 U6974 ( .I(n21929), .ZN(n36721) );
  NAND2_X1 U6975 ( .A1(n21787), .A2(n18205), .ZN(n17966) );
  CLKBUF_X1 U6979 ( .I(n21669), .Z(n31222) );
  INV_X1 U6983 ( .I(n21582), .ZN(n19579) );
  NAND2_X1 U6985 ( .A1(n21274), .A2(n7536), .ZN(n38496) );
  CLKBUF_X1 U6988 ( .I(n32820), .Z(n39594) );
  CLKBUF_X2 U6991 ( .I(n33999), .Z(n39192) );
  NOR2_X1 U6993 ( .A1(n19403), .A2(n19554), .ZN(n19553) );
  NAND2_X1 U7000 ( .A1(n19084), .A2(n12754), .ZN(n2643) );
  AOI21_X1 U7004 ( .A1(n21820), .A2(n39594), .B(n1349), .ZN(n14734) );
  CLKBUF_X1 U7007 ( .I(n21721), .Z(n32704) );
  CLKBUF_X4 U7009 ( .I(n3839), .Z(n3562) );
  CLKBUF_X1 U7010 ( .I(n21644), .Z(n18112) );
  NOR2_X1 U7013 ( .A1(n21804), .A2(n36735), .ZN(n10127) );
  NAND2_X1 U7019 ( .A1(n21555), .A2(n10211), .ZN(n10144) );
  NAND2_X1 U7021 ( .A1(n21713), .A2(n19542), .ZN(n21531) );
  INV_X1 U7030 ( .I(n21854), .ZN(n21852) );
  NAND3_X1 U7036 ( .A1(n1156), .A2(n38241), .A3(n1345), .ZN(n7963) );
  NAND2_X1 U7040 ( .A1(n14928), .A2(n22315), .ZN(n19136) );
  INV_X1 U7044 ( .I(n37963), .ZN(n37962) );
  CLKBUF_X2 U7047 ( .I(n36728), .Z(n21783) );
  NAND2_X1 U7054 ( .A1(n30824), .A2(n3564), .ZN(n39785) );
  NAND2_X1 U7059 ( .A1(n6101), .A2(n21850), .ZN(n6098) );
  NAND2_X1 U7061 ( .A1(n5391), .A2(n5392), .ZN(n13438) );
  INV_X2 U7066 ( .I(n22229), .ZN(n1675) );
  INV_X1 U7067 ( .I(n22316), .ZN(n915) );
  CLKBUF_X4 U7073 ( .I(n21488), .Z(n21893) );
  BUF_X2 U7074 ( .I(n22292), .Z(n33571) );
  OAI21_X1 U7079 ( .A1(n22176), .A2(n4613), .B(n22335), .ZN(n21298) );
  OAI21_X1 U7083 ( .A1(n11091), .A2(n39075), .B(n1680), .ZN(n11142) );
  NAND2_X1 U7084 ( .A1(n22365), .A2(n7357), .ZN(n22007) );
  CLKBUF_X2 U7087 ( .I(n15350), .Z(n36227) );
  NOR2_X1 U7093 ( .A1(n37358), .A2(n33886), .ZN(n19777) );
  CLKBUF_X4 U7104 ( .I(n5929), .Z(n5075) );
  AOI21_X1 U7108 ( .A1(n133), .A2(n17897), .B(n7613), .ZN(n20254) );
  INV_X2 U7112 ( .I(n4613), .ZN(n22101) );
  NOR2_X1 U7117 ( .A1(n6347), .A2(n2257), .ZN(n2816) );
  AOI21_X1 U7128 ( .A1(n915), .A2(n22317), .B(n9824), .ZN(n12433) );
  NAND2_X1 U7131 ( .A1(n11171), .A2(n36397), .ZN(n19385) );
  NAND2_X1 U7134 ( .A1(n39151), .A2(n17723), .ZN(n12091) );
  OAI22_X1 U7137 ( .A1(n18429), .A2(n20623), .B1(n22365), .B2(n22366), .ZN(
        n11878) );
  NAND2_X1 U7138 ( .A1(n12365), .A2(n22324), .ZN(n37918) );
  NAND3_X1 U7141 ( .A1(n22061), .A2(n22178), .A3(n19261), .ZN(n16259) );
  INV_X1 U7143 ( .I(n22511), .ZN(n22695) );
  CLKBUF_X1 U7146 ( .I(n22621), .Z(n39654) );
  INV_X1 U7152 ( .I(n15871), .ZN(n22677) );
  INV_X1 U7153 ( .I(n15439), .ZN(n38920) );
  OAI21_X1 U7157 ( .A1(n16346), .A2(n16345), .B(n15439), .ZN(n6048) );
  NAND2_X1 U7161 ( .A1(n22255), .A2(n20308), .ZN(n17407) );
  INV_X1 U7162 ( .I(n7510), .ZN(n10384) );
  INV_X1 U7172 ( .I(n22689), .ZN(n3233) );
  INV_X1 U7180 ( .I(n22435), .ZN(n39047) );
  NAND2_X1 U7185 ( .A1(n33925), .A2(n14409), .ZN(n19724) );
  NAND2_X1 U7186 ( .A1(n10383), .A2(n15794), .ZN(n13719) );
  NAND3_X1 U7187 ( .A1(n20439), .A2(n17127), .A3(n1989), .ZN(n3289) );
  NAND2_X1 U7188 ( .A1(n14524), .A2(n5907), .ZN(n22799) );
  NAND2_X1 U7196 ( .A1(n20957), .A2(n23079), .ZN(n32358) );
  OAI22_X1 U7199 ( .A1(n15678), .A2(n781), .B1(n22895), .B2(n35918), .ZN(
        n14544) );
  NAND2_X1 U7201 ( .A1(n33935), .A2(n8197), .ZN(n7804) );
  NOR2_X1 U7205 ( .A1(n15455), .A2(n14089), .ZN(n22948) );
  INV_X2 U7208 ( .I(n19966), .ZN(n1648) );
  NOR2_X1 U7209 ( .A1(n8628), .A2(n16174), .ZN(n34522) );
  CLKBUF_X2 U7215 ( .I(n23080), .Z(n4846) );
  INV_X1 U7220 ( .I(n38282), .ZN(n22889) );
  CLKBUF_X2 U7226 ( .I(n23132), .Z(n17578) );
  INV_X1 U7230 ( .I(n33972), .ZN(n22931) );
  AOI21_X1 U7238 ( .A1(n17131), .A2(n17127), .B(n39810), .ZN(n18481) );
  CLKBUF_X1 U7244 ( .I(n23188), .Z(n39266) );
  INV_X2 U7245 ( .I(n22802), .ZN(n1645) );
  NAND2_X1 U7246 ( .A1(n22949), .A2(n37108), .ZN(n22722) );
  AOI21_X1 U7248 ( .A1(n23166), .A2(n22975), .B(n36554), .ZN(n22976) );
  NOR2_X1 U7250 ( .A1(n38019), .A2(n4773), .ZN(n37913) );
  INV_X2 U7252 ( .I(n14409), .ZN(n13946) );
  OAI21_X1 U7253 ( .A1(n22802), .A2(n32228), .B(n19134), .ZN(n9798) );
  NAND2_X1 U7254 ( .A1(n8676), .A2(n14804), .ZN(n33585) );
  NAND2_X1 U7263 ( .A1(n9797), .A2(n20518), .ZN(n14744) );
  AOI22_X1 U7271 ( .A1(n23044), .A2(n22368), .B1(n1989), .B2(n5806), .ZN(n5805) );
  AOI21_X1 U7274 ( .A1(n10378), .A2(n10377), .B(n8730), .ZN(n37840) );
  NAND2_X1 U7275 ( .A1(n22993), .A2(n22994), .ZN(n23067) );
  CLKBUF_X2 U7283 ( .I(n20077), .Z(n39418) );
  INV_X1 U7286 ( .I(n14561), .ZN(n23212) );
  INV_X1 U7290 ( .I(n37043), .ZN(n9543) );
  INV_X1 U7305 ( .I(n18481), .ZN(n37792) );
  OAI22_X1 U7306 ( .A1(n5658), .A2(n5657), .B1(n23197), .B2(n12245), .ZN(n327)
         );
  NAND2_X1 U7323 ( .A1(n1304), .A2(n20418), .ZN(n30789) );
  INV_X1 U7325 ( .I(n9823), .ZN(n18284) );
  INV_X1 U7327 ( .I(n23456), .ZN(n23293) );
  NAND3_X1 U7333 ( .A1(n1043), .A2(n1146), .A3(n31838), .ZN(n13078) );
  AOI21_X1 U7336 ( .A1(n936), .A2(n23020), .B(n1046), .ZN(n35939) );
  CLKBUF_X4 U7345 ( .I(n22005), .Z(n23111) );
  OAI21_X1 U7346 ( .A1(n38248), .A2(n1136), .B(n9321), .ZN(n38376) );
  NAND3_X1 U7350 ( .A1(n1632), .A2(n21247), .A3(n23602), .ZN(n23604) );
  INV_X2 U7352 ( .I(n10334), .ZN(n1144) );
  AOI21_X1 U7353 ( .A1(n23401), .A2(n16047), .B(n38353), .ZN(n12639) );
  OAI21_X1 U7355 ( .A1(n23358), .A2(n23250), .B(n33864), .ZN(n31055) );
  INV_X1 U7358 ( .I(n19005), .ZN(n21051) );
  INV_X1 U7359 ( .I(n37354), .ZN(n36635) );
  INV_X1 U7362 ( .I(n35001), .ZN(n38299) );
  NAND2_X1 U7366 ( .A1(n16047), .A2(n23400), .ZN(n37924) );
  AOI21_X1 U7372 ( .A1(n18939), .A2(n36564), .B(n30456), .ZN(n38373) );
  INV_X1 U7374 ( .I(n15353), .ZN(n5759) );
  NAND3_X1 U7375 ( .A1(n23370), .A2(n9823), .A3(n1140), .ZN(n4287) );
  NAND2_X1 U7380 ( .A1(n23493), .A2(n23315), .ZN(n22966) );
  NOR2_X1 U7381 ( .A1(n38535), .A2(n37463), .ZN(n20818) );
  NOR3_X1 U7382 ( .A1(n1290), .A2(n39194), .A3(n13414), .ZN(n9772) );
  OAI21_X1 U7389 ( .A1(n1304), .A2(n30499), .B(n12638), .ZN(n18917) );
  NAND2_X1 U7396 ( .A1(n19869), .A2(n18850), .ZN(n23009) );
  NAND2_X1 U7401 ( .A1(n20418), .A2(n36810), .ZN(n20776) );
  CLKBUF_X2 U7408 ( .I(n12966), .Z(n38881) );
  NAND2_X1 U7409 ( .A1(n4525), .A2(n38611), .ZN(n35302) );
  INV_X2 U7410 ( .I(n23749), .ZN(n10763) );
  INV_X1 U7419 ( .I(n23515), .ZN(n1293) );
  CLKBUF_X4 U7423 ( .I(n18681), .Z(n32858) );
  NOR2_X1 U7424 ( .A1(n16013), .A2(n23619), .ZN(n23455) );
  AOI21_X1 U7431 ( .A1(n37523), .A2(n23350), .B(n31906), .ZN(n38754) );
  AOI21_X1 U7432 ( .A1(n23321), .A2(n16299), .B(n23320), .ZN(n23322) );
  CLKBUF_X2 U7435 ( .I(n23967), .Z(n35561) );
  INV_X1 U7441 ( .I(n6559), .ZN(n36143) );
  NAND2_X1 U7447 ( .A1(n12597), .A2(n23303), .ZN(n32406) );
  INV_X1 U7449 ( .I(n4117), .ZN(n7833) );
  CLKBUF_X4 U7452 ( .I(n12362), .Z(n5116) );
  INV_X1 U7453 ( .I(n23943), .ZN(n30688) );
  INV_X1 U7454 ( .I(n23729), .ZN(n36068) );
  NOR2_X1 U7459 ( .A1(n9193), .A2(n39648), .ZN(n10589) );
  INV_X1 U7468 ( .I(n12799), .ZN(n11794) );
  NOR2_X1 U7469 ( .A1(n19656), .A2(n23976), .ZN(n2223) );
  CLKBUF_X2 U7471 ( .I(n24052), .Z(n39310) );
  NOR2_X1 U7475 ( .A1(n24235), .A2(n10477), .ZN(n32787) );
  NAND2_X1 U7478 ( .A1(n23819), .A2(n34561), .ZN(n36003) );
  NAND2_X1 U7480 ( .A1(n20404), .A2(n37230), .ZN(n34330) );
  NAND2_X1 U7481 ( .A1(n19857), .A2(n24271), .ZN(n38595) );
  INV_X1 U7485 ( .I(n1131), .ZN(n6465) );
  NAND2_X1 U7486 ( .A1(n4880), .A2(n21043), .ZN(n4286) );
  NAND2_X1 U7488 ( .A1(n39706), .A2(n94), .ZN(n7772) );
  NOR2_X1 U7493 ( .A1(n32899), .A2(n4880), .ZN(n37580) );
  INV_X1 U7497 ( .I(n39605), .ZN(n37849) );
  NAND2_X1 U7499 ( .A1(n24271), .A2(n11795), .ZN(n24272) );
  NAND2_X1 U7503 ( .A1(n38473), .A2(n1130), .ZN(n38472) );
  NAND2_X1 U7507 ( .A1(n2348), .A2(n11585), .ZN(n36561) );
  NOR2_X1 U7509 ( .A1(n24458), .A2(n38886), .ZN(n35854) );
  NOR2_X1 U7510 ( .A1(n24390), .A2(n9963), .ZN(n24187) );
  INV_X1 U7513 ( .I(n24164), .ZN(n24484) );
  AOI21_X1 U7514 ( .A1(n1128), .A2(n1130), .B(n38032), .ZN(n8360) );
  NOR2_X1 U7515 ( .A1(n24329), .A2(n24328), .ZN(n31443) );
  INV_X1 U7518 ( .I(n24467), .ZN(n1600) );
  NOR2_X1 U7527 ( .A1(n39067), .A2(n24461), .ZN(n20395) );
  NAND2_X1 U7529 ( .A1(n2395), .A2(n2393), .ZN(n2400) );
  NOR2_X1 U7530 ( .A1(n1275), .A2(n39699), .ZN(n34133) );
  OAI22_X1 U7532 ( .A1(n1601), .A2(n24309), .B1(n19745), .B2(n24445), .ZN(
        n24137) );
  OAI21_X1 U7535 ( .A1(n16590), .A2(n1594), .B(n24412), .ZN(n12425) );
  INV_X1 U7542 ( .I(n18830), .ZN(n24382) );
  INV_X1 U7545 ( .I(n12804), .ZN(n24399) );
  NAND2_X1 U7550 ( .A1(n24650), .A2(n37477), .ZN(n15850) );
  INV_X2 U7552 ( .I(n17693), .ZN(n1586) );
  NOR2_X1 U7554 ( .A1(n35952), .A2(n32093), .ZN(n34372) );
  NAND2_X1 U7555 ( .A1(n18721), .A2(n33104), .ZN(n17811) );
  OAI21_X1 U7557 ( .A1(n14617), .A2(n18551), .B(n24464), .ZN(n18550) );
  NAND2_X1 U7558 ( .A1(n10815), .A2(n37994), .ZN(n5138) );
  NAND2_X1 U7560 ( .A1(n19566), .A2(n205), .ZN(n24157) );
  NOR2_X1 U7565 ( .A1(n12665), .A2(n36154), .ZN(n34656) );
  NAND3_X1 U7566 ( .A1(n24442), .A2(n24443), .A3(n250), .ZN(n5066) );
  NOR2_X1 U7567 ( .A1(n3226), .A2(n24400), .ZN(n32484) );
  NAND2_X1 U7573 ( .A1(n4050), .A2(n2989), .ZN(n13228) );
  AOI22_X1 U7574 ( .A1(n14241), .A2(n36340), .B1(n24792), .B2(n19901), .ZN(
        n15849) );
  INV_X1 U7575 ( .I(n24674), .ZN(n13128) );
  NAND3_X1 U7579 ( .A1(n958), .A2(n24717), .A3(n24719), .ZN(n30507) );
  INV_X1 U7581 ( .I(n7529), .ZN(n24818) );
  NOR2_X1 U7582 ( .A1(n30554), .A2(n1577), .ZN(n30947) );
  CLKBUF_X2 U7586 ( .I(n19294), .Z(n36296) );
  AOI22_X1 U7587 ( .A1(n11053), .A2(n5431), .B1(n33012), .B2(n24826), .ZN(
        n38044) );
  NAND2_X1 U7590 ( .A1(n32882), .A2(n24746), .ZN(n13735) );
  NAND2_X1 U7591 ( .A1(n24789), .A2(n20039), .ZN(n8428) );
  NOR2_X1 U7595 ( .A1(n24897), .A2(n38317), .ZN(n38475) );
  INV_X1 U7598 ( .I(n21310), .ZN(n11169) );
  INV_X2 U7599 ( .I(n7769), .ZN(n38317) );
  BUF_X2 U7603 ( .I(n30464), .Z(n9921) );
  NOR3_X1 U7604 ( .A1(n1284), .A2(n24300), .A3(n8581), .ZN(n24185) );
  INV_X1 U7607 ( .I(n6066), .ZN(n5261) );
  INV_X1 U7609 ( .I(n7250), .ZN(n11319) );
  OAI21_X1 U7612 ( .A1(n24770), .A2(n8173), .B(n5495), .ZN(n5494) );
  NAND2_X1 U7613 ( .A1(n6491), .A2(n34526), .ZN(n31361) );
  INV_X1 U7626 ( .I(n25080), .ZN(n25124) );
  INV_X1 U7627 ( .I(n24545), .ZN(n24783) );
  OAI22_X1 U7628 ( .A1(n24798), .A2(n33409), .B1(n24800), .B2(n24799), .ZN(
        n3878) );
  NOR2_X1 U7630 ( .A1(n443), .A2(n36920), .ZN(n442) );
  AOI21_X1 U7635 ( .A1(n1122), .A2(n14857), .B(n14265), .ZN(n32400) );
  OAI21_X1 U7639 ( .A1(n37983), .A2(n16196), .B(n39279), .ZN(n7248) );
  INV_X1 U7640 ( .I(n24719), .ZN(n24721) );
  NAND2_X1 U7642 ( .A1(n1845), .A2(n933), .ZN(n1844) );
  INV_X1 U7643 ( .I(n24417), .ZN(n1559) );
  INV_X1 U7646 ( .I(n12233), .ZN(n32896) );
  CLKBUF_X2 U7648 ( .I(n24997), .Z(n38641) );
  INV_X1 U7650 ( .I(n25284), .ZN(n1556) );
  INV_X1 U7651 ( .I(n25272), .ZN(n39655) );
  OAI21_X1 U7652 ( .A1(n17100), .A2(n16540), .B(n16539), .ZN(n2530) );
  NAND2_X1 U7662 ( .A1(n24651), .A2(n24868), .ZN(n24652) );
  NAND2_X1 U7664 ( .A1(n21049), .A2(n24841), .ZN(n16746) );
  INV_X1 U7666 ( .I(n25210), .ZN(n4796) );
  INV_X1 U7669 ( .I(n25317), .ZN(n38430) );
  INV_X1 U7671 ( .I(n25196), .ZN(n38712) );
  INV_X1 U7674 ( .I(n32349), .ZN(n5433) );
  INV_X1 U7675 ( .I(n20304), .ZN(n35472) );
  INV_X1 U7680 ( .I(n36039), .ZN(n12251) );
  NAND2_X1 U7684 ( .A1(n25616), .A2(n18031), .ZN(n38625) );
  INV_X1 U7687 ( .I(n18810), .ZN(n38425) );
  NAND2_X1 U7692 ( .A1(n33268), .A2(n25361), .ZN(n149) );
  INV_X2 U7698 ( .I(n10055), .ZN(n38686) );
  NAND2_X1 U7699 ( .A1(n36991), .A2(n25513), .ZN(n38730) );
  NOR2_X1 U7700 ( .A1(n31359), .A2(n31358), .ZN(n831) );
  INV_X1 U7703 ( .I(n12944), .ZN(n12748) );
  OAI21_X1 U7706 ( .A1(n25527), .A2(n16933), .B(n19701), .ZN(n10788) );
  INV_X1 U7707 ( .I(n3451), .ZN(n32495) );
  NAND2_X1 U7708 ( .A1(n25365), .A2(n2576), .ZN(n20881) );
  NOR2_X1 U7716 ( .A1(n25328), .A2(n2803), .ZN(n19927) );
  NOR2_X1 U7717 ( .A1(n1252), .A2(n24963), .ZN(n39223) );
  AOI21_X1 U7732 ( .A1(n1531), .A2(n25692), .B(n8014), .ZN(n12779) );
  NAND2_X1 U7733 ( .A1(n36792), .A2(n16677), .ZN(n36475) );
  NOR2_X1 U7734 ( .A1(n1548), .A2(n32654), .ZN(n16739) );
  NOR2_X1 U7737 ( .A1(n178), .A2(n25670), .ZN(n12983) );
  CLKBUF_X4 U7742 ( .I(n15566), .Z(n39061) );
  INV_X2 U7743 ( .I(n826), .ZN(n21302) );
  NOR3_X1 U7748 ( .A1(n39061), .A2(n14413), .A3(n13129), .ZN(n18842) );
  AOI22_X1 U7751 ( .A1(n38732), .A2(n5042), .B1(n13461), .B2(n36486), .ZN(
        n15790) );
  CLKBUF_X2 U7754 ( .I(n36105), .Z(n34583) );
  OAI21_X1 U7756 ( .A1(n33130), .A2(n21042), .B(n39053), .ZN(n25497) );
  BUF_X2 U7758 ( .I(n25322), .Z(n25484) );
  INV_X1 U7760 ( .I(n13717), .ZN(n35015) );
  INV_X1 U7767 ( .I(n19644), .ZN(n12896) );
  OAI22_X1 U7772 ( .A1(n25603), .A2(n14708), .B1(n8739), .B2(n10814), .ZN(
        n35467) );
  NAND2_X1 U7773 ( .A1(n9336), .A2(n25644), .ZN(n9335) );
  AOI21_X1 U7775 ( .A1(n541), .A2(n16114), .B(n25517), .ZN(n16113) );
  NAND3_X1 U7777 ( .A1(n541), .A2(n11874), .A3(n1249), .ZN(n25621) );
  NAND2_X1 U7778 ( .A1(n16200), .A2(n26042), .ZN(n32468) );
  NOR2_X1 U7780 ( .A1(n926), .A2(n26055), .ZN(n13732) );
  AOI21_X1 U7781 ( .A1(n6844), .A2(n6845), .B(n1377), .ZN(n3219) );
  INV_X1 U7783 ( .I(n25915), .ZN(n5982) );
  NAND2_X1 U7784 ( .A1(n24535), .A2(n25647), .ZN(n33056) );
  AOI21_X1 U7786 ( .A1(n37336), .A2(n39160), .B(n911), .ZN(n38477) );
  INV_X1 U7788 ( .I(n35648), .ZN(n26103) );
  CLKBUF_X2 U7795 ( .I(n9743), .Z(n424) );
  INV_X2 U7797 ( .I(n12548), .ZN(n32690) );
  CLKBUF_X1 U7798 ( .I(n26086), .Z(n4772) );
  INV_X1 U7799 ( .I(n25870), .ZN(n25871) );
  NOR3_X1 U7800 ( .A1(n36906), .A2(n7767), .A3(n37393), .ZN(n30283) );
  OAI21_X1 U7802 ( .A1(n11624), .A2(n11552), .B(n18406), .ZN(n11623) );
  CLKBUF_X2 U7803 ( .I(n26092), .Z(n33237) );
  NAND2_X1 U7806 ( .A1(n4512), .A2(n4511), .ZN(n37821) );
  INV_X1 U7808 ( .I(n17455), .ZN(n16376) );
  INV_X1 U7812 ( .I(n11533), .ZN(n13391) );
  OAI21_X1 U7813 ( .A1(n34206), .A2(n2424), .B(n11858), .ZN(n17188) );
  NOR2_X1 U7814 ( .A1(n26331), .A2(n1240), .ZN(n24967) );
  NAND2_X1 U7816 ( .A1(n9294), .A2(n34743), .ZN(n34742) );
  OAI22_X1 U7817 ( .A1(n12002), .A2(n37072), .B1(n4191), .B2(n929), .ZN(n4189)
         );
  INV_X1 U7820 ( .I(n19648), .ZN(n39183) );
  INV_X2 U7823 ( .I(n37476), .ZN(n1506) );
  CLKBUF_X2 U7825 ( .I(n32106), .Z(n39793) );
  INV_X1 U7827 ( .I(n16294), .ZN(n37448) );
  CLKBUF_X2 U7829 ( .I(n26334), .Z(n38279) );
  CLKBUF_X4 U7841 ( .I(n6571), .Z(n39172) );
  CLKBUF_X2 U7844 ( .I(n26161), .Z(n38753) );
  INV_X1 U7846 ( .I(n26205), .ZN(n38028) );
  INV_X1 U7850 ( .I(n32386), .ZN(n7726) );
  CLKBUF_X2 U7853 ( .I(n34768), .Z(n39032) );
  NAND2_X1 U7857 ( .A1(n35967), .A2(n14355), .ZN(n3351) );
  NAND2_X1 U7860 ( .A1(n13110), .A2(n39825), .ZN(n3368) );
  INV_X1 U7862 ( .I(n19448), .ZN(n26830) );
  INV_X1 U7867 ( .I(n26385), .ZN(n34648) );
  NAND3_X1 U7869 ( .A1(n19972), .A2(n1234), .A3(n9117), .ZN(n26907) );
  INV_X1 U7871 ( .I(n26627), .ZN(n18226) );
  INV_X2 U7873 ( .I(n26830), .ZN(n1231) );
  INV_X1 U7876 ( .I(n26877), .ZN(n30724) );
  NAND2_X1 U7879 ( .A1(n14394), .A2(n1234), .ZN(n31220) );
  CLKBUF_X2 U7880 ( .I(n7742), .Z(n33279) );
  INV_X1 U7881 ( .I(n10187), .ZN(n38775) );
  AND3_X1 U7882 ( .A1(n10479), .A2(n37289), .A3(n11696), .Z(n37139) );
  INV_X2 U7886 ( .I(n26852), .ZN(n26614) );
  OAI21_X1 U7887 ( .A1(n26909), .A2(n26908), .B(n19972), .ZN(n26911) );
  NAND2_X1 U7890 ( .A1(n14079), .A2(n39564), .ZN(n15341) );
  NAND2_X1 U7894 ( .A1(n38776), .A2(n26709), .ZN(n9619) );
  BUF_X2 U7898 ( .I(n26832), .Z(n19225) );
  CLKBUF_X4 U7899 ( .I(n26839), .Z(n32345) );
  NAND2_X1 U7901 ( .A1(n30724), .A2(n30725), .ZN(n38778) );
  INV_X1 U7904 ( .I(n20704), .ZN(n26797) );
  CLKBUF_X4 U7906 ( .I(n18135), .Z(n13757) );
  AOI21_X1 U7907 ( .A1(n26840), .A2(n37103), .B(n32345), .ZN(n20754) );
  OAI21_X1 U7908 ( .A1(n948), .A2(n26696), .B(n1495), .ZN(n16708) );
  NOR2_X1 U7910 ( .A1(n37289), .A2(n11696), .ZN(n6312) );
  CLKBUF_X4 U7911 ( .I(n14383), .Z(n36344) );
  CLKBUF_X2 U7917 ( .I(n26935), .Z(n38120) );
  OAI21_X1 U7918 ( .A1(n26758), .A2(n12755), .B(n12767), .ZN(n12766) );
  NAND2_X1 U7924 ( .A1(n15411), .A2(n17158), .ZN(n11467) );
  NOR2_X1 U7927 ( .A1(n11696), .A2(n17515), .ZN(n13487) );
  INV_X1 U7930 ( .I(n35485), .ZN(n37654) );
  INV_X1 U7931 ( .I(n1492), .ZN(n21091) );
  INV_X1 U7938 ( .I(n4272), .ZN(n37653) );
  AND3_X1 U7939 ( .A1(n18054), .A2(n36344), .A3(n2158), .Z(n36583) );
  AND2_X1 U7940 ( .A1(n1092), .A2(n38002), .Z(n3962) );
  CLKBUF_X1 U7942 ( .I(n9618), .Z(n38577) );
  NAND3_X1 U7943 ( .A1(n14825), .A2(n16834), .A3(n6615), .ZN(n14824) );
  NAND2_X1 U7945 ( .A1(n26672), .A2(n3328), .ZN(n17260) );
  CLKBUF_X2 U7946 ( .I(n9188), .Z(n35282) );
  INV_X1 U7948 ( .I(n27363), .ZN(n1484) );
  OAI21_X1 U7956 ( .A1(n14521), .A2(n19505), .B(n26804), .ZN(n19504) );
  NAND2_X1 U7960 ( .A1(n27278), .A2(n9875), .ZN(n38306) );
  INV_X1 U7962 ( .I(n27131), .ZN(n19557) );
  INV_X1 U7968 ( .I(n32205), .ZN(n27053) );
  CLKBUF_X1 U7970 ( .I(n27213), .Z(n38926) );
  INV_X1 U7972 ( .I(n27392), .ZN(n13699) );
  NOR2_X1 U7973 ( .A1(n36989), .A2(n4034), .ZN(n27170) );
  NAND2_X1 U7978 ( .A1(n27150), .A2(n27149), .ZN(n32942) );
  NOR2_X1 U7979 ( .A1(n11162), .A2(n20057), .ZN(n9926) );
  NOR2_X1 U7989 ( .A1(n2035), .A2(n27402), .ZN(n11090) );
  NOR2_X1 U7992 ( .A1(n31875), .A2(n16170), .ZN(n37771) );
  NOR2_X1 U7993 ( .A1(n13278), .A2(n4272), .ZN(n27220) );
  INV_X1 U7997 ( .I(n20190), .ZN(n27015) );
  CLKBUF_X4 U7998 ( .I(n36177), .Z(n35990) );
  OR3_X1 U7999 ( .A1(n27337), .A2(n19326), .A3(n7096), .Z(n31735) );
  INV_X2 U8000 ( .I(n27320), .ZN(n27391) );
  NAND2_X1 U8001 ( .A1(n5027), .A2(n7096), .ZN(n35681) );
  NAND2_X1 U8007 ( .A1(n14261), .A2(n5675), .ZN(n33403) );
  OAI21_X1 U8008 ( .A1(n39532), .A2(n39531), .B(n6191), .ZN(n39730) );
  NOR2_X1 U8010 ( .A1(n2522), .A2(n1891), .ZN(n2304) );
  OAI21_X1 U8012 ( .A1(n11767), .A2(n36762), .B(n27449), .ZN(n8644) );
  NAND2_X1 U8013 ( .A1(n27232), .A2(n30671), .ZN(n18350) );
  OAI21_X1 U8014 ( .A1(n37801), .A2(n27092), .B(n16043), .ZN(n16045) );
  NAND2_X1 U8015 ( .A1(n32631), .A2(n7312), .ZN(n35158) );
  CLKBUF_X2 U8018 ( .I(n5588), .Z(n35485) );
  INV_X1 U8019 ( .I(n27304), .ZN(n27585) );
  BUF_X2 U8020 ( .I(n27404), .Z(n33803) );
  NAND3_X1 U8022 ( .A1(n34387), .A2(n31875), .A3(n4743), .ZN(n38637) );
  NAND2_X1 U8026 ( .A1(n27401), .A2(n33335), .ZN(n26845) );
  OAI21_X1 U8027 ( .A1(n38630), .A2(n27314), .B(n4434), .ZN(n4490) );
  INV_X2 U8028 ( .I(n6533), .ZN(n6534) );
  NOR2_X1 U8033 ( .A1(n13294), .A2(n39414), .ZN(n3921) );
  NOR2_X1 U8038 ( .A1(n27172), .A2(n19062), .ZN(n38144) );
  CLKBUF_X2 U8049 ( .I(n37881), .Z(n37499) );
  INV_X1 U8052 ( .I(n31778), .ZN(n27531) );
  CLKBUF_X4 U8054 ( .I(n11694), .Z(n282) );
  CLKBUF_X1 U8057 ( .I(n27810), .Z(n31320) );
  INV_X1 U8058 ( .I(n27725), .ZN(n37327) );
  INV_X1 U8061 ( .I(n27712), .ZN(n31137) );
  INV_X1 U8065 ( .I(n762), .ZN(n6365) );
  CLKBUF_X2 U8066 ( .I(n27498), .Z(n37639) );
  CLKBUF_X2 U8067 ( .I(n27566), .Z(n34902) );
  INV_X1 U8068 ( .I(n27547), .ZN(n11155) );
  INV_X1 U8069 ( .I(n35469), .ZN(n37418) );
  INV_X2 U8070 ( .I(n14426), .ZN(n1759) );
  INV_X1 U8082 ( .I(n27692), .ZN(n6642) );
  NOR2_X1 U8085 ( .A1(n20053), .A2(n15925), .ZN(n5940) );
  NAND2_X1 U8088 ( .A1(n11512), .A2(n17447), .ZN(n15364) );
  OR2_X1 U8090 ( .A1(n3771), .A2(n3770), .Z(n28234) );
  BUF_X2 U8094 ( .I(n20774), .Z(n39571) );
  INV_X2 U8095 ( .I(n14399), .ZN(n28273) );
  INV_X1 U8098 ( .I(n8078), .ZN(n28220) );
  INV_X1 U8099 ( .I(n1212), .ZN(n1450) );
  CLKBUF_X2 U8100 ( .I(n8080), .Z(n4649) );
  NAND2_X1 U8106 ( .A1(n288), .A2(n31571), .ZN(n37784) );
  INV_X1 U8108 ( .I(n36197), .ZN(n36954) );
  CLKBUF_X1 U8110 ( .I(n2980), .Z(n2262) );
  NOR2_X1 U8111 ( .A1(n28079), .A2(n7872), .ZN(n28080) );
  INV_X2 U8114 ( .I(n14480), .ZN(n16869) );
  CLKBUF_X2 U8116 ( .I(n9516), .Z(n156) );
  NOR2_X1 U8122 ( .A1(n36979), .A2(n14376), .ZN(n35146) );
  NAND2_X1 U8123 ( .A1(n16065), .A2(n28221), .ZN(n9702) );
  CLKBUF_X4 U8126 ( .I(n33958), .Z(n12260) );
  NAND2_X1 U8127 ( .A1(n6643), .A2(n16065), .ZN(n9024) );
  NOR2_X1 U8129 ( .A1(n28212), .A2(n12192), .ZN(n37642) );
  NOR3_X1 U8131 ( .A1(n6733), .A2(n28089), .A3(n8149), .ZN(n5160) );
  NAND2_X1 U8133 ( .A1(n2982), .A2(n2740), .ZN(n2981) );
  INV_X2 U8134 ( .I(n16363), .ZN(n17532) );
  NAND2_X1 U8136 ( .A1(n20663), .A2(n28269), .ZN(n20470) );
  INV_X1 U8138 ( .I(n28049), .ZN(n28139) );
  CLKBUF_X2 U8145 ( .I(n3158), .Z(n37451) );
  CLKBUF_X2 U8146 ( .I(n16500), .Z(n16154) );
  NOR2_X1 U8147 ( .A1(n28249), .A2(n3032), .ZN(n30366) );
  NOR2_X1 U8148 ( .A1(n35694), .A2(n16576), .ZN(n18379) );
  OAI21_X1 U8151 ( .A1(n28217), .A2(n987), .B(n16971), .ZN(n28083) );
  AOI21_X1 U8153 ( .A1(n1200), .A2(n12406), .B(n1074), .ZN(n27743) );
  OAI21_X1 U8157 ( .A1(n10756), .A2(n13059), .B(n33405), .ZN(n5864) );
  NAND2_X1 U8160 ( .A1(n15691), .A2(n15693), .ZN(n34480) );
  INV_X1 U8165 ( .I(n28753), .ZN(n31924) );
  NAND2_X1 U8170 ( .A1(n3598), .A2(n28575), .ZN(n2704) );
  NAND3_X1 U8171 ( .A1(n34516), .A2(n27983), .A3(n34515), .ZN(n38155) );
  NAND2_X1 U8172 ( .A1(n35357), .A2(n28807), .ZN(n8637) );
  NAND2_X1 U8174 ( .A1(n28546), .A2(n28729), .ZN(n9056) );
  CLKBUF_X1 U8175 ( .I(n28591), .Z(n35888) );
  AOI21_X1 U8177 ( .A1(n36788), .A2(n35173), .B(n28611), .ZN(n12891) );
  NOR2_X1 U8184 ( .A1(n32759), .A2(n1882), .ZN(n28708) );
  OAI21_X1 U8185 ( .A1(n19946), .A2(n34170), .B(n4724), .ZN(n28091) );
  INV_X2 U8192 ( .I(n28620), .ZN(n28339) );
  NOR2_X1 U8194 ( .A1(n1874), .A2(n30581), .ZN(n34305) );
  INV_X2 U8195 ( .I(n33765), .ZN(n19349) );
  NAND2_X1 U8200 ( .A1(n28758), .A2(n978), .ZN(n9017) );
  NOR2_X1 U8204 ( .A1(n12237), .A2(n5383), .ZN(n2333) );
  CLKBUF_X4 U8205 ( .I(n9597), .Z(n2022) );
  AND2_X1 U8207 ( .A1(n13727), .A2(n13726), .Z(n38172) );
  INV_X1 U8209 ( .I(n34651), .ZN(n31147) );
  NOR3_X1 U8210 ( .A1(n30953), .A2(n977), .A3(n28746), .ZN(n18626) );
  NOR2_X1 U8212 ( .A1(n28312), .A2(n5418), .ZN(n4969) );
  INV_X2 U8213 ( .I(n28496), .ZN(n7454) );
  INV_X1 U8214 ( .I(n28559), .ZN(n28655) );
  INV_X1 U8216 ( .I(n1184), .ZN(n34739) );
  OAI21_X1 U8218 ( .A1(n13237), .A2(n34915), .B(n28758), .ZN(n8449) );
  NAND2_X1 U8220 ( .A1(n38857), .A2(n38856), .ZN(n28565) );
  NAND2_X1 U8225 ( .A1(n13891), .A2(n17800), .ZN(n13893) );
  NAND2_X1 U8231 ( .A1(n28605), .A2(n8349), .ZN(n10758) );
  CLKBUF_X2 U8232 ( .I(n7429), .Z(n37956) );
  CLKBUF_X2 U8233 ( .I(n29057), .Z(n39631) );
  CLKBUF_X2 U8234 ( .I(n28971), .Z(n19405) );
  NAND2_X1 U8236 ( .A1(n35804), .A2(n35805), .ZN(n13965) );
  NOR3_X1 U8238 ( .A1(n39332), .A2(n13598), .A3(n31888), .ZN(n38608) );
  CLKBUF_X4 U8239 ( .I(n29144), .Z(n36905) );
  NAND2_X1 U8240 ( .A1(n1184), .A2(n9106), .ZN(n9109) );
  INV_X1 U8242 ( .I(n20465), .ZN(n38679) );
  CLKBUF_X2 U8243 ( .I(n15157), .Z(n15156) );
  INV_X1 U8248 ( .I(n29645), .ZN(n37304) );
  NOR2_X1 U8252 ( .A1(n29200), .A2(n15153), .ZN(n11885) );
  OAI21_X1 U8254 ( .A1(n30238), .A2(n9394), .B(n15651), .ZN(n33267) );
  NAND2_X1 U8255 ( .A1(n14449), .A2(n32906), .ZN(n29265) );
  NAND2_X1 U8257 ( .A1(n29459), .A2(n36275), .ZN(n36893) );
  INV_X1 U8258 ( .I(n19896), .ZN(n20429) );
  INV_X1 U8262 ( .I(n33368), .ZN(n18947) );
  CLKBUF_X2 U8264 ( .I(n14403), .Z(n8677) );
  INV_X2 U8265 ( .I(n14158), .ZN(n1183) );
  NAND2_X1 U8266 ( .A1(n1183), .A2(n14600), .ZN(n29861) );
  CLKBUF_X2 U8269 ( .I(n12940), .Z(n39585) );
  INV_X2 U8271 ( .I(n29059), .ZN(n39392) );
  NAND2_X1 U8276 ( .A1(n29452), .A2(n9993), .ZN(n28900) );
  INV_X2 U8279 ( .I(n37061), .ZN(n21269) );
  NOR2_X1 U8281 ( .A1(n19734), .A2(n29642), .ZN(n36102) );
  AOI21_X1 U8283 ( .A1(n28864), .A2(n14428), .B(n18947), .ZN(n9885) );
  CLKBUF_X4 U8285 ( .I(n17698), .Z(n1962) );
  NOR2_X1 U8288 ( .A1(n10610), .A2(n29815), .ZN(n39017) );
  INV_X1 U8289 ( .I(n16224), .ZN(n29938) );
  OAI21_X1 U8292 ( .A1(n16060), .A2(n8529), .B(n4255), .ZN(n37531) );
  NAND2_X1 U8295 ( .A1(n1181), .A2(n29185), .ZN(n14184) );
  CLKBUF_X2 U8297 ( .I(n29381), .Z(n12876) );
  NAND2_X1 U8301 ( .A1(n2792), .A2(n15189), .ZN(n7015) );
  INV_X2 U8302 ( .I(n4083), .ZN(n19476) );
  OAI21_X1 U8307 ( .A1(n28822), .A2(n30046), .B(n28825), .ZN(n11404) );
  NAND2_X1 U8309 ( .A1(n19162), .A2(n14892), .ZN(n30237) );
  NAND2_X1 U8310 ( .A1(n38163), .A2(n30128), .ZN(n11845) );
  CLKBUF_X1 U8311 ( .I(n29532), .Z(n39178) );
  NAND2_X1 U8312 ( .A1(n29437), .A2(n18502), .ZN(n29434) );
  NAND2_X1 U8313 ( .A1(n36101), .A2(n36100), .ZN(n19175) );
  INV_X1 U8321 ( .I(n29971), .ZN(n32129) );
  NOR2_X1 U8324 ( .A1(n11845), .A2(n17192), .ZN(n35625) );
  CLKBUF_X1 U8325 ( .I(n29535), .Z(n37605) );
  NOR2_X1 U8326 ( .A1(n19090), .A2(n16233), .ZN(n29275) );
  INV_X1 U8329 ( .I(n29410), .ZN(n29416) );
  OAI21_X1 U8335 ( .A1(n18793), .A2(n18794), .B(n33128), .ZN(n32452) );
  BUF_X2 U8338 ( .I(n18241), .Z(n3896) );
  CLKBUF_X1 U8343 ( .I(Key[140]), .Z(n29522) );
  INV_X1 U8345 ( .I(n29680), .ZN(n34239) );
  AOI22_X1 U8346 ( .A1(n13277), .A2(n29355), .B1(n29356), .B2(n13981), .ZN(
        n37262) );
  OAI21_X1 U8350 ( .A1(n32768), .A2(n32767), .B(n29362), .ZN(n37273) );
  INV_X1 U8355 ( .I(n29334), .ZN(n39482) );
  INV_X1 U8356 ( .I(n29442), .ZN(n1377) );
  AOI21_X1 U8361 ( .A1(n29790), .A2(n29791), .B(n37781), .ZN(n20939) );
  INV_X1 U8362 ( .I(n19674), .ZN(n1051) );
  OR2_X1 U8367 ( .A1(n14349), .A2(n11344), .Z(n37113) );
  NAND2_X1 U8370 ( .A1(n15573), .A2(n6067), .ZN(n37114) );
  AND2_X2 U8373 ( .A1(n24698), .A2(n24903), .Z(n37115) );
  OR2_X2 U8381 ( .A1(n11404), .A2(n35183), .Z(n37117) );
  AND2_X2 U8383 ( .A1(n6876), .A2(n35228), .Z(n37118) );
  AND2_X1 U8384 ( .A1(n5314), .A2(n16246), .Z(n37119) );
  AND3_X1 U8389 ( .A1(n28149), .A2(n37754), .A3(n1076), .Z(n37120) );
  XNOR2_X1 U8391 ( .A1(n15102), .A2(n19851), .ZN(n37121) );
  OR2_X1 U8393 ( .A1(n24169), .A2(n20457), .Z(n37122) );
  AND2_X1 U8396 ( .A1(n1408), .A2(n29780), .Z(n37123) );
  AND2_X2 U8397 ( .A1(n32472), .A2(n35705), .Z(n37125) );
  OR2_X1 U8399 ( .A1(n14560), .A2(n38229), .Z(n37127) );
  OR2_X2 U8400 ( .A1(n38636), .A2(n38635), .Z(n37129) );
  OR2_X1 U8409 ( .A1(n2761), .A2(n35299), .Z(n37130) );
  OR2_X1 U8411 ( .A1(n446), .A2(n14212), .Z(n37132) );
  OR2_X2 U8414 ( .A1(n2741), .A2(n37896), .Z(n37134) );
  AND2_X2 U8415 ( .A1(n31005), .A2(n33933), .Z(n37137) );
  OR2_X1 U8418 ( .A1(n22920), .A2(n9725), .Z(n37138) );
  AND2_X1 U8419 ( .A1(n22995), .A2(n19288), .Z(n37141) );
  AND2_X1 U8420 ( .A1(n27284), .A2(n30851), .Z(n37143) );
  AND2_X1 U8422 ( .A1(n38578), .A2(n27267), .Z(n37144) );
  AND3_X1 U8426 ( .A1(n15209), .A2(n1393), .A3(n29571), .Z(n37145) );
  AND2_X2 U8428 ( .A1(n29346), .A2(n29241), .Z(n37146) );
  XOR2_X1 U8430 ( .A1(n27851), .A2(n19940), .Z(n37147) );
  XNOR2_X1 U8432 ( .A1(n23933), .A2(n29432), .ZN(n37148) );
  XOR2_X1 U8436 ( .A1(n17310), .A2(n19763), .Z(n37149) );
  AND2_X1 U8437 ( .A1(n26329), .A2(n26092), .Z(n37150) );
  INV_X1 U8438 ( .I(n15466), .ZN(n21930) );
  OR2_X2 U8440 ( .A1(n38507), .A2(n32691), .Z(n37151) );
  AND2_X2 U8442 ( .A1(n19434), .A2(n19238), .Z(n37152) );
  OR2_X1 U8447 ( .A1(n26901), .A2(n34005), .Z(n37153) );
  AND2_X1 U8449 ( .A1(n21893), .A2(n21894), .Z(n37155) );
  AND2_X1 U8450 ( .A1(n8155), .A2(n18870), .Z(n37156) );
  NOR2_X1 U8452 ( .A1(n1445), .A2(n17755), .ZN(n37159) );
  AND2_X2 U8457 ( .A1(n39061), .A2(n20838), .Z(n37160) );
  AND2_X2 U8458 ( .A1(n9875), .A2(n15284), .Z(n37162) );
  AND2_X2 U8459 ( .A1(n22317), .A2(n22316), .Z(n37163) );
  NOR2_X1 U8461 ( .A1(n38202), .A2(n20056), .ZN(n37164) );
  CLKBUF_X2 U8465 ( .I(n19326), .Z(n5027) );
  INV_X1 U8468 ( .I(n10006), .ZN(n14428) );
  AND2_X1 U8472 ( .A1(n25566), .A2(n5166), .Z(n37165) );
  AND3_X1 U8474 ( .A1(n24310), .A2(n1289), .A3(n250), .Z(n37166) );
  AND2_X1 U8477 ( .A1(n23128), .A2(n5380), .Z(n37167) );
  OR3_X1 U8479 ( .A1(n34783), .A2(n24234), .A3(n30311), .Z(n37168) );
  AND2_X1 U8482 ( .A1(n5124), .A2(n5063), .Z(n37169) );
  AND2_X1 U8484 ( .A1(n39406), .A2(n35137), .Z(n37171) );
  NOR2_X1 U8491 ( .A1(n33949), .A2(n13286), .ZN(n37173) );
  AND3_X1 U8492 ( .A1(n1016), .A2(n26032), .A3(n3345), .Z(n37175) );
  OR2_X1 U8496 ( .A1(n21618), .A2(n1049), .Z(n37176) );
  AND2_X1 U8499 ( .A1(n16860), .A2(n39676), .Z(n37178) );
  AND2_X1 U8500 ( .A1(n3631), .A2(n18815), .Z(n37179) );
  OR2_X2 U8501 ( .A1(n32134), .A2(n37025), .Z(n37183) );
  OR2_X2 U8502 ( .A1(n25587), .A2(n4603), .Z(n37184) );
  AND2_X1 U8503 ( .A1(n18667), .A2(n777), .Z(n37185) );
  AND2_X1 U8506 ( .A1(n4542), .A2(n8692), .Z(n37190) );
  OR2_X1 U8508 ( .A1(n18114), .A2(n6337), .Z(n37193) );
  XNOR2_X1 U8509 ( .A1(n22492), .A2(n30101), .ZN(n37194) );
  XNOR2_X1 U8510 ( .A1(n27499), .A2(n28910), .ZN(n37195) );
  INV_X1 U8513 ( .I(n18757), .ZN(n19850) );
  CLKBUF_X2 U8514 ( .I(n18757), .Z(n16302) );
  INV_X1 U8519 ( .I(n19677), .ZN(n37443) );
  OR2_X1 U8520 ( .A1(n17931), .A2(n13029), .Z(n37196) );
  XNOR2_X1 U8526 ( .A1(n8312), .A2(n10558), .ZN(n37197) );
  OR2_X2 U8527 ( .A1(n27153), .A2(n27408), .Z(n37198) );
  CLKBUF_X2 U8530 ( .I(n21871), .Z(n19650) );
  INV_X1 U8532 ( .I(n21871), .ZN(n21756) );
  XOR2_X1 U8534 ( .A1(Plaintext[64]), .A2(Key[64]), .Z(n37200) );
  AND2_X2 U8535 ( .A1(n5089), .A2(n34644), .Z(n37201) );
  AND2_X1 U8536 ( .A1(n28726), .A2(n12237), .Z(n37203) );
  AND3_X2 U8538 ( .A1(n34516), .A2(n27983), .A3(n34515), .Z(n37204) );
  AND2_X1 U8540 ( .A1(n27397), .A2(n2522), .Z(n37205) );
  INV_X1 U8544 ( .I(n5126), .ZN(n30621) );
  INV_X2 U8547 ( .I(n12754), .ZN(n21942) );
  XNOR2_X1 U8555 ( .A1(n9151), .A2(n7018), .ZN(n37206) );
  NOR2_X1 U8560 ( .A1(n20346), .A2(n7644), .ZN(n37207) );
  AND2_X2 U8561 ( .A1(n23227), .A2(n23533), .Z(n37208) );
  AND2_X2 U8562 ( .A1(n12617), .A2(n19481), .Z(n37209) );
  OR2_X2 U8566 ( .A1(n30845), .A2(n7529), .Z(n37210) );
  INV_X2 U8567 ( .I(n31307), .ZN(n12943) );
  INV_X1 U8571 ( .I(n38948), .ZN(n15145) );
  AND3_X1 U8575 ( .A1(n19740), .A2(n37819), .A3(n37613), .Z(n37211) );
  OR2_X2 U8579 ( .A1(n10980), .A2(n16502), .Z(n37212) );
  CLKBUF_X1 U8586 ( .I(n10980), .Z(n36395) );
  INV_X1 U8590 ( .I(n27820), .ZN(n37855) );
  XNOR2_X1 U8591 ( .A1(n22584), .A2(n5235), .ZN(n37214) );
  NOR2_X1 U8592 ( .A1(n3510), .A2(n32956), .ZN(n39714) );
  NAND2_X1 U8593 ( .A1(n39714), .A2(n24912), .ZN(n37215) );
  AND2_X2 U8595 ( .A1(n17074), .A2(n10632), .Z(n37216) );
  OR2_X2 U8597 ( .A1(n21370), .A2(n21369), .Z(n37217) );
  INV_X1 U8608 ( .I(n23201), .ZN(n19524) );
  INV_X1 U8609 ( .I(n34200), .ZN(n7266) );
  XOR2_X1 U8618 ( .A1(n5835), .A2(n35286), .Z(n37218) );
  OR2_X1 U8622 ( .A1(n23192), .A2(n1147), .Z(n37219) );
  OR2_X1 U8625 ( .A1(n9835), .A2(n23475), .Z(n37220) );
  XOR2_X1 U8626 ( .A1(n23952), .A2(n30122), .Z(n37221) );
  XNOR2_X1 U8630 ( .A1(n32239), .A2(n16320), .ZN(n37222) );
  XNOR2_X1 U8634 ( .A1(n11372), .A2(n39183), .ZN(n37223) );
  XNOR2_X1 U8643 ( .A1(n23888), .A2(n23808), .ZN(n37224) );
  AND2_X1 U8646 ( .A1(n1290), .A2(n39194), .Z(n37225) );
  AND2_X1 U8647 ( .A1(n22295), .A2(n16880), .Z(n37226) );
  XNOR2_X1 U8651 ( .A1(n6156), .A2(n30451), .ZN(n37227) );
  NAND2_X1 U8652 ( .A1(n37016), .A2(n37411), .ZN(n37228) );
  INV_X1 U8657 ( .I(n25574), .ZN(n1113) );
  AND2_X2 U8660 ( .A1(n24369), .A2(n24192), .Z(n37229) );
  XNOR2_X1 U8665 ( .A1(n7920), .A2(n31869), .ZN(n37230) );
  XNOR2_X1 U8673 ( .A1(n4302), .A2(n36171), .ZN(n37231) );
  XOR2_X1 U8674 ( .A1(n37816), .A2(n39044), .Z(n37232) );
  INV_X1 U8675 ( .I(n39681), .ZN(n19565) );
  INV_X2 U8677 ( .I(n31722), .ZN(n16990) );
  OR2_X1 U8678 ( .A1(n3760), .A2(n30464), .Z(n37233) );
  XOR2_X1 U8679 ( .A1(n11321), .A2(n19919), .Z(n37234) );
  INV_X2 U8680 ( .I(n5634), .ZN(n37983) );
  CLKBUF_X1 U8681 ( .I(n36798), .Z(n39048) );
  CLKBUF_X2 U8689 ( .I(n21301), .Z(n15541) );
  INV_X1 U8694 ( .I(n21301), .ZN(n37553) );
  INV_X2 U8699 ( .I(n840), .ZN(n19889) );
  XNOR2_X1 U8702 ( .A1(n5118), .A2(n6877), .ZN(n37235) );
  XOR2_X1 U8703 ( .A1(n34469), .A2(n29371), .Z(n37236) );
  OR2_X2 U8713 ( .A1(n33949), .A2(n25322), .Z(n37237) );
  OR2_X2 U8714 ( .A1(n14045), .A2(n730), .Z(n37238) );
  AND2_X2 U8730 ( .A1(n11003), .A2(n840), .Z(n37239) );
  INV_X1 U8731 ( .I(n17237), .ZN(n36391) );
  CLKBUF_X4 U8742 ( .I(n17237), .Z(n38238) );
  XNOR2_X1 U8747 ( .A1(n21044), .A2(n27634), .ZN(n37240) );
  INV_X2 U8797 ( .I(n1235), .ZN(n11513) );
  AND2_X2 U8800 ( .A1(n8988), .A2(n8798), .Z(n37241) );
  XNOR2_X1 U8801 ( .A1(n27499), .A2(n27178), .ZN(n37242) );
  XNOR2_X1 U8805 ( .A1(n27681), .A2(n27680), .ZN(n37243) );
  OR2_X1 U8807 ( .A1(n33491), .A2(n35260), .Z(n37244) );
  OR2_X2 U8809 ( .A1(n9658), .A2(n32563), .Z(n37245) );
  XNOR2_X1 U8810 ( .A1(n20713), .A2(n6133), .ZN(n37247) );
  OR3_X1 U8814 ( .A1(n28683), .A2(n1414), .A3(n1196), .Z(n37248) );
  AND2_X1 U8821 ( .A1(n28698), .A2(n28695), .Z(n37249) );
  CLKBUF_X4 U8822 ( .I(n26906), .Z(n1234) );
  INV_X1 U8823 ( .I(n13891), .ZN(n6703) );
  INV_X1 U8825 ( .I(n11375), .ZN(n14152) );
  INV_X1 U8833 ( .I(n14411), .ZN(n13492) );
  NOR2_X1 U8837 ( .A1(n10461), .A2(n35427), .ZN(n37250) );
  AND2_X2 U8843 ( .A1(n20056), .A2(n15047), .Z(n37251) );
  XNOR2_X1 U8845 ( .A1(n15745), .A2(n1710), .ZN(n37252) );
  INV_X1 U8848 ( .I(n29247), .ZN(n4905) );
  OR2_X1 U8850 ( .A1(n31595), .A2(n30057), .Z(n37253) );
  XNOR2_X1 U8851 ( .A1(n29095), .A2(n19683), .ZN(n37254) );
  AND2_X1 U8852 ( .A1(n36935), .A2(n31554), .Z(n37255) );
  AND2_X2 U8861 ( .A1(n11491), .A2(n11492), .Z(n37256) );
  INV_X1 U8866 ( .I(n10422), .ZN(n14449) );
  AND2_X1 U8869 ( .A1(n3159), .A2(n32932), .Z(n37257) );
  INV_X1 U8870 ( .I(n30221), .ZN(n30158) );
  AND2_X1 U8871 ( .A1(n29627), .A2(n29626), .Z(n37258) );
  XOR2_X1 U8885 ( .A1(n13248), .A2(n13246), .Z(n37259) );
  NOR3_X2 U8887 ( .A1(n38542), .A2(n8491), .A3(n35684), .ZN(n33737) );
  XOR2_X1 U8889 ( .A1(n31775), .A2(n29282), .Z(n34586) );
  NAND2_X2 U8891 ( .A1(n35885), .A2(n3795), .ZN(n31775) );
  XOR2_X1 U8894 ( .A1(n15532), .A2(n37260), .Z(n33701) );
  XOR2_X1 U8895 ( .A1(n23973), .A2(n37261), .Z(n37260) );
  NAND2_X2 U8896 ( .A1(n3076), .A2(n31861), .ZN(n31637) );
  XOR2_X1 U8901 ( .A1(n37262), .A2(n1717), .Z(Ciphertext[30]) );
  XOR2_X1 U8902 ( .A1(n4622), .A2(n37112), .Z(n34165) );
  NAND2_X2 U8905 ( .A1(n25377), .A2(n36900), .ZN(n4622) );
  XOR2_X1 U8906 ( .A1(n23700), .A2(n13074), .Z(n13871) );
  XNOR2_X1 U8908 ( .A1(n23832), .A2(n23938), .ZN(n23700) );
  NAND2_X1 U8909 ( .A1(n10404), .A2(n34685), .ZN(n25370) );
  NAND2_X2 U8912 ( .A1(n16767), .A2(n36897), .ZN(n34685) );
  INV_X2 U8914 ( .I(n11145), .ZN(n25513) );
  NAND2_X2 U8923 ( .A1(n37346), .A2(n32942), .ZN(n34838) );
  OAI22_X2 U8927 ( .A1(n32255), .A2(n8221), .B1(n8223), .B2(n20648), .ZN(
        n37378) );
  XOR2_X1 U8931 ( .A1(n22619), .A2(n22759), .Z(n8068) );
  XOR2_X1 U8932 ( .A1(n5171), .A2(n22371), .Z(n22759) );
  CLKBUF_X4 U8934 ( .I(n15218), .Z(n37589) );
  NAND2_X2 U8938 ( .A1(n29845), .A2(n37263), .ZN(n2346) );
  NAND3_X2 U8939 ( .A1(n29908), .A2(n29954), .A3(n29863), .ZN(n37263) );
  XOR2_X1 U8941 ( .A1(n30856), .A2(n8729), .Z(n28970) );
  AOI21_X2 U8943 ( .A1(n15829), .A2(n19690), .B(n24219), .ZN(n24565) );
  XNOR2_X1 U8950 ( .A1(n9930), .A2(n28982), .ZN(n29066) );
  NAND2_X2 U8951 ( .A1(n4196), .A2(n4197), .ZN(n28982) );
  NAND2_X1 U8958 ( .A1(n4745), .A2(n4746), .ZN(n33036) );
  BUF_X4 U8963 ( .I(n19857), .Z(n37264) );
  NAND2_X1 U8966 ( .A1(n12065), .A2(n37604), .ZN(n18469) );
  XOR2_X1 U8967 ( .A1(n15442), .A2(n37053), .Z(n11927) );
  INV_X2 U8969 ( .I(n36743), .ZN(n37053) );
  XOR2_X1 U8973 ( .A1(n18012), .A2(n13155), .Z(n36743) );
  NOR2_X2 U8975 ( .A1(n38911), .A2(n2886), .ZN(n37031) );
  NAND2_X2 U8980 ( .A1(n37265), .A2(n39179), .ZN(n7542) );
  NOR2_X2 U8982 ( .A1(n36307), .A2(n36306), .ZN(n37265) );
  XOR2_X1 U8983 ( .A1(n37381), .A2(n10592), .Z(n36435) );
  NAND2_X2 U8984 ( .A1(n27233), .A2(n12306), .ZN(n27434) );
  NAND2_X2 U8990 ( .A1(n35321), .A2(n3136), .ZN(n27233) );
  NAND2_X2 U8993 ( .A1(n1294), .A2(n2182), .ZN(n37266) );
  NAND2_X2 U8994 ( .A1(n7034), .A2(n7033), .ZN(n24746) );
  INV_X2 U8997 ( .I(n14353), .ZN(n14668) );
  NAND2_X2 U9000 ( .A1(n17926), .A2(n14354), .ZN(n14353) );
  INV_X2 U9001 ( .I(n31673), .ZN(n37267) );
  XOR2_X1 U9002 ( .A1(n37268), .A2(n12014), .Z(n35796) );
  XOR2_X1 U9007 ( .A1(n30653), .A2(n31073), .Z(n37268) );
  XOR2_X1 U9008 ( .A1(n10792), .A2(n25303), .Z(n25102) );
  OAI22_X2 U9009 ( .A1(n24128), .A2(n18114), .B1(n24127), .B2(n6337), .ZN(
        n10792) );
  NAND2_X2 U9014 ( .A1(n910), .A2(n11034), .ZN(n2865) );
  OAI22_X2 U9015 ( .A1(n7513), .A2(n11548), .B1(n25365), .B2(n36345), .ZN(
        n11034) );
  OAI21_X1 U9016 ( .A1(n1140), .A2(n18090), .B(n23299), .ZN(n31052) );
  NAND2_X2 U9020 ( .A1(n27357), .A2(n35198), .ZN(n27066) );
  NAND2_X2 U9021 ( .A1(n6376), .A2(n5560), .ZN(n27357) );
  XOR2_X1 U9025 ( .A1(n12296), .A2(n37269), .Z(n35645) );
  XOR2_X1 U9026 ( .A1(n25083), .A2(n37498), .Z(n37269) );
  XOR2_X1 U9028 ( .A1(n22549), .A2(n22647), .Z(n22736) );
  NAND2_X2 U9030 ( .A1(n22105), .A2(n22104), .ZN(n22647) );
  NAND2_X1 U9032 ( .A1(n38079), .A2(n19061), .ZN(n4463) );
  NAND2_X2 U9033 ( .A1(n37270), .A2(n5625), .ZN(n5623) );
  NAND2_X2 U9034 ( .A1(n31702), .A2(n5361), .ZN(n32354) );
  OR2_X1 U9037 ( .A1(n7317), .A2(n35138), .Z(n2940) );
  NAND3_X1 U9045 ( .A1(n25999), .A2(n2940), .A3(n19121), .ZN(n38342) );
  AOI22_X2 U9060 ( .A1(n1604), .A2(n37271), .B1(n37480), .B2(n33289), .ZN(
        n15829) );
  NAND2_X1 U9061 ( .A1(n35954), .A2(n12950), .ZN(n37271) );
  XOR2_X1 U9064 ( .A1(n22475), .A2(n9873), .Z(n7942) );
  AOI21_X2 U9071 ( .A1(n5878), .A2(n5877), .B(n5874), .ZN(n22475) );
  INV_X2 U9073 ( .I(n28163), .ZN(n2877) );
  XOR2_X1 U9075 ( .A1(n11730), .A2(n27748), .Z(n31880) );
  OAI22_X1 U9084 ( .A1(n961), .A2(n20418), .B1(n32471), .B2(n23399), .ZN(
        n22873) );
  OAI21_X2 U9085 ( .A1(n18413), .A2(n37272), .B(n1056), .ZN(n33476) );
  NOR2_X1 U9087 ( .A1(n29998), .A2(n30041), .ZN(n37272) );
  XOR2_X1 U9091 ( .A1(n37273), .A2(n29363), .Z(Ciphertext[33]) );
  AOI21_X2 U9093 ( .A1(n4075), .A2(n34652), .B(n37274), .ZN(n4073) );
  AND2_X1 U9096 ( .A1(n14089), .A2(n17210), .Z(n17459) );
  NOR2_X2 U9097 ( .A1(n37275), .A2(n3624), .ZN(n24813) );
  XOR2_X1 U9098 ( .A1(n21096), .A2(n34809), .Z(n19458) );
  XOR2_X1 U9100 ( .A1(n37280), .A2(n13568), .Z(n36822) );
  XOR2_X1 U9106 ( .A1(n8865), .A2(n557), .Z(n37280) );
  OAI21_X1 U9108 ( .A1(n27951), .A2(n20739), .B(n12303), .ZN(n37895) );
  XOR2_X1 U9109 ( .A1(n36522), .A2(n19933), .Z(n12935) );
  NAND2_X2 U9112 ( .A1(n8234), .A2(n8235), .ZN(n36522) );
  XOR2_X1 U9115 ( .A1(n27668), .A2(n18548), .Z(n18547) );
  XOR2_X1 U9118 ( .A1(n4934), .A2(n27802), .Z(n27668) );
  INV_X2 U9119 ( .I(n26026), .ZN(n26525) );
  OR2_X1 U9120 ( .A1(n28661), .A2(n28660), .Z(n34176) );
  XOR2_X1 U9123 ( .A1(n26514), .A2(n10965), .Z(n26375) );
  NOR2_X2 U9126 ( .A1(n14722), .A2(n21307), .ZN(n26514) );
  NAND2_X2 U9130 ( .A1(n9916), .A2(n25936), .ZN(n25812) );
  NAND3_X2 U9131 ( .A1(n10936), .A2(n10935), .A3(n10313), .ZN(n9916) );
  NAND2_X2 U9132 ( .A1(n33546), .A2(n15667), .ZN(n27508) );
  NOR2_X2 U9133 ( .A1(n37281), .A2(n36801), .ZN(n37522) );
  AOI21_X2 U9134 ( .A1(n24227), .A2(n18573), .B(n4601), .ZN(n10648) );
  NAND2_X2 U9136 ( .A1(n1029), .A2(n2634), .ZN(n24227) );
  NAND2_X2 U9141 ( .A1(n19438), .A2(n25567), .ZN(n5356) );
  NAND2_X1 U9147 ( .A1(n5354), .A2(n25724), .ZN(n19438) );
  XOR2_X1 U9149 ( .A1(n37593), .A2(n11105), .Z(n2068) );
  NAND2_X2 U9152 ( .A1(n10269), .A2(n10270), .ZN(n37593) );
  XOR2_X1 U9155 ( .A1(n37282), .A2(n33758), .Z(n39326) );
  XOR2_X1 U9158 ( .A1(n37855), .A2(n3114), .Z(n37282) );
  AOI22_X2 U9161 ( .A1(n37915), .A2(n37914), .B1(n38319), .B2(n30237), .ZN(
        n38204) );
  NAND2_X2 U9164 ( .A1(n34853), .A2(n27306), .ZN(n26790) );
  XOR2_X1 U9165 ( .A1(n34237), .A2(n26485), .Z(n38968) );
  NAND3_X2 U9166 ( .A1(n36458), .A2(n38632), .A3(n38633), .ZN(n26485) );
  XOR2_X1 U9168 ( .A1(n27655), .A2(n27654), .Z(n11358) );
  XOR2_X1 U9169 ( .A1(n27637), .A2(n27729), .Z(n27655) );
  NAND2_X2 U9170 ( .A1(n38766), .A2(n37283), .ZN(n28400) );
  AOI22_X2 U9171 ( .A1(n10084), .A2(n38666), .B1(n1202), .B2(n12038), .ZN(
        n37283) );
  XOR2_X1 U9173 ( .A1(n29147), .A2(n6758), .Z(n29258) );
  NAND2_X2 U9179 ( .A1(n28304), .A2(n28305), .ZN(n6758) );
  XOR2_X1 U9181 ( .A1(n27668), .A2(n7416), .Z(n7864) );
  XOR2_X1 U9183 ( .A1(n27504), .A2(n27492), .Z(n7416) );
  NOR3_X2 U9194 ( .A1(n33395), .A2(n586), .A3(n26053), .ZN(n34310) );
  XNOR2_X1 U9196 ( .A1(n25087), .A2(n14643), .ZN(n38109) );
  OAI22_X2 U9201 ( .A1(n37284), .A2(n33963), .B1(n10568), .B2(n20251), .ZN(
        n20274) );
  NOR2_X2 U9202 ( .A1(n14539), .A2(n18007), .ZN(n37284) );
  NOR3_X1 U9205 ( .A1(n26018), .A2(n2349), .A3(n26054), .ZN(n2621) );
  NAND2_X2 U9206 ( .A1(n9788), .A2(n37711), .ZN(n26018) );
  NAND4_X2 U9207 ( .A1(n9806), .A2(n12452), .A3(n30401), .A4(n31495), .ZN(
        n38067) );
  NAND2_X1 U9209 ( .A1(n35381), .A2(n6191), .ZN(n35380) );
  NOR2_X1 U9210 ( .A1(n38051), .A2(n19151), .ZN(n29499) );
  XOR2_X1 U9212 ( .A1(n15091), .A2(n15090), .Z(n17425) );
  XOR2_X1 U9214 ( .A1(n26536), .A2(n26539), .Z(n8021) );
  XOR2_X1 U9215 ( .A1(n5241), .A2(n26163), .Z(n26539) );
  OR2_X1 U9218 ( .A1(n27218), .A2(n15616), .Z(n13231) );
  NAND2_X1 U9220 ( .A1(n28724), .A2(n28360), .ZN(n37285) );
  XOR2_X1 U9222 ( .A1(n26160), .A2(n26484), .Z(n13426) );
  XOR2_X1 U9223 ( .A1(n38514), .A2(n26448), .Z(n26160) );
  NAND2_X1 U9225 ( .A1(n32861), .A2(n37002), .ZN(n38482) );
  NOR2_X2 U9228 ( .A1(n37287), .A2(n37286), .ZN(n31769) );
  INV_X2 U9234 ( .I(n26893), .ZN(n37289) );
  XOR2_X1 U9236 ( .A1(n27612), .A2(n27469), .Z(n37668) );
  XOR2_X1 U9242 ( .A1(n37833), .A2(n5900), .Z(n27612) );
  OAI22_X2 U9245 ( .A1(n26700), .A2(n19951), .B1(n36244), .B2(n10440), .ZN(
        n26178) );
  XOR2_X1 U9246 ( .A1(n37290), .A2(n7734), .Z(n9133) );
  XOR2_X1 U9248 ( .A1(n23716), .A2(n23725), .Z(n37290) );
  AOI21_X2 U9249 ( .A1(n5906), .A2(n1440), .B(n37291), .ZN(n6426) );
  OAI22_X1 U9250 ( .A1(n5905), .A2(n8522), .B1(n18696), .B2(n5266), .ZN(n37291) );
  NOR2_X1 U9251 ( .A1(n920), .A2(n37632), .ZN(n11567) );
  AOI22_X2 U9257 ( .A1(n38237), .A2(n38236), .B1(n12657), .B2(n18043), .ZN(
        n37632) );
  NAND3_X2 U9259 ( .A1(n38093), .A2(n27203), .A3(n37292), .ZN(n27792) );
  NAND3_X1 U9264 ( .A1(n16946), .A2(n27201), .A3(n14881), .ZN(n37292) );
  NOR2_X2 U9265 ( .A1(n39291), .A2(n25921), .ZN(n34339) );
  NAND2_X2 U9268 ( .A1(n5908), .A2(n26215), .ZN(n25921) );
  NOR2_X2 U9274 ( .A1(n14469), .A2(n37293), .ZN(n7424) );
  OAI22_X2 U9276 ( .A1(n26858), .A2(n8103), .B1(n11651), .B2(n11652), .ZN(
        n37293) );
  INV_X4 U9277 ( .I(n23381), .ZN(n33864) );
  OAI22_X2 U9280 ( .A1(n4099), .A2(n4100), .B1(n4102), .B2(n23057), .ZN(n23381) );
  XOR2_X1 U9281 ( .A1(n22538), .A2(n37294), .Z(n37459) );
  XOR2_X1 U9285 ( .A1(n22534), .A2(n22533), .Z(n37294) );
  BUF_X2 U9291 ( .I(n28772), .Z(n37295) );
  XOR2_X1 U9294 ( .A1(n4077), .A2(n26417), .Z(n3161) );
  NAND2_X2 U9297 ( .A1(n7317), .A2(n35138), .ZN(n26000) );
  OR2_X2 U9303 ( .A1(n5929), .A2(n8882), .Z(n8089) );
  NAND3_X2 U9307 ( .A1(n38481), .A2(n38482), .A3(n26789), .ZN(n27542) );
  OAI21_X2 U9308 ( .A1(n6585), .A2(n24175), .B(n24228), .ZN(n37601) );
  XOR2_X1 U9310 ( .A1(n9122), .A2(n23882), .Z(n9121) );
  XOR2_X1 U9311 ( .A1(n37932), .A2(n23890), .Z(n23882) );
  INV_X2 U9316 ( .I(n2030), .ZN(n38282) );
  XOR2_X1 U9318 ( .A1(n37296), .A2(n25323), .Z(n25174) );
  NOR2_X2 U9320 ( .A1(n17474), .A2(n17473), .ZN(n25323) );
  INV_X2 U9323 ( .I(n24857), .ZN(n37296) );
  XOR2_X1 U9325 ( .A1(n37297), .A2(n18359), .Z(n32128) );
  XOR2_X1 U9326 ( .A1(n22627), .A2(n22628), .Z(n37297) );
  OAI22_X2 U9331 ( .A1(n33359), .A2(n17989), .B1(n4200), .B2(n17499), .ZN(
        n4199) );
  NAND2_X1 U9333 ( .A1(n38063), .A2(n29626), .ZN(n37298) );
  NAND3_X2 U9335 ( .A1(n28326), .A2(n30389), .A3(n28325), .ZN(n3927) );
  NAND2_X2 U9339 ( .A1(n36860), .A2(n7872), .ZN(n30389) );
  XOR2_X1 U9340 ( .A1(n26527), .A2(n37299), .Z(n2754) );
  XOR2_X1 U9343 ( .A1(n1506), .A2(n26587), .Z(n37299) );
  NOR2_X2 U9344 ( .A1(n1244), .A2(n26055), .ZN(n26053) );
  OAI21_X2 U9346 ( .A1(n1320), .A2(n8491), .B(n22935), .ZN(n13542) );
  INV_X2 U9348 ( .I(n31558), .ZN(n8491) );
  XOR2_X1 U9349 ( .A1(n628), .A2(n31559), .Z(n31558) );
  NAND2_X2 U9359 ( .A1(n15763), .A2(n21091), .ZN(n4579) );
  OAI22_X2 U9361 ( .A1(n12065), .A2(n7305), .B1(n2140), .B2(n33952), .ZN(
        n15763) );
  NAND2_X2 U9362 ( .A1(n21067), .A2(n21066), .ZN(n23885) );
  NAND2_X2 U9363 ( .A1(n23520), .A2(n10024), .ZN(n21067) );
  XOR2_X1 U9364 ( .A1(n8021), .A2(n8020), .Z(n19298) );
  XOR2_X1 U9366 ( .A1(n9861), .A2(n19751), .Z(n33924) );
  OAI22_X2 U9369 ( .A1(n24254), .A2(n34055), .B1(n34141), .B2(n21049), .ZN(
        n9861) );
  XOR2_X1 U9370 ( .A1(n9548), .A2(n9549), .Z(n9383) );
  NAND3_X2 U9371 ( .A1(n35145), .A2(n2495), .A3(n2496), .ZN(n692) );
  NAND2_X2 U9373 ( .A1(n20458), .A2(n15258), .ZN(n37732) );
  NAND2_X1 U9380 ( .A1(n4001), .A2(n1545), .ZN(n4468) );
  XOR2_X1 U9385 ( .A1(n37301), .A2(n38712), .Z(n38711) );
  XOR2_X1 U9388 ( .A1(n37357), .A2(n25083), .Z(n37301) );
  XOR2_X1 U9390 ( .A1(n16743), .A2(n31767), .Z(n34365) );
  NAND2_X2 U9391 ( .A1(n36467), .A2(n8485), .ZN(n16743) );
  NAND3_X2 U9393 ( .A1(n946), .A2(n26695), .A3(n10338), .ZN(n142) );
  NAND2_X2 U9397 ( .A1(n37550), .A2(n5533), .ZN(n5024) );
  NAND2_X1 U9398 ( .A1(n22323), .A2(n22322), .ZN(n37302) );
  OAI22_X2 U9400 ( .A1(n28618), .A2(n30858), .B1(n2500), .B2(n28655), .ZN(
        n29137) );
  NOR2_X2 U9401 ( .A1(n2678), .A2(n11034), .ZN(n25925) );
  NAND2_X2 U9405 ( .A1(n6965), .A2(n32615), .ZN(n2678) );
  NAND2_X2 U9407 ( .A1(n37305), .A2(n3722), .ZN(n34603) );
  NAND3_X2 U9408 ( .A1(n36251), .A2(n5309), .A3(n1653), .ZN(n37305) );
  BUF_X2 U9410 ( .I(n37730), .Z(n37306) );
  XOR2_X1 U9412 ( .A1(n27631), .A2(n37307), .Z(n31778) );
  XOR2_X1 U9413 ( .A1(n10582), .A2(n25201), .Z(n10583) );
  INV_X2 U9414 ( .I(n30279), .ZN(n19466) );
  NOR2_X2 U9415 ( .A1(n13201), .A2(n13200), .ZN(n25133) );
  OR2_X1 U9418 ( .A1(n37308), .A2(n23461), .Z(n3174) );
  OAI21_X2 U9419 ( .A1(n37310), .A2(n37309), .B(n12711), .ZN(n39521) );
  INV_X2 U9420 ( .I(n28680), .ZN(n37311) );
  XOR2_X1 U9422 ( .A1(n27677), .A2(n8874), .Z(n8873) );
  XOR2_X1 U9424 ( .A1(n8875), .A2(n39442), .Z(n8874) );
  XOR2_X1 U9426 ( .A1(n37313), .A2(n17646), .Z(Ciphertext[168]) );
  AOI22_X1 U9432 ( .A1(n30135), .A2(n30144), .B1(n30134), .B2(n30133), .ZN(
        n37313) );
  NOR2_X2 U9434 ( .A1(n19657), .A2(n37251), .ZN(n27686) );
  XOR2_X1 U9439 ( .A1(n37314), .A2(n23921), .Z(n32472) );
  XOR2_X1 U9440 ( .A1(n5441), .A2(n5442), .Z(n37314) );
  OAI21_X2 U9442 ( .A1(n2464), .A2(n21148), .B(n37315), .ZN(n19279) );
  OAI21_X2 U9449 ( .A1(n5572), .A2(n33077), .B(n37316), .ZN(n37315) );
  NOR2_X2 U9450 ( .A1(n32507), .A2(n37125), .ZN(n37316) );
  XOR2_X1 U9452 ( .A1(n2618), .A2(n37317), .Z(n30982) );
  XOR2_X1 U9453 ( .A1(n34149), .A2(n25314), .Z(n37317) );
  NAND2_X2 U9454 ( .A1(n26608), .A2(n21317), .ZN(n27449) );
  XOR2_X1 U9455 ( .A1(n14312), .A2(n11215), .Z(n5322) );
  XOR2_X1 U9457 ( .A1(n4956), .A2(n23832), .Z(n14312) );
  NAND2_X2 U9458 ( .A1(n27263), .A2(n36969), .ZN(n27265) );
  XOR2_X1 U9459 ( .A1(n12196), .A2(n34250), .Z(n15412) );
  OAI22_X2 U9460 ( .A1(n37732), .A2(n21124), .B1(n37229), .B2(n20083), .ZN(
        n24650) );
  AOI22_X2 U9461 ( .A1(n9071), .A2(n9073), .B1(n18845), .B2(n355), .ZN(n37498)
         );
  INV_X1 U9462 ( .I(n28719), .ZN(n37561) );
  NOR2_X2 U9463 ( .A1(n29413), .A2(n29409), .ZN(n20724) );
  AOI22_X2 U9468 ( .A1(n29379), .A2(n6314), .B1(n17295), .B2(n16876), .ZN(
        n29413) );
  INV_X2 U9470 ( .I(n4322), .ZN(n31192) );
  NAND2_X2 U9472 ( .A1(n25384), .A2(n12996), .ZN(n4322) );
  NOR3_X2 U9475 ( .A1(n31483), .A2(n37318), .A3(n32504), .ZN(n37989) );
  INV_X1 U9479 ( .I(n38941), .ZN(n29600) );
  OAI21_X2 U9489 ( .A1(n5035), .A2(n35663), .B(n3923), .ZN(n35998) );
  AOI22_X2 U9499 ( .A1(n39448), .A2(n37598), .B1(n19719), .B2(n36203), .ZN(
        n35663) );
  AOI22_X2 U9505 ( .A1(n2462), .A2(n2461), .B1(n25437), .B2(n25562), .ZN(n8096) );
  OAI22_X2 U9506 ( .A1(n6505), .A2(n28376), .B1(n32012), .B2(n28448), .ZN(
        n32866) );
  NOR2_X2 U9509 ( .A1(n3899), .A2(n39020), .ZN(n28376) );
  NOR2_X2 U9510 ( .A1(n36583), .A2(n36582), .ZN(n998) );
  AND2_X1 U9511 ( .A1(n6892), .A2(n12527), .Z(n28336) );
  XNOR2_X1 U9514 ( .A1(n25272), .A2(n2064), .ZN(n37324) );
  BUF_X4 U9516 ( .I(n18967), .Z(n34000) );
  NAND3_X2 U9523 ( .A1(n37321), .A2(n4543), .A3(n37320), .ZN(n24034) );
  NAND2_X2 U9525 ( .A1(n13603), .A2(n33080), .ZN(n37321) );
  NOR2_X2 U9532 ( .A1(n39303), .A2(n37108), .ZN(n22950) );
  XOR2_X1 U9534 ( .A1(n2065), .A2(n37324), .Z(n37662) );
  XOR2_X1 U9536 ( .A1(n37325), .A2(n287), .Z(n1961) );
  XOR2_X1 U9538 ( .A1(n38133), .A2(n33715), .Z(n37325) );
  XOR2_X1 U9539 ( .A1(n37326), .A2(n14031), .Z(n38470) );
  XOR2_X1 U9540 ( .A1(n37427), .A2(n37327), .Z(n37326) );
  OAI21_X2 U9541 ( .A1(n13536), .A2(n13538), .B(n13535), .ZN(n37393) );
  XOR2_X1 U9545 ( .A1(n15686), .A2(n37328), .Z(n16186) );
  XOR2_X1 U9546 ( .A1(n25208), .A2(n17595), .Z(n37328) );
  NAND3_X2 U9547 ( .A1(n37330), .A2(n14232), .A3(n37329), .ZN(n39382) );
  INV_X2 U9548 ( .I(n28272), .ZN(n37329) );
  NAND2_X2 U9550 ( .A1(n1759), .A2(n11628), .ZN(n37330) );
  NAND2_X2 U9551 ( .A1(n11252), .A2(n11251), .ZN(n6904) );
  INV_X2 U9553 ( .I(n37331), .ZN(n38084) );
  NAND2_X2 U9566 ( .A1(n13780), .A2(n11613), .ZN(n37331) );
  INV_X1 U9573 ( .I(n3441), .ZN(n39501) );
  NOR2_X2 U9575 ( .A1(n11560), .A2(n37332), .ZN(n6559) );
  OAI22_X2 U9588 ( .A1(n23338), .A2(n21293), .B1(n12870), .B2(n23474), .ZN(
        n37332) );
  OAI21_X2 U9592 ( .A1(n13206), .A2(n5569), .B(n37333), .ZN(n17508) );
  NAND2_X2 U9597 ( .A1(n15743), .A2(n32590), .ZN(n37333) );
  XOR2_X1 U9599 ( .A1(n23786), .A2(n23785), .Z(n6092) );
  NAND2_X2 U9601 ( .A1(n26003), .A2(n38507), .ZN(n25854) );
  NAND2_X2 U9603 ( .A1(n37334), .A2(n34762), .ZN(n3903) );
  BUF_X2 U9605 ( .I(n22849), .Z(n37335) );
  AOI21_X2 U9607 ( .A1(n13690), .A2(n10883), .B(n1429), .ZN(n9692) );
  INV_X4 U9611 ( .I(n27624), .ZN(n35694) );
  BUF_X2 U9612 ( .I(n39061), .Z(n37336) );
  NOR2_X2 U9614 ( .A1(n38755), .A2(n38939), .ZN(n38211) );
  XOR2_X1 U9615 ( .A1(n23965), .A2(n11383), .Z(n1971) );
  NAND2_X2 U9621 ( .A1(n2950), .A2(n23345), .ZN(n23965) );
  NOR2_X1 U9624 ( .A1(n39696), .A2(n18144), .ZN(n38906) );
  XOR2_X1 U9625 ( .A1(n37337), .A2(n7729), .Z(n27903) );
  XOR2_X1 U9626 ( .A1(n37540), .A2(n1859), .Z(n37337) );
  NAND3_X2 U9627 ( .A1(n17754), .A2(n27147), .A3(n27434), .ZN(n37346) );
  OR2_X1 U9628 ( .A1(n24699), .A2(n24698), .Z(n35735) );
  NAND2_X2 U9637 ( .A1(n24712), .A2(n24903), .ZN(n24699) );
  NAND2_X2 U9640 ( .A1(n10907), .A2(n28686), .ZN(n18035) );
  NAND2_X2 U9641 ( .A1(n35496), .A2(n12349), .ZN(n10907) );
  NOR2_X2 U9645 ( .A1(n12925), .A2(n22899), .ZN(n22902) );
  INV_X4 U9646 ( .I(n39127), .ZN(n13491) );
  INV_X2 U9649 ( .I(n17727), .ZN(n1659) );
  NAND2_X2 U9652 ( .A1(n9391), .A2(n9392), .ZN(n17727) );
  NOR2_X2 U9653 ( .A1(n11676), .A2(n27910), .ZN(n12038) );
  NAND2_X2 U9662 ( .A1(n37669), .A2(n25608), .ZN(n19258) );
  AOI22_X2 U9667 ( .A1(n25872), .A2(n32520), .B1(n25871), .B2(n17501), .ZN(
        n37742) );
  XOR2_X1 U9668 ( .A1(n26340), .A2(n26227), .Z(n12014) );
  NOR2_X2 U9671 ( .A1(n12709), .A2(n12708), .ZN(n26340) );
  BUF_X2 U9672 ( .I(n39442), .Z(n37338) );
  NAND3_X2 U9674 ( .A1(n37339), .A2(n5902), .A3(n5901), .ZN(n17696) );
  XOR2_X1 U9676 ( .A1(n20044), .A2(n19343), .Z(n31673) );
  XOR2_X1 U9679 ( .A1(n12299), .A2(n33120), .Z(n15988) );
  XOR2_X1 U9681 ( .A1(n12805), .A2(n37340), .Z(n33934) );
  XOR2_X1 U9682 ( .A1(n39047), .A2(n22436), .Z(n37340) );
  XOR2_X1 U9686 ( .A1(n25204), .A2(n39582), .Z(n38736) );
  BUF_X2 U9689 ( .I(n10054), .Z(n37341) );
  XOR2_X1 U9694 ( .A1(n27526), .A2(n27813), .Z(n3474) );
  XOR2_X1 U9695 ( .A1(n13802), .A2(n27617), .Z(n27526) );
  NAND2_X2 U9697 ( .A1(n38604), .A2(n4997), .ZN(n14234) );
  XOR2_X1 U9699 ( .A1(n31293), .A2(n26279), .Z(n10668) );
  NAND2_X2 U9702 ( .A1(n38122), .A2(n34499), .ZN(n26279) );
  INV_X2 U9709 ( .I(n37342), .ZN(n3873) );
  XNOR2_X1 U9711 ( .A1(n3732), .A2(n38706), .ZN(n37342) );
  NAND2_X2 U9713 ( .A1(n37343), .A2(n22952), .ZN(n10480) );
  OAI21_X2 U9715 ( .A1(n22948), .A2(n17459), .B(n23138), .ZN(n37343) );
  XOR2_X1 U9716 ( .A1(n38639), .A2(n37344), .Z(n18732) );
  XOR2_X1 U9718 ( .A1(n10562), .A2(n8723), .Z(n37344) );
  INV_X2 U9720 ( .I(n34969), .ZN(n27411) );
  NAND3_X2 U9722 ( .A1(n7362), .A2(n25428), .A3(n20358), .ZN(n11148) );
  XOR2_X1 U9723 ( .A1(n37345), .A2(n26403), .Z(n26410) );
  XOR2_X1 U9724 ( .A1(n26405), .A2(n26402), .Z(n37345) );
  NAND2_X2 U9725 ( .A1(n10480), .A2(n8668), .ZN(n23620) );
  OR2_X1 U9727 ( .A1(n23572), .A2(n12154), .Z(n32362) );
  OAI21_X2 U9728 ( .A1(n28129), .A2(n31942), .B(n10287), .ZN(n28464) );
  XOR2_X1 U9734 ( .A1(n22720), .A2(n17612), .Z(n37382) );
  XOR2_X1 U9735 ( .A1(n16226), .A2(n39528), .Z(n17612) );
  XOR2_X1 U9739 ( .A1(n37347), .A2(n11072), .Z(n3827) );
  XOR2_X1 U9742 ( .A1(n14454), .A2(n23985), .Z(n35601) );
  OAI21_X2 U9743 ( .A1(n24182), .A2(n19739), .B(n1587), .ZN(n12279) );
  NOR2_X1 U9749 ( .A1(n12138), .A2(n35164), .ZN(n19739) );
  INV_X2 U9753 ( .I(n29377), .ZN(n31521) );
  NAND2_X2 U9754 ( .A1(n3697), .A2(n35952), .ZN(n38801) );
  NAND2_X2 U9756 ( .A1(n33529), .A2(n4184), .ZN(n3697) );
  INV_X1 U9759 ( .I(n39788), .ZN(n7224) );
  AND2_X1 U9761 ( .A1(n39788), .A2(n13414), .Z(n39803) );
  NAND2_X1 U9764 ( .A1(n29611), .A2(n32980), .ZN(n20126) );
  NOR2_X1 U9767 ( .A1(n25564), .A2(n25563), .ZN(n37584) );
  NAND2_X2 U9773 ( .A1(n12363), .A2(n12364), .ZN(n33132) );
  XOR2_X1 U9774 ( .A1(n26242), .A2(n26243), .Z(n37347) );
  OAI22_X2 U9775 ( .A1(n4433), .A2(n35887), .B1(n299), .B2(n4013), .ZN(n38416)
         );
  AOI22_X2 U9778 ( .A1(n19495), .A2(n1254), .B1(n9815), .B2(n33491), .ZN(n4013) );
  AOI22_X2 U9779 ( .A1(n37244), .A2(n37348), .B1(n25597), .B2(n20515), .ZN(
        n20381) );
  NOR2_X2 U9780 ( .A1(n37350), .A2(n5503), .ZN(n37559) );
  AOI21_X2 U9781 ( .A1(n13437), .A2(n6604), .B(n5392), .ZN(n37350) );
  NOR3_X2 U9782 ( .A1(n31607), .A2(n36844), .A3(n28246), .ZN(n15087) );
  OAI21_X2 U9783 ( .A1(n4152), .A2(n4153), .B(n28102), .ZN(n20020) );
  OAI22_X2 U9794 ( .A1(n36574), .A2(n36575), .B1(n15183), .B2(n3356), .ZN(
        n32253) );
  XOR2_X1 U9796 ( .A1(n19024), .A2(n6177), .Z(n17486) );
  AOI22_X2 U9798 ( .A1(n32109), .A2(n13731), .B1(n34524), .B2(n25424), .ZN(
        n4660) );
  XOR2_X1 U9801 ( .A1(n25239), .A2(n19064), .Z(n20365) );
  XOR2_X1 U9802 ( .A1(n17653), .A2(n1261), .Z(n19064) );
  XOR2_X1 U9805 ( .A1(n13199), .A2(n3475), .Z(n35987) );
  OR2_X1 U9806 ( .A1(n23202), .A2(n2430), .Z(n11704) );
  BUF_X2 U9809 ( .I(n686), .Z(n37351) );
  NAND2_X2 U9817 ( .A1(n38049), .A2(n36927), .ZN(n23873) );
  XOR2_X1 U9828 ( .A1(n20698), .A2(n7728), .Z(n25268) );
  OAI22_X2 U9834 ( .A1(n20806), .A2(n20696), .B1(n19507), .B2(n20807), .ZN(
        n20698) );
  XOR2_X1 U9837 ( .A1(n37353), .A2(n37352), .Z(n791) );
  XOR2_X1 U9843 ( .A1(n36461), .A2(n1374), .Z(n37353) );
  NAND2_X1 U9844 ( .A1(n35809), .A2(n29898), .ZN(n19540) );
  NOR2_X2 U9847 ( .A1(n38408), .A2(n1627), .ZN(n37354) );
  NOR2_X1 U9848 ( .A1(n37356), .A2(n30087), .ZN(n30084) );
  BUF_X2 U9859 ( .I(n34564), .Z(n37357) );
  NAND2_X2 U9860 ( .A1(n39499), .A2(n8196), .ZN(n13400) );
  OAI21_X1 U9863 ( .A1(n33516), .A2(n12218), .B(n1198), .ZN(n38804) );
  XOR2_X1 U9870 ( .A1(n8404), .A2(n8403), .Z(n17755) );
  XOR2_X1 U9872 ( .A1(n27748), .A2(n27716), .Z(n8404) );
  NAND2_X2 U9875 ( .A1(n4388), .A2(n21980), .ZN(n37358) );
  NAND2_X2 U9876 ( .A1(n37942), .A2(n37359), .ZN(n29270) );
  NAND2_X2 U9877 ( .A1(n37360), .A2(n21021), .ZN(n495) );
  AOI22_X2 U9878 ( .A1(n37549), .A2(n11336), .B1(n11339), .B2(n1093), .ZN(
        n37360) );
  XOR2_X1 U9882 ( .A1(n30950), .A2(n1668), .Z(n17854) );
  NAND3_X1 U9883 ( .A1(n1170), .A2(n6623), .A3(n18897), .ZN(n7270) );
  NAND2_X2 U9884 ( .A1(n35570), .A2(n37361), .ZN(n12168) );
  NOR2_X2 U9886 ( .A1(n33912), .A2(n33913), .ZN(n37361) );
  AOI22_X2 U9891 ( .A1(n1027), .A2(n24556), .B1(n24528), .B2(n12159), .ZN(
        n39120) );
  NOR2_X2 U9892 ( .A1(n24811), .A2(n12159), .ZN(n24556) );
  XOR2_X1 U9893 ( .A1(n11369), .A2(n37362), .Z(n14332) );
  XOR2_X1 U9897 ( .A1(n25302), .A2(n33005), .Z(n37362) );
  NAND2_X2 U9902 ( .A1(n20966), .A2(n37363), .ZN(n28396) );
  NAND3_X1 U9903 ( .A1(n11353), .A2(n9534), .A3(n27666), .ZN(n37363) );
  NAND2_X1 U9905 ( .A1(n11820), .A2(n9369), .ZN(n33203) );
  NAND2_X2 U9906 ( .A1(n11818), .A2(n37798), .ZN(n11820) );
  XOR2_X1 U9907 ( .A1(n22686), .A2(n22688), .Z(n16755) );
  XOR2_X1 U9908 ( .A1(n22657), .A2(n22776), .Z(n22688) );
  NOR2_X2 U9912 ( .A1(n15433), .A2(n15434), .ZN(n15368) );
  NOR2_X2 U9913 ( .A1(n30485), .A2(n3718), .ZN(n15433) );
  NAND2_X2 U9914 ( .A1(n37364), .A2(n16369), .ZN(n10570) );
  NAND3_X2 U9917 ( .A1(n23116), .A2(n23117), .A3(n12289), .ZN(n37364) );
  OR2_X1 U9925 ( .A1(n39678), .A2(n5227), .Z(n13016) );
  NAND2_X2 U9926 ( .A1(n20507), .A2(n37365), .ZN(n9030) );
  INV_X2 U9927 ( .I(n37366), .ZN(n20541) );
  XNOR2_X1 U9928 ( .A1(n10390), .A2(n10391), .ZN(n37366) );
  XOR2_X1 U9930 ( .A1(n37367), .A2(n23954), .Z(n2229) );
  XOR2_X1 U9931 ( .A1(n14345), .A2(n18160), .Z(n37367) );
  NAND2_X1 U9938 ( .A1(n10764), .A2(n37746), .ZN(n5326) );
  AOI22_X2 U9940 ( .A1(n37177), .A2(n37368), .B1(n6496), .B2(n37021), .ZN(
        n17980) );
  INV_X2 U9941 ( .I(n30000), .ZN(n37368) );
  XOR2_X1 U9943 ( .A1(n37369), .A2(n21226), .Z(Ciphertext[5]) );
  AOI22_X1 U9944 ( .A1(n9807), .A2(n29209), .B1(n18039), .B2(n11972), .ZN(
        n37369) );
  NAND3_X2 U9948 ( .A1(n39402), .A2(n32235), .A3(n37370), .ZN(n14193) );
  NAND3_X1 U9951 ( .A1(n941), .A2(n18603), .A3(n34120), .ZN(n37370) );
  NAND2_X2 U9955 ( .A1(n15586), .A2(n37371), .ZN(n32765) );
  NOR2_X2 U9960 ( .A1(n39712), .A2(n39713), .ZN(n37371) );
  INV_X2 U9974 ( .I(n36058), .ZN(n19593) );
  NOR2_X2 U9975 ( .A1(n31626), .A2(n26135), .ZN(n37372) );
  NOR2_X1 U9976 ( .A1(n6246), .A2(n4211), .ZN(n37373) );
  XOR2_X1 U9977 ( .A1(n31043), .A2(n881), .Z(n28025) );
  XOR2_X1 U9980 ( .A1(n37650), .A2(n11349), .Z(n11482) );
  AND2_X1 U9982 ( .A1(n37103), .A2(n26839), .Z(n21171) );
  XOR2_X1 U9983 ( .A1(n10221), .A2(n9151), .Z(n26208) );
  NAND2_X2 U9984 ( .A1(n6219), .A2(n1851), .ZN(n9151) );
  XOR2_X1 U9988 ( .A1(n38703), .A2(n39698), .Z(n31582) );
  XOR2_X1 U9989 ( .A1(n19289), .A2(n28821), .Z(n26566) );
  OAI21_X2 U9992 ( .A1(n20612), .A2(n20611), .B(n11848), .ZN(n8699) );
  NAND2_X2 U9993 ( .A1(n39227), .A2(n38203), .ZN(n28430) );
  NAND2_X1 U9994 ( .A1(n28267), .A2(n1206), .ZN(n18665) );
  XOR2_X1 U9995 ( .A1(n37379), .A2(n5801), .Z(n14751) );
  XOR2_X1 U9996 ( .A1(n25161), .A2(n5800), .Z(n37379) );
  XOR2_X1 U10001 ( .A1(n27655), .A2(n11564), .Z(n11563) );
  XOR2_X1 U10006 ( .A1(n25115), .A2(n24985), .Z(n25072) );
  OAI22_X2 U10007 ( .A1(n11199), .A2(n11198), .B1(n1842), .B2(n24528), .ZN(
        n25115) );
  INV_X2 U10010 ( .I(n29204), .ZN(n29208) );
  XOR2_X1 U10012 ( .A1(n33921), .A2(n37380), .Z(n36730) );
  INV_X1 U10017 ( .I(n19894), .ZN(n37380) );
  NAND2_X2 U10018 ( .A1(n39077), .A2(n25451), .ZN(n37730) );
  NOR2_X1 U10019 ( .A1(n18077), .A2(n10004), .ZN(n25045) );
  BUF_X4 U10020 ( .I(n11676), .Z(n38666) );
  INV_X2 U10023 ( .I(n7099), .ZN(n19465) );
  XNOR2_X1 U10027 ( .A1(n7102), .A2(n7100), .ZN(n7099) );
  NAND2_X2 U10029 ( .A1(n18929), .A2(n5061), .ZN(n22296) );
  NAND2_X2 U10030 ( .A1(n37559), .A2(n5504), .ZN(n18929) );
  XOR2_X1 U10044 ( .A1(n37053), .A2(n3330), .Z(n37381) );
  XOR2_X1 U10047 ( .A1(n33533), .A2(n27864), .Z(n27598) );
  NAND2_X2 U10048 ( .A1(n39565), .A2(n12017), .ZN(n33533) );
  XOR2_X1 U10053 ( .A1(n36756), .A2(n37382), .Z(n14381) );
  XOR2_X1 U10059 ( .A1(n13977), .A2(n23917), .Z(n6988) );
  XOR2_X1 U10063 ( .A1(n35181), .A2(n39209), .Z(n23917) );
  INV_X2 U10067 ( .I(n37383), .ZN(n25611) );
  XNOR2_X1 U10070 ( .A1(n10615), .A2(n1896), .ZN(n37383) );
  OR2_X1 U10071 ( .A1(n32898), .A2(n35686), .Z(n36280) );
  NOR2_X1 U10072 ( .A1(n27299), .A2(n34717), .ZN(n37385) );
  XOR2_X1 U10074 ( .A1(n26460), .A2(n26498), .Z(n26150) );
  NAND2_X2 U10075 ( .A1(n9983), .A2(n34481), .ZN(n26460) );
  NOR2_X2 U10078 ( .A1(n4824), .A2(n38779), .ZN(n13534) );
  OAI22_X2 U10081 ( .A1(n14736), .A2(n14696), .B1(n7904), .B2(n27902), .ZN(
        n38220) );
  AOI22_X2 U10082 ( .A1(n985), .A2(n1208), .B1(n759), .B2(n1439), .ZN(n27902)
         );
  XOR2_X1 U10084 ( .A1(n19642), .A2(n14264), .Z(n27712) );
  NAND2_X2 U10087 ( .A1(n35037), .A2(n9491), .ZN(n14264) );
  XOR2_X1 U10091 ( .A1(n11372), .A2(n39073), .Z(n2106) );
  NAND2_X2 U10097 ( .A1(n18890), .A2(n18889), .ZN(n39073) );
  NAND3_X2 U10099 ( .A1(n21979), .A2(n21978), .A3(n19654), .ZN(n22586) );
  NAND2_X2 U10108 ( .A1(n36525), .A2(n37386), .ZN(n12527) );
  AOI22_X2 U10113 ( .A1(n39399), .A2(n28115), .B1(n15993), .B2(n13457), .ZN(
        n37386) );
  NOR2_X2 U10127 ( .A1(n37387), .A2(n21356), .ZN(n22497) );
  AOI21_X2 U10128 ( .A1(n21354), .A2(n39368), .B(n39716), .ZN(n37387) );
  NOR2_X2 U10132 ( .A1(n21666), .A2(n21436), .ZN(n21359) );
  XOR2_X1 U10133 ( .A1(n27793), .A2(n27795), .Z(n15723) );
  XOR2_X1 U10136 ( .A1(n27776), .A2(n38964), .Z(n27793) );
  INV_X1 U10146 ( .I(n10992), .ZN(n37453) );
  INV_X1 U10150 ( .I(n37388), .ZN(n5817) );
  INV_X4 U10157 ( .I(n20597), .ZN(n978) );
  NAND2_X2 U10158 ( .A1(n10720), .A2(n2023), .ZN(n20597) );
  NOR2_X2 U10159 ( .A1(n35192), .A2(n38614), .ZN(n11108) );
  NAND2_X2 U10163 ( .A1(n37516), .A2(n6860), .ZN(n38614) );
  NAND2_X2 U10164 ( .A1(n30191), .A2(n30241), .ZN(n9173) );
  INV_X2 U10173 ( .I(n35893), .ZN(n37389) );
  OR2_X1 U10174 ( .A1(n35128), .A2(n37389), .Z(n38634) );
  NOR2_X2 U10178 ( .A1(n16576), .A2(n28153), .ZN(n28004) );
  XOR2_X1 U10182 ( .A1(n16342), .A2(n24049), .Z(n31636) );
  INV_X2 U10189 ( .I(n3903), .ZN(n28666) );
  NOR3_X2 U10190 ( .A1(n9676), .A2(n37390), .A3(n14160), .ZN(n37952) );
  NOR2_X2 U10195 ( .A1(n11717), .A2(n28402), .ZN(n28772) );
  OAI21_X2 U10196 ( .A1(n7984), .A2(n32186), .B(n7983), .ZN(n11717) );
  XOR2_X1 U10199 ( .A1(n7848), .A2(n30090), .Z(n2036) );
  NAND2_X2 U10201 ( .A1(n37719), .A2(n38818), .ZN(n7848) );
  XOR2_X1 U10202 ( .A1(n37391), .A2(n27784), .Z(n11823) );
  XOR2_X1 U10204 ( .A1(n9162), .A2(n36861), .Z(n37391) );
  INV_X4 U10206 ( .I(n15573), .ZN(n37981) );
  XNOR2_X1 U10207 ( .A1(n19187), .A2(n33439), .ZN(n37394) );
  NOR2_X2 U10208 ( .A1(n37392), .A2(n7880), .ZN(n7882) );
  XOR2_X1 U10209 ( .A1(n32994), .A2(n37394), .Z(n34764) );
  NAND2_X2 U10214 ( .A1(n37396), .A2(n37395), .ZN(n34141) );
  INV_X2 U10224 ( .I(n24639), .ZN(n37395) );
  INV_X2 U10225 ( .I(n34906), .ZN(n37396) );
  XOR2_X1 U10230 ( .A1(n10526), .A2(n9611), .Z(n37738) );
  NAND2_X2 U10231 ( .A1(n1919), .A2(n1917), .ZN(n10526) );
  NOR2_X2 U10232 ( .A1(n2202), .A2(n3683), .ZN(n39441) );
  AOI21_X1 U10233 ( .A1(n37423), .A2(n29679), .B(n9610), .ZN(n36168) );
  INV_X1 U10234 ( .I(n39268), .ZN(n37539) );
  XOR2_X1 U10237 ( .A1(n22754), .A2(n7358), .Z(n9449) );
  NAND3_X2 U10239 ( .A1(n37397), .A2(n25874), .A3(n6222), .ZN(n25878) );
  NAND2_X2 U10243 ( .A1(n32974), .A2(n36546), .ZN(n37397) );
  OR3_X1 U10244 ( .A1(n10436), .A2(n37815), .A3(n8452), .Z(n4566) );
  NAND2_X2 U10246 ( .A1(n38014), .A2(n27685), .ZN(n9848) );
  OAI21_X2 U10249 ( .A1(n19546), .A2(n35839), .B(n37398), .ZN(n21774) );
  XOR2_X1 U10251 ( .A1(n37400), .A2(n1738), .Z(Ciphertext[184]) );
  NOR2_X1 U10252 ( .A1(n15419), .A2(n39139), .ZN(n37400) );
  OAI21_X2 U10254 ( .A1(n37401), .A2(n15605), .B(n30238), .ZN(n5054) );
  INV_X2 U10257 ( .I(n29200), .ZN(n37401) );
  NAND2_X2 U10276 ( .A1(n892), .A2(n30154), .ZN(n29200) );
  OAI22_X2 U10284 ( .A1(n37178), .A2(n11945), .B1(n20884), .B2(n34117), .ZN(
        n26157) );
  OAI21_X2 U10285 ( .A1(n4317), .A2(n4318), .B(n4316), .ZN(n35727) );
  NAND2_X2 U10287 ( .A1(n5527), .A2(n33015), .ZN(n4317) );
  XOR2_X1 U10288 ( .A1(n26466), .A2(n26465), .Z(n10112) );
  XOR2_X1 U10290 ( .A1(n26394), .A2(n37024), .Z(n26465) );
  NOR2_X1 U10291 ( .A1(n37584), .A2(n25560), .ZN(n37663) );
  NAND2_X2 U10294 ( .A1(n37402), .A2(n505), .ZN(n37486) );
  NAND2_X2 U10295 ( .A1(n12428), .A2(n29451), .ZN(n37402) );
  OAI21_X2 U10307 ( .A1(n38594), .A2(n24274), .B(n7279), .ZN(n37717) );
  AOI21_X2 U10311 ( .A1(n1823), .A2(n20494), .B(n38970), .ZN(n35549) );
  XOR2_X1 U10321 ( .A1(n334), .A2(n16610), .Z(n26497) );
  OAI21_X2 U10325 ( .A1(n37821), .A2(n39781), .B(n13756), .ZN(n16610) );
  XOR2_X1 U10332 ( .A1(n5484), .A2(n38791), .Z(n2391) );
  XOR2_X1 U10335 ( .A1(n27864), .A2(n37403), .Z(n27757) );
  INV_X2 U10337 ( .I(n27738), .ZN(n37403) );
  OAI22_X2 U10341 ( .A1(n18438), .A2(n12108), .B1(n4490), .B2(n18436), .ZN(
        n27738) );
  AOI21_X2 U10355 ( .A1(n37918), .A2(n37919), .B(n37404), .ZN(n22588) );
  OAI22_X2 U10366 ( .A1(n37113), .A2(n18253), .B1(n17976), .B2(n1683), .ZN(
        n37404) );
  XOR2_X1 U10370 ( .A1(n32776), .A2(n20586), .Z(n17344) );
  AOI22_X2 U10371 ( .A1(n2156), .A2(n37200), .B1(n2154), .B2(n1349), .ZN(n2153) );
  NAND2_X2 U10372 ( .A1(n37487), .A2(n18562), .ZN(n37603) );
  XOR2_X1 U10374 ( .A1(n10525), .A2(n22452), .Z(n5516) );
  NAND2_X2 U10377 ( .A1(n4495), .A2(n4494), .ZN(n10525) );
  OR2_X1 U10378 ( .A1(n11164), .A2(n8743), .Z(n37557) );
  NAND2_X2 U10380 ( .A1(n6491), .A2(n6492), .ZN(n6490) );
  OAI21_X1 U10381 ( .A1(n29884), .A2(n17286), .B(n37405), .ZN(n17748) );
  NAND3_X2 U10382 ( .A1(n29883), .A2(n15773), .A3(n6720), .ZN(n37405) );
  XOR2_X1 U10384 ( .A1(n37406), .A2(n10107), .Z(n23083) );
  XOR2_X1 U10385 ( .A1(n22446), .A2(n21206), .Z(n37406) );
  XOR2_X1 U10386 ( .A1(n23946), .A2(n23947), .Z(n23948) );
  XOR2_X1 U10387 ( .A1(n35376), .A2(n10526), .Z(n23947) );
  XOR2_X1 U10388 ( .A1(n29243), .A2(n28824), .Z(n3707) );
  XOR2_X1 U10389 ( .A1(n29042), .A2(n39739), .Z(n29243) );
  OR2_X1 U10391 ( .A1(n31272), .A2(n20070), .Z(n39692) );
  XOR2_X1 U10393 ( .A1(n22710), .A2(n1322), .Z(n39215) );
  XOR2_X1 U10402 ( .A1(n37407), .A2(n19800), .Z(Ciphertext[87]) );
  NAND3_X1 U10414 ( .A1(n2111), .A2(n2110), .A3(n3118), .ZN(n37407) );
  NAND2_X2 U10416 ( .A1(n37408), .A2(n7717), .ZN(n28433) );
  NAND2_X2 U10417 ( .A1(n39419), .A2(n34863), .ZN(n37408) );
  OAI21_X2 U10427 ( .A1(n1564), .A2(n24816), .B(n33012), .ZN(n6408) );
  INV_X2 U10428 ( .I(n36191), .ZN(n1633) );
  NAND2_X2 U10431 ( .A1(n12698), .A2(n12697), .ZN(n36191) );
  NAND2_X2 U10434 ( .A1(n37409), .A2(n27176), .ZN(n27499) );
  OAI22_X2 U10494 ( .A1(n30732), .A2(n27174), .B1(n34562), .B2(n19132), .ZN(
        n37409) );
  NAND2_X2 U10498 ( .A1(n37892), .A2(n37410), .ZN(n39423) );
  AOI21_X2 U10503 ( .A1(n28015), .A2(n7326), .B(n20164), .ZN(n37410) );
  OAI21_X1 U10506 ( .A1(n16590), .A2(n16366), .B(n18920), .ZN(n24100) );
  INV_X2 U10508 ( .I(n32898), .ZN(n37411) );
  AND2_X1 U10509 ( .A1(n37016), .A2(n37411), .Z(n24644) );
  XOR2_X1 U10511 ( .A1(n10941), .A2(n37412), .Z(n10940) );
  XOR2_X1 U10512 ( .A1(n33524), .A2(n23727), .Z(n37412) );
  OAI21_X1 U10517 ( .A1(n37414), .A2(n9586), .B(n37413), .ZN(n28063) );
  NAND2_X1 U10520 ( .A1(n18722), .A2(n32820), .ZN(n2155) );
  XOR2_X1 U10523 ( .A1(Plaintext[61]), .A2(Key[61]), .Z(n32820) );
  NOR2_X2 U10524 ( .A1(n20267), .A2(n36620), .ZN(n11476) );
  XOR2_X1 U10525 ( .A1(n20341), .A2(n37243), .Z(n38381) );
  XOR2_X1 U10527 ( .A1(n37415), .A2(n17140), .Z(n38111) );
  XOR2_X1 U10528 ( .A1(n17850), .A2(n11525), .Z(n37415) );
  NAND2_X2 U10530 ( .A1(n11697), .A2(n18036), .ZN(n3664) );
  NOR2_X2 U10531 ( .A1(n15975), .A2(n3234), .ZN(n11697) );
  XOR2_X1 U10533 ( .A1(n33252), .A2(n26379), .Z(n26521) );
  NAND2_X2 U10534 ( .A1(n38131), .A2(n5161), .ZN(n33252) );
  INV_X2 U10535 ( .I(n24469), .ZN(n38303) );
  AND2_X1 U10536 ( .A1(n24469), .A2(n38839), .Z(n8916) );
  NOR2_X2 U10538 ( .A1(n26089), .A2(n37416), .ZN(n5164) );
  NOR2_X1 U10539 ( .A1(n32424), .A2(n7577), .ZN(n34996) );
  NAND2_X2 U10541 ( .A1(n37417), .A2(n1076), .ZN(n11279) );
  NAND2_X2 U10545 ( .A1(n37419), .A2(n274), .ZN(n37417) );
  NAND2_X2 U10548 ( .A1(n36954), .A2(n28278), .ZN(n37419) );
  XOR2_X1 U10549 ( .A1(n26231), .A2(n37476), .Z(n26311) );
  NAND2_X2 U10551 ( .A1(n3332), .A2(n26188), .ZN(n26231) );
  XOR2_X1 U10553 ( .A1(n37420), .A2(n24931), .Z(n32639) );
  XOR2_X1 U10555 ( .A1(n2653), .A2(n29051), .Z(n37420) );
  XOR2_X1 U10556 ( .A1(n19156), .A2(n25292), .Z(n36138) );
  INV_X1 U10557 ( .I(n38909), .ZN(n34156) );
  OR2_X1 U10559 ( .A1(n38909), .A2(n25345), .Z(n18217) );
  BUF_X2 U10564 ( .I(n16048), .Z(n35001) );
  BUF_X2 U10566 ( .I(n19593), .Z(n37421) );
  XOR2_X1 U10569 ( .A1(n37422), .A2(n38870), .Z(n38259) );
  XOR2_X1 U10576 ( .A1(n27725), .A2(n37242), .Z(n37422) );
  XOR2_X1 U10577 ( .A1(n26569), .A2(n39691), .Z(n32844) );
  NAND2_X1 U10583 ( .A1(n37493), .A2(n18478), .ZN(n32574) );
  BUF_X4 U10585 ( .I(n20936), .Z(n35537) );
  NAND2_X1 U10586 ( .A1(n29674), .A2(n14522), .ZN(n37423) );
  XOR2_X1 U10588 ( .A1(n5789), .A2(n37424), .Z(n3675) );
  XOR2_X1 U10601 ( .A1(n8003), .A2(n11102), .Z(n37424) );
  AOI21_X2 U10604 ( .A1(n10735), .A2(n27307), .B(n37425), .ZN(n5750) );
  NOR2_X1 U10607 ( .A1(n14041), .A2(n17166), .ZN(n37425) );
  NAND2_X2 U10610 ( .A1(n36222), .A2(n27306), .ZN(n14041) );
  NAND2_X2 U10620 ( .A1(n16129), .A2(n14420), .ZN(n22277) );
  OR2_X1 U10623 ( .A1(n309), .A2(n28771), .Z(n35776) );
  XOR2_X1 U10624 ( .A1(n23563), .A2(n37426), .Z(n35300) );
  XOR2_X1 U10627 ( .A1(n39239), .A2(n23562), .Z(n37426) );
  XOR2_X1 U10628 ( .A1(n35220), .A2(n10791), .Z(n3589) );
  NAND2_X2 U10629 ( .A1(n14874), .A2(n24754), .ZN(n10791) );
  NOR2_X1 U10634 ( .A1(n3169), .A2(n3170), .ZN(n38757) );
  NAND2_X2 U10637 ( .A1(n14082), .A2(n25674), .ZN(n14083) );
  NOR2_X2 U10638 ( .A1(n11596), .A2(n11594), .ZN(n12141) );
  AOI21_X2 U10640 ( .A1(n11597), .A2(n29317), .B(n29263), .ZN(n11596) );
  AND3_X1 U10644 ( .A1(n12235), .A2(n18466), .A3(n19658), .Z(n4785) );
  XOR2_X1 U10645 ( .A1(n27549), .A2(n27679), .Z(n27725) );
  NAND2_X2 U10647 ( .A1(n16751), .A2(n15945), .ZN(n25097) );
  NAND3_X2 U10649 ( .A1(n16990), .A2(n38738), .A3(n38942), .ZN(n16751) );
  XOR2_X1 U10652 ( .A1(n19561), .A2(n27823), .Z(n13035) );
  NAND2_X2 U10653 ( .A1(n34989), .A2(n33016), .ZN(n19561) );
  BUF_X2 U10655 ( .I(n18595), .Z(n37428) );
  XOR2_X1 U10656 ( .A1(n31240), .A2(n23937), .Z(n34439) );
  XOR2_X1 U10658 ( .A1(n39412), .A2(n23938), .Z(n31240) );
  NAND2_X2 U10660 ( .A1(n37429), .A2(n22032), .ZN(n22348) );
  OAI21_X2 U10661 ( .A1(n19012), .A2(n7916), .B(n19011), .ZN(n37429) );
  OAI21_X1 U10662 ( .A1(n36548), .A2(n29627), .B(n35405), .ZN(n37430) );
  NAND2_X2 U10665 ( .A1(n12543), .A2(n18960), .ZN(n28652) );
  AOI21_X2 U10672 ( .A1(n27115), .A2(n33088), .B(n19334), .ZN(n37433) );
  NOR2_X2 U10674 ( .A1(n37435), .A2(n16132), .ZN(n12396) );
  XOR2_X1 U10675 ( .A1(n37874), .A2(n31515), .Z(n21186) );
  AOI21_X2 U10679 ( .A1(n13028), .A2(n28653), .B(n13027), .ZN(n37874) );
  NAND3_X2 U10681 ( .A1(n38536), .A2(n38534), .A3(n38252), .ZN(n21066) );
  XOR2_X1 U10689 ( .A1(n31137), .A2(n18650), .Z(n5566) );
  XOR2_X1 U10691 ( .A1(n27687), .A2(n19606), .Z(n18650) );
  XOR2_X1 U10692 ( .A1(n22635), .A2(n37434), .Z(n17430) );
  XOR2_X1 U10693 ( .A1(n36641), .A2(n22620), .Z(n37434) );
  AOI21_X2 U10694 ( .A1(n2751), .A2(n5674), .B(n34310), .ZN(n37476) );
  OR2_X2 U10695 ( .A1(n37104), .A2(n26988), .Z(n26989) );
  OR2_X1 U10697 ( .A1(n29885), .A2(n6720), .Z(n29884) );
  OAI22_X2 U10701 ( .A1(n32539), .A2(n35342), .B1(n17148), .B2(n19093), .ZN(
        n6720) );
  NAND2_X2 U10702 ( .A1(n30191), .A2(n30245), .ZN(n35391) );
  INV_X2 U10703 ( .I(n883), .ZN(n1070) );
  XNOR2_X1 U10704 ( .A1(n4362), .A2(n4364), .ZN(n883) );
  XOR2_X1 U10708 ( .A1(n39100), .A2(n30648), .Z(n33621) );
  AOI22_X2 U10709 ( .A1(n33510), .A2(n14480), .B1(n17447), .B2(n28093), .ZN(
        n28129) );
  OAI22_X2 U10710 ( .A1(n18527), .A2(n14594), .B1(n20230), .B2(n33196), .ZN(
        n37435) );
  NAND2_X2 U10711 ( .A1(n38435), .A2(n34799), .ZN(n12306) );
  XOR2_X1 U10714 ( .A1(n37436), .A2(n37380), .Z(Ciphertext[35]) );
  NOR2_X1 U10715 ( .A1(n15957), .A2(n15956), .ZN(n37436) );
  XOR2_X1 U10719 ( .A1(n17159), .A2(n12231), .Z(n13724) );
  XOR2_X1 U10720 ( .A1(n37437), .A2(n19681), .Z(Ciphertext[14]) );
  NAND2_X1 U10721 ( .A1(n15027), .A2(n15026), .ZN(n37437) );
  INV_X4 U10723 ( .I(n25611), .ZN(n34010) );
  XOR2_X1 U10724 ( .A1(n15078), .A2(n26260), .Z(n15077) );
  INV_X2 U10725 ( .I(n26412), .ZN(n15078) );
  XOR2_X1 U10727 ( .A1(n26519), .A2(n26259), .Z(n26412) );
  XOR2_X1 U10729 ( .A1(n37438), .A2(n9315), .Z(n37829) );
  XOR2_X1 U10730 ( .A1(n27774), .A2(n13703), .Z(n37438) );
  NOR2_X2 U10737 ( .A1(n35434), .A2(n37439), .ZN(n4184) );
  AOI21_X2 U10738 ( .A1(n10013), .A2(n24847), .B(n19630), .ZN(n24730) );
  NAND2_X2 U10740 ( .A1(n37168), .A2(n13625), .ZN(n24847) );
  AOI21_X2 U10749 ( .A1(n36590), .A2(n1408), .B(n37440), .ZN(n2013) );
  NOR3_X1 U10757 ( .A1(n1962), .A2(n20866), .A3(n20673), .ZN(n37440) );
  XOR2_X1 U10758 ( .A1(n26379), .A2(n19902), .Z(n26380) );
  NAND2_X2 U10760 ( .A1(n21265), .A2(n34742), .ZN(n26379) );
  XOR2_X1 U10763 ( .A1(n9858), .A2(n17890), .Z(n26376) );
  NAND2_X2 U10764 ( .A1(n10016), .A2(n12941), .ZN(n9858) );
  NAND2_X2 U10766 ( .A1(n34217), .A2(n16250), .ZN(n25990) );
  NAND2_X2 U10771 ( .A1(n20337), .A2(n37441), .ZN(n25951) );
  NAND2_X2 U10772 ( .A1(n25564), .A2(n39458), .ZN(n37441) );
  XOR2_X1 U10773 ( .A1(n4624), .A2(n22488), .Z(n22760) );
  NAND2_X2 U10776 ( .A1(n3267), .A2(n3265), .ZN(n4624) );
  XOR2_X1 U10779 ( .A1(n37442), .A2(n8826), .Z(n37587) );
  XOR2_X1 U10783 ( .A1(n31773), .A2(n23801), .Z(n37442) );
  NOR3_X1 U10785 ( .A1(n27288), .A2(n34279), .A3(n39417), .ZN(n36314) );
  NAND2_X2 U10786 ( .A1(n4641), .A2(n36538), .ZN(n39417) );
  NOR2_X2 U10787 ( .A1(n35119), .A2(n35118), .ZN(n15945) );
  OR2_X1 U10791 ( .A1(n31760), .A2(n13872), .Z(n39273) );
  XOR2_X1 U10793 ( .A1(n36423), .A2(n38569), .Z(n31760) );
  INV_X2 U10795 ( .I(n38880), .ZN(n1612) );
  XOR2_X1 U10797 ( .A1(n38880), .A2(n37443), .Z(n23357) );
  NAND2_X2 U10802 ( .A1(n39276), .A2(n2933), .ZN(n38880) );
  NOR2_X2 U10805 ( .A1(n12966), .A2(n7225), .ZN(n39788) );
  NOR2_X2 U10810 ( .A1(n23137), .A2(n23136), .ZN(n12966) );
  OAI22_X2 U10814 ( .A1(n7209), .A2(n17067), .B1(n20795), .B2(n7210), .ZN(
        n35893) );
  NAND2_X1 U10815 ( .A1(n14900), .A2(n2500), .ZN(n14001) );
  AOI22_X2 U10817 ( .A1(n31353), .A2(n15792), .B1(n28560), .B2(n28617), .ZN(
        n2500) );
  OAI21_X2 U10818 ( .A1(n37444), .A2(n36643), .B(n31942), .ZN(n18223) );
  NOR2_X2 U10820 ( .A1(n13366), .A2(n36517), .ZN(n37444) );
  NAND2_X1 U10821 ( .A1(n8651), .A2(n19448), .ZN(n16049) );
  XOR2_X1 U10823 ( .A1(n10076), .A2(n26520), .Z(n26258) );
  OAI21_X2 U10824 ( .A1(n14579), .A2(n15177), .B(n33764), .ZN(n10076) );
  AND2_X1 U10830 ( .A1(n37934), .A2(n37651), .Z(n14645) );
  AOI21_X2 U10831 ( .A1(n7239), .A2(n7237), .B(n7234), .ZN(n33263) );
  XOR2_X1 U10832 ( .A1(n37446), .A2(n29282), .Z(Ciphertext[21]) );
  NAND3_X1 U10837 ( .A1(n29280), .A2(n29281), .A3(n29279), .ZN(n37446) );
  XOR2_X1 U10839 ( .A1(n8402), .A2(n35986), .Z(n27716) );
  XOR2_X1 U10840 ( .A1(n37447), .A2(n1714), .Z(Ciphertext[121]) );
  AOI22_X1 U10841 ( .A1(n29877), .A2(n29876), .B1(n29880), .B2(n29889), .ZN(
        n37447) );
  INV_X4 U10842 ( .I(n1548), .ZN(n33022) );
  NAND2_X1 U10851 ( .A1(n1284), .A2(n17081), .ZN(n38097) );
  XOR2_X1 U10854 ( .A1(n35721), .A2(n37448), .Z(n39611) );
  INV_X4 U10856 ( .I(n2678), .ZN(n2534) );
  INV_X4 U10859 ( .I(n32802), .ZN(n39258) );
  INV_X4 U10860 ( .I(n8131), .ZN(n35357) );
  NAND2_X2 U10862 ( .A1(n33059), .A2(n6588), .ZN(n8131) );
  XOR2_X1 U10864 ( .A1(n10329), .A2(n25180), .Z(n10333) );
  XOR2_X1 U10879 ( .A1(n1259), .A2(n11698), .Z(n10329) );
  NAND2_X1 U10880 ( .A1(n38906), .A2(n30799), .ZN(n28184) );
  OR2_X1 U10881 ( .A1(n10266), .A2(n19435), .Z(n12349) );
  NAND2_X1 U10889 ( .A1(n33646), .A2(n20879), .ZN(n34285) );
  NOR2_X1 U10890 ( .A1(n38568), .A2(n37903), .ZN(n12776) );
  NAND2_X1 U10891 ( .A1(n24273), .A2(n24272), .ZN(n35959) );
  XOR2_X1 U10895 ( .A1(n22748), .A2(n12901), .Z(n12898) );
  XOR2_X1 U10899 ( .A1(n22411), .A2(n22430), .Z(n22748) );
  NAND2_X2 U10900 ( .A1(n19476), .A2(n1755), .ZN(n30720) );
  NAND2_X2 U10901 ( .A1(n31312), .A2(n37449), .ZN(n34533) );
  OR2_X1 U10904 ( .A1(n26019), .A2(n26020), .Z(n37449) );
  NAND3_X2 U10905 ( .A1(n37450), .A2(n2130), .A3(n2129), .ZN(n36496) );
  NAND2_X1 U10906 ( .A1(n26624), .A2(n35764), .ZN(n37450) );
  XOR2_X1 U10910 ( .A1(n17908), .A2(n22486), .Z(n19781) );
  XOR2_X1 U10911 ( .A1(n22485), .A2(n22484), .Z(n17908) );
  INV_X1 U10912 ( .I(n39769), .ZN(n34070) );
  NAND2_X2 U10913 ( .A1(n19544), .A2(n12081), .ZN(n39769) );
  XOR2_X1 U10914 ( .A1(n22392), .A2(n1660), .Z(n38118) );
  NAND3_X2 U10916 ( .A1(n37453), .A2(n38855), .A3(n37452), .ZN(n37927) );
  NAND2_X1 U10919 ( .A1(n5383), .A2(n12527), .ZN(n37452) );
  NAND3_X2 U10929 ( .A1(n32283), .A2(n34664), .A3(n2356), .ZN(n16094) );
  NAND2_X2 U10934 ( .A1(n14052), .A2(n8499), .ZN(n35981) );
  AOI22_X2 U10935 ( .A1(n38047), .A2(n20981), .B1(n27286), .B2(n10284), .ZN(
        n27501) );
  NAND2_X2 U10938 ( .A1(n465), .A2(n8758), .ZN(n15423) );
  OAI22_X2 U10939 ( .A1(n10487), .A2(n22344), .B1(n22170), .B2(n22342), .ZN(
        n347) );
  NAND2_X2 U10941 ( .A1(n37455), .A2(n26835), .ZN(n8105) );
  NAND2_X2 U10942 ( .A1(n26722), .A2(n9269), .ZN(n37455) );
  INV_X1 U10945 ( .I(n2437), .ZN(n38076) );
  NOR2_X1 U10948 ( .A1(n34430), .A2(n24394), .ZN(n21319) );
  XOR2_X1 U10949 ( .A1(n19536), .A2(n23861), .Z(n23688) );
  AOI21_X2 U10951 ( .A1(n23447), .A2(n2084), .B(n10078), .ZN(n23861) );
  NAND3_X1 U10952 ( .A1(n30230), .A2(n30228), .A3(n30229), .ZN(n37636) );
  NAND2_X2 U10953 ( .A1(n36243), .A2(n35535), .ZN(n19203) );
  XOR2_X1 U10956 ( .A1(n37456), .A2(n9994), .Z(n4786) );
  XOR2_X1 U10957 ( .A1(n13176), .A2(n11479), .Z(n37456) );
  NAND2_X2 U10959 ( .A1(n24138), .A2(n24139), .ZN(n39279) );
  OR2_X1 U10960 ( .A1(n24639), .A2(n24250), .Z(n20800) );
  NOR2_X1 U10962 ( .A1(n9758), .A2(n30445), .ZN(n14916) );
  OAI22_X2 U10965 ( .A1(n2769), .A2(n2768), .B1(n2767), .B2(n36225), .ZN(
        n16180) );
  XOR2_X1 U10969 ( .A1(n38989), .A2(n21154), .Z(n233) );
  OAI22_X2 U10978 ( .A1(n36624), .A2(n4636), .B1(n4132), .B2(n17353), .ZN(
        n17624) );
  INV_X4 U10981 ( .I(n2747), .ZN(n38794) );
  XOR2_X1 U10983 ( .A1(n20501), .A2(n37457), .Z(n14000) );
  XOR2_X1 U10984 ( .A1(n10153), .A2(n31999), .Z(n37457) );
  NOR2_X2 U10986 ( .A1(n21627), .A2(n10085), .ZN(n7357) );
  XOR2_X1 U10987 ( .A1(n18051), .A2(n8833), .Z(n4077) );
  NOR2_X2 U10991 ( .A1(n38672), .A2(n31831), .ZN(n8833) );
  AOI21_X1 U10993 ( .A1(n5424), .A2(n3538), .B(n17583), .ZN(n39555) );
  NAND3_X2 U10994 ( .A1(n32374), .A2(n3461), .A3(n28075), .ZN(n17583) );
  INV_X2 U10995 ( .I(n16180), .ZN(n30111) );
  XOR2_X1 U10996 ( .A1(n23885), .A2(n24025), .Z(n23743) );
  AOI21_X2 U11002 ( .A1(n22873), .A2(n16047), .B(n37458), .ZN(n23623) );
  OAI22_X2 U11004 ( .A1(n22872), .A2(n16047), .B1(n20776), .B2(n961), .ZN(
        n37458) );
  INV_X2 U11007 ( .I(n37459), .ZN(n23162) );
  XOR2_X1 U11008 ( .A1(n37461), .A2(n10396), .Z(n13862) );
  XOR2_X1 U11010 ( .A1(n15164), .A2(n36656), .Z(n37461) );
  XOR2_X1 U11014 ( .A1(n27580), .A2(n29805), .Z(n10399) );
  NAND2_X2 U11016 ( .A1(n37978), .A2(n33160), .ZN(n27580) );
  NAND2_X2 U11019 ( .A1(n31362), .A2(n692), .ZN(n25954) );
  NOR3_X1 U11027 ( .A1(n39048), .A2(n31133), .A3(n25820), .ZN(n25821) );
  NOR2_X2 U11029 ( .A1(n37464), .A2(n36682), .ZN(n7291) );
  NOR2_X1 U11030 ( .A1(n2967), .A2(n2968), .ZN(n37464) );
  XNOR2_X1 U11036 ( .A1(n15368), .A2(n6026), .ZN(n39259) );
  NAND2_X1 U11037 ( .A1(n9415), .A2(n27428), .ZN(n17718) );
  INV_X2 U11038 ( .I(n35427), .ZN(n27428) );
  NAND2_X2 U11042 ( .A1(n37766), .A2(n39508), .ZN(n35427) );
  NAND2_X2 U11051 ( .A1(n37734), .A2(n30220), .ZN(n29202) );
  OAI21_X2 U11053 ( .A1(n37250), .A2(n37465), .B(n27228), .ZN(n27592) );
  OR2_X1 U11054 ( .A1(n29208), .A2(n15535), .Z(n29207) );
  XNOR2_X1 U11055 ( .A1(n38192), .A2(n7247), .ZN(n9960) );
  NAND2_X2 U11056 ( .A1(n7243), .A2(n7241), .ZN(n7247) );
  INV_X2 U11059 ( .I(n38848), .ZN(n34720) );
  NAND2_X2 U11061 ( .A1(n37975), .A2(n37472), .ZN(n38848) );
  XOR2_X1 U11062 ( .A1(n25206), .A2(n25208), .Z(n6658) );
  BUF_X2 U11063 ( .I(n34345), .Z(n37466) );
  NAND2_X2 U11068 ( .A1(n39533), .A2(n38373), .ZN(n23982) );
  OR2_X2 U11071 ( .A1(n39639), .A2(n20361), .Z(n21854) );
  NAND2_X1 U11080 ( .A1(n15376), .A2(n19599), .ZN(n39740) );
  INV_X2 U11083 ( .I(n9387), .ZN(n8792) );
  NAND2_X2 U11084 ( .A1(n7998), .A2(n7999), .ZN(n9387) );
  NAND2_X1 U11086 ( .A1(n10019), .A2(n37999), .ZN(n24689) );
  NAND2_X2 U11087 ( .A1(n37468), .A2(n37467), .ZN(n24412) );
  INV_X1 U11090 ( .I(n31403), .ZN(n37467) );
  INV_X2 U11093 ( .I(n24408), .ZN(n37468) );
  XOR2_X1 U11097 ( .A1(n19600), .A2(n7032), .Z(n7031) );
  NAND2_X2 U11098 ( .A1(n37114), .A2(n37469), .ZN(n6068) );
  NOR2_X2 U11108 ( .A1(n4369), .A2(n37470), .ZN(n37469) );
  NOR2_X2 U11111 ( .A1(n28639), .A2(n39355), .ZN(n37470) );
  NOR2_X2 U11112 ( .A1(n37471), .A2(n8963), .ZN(n4584) );
  NOR2_X2 U11116 ( .A1(n1495), .A2(n8311), .ZN(n37471) );
  NAND2_X2 U11125 ( .A1(n9218), .A2(n20326), .ZN(n20605) );
  XOR2_X1 U11127 ( .A1(n25164), .A2(n8240), .Z(n31151) );
  XOR2_X1 U11132 ( .A1(n13076), .A2(n15625), .Z(n25164) );
  XOR2_X1 U11133 ( .A1(n29140), .A2(n29139), .Z(n5347) );
  OAI22_X1 U11138 ( .A1(n30080), .A2(n30070), .B1(n6453), .B2(n30066), .ZN(
        n30730) );
  NOR2_X2 U11143 ( .A1(n4168), .A2(n4379), .ZN(n30080) );
  NAND2_X2 U11145 ( .A1(n39194), .A2(n9862), .ZN(n23441) );
  NAND2_X2 U11148 ( .A1(n3047), .A2(n3046), .ZN(n39194) );
  NAND2_X1 U11152 ( .A1(n36669), .A2(n13610), .ZN(n39735) );
  AOI21_X1 U11157 ( .A1(n7797), .A2(n37473), .B(n7792), .ZN(n32903) );
  NAND2_X1 U11159 ( .A1(n7795), .A2(n7796), .ZN(n37473) );
  AND2_X1 U11160 ( .A1(n18164), .A2(n32622), .Z(n11646) );
  XOR2_X1 U11161 ( .A1(n4341), .A2(n29289), .Z(n17957) );
  NAND2_X2 U11163 ( .A1(n6093), .A2(n12342), .ZN(n4341) );
  NAND2_X1 U11166 ( .A1(n38595), .A2(n38115), .ZN(n38594) );
  NOR2_X2 U11174 ( .A1(n39513), .A2(n37475), .ZN(n37474) );
  INV_X2 U11182 ( .I(n38674), .ZN(n37475) );
  BUF_X4 U11183 ( .I(n3455), .Z(n38437) );
  NOR2_X2 U11184 ( .A1(n4155), .A2(n19750), .ZN(n4927) );
  NAND2_X2 U11187 ( .A1(n11890), .A2(n10254), .ZN(n4155) );
  NAND2_X2 U11188 ( .A1(n6913), .A2(n6912), .ZN(n39196) );
  INV_X4 U11192 ( .I(n19465), .ZN(n37604) );
  XOR2_X1 U11199 ( .A1(n6535), .A2(n6537), .Z(n11428) );
  AOI21_X1 U11201 ( .A1(n37819), .A2(n37613), .B(n19740), .ZN(n12526) );
  OAI21_X2 U11202 ( .A1(n20628), .A2(n20626), .B(n14486), .ZN(n37613) );
  NOR2_X1 U11209 ( .A1(n9547), .A2(n626), .ZN(n6483) );
  INV_X2 U11210 ( .I(n32518), .ZN(n626) );
  XOR2_X1 U11211 ( .A1(n6988), .A2(n6985), .Z(n32518) );
  NAND2_X1 U11214 ( .A1(n6645), .A2(n37478), .ZN(n3723) );
  NAND2_X2 U11220 ( .A1(n6646), .A2(n38725), .ZN(n37478) );
  XOR2_X1 U11224 ( .A1(n25089), .A2(n37479), .Z(n36537) );
  XOR2_X1 U11226 ( .A1(n39320), .A2(n15912), .Z(n37479) );
  XOR2_X1 U11227 ( .A1(n1555), .A2(n25241), .Z(n25089) );
  XOR2_X1 U11232 ( .A1(n38710), .A2(n29817), .Z(n29936) );
  XOR2_X1 U11233 ( .A1(n29043), .A2(n31782), .Z(n29817) );
  XOR2_X1 U11234 ( .A1(n23776), .A2(n23829), .Z(n24058) );
  NAND3_X2 U11236 ( .A1(n23239), .A2(n23241), .A3(n23240), .ZN(n23776) );
  NAND2_X2 U11237 ( .A1(n9823), .A2(n23238), .ZN(n23460) );
  NAND2_X2 U11239 ( .A1(n35347), .A2(n14875), .ZN(n9823) );
  NAND2_X2 U11240 ( .A1(n30775), .A2(n23873), .ZN(n6583) );
  NAND2_X2 U11242 ( .A1(n35278), .A2(n35279), .ZN(n30775) );
  NAND2_X2 U11247 ( .A1(n11852), .A2(n4058), .ZN(n21925) );
  XOR2_X1 U11249 ( .A1(n11099), .A2(n32127), .Z(n36253) );
  XOR2_X1 U11251 ( .A1(n18498), .A2(n39614), .Z(n11099) );
  XOR2_X1 U11253 ( .A1(n1895), .A2(n11950), .Z(n1897) );
  NAND2_X2 U11254 ( .A1(n198), .A2(n199), .ZN(n1895) );
  NOR2_X2 U11255 ( .A1(n37482), .A2(n37481), .ZN(n7144) );
  NOR2_X2 U11258 ( .A1(n23229), .A2(n23749), .ZN(n37481) );
  XOR2_X1 U11261 ( .A1(n22601), .A2(n37466), .Z(n13652) );
  AOI21_X2 U11263 ( .A1(n5557), .A2(n8518), .B(n5556), .ZN(n34345) );
  NAND2_X1 U11266 ( .A1(n39638), .A2(n14170), .ZN(n26860) );
  XOR2_X1 U11269 ( .A1(n39612), .A2(n39611), .Z(n39638) );
  INV_X2 U11270 ( .I(n37483), .ZN(n10642) );
  XNOR2_X1 U11273 ( .A1(n11099), .A2(n32127), .ZN(n37483) );
  NAND2_X2 U11274 ( .A1(n37485), .A2(n37506), .ZN(n9859) );
  AND2_X1 U11275 ( .A1(n14840), .A2(n25369), .Z(n37485) );
  NAND2_X2 U11279 ( .A1(n37486), .A2(n2132), .ZN(n29473) );
  INV_X2 U11281 ( .I(n36177), .ZN(n27372) );
  NAND2_X2 U11283 ( .A1(n33853), .A2(n3255), .ZN(n36177) );
  NAND3_X1 U11285 ( .A1(n24788), .A2(n8430), .A3(n18148), .ZN(n18564) );
  XOR2_X1 U11287 ( .A1(n6403), .A2(n33231), .Z(n6402) );
  NOR3_X2 U11288 ( .A1(n3644), .A2(n38448), .A3(n1049), .ZN(n10743) );
  INV_X4 U11289 ( .I(n2654), .ZN(n3644) );
  NOR2_X2 U11290 ( .A1(n34059), .A2(n35860), .ZN(n2654) );
  NAND2_X2 U11291 ( .A1(n32614), .A2(n38967), .ZN(n18850) );
  XOR2_X1 U11292 ( .A1(n5116), .A2(n24076), .Z(n10683) );
  NAND2_X1 U11295 ( .A1(n11196), .A2(n24447), .ZN(n38312) );
  NAND3_X2 U11297 ( .A1(n35753), .A2(n10842), .A3(n10841), .ZN(n12362) );
  XOR2_X1 U11300 ( .A1(n37489), .A2(n15311), .Z(n10860) );
  XOR2_X1 U11302 ( .A1(n13236), .A2(n10862), .Z(n37489) );
  AOI22_X2 U11303 ( .A1(n30862), .A2(n24723), .B1(n32398), .B2(n4323), .ZN(
        n18600) );
  OAI22_X2 U11304 ( .A1(n24723), .A2(n24717), .B1(n5056), .B2(n24719), .ZN(
        n4323) );
  NAND2_X2 U11308 ( .A1(n34317), .A2(n37490), .ZN(n16226) );
  OAI21_X2 U11309 ( .A1(n22235), .A2(n19261), .B(n18064), .ZN(n37491) );
  XOR2_X1 U11310 ( .A1(n37492), .A2(n29157), .Z(n8443) );
  XOR2_X1 U11317 ( .A1(n16334), .A2(n5041), .Z(n37492) );
  OAI22_X2 U11320 ( .A1(n38357), .A2(n39800), .B1(n25379), .B2(n19863), .ZN(
        n38356) );
  XOR2_X1 U11325 ( .A1(n23685), .A2(n19953), .Z(n4327) );
  NAND3_X2 U11327 ( .A1(n4287), .A2(n4290), .A3(n4288), .ZN(n23685) );
  XOR2_X1 U11336 ( .A1(n26324), .A2(n26247), .Z(n2069) );
  XOR2_X1 U11345 ( .A1(n26554), .A2(n7402), .Z(n26247) );
  NAND2_X2 U11346 ( .A1(n23333), .A2(n17167), .ZN(n37493) );
  AND2_X1 U11347 ( .A1(n36685), .A2(n28591), .Z(n4833) );
  NAND3_X2 U11352 ( .A1(n17), .A2(n28162), .A3(n11742), .ZN(n36685) );
  XOR2_X1 U11355 ( .A1(n17462), .A2(n23675), .Z(n24019) );
  NAND2_X2 U11356 ( .A1(n10570), .A2(n23118), .ZN(n17462) );
  NAND2_X2 U11358 ( .A1(n23094), .A2(n6466), .ZN(n7026) );
  NOR2_X2 U11362 ( .A1(n9586), .A2(n28430), .ZN(n39190) );
  INV_X2 U11364 ( .I(n32472), .ZN(n585) );
  XOR2_X1 U11365 ( .A1(n38781), .A2(n37494), .Z(n38597) );
  XOR2_X1 U11366 ( .A1(n742), .A2(n37223), .Z(n37494) );
  AOI21_X2 U11368 ( .A1(n1521), .A2(n930), .B(n7258), .ZN(n36568) );
  XOR2_X1 U11374 ( .A1(n10926), .A2(n10928), .Z(n20838) );
  NAND2_X1 U11377 ( .A1(n18694), .A2(n38477), .ZN(n38476) );
  XOR2_X1 U11380 ( .A1(n2896), .A2(n24552), .Z(n33946) );
  NAND2_X2 U11381 ( .A1(n4159), .A2(n31080), .ZN(n16182) );
  INV_X1 U11382 ( .I(n29856), .ZN(n37497) );
  NAND2_X2 U11384 ( .A1(n23390), .A2(n16013), .ZN(n23453) );
  XOR2_X1 U11389 ( .A1(n37495), .A2(n18751), .Z(n22781) );
  XOR2_X1 U11393 ( .A1(n33862), .A2(n22776), .Z(n37495) );
  XOR2_X1 U11395 ( .A1(n10370), .A2(n10722), .Z(n10371) );
  AOI21_X2 U11403 ( .A1(n12638), .A2(n12639), .B(n36241), .ZN(n10370) );
  INV_X2 U11408 ( .I(n13379), .ZN(n3988) );
  OAI21_X2 U11410 ( .A1(n36914), .A2(n34470), .B(n27982), .ZN(n13379) );
  NOR3_X1 U11415 ( .A1(n22925), .A2(n6327), .A3(n38229), .ZN(n32753) );
  XOR2_X1 U11416 ( .A1(n17159), .A2(n17493), .Z(n9923) );
  XOR2_X1 U11420 ( .A1(n1065), .A2(n15581), .Z(n17493) );
  XOR2_X1 U11423 ( .A1(n36916), .A2(n10132), .Z(n28262) );
  OAI21_X2 U11427 ( .A1(n33706), .A2(n23084), .B(n37496), .ZN(n3713) );
  AOI22_X2 U11431 ( .A1(n23184), .A2(n14396), .B1(n14725), .B2(n35567), .ZN(
        n37496) );
  AOI22_X1 U11434 ( .A1(n37497), .A2(n1054), .B1(n5579), .B2(n29858), .ZN(
        n19872) );
  NAND2_X2 U11438 ( .A1(n2347), .A2(n3861), .ZN(n29856) );
  NAND2_X2 U11442 ( .A1(n39538), .A2(n31937), .ZN(n36058) );
  NAND2_X2 U11443 ( .A1(n6921), .A2(n6920), .ZN(n30033) );
  XOR2_X1 U11445 ( .A1(n23590), .A2(n39209), .Z(n17775) );
  NAND2_X2 U11446 ( .A1(n38025), .A2(n38024), .ZN(n39209) );
  XOR2_X1 U11449 ( .A1(n27837), .A2(n27719), .Z(n18048) );
  XOR2_X1 U11450 ( .A1(n1468), .A2(n35229), .Z(n27719) );
  NAND2_X1 U11452 ( .A1(n21039), .A2(n17400), .ZN(n25958) );
  NAND3_X1 U11457 ( .A1(n35333), .A2(n5908), .A3(n26039), .ZN(n36766) );
  NAND2_X2 U11460 ( .A1(n25464), .A2(n34877), .ZN(n35333) );
  AOI22_X2 U11462 ( .A1(n17191), .A2(n28755), .B1(n32791), .B2(n16691), .ZN(
        n14971) );
  AOI22_X2 U11467 ( .A1(n34465), .A2(n34464), .B1(n1546), .B2(n25501), .ZN(
        n25288) );
  OAI22_X2 U11469 ( .A1(n6592), .A2(n37025), .B1(n14081), .B2(n25434), .ZN(
        n25501) );
  NAND3_X2 U11474 ( .A1(n2682), .A2(n2683), .A3(n23386), .ZN(n2685) );
  XOR2_X1 U11475 ( .A1(n6984), .A2(n25), .Z(n34397) );
  XOR2_X1 U11478 ( .A1(n27698), .A2(n27667), .Z(n27001) );
  XOR2_X1 U11483 ( .A1(n19396), .A2(n9315), .Z(n27698) );
  INV_X2 U11484 ( .I(n28089), .ZN(n8207) );
  NOR3_X1 U11485 ( .A1(n36796), .A2(n11614), .A3(n8743), .ZN(n27653) );
  INV_X4 U11486 ( .I(n3669), .ZN(n17501) );
  NAND2_X2 U11488 ( .A1(n35710), .A2(n39486), .ZN(n3669) );
  NAND2_X2 U11490 ( .A1(n37643), .A2(n19615), .ZN(n26824) );
  INV_X2 U11494 ( .I(n37501), .ZN(n12663) );
  XNOR2_X1 U11495 ( .A1(n11235), .A2(n11237), .ZN(n37501) );
  INV_X2 U11496 ( .I(n26328), .ZN(n1515) );
  NAND2_X2 U11498 ( .A1(n11533), .A2(n33258), .ZN(n26328) );
  NAND2_X1 U11500 ( .A1(n15290), .A2(n23173), .ZN(n6645) );
  NAND2_X2 U11504 ( .A1(n36911), .A2(n5101), .ZN(n8260) );
  INV_X2 U11510 ( .I(n28389), .ZN(n34702) );
  NOR2_X1 U11511 ( .A1(n28081), .A2(n28080), .ZN(n28082) );
  NAND2_X2 U11512 ( .A1(n37503), .A2(n3904), .ZN(n39020) );
  NAND3_X2 U11513 ( .A1(n37960), .A2(n15334), .A3(n39235), .ZN(n37503) );
  NAND2_X2 U11515 ( .A1(n37504), .A2(n24481), .ZN(n19713) );
  XOR2_X1 U11518 ( .A1(n4436), .A2(n37505), .Z(n39427) );
  XOR2_X1 U11519 ( .A1(n22600), .A2(n3528), .Z(n37505) );
  XOR2_X1 U11521 ( .A1(n1616), .A2(n38468), .Z(n6468) );
  NOR2_X2 U11522 ( .A1(n38794), .A2(n934), .ZN(n15527) );
  NAND2_X1 U11525 ( .A1(n25368), .A2(n17855), .ZN(n37506) );
  NAND3_X2 U11526 ( .A1(n36918), .A2(n37507), .A3(n34881), .ZN(n33038) );
  NAND2_X1 U11530 ( .A1(n18325), .A2(n18326), .ZN(n37507) );
  NAND2_X1 U11537 ( .A1(n29380), .A2(n13302), .ZN(n13942) );
  BUF_X2 U11538 ( .I(n27395), .Z(n37508) );
  INV_X2 U11539 ( .I(n8899), .ZN(n22300) );
  NAND2_X2 U11541 ( .A1(n21), .A2(n4391), .ZN(n8899) );
  NOR2_X2 U11542 ( .A1(n35560), .A2(n32045), .ZN(n24612) );
  NAND2_X2 U11547 ( .A1(n37509), .A2(n34811), .ZN(n2305) );
  NAND2_X2 U11549 ( .A1(n9202), .A2(n1890), .ZN(n37509) );
  XOR2_X1 U11552 ( .A1(n23714), .A2(n2145), .Z(n23725) );
  NOR2_X2 U11553 ( .A1(n33775), .A2(n2086), .ZN(n2145) );
  NAND2_X2 U11554 ( .A1(n39668), .A2(n9941), .ZN(n22298) );
  AOI21_X2 U11556 ( .A1(n28399), .A2(n28755), .B(n37510), .ZN(n28610) );
  AOI21_X2 U11558 ( .A1(n12312), .A2(n12313), .B(n28755), .ZN(n37510) );
  NAND3_X2 U11559 ( .A1(n35963), .A2(n23444), .A3(n4207), .ZN(n2087) );
  XOR2_X1 U11561 ( .A1(n29306), .A2(n28948), .Z(n29257) );
  OAI21_X2 U11562 ( .A1(n27958), .A2(n28490), .B(n27957), .ZN(n29306) );
  XOR2_X1 U11567 ( .A1(n33645), .A2(n26487), .Z(n26370) );
  NAND2_X2 U11569 ( .A1(n39633), .A2(n39822), .ZN(n26487) );
  XOR2_X1 U11570 ( .A1(n23952), .A2(n23775), .Z(n23904) );
  AOI21_X2 U11572 ( .A1(n6052), .A2(n23394), .B(n23393), .ZN(n23952) );
  XOR2_X1 U11573 ( .A1(n37511), .A2(n10478), .Z(n14463) );
  XOR2_X1 U11575 ( .A1(n10887), .A2(n10888), .Z(n37511) );
  AND2_X1 U11581 ( .A1(n15359), .A2(n7696), .Z(n17948) );
  XOR2_X1 U11585 ( .A1(n38054), .A2(n18923), .Z(n34120) );
  NOR2_X2 U11589 ( .A1(n12663), .A2(n16500), .ZN(n39127) );
  INV_X2 U11590 ( .I(n16489), .ZN(n26639) );
  XOR2_X1 U11591 ( .A1(n3995), .A2(n35017), .Z(n16489) );
  NAND2_X2 U11592 ( .A1(n26109), .A2(n13712), .ZN(n16860) );
  XOR2_X1 U11595 ( .A1(n26495), .A2(n11935), .Z(n4205) );
  NAND2_X2 U11598 ( .A1(n38249), .A2(n1647), .ZN(n3813) );
  XNOR2_X1 U11599 ( .A1(n25026), .A2(n18600), .ZN(n25166) );
  XOR2_X1 U11600 ( .A1(n37513), .A2(n4238), .Z(n3229) );
  INV_X1 U11602 ( .I(n17837), .ZN(n37513) );
  XOR2_X1 U11603 ( .A1(n1261), .A2(n15102), .Z(n17837) );
  NAND2_X1 U11605 ( .A1(n1094), .A2(n37054), .ZN(n26858) );
  INV_X1 U11606 ( .I(n25198), .ZN(n37658) );
  NOR2_X2 U11609 ( .A1(n37135), .A2(n37514), .ZN(n38397) );
  NAND2_X2 U11611 ( .A1(n6466), .A2(n31183), .ZN(n22836) );
  OAI22_X2 U11613 ( .A1(n39317), .A2(n37515), .B1(n24547), .B2(n37067), .ZN(
        n19691) );
  NOR2_X2 U11614 ( .A1(n37717), .A2(n11494), .ZN(n32091) );
  NAND2_X1 U11615 ( .A1(n33289), .A2(n12950), .ZN(n24205) );
  NOR2_X2 U11617 ( .A1(n37518), .A2(n37517), .ZN(n37516) );
  NAND3_X2 U11619 ( .A1(n37519), .A2(n19111), .A3(n31583), .ZN(n19109) );
  NAND2_X2 U11625 ( .A1(n38580), .A2(n32720), .ZN(n37519) );
  XOR2_X1 U11626 ( .A1(n17566), .A2(n22449), .Z(n17565) );
  XOR2_X1 U11634 ( .A1(n33736), .A2(n22743), .Z(n22449) );
  OAI21_X1 U11635 ( .A1(n31598), .A2(n967), .B(n10848), .ZN(n10847) );
  XOR2_X1 U11640 ( .A1(n15912), .A2(n25182), .Z(n19072) );
  NAND2_X2 U11641 ( .A1(n18458), .A2(n24652), .ZN(n15912) );
  CLKBUF_X4 U11642 ( .I(n17114), .Z(n37661) );
  OAI22_X2 U11645 ( .A1(n25927), .A2(n2029), .B1(n25928), .B2(n2561), .ZN(
        n26084) );
  AOI22_X2 U11646 ( .A1(n30059), .A2(n30000), .B1(n16353), .B2(n30057), .ZN(
        n32548) );
  XOR2_X1 U11649 ( .A1(n37520), .A2(n710), .Z(n10181) );
  XOR2_X1 U11653 ( .A1(n23671), .A2(n37521), .Z(n37520) );
  INV_X2 U11659 ( .I(n7148), .ZN(n37521) );
  XOR2_X1 U11660 ( .A1(n37874), .A2(n296), .Z(n29043) );
  OAI21_X2 U11666 ( .A1(n28177), .A2(n38311), .B(n35961), .ZN(n296) );
  XOR2_X1 U11670 ( .A1(n4077), .A2(n7101), .Z(n7100) );
  NOR2_X1 U11671 ( .A1(n8599), .A2(n8600), .ZN(n8598) );
  NAND2_X2 U11675 ( .A1(n37522), .A2(n37140), .ZN(n14496) );
  NAND2_X2 U11677 ( .A1(n37604), .A2(n37524), .ZN(n10901) );
  INV_X1 U11678 ( .I(n26885), .ZN(n37524) );
  BUF_X2 U11679 ( .I(n20128), .Z(n37525) );
  AND2_X1 U11680 ( .A1(n23060), .A2(n37922), .Z(n39004) );
  XOR2_X1 U11681 ( .A1(n11752), .A2(n6523), .Z(n8502) );
  OAI21_X2 U11683 ( .A1(n2421), .A2(n4854), .B(n8161), .ZN(n6523) );
  XOR2_X1 U11684 ( .A1(n37526), .A2(n39245), .Z(n34587) );
  XOR2_X1 U11685 ( .A1(n11502), .A2(n27790), .Z(n37526) );
  XOR2_X1 U11687 ( .A1(n37527), .A2(n29168), .Z(n33716) );
  XOR2_X1 U11688 ( .A1(n32073), .A2(n29167), .Z(n37527) );
  AND2_X1 U11689 ( .A1(n19326), .A2(n27131), .Z(n8486) );
  NAND2_X2 U11692 ( .A1(n14216), .A2(n13607), .ZN(n17287) );
  XOR2_X1 U11694 ( .A1(n37529), .A2(n29206), .Z(Ciphertext[4]) );
  NAND2_X1 U11698 ( .A1(n2569), .A2(n36862), .ZN(n37529) );
  INV_X4 U11704 ( .I(n28400), .ZN(n12537) );
  NOR2_X1 U11705 ( .A1(n974), .A2(n28400), .ZN(n36465) );
  XOR2_X1 U11708 ( .A1(n37530), .A2(n23943), .Z(n15860) );
  XOR2_X1 U11711 ( .A1(n39408), .A2(n36461), .Z(n37530) );
  XOR2_X1 U11712 ( .A1(n33473), .A2(n37532), .Z(n9214) );
  XOR2_X1 U11713 ( .A1(n26522), .A2(n26344), .Z(n37532) );
  XOR2_X1 U11714 ( .A1(n37533), .A2(n36040), .Z(Ciphertext[51]) );
  AOI22_X1 U11719 ( .A1(n6340), .A2(n6343), .B1(n6339), .B2(n13433), .ZN(
        n37533) );
  XOR2_X1 U11721 ( .A1(n10214), .A2(n10939), .Z(n36002) );
  NOR2_X2 U11725 ( .A1(n37534), .A2(n12239), .ZN(n39588) );
  NOR3_X2 U11726 ( .A1(n1146), .A2(n8569), .A3(n9699), .ZN(n37534) );
  OAI22_X2 U11729 ( .A1(n1337), .A2(n2709), .B1(n22022), .B2(n32434), .ZN(
        n39455) );
  INV_X2 U11733 ( .I(n22086), .ZN(n1337) );
  OAI21_X2 U11734 ( .A1(n21491), .A2(n3670), .B(n38091), .ZN(n22086) );
  XOR2_X1 U11735 ( .A1(n31568), .A2(n37038), .Z(n15978) );
  NOR2_X2 U11736 ( .A1(n15525), .A2(n15526), .ZN(n37038) );
  NAND4_X1 U11737 ( .A1(n29472), .A2(n29473), .A3(n29469), .A4(n29470), .ZN(
        n6342) );
  XOR2_X1 U11744 ( .A1(n10794), .A2(n29833), .Z(n32200) );
  AOI22_X2 U11746 ( .A1(n7869), .A2(n28539), .B1(n4228), .B2(n28538), .ZN(
        n10794) );
  NAND2_X2 U11753 ( .A1(n5304), .A2(n5303), .ZN(n38976) );
  AOI22_X2 U11754 ( .A1(n5551), .A2(n5132), .B1(n21916), .B2(n5391), .ZN(n5304) );
  XOR2_X1 U11759 ( .A1(n26569), .A2(n26466), .Z(n26313) );
  XOR2_X1 U11761 ( .A1(n26421), .A2(n20600), .Z(n26466) );
  NAND2_X2 U11764 ( .A1(n17826), .A2(n32797), .ZN(n38466) );
  NOR2_X2 U11766 ( .A1(n37535), .A2(n9233), .ZN(n36889) );
  AOI21_X2 U11768 ( .A1(n29993), .A2(n4095), .B(n3693), .ZN(n37535) );
  OAI22_X2 U11771 ( .A1(n37536), .A2(n3363), .B1(n23525), .B2(n36103), .ZN(
        n18540) );
  NAND2_X2 U11775 ( .A1(n3366), .A2(n30835), .ZN(n37536) );
  OAI21_X2 U11776 ( .A1(n37538), .A2(n31845), .B(n37537), .ZN(n23859) );
  NOR2_X2 U11777 ( .A1(n957), .A2(n38777), .ZN(n37538) );
  NAND2_X2 U11779 ( .A1(n37541), .A2(n16121), .ZN(n15841) );
  NAND2_X1 U11782 ( .A1(n36968), .A2(n16252), .ZN(n37541) );
  NAND2_X2 U11783 ( .A1(n3862), .A2(n19288), .ZN(n17928) );
  OAI22_X2 U11791 ( .A1(n14817), .A2(n22993), .B1(n22929), .B2(n20449), .ZN(
        n3862) );
  NAND2_X2 U11793 ( .A1(n30107), .A2(n35187), .ZN(n30112) );
  NAND2_X2 U11802 ( .A1(n33070), .A2(n4073), .ZN(n30107) );
  XOR2_X1 U11804 ( .A1(n26155), .A2(n26503), .Z(n17171) );
  OR2_X1 U11812 ( .A1(n875), .A2(n26934), .Z(n34918) );
  AOI21_X1 U11813 ( .A1(n9512), .A2(n30986), .B(n9454), .ZN(n37760) );
  INV_X2 U11815 ( .I(n8050), .ZN(n451) );
  NAND2_X2 U11816 ( .A1(n14278), .A2(n11956), .ZN(n8050) );
  NAND2_X2 U11818 ( .A1(n28344), .A2(n28346), .ZN(n28716) );
  NOR2_X2 U11822 ( .A1(n24328), .A2(n1607), .ZN(n6585) );
  NAND2_X2 U11826 ( .A1(n39664), .A2(n37460), .ZN(n16921) );
  NAND2_X2 U11829 ( .A1(n27346), .A2(n27345), .ZN(n9185) );
  OAI21_X2 U11835 ( .A1(n4668), .A2(n5027), .B(n4667), .ZN(n27346) );
  AOI22_X2 U11839 ( .A1(n3708), .A2(n23523), .B1(n34959), .B2(n5258), .ZN(
        n23589) );
  NAND2_X2 U11841 ( .A1(n35361), .A2(n30815), .ZN(n3708) );
  XOR2_X1 U11844 ( .A1(n26462), .A2(n19973), .Z(n10113) );
  XOR2_X1 U11847 ( .A1(n1505), .A2(n12649), .Z(n26462) );
  XOR2_X1 U11849 ( .A1(n3501), .A2(n27745), .Z(n14977) );
  XOR2_X1 U11852 ( .A1(n37542), .A2(n25185), .Z(n10926) );
  XOR2_X1 U11855 ( .A1(n25184), .A2(n39146), .Z(n37542) );
  XOR2_X1 U11858 ( .A1(n10100), .A2(n1614), .Z(n39344) );
  NAND2_X1 U11860 ( .A1(n15919), .A2(n32690), .ZN(n38866) );
  INV_X2 U11862 ( .I(n11219), .ZN(n39126) );
  NAND3_X2 U11865 ( .A1(n38734), .A2(n34535), .A3(n27398), .ZN(n35243) );
  NAND2_X2 U11869 ( .A1(n10856), .A2(n37543), .ZN(n29050) );
  AOI22_X2 U11873 ( .A1(n38275), .A2(n18996), .B1(n36663), .B2(n36076), .ZN(
        n37543) );
  NAND2_X2 U11874 ( .A1(n37545), .A2(n37544), .ZN(n37915) );
  INV_X2 U11877 ( .I(n777), .ZN(n37544) );
  XOR2_X1 U11878 ( .A1(n11250), .A2(n37546), .Z(n32474) );
  XOR2_X1 U11890 ( .A1(n27812), .A2(n27813), .Z(n37546) );
  NAND2_X1 U11893 ( .A1(n20923), .A2(n12754), .ZN(n21606) );
  NAND2_X2 U11895 ( .A1(n37548), .A2(n37547), .ZN(n36810) );
  OAI21_X2 U11897 ( .A1(n22869), .A2(n22870), .B(n16963), .ZN(n37547) );
  XOR2_X1 U11901 ( .A1(n26205), .A2(n26462), .Z(n3780) );
  AOI21_X2 U11904 ( .A1(n14146), .A2(n10290), .B(n13677), .ZN(n14145) );
  NOR2_X2 U11906 ( .A1(n1014), .A2(n31205), .ZN(n10290) );
  AND2_X1 U11910 ( .A1(n23493), .A2(n34603), .Z(n37906) );
  NOR2_X1 U11911 ( .A1(n9452), .A2(n37760), .ZN(n9513) );
  NOR2_X1 U11912 ( .A1(n12331), .A2(n22929), .ZN(n22991) );
  INV_X2 U11916 ( .I(n12100), .ZN(n12331) );
  XOR2_X1 U11917 ( .A1(n12102), .A2(n9595), .Z(n12100) );
  NAND2_X1 U11919 ( .A1(n37557), .A2(n28503), .ZN(n37556) );
  NOR2_X2 U11920 ( .A1(n36912), .A2(n39426), .ZN(n37550) );
  NOR2_X2 U11921 ( .A1(n35781), .A2(n37551), .ZN(n38478) );
  AND2_X1 U11926 ( .A1(n25882), .A2(n840), .Z(n31471) );
  XOR2_X1 U11927 ( .A1(n38022), .A2(n5841), .Z(n23807) );
  NAND2_X2 U11928 ( .A1(n37625), .A2(n10853), .ZN(n9875) );
  OR2_X1 U11930 ( .A1(n39417), .A2(n39628), .Z(n36984) );
  NAND3_X2 U11933 ( .A1(n17191), .A2(n28756), .A3(n28398), .ZN(n17190) );
  INV_X1 U11934 ( .I(n14369), .ZN(n1552) );
  AND2_X2 U11936 ( .A1(n14369), .A2(n37553), .Z(n25603) );
  XOR2_X1 U11942 ( .A1(n8713), .A2(n31075), .Z(n14369) );
  OAI21_X1 U11943 ( .A1(n17369), .A2(n29662), .B(n29660), .ZN(n32290) );
  INV_X1 U11945 ( .I(n29641), .ZN(n17369) );
  AOI22_X2 U11947 ( .A1(n29638), .A2(n29761), .B1(n29637), .B2(n1178), .ZN(
        n29641) );
  XOR2_X1 U11948 ( .A1(n9939), .A2(n15592), .Z(n7076) );
  XOR2_X1 U11949 ( .A1(n589), .A2(n14835), .Z(n14834) );
  XOR2_X1 U11954 ( .A1(n3342), .A2(n34375), .Z(n589) );
  XOR2_X1 U11955 ( .A1(n37554), .A2(n14147), .Z(n13091) );
  XOR2_X1 U11959 ( .A1(n27790), .A2(n39410), .Z(n37554) );
  XOR2_X1 U11962 ( .A1(n26356), .A2(n26357), .Z(n20082) );
  NAND2_X2 U11970 ( .A1(n1849), .A2(n1850), .ZN(n26356) );
  AND2_X1 U11971 ( .A1(n6056), .A2(n4382), .Z(n25792) );
  OAI22_X2 U11973 ( .A1(n37555), .A2(n6698), .B1(n6697), .B2(n28178), .ZN(
        n28966) );
  NAND2_X2 U11980 ( .A1(n6684), .A2(n1637), .ZN(n9346) );
  XOR2_X1 U11981 ( .A1(n25280), .A2(n6185), .Z(n10582) );
  AOI21_X2 U11982 ( .A1(n20505), .A2(n3630), .B(n3629), .ZN(n25280) );
  XOR2_X1 U11983 ( .A1(n36366), .A2(n26502), .Z(n26512) );
  OAI22_X2 U11984 ( .A1(n38084), .A2(n13891), .B1(n37558), .B2(n37556), .ZN(
        n29041) );
  NAND2_X2 U11988 ( .A1(n36798), .A2(n598), .ZN(n25822) );
  AOI22_X2 U11990 ( .A1(n12931), .A2(n9439), .B1(n9440), .B2(n38338), .ZN(n598) );
  NOR2_X2 U11992 ( .A1(n4941), .A2(n30837), .ZN(n28503) );
  NAND2_X2 U11995 ( .A1(n18131), .A2(n31087), .ZN(n4941) );
  NAND2_X1 U12003 ( .A1(n12675), .A2(n13811), .ZN(n38959) );
  AND2_X2 U12006 ( .A1(n18342), .A2(n24271), .Z(n18698) );
  NOR2_X2 U12009 ( .A1(n2522), .A2(n1081), .ZN(n2519) );
  NOR2_X2 U12015 ( .A1(n12081), .A2(n19544), .ZN(n39393) );
  NAND2_X2 U12016 ( .A1(n37788), .A2(n37562), .ZN(n27438) );
  NAND2_X2 U12022 ( .A1(n34820), .A2(n37563), .ZN(n8966) );
  OAI21_X2 U12024 ( .A1(n30944), .A2(n31490), .B(n305), .ZN(n37563) );
  XOR2_X1 U12026 ( .A1(n26246), .A2(n26245), .Z(n26324) );
  NOR2_X2 U12027 ( .A1(n4884), .A2(n25531), .ZN(n26246) );
  NAND3_X2 U12028 ( .A1(n37028), .A2(n25916), .A3(n1016), .ZN(n25917) );
  BUF_X2 U12029 ( .I(n3937), .Z(n4001) );
  OAI21_X1 U12032 ( .A1(n25644), .A2(n25666), .B(n4468), .ZN(n4466) );
  OR2_X1 U12034 ( .A1(n5062), .A2(n28197), .Z(n33804) );
  OR2_X1 U12036 ( .A1(n12924), .A2(n36396), .Z(n18997) );
  XOR2_X1 U12037 ( .A1(n29829), .A2(n29081), .Z(n28893) );
  OAI21_X2 U12038 ( .A1(n27033), .A2(n37205), .B(n27032), .ZN(n27774) );
  NAND2_X1 U12042 ( .A1(n35380), .A2(n4700), .ZN(n37657) );
  OAI21_X2 U12046 ( .A1(n299), .A2(n17613), .B(n20381), .ZN(n35903) );
  XOR2_X1 U12051 ( .A1(n37564), .A2(n19498), .Z(Ciphertext[100]) );
  NAND2_X1 U12053 ( .A1(n29749), .A2(n31477), .ZN(n37564) );
  NAND2_X1 U12054 ( .A1(n32802), .A2(n24900), .ZN(n17475) );
  NAND2_X1 U12059 ( .A1(n29632), .A2(n1398), .ZN(n37565) );
  XOR2_X1 U12064 ( .A1(n26141), .A2(n21086), .Z(n34966) );
  OAI21_X2 U12065 ( .A1(n3044), .A2(n38073), .B(n37566), .ZN(n35925) );
  NAND3_X2 U12066 ( .A1(n37737), .A2(n39279), .A3(n34011), .ZN(n37566) );
  NAND3_X2 U12067 ( .A1(n19400), .A2(n39389), .A3(n37051), .ZN(n13535) );
  NAND2_X1 U12069 ( .A1(n36177), .A2(n9267), .ZN(n38788) );
  XOR2_X1 U12079 ( .A1(n37567), .A2(n31062), .Z(Ciphertext[62]) );
  NAND3_X2 U12083 ( .A1(n28905), .A2(n28906), .A3(n28907), .ZN(n37567) );
  XOR2_X1 U12085 ( .A1(n35062), .A2(n23930), .Z(n23787) );
  NOR2_X1 U12086 ( .A1(n14278), .A2(n11956), .ZN(n34567) );
  OAI21_X2 U12089 ( .A1(n6160), .A2(n31275), .B(n31785), .ZN(n11956) );
  NAND2_X2 U12093 ( .A1(n4579), .A2(n4580), .ZN(n15135) );
  XOR2_X1 U12099 ( .A1(n37568), .A2(n34017), .Z(Ciphertext[11]) );
  AOI22_X1 U12100 ( .A1(n29226), .A2(n35264), .B1(n1378), .B2(n12691), .ZN(
        n37568) );
  XOR2_X1 U12121 ( .A1(n9874), .A2(n22572), .Z(n22625) );
  XOR2_X1 U12125 ( .A1(n33194), .A2(n26548), .Z(n26408) );
  NAND2_X2 U12129 ( .A1(n25984), .A2(n25983), .ZN(n26548) );
  XOR2_X1 U12130 ( .A1(n6559), .A2(n6560), .Z(n23785) );
  OAI21_X2 U12134 ( .A1(n37569), .A2(n17674), .B(n10763), .ZN(n17673) );
  XOR2_X1 U12140 ( .A1(n37038), .A2(n31181), .Z(n25180) );
  NAND2_X2 U12141 ( .A1(n37570), .A2(n19702), .ZN(n38713) );
  AOI21_X2 U12143 ( .A1(n25527), .A2(n19701), .B(n1539), .ZN(n37570) );
  NOR2_X1 U12148 ( .A1(n33266), .A2(n39026), .ZN(n38257) );
  NOR2_X2 U12150 ( .A1(n3190), .A2(n7950), .ZN(n3441) );
  XOR2_X1 U12151 ( .A1(n1260), .A2(n12297), .Z(n12296) );
  AOI22_X2 U12161 ( .A1(n24701), .A2(n6791), .B1(n24270), .B2(n24530), .ZN(
        n25259) );
  XOR2_X1 U12163 ( .A1(n29096), .A2(n37571), .Z(n12157) );
  INV_X2 U12168 ( .I(n14956), .ZN(n37571) );
  OAI21_X2 U12169 ( .A1(n37572), .A2(n23372), .B(n38623), .ZN(n13395) );
  OAI21_X2 U12173 ( .A1(n34386), .A2(n32061), .B(n37573), .ZN(n37572) );
  NAND2_X2 U12174 ( .A1(n34386), .A2(n23370), .ZN(n37573) );
  NOR2_X1 U12177 ( .A1(n13432), .A2(n13431), .ZN(n37620) );
  XOR2_X1 U12179 ( .A1(n16805), .A2(n37574), .Z(n32822) );
  XOR2_X1 U12180 ( .A1(n37860), .A2(n767), .Z(n37574) );
  NOR2_X2 U12182 ( .A1(n11470), .A2(n11208), .ZN(n18960) );
  NAND3_X2 U12186 ( .A1(n9303), .A2(n25756), .A3(n12931), .ZN(n37949) );
  XOR2_X1 U12188 ( .A1(n25324), .A2(n24931), .Z(n24946) );
  NAND2_X2 U12190 ( .A1(n19356), .A2(n24706), .ZN(n25324) );
  NAND2_X2 U12193 ( .A1(n37575), .A2(n7488), .ZN(n32691) );
  NOR2_X2 U12196 ( .A1(n36302), .A2(n19927), .ZN(n37575) );
  XOR2_X1 U12209 ( .A1(n38455), .A2(n11402), .Z(n3785) );
  XOR2_X1 U12211 ( .A1(n27483), .A2(n27535), .Z(n36628) );
  NAND2_X2 U12212 ( .A1(n29895), .A2(n37576), .ZN(n19097) );
  OAI21_X2 U12213 ( .A1(n32498), .A2(n32499), .B(n17240), .ZN(n37576) );
  NOR2_X1 U12217 ( .A1(n30747), .A2(n1178), .ZN(n15376) );
  BUF_X4 U12219 ( .I(n25324), .Z(n37943) );
  XOR2_X1 U12221 ( .A1(n18498), .A2(n27865), .Z(n33642) );
  XOR2_X1 U12229 ( .A1(n27737), .A2(n27736), .Z(n27865) );
  AOI21_X2 U12230 ( .A1(n37578), .A2(n37577), .B(n14652), .ZN(n28896) );
  NOR2_X2 U12231 ( .A1(n28438), .A2(n37579), .ZN(n37578) );
  NAND2_X2 U12232 ( .A1(n35123), .A2(n38078), .ZN(n38816) );
  XOR2_X1 U12233 ( .A1(n27722), .A2(n27721), .Z(n36603) );
  XOR2_X1 U12237 ( .A1(n27593), .A2(n27703), .Z(n27722) );
  OAI21_X2 U12238 ( .A1(n1011), .A2(n1243), .B(n30629), .ZN(n11980) );
  OAI21_X2 U12247 ( .A1(n13534), .A2(n13533), .B(n12705), .ZN(n30629) );
  XOR2_X1 U12249 ( .A1(n27777), .A2(n27511), .Z(n608) );
  NAND2_X2 U12254 ( .A1(n27052), .A2(n27051), .ZN(n27777) );
  NAND2_X1 U12258 ( .A1(n8820), .A2(n8822), .ZN(n11514) );
  NAND2_X2 U12262 ( .A1(n17231), .A2(n17232), .ZN(n25801) );
  OAI21_X2 U12264 ( .A1(n36344), .A2(n26857), .B(n1491), .ZN(n34985) );
  XOR2_X1 U12266 ( .A1(n33578), .A2(n2222), .Z(n6226) );
  NAND2_X2 U12268 ( .A1(n19636), .A2(n19637), .ZN(n25387) );
  NAND2_X2 U12270 ( .A1(n11496), .A2(n24741), .ZN(n19636) );
  XOR2_X1 U12272 ( .A1(n1184), .A2(n14941), .Z(n29126) );
  BUF_X4 U12273 ( .I(n15988), .Z(n1006) );
  NOR2_X2 U12276 ( .A1(n37581), .A2(n6423), .ZN(n23310) );
  NOR2_X2 U12278 ( .A1(n16416), .A2(n23013), .ZN(n37581) );
  BUF_X2 U12280 ( .I(n36571), .Z(n37582) );
  NAND2_X2 U12281 ( .A1(n37583), .A2(n6509), .ZN(n7565) );
  NOR2_X2 U12283 ( .A1(n18698), .A2(n37264), .ZN(n37583) );
  XOR2_X1 U12284 ( .A1(n25016), .A2(n35900), .Z(n9939) );
  NAND2_X2 U12288 ( .A1(n8108), .A2(n11738), .ZN(n25016) );
  BUF_X2 U12291 ( .I(n19728), .Z(n37585) );
  NOR2_X2 U12297 ( .A1(n29468), .A2(n9105), .ZN(n12369) );
  NOR2_X2 U12299 ( .A1(n39060), .A2(n8924), .ZN(n29468) );
  OAI21_X2 U12301 ( .A1(n12167), .A2(n29644), .B(n37586), .ZN(n10030) );
  NAND2_X2 U12305 ( .A1(n37743), .A2(n29645), .ZN(n37586) );
  INV_X2 U12312 ( .I(n37587), .ZN(n35233) );
  XOR2_X1 U12315 ( .A1(n9555), .A2(n6455), .Z(n37588) );
  XOR2_X1 U12319 ( .A1(n10498), .A2(n8793), .Z(n9266) );
  AOI22_X2 U12322 ( .A1(n10901), .A2(n10903), .B1(n39302), .B2(n10902), .ZN(
        n37625) );
  XOR2_X1 U12325 ( .A1(n17757), .A2(n26463), .Z(n12145) );
  NOR3_X2 U12326 ( .A1(n13440), .A2(n18314), .A3(n17297), .ZN(n26463) );
  NOR2_X2 U12327 ( .A1(n37591), .A2(n37590), .ZN(n38965) );
  NAND3_X1 U12328 ( .A1(n16633), .A2(n4410), .A3(n37235), .ZN(n37592) );
  AND2_X1 U12330 ( .A1(n26642), .A2(n26644), .Z(n39179) );
  NAND2_X2 U12334 ( .A1(n9694), .A2(n26031), .ZN(n25915) );
  NAND2_X2 U12338 ( .A1(n34260), .A2(n25605), .ZN(n9694) );
  AOI21_X2 U12339 ( .A1(n31516), .A2(n30747), .B(n19599), .ZN(n30746) );
  NOR2_X1 U12341 ( .A1(n9893), .A2(n14369), .ZN(n12616) );
  XOR2_X1 U12342 ( .A1(n25102), .A2(n10611), .Z(n37998) );
  NOR2_X2 U12348 ( .A1(n3509), .A2(n36450), .ZN(n2561) );
  NAND2_X2 U12351 ( .A1(n7466), .A2(n39380), .ZN(n3509) );
  NAND2_X2 U12353 ( .A1(n167), .A2(n19425), .ZN(n26943) );
  INV_X2 U12354 ( .I(n35176), .ZN(n19272) );
  XOR2_X1 U12357 ( .A1(n37594), .A2(n37639), .Z(n39750) );
  XOR2_X1 U12359 ( .A1(n33587), .A2(n27556), .Z(n37594) );
  INV_X2 U12361 ( .I(n5745), .ZN(n11083) );
  OR2_X1 U12362 ( .A1(n17119), .A2(n39810), .Z(n17128) );
  OR2_X1 U12364 ( .A1(n18682), .A2(n16528), .Z(n18478) );
  XOR2_X1 U12367 ( .A1(n37595), .A2(n1371), .Z(Ciphertext[112]) );
  NOR3_X1 U12369 ( .A1(n36410), .A2(n36365), .A3(n6650), .ZN(n37595) );
  NAND2_X2 U12372 ( .A1(n12178), .A2(n20845), .ZN(n28500) );
  OR2_X1 U12375 ( .A1(n12682), .A2(n3873), .Z(n26859) );
  XOR2_X1 U12381 ( .A1(n26486), .A2(n10668), .Z(n3732) );
  XOR2_X1 U12382 ( .A1(n26542), .A2(n35214), .Z(n26486) );
  OAI21_X2 U12384 ( .A1(n3631), .A2(n3699), .B(n3698), .ZN(n28924) );
  NAND2_X2 U12391 ( .A1(n37596), .A2(n30372), .ZN(n31362) );
  XOR2_X1 U12392 ( .A1(n11116), .A2(n15202), .Z(n11115) );
  XOR2_X1 U12394 ( .A1(n25166), .A2(n25007), .Z(n3495) );
  INV_X2 U12401 ( .I(n18870), .ZN(n17346) );
  NOR2_X1 U12403 ( .A1(n35881), .A2(n5392), .ZN(n21916) );
  NAND2_X2 U12418 ( .A1(n37597), .A2(n12249), .ZN(n14283) );
  NAND2_X2 U12419 ( .A1(n37967), .A2(n1127), .ZN(n37597) );
  OR2_X1 U12422 ( .A1(n38976), .A2(n30800), .Z(n20756) );
  BUF_X2 U12424 ( .I(n34977), .Z(n37598) );
  NAND2_X2 U12429 ( .A1(n19340), .A2(n37599), .ZN(n25924) );
  NAND2_X2 U12435 ( .A1(n25803), .A2(n16407), .ZN(n37599) );
  XOR2_X1 U12437 ( .A1(n37600), .A2(n20819), .Z(n29196) );
  XOR2_X1 U12440 ( .A1(n28502), .A2(n29105), .Z(n37600) );
  INV_X2 U12441 ( .I(n29626), .ZN(n29618) );
  NAND3_X2 U12442 ( .A1(n34097), .A2(n8996), .A3(n8999), .ZN(n29626) );
  NAND2_X2 U12448 ( .A1(n36986), .A2(n2774), .ZN(n34599) );
  NAND2_X2 U12450 ( .A1(n37601), .A2(n24167), .ZN(n10980) );
  XOR2_X1 U12456 ( .A1(n10215), .A2(n21253), .Z(n8923) );
  AOI22_X2 U12467 ( .A1(n29557), .A2(n29558), .B1(n29559), .B2(n29560), .ZN(
        n21158) );
  XOR2_X1 U12468 ( .A1(n28835), .A2(n29816), .Z(n10899) );
  XOR2_X1 U12469 ( .A1(n36928), .A2(n296), .Z(n28835) );
  XOR2_X1 U12471 ( .A1(n23732), .A2(n714), .Z(n37834) );
  XOR2_X1 U12474 ( .A1(n23888), .A2(n23886), .Z(n23732) );
  INV_X2 U12475 ( .I(n29124), .ZN(n38610) );
  NAND2_X2 U12478 ( .A1(n37759), .A2(n36313), .ZN(n29124) );
  NOR2_X2 U12481 ( .A1(n10171), .A2(n15135), .ZN(n26791) );
  XOR2_X1 U12483 ( .A1(n26441), .A2(n4622), .Z(n26254) );
  NOR2_X2 U12484 ( .A1(n34413), .A2(n11010), .ZN(n26441) );
  XOR2_X1 U12485 ( .A1(n37602), .A2(n26374), .Z(n26272) );
  XOR2_X1 U12488 ( .A1(n32442), .A2(n13814), .Z(n37602) );
  OR2_X2 U12490 ( .A1(n2616), .A2(n17351), .Z(n7267) );
  OAI21_X2 U12493 ( .A1(n27026), .A2(n27174), .B(n37603), .ZN(n7808) );
  AND2_X1 U12495 ( .A1(n5392), .A2(n21912), .Z(n21913) );
  OAI22_X1 U12497 ( .A1(n30110), .A2(n10118), .B1(n30111), .B2(n30112), .ZN(
        n39578) );
  OAI22_X2 U12498 ( .A1(n37604), .A2(n12066), .B1(n12065), .B2(n2140), .ZN(
        n7861) );
  BUF_X4 U12499 ( .I(n15579), .Z(n34386) );
  OR3_X1 U12503 ( .A1(n27969), .A2(n14451), .A3(n19366), .Z(n20919) );
  XOR2_X1 U12512 ( .A1(n7061), .A2(n7059), .Z(n19764) );
  XOR2_X1 U12513 ( .A1(n27842), .A2(n27754), .Z(n27524) );
  NOR2_X2 U12514 ( .A1(n27060), .A2(n27061), .ZN(n27842) );
  NAND3_X1 U12515 ( .A1(n28498), .A2(n33591), .A3(n28497), .ZN(n12178) );
  NAND2_X2 U12529 ( .A1(n35491), .A2(n1882), .ZN(n28498) );
  NOR2_X2 U12530 ( .A1(n37607), .A2(n37606), .ZN(n20454) );
  OAI22_X2 U12536 ( .A1(n19276), .A2(n7676), .B1(n27118), .B2(n32976), .ZN(
        n37606) );
  AOI21_X1 U12538 ( .A1(n20455), .A2(n27006), .B(n35184), .ZN(n37607) );
  XOR2_X1 U12543 ( .A1(n8474), .A2(n28988), .Z(n10541) );
  XOR2_X1 U12544 ( .A1(n31615), .A2(n28500), .Z(n28988) );
  NAND2_X2 U12545 ( .A1(n26657), .A2(n37608), .ZN(n7975) );
  AOI22_X2 U12553 ( .A1(n13645), .A2(n26701), .B1(n13644), .B2(n36244), .ZN(
        n37608) );
  XOR2_X1 U12558 ( .A1(n10153), .A2(n37609), .Z(n7980) );
  XOR2_X1 U12560 ( .A1(n33812), .A2(n38209), .Z(n37609) );
  XOR2_X1 U12562 ( .A1(n10792), .A2(n16900), .Z(n25251) );
  AOI22_X2 U12573 ( .A1(n35180), .A2(n29525), .B1(n29527), .B2(n29531), .ZN(
        n29536) );
  AOI21_X2 U12574 ( .A1(n14780), .A2(n24275), .B(n364), .ZN(n2616) );
  NAND2_X2 U12576 ( .A1(n39250), .A2(n10321), .ZN(n26097) );
  XOR2_X1 U12578 ( .A1(n5609), .A2(n37610), .Z(n5732) );
  XOR2_X1 U12579 ( .A1(n17910), .A2(n3734), .Z(n37610) );
  XOR2_X1 U12580 ( .A1(n37611), .A2(n39103), .Z(n13429) );
  XOR2_X1 U12581 ( .A1(n5913), .A2(n5915), .Z(n37611) );
  BUF_X2 U12582 ( .I(n7935), .Z(n37612) );
  XOR2_X1 U12584 ( .A1(n22774), .A2(n22494), .Z(n387) );
  XOR2_X1 U12585 ( .A1(n22600), .A2(n13704), .Z(n22774) );
  XOR2_X1 U12588 ( .A1(n12069), .A2(n13800), .Z(n39171) );
  NAND3_X2 U12595 ( .A1(n3221), .A2(n11465), .A3(n16791), .ZN(n29289) );
  XOR2_X1 U12597 ( .A1(n36743), .A2(n26184), .Z(n32339) );
  XOR2_X1 U12601 ( .A1(n17048), .A2(n26567), .Z(n26184) );
  AND2_X1 U12606 ( .A1(n32284), .A2(n35777), .Z(n37615) );
  OAI22_X2 U12607 ( .A1(n29541), .A2(n1394), .B1(n29546), .B2(n29558), .ZN(
        n29560) );
  NAND2_X2 U12619 ( .A1(n37645), .A2(n37616), .ZN(n25971) );
  XOR2_X1 U12621 ( .A1(n18975), .A2(n26386), .Z(n18974) );
  XOR2_X1 U12628 ( .A1(n26511), .A2(n26224), .Z(n26386) );
  INV_X2 U12631 ( .I(n20877), .ZN(n24017) );
  XOR2_X1 U12635 ( .A1(n23778), .A2(n37617), .Z(n20877) );
  INV_X2 U12636 ( .I(n23899), .ZN(n37617) );
  XOR2_X1 U12640 ( .A1(n8303), .A2(n28886), .Z(n29151) );
  OAI21_X2 U12641 ( .A1(n21026), .A2(n28298), .B(n21024), .ZN(n8303) );
  XOR2_X1 U12646 ( .A1(n31524), .A2(n31127), .Z(n38772) );
  NAND2_X2 U12647 ( .A1(n32758), .A2(n11719), .ZN(n31524) );
  OR2_X2 U12654 ( .A1(n10111), .A2(n20891), .Z(n26926) );
  XOR2_X1 U12655 ( .A1(n16647), .A2(n9590), .Z(n39443) );
  NAND3_X2 U12657 ( .A1(n18352), .A2(n37618), .A3(n18353), .ZN(n33645) );
  NAND2_X2 U12658 ( .A1(n37619), .A2(n12537), .ZN(n34171) );
  INV_X2 U12659 ( .I(n32146), .ZN(n37619) );
  XOR2_X1 U12663 ( .A1(n37620), .A2(n33184), .Z(Ciphertext[48]) );
  OAI22_X2 U12667 ( .A1(n17066), .A2(n24383), .B1(n18907), .B2(n18402), .ZN(
        n20795) );
  OAI21_X2 U12669 ( .A1(n30357), .A2(n15389), .B(n37621), .ZN(n28245) );
  NAND2_X2 U12671 ( .A1(n15389), .A2(n28240), .ZN(n37621) );
  NOR2_X1 U12673 ( .A1(n39554), .A2(n18668), .ZN(n19034) );
  BUF_X2 U12675 ( .I(n28159), .Z(n37623) );
  XOR2_X1 U12680 ( .A1(n4999), .A2(n5646), .Z(n11543) );
  XOR2_X1 U12685 ( .A1(n17563), .A2(n8113), .Z(n6403) );
  OAI22_X2 U12688 ( .A1(n27057), .A2(n27368), .B1(n27056), .B2(n33050), .ZN(
        n27511) );
  NOR2_X1 U12689 ( .A1(n31788), .A2(n30154), .ZN(n34065) );
  AOI21_X2 U12690 ( .A1(n28149), .A2(n27622), .B(n17753), .ZN(n37626) );
  NAND2_X2 U12698 ( .A1(n21144), .A2(n27276), .ZN(n27059) );
  XOR2_X1 U12703 ( .A1(n27645), .A2(n27494), .Z(n10498) );
  XOR2_X1 U12704 ( .A1(n14808), .A2(n10997), .Z(n27645) );
  INV_X2 U12713 ( .I(n11126), .ZN(n37624) );
  NAND2_X2 U12717 ( .A1(n13179), .A2(n37626), .ZN(n8743) );
  XOR2_X1 U12718 ( .A1(n12865), .A2(n37627), .Z(n5291) );
  XOR2_X1 U12719 ( .A1(n16857), .A2(n33587), .Z(n37627) );
  NOR3_X1 U12720 ( .A1(n15004), .A2(n8493), .A3(n19604), .ZN(n31369) );
  NOR2_X2 U12721 ( .A1(n19454), .A2(n37628), .ZN(n34378) );
  OAI22_X1 U12724 ( .A1(n6692), .A2(n8529), .B1(n29937), .B2(n29935), .ZN(
        n37628) );
  OR2_X1 U12725 ( .A1(n3873), .A2(n14415), .Z(n5263) );
  XOR2_X1 U12727 ( .A1(n34812), .A2(n27554), .Z(n11236) );
  NAND2_X2 U12729 ( .A1(n2303), .A2(n2305), .ZN(n27554) );
  NAND2_X1 U12732 ( .A1(n34008), .A2(n27932), .ZN(n8056) );
  NAND3_X2 U12737 ( .A1(n37630), .A2(n11455), .A3(n11456), .ZN(n22740) );
  NAND2_X1 U12739 ( .A1(n3137), .A2(n11234), .ZN(n37630) );
  XOR2_X1 U12743 ( .A1(n37631), .A2(n39071), .Z(n13540) );
  XOR2_X1 U12745 ( .A1(n3932), .A2(n8884), .Z(n37631) );
  INV_X2 U12748 ( .I(n3937), .ZN(n20441) );
  NAND2_X2 U12750 ( .A1(n37633), .A2(n8289), .ZN(n31663) );
  OAI21_X2 U12753 ( .A1(n33020), .A2(n33981), .B(n28265), .ZN(n37633) );
  AOI22_X2 U12755 ( .A1(n9068), .A2(n24297), .B1(n12248), .B2(n37634), .ZN(
        n19499) );
  NAND3_X2 U12759 ( .A1(n37635), .A2(n4360), .A3(n4361), .ZN(n15266) );
  INV_X4 U12762 ( .I(n19771), .ZN(n28742) );
  NAND2_X2 U12764 ( .A1(n34965), .A2(n406), .ZN(n19771) );
  NAND3_X2 U12765 ( .A1(n20994), .A2(n30231), .A3(n37636), .ZN(n30249) );
  XOR2_X1 U12766 ( .A1(n37899), .A2(n17850), .Z(n17518) );
  OAI21_X1 U12767 ( .A1(n36649), .A2(n38830), .B(n37805), .ZN(n38832) );
  NAND2_X1 U12768 ( .A1(n38832), .A2(n38746), .ZN(n9734) );
  XNOR2_X1 U12770 ( .A1(n27703), .A2(n27595), .ZN(n27831) );
  NAND2_X2 U12773 ( .A1(n8601), .A2(n13792), .ZN(n27595) );
  OAI22_X2 U12774 ( .A1(n2338), .A2(n37671), .B1(n3235), .B2(n39298), .ZN(
        n6160) );
  NAND3_X1 U12777 ( .A1(n2803), .A2(n25484), .A3(n3985), .ZN(n36459) );
  XOR2_X1 U12778 ( .A1(n28967), .A2(n9035), .Z(n37973) );
  NOR2_X2 U12782 ( .A1(n37638), .A2(n37637), .ZN(n28967) );
  INV_X2 U12785 ( .I(n17132), .ZN(n38060) );
  NAND2_X2 U12787 ( .A1(n7914), .A2(n28547), .ZN(n35326) );
  NAND2_X2 U12788 ( .A1(n7251), .A2(n11956), .ZN(n7914) );
  BUF_X2 U12790 ( .I(n14415), .Z(n278) );
  INV_X2 U12791 ( .I(n35657), .ZN(n2870) );
  NAND2_X1 U12792 ( .A1(n12869), .A2(n12552), .ZN(n34826) );
  AOI21_X2 U12794 ( .A1(n5365), .A2(n7612), .B(n36407), .ZN(n31702) );
  INV_X1 U12798 ( .I(n27390), .ZN(n37641) );
  NOR2_X1 U12800 ( .A1(n30358), .A2(n37641), .ZN(n38146) );
  BUF_X2 U12802 ( .I(n38742), .Z(n37643) );
  OAI22_X2 U12803 ( .A1(n6691), .A2(n23060), .B1(n37629), .B2(n22925), .ZN(
        n14743) );
  XOR2_X1 U12805 ( .A1(n37644), .A2(n30170), .Z(Ciphertext[175]) );
  NOR2_X2 U12806 ( .A1(n38029), .A2(n7339), .ZN(n37645) );
  XOR2_X1 U12810 ( .A1(n8505), .A2(n37646), .Z(n9945) );
  XOR2_X1 U12811 ( .A1(n33248), .A2(n24055), .Z(n37646) );
  NAND2_X2 U12812 ( .A1(n25667), .A2(n37647), .ZN(n25936) );
  INV_X2 U12814 ( .I(n5768), .ZN(n5124) );
  NAND2_X2 U12815 ( .A1(n24584), .A2(n24583), .ZN(n5768) );
  NAND3_X1 U12816 ( .A1(n37648), .A2(n10642), .A3(n28074), .ZN(n3461) );
  NAND2_X2 U12817 ( .A1(n28273), .A2(n988), .ZN(n37648) );
  NOR2_X1 U12834 ( .A1(n19615), .A2(n38742), .ZN(n26769) );
  XOR2_X1 U12836 ( .A1(n35222), .A2(n29088), .Z(n29001) );
  NAND2_X2 U12837 ( .A1(n6370), .A2(n6371), .ZN(n29088) );
  NAND2_X2 U12838 ( .A1(n13213), .A2(n19918), .ZN(n27118) );
  NAND2_X2 U12840 ( .A1(n38871), .A2(n13890), .ZN(n29820) );
  NOR2_X2 U12841 ( .A1(n38924), .A2(n36834), .ZN(n38871) );
  XOR2_X1 U12842 ( .A1(n3560), .A2(n1938), .Z(n3559) );
  XOR2_X1 U12844 ( .A1(n28987), .A2(n39233), .Z(n37650) );
  XOR2_X1 U12845 ( .A1(n7374), .A2(n36510), .Z(n36931) );
  NAND2_X2 U12847 ( .A1(n13860), .A2(n37030), .ZN(n1746) );
  INV_X2 U12853 ( .I(n5227), .ZN(n12394) );
  XNOR2_X1 U12857 ( .A1(n5228), .A2(n5229), .ZN(n5227) );
  NAND2_X2 U12859 ( .A1(n23225), .A2(n14365), .ZN(n37851) );
  XOR2_X1 U12860 ( .A1(n19071), .A2(n37221), .Z(n16942) );
  XOR2_X1 U12863 ( .A1(n35936), .A2(n15202), .Z(n19071) );
  BUF_X2 U12865 ( .I(n24408), .Z(n37651) );
  INV_X2 U12870 ( .I(n37656), .ZN(n38130) );
  NAND3_X2 U12871 ( .A1(n23169), .A2(n36554), .A3(n23167), .ZN(n37656) );
  NAND2_X2 U12876 ( .A1(n37657), .A2(n17500), .ZN(n21110) );
  XOR2_X1 U12878 ( .A1(n8302), .A2(n35241), .Z(n9947) );
  NAND2_X2 U12879 ( .A1(n23081), .A2(n3145), .ZN(n23566) );
  XOR2_X1 U12883 ( .A1(n37658), .A2(n37037), .Z(n32118) );
  XOR2_X1 U12884 ( .A1(n3110), .A2(n25151), .Z(n25198) );
  NOR3_X2 U12888 ( .A1(n21887), .A2(n21889), .A3(n16302), .ZN(n15812) );
  XOR2_X1 U12889 ( .A1(n25063), .A2(n18543), .Z(n3292) );
  XOR2_X1 U12891 ( .A1(n25133), .A2(n24857), .Z(n18543) );
  AOI22_X2 U12893 ( .A1(n5791), .A2(n31829), .B1(n5790), .B2(n17556), .ZN(
        n2932) );
  NAND2_X2 U12901 ( .A1(n20153), .A2(n13545), .ZN(n25483) );
  AOI22_X1 U12906 ( .A1(n23256), .A2(n23515), .B1(n4638), .B2(n4637), .ZN(
        n36279) );
  XNOR2_X1 U12908 ( .A1(n15368), .A2(n37833), .ZN(n39186) );
  XOR2_X1 U12920 ( .A1(n13852), .A2(n8475), .Z(n8474) );
  AOI21_X2 U12923 ( .A1(n35621), .A2(n10758), .B(n10757), .ZN(n13852) );
  BUF_X2 U12926 ( .I(n35920), .Z(n37660) );
  NOR2_X2 U12928 ( .A1(n35449), .A2(n18909), .ZN(n4636) );
  XOR2_X1 U12933 ( .A1(n38581), .A2(n24924), .Z(n25191) );
  NAND2_X2 U12936 ( .A1(n39496), .A2(n17267), .ZN(n38581) );
  AOI21_X1 U12937 ( .A1(n29593), .A2(n38420), .B(n31374), .ZN(n38941) );
  NOR2_X1 U12940 ( .A1(n63), .A2(n29946), .ZN(n14592) );
  INV_X2 U12945 ( .I(n2792), .ZN(n6652) );
  INV_X2 U12948 ( .I(n37662), .ZN(n25718) );
  NAND2_X2 U12956 ( .A1(n37663), .A2(n1855), .ZN(n26125) );
  NAND2_X2 U12957 ( .A1(n1425), .A2(n5418), .ZN(n28365) );
  AOI21_X2 U12960 ( .A1(n37664), .A2(n38073), .B(n35925), .ZN(n10012) );
  NAND3_X2 U12962 ( .A1(n28146), .A2(n28145), .A3(n28144), .ZN(n28686) );
  XOR2_X1 U12970 ( .A1(n22391), .A2(n22542), .Z(n20294) );
  NAND2_X2 U12974 ( .A1(n10744), .A2(n10742), .ZN(n22391) );
  INV_X2 U12981 ( .I(n16237), .ZN(n1477) );
  NAND2_X2 U12982 ( .A1(n30617), .A2(n39542), .ZN(n16237) );
  XOR2_X1 U12983 ( .A1(n6318), .A2(n37666), .Z(n20726) );
  XOR2_X1 U12987 ( .A1(n37665), .A2(n19786), .Z(Ciphertext[148]) );
  NAND4_X2 U12990 ( .A1(n30075), .A2(n30072), .A3(n30074), .A4(n30073), .ZN(
        n37665) );
  OAI21_X2 U12992 ( .A1(n30043), .A2(n29998), .B(n29997), .ZN(n35649) );
  OAI21_X2 U12993 ( .A1(n35653), .A2(n20125), .B(n35649), .ZN(n6919) );
  INV_X2 U12994 ( .I(n3815), .ZN(n30077) );
  NAND2_X2 U12995 ( .A1(n34378), .A2(n31499), .ZN(n3815) );
  XOR2_X1 U13000 ( .A1(n6316), .A2(n20727), .Z(n37666) );
  OR2_X1 U13006 ( .A1(n25309), .A2(n825), .Z(n18233) );
  XOR2_X1 U13014 ( .A1(n37667), .A2(n27706), .Z(n20511) );
  XOR2_X1 U13016 ( .A1(n20513), .A2(n35177), .Z(n37667) );
  XOR2_X1 U13018 ( .A1(n37668), .A2(n6991), .Z(n5899) );
  XOR2_X1 U13019 ( .A1(n6522), .A2(n26500), .Z(n3995) );
  NAND2_X1 U13021 ( .A1(n18234), .A2(n18233), .ZN(n37669) );
  XOR2_X1 U13031 ( .A1(n9030), .A2(n30913), .Z(n6522) );
  XOR2_X1 U13032 ( .A1(n22789), .A2(n20335), .Z(n22522) );
  NOR2_X2 U13035 ( .A1(n11440), .A2(n11439), .ZN(n22789) );
  NOR2_X2 U13038 ( .A1(n31769), .A2(n18776), .ZN(n39424) );
  NAND3_X2 U13053 ( .A1(n39083), .A2(n30213), .A3(n14387), .ZN(n39142) );
  NAND2_X2 U13060 ( .A1(n13488), .A2(n36769), .ZN(n6533) );
  OAI21_X2 U13063 ( .A1(n18743), .A2(n32131), .B(n19061), .ZN(n39249) );
  NAND2_X2 U13067 ( .A1(n39249), .A2(n4570), .ZN(n30908) );
  XOR2_X1 U13070 ( .A1(n5395), .A2(n37786), .Z(n8148) );
  NAND2_X2 U13071 ( .A1(n39222), .A2(n37670), .ZN(n27211) );
  NAND2_X1 U13073 ( .A1(n35612), .A2(n35613), .ZN(n37670) );
  NOR2_X2 U13074 ( .A1(n33407), .A2(n3057), .ZN(n38398) );
  INV_X4 U13076 ( .I(n3697), .ZN(n4225) );
  NAND3_X1 U13078 ( .A1(n6839), .A2(n12975), .A3(n19942), .ZN(n24088) );
  XOR2_X1 U13087 ( .A1(n22763), .A2(n9982), .Z(n22713) );
  AOI22_X2 U13091 ( .A1(n22186), .A2(n35652), .B1(n22188), .B2(n22187), .ZN(
        n22763) );
  NOR2_X2 U13092 ( .A1(n23162), .A2(n23163), .ZN(n22869) );
  XOR2_X1 U13096 ( .A1(n2370), .A2(n2372), .Z(n11573) );
  NOR2_X2 U13099 ( .A1(n39264), .A2(n13197), .ZN(n13196) );
  NOR2_X2 U13102 ( .A1(n5140), .A2(n37672), .ZN(n6756) );
  OAI21_X2 U13103 ( .A1(n1054), .A2(n29859), .B(n11898), .ZN(n11897) );
  XOR2_X1 U13104 ( .A1(n37673), .A2(n22457), .Z(n19002) );
  XOR2_X1 U13107 ( .A1(n36641), .A2(n1656), .Z(n37673) );
  BUF_X2 U13111 ( .I(n23149), .Z(n37674) );
  XOR2_X1 U13112 ( .A1(n37675), .A2(n9994), .Z(n10959) );
  XOR2_X1 U13113 ( .A1(n39520), .A2(n29098), .Z(n37675) );
  XOR2_X1 U13117 ( .A1(n437), .A2(n32959), .Z(n35260) );
  XOR2_X1 U13122 ( .A1(n19074), .A2(n19073), .Z(n32959) );
  XOR2_X1 U13126 ( .A1(n37676), .A2(n35969), .Z(n30736) );
  XOR2_X1 U13127 ( .A1(n16523), .A2(n23961), .Z(n37676) );
  NAND2_X1 U13128 ( .A1(n28626), .A2(n7914), .ZN(n18125) );
  NAND2_X2 U13135 ( .A1(n38065), .A2(n32681), .ZN(n28626) );
  INV_X4 U13137 ( .I(n3642), .ZN(n7258) );
  NAND2_X2 U13143 ( .A1(n14300), .A2(n34297), .ZN(n3642) );
  NAND2_X2 U13144 ( .A1(n15896), .A2(n37677), .ZN(n18743) );
  AOI22_X2 U13150 ( .A1(n9423), .A2(n18870), .B1(n17346), .B2(n8155), .ZN(
        n37677) );
  NOR2_X2 U13153 ( .A1(n37589), .A2(n4473), .ZN(n22683) );
  XOR2_X1 U13154 ( .A1(n28990), .A2(n9787), .Z(n9786) );
  XOR2_X1 U13159 ( .A1(n10080), .A2(n10079), .Z(n28990) );
  INV_X2 U13160 ( .I(n7703), .ZN(n37678) );
  OR2_X1 U13161 ( .A1(n13359), .A2(n37678), .Z(n9466) );
  NAND2_X2 U13162 ( .A1(n37679), .A2(n38010), .ZN(n13458) );
  OAI21_X2 U13164 ( .A1(n21223), .A2(n28249), .B(n28115), .ZN(n37679) );
  OAI21_X1 U13165 ( .A1(n12189), .A2(n10677), .B(n6648), .ZN(n10177) );
  XOR2_X1 U13167 ( .A1(n12441), .A2(n19096), .Z(n24560) );
  XOR2_X1 U13168 ( .A1(n37680), .A2(n19342), .Z(n11627) );
  XOR2_X1 U13170 ( .A1(n7118), .A2(n7119), .Z(n37680) );
  XOR2_X1 U13171 ( .A1(n8670), .A2(n33851), .Z(n13099) );
  XOR2_X1 U13174 ( .A1(n37681), .A2(n15046), .Z(Ciphertext[69]) );
  NOR3_X1 U13176 ( .A1(n39340), .A2(n29569), .A3(n37145), .ZN(n37681) );
  XOR2_X1 U13180 ( .A1(n6435), .A2(n34492), .Z(n28040) );
  NAND2_X2 U13182 ( .A1(n14788), .A2(n31717), .ZN(n5457) );
  OAI22_X2 U13186 ( .A1(n18616), .A2(n15062), .B1(n38320), .B2(n38319), .ZN(
        n14788) );
  NAND2_X2 U13187 ( .A1(n18166), .A2(n22408), .ZN(n7644) );
  XOR2_X1 U13195 ( .A1(n37682), .A2(n29169), .Z(n16371) );
  XOR2_X1 U13199 ( .A1(n38058), .A2(n29038), .Z(n37682) );
  XOR2_X1 U13202 ( .A1(n26302), .A2(n26303), .Z(n38188) );
  XOR2_X1 U13203 ( .A1(n26449), .A2(n26301), .Z(n26302) );
  BUF_X2 U13204 ( .I(n7660), .Z(n37683) );
  NAND3_X2 U13211 ( .A1(n5775), .A2(n5774), .A3(n5771), .ZN(n27537) );
  OAI22_X2 U13212 ( .A1(n13275), .A2(n2254), .B1(n38492), .B2(n2253), .ZN(
        n16048) );
  INV_X2 U13216 ( .I(n7500), .ZN(n14473) );
  NAND2_X2 U13222 ( .A1(n12290), .A2(n26688), .ZN(n26982) );
  OAI21_X2 U13226 ( .A1(n37684), .A2(n24862), .B(n524), .ZN(n15001) );
  NAND2_X2 U13229 ( .A1(n37685), .A2(n8217), .ZN(n8475) );
  NAND2_X1 U13233 ( .A1(n31077), .A2(n8216), .ZN(n37685) );
  XOR2_X1 U13235 ( .A1(n37686), .A2(n19808), .Z(Ciphertext[109]) );
  OAI22_X1 U13237 ( .A1(n39062), .A2(n3612), .B1(n3611), .B2(n29813), .ZN(
        n37686) );
  BUF_X2 U13239 ( .I(n24589), .Z(n37687) );
  XOR2_X1 U13249 ( .A1(n39163), .A2(n38175), .Z(n13074) );
  INV_X4 U13256 ( .I(n24590), .ZN(n24717) );
  NAND2_X2 U13258 ( .A1(n16882), .A2(n16881), .ZN(n24590) );
  NOR2_X2 U13260 ( .A1(n37688), .A2(n19278), .ZN(n20657) );
  NAND2_X2 U13261 ( .A1(n19942), .A2(n24221), .ZN(n20119) );
  NOR2_X2 U13264 ( .A1(n4686), .A2(n6891), .ZN(n34658) );
  NOR2_X2 U13271 ( .A1(n14377), .A2(n19179), .ZN(n4686) );
  NAND2_X2 U13272 ( .A1(n38141), .A2(n2792), .ZN(n29800) );
  AOI22_X2 U13277 ( .A1(n6649), .A2(n19393), .B1(n28960), .B2(n972), .ZN(
        n15189) );
  XOR2_X1 U13278 ( .A1(n30776), .A2(n37689), .Z(n26665) );
  XOR2_X1 U13280 ( .A1(n26375), .A2(n26166), .Z(n37689) );
  XNOR2_X1 U13282 ( .A1(n25310), .A2(n6996), .ZN(n37968) );
  NOR2_X1 U13284 ( .A1(n32111), .A2(n8784), .ZN(n31079) );
  AOI21_X2 U13285 ( .A1(n15767), .A2(n31133), .B(n37690), .ZN(n16525) );
  OAI21_X2 U13286 ( .A1(n31626), .A2(n31133), .B(n25822), .ZN(n37690) );
  NAND2_X2 U13300 ( .A1(n17616), .A2(n7585), .ZN(n27395) );
  NAND3_X1 U13304 ( .A1(n19362), .A2(n29517), .A3(n18384), .ZN(n29521) );
  XOR2_X1 U13307 ( .A1(n10611), .A2(n18428), .Z(n32126) );
  OR2_X1 U13310 ( .A1(n27624), .A2(n31121), .Z(n18131) );
  NAND2_X2 U13311 ( .A1(n17538), .A2(n5405), .ZN(n32851) );
  OAI22_X2 U13316 ( .A1(n6606), .A2(n26932), .B1(n4411), .B2(n5274), .ZN(
        n17538) );
  XOR2_X1 U13317 ( .A1(n23737), .A2(n37691), .Z(n34933) );
  INV_X2 U13318 ( .I(n23709), .ZN(n37691) );
  XOR2_X1 U13323 ( .A1(n13617), .A2(n14289), .Z(n23709) );
  OR2_X1 U13329 ( .A1(n18790), .A2(n10810), .Z(n24371) );
  NAND2_X2 U13331 ( .A1(n37692), .A2(n23539), .ZN(n5181) );
  OAI22_X2 U13334 ( .A1(n23537), .A2(n31332), .B1(n23538), .B2(n12289), .ZN(
        n37692) );
  NAND2_X2 U13338 ( .A1(n37693), .A2(n35005), .ZN(n28621) );
  OR2_X1 U13342 ( .A1(n28232), .A2(n876), .Z(n37693) );
  BUF_X4 U13345 ( .I(n5554), .Z(n36911) );
  CLKBUF_X4 U13346 ( .I(n11569), .Z(n6747) );
  XOR2_X1 U13349 ( .A1(n7125), .A2(n7128), .Z(n32010) );
  NAND2_X2 U13352 ( .A1(n37694), .A2(n39128), .ZN(n6355) );
  NOR2_X1 U13353 ( .A1(n34028), .A2(n36052), .ZN(n36004) );
  NOR2_X2 U13354 ( .A1(n23476), .A2(n21293), .ZN(n35917) );
  NAND2_X2 U13359 ( .A1(n15176), .A2(n38600), .ZN(n23476) );
  NAND3_X2 U13361 ( .A1(n4857), .A2(n37897), .A3(n37695), .ZN(n9108) );
  NAND2_X1 U13362 ( .A1(n11490), .A2(n12537), .ZN(n37695) );
  NAND2_X2 U13364 ( .A1(n446), .A2(n38953), .ZN(n25988) );
  NOR2_X2 U13369 ( .A1(n36720), .A2(n23505), .ZN(n7885) );
  NAND2_X2 U13372 ( .A1(n37696), .A2(n8263), .ZN(n35795) );
  INV_X2 U13373 ( .I(n37697), .ZN(n19990) );
  XNOR2_X1 U13374 ( .A1(n8937), .A2(n38000), .ZN(n37697) );
  NAND2_X2 U13376 ( .A1(n19175), .A2(n38101), .ZN(n31899) );
  BUF_X2 U13377 ( .I(n18209), .Z(n6691) );
  AOI22_X2 U13379 ( .A1(n35048), .A2(n35049), .B1(n24743), .B2(n24744), .ZN(
        n3111) );
  NOR2_X2 U13380 ( .A1(n16999), .A2(n39317), .ZN(n24744) );
  NOR2_X2 U13385 ( .A1(n14993), .A2(n23597), .ZN(n23680) );
  NAND2_X2 U13386 ( .A1(n12373), .A2(n26639), .ZN(n3992) );
  NAND2_X2 U13391 ( .A1(n36726), .A2(n37698), .ZN(n20418) );
  NAND3_X2 U13394 ( .A1(n23061), .A2(n18637), .A3(n20518), .ZN(n37698) );
  BUF_X4 U13395 ( .I(n23142), .Z(n37984) );
  NAND2_X2 U13396 ( .A1(n3077), .A2(n3561), .ZN(n33609) );
  NAND2_X2 U13401 ( .A1(n8766), .A2(n37948), .ZN(n3077) );
  NOR2_X2 U13404 ( .A1(n10474), .A2(n35956), .ZN(n10473) );
  BUF_X2 U13412 ( .I(n19152), .Z(n37699) );
  OAI21_X2 U13417 ( .A1(n34000), .A2(n1962), .B(n37700), .ZN(n39736) );
  AOI21_X2 U13421 ( .A1(n1962), .A2(n20673), .B(n29781), .ZN(n37700) );
  XOR2_X1 U13423 ( .A1(n39760), .A2(n33672), .Z(n23781) );
  INV_X4 U13424 ( .I(n8287), .ZN(n1385) );
  OR2_X1 U13425 ( .A1(n19713), .A2(n37016), .Z(n7830) );
  BUF_X2 U13427 ( .I(n23714), .Z(n37701) );
  XOR2_X1 U13442 ( .A1(n33041), .A2(n1184), .Z(n2032) );
  XOR2_X1 U13443 ( .A1(n12534), .A2(n19862), .Z(n25046) );
  NAND3_X2 U13446 ( .A1(n38331), .A2(n24534), .A3(n37931), .ZN(n19862) );
  NOR2_X1 U13450 ( .A1(n37724), .A2(n10813), .ZN(n37988) );
  INV_X1 U13455 ( .I(n14742), .ZN(n38335) );
  INV_X1 U13457 ( .I(n29009), .ZN(n37729) );
  XOR2_X1 U13460 ( .A1(n22752), .A2(n22581), .Z(n5233) );
  XNOR2_X1 U13462 ( .A1(n5849), .A2(n5851), .ZN(n38445) );
  XOR2_X1 U13464 ( .A1(n14285), .A2(n14533), .Z(n5851) );
  NOR2_X2 U13466 ( .A1(n38695), .A2(n37702), .ZN(n32136) );
  OAI22_X2 U13468 ( .A1(n4702), .A2(n9101), .B1(n16902), .B2(n1035), .ZN(
        n37702) );
  XOR2_X1 U13470 ( .A1(n11695), .A2(n28997), .Z(n29294) );
  NAND2_X2 U13471 ( .A1(n39104), .A2(n13784), .ZN(n28997) );
  OAI21_X1 U13476 ( .A1(n26819), .A2(n7195), .B(n30859), .ZN(n26283) );
  NAND2_X2 U13478 ( .A1(n37705), .A2(n23305), .ZN(n18849) );
  XOR2_X1 U13479 ( .A1(n11161), .A2(n39719), .Z(n36064) );
  NAND2_X2 U13481 ( .A1(n37706), .A2(n19460), .ZN(n32646) );
  NAND2_X1 U13484 ( .A1(n30615), .A2(n30613), .ZN(n37706) );
  XOR2_X1 U13486 ( .A1(n27679), .A2(n27633), .Z(n27765) );
  NAND2_X2 U13489 ( .A1(n27038), .A2(n18861), .ZN(n27679) );
  XOR2_X1 U13490 ( .A1(n16085), .A2(n27726), .Z(n8563) );
  XOR2_X1 U13492 ( .A1(n12556), .A2(n4885), .Z(n27726) );
  BUF_X4 U13494 ( .I(n2046), .Z(n1989) );
  XOR2_X1 U13499 ( .A1(n7942), .A2(n37707), .Z(n3476) );
  XOR2_X1 U13501 ( .A1(n3478), .A2(n359), .Z(n37707) );
  NAND2_X2 U13502 ( .A1(n15946), .A2(n39521), .ZN(n30913) );
  NOR2_X1 U13508 ( .A1(n29810), .A2(n29803), .ZN(n3614) );
  NAND2_X2 U13509 ( .A1(n28923), .A2(n28924), .ZN(n29810) );
  NAND2_X2 U13511 ( .A1(n37708), .A2(n38640), .ZN(n17756) );
  OAI21_X2 U13515 ( .A1(n37803), .A2(n31270), .B(n6849), .ZN(n30684) );
  NAND2_X2 U13519 ( .A1(n37709), .A2(n38484), .ZN(n22376) );
  NAND2_X1 U13526 ( .A1(n36090), .A2(n7852), .ZN(n8580) );
  NAND2_X1 U13536 ( .A1(n10004), .A2(n1257), .ZN(n37712) );
  INV_X1 U13549 ( .I(n18249), .ZN(n37713) );
  XOR2_X1 U13551 ( .A1(n14264), .A2(n13245), .Z(n10129) );
  INV_X1 U13552 ( .I(n38785), .ZN(n38784) );
  XOR2_X1 U13553 ( .A1(n28842), .A2(n8371), .Z(n1914) );
  XOR2_X1 U13558 ( .A1(n29147), .A2(n1915), .Z(n8371) );
  NAND2_X2 U13559 ( .A1(n37714), .A2(n2342), .ZN(n2634) );
  NOR2_X2 U13561 ( .A1(n15898), .A2(n33500), .ZN(n37714) );
  NAND2_X2 U13565 ( .A1(n9508), .A2(n19508), .ZN(n33855) );
  XOR2_X1 U13571 ( .A1(n37715), .A2(n23921), .Z(n11699) );
  XOR2_X1 U13572 ( .A1(n8904), .A2(n39177), .Z(n37715) );
  XOR2_X1 U13574 ( .A1(n4123), .A2(n4210), .Z(n4209) );
  NAND2_X2 U13576 ( .A1(n30877), .A2(n30354), .ZN(n4210) );
  NAND2_X2 U13577 ( .A1(n33461), .A2(n5619), .ZN(n31612) );
  AND2_X2 U13579 ( .A1(n25639), .A2(n25669), .Z(n3101) );
  XOR2_X1 U13580 ( .A1(n39219), .A2(n29294), .Z(n15091) );
  XOR2_X1 U13591 ( .A1(n2126), .A2(n5246), .Z(n7582) );
  NAND2_X2 U13595 ( .A1(n36795), .A2(n3909), .ZN(n2126) );
  AOI21_X1 U13600 ( .A1(n14337), .A2(n29722), .B(n29719), .ZN(n29705) );
  AOI22_X2 U13604 ( .A1(n32192), .A2(n4448), .B1(n29703), .B2(n4447), .ZN(
        n29722) );
  INV_X1 U13607 ( .I(n32228), .ZN(n1655) );
  AND2_X1 U13608 ( .A1(n32228), .A2(n19840), .Z(n32202) );
  OAI22_X2 U13609 ( .A1(n2772), .A2(n8942), .B1(n5628), .B2(n8707), .ZN(n31325) );
  AOI22_X2 U13613 ( .A1(n29430), .A2(n37716), .B1(n35517), .B2(n34194), .ZN(
        n18502) );
  NAND2_X1 U13617 ( .A1(n15089), .A2(n29497), .ZN(n37716) );
  XOR2_X1 U13623 ( .A1(n37718), .A2(n38875), .Z(n9791) );
  XOR2_X1 U13625 ( .A1(n11730), .A2(n39515), .Z(n37718) );
  INV_X2 U13632 ( .I(n10216), .ZN(n2182) );
  NAND3_X2 U13633 ( .A1(n39588), .A2(n13077), .A3(n13078), .ZN(n10216) );
  INV_X2 U13634 ( .I(n33949), .ZN(n36162) );
  OAI21_X2 U13637 ( .A1(n35788), .A2(n35789), .B(n19827), .ZN(n37719) );
  XOR2_X1 U13641 ( .A1(n4077), .A2(n37720), .Z(n4081) );
  XOR2_X1 U13643 ( .A1(n30913), .A2(n1238), .Z(n37720) );
  XOR2_X1 U13651 ( .A1(n37721), .A2(n12972), .Z(n10872) );
  NAND2_X2 U13655 ( .A1(n36966), .A2(n31446), .ZN(n12972) );
  NAND2_X2 U13659 ( .A1(n29781), .A2(n29777), .ZN(n39154) );
  NAND2_X2 U13660 ( .A1(n39154), .A2(n29779), .ZN(n38574) );
  XOR2_X1 U13662 ( .A1(n37723), .A2(n37722), .Z(n12334) );
  XOR2_X1 U13663 ( .A1(n4815), .A2(n27641), .Z(n37722) );
  XOR2_X1 U13666 ( .A1(n27642), .A2(n20641), .Z(n37723) );
  OAI22_X2 U13667 ( .A1(n17502), .A2(n7915), .B1(n32747), .B2(n32520), .ZN(
        n10458) );
  XOR2_X1 U13672 ( .A1(n29037), .A2(n37725), .Z(n38136) );
  XOR2_X1 U13674 ( .A1(n37726), .A2(n14956), .Z(n37725) );
  AOI21_X2 U13679 ( .A1(n36701), .A2(n36011), .B(n1695), .ZN(n37763) );
  XNOR2_X1 U13682 ( .A1(n33756), .A2(n32646), .ZN(n514) );
  NAND2_X2 U13683 ( .A1(n29010), .A2(n37728), .ZN(n37727) );
  INV_X2 U13684 ( .I(n20525), .ZN(n37728) );
  BUF_X4 U13687 ( .I(n25319), .Z(n39491) );
  INV_X2 U13688 ( .I(n37731), .ZN(n21768) );
  XNOR2_X1 U13691 ( .A1(Key[161]), .A2(Plaintext[161]), .ZN(n37731) );
  OAI21_X2 U13694 ( .A1(n23302), .A2(n32017), .B(n23489), .ZN(n529) );
  BUF_X2 U13699 ( .I(n30186), .Z(n37734) );
  NAND2_X2 U13702 ( .A1(n34205), .A2(n37735), .ZN(n30358) );
  OAI21_X2 U13706 ( .A1(n37173), .A2(n37736), .B(n36133), .ZN(n36460) );
  NOR2_X2 U13708 ( .A1(n36162), .A2(n3985), .ZN(n37736) );
  INV_X4 U13709 ( .I(n36385), .ZN(n1271) );
  NAND2_X2 U13712 ( .A1(n13706), .A2(n13709), .ZN(n36385) );
  XOR2_X1 U13713 ( .A1(n27723), .A2(n27635), .Z(n7022) );
  XOR2_X1 U13715 ( .A1(n27829), .A2(n27595), .Z(n27723) );
  NAND3_X2 U13717 ( .A1(n38960), .A2(n19584), .A3(n24443), .ZN(n24313) );
  XOR2_X1 U13731 ( .A1(n37738), .A2(n23789), .Z(n23926) );
  NAND2_X2 U13737 ( .A1(n32025), .A2(n23093), .ZN(n23568) );
  NOR2_X2 U13739 ( .A1(n12050), .A2(n37739), .ZN(n24668) );
  AND2_X1 U13756 ( .A1(n13040), .A2(n5954), .Z(n37739) );
  NOR2_X2 U13760 ( .A1(n31144), .A2(n37740), .ZN(n31143) );
  NOR3_X2 U13761 ( .A1(n1570), .A2(n24750), .A3(n38182), .ZN(n37740) );
  XOR2_X1 U13763 ( .A1(n24039), .A2(n24028), .Z(n36760) );
  XOR2_X1 U13765 ( .A1(n17925), .A2(n35235), .Z(n24028) );
  AOI22_X2 U13775 ( .A1(n39260), .A2(n37102), .B1(n38138), .B2(n10340), .ZN(
        n35750) );
  AOI21_X2 U13777 ( .A1(n23360), .A2(n23359), .B(n31594), .ZN(n38650) );
  INV_X2 U13778 ( .I(n281), .ZN(n28143) );
  XOR2_X1 U13779 ( .A1(n11856), .A2(n37741), .Z(n16699) );
  XOR2_X1 U13780 ( .A1(n25251), .A2(n10215), .Z(n37741) );
  NAND2_X2 U13782 ( .A1(n9499), .A2(n37742), .ZN(n10225) );
  XOR2_X1 U13783 ( .A1(n29824), .A2(n28852), .Z(n13381) );
  NAND2_X2 U13786 ( .A1(n35574), .A2(n12607), .ZN(n29824) );
  NAND3_X1 U13789 ( .A1(n28671), .A2(n28674), .A3(n18883), .ZN(n15959) );
  XOR2_X1 U13791 ( .A1(n20095), .A2(n15545), .Z(n38081) );
  NOR2_X1 U13793 ( .A1(n35368), .A2(n13620), .ZN(n13618) );
  XOR2_X1 U13798 ( .A1(n27759), .A2(n27760), .Z(n36863) );
  XOR2_X1 U13801 ( .A1(n38937), .A2(n17349), .Z(n27759) );
  OR2_X1 U13804 ( .A1(n26724), .A2(n26832), .Z(n26679) );
  OAI21_X2 U13805 ( .A1(n21587), .A2(n14499), .B(n8597), .ZN(n21413) );
  NOR2_X2 U13808 ( .A1(n20979), .A2(n29642), .ZN(n37743) );
  XOR2_X1 U13809 ( .A1(n37744), .A2(n8502), .Z(n39027) );
  XOR2_X1 U13812 ( .A1(n33812), .A2(n38495), .Z(n37744) );
  INV_X2 U13814 ( .I(n32134), .ZN(n6592) );
  XOR2_X1 U13821 ( .A1(n13920), .A2(n6595), .Z(n32134) );
  OAI22_X2 U13822 ( .A1(n19590), .A2(n16200), .B1(n1518), .B2(n32469), .ZN(
        n37745) );
  XOR2_X1 U13827 ( .A1(n29098), .A2(n28916), .Z(n28878) );
  XOR2_X1 U13829 ( .A1(n18305), .A2(n15745), .Z(n29098) );
  XOR2_X1 U13832 ( .A1(n27459), .A2(n27715), .Z(n14359) );
  XOR2_X1 U13837 ( .A1(n31551), .A2(n34963), .Z(n27459) );
  XOR2_X1 U13838 ( .A1(n23878), .A2(n20877), .Z(n2596) );
  XOR2_X1 U13840 ( .A1(n1617), .A2(n24079), .Z(n23878) );
  NAND2_X2 U13844 ( .A1(n31640), .A2(n5787), .ZN(n10764) );
  XOR2_X1 U13847 ( .A1(n26558), .A2(n3152), .Z(n3151) );
  NAND2_X2 U13848 ( .A1(n37747), .A2(n35670), .ZN(n31937) );
  NAND2_X2 U13850 ( .A1(n34504), .A2(n1602), .ZN(n37747) );
  XOR2_X1 U13855 ( .A1(n23975), .A2(n23742), .Z(n11119) );
  OAI21_X2 U13859 ( .A1(n19246), .A2(n39045), .B(n37749), .ZN(n17931) );
  NOR2_X2 U13860 ( .A1(n37750), .A2(n15452), .ZN(n1627) );
  XOR2_X1 U13861 ( .A1(n25144), .A2(n25318), .Z(n32532) );
  NAND3_X1 U13864 ( .A1(n38012), .A2(n5038), .A3(n39350), .ZN(n20191) );
  XNOR2_X1 U13865 ( .A1(n22470), .A2(n22567), .ZN(n37869) );
  AOI22_X2 U13878 ( .A1(n20013), .A2(n24664), .B1(n37751), .B2(n2340), .ZN(
        n16051) );
  NOR2_X2 U13879 ( .A1(n35578), .A2(n38523), .ZN(n37751) );
  XOR2_X1 U13883 ( .A1(n16900), .A2(n33271), .Z(n10611) );
  NAND2_X2 U13884 ( .A1(n7396), .A2(n4729), .ZN(n16900) );
  INV_X1 U13885 ( .I(n20010), .ZN(n37753) );
  NOR3_X2 U13886 ( .A1(n36662), .A2(n3411), .A3(n3410), .ZN(n3409) );
  XOR2_X1 U13891 ( .A1(n7553), .A2(n26570), .Z(n18738) );
  XOR2_X1 U13894 ( .A1(n26571), .A2(n6177), .Z(n7553) );
  AOI22_X2 U13895 ( .A1(n7479), .A2(n10702), .B1(n19544), .B2(n11677), .ZN(
        n3463) );
  NOR2_X2 U13905 ( .A1(n34264), .A2(n4215), .ZN(n26029) );
  XOR2_X1 U13906 ( .A1(n11050), .A2(n37755), .Z(n38026) );
  XOR2_X1 U13910 ( .A1(n37889), .A2(n35257), .Z(n37755) );
  XOR2_X1 U13919 ( .A1(n7981), .A2(n37756), .Z(n23682) );
  XOR2_X1 U13920 ( .A1(n24058), .A2(n17398), .Z(n37756) );
  INV_X2 U13928 ( .I(n4599), .ZN(n33561) );
  OR2_X1 U13930 ( .A1(n1265), .A2(n24737), .Z(n38738) );
  OAI21_X2 U13937 ( .A1(n2581), .A2(n25466), .B(n35271), .ZN(n36499) );
  NOR2_X2 U13948 ( .A1(n220), .A2(n591), .ZN(n2581) );
  BUF_X2 U13949 ( .I(n35534), .Z(n37757) );
  OAI22_X2 U13953 ( .A1(n33325), .A2(n28457), .B1(n1823), .B2(n28458), .ZN(
        n37759) );
  NAND3_X1 U13954 ( .A1(n25999), .A2(n31362), .A3(n35138), .ZN(n2493) );
  OAI21_X2 U13958 ( .A1(n8698), .A2(n35749), .B(n14041), .ZN(n8697) );
  NAND2_X1 U13959 ( .A1(n34069), .A2(n28276), .ZN(n35844) );
  OR2_X1 U13964 ( .A1(n2654), .A2(n36371), .Z(n30893) );
  OAI21_X2 U13965 ( .A1(n8154), .A2(n17194), .B(n19222), .ZN(n9367) );
  BUF_X4 U13967 ( .I(n39477), .Z(n38519) );
  XOR2_X1 U13969 ( .A1(n37761), .A2(n39559), .Z(Ciphertext[46]) );
  AOI22_X1 U13971 ( .A1(n15132), .A2(n15131), .B1(n15128), .B2(n15127), .ZN(
        n37761) );
  XOR2_X1 U13975 ( .A1(n23891), .A2(n23892), .Z(n23897) );
  XOR2_X1 U13977 ( .A1(n24061), .A2(n23808), .Z(n23891) );
  NOR2_X2 U13978 ( .A1(n11247), .A2(n25759), .ZN(n38584) );
  NAND2_X2 U13989 ( .A1(n37762), .A2(n25443), .ZN(n11734) );
  NAND3_X2 U13996 ( .A1(n37949), .A2(n30399), .A3(n9305), .ZN(n37762) );
  INV_X1 U13997 ( .I(n37763), .ZN(n11987) );
  XOR2_X1 U13999 ( .A1(n37765), .A2(n37764), .Z(n18220) );
  XOR2_X1 U14000 ( .A1(n487), .A2(n7337), .Z(n37765) );
  XOR2_X1 U14008 ( .A1(n22527), .A2(n1368), .Z(n39693) );
  OAI22_X2 U14012 ( .A1(n7105), .A2(n20376), .B1(n31953), .B2(n7104), .ZN(
        n22527) );
  XOR2_X1 U14018 ( .A1(n17606), .A2(n13935), .Z(n24955) );
  INV_X2 U14022 ( .I(n38385), .ZN(n38905) );
  XOR2_X1 U14032 ( .A1(n3917), .A2(n38385), .Z(n3773) );
  NOR2_X2 U14062 ( .A1(n35018), .A2(n31816), .ZN(n38385) );
  XOR2_X1 U14072 ( .A1(n26254), .A2(n15010), .Z(n21085) );
  XOR2_X1 U14074 ( .A1(n8634), .A2(n23807), .Z(n30891) );
  XOR2_X1 U14075 ( .A1(n24030), .A2(n238), .Z(n8634) );
  AOI22_X2 U14078 ( .A1(n9672), .A2(n23522), .B1(n36878), .B2(n9190), .ZN(
        n35885) );
  XOR2_X1 U14079 ( .A1(n37767), .A2(n4270), .Z(n3585) );
  XOR2_X1 U14083 ( .A1(n3475), .A2(n22711), .Z(n37767) );
  INV_X4 U14085 ( .I(n2616), .ZN(n16841) );
  AOI21_X2 U14097 ( .A1(n37142), .A2(n21472), .B(n37768), .ZN(n22250) );
  AOI22_X1 U14101 ( .A1(n21617), .A2(n18293), .B1(n19372), .B2(n917), .ZN(
        n37768) );
  XOR2_X1 U14106 ( .A1(n26518), .A2(n31293), .Z(n26221) );
  NAND2_X2 U14108 ( .A1(n16952), .A2(n25914), .ZN(n26518) );
  XOR2_X1 U14111 ( .A1(n11602), .A2(n34911), .Z(n15566) );
  INV_X2 U14116 ( .I(n37769), .ZN(n38166) );
  NAND3_X2 U14117 ( .A1(n29597), .A2(n29596), .A3(n29595), .ZN(n37769) );
  INV_X1 U14126 ( .I(n19997), .ZN(n37770) );
  NOR2_X2 U14127 ( .A1(n38368), .A2(n5385), .ZN(n34632) );
  INV_X4 U14129 ( .I(n29452), .ZN(n14151) );
  XOR2_X1 U14131 ( .A1(n29041), .A2(n28966), .Z(n29090) );
  XOR2_X1 U14132 ( .A1(n31599), .A2(n23965), .Z(n8400) );
  AOI21_X2 U14133 ( .A1(n23356), .A2(n39534), .B(n33696), .ZN(n31599) );
  XOR2_X1 U14134 ( .A1(n17703), .A2(n14603), .Z(n8888) );
  XOR2_X1 U14135 ( .A1(n6435), .A2(n37951), .Z(n17703) );
  NAND2_X2 U14140 ( .A1(n5209), .A2(n10373), .ZN(n7328) );
  NAND2_X2 U14147 ( .A1(n35248), .A2(n36105), .ZN(n12944) );
  NOR2_X2 U14148 ( .A1(n12406), .A2(n14397), .ZN(n27870) );
  NAND2_X2 U14153 ( .A1(n7751), .A2(n19168), .ZN(n33747) );
  XOR2_X1 U14161 ( .A1(n35222), .A2(n18362), .Z(n3140) );
  BUF_X2 U14166 ( .I(n14260), .Z(n37833) );
  XOR2_X1 U14167 ( .A1(n18808), .A2(n37772), .Z(n36962) );
  XOR2_X1 U14169 ( .A1(n31293), .A2(n39662), .Z(n37772) );
  BUF_X2 U14171 ( .I(n10764), .Z(n32520) );
  XOR2_X1 U14172 ( .A1(n16566), .A2(n26508), .Z(n4572) );
  NAND2_X2 U14176 ( .A1(n37773), .A2(n29771), .ZN(n15867) );
  NAND2_X1 U14181 ( .A1(n20895), .A2(n20894), .ZN(n37773) );
  AND2_X1 U14190 ( .A1(n11970), .A2(n37774), .Z(n11969) );
  XOR2_X1 U14193 ( .A1(n37995), .A2(n26510), .Z(n33750) );
  NAND2_X2 U14194 ( .A1(n25918), .A2(n25917), .ZN(n26510) );
  XOR2_X1 U14197 ( .A1(n24023), .A2(n24065), .Z(n17563) );
  NOR2_X2 U14201 ( .A1(n37777), .A2(n37776), .ZN(n34639) );
  INV_X2 U14202 ( .I(n39423), .ZN(n37776) );
  NOR2_X2 U14204 ( .A1(n37976), .A2(n11797), .ZN(n16057) );
  XOR2_X1 U14205 ( .A1(n25315), .A2(n17606), .Z(n2618) );
  XOR2_X1 U14208 ( .A1(n25296), .A2(n25196), .Z(n25315) );
  NOR2_X2 U14210 ( .A1(n6747), .A2(n1545), .ZN(n25666) );
  NAND2_X1 U14212 ( .A1(n37539), .A2(n39196), .ZN(n6186) );
  XOR2_X1 U14213 ( .A1(n37778), .A2(n4564), .Z(n16445) );
  XOR2_X1 U14214 ( .A1(n21257), .A2(n4563), .Z(n37778) );
  XOR2_X1 U14215 ( .A1(n14297), .A2(n12101), .Z(n30842) );
  XOR2_X1 U14218 ( .A1(n22439), .A2(n1668), .Z(n14297) );
  AOI21_X2 U14219 ( .A1(n6184), .A2(n6183), .B(n6189), .ZN(n6185) );
  NAND2_X2 U14221 ( .A1(n31200), .A2(n37779), .ZN(n23976) );
  AND2_X1 U14222 ( .A1(n9694), .A2(n4553), .Z(n19898) );
  XOR2_X1 U14226 ( .A1(n9274), .A2(n2815), .Z(n18383) );
  OAI21_X2 U14230 ( .A1(n29775), .A2(n18222), .B(n37780), .ZN(n29797) );
  NOR2_X2 U14232 ( .A1(n18221), .A2(n17912), .ZN(n37780) );
  NAND2_X1 U14235 ( .A1(n28017), .A2(n31494), .ZN(n37785) );
  XOR2_X1 U14236 ( .A1(n27718), .A2(n5394), .Z(n37786) );
  XOR2_X1 U14242 ( .A1(n404), .A2(n37787), .Z(n20945) );
  XOR2_X1 U14243 ( .A1(n29000), .A2(n37256), .Z(n37787) );
  OAI21_X2 U14249 ( .A1(n3742), .A2(n34249), .B(n32256), .ZN(n37788) );
  NAND2_X1 U14250 ( .A1(n30465), .A2(n6747), .ZN(n20440) );
  AOI21_X2 U14252 ( .A1(n8752), .A2(n22401), .B(n8750), .ZN(n35824) );
  OAI21_X2 U14253 ( .A1(n21497), .A2(n38878), .B(n21309), .ZN(n37789) );
  XOR2_X1 U14254 ( .A1(n9576), .A2(n2055), .Z(n19973) );
  NAND2_X2 U14255 ( .A1(n5679), .A2(n5683), .ZN(n2055) );
  XOR2_X1 U14257 ( .A1(n37790), .A2(n33429), .Z(n19170) );
  XOR2_X1 U14262 ( .A1(n3787), .A2(n38440), .Z(n37790) );
  NAND3_X2 U14266 ( .A1(n7014), .A2(n7012), .A3(n7013), .ZN(n35232) );
  NAND2_X2 U14267 ( .A1(n38574), .A2(n481), .ZN(n2560) );
  AOI22_X2 U14274 ( .A1(n37792), .A2(n37791), .B1(n22368), .B2(n17319), .ZN(
        n16528) );
  XOR2_X1 U14279 ( .A1(n28888), .A2(n17325), .Z(n39247) );
  INV_X2 U14281 ( .I(n8787), .ZN(n28494) );
  NAND3_X2 U14282 ( .A1(n28352), .A2(n12885), .A3(n28349), .ZN(n8787) );
  NAND2_X1 U14283 ( .A1(n35551), .A2(n19693), .ZN(n35695) );
  NOR2_X1 U14284 ( .A1(n20943), .A2(n20351), .ZN(n37793) );
  XOR2_X1 U14287 ( .A1(n26255), .A2(n5848), .Z(n26417) );
  NAND2_X2 U14291 ( .A1(n30967), .A2(n31630), .ZN(n5241) );
  BUF_X2 U14293 ( .I(n2803), .Z(n37795) );
  XOR2_X1 U14294 ( .A1(n24061), .A2(n23762), .Z(n23944) );
  OAI22_X2 U14295 ( .A1(n17787), .A2(n14649), .B1(n17788), .B2(n38252), .ZN(
        n24061) );
  XOR2_X1 U14297 ( .A1(n27542), .A2(n13374), .Z(n27654) );
  AOI22_X2 U14298 ( .A1(n10356), .A2(n10357), .B1(n10358), .B2(n1474), .ZN(
        n13374) );
  XOR2_X1 U14299 ( .A1(n28878), .A2(n34773), .Z(n18967) );
  AOI22_X2 U14302 ( .A1(n15918), .A2(n4434), .B1(n27410), .B2(n15917), .ZN(
        n4462) );
  NAND2_X1 U14306 ( .A1(n1414), .A2(n38629), .ZN(n28480) );
  NAND2_X2 U14312 ( .A1(n20020), .A2(n28104), .ZN(n38629) );
  AOI22_X2 U14316 ( .A1(n24165), .A2(n39156), .B1(n1282), .B2(n23704), .ZN(
        n24584) );
  NOR2_X1 U14321 ( .A1(n6331), .A2(n20601), .ZN(n23704) );
  XOR2_X1 U14325 ( .A1(n2445), .A2(n39550), .Z(n7500) );
  XOR2_X1 U14326 ( .A1(n6987), .A2(n37796), .Z(n15935) );
  XOR2_X1 U14329 ( .A1(n1614), .A2(n13978), .Z(n37796) );
  XOR2_X1 U14331 ( .A1(n25173), .A2(n25172), .Z(n36959) );
  XOR2_X1 U14332 ( .A1(n25214), .A2(n8183), .Z(n25173) );
  XOR2_X1 U14335 ( .A1(n26399), .A2(n15595), .Z(n13658) );
  XOR2_X1 U14336 ( .A1(n26117), .A2(n31965), .Z(n15595) );
  AND2_X1 U14341 ( .A1(n15284), .A2(n39484), .Z(n26694) );
  NAND2_X2 U14355 ( .A1(n38232), .A2(n31406), .ZN(n15284) );
  NAND2_X2 U14356 ( .A1(n38805), .A2(n37797), .ZN(n29439) );
  OAI21_X2 U14358 ( .A1(n25347), .A2(n4013), .B(n25346), .ZN(n31115) );
  NAND2_X2 U14359 ( .A1(n3337), .A2(n13861), .ZN(n13860) );
  NOR2_X2 U14365 ( .A1(n3784), .A2(n13855), .ZN(n3337) );
  NAND2_X2 U14373 ( .A1(n26928), .A2(n26927), .ZN(n37798) );
  AOI21_X2 U14374 ( .A1(n19993), .A2(n16790), .B(n34000), .ZN(n16845) );
  NAND3_X2 U14378 ( .A1(n4931), .A2(n5702), .A3(n33972), .ZN(n37982) );
  XOR2_X1 U14379 ( .A1(n37799), .A2(n19890), .Z(Ciphertext[43]) );
  NAND3_X1 U14387 ( .A1(n12340), .A2(n12339), .A3(n12321), .ZN(n37799) );
  XOR2_X1 U14390 ( .A1(n37800), .A2(n14715), .Z(n25598) );
  XOR2_X1 U14392 ( .A1(n720), .A2(n25002), .Z(n37800) );
  OAI21_X1 U14394 ( .A1(n4576), .A2(n23426), .B(n32024), .ZN(n37802) );
  XOR2_X1 U14397 ( .A1(n27501), .A2(n12341), .Z(n27760) );
  AOI22_X2 U14400 ( .A1(n8268), .A2(n1625), .B1(n23531), .B2(n8269), .ZN(
        n33462) );
  AND2_X1 U14403 ( .A1(n25597), .A2(n1254), .Z(n33407) );
  NAND2_X1 U14408 ( .A1(n4613), .A2(n4342), .ZN(n37805) );
  INV_X2 U14410 ( .I(n6691), .ZN(n36724) );
  XOR2_X1 U14413 ( .A1(n37806), .A2(n29974), .Z(Ciphertext[135]) );
  NAND3_X2 U14415 ( .A1(n32570), .A2(n7270), .A3(n7271), .ZN(n37806) );
  XOR2_X1 U14423 ( .A1(n29094), .A2(n29255), .Z(n14981) );
  NAND3_X2 U14424 ( .A1(n7752), .A2(n9269), .A3(n16970), .ZN(n20094) );
  AND2_X1 U14426 ( .A1(n4613), .A2(n22337), .Z(n22102) );
  OAI21_X1 U14428 ( .A1(n19442), .A2(n14000), .B(n35197), .ZN(n11421) );
  XOR2_X1 U14430 ( .A1(n37807), .A2(n27844), .Z(n38054) );
  XOR2_X1 U14437 ( .A1(n15421), .A2(n27554), .Z(n37807) );
  OR2_X1 U14441 ( .A1(n23517), .A2(n39001), .Z(n38536) );
  XOR2_X1 U14445 ( .A1(n37808), .A2(n26201), .Z(n26770) );
  XOR2_X1 U14446 ( .A1(n32934), .A2(n26200), .Z(n37808) );
  OR2_X1 U14450 ( .A1(n24747), .A2(n24601), .Z(n19999) );
  NAND2_X2 U14453 ( .A1(n16196), .A2(n37983), .ZN(n24747) );
  NOR2_X2 U14454 ( .A1(n23201), .A2(n35576), .ZN(n15200) );
  NAND2_X2 U14455 ( .A1(n37810), .A2(n3437), .ZN(n22196) );
  NAND2_X1 U14458 ( .A1(n20844), .A2(n9316), .ZN(n37810) );
  XOR2_X1 U14459 ( .A1(n31445), .A2(n37811), .Z(n10665) );
  XOR2_X1 U14462 ( .A1(n25171), .A2(n16555), .Z(n37811) );
  AOI21_X2 U14463 ( .A1(n29202), .A2(n33488), .B(n37813), .ZN(n39829) );
  NOR2_X1 U14464 ( .A1(n10779), .A2(n1436), .ZN(n38764) );
  BUF_X2 U14465 ( .I(n36150), .Z(n37815) );
  XOR2_X1 U14466 ( .A1(n4305), .A2(n39725), .Z(n37816) );
  OR2_X1 U14467 ( .A1(n5886), .A2(n26048), .Z(n8898) );
  INV_X2 U14474 ( .I(n29220), .ZN(n13107) );
  NAND2_X2 U14475 ( .A1(n32189), .A2(n38071), .ZN(n29220) );
  NAND2_X2 U14476 ( .A1(n16348), .A2(n16347), .ZN(n19094) );
  NAND2_X2 U14478 ( .A1(n17557), .A2(n2458), .ZN(n16348) );
  AOI22_X2 U14480 ( .A1(n9508), .A2(n5471), .B1(n18816), .B2(n5570), .ZN(n3247) );
  XOR2_X1 U14481 ( .A1(n3015), .A2(n25292), .Z(n8003) );
  NOR2_X2 U14483 ( .A1(n2905), .A2(n2903), .ZN(n25292) );
  AND2_X1 U14487 ( .A1(n11145), .A2(n14332), .Z(n32536) );
  NAND3_X1 U14488 ( .A1(n32783), .A2(n13714), .A3(n15597), .ZN(n32235) );
  AND2_X1 U14491 ( .A1(n2117), .A2(n32310), .Z(n24314) );
  NOR2_X1 U14494 ( .A1(n13005), .A2(n19249), .ZN(n38995) );
  INV_X2 U14500 ( .I(n25860), .ZN(n1520) );
  XOR2_X1 U14501 ( .A1(n17399), .A2(n3126), .Z(n3117) );
  XOR2_X1 U14505 ( .A1(n29045), .A2(n30964), .Z(n17399) );
  XOR2_X1 U14508 ( .A1(n37817), .A2(n23913), .Z(n31505) );
  XOR2_X1 U14509 ( .A1(n10312), .A2(n1619), .Z(n37817) );
  AOI21_X2 U14512 ( .A1(n34608), .A2(n37818), .B(n36314), .ZN(n38318) );
  NAND2_X2 U14515 ( .A1(n35745), .A2(n31433), .ZN(n37818) );
  XOR2_X1 U14516 ( .A1(n16296), .A2(n23939), .Z(n8904) );
  NAND2_X2 U14519 ( .A1(n39218), .A2(n23322), .ZN(n16296) );
  OR2_X1 U14521 ( .A1(n8395), .A2(n8604), .Z(n8291) );
  OAI21_X1 U14522 ( .A1(n38830), .A2(n20391), .B(n22058), .ZN(n16403) );
  XOR2_X1 U14525 ( .A1(n34544), .A2(n27646), .Z(n18474) );
  XOR2_X1 U14526 ( .A1(n6960), .A2(n37820), .Z(n36847) );
  XOR2_X1 U14527 ( .A1(n26234), .A2(n17396), .Z(n37820) );
  NAND3_X2 U14529 ( .A1(n8491), .A2(n1042), .A3(n35684), .ZN(n10437) );
  NAND2_X2 U14536 ( .A1(n23255), .A2(n33702), .ZN(n19536) );
  NAND2_X1 U14537 ( .A1(n24371), .A2(n24370), .ZN(n13070) );
  XOR2_X1 U14538 ( .A1(n39804), .A2(n16898), .Z(n14106) );
  NOR2_X2 U14539 ( .A1(n21338), .A2(n19216), .ZN(n39804) );
  XOR2_X1 U14542 ( .A1(n8852), .A2(n31127), .Z(n29153) );
  OAI21_X2 U14544 ( .A1(n38127), .A2(n28759), .B(n8449), .ZN(n8852) );
  XOR2_X1 U14545 ( .A1(n34998), .A2(n5703), .Z(n35724) );
  XOR2_X1 U14546 ( .A1(n37998), .A2(n39744), .Z(n32556) );
  XOR2_X1 U14547 ( .A1(n38585), .A2(n2712), .Z(n30503) );
  XOR2_X1 U14548 ( .A1(n6719), .A2(n14307), .Z(n29038) );
  NAND2_X2 U14549 ( .A1(n38077), .A2(n4005), .ZN(n14307) );
  XNOR2_X1 U14550 ( .A1(n1010), .A2(n5084), .ZN(n26420) );
  NAND2_X2 U14554 ( .A1(n8380), .A2(n8381), .ZN(n5625) );
  NAND2_X2 U14556 ( .A1(n8383), .A2(n8385), .ZN(n8380) );
  NOR2_X2 U14562 ( .A1(n37823), .A2(n37822), .ZN(n17249) );
  INV_X1 U14564 ( .I(n5131), .ZN(n37822) );
  INV_X2 U14566 ( .I(n21912), .ZN(n37823) );
  NAND2_X2 U14571 ( .A1(n37824), .A2(n15201), .ZN(n8693) );
  OAI21_X2 U14575 ( .A1(n15200), .A2(n15199), .B(n22849), .ZN(n37824) );
  XOR2_X1 U14577 ( .A1(n37825), .A2(n19676), .Z(Ciphertext[177]) );
  XOR2_X1 U14579 ( .A1(n13917), .A2(n25267), .Z(n14955) );
  OAI21_X2 U14589 ( .A1(n36485), .A2(n24113), .B(n24101), .ZN(n13316) );
  OAI21_X2 U14593 ( .A1(n16890), .A2(n2498), .B(n692), .ZN(n39164) );
  XOR2_X1 U14594 ( .A1(n4929), .A2(n14953), .Z(n11092) );
  INV_X2 U14595 ( .I(n38630), .ZN(n35287) );
  NAND2_X2 U14596 ( .A1(n37827), .A2(n37826), .ZN(n38630) );
  OAI21_X2 U14598 ( .A1(n30699), .A2(n37737), .B(n2549), .ZN(n10894) );
  BUF_X2 U14599 ( .I(n28219), .Z(n37828) );
  NAND2_X2 U14600 ( .A1(n8817), .A2(n8814), .ZN(n13056) );
  INV_X2 U14605 ( .I(n32622), .ZN(n841) );
  NAND2_X2 U14608 ( .A1(n38397), .A2(n37220), .ZN(n11383) );
  AOI21_X1 U14609 ( .A1(n24467), .A2(n18345), .B(n37259), .ZN(n35774) );
  XOR2_X1 U14610 ( .A1(n37829), .A2(n16806), .Z(n16804) );
  XOR2_X1 U14611 ( .A1(n25113), .A2(n25189), .Z(n25208) );
  OAI22_X2 U14612 ( .A1(n14797), .A2(n14796), .B1(n37246), .B2(n14795), .ZN(
        n37881) );
  XOR2_X1 U14614 ( .A1(n11887), .A2(n11615), .Z(n9023) );
  XOR2_X1 U14615 ( .A1(n13617), .A2(n23903), .Z(n11887) );
  OAI22_X2 U14618 ( .A1(n36021), .A2(n33449), .B1(n37831), .B2(n37830), .ZN(
        n3649) );
  NOR2_X2 U14624 ( .A1(n24609), .A2(n39704), .ZN(n37831) );
  XOR2_X1 U14626 ( .A1(n25257), .A2(n37832), .Z(n25122) );
  XOR2_X1 U14635 ( .A1(n25224), .A2(n25116), .Z(n37832) );
  NOR2_X2 U14646 ( .A1(n24327), .A2(n2396), .ZN(n24175) );
  XOR2_X1 U14648 ( .A1(n37834), .A2(n2402), .Z(n39362) );
  NAND2_X2 U14649 ( .A1(n36945), .A2(n39670), .ZN(n37957) );
  NAND2_X2 U14650 ( .A1(n37835), .A2(n32999), .ZN(n26498) );
  NOR2_X1 U14651 ( .A1(n37893), .A2(n17954), .ZN(n37835) );
  NOR2_X2 U14655 ( .A1(n37836), .A2(n31074), .ZN(n16524) );
  NOR2_X2 U14656 ( .A1(n31951), .A2(n36888), .ZN(n37836) );
  NOR2_X2 U14657 ( .A1(n18540), .A2(n19227), .ZN(n10722) );
  INV_X2 U14660 ( .I(n39401), .ZN(n37839) );
  XOR2_X1 U14665 ( .A1(n16054), .A2(n38147), .Z(n34649) );
  AOI22_X2 U14666 ( .A1(n37733), .A2(n37841), .B1(n24314), .B2(n7883), .ZN(
        n8961) );
  NAND2_X2 U14667 ( .A1(n38366), .A2(n33077), .ZN(n37841) );
  INV_X4 U14668 ( .I(n12931), .ZN(n38338) );
  XOR2_X1 U14669 ( .A1(n35707), .A2(n33038), .Z(n828) );
  AOI21_X2 U14678 ( .A1(n11942), .A2(n3879), .B(n3878), .ZN(n35707) );
  OAI22_X2 U14679 ( .A1(n24755), .A2(n37852), .B1(n19420), .B2(n1577), .ZN(
        n17963) );
  NOR2_X2 U14684 ( .A1(n933), .A2(n36385), .ZN(n37852) );
  XOR2_X1 U14685 ( .A1(n23697), .A2(n31775), .Z(n23913) );
  NAND2_X2 U14686 ( .A1(n22825), .A2(n22824), .ZN(n23697) );
  XOR2_X1 U14687 ( .A1(n34440), .A2(n32646), .Z(n17651) );
  INV_X2 U14690 ( .I(n37843), .ZN(n35954) );
  XNOR2_X1 U14697 ( .A1(n12921), .A2(n12920), .ZN(n37843) );
  NAND2_X1 U14699 ( .A1(n22823), .A2(n1630), .ZN(n38266) );
  INV_X4 U14700 ( .I(n6945), .ZN(n13150) );
  XOR2_X1 U14704 ( .A1(n22669), .A2(n30406), .Z(n30898) );
  XOR2_X1 U14705 ( .A1(n18595), .A2(n22728), .Z(n22669) );
  NAND2_X2 U14710 ( .A1(n5330), .A2(n37846), .ZN(n7445) );
  NAND2_X2 U14711 ( .A1(n32322), .A2(n37847), .ZN(n37846) );
  NAND2_X2 U14712 ( .A1(n37849), .A2(n37848), .ZN(n37847) );
  INV_X2 U14713 ( .I(n1125), .ZN(n37848) );
  INV_X4 U14716 ( .I(n30059), .ZN(n1403) );
  XOR2_X1 U14717 ( .A1(n37850), .A2(n11976), .Z(n12187) );
  XOR2_X1 U14719 ( .A1(n27790), .A2(n27789), .Z(n37850) );
  XOR2_X1 U14720 ( .A1(n29039), .A2(n29108), .Z(n28895) );
  XOR2_X1 U14721 ( .A1(n973), .A2(n17039), .Z(n29108) );
  OAI21_X2 U14723 ( .A1(n37851), .A2(n23335), .B(n20421), .ZN(n19846) );
  XOR2_X1 U14733 ( .A1(n26376), .A2(n20425), .Z(n20424) );
  XOR2_X1 U14734 ( .A1(n33178), .A2(n2281), .Z(n19652) );
  NAND2_X2 U14735 ( .A1(n13196), .A2(n13194), .ZN(n11533) );
  NAND3_X2 U14737 ( .A1(n21501), .A2(n39705), .A3(n37853), .ZN(n22332) );
  NAND2_X1 U14738 ( .A1(n39627), .A2(n21499), .ZN(n37853) );
  NOR2_X2 U14740 ( .A1(n33561), .A2(n26818), .ZN(n39054) );
  XOR2_X1 U14741 ( .A1(n39058), .A2(n33486), .Z(n4599) );
  INV_X1 U14744 ( .I(n10213), .ZN(n34553) );
  XNOR2_X1 U14746 ( .A1(n19152), .A2(n10213), .ZN(n10939) );
  NOR2_X2 U14749 ( .A1(n39801), .A2(n4479), .ZN(n10213) );
  NAND2_X2 U14750 ( .A1(n1944), .A2(n28612), .ZN(n5928) );
  XOR2_X1 U14753 ( .A1(n32106), .A2(n26278), .Z(n7661) );
  NAND2_X2 U14761 ( .A1(n5101), .A2(n37854), .ZN(n38689) );
  INV_X4 U14763 ( .I(n34217), .ZN(n38953) );
  NOR2_X2 U14764 ( .A1(n28093), .A2(n9266), .ZN(n36643) );
  NAND2_X2 U14765 ( .A1(n26759), .A2(n12755), .ZN(n12767) );
  NOR2_X2 U14768 ( .A1(n37098), .A2(n37856), .ZN(n26759) );
  NOR2_X2 U14771 ( .A1(n19232), .A2(n34603), .ZN(n4149) );
  NAND2_X2 U14778 ( .A1(n21195), .A2(n37857), .ZN(n29336) );
  OR2_X2 U14781 ( .A1(n11657), .A2(n7923), .Z(n25625) );
  XOR2_X1 U14783 ( .A1(n27477), .A2(n35190), .Z(n37860) );
  XOR2_X1 U14785 ( .A1(n22710), .A2(n10558), .Z(n35835) );
  OR2_X1 U14787 ( .A1(n19142), .A2(n6402), .Z(n16902) );
  OAI21_X2 U14788 ( .A1(n31921), .A2(n5953), .B(n39413), .ZN(n24583) );
  XOR2_X1 U14790 ( .A1(n6559), .A2(n37861), .Z(n18080) );
  NOR2_X2 U14795 ( .A1(n31404), .A2(n37862), .ZN(n10343) );
  XOR2_X1 U14801 ( .A1(n11721), .A2(n3488), .Z(n39552) );
  INV_X4 U14802 ( .I(n21401), .ZN(n20037) );
  NAND2_X2 U14805 ( .A1(n36275), .A2(n37614), .ZN(n18216) );
  AOI21_X2 U14808 ( .A1(n5124), .A2(n37640), .B(n37475), .ZN(n6619) );
  BUF_X2 U14809 ( .I(n31664), .Z(n37863) );
  XOR2_X1 U14814 ( .A1(n3824), .A2(n37864), .Z(n38770) );
  XOR2_X1 U14816 ( .A1(n10083), .A2(n16368), .Z(n37864) );
  NOR2_X2 U14817 ( .A1(n34892), .A2(n3449), .ZN(n26952) );
  XOR2_X1 U14824 ( .A1(n37865), .A2(n26338), .Z(n38009) );
  XOR2_X1 U14827 ( .A1(n10965), .A2(n19681), .Z(n37865) );
  NAND3_X2 U14828 ( .A1(n34116), .A2(n1777), .A3(n1781), .ZN(n31565) );
  XOR2_X1 U14837 ( .A1(n18490), .A2(n29509), .Z(n20956) );
  NAND3_X2 U14838 ( .A1(n18745), .A2(n25896), .A3(n34565), .ZN(n18490) );
  NAND3_X2 U14840 ( .A1(n35398), .A2(n35397), .A3(n5839), .ZN(n23714) );
  INV_X1 U14843 ( .I(n8080), .ZN(n16115) );
  NOR2_X1 U14847 ( .A1(n37867), .A2(n37866), .ZN(n11650) );
  INV_X1 U14848 ( .I(n20632), .ZN(n37866) );
  NAND2_X1 U14849 ( .A1(n20774), .A2(n8080), .ZN(n37867) );
  XOR2_X1 U14851 ( .A1(n7864), .A2(n7865), .Z(n8080) );
  NAND2_X2 U14852 ( .A1(n5231), .A2(n37868), .ZN(n12324) );
  NAND2_X1 U14853 ( .A1(n39075), .A2(n37226), .ZN(n37868) );
  NAND3_X2 U14854 ( .A1(n27381), .A2(n27382), .A3(n32913), .ZN(n4934) );
  NOR2_X2 U14857 ( .A1(n1962), .A2(n33964), .ZN(n2456) );
  XOR2_X1 U14860 ( .A1(n37870), .A2(n37869), .Z(n37929) );
  XOR2_X1 U14863 ( .A1(n32972), .A2(n11437), .Z(n37870) );
  INV_X4 U14866 ( .I(n35932), .ZN(n23505) );
  XOR2_X1 U14868 ( .A1(n26432), .A2(n32095), .Z(n26454) );
  NAND2_X2 U14869 ( .A1(n11270), .A2(n11269), .ZN(n26432) );
  NAND2_X2 U14871 ( .A1(n18729), .A2(n37871), .ZN(n11974) );
  AOI22_X2 U14875 ( .A1(n18728), .A2(n36237), .B1(n22229), .B2(n22230), .ZN(
        n37871) );
  NOR2_X1 U14877 ( .A1(n30629), .A2(n36404), .ZN(n8377) );
  OAI21_X2 U14882 ( .A1(n28594), .A2(n31088), .B(n37872), .ZN(n6810) );
  NAND2_X2 U14883 ( .A1(n28700), .A2(n38669), .ZN(n37872) );
  XOR2_X1 U14887 ( .A1(n22500), .A2(n22509), .Z(n22635) );
  NAND2_X2 U14890 ( .A1(n39275), .A2(n19284), .ZN(n22500) );
  XOR2_X1 U14891 ( .A1(n10658), .A2(n35027), .Z(n7666) );
  XOR2_X1 U14895 ( .A1(n15157), .A2(n28943), .Z(n3126) );
  NAND3_X2 U14899 ( .A1(n16183), .A2(n3128), .A3(n28709), .ZN(n15157) );
  AND2_X1 U14901 ( .A1(n3850), .A2(n1890), .Z(n38910) );
  NAND2_X1 U14902 ( .A1(n38345), .A2(n8085), .ZN(n34891) );
  NAND2_X2 U14905 ( .A1(n31364), .A2(n11588), .ZN(n7225) );
  XOR2_X1 U14907 ( .A1(n4366), .A2(n38816), .Z(n16085) );
  NOR2_X1 U14909 ( .A1(n2500), .A2(n28442), .ZN(n14002) );
  NAND2_X2 U14913 ( .A1(n14660), .A2(n37873), .ZN(n26223) );
  AOI22_X2 U14923 ( .A1(n11633), .A2(n31133), .B1(n7732), .B2(n1018), .ZN(
        n37873) );
  OAI21_X2 U14926 ( .A1(n34601), .A2(n37875), .B(n5263), .ZN(n1788) );
  NOR2_X2 U14934 ( .A1(n32256), .A2(n2735), .ZN(n37875) );
  OAI21_X2 U14936 ( .A1(n12926), .A2(n15755), .B(n33944), .ZN(n36016) );
  NAND2_X2 U14939 ( .A1(n20572), .A2(n38365), .ZN(n28285) );
  INV_X1 U14941 ( .I(n9956), .ZN(n38414) );
  NAND2_X2 U14943 ( .A1(n11736), .A2(n33417), .ZN(n19061) );
  NOR2_X2 U14944 ( .A1(n14201), .A2(n32917), .ZN(n33417) );
  XOR2_X1 U14945 ( .A1(n37876), .A2(n37240), .Z(n34610) );
  XOR2_X1 U14946 ( .A1(n27635), .A2(n379), .Z(n37876) );
  XOR2_X1 U14949 ( .A1(n22600), .A2(n22561), .Z(n22609) );
  AOI22_X2 U14950 ( .A1(n9523), .A2(n22239), .B1(n16888), .B2(n9521), .ZN(
        n22600) );
  NOR2_X1 U14951 ( .A1(n32594), .A2(n38611), .ZN(n38892) );
  XOR2_X1 U14962 ( .A1(n37877), .A2(n4064), .Z(n8057) );
  XOR2_X1 U14963 ( .A1(n27459), .A2(n38121), .Z(n37877) );
  NAND2_X2 U14964 ( .A1(n7), .A2(n39036), .ZN(n31767) );
  NAND2_X2 U14967 ( .A1(n29644), .A2(n37878), .ZN(n33643) );
  NAND2_X2 U14969 ( .A1(n29643), .A2(n37879), .ZN(n37878) );
  NAND2_X2 U14971 ( .A1(n33630), .A2(n25907), .ZN(n26402) );
  NAND2_X2 U14974 ( .A1(n32574), .A2(n32573), .ZN(n15202) );
  NOR2_X1 U14978 ( .A1(n15174), .A2(n29551), .ZN(n21177) );
  BUF_X2 U14981 ( .I(n33047), .Z(n37880) );
  OR2_X2 U14984 ( .A1(n14383), .A2(n860), .Z(n26946) );
  INV_X4 U14987 ( .I(n17887), .ZN(n6514) );
  NAND2_X2 U14989 ( .A1(n3545), .A2(n3544), .ZN(n17887) );
  NAND2_X1 U14990 ( .A1(n11521), .A2(n8194), .ZN(n36584) );
  XOR2_X1 U14994 ( .A1(n38180), .A2(n37882), .Z(n751) );
  NOR2_X2 U14998 ( .A1(n12456), .A2(n12458), .ZN(n38180) );
  XOR2_X1 U15000 ( .A1(n24926), .A2(n25181), .Z(n6352) );
  NOR2_X2 U15007 ( .A1(n7350), .A2(n12643), .ZN(n24926) );
  XOR2_X1 U15010 ( .A1(n5473), .A2(n5472), .Z(n5518) );
  AOI22_X2 U15011 ( .A1(n31030), .A2(n28463), .B1(n34312), .B2(n30757), .ZN(
        n28791) );
  NAND2_X2 U15012 ( .A1(n33022), .A2(n19452), .ZN(n25697) );
  XOR2_X1 U15013 ( .A1(n11189), .A2(n37094), .Z(n11192) );
  XOR2_X1 U15015 ( .A1(n37884), .A2(n20536), .Z(n11188) );
  XOR2_X1 U15018 ( .A1(n5553), .A2(n39512), .Z(n37884) );
  NAND2_X2 U15019 ( .A1(n11669), .A2(n7577), .ZN(n32832) );
  OAI22_X2 U15022 ( .A1(n30145), .A2(n35234), .B1(n18241), .B2(n30132), .ZN(
        n29015) );
  NAND2_X2 U15024 ( .A1(n7366), .A2(n22896), .ZN(n23456) );
  NOR2_X1 U15033 ( .A1(n3356), .A2(n1106), .ZN(n3360) );
  NOR2_X2 U15035 ( .A1(n37120), .A2(n37885), .ZN(n36705) );
  NOR2_X1 U15036 ( .A1(n274), .A2(n28150), .ZN(n37885) );
  NOR2_X1 U15037 ( .A1(n28616), .A2(n180), .ZN(n28454) );
  NAND2_X2 U15040 ( .A1(n34871), .A2(n14330), .ZN(n180) );
  NAND2_X2 U15041 ( .A1(n38957), .A2(n28170), .ZN(n28676) );
  XOR2_X1 U15044 ( .A1(n28891), .A2(n6433), .Z(n29159) );
  NAND3_X2 U15047 ( .A1(n15630), .A2(n28678), .A3(n15629), .ZN(n6433) );
  NAND2_X2 U15053 ( .A1(n1445), .A2(n34166), .ZN(n38743) );
  AOI21_X2 U15057 ( .A1(n16353), .A2(n30057), .B(n30059), .ZN(n3045) );
  XOR2_X1 U15060 ( .A1(n4413), .A2(n22741), .Z(n7358) );
  NAND2_X2 U15064 ( .A1(n35727), .A2(n20123), .ZN(n4413) );
  INV_X2 U15068 ( .I(n26255), .ZN(n1505) );
  NAND3_X2 U15071 ( .A1(n38866), .A2(n30468), .A3(n16612), .ZN(n26255) );
  AOI21_X2 U15073 ( .A1(n15790), .A2(n15791), .B(n15789), .ZN(n12548) );
  OAI21_X2 U15078 ( .A1(n38387), .A2(n9888), .B(n37886), .ZN(n7852) );
  NAND2_X1 U15080 ( .A1(n37887), .A2(n2597), .ZN(n37886) );
  NOR2_X1 U15082 ( .A1(n15049), .A2(n38702), .ZN(n37887) );
  XOR2_X1 U15083 ( .A1(n14136), .A2(n37888), .Z(n16907) );
  XOR2_X1 U15085 ( .A1(n29055), .A2(n29056), .Z(n37888) );
  NAND2_X1 U15086 ( .A1(n29265), .A2(n1406), .ZN(n37942) );
  XOR2_X1 U15091 ( .A1(n16610), .A2(n29432), .Z(n37889) );
  XOR2_X1 U15094 ( .A1(n15916), .A2(n16324), .Z(n23954) );
  AOI21_X2 U15097 ( .A1(n15799), .A2(n18762), .B(n15949), .ZN(n15916) );
  NOR2_X1 U15098 ( .A1(n17692), .A2(n17691), .ZN(n39645) );
  NAND3_X1 U15107 ( .A1(n6487), .A2(n3947), .A3(n6486), .ZN(n32460) );
  AOI22_X2 U15114 ( .A1(n31498), .A2(n9295), .B1(n27374), .B2(n27266), .ZN(
        n27749) );
  XOR2_X1 U15120 ( .A1(n3889), .A2(n27677), .Z(n3886) );
  NAND3_X1 U15121 ( .A1(n13191), .A2(n36371), .A3(n2654), .ZN(n11455) );
  BUF_X4 U15122 ( .I(n1033), .Z(n39156) );
  NAND2_X2 U15124 ( .A1(n17227), .A2(n27046), .ZN(n18195) );
  AOI22_X2 U15125 ( .A1(n34170), .A2(n19946), .B1(n37186), .B2(n28131), .ZN(
        n37892) );
  OAI21_X2 U15129 ( .A1(n37167), .A2(n23127), .B(n34124), .ZN(n9862) );
  NAND2_X2 U15133 ( .A1(n1302), .A2(n5487), .ZN(n18312) );
  NAND2_X1 U15134 ( .A1(n26902), .A2(n19673), .ZN(n37900) );
  NAND2_X1 U15135 ( .A1(n37077), .A2(n27018), .ZN(n39503) );
  OAI21_X2 U15137 ( .A1(n13261), .A2(n29377), .B(n29453), .ZN(n29379) );
  XOR2_X1 U15139 ( .A1(n13703), .A2(n27631), .Z(n31731) );
  AOI21_X2 U15142 ( .A1(n30678), .A2(n4231), .B(n30416), .ZN(n27631) );
  XOR2_X1 U15144 ( .A1(n26571), .A2(n12838), .Z(n26197) );
  NOR2_X2 U15147 ( .A1(n18631), .A2(n18630), .ZN(n12838) );
  AND2_X1 U15148 ( .A1(n32377), .A2(n6945), .Z(n13830) );
  XOR2_X1 U15149 ( .A1(n32660), .A2(n30976), .Z(n37934) );
  BUF_X4 U15153 ( .I(n26556), .Z(n11667) );
  NOR2_X1 U15155 ( .A1(n36352), .A2(n3013), .ZN(n37893) );
  NAND2_X2 U15156 ( .A1(n37894), .A2(n39566), .ZN(n27858) );
  NAND2_X1 U15158 ( .A1(n17718), .A2(n17719), .ZN(n37894) );
  XOR2_X1 U15162 ( .A1(n25318), .A2(n25320), .Z(n12330) );
  NAND2_X2 U15166 ( .A1(n33043), .A2(n2530), .ZN(n25318) );
  NAND2_X2 U15174 ( .A1(n13782), .A2(n30766), .ZN(n30845) );
  XOR2_X1 U15175 ( .A1(n24036), .A2(n18849), .Z(n23756) );
  OAI22_X2 U15176 ( .A1(n21040), .A2(n17458), .B1(n15524), .B2(n4382), .ZN(
        n11668) );
  OR2_X1 U15177 ( .A1(n23198), .A2(n32856), .Z(n8462) );
  NAND3_X1 U15179 ( .A1(n9107), .A2(n9878), .A3(n37619), .ZN(n37897) );
  OAI22_X2 U15183 ( .A1(n22275), .A2(n35771), .B1(n16772), .B2(n14196), .ZN(
        n13785) );
  BUF_X2 U15194 ( .I(n32535), .Z(n37898) );
  AOI21_X1 U15195 ( .A1(n34299), .A2(n8988), .B(n35767), .ZN(n6383) );
  INV_X2 U15197 ( .I(n19477), .ZN(n35767) );
  NAND2_X2 U15202 ( .A1(n11514), .A2(n11516), .ZN(n19477) );
  OAI21_X2 U15204 ( .A1(n10753), .A2(n31780), .B(n1548), .ZN(n32481) );
  INV_X2 U15207 ( .I(n26808), .ZN(n26810) );
  XOR2_X1 U15208 ( .A1(n6033), .A2(n29666), .Z(n13229) );
  NAND2_X2 U15213 ( .A1(n38318), .A2(n13231), .ZN(n6033) );
  NOR2_X1 U15214 ( .A1(n35264), .A2(n36910), .ZN(n36976) );
  INV_X4 U15215 ( .I(n16559), .ZN(n19893) );
  AOI22_X2 U15216 ( .A1(n7945), .A2(n1072), .B1(n6788), .B2(n7946), .ZN(n7324)
         );
  XOR2_X1 U15217 ( .A1(n8897), .A2(n33133), .Z(n10009) );
  AND2_X1 U15221 ( .A1(n32566), .A2(n33593), .Z(n3690) );
  NAND2_X2 U15227 ( .A1(n3102), .A2(n8685), .ZN(n32566) );
  NAND2_X2 U15228 ( .A1(n16182), .A2(n23482), .ZN(n38691) );
  NAND2_X2 U15229 ( .A1(n19414), .A2(n14632), .ZN(n9686) );
  XOR2_X1 U15231 ( .A1(n38815), .A2(n38814), .Z(n13872) );
  NAND2_X2 U15234 ( .A1(n31079), .A2(n15534), .ZN(n39163) );
  NOR2_X2 U15235 ( .A1(n37900), .A2(n35311), .ZN(n9956) );
  NAND2_X1 U15236 ( .A1(n39569), .A2(n929), .ZN(n4512) );
  NAND2_X2 U15241 ( .A1(n8843), .A2(n15365), .ZN(n31679) );
  OAI21_X2 U15243 ( .A1(n38527), .A2(n38528), .B(n35761), .ZN(n8843) );
  INV_X2 U15246 ( .I(n28758), .ZN(n1426) );
  OR2_X1 U15247 ( .A1(n28758), .A2(n20597), .Z(n8850) );
  INV_X4 U15249 ( .I(n9855), .ZN(n11807) );
  NAND2_X2 U15250 ( .A1(n32826), .A2(n32827), .ZN(n9855) );
  NAND2_X2 U15251 ( .A1(n36374), .A2(n37901), .ZN(n32854) );
  NAND3_X2 U15255 ( .A1(n13585), .A2(n25762), .A3(n25761), .ZN(n19450) );
  OAI22_X2 U15256 ( .A1(n548), .A2(n33401), .B1(n1119), .B2(n18858), .ZN(
        n13637) );
  AOI22_X2 U15259 ( .A1(n17754), .A2(n27235), .B1(n36234), .B2(n27233), .ZN(
        n35902) );
  XOR2_X1 U15260 ( .A1(n26411), .A2(n16216), .Z(n14770) );
  XOR2_X1 U15261 ( .A1(n26532), .A2(n26591), .Z(n26411) );
  XOR2_X1 U15265 ( .A1(n34800), .A2(n33364), .Z(n3771) );
  XOR2_X1 U15266 ( .A1(n828), .A2(n25191), .Z(n15686) );
  XOR2_X1 U15267 ( .A1(n140), .A2(n36363), .Z(n34213) );
  XOR2_X1 U15271 ( .A1(n29126), .A2(n2142), .Z(n2005) );
  AND2_X1 U15272 ( .A1(n23613), .A2(n1627), .Z(n32294) );
  NAND2_X1 U15276 ( .A1(n30453), .A2(n33356), .ZN(n35018) );
  OAI21_X1 U15278 ( .A1(n39806), .A2(n2830), .B(n32193), .ZN(n1743) );
  NAND2_X2 U15280 ( .A1(n15579), .A2(n23237), .ZN(n23459) );
  NOR2_X2 U15284 ( .A1(n327), .A2(n32850), .ZN(n15579) );
  XOR2_X1 U15285 ( .A1(n23794), .A2(n23671), .Z(n17398) );
  NAND2_X2 U15287 ( .A1(n6141), .A2(n6139), .ZN(n23671) );
  NOR2_X1 U15291 ( .A1(n39510), .A2(n37902), .ZN(n38462) );
  OAI22_X1 U15292 ( .A1(n18424), .A2(n30144), .B1(n30143), .B2(n18588), .ZN(
        n37902) );
  OAI21_X2 U15293 ( .A1(n37981), .A2(n37880), .B(n4369), .ZN(n38504) );
  XOR2_X1 U15295 ( .A1(n32239), .A2(n17463), .Z(n8299) );
  NAND2_X2 U15297 ( .A1(n36429), .A2(n3031), .ZN(n32239) );
  NAND2_X1 U15298 ( .A1(n15575), .A2(n18827), .ZN(n25866) );
  NAND2_X2 U15301 ( .A1(n32658), .A2(n17740), .ZN(n15575) );
  XOR2_X1 U15304 ( .A1(n15676), .A2(n35240), .Z(n36383) );
  INV_X2 U15306 ( .I(n17989), .ZN(n14024) );
  NAND2_X1 U15313 ( .A1(n20555), .A2(n35687), .ZN(n22809) );
  INV_X4 U15315 ( .I(n23198), .ZN(n38283) );
  BUF_X2 U15321 ( .I(n2576), .Z(n37905) );
  NOR2_X2 U15327 ( .A1(n39584), .A2(n34399), .ZN(n38956) );
  XOR2_X1 U15328 ( .A1(n31633), .A2(n17581), .Z(n12138) );
  NAND2_X2 U15330 ( .A1(n1177), .A2(n1399), .ZN(n12955) );
  OAI22_X2 U15334 ( .A1(n37906), .A2(n23416), .B1(n23418), .B2(n36130), .ZN(
        n3521) );
  XOR2_X1 U15339 ( .A1(n23677), .A2(n23947), .Z(n1791) );
  NAND2_X1 U15341 ( .A1(n15223), .A2(n16430), .ZN(n38182) );
  NAND2_X2 U15343 ( .A1(n5146), .A2(n39174), .ZN(n5171) );
  NOR2_X2 U15346 ( .A1(n7170), .A2(n37907), .ZN(n7168) );
  NOR2_X2 U15347 ( .A1(n8120), .A2(n11807), .ZN(n37907) );
  XOR2_X1 U15348 ( .A1(n13531), .A2(n25316), .Z(n39315) );
  XOR2_X1 U15356 ( .A1(n4592), .A2(n32190), .Z(n18655) );
  INV_X2 U15357 ( .I(n29803), .ZN(n966) );
  INV_X2 U15363 ( .I(n5869), .ZN(n4411) );
  XOR2_X1 U15370 ( .A1(n5312), .A2(n32915), .Z(n5869) );
  NAND3_X2 U15372 ( .A1(n8041), .A2(n18721), .A3(n8042), .ZN(n33102) );
  XOR2_X1 U15376 ( .A1(n27642), .A2(n27861), .Z(n17276) );
  XOR2_X1 U15378 ( .A1(n27828), .A2(n27766), .Z(n27861) );
  XOR2_X1 U15380 ( .A1(n37908), .A2(n13172), .Z(n23132) );
  XOR2_X1 U15382 ( .A1(n13174), .A2(n22658), .Z(n37908) );
  XOR2_X1 U15385 ( .A1(n17612), .A2(n37909), .Z(n32662) );
  XOR2_X1 U15386 ( .A1(n2585), .A2(n963), .Z(n37909) );
  XOR2_X1 U15387 ( .A1(n29297), .A2(n28967), .Z(n29033) );
  XOR2_X1 U15392 ( .A1(n7848), .A2(n29166), .Z(n29297) );
  XOR2_X1 U15396 ( .A1(n16709), .A2(n37910), .Z(n6848) );
  XOR2_X1 U15397 ( .A1(n282), .A2(n27825), .Z(n37910) );
  NAND2_X2 U15398 ( .A1(n15701), .A2(n15775), .ZN(n13386) );
  XOR2_X1 U15402 ( .A1(n22703), .A2(n17756), .Z(n18001) );
  NAND2_X2 U15403 ( .A1(n21452), .A2(n21453), .ZN(n22703) );
  XOR2_X1 U15404 ( .A1(n12570), .A2(n37912), .Z(n12200) );
  XOR2_X1 U15407 ( .A1(n20509), .A2(n23894), .Z(n12570) );
  INV_X1 U15408 ( .I(n24039), .ZN(n37912) );
  OR2_X1 U15415 ( .A1(n24271), .A2(n18342), .Z(n38115) );
  NAND2_X2 U15416 ( .A1(n37970), .A2(n37913), .ZN(n23251) );
  AND2_X1 U15420 ( .A1(n2840), .A2(n22042), .Z(n10623) );
  NOR2_X2 U15429 ( .A1(n7636), .A2(n37920), .ZN(n37919) );
  INV_X2 U15437 ( .I(n18253), .ZN(n37920) );
  NOR2_X2 U15441 ( .A1(n18637), .A2(n23060), .ZN(n18636) );
  NAND2_X2 U15446 ( .A1(n37922), .A2(n37921), .ZN(n18637) );
  INV_X1 U15448 ( .I(n18209), .ZN(n37921) );
  XOR2_X1 U15454 ( .A1(n15532), .A2(n23971), .Z(n20615) );
  AOI21_X2 U15460 ( .A1(n28216), .A2(n28219), .B(n28217), .ZN(n16467) );
  NAND2_X2 U15461 ( .A1(n987), .A2(n16631), .ZN(n28219) );
  NOR2_X2 U15462 ( .A1(n23522), .A2(n3708), .ZN(n23318) );
  AOI21_X1 U15464 ( .A1(n16869), .A2(n33510), .B(n28214), .ZN(n16868) );
  XOR2_X1 U15467 ( .A1(n4136), .A2(n13939), .Z(n4135) );
  NAND2_X2 U15471 ( .A1(n11491), .A2(n11492), .ZN(n31515) );
  XOR2_X1 U15478 ( .A1(n28500), .A2(n28886), .Z(n29105) );
  OAI21_X2 U15480 ( .A1(n3877), .A2(n8878), .B(n37925), .ZN(n3874) );
  OAI21_X2 U15481 ( .A1(n15620), .A2(n34060), .B(n10882), .ZN(n37925) );
  BUF_X2 U15483 ( .I(n31305), .Z(n37926) );
  XOR2_X1 U15484 ( .A1(n37247), .A2(n6134), .Z(n38467) );
  XOR2_X1 U15486 ( .A1(n11319), .A2(n15930), .Z(n6458) );
  AND2_X2 U15488 ( .A1(n8479), .A2(n35476), .Z(n26805) );
  XOR2_X1 U15492 ( .A1(n3320), .A2(n27475), .Z(n18846) );
  XOR2_X1 U15493 ( .A1(n7910), .A2(n16162), .Z(n27475) );
  NOR3_X1 U15495 ( .A1(n26220), .A2(n2000), .A3(n26839), .ZN(n16298) );
  OAI22_X1 U15496 ( .A1(n29276), .A2(n17773), .B1(n13886), .B2(n29275), .ZN(
        n5088) );
  NAND2_X2 U15500 ( .A1(n7088), .A2(n29125), .ZN(n33833) );
  NAND2_X2 U15501 ( .A1(n37248), .A2(n13823), .ZN(n29125) );
  NAND3_X2 U15502 ( .A1(n37927), .A2(n38062), .A3(n38061), .ZN(n29057) );
  XOR2_X1 U15505 ( .A1(n8003), .A2(n37928), .Z(n135) );
  XOR2_X1 U15508 ( .A1(n16673), .A2(n25225), .Z(n37928) );
  AOI21_X2 U15509 ( .A1(n37890), .A2(n27372), .B(n16042), .ZN(n13526) );
  INV_X2 U15511 ( .I(n16040), .ZN(n16042) );
  NOR2_X2 U15513 ( .A1(n17795), .A2(n27123), .ZN(n16040) );
  NOR2_X2 U15515 ( .A1(n20035), .A2(n31798), .ZN(n23590) );
  NAND2_X1 U15519 ( .A1(n4190), .A2(n10834), .ZN(n26012) );
  NAND2_X2 U15521 ( .A1(n4018), .A2(n9335), .ZN(n4190) );
  INV_X2 U15523 ( .I(n37929), .ZN(n33972) );
  XOR2_X1 U15524 ( .A1(n5289), .A2(n15960), .Z(n5320) );
  NAND2_X2 U15528 ( .A1(n5287), .A2(n33190), .ZN(n5289) );
  NAND2_X2 U15529 ( .A1(n7892), .A2(n14869), .ZN(n16548) );
  NAND3_X1 U15530 ( .A1(n24806), .A2(n1026), .A3(n19565), .ZN(n37931) );
  INV_X2 U15531 ( .I(n18035), .ZN(n28425) );
  BUF_X4 U15534 ( .I(n21660), .Z(n39627) );
  NOR2_X2 U15535 ( .A1(n209), .A2(n1424), .ZN(n12398) );
  NAND2_X2 U15536 ( .A1(n14107), .A2(n23252), .ZN(n23890) );
  INV_X2 U15540 ( .I(n32239), .ZN(n37932) );
  XOR2_X1 U15545 ( .A1(n25204), .A2(n25114), .Z(n15758) );
  NOR2_X2 U15550 ( .A1(n13637), .A2(n13638), .ZN(n25204) );
  XOR2_X1 U15552 ( .A1(n5761), .A2(n5760), .Z(n12758) );
  NAND2_X2 U15556 ( .A1(n31862), .A2(n32607), .ZN(n27383) );
  NAND2_X2 U15558 ( .A1(n37933), .A2(n39734), .ZN(n10118) );
  NAND3_X2 U15559 ( .A1(n39416), .A2(n3958), .A3(n38883), .ZN(n37933) );
  NAND2_X2 U15561 ( .A1(n39216), .A2(n20671), .ZN(n27205) );
  NOR2_X2 U15568 ( .A1(n27139), .A2(n27140), .ZN(n27197) );
  OAI22_X2 U15570 ( .A1(n19433), .A2(n26692), .B1(n26691), .B2(n39825), .ZN(
        n27139) );
  XOR2_X1 U15571 ( .A1(n37935), .A2(n19815), .Z(Ciphertext[151]) );
  OAI22_X1 U15574 ( .A1(n28658), .A2(n28657), .B1(n17977), .B2(n1197), .ZN(
        n31705) );
  NAND3_X2 U15579 ( .A1(n2338), .A2(n20184), .A3(n16154), .ZN(n2023) );
  XOR2_X1 U15580 ( .A1(n4282), .A2(n38659), .Z(n16931) );
  NAND2_X1 U15582 ( .A1(n36060), .A2(n36059), .ZN(n39388) );
  OAI21_X2 U15583 ( .A1(n29867), .A2(n29843), .B(n29869), .ZN(n20894) );
  XOR2_X1 U15589 ( .A1(n1503), .A2(n26584), .Z(n26482) );
  NAND3_X2 U15591 ( .A1(n13103), .A2(n25827), .A3(n25828), .ZN(n26584) );
  INV_X2 U15593 ( .I(n37937), .ZN(n26249) );
  XNOR2_X1 U15597 ( .A1(n2069), .A2(n2066), .ZN(n37937) );
  OAI22_X2 U15601 ( .A1(n20370), .A2(n29629), .B1(n20371), .B2(n13441), .ZN(
        n20369) );
  CLKBUF_X4 U15607 ( .I(n33424), .Z(n38275) );
  INV_X1 U15608 ( .I(n21790), .ZN(n37939) );
  XNOR2_X1 U15616 ( .A1(n17804), .A2(n8796), .ZN(n38558) );
  NAND2_X2 U15617 ( .A1(n38737), .A2(n29103), .ZN(n29236) );
  NAND2_X2 U15619 ( .A1(n38034), .A2(n33102), .ZN(n38918) );
  INV_X1 U15622 ( .I(n9935), .ZN(n37940) );
  NAND2_X1 U15623 ( .A1(n37940), .A2(n36076), .ZN(n5642) );
  XOR2_X1 U15624 ( .A1(n17957), .A2(n37941), .Z(n10812) );
  XOR2_X1 U15628 ( .A1(n3223), .A2(n29050), .Z(n37941) );
  OR2_X1 U15632 ( .A1(n26029), .A2(n18320), .Z(n25804) );
  NAND2_X2 U15634 ( .A1(n8407), .A2(n26041), .ZN(n25825) );
  NAND2_X2 U15635 ( .A1(n25814), .A2(n25813), .ZN(n26023) );
  NAND3_X1 U15636 ( .A1(n29278), .A2(n29284), .A3(n1379), .ZN(n29279) );
  INV_X2 U15648 ( .I(n19518), .ZN(n35618) );
  NAND3_X2 U15652 ( .A1(n5024), .A2(n5023), .A3(n13438), .ZN(n19518) );
  NAND2_X1 U15655 ( .A1(n7305), .A2(n19465), .ZN(n14427) );
  XOR2_X1 U15656 ( .A1(n3703), .A2(n3668), .Z(n31725) );
  XOR2_X1 U15658 ( .A1(n15013), .A2(n22664), .Z(n15012) );
  XOR2_X1 U15659 ( .A1(n37944), .A2(n3404), .Z(n18860) );
  XOR2_X1 U15672 ( .A1(n27765), .A2(n37991), .Z(n37944) );
  XOR2_X1 U15673 ( .A1(n20303), .A2(n24949), .Z(n25158) );
  XOR2_X1 U15674 ( .A1(n20304), .A2(n24946), .Z(n20303) );
  XOR2_X1 U15679 ( .A1(n35243), .A2(n20483), .Z(n38069) );
  NAND2_X2 U15684 ( .A1(n24875), .A2(n1580), .ZN(n9213) );
  XOR2_X1 U15686 ( .A1(n37945), .A2(n29411), .Z(Ciphertext[40]) );
  NAND3_X2 U15691 ( .A1(n7733), .A2(n15042), .A3(n14517), .ZN(n37945) );
  INV_X2 U15693 ( .I(n25177), .ZN(n1557) );
  NAND2_X2 U15695 ( .A1(n32268), .A2(n24871), .ZN(n25177) );
  AOI21_X2 U15698 ( .A1(n11094), .A2(n28772), .B(n37946), .ZN(n11389) );
  NOR3_X2 U15703 ( .A1(n5662), .A2(n31418), .A3(n10618), .ZN(n37946) );
  XOR2_X1 U15704 ( .A1(n17250), .A2(n37947), .Z(n5317) );
  XOR2_X1 U15705 ( .A1(n31550), .A2(n29070), .Z(n37947) );
  NAND3_X2 U15711 ( .A1(n8769), .A2(n38001), .A3(n2771), .ZN(n37948) );
  AND2_X1 U15712 ( .A1(n12682), .A2(n3873), .Z(n2735) );
  NAND2_X2 U15713 ( .A1(n37950), .A2(n14192), .ZN(n35151) );
  AND2_X1 U15714 ( .A1(n14262), .A2(n25643), .Z(n37950) );
  NOR2_X2 U15719 ( .A1(n6127), .A2(n15268), .ZN(n12628) );
  NAND2_X1 U15721 ( .A1(n32418), .A2(n18529), .ZN(n27873) );
  AOI21_X2 U15722 ( .A1(n36269), .A2(n37368), .B(n3045), .ZN(n3600) );
  XNOR2_X1 U15728 ( .A1(n27516), .A2(n27566), .ZN(n13883) );
  XOR2_X1 U15732 ( .A1(n37952), .A2(n20420), .Z(Ciphertext[117]) );
  BUF_X4 U15733 ( .I(n16040), .Z(n1475) );
  XOR2_X1 U15734 ( .A1(n11739), .A2(n19851), .Z(n6746) );
  NAND2_X2 U15736 ( .A1(n3348), .A2(n430), .ZN(n11739) );
  NOR2_X2 U15737 ( .A1(n39235), .A2(n17770), .ZN(n34446) );
  NAND2_X2 U15748 ( .A1(n9514), .A2(n7904), .ZN(n17770) );
  INV_X2 U15749 ( .I(n26015), .ZN(n26120) );
  OAI22_X2 U15750 ( .A1(n15254), .A2(n25501), .B1(n15647), .B2(n37183), .ZN(
        n26015) );
  XOR2_X1 U15759 ( .A1(n37953), .A2(n28793), .Z(n28796) );
  XOR2_X1 U15760 ( .A1(n29260), .A2(n36990), .Z(n37953) );
  OR2_X1 U15766 ( .A1(n686), .A2(n21912), .Z(n3692) );
  OR2_X1 U15767 ( .A1(n39444), .A2(n19223), .Z(n25502) );
  XOR2_X1 U15771 ( .A1(n27749), .A2(n27537), .Z(n27665) );
  NOR2_X2 U15773 ( .A1(n38860), .A2(n36791), .ZN(n31371) );
  XOR2_X1 U15782 ( .A1(n28873), .A2(n10430), .Z(n13315) );
  XNOR2_X1 U15785 ( .A1(n25170), .A2(n25285), .ZN(n31445) );
  XOR2_X1 U15791 ( .A1(n25284), .A2(n9701), .Z(n25170) );
  NAND2_X2 U15792 ( .A1(n12733), .A2(n37954), .ZN(n30379) );
  INV_X2 U15793 ( .I(n2394), .ZN(n37954) );
  XOR2_X1 U15799 ( .A1(n35177), .A2(n38964), .Z(n10866) );
  NAND2_X2 U15803 ( .A1(n36639), .A2(n35603), .ZN(n35177) );
  INV_X2 U15805 ( .I(n26946), .ZN(n14135) );
  XOR2_X1 U15806 ( .A1(n6774), .A2(n15782), .Z(n29943) );
  XOR2_X1 U15807 ( .A1(n15930), .A2(n17078), .Z(n13763) );
  AOI22_X2 U15809 ( .A1(n38424), .A2(n33705), .B1(n21028), .B2(n24750), .ZN(
        n15930) );
  AND2_X1 U15811 ( .A1(n15049), .A2(n2597), .Z(n36621) );
  NOR2_X2 U15812 ( .A1(n10883), .A2(n28685), .ZN(n9935) );
  INV_X4 U15813 ( .I(n7291), .ZN(n38305) );
  NAND2_X2 U15814 ( .A1(n32206), .A2(n5665), .ZN(n10883) );
  NAND2_X2 U15815 ( .A1(n1441), .A2(n1438), .ZN(n37960) );
  NAND2_X2 U15817 ( .A1(n33713), .A2(n31202), .ZN(n22293) );
  NAND2_X2 U15818 ( .A1(n3323), .A2(n3327), .ZN(n20397) );
  XOR2_X1 U15819 ( .A1(n26313), .A2(n26312), .Z(n26809) );
  XOR2_X1 U15821 ( .A1(n34686), .A2(n13608), .Z(n13787) );
  AND2_X2 U15826 ( .A1(n37961), .A2(n7245), .Z(n7250) );
  OAI21_X1 U15827 ( .A1(n3374), .A2(n16745), .B(n7044), .ZN(n37961) );
  NAND3_X2 U15835 ( .A1(n19575), .A2(n26946), .A3(n26857), .ZN(n36942) );
  NAND2_X2 U15836 ( .A1(n23767), .A2(n23796), .ZN(n33987) );
  AOI21_X2 U15839 ( .A1(n37962), .A2(n4298), .B(n9040), .ZN(n4297) );
  OAI21_X2 U15840 ( .A1(n19545), .A2(n21804), .B(n36735), .ZN(n37963) );
  NAND2_X2 U15845 ( .A1(n12620), .A2(n12618), .ZN(n12617) );
  NAND2_X2 U15850 ( .A1(n7008), .A2(n35232), .ZN(n21213) );
  NOR2_X1 U15851 ( .A1(n24829), .A2(n20128), .ZN(n15688) );
  NAND2_X2 U15852 ( .A1(n24625), .A2(n10421), .ZN(n20128) );
  XOR2_X1 U15854 ( .A1(n37964), .A2(n13313), .Z(n13312) );
  XOR2_X1 U15856 ( .A1(n38290), .A2(n37965), .Z(n37964) );
  INV_X2 U15857 ( .I(n19035), .ZN(n37965) );
  INV_X4 U15858 ( .I(n15049), .ZN(n38404) );
  XOR2_X1 U15859 ( .A1(n28830), .A2(n7744), .Z(n29029) );
  NAND2_X2 U15860 ( .A1(n34753), .A2(n31887), .ZN(n28830) );
  OR2_X1 U15864 ( .A1(n21497), .A2(n14418), .Z(n15707) );
  BUF_X2 U15865 ( .I(n33514), .Z(n37966) );
  NAND3_X2 U15866 ( .A1(n25435), .A2(n39269), .A3(n4467), .ZN(n12893) );
  OR2_X2 U15867 ( .A1(n13561), .A2(n14381), .Z(n22816) );
  NAND2_X2 U15868 ( .A1(n34883), .A2(n38102), .ZN(n26532) );
  XOR2_X1 U15869 ( .A1(n24935), .A2(n24999), .Z(n20618) );
  NAND3_X2 U15870 ( .A1(n14782), .A2(n9912), .A3(n15689), .ZN(n24999) );
  XOR2_X1 U15872 ( .A1(n821), .A2(n37968), .Z(n35077) );
  XOR2_X1 U15876 ( .A1(n37969), .A2(n32309), .Z(n39710) );
  XOR2_X1 U15882 ( .A1(n5848), .A2(n29602), .Z(n37969) );
  OR2_X1 U15887 ( .A1(n19590), .A2(n26042), .Z(n25828) );
  NAND3_X2 U15889 ( .A1(n22962), .A2(n23020), .A3(n10507), .ZN(n37970) );
  INV_X1 U15890 ( .I(n28647), .ZN(n30951) );
  OAI21_X2 U15891 ( .A1(n9099), .A2(n37971), .B(n9098), .ZN(n7974) );
  AOI22_X2 U15895 ( .A1(n14807), .A2(n26661), .B1(n39342), .B2(n14458), .ZN(
        n37971) );
  NAND2_X1 U15900 ( .A1(n6876), .A2(n21101), .ZN(n5773) );
  NAND2_X2 U15903 ( .A1(n34001), .A2(n27363), .ZN(n6876) );
  NAND2_X2 U15904 ( .A1(n37972), .A2(n19812), .ZN(n22573) );
  NAND2_X2 U15909 ( .A1(n17896), .A2(n17898), .ZN(n37972) );
  XOR2_X1 U15913 ( .A1(n37973), .A2(n29001), .Z(n32718) );
  NAND2_X1 U15914 ( .A1(n18199), .A2(n13029), .ZN(n23351) );
  NAND2_X2 U15915 ( .A1(n35067), .A2(n22846), .ZN(n18199) );
  XOR2_X1 U15918 ( .A1(n12393), .A2(n37974), .Z(n22639) );
  INV_X2 U15931 ( .I(n8312), .ZN(n37974) );
  OAI22_X2 U15932 ( .A1(n7816), .A2(n916), .B1(n7815), .B2(n7814), .ZN(n8312)
         );
  XOR2_X1 U15939 ( .A1(n25189), .A2(n20707), .Z(n25317) );
  NAND2_X2 U15944 ( .A1(n38083), .A2(n471), .ZN(n25189) );
  AOI21_X2 U15946 ( .A1(n5254), .A2(n1034), .B(n7657), .ZN(n37975) );
  NAND2_X2 U15947 ( .A1(n37977), .A2(n20583), .ZN(n36908) );
  XOR2_X1 U15950 ( .A1(n36515), .A2(n24054), .Z(n798) );
  NAND3_X1 U15955 ( .A1(n7251), .A2(n32682), .A3(n36935), .ZN(n8048) );
  XOR2_X1 U15956 ( .A1(n26597), .A2(n13232), .Z(n11600) );
  XOR2_X1 U15957 ( .A1(n38137), .A2(n10776), .Z(n26597) );
  NAND2_X2 U15960 ( .A1(n35709), .A2(n31060), .ZN(n29803) );
  NAND3_X1 U15962 ( .A1(n23013), .A2(n4573), .A3(n39527), .ZN(n16400) );
  XOR2_X1 U15963 ( .A1(n26574), .A2(n26575), .Z(n36864) );
  AND2_X1 U15966 ( .A1(n21232), .A2(n27028), .Z(n37978) );
  NAND3_X1 U15967 ( .A1(n18408), .A2(n22274), .A3(n22151), .ZN(n22152) );
  XOR2_X1 U15968 ( .A1(n37979), .A2(n12322), .Z(n36868) );
  XOR2_X1 U15971 ( .A1(n39118), .A2(n35639), .Z(n37979) );
  NOR2_X2 U15974 ( .A1(n19228), .A2(n37980), .ZN(n2273) );
  NAND2_X2 U15976 ( .A1(n5249), .A2(n5248), .ZN(n26031) );
  XOR2_X1 U15977 ( .A1(n5241), .A2(n37261), .Z(n484) );
  NOR2_X2 U15978 ( .A1(n37981), .A2(n28639), .ZN(n35788) );
  XOR2_X1 U15983 ( .A1(n9185), .A2(n3963), .Z(n3501) );
  XOR2_X1 U15987 ( .A1(n12310), .A2(n12311), .Z(n25421) );
  NAND3_X2 U15989 ( .A1(n6900), .A2(n6903), .A3(n37982), .ZN(n38981) );
  XOR2_X1 U15990 ( .A1(n27688), .A2(n27502), .Z(n10540) );
  XOR2_X1 U15991 ( .A1(n20706), .A2(n13245), .Z(n27688) );
  NOR2_X2 U15993 ( .A1(n30778), .A2(n13034), .ZN(n39486) );
  OR2_X1 U16002 ( .A1(n31014), .A2(n17095), .Z(n27334) );
  NAND2_X2 U16007 ( .A1(n34309), .A2(n12391), .ZN(n26329) );
  NAND2_X2 U16008 ( .A1(n15867), .A2(n29792), .ZN(n29795) );
  OAI22_X2 U16010 ( .A1(n3693), .A2(n3986), .B1(n20616), .B2(n775), .ZN(n31326) );
  NOR3_X1 U16019 ( .A1(n1531), .A2(n33446), .A3(n39678), .ZN(n9944) );
  XOR2_X1 U16022 ( .A1(n18399), .A2(n1051), .Z(n295) );
  NAND2_X2 U16030 ( .A1(n6785), .A2(n6784), .ZN(n18399) );
  OAI21_X2 U16032 ( .A1(n9656), .A2(n24717), .B(n24719), .ZN(n37985) );
  NAND2_X2 U16034 ( .A1(n37986), .A2(n19951), .ZN(n36538) );
  NAND2_X2 U16038 ( .A1(n30539), .A2(n26702), .ZN(n37986) );
  NOR2_X1 U16039 ( .A1(n26872), .A2(n5935), .ZN(n35345) );
  NAND2_X1 U16046 ( .A1(n37988), .A2(n37987), .ZN(n372) );
  NAND2_X1 U16047 ( .A1(n1385), .A2(n30128), .ZN(n37987) );
  NOR3_X2 U16048 ( .A1(n707), .A2(n7315), .A3(n684), .ZN(n10650) );
  AOI21_X1 U16050 ( .A1(n12617), .A2(n35534), .B(n19481), .ZN(n34373) );
  NAND2_X2 U16051 ( .A1(n39492), .A2(n11156), .ZN(n19481) );
  NAND2_X2 U16053 ( .A1(n31253), .A2(n7397), .ZN(n6191) );
  NAND2_X2 U16054 ( .A1(n37989), .A2(n6934), .ZN(n25086) );
  OAI21_X2 U16055 ( .A1(n34047), .A2(n31743), .B(n37990), .ZN(n3082) );
  XOR2_X1 U16056 ( .A1(n31807), .A2(n38069), .Z(n37991) );
  OR2_X2 U16057 ( .A1(n11481), .A2(n12770), .Z(n9080) );
  OR2_X1 U16060 ( .A1(n20596), .A2(n293), .Z(n19756) );
  NAND2_X1 U16063 ( .A1(n23131), .A2(n22674), .ZN(n22800) );
  NAND2_X2 U16068 ( .A1(n23226), .A2(n23337), .ZN(n23534) );
  NAND3_X2 U16071 ( .A1(n20191), .A2(n22708), .A3(n16400), .ZN(n23226) );
  INV_X2 U16075 ( .I(n19094), .ZN(n38921) );
  NAND2_X2 U16079 ( .A1(n5716), .A2(n37992), .ZN(n31722) );
  NOR2_X2 U16081 ( .A1(n4784), .A2(n4785), .ZN(n37992) );
  BUF_X2 U16091 ( .I(n37051), .Z(n37993) );
  INV_X2 U16092 ( .I(n33750), .ZN(n16566) );
  OAI22_X2 U16099 ( .A1(n33001), .A2(n32948), .B1(n36711), .B2(n38092), .ZN(
        n38187) );
  INV_X2 U16101 ( .I(n25978), .ZN(n37997) );
  CLKBUF_X4 U16105 ( .I(n36509), .Z(n39632) );
  NAND3_X1 U16113 ( .A1(n37153), .A2(n38643), .A3(n26645), .ZN(n38831) );
  XOR2_X1 U16121 ( .A1(n38736), .A2(n25207), .Z(n31724) );
  XOR2_X1 U16123 ( .A1(n25241), .A2(n25181), .Z(n25183) );
  AOI21_X2 U16127 ( .A1(n24657), .A2(n24656), .B(n14781), .ZN(n25241) );
  NAND2_X1 U16129 ( .A1(n10940), .A2(n15873), .ZN(n31184) );
  XOR2_X1 U16131 ( .A1(n24055), .A2(n14312), .Z(n38000) );
  BUF_X2 U16133 ( .I(n26625), .Z(n38002) );
  XOR2_X1 U16137 ( .A1(n7416), .A2(n869), .Z(n34358) );
  NAND2_X1 U16138 ( .A1(n4772), .A2(n36546), .ZN(n6831) );
  NAND2_X2 U16148 ( .A1(n7540), .A2(n12995), .ZN(n36546) );
  XOR2_X1 U16149 ( .A1(n38003), .A2(n1050), .Z(Ciphertext[180]) );
  AOI22_X1 U16153 ( .A1(n30201), .A2(n14387), .B1(n32263), .B2(n36738), .ZN(
        n38003) );
  AND2_X1 U16157 ( .A1(n26933), .A2(n4411), .Z(n5720) );
  XOR2_X1 U16161 ( .A1(n38005), .A2(n29239), .Z(Ciphertext[17]) );
  AOI22_X1 U16163 ( .A1(n35185), .A2(n15482), .B1(n15483), .B2(n29237), .ZN(
        n38005) );
  OR2_X1 U16164 ( .A1(n29241), .A2(n13815), .Z(n9716) );
  OAI22_X2 U16169 ( .A1(n6619), .A2(n5030), .B1(n37640), .B2(n37212), .ZN(
        n8605) );
  INV_X2 U16170 ( .I(n27774), .ZN(n4366) );
  NAND2_X2 U16171 ( .A1(n4120), .A2(n4119), .ZN(n13807) );
  XOR2_X1 U16177 ( .A1(n4560), .A2(n38006), .Z(n19167) );
  XOR2_X1 U16190 ( .A1(n4558), .A2(n4559), .Z(n38006) );
  INV_X2 U16191 ( .I(n17876), .ZN(n20498) );
  OAI22_X2 U16205 ( .A1(n29693), .A2(n29843), .B1(n17877), .B2(n29867), .ZN(
        n17876) );
  OAI21_X2 U16209 ( .A1(n38008), .A2(n38007), .B(n8623), .ZN(n57) );
  NOR2_X2 U16210 ( .A1(n8621), .A2(n8622), .ZN(n38008) );
  INV_X2 U16212 ( .I(n30217), .ZN(n14869) );
  OAI22_X2 U16214 ( .A1(n31025), .A2(n4807), .B1(n2322), .B2(n2321), .ZN(
        n30217) );
  XOR2_X1 U16215 ( .A1(n20715), .A2(n24060), .Z(n20516) );
  NOR2_X1 U16216 ( .A1(n27199), .A2(n4353), .ZN(n27030) );
  INV_X2 U16217 ( .I(n27395), .ZN(n27199) );
  NOR2_X1 U16218 ( .A1(n24279), .A2(n17911), .ZN(n34046) );
  XOR2_X1 U16219 ( .A1(n38009), .A2(n26419), .Z(n34580) );
  NAND2_X1 U16221 ( .A1(n35098), .A2(n33514), .ZN(n36007) );
  OAI21_X2 U16223 ( .A1(n7890), .A2(n25366), .B(n38662), .ZN(n33514) );
  NAND3_X2 U16230 ( .A1(n34654), .A2(n17813), .A3(n22029), .ZN(n9127) );
  NOR2_X2 U16231 ( .A1(n1535), .A2(n32775), .ZN(n25466) );
  BUF_X2 U16239 ( .I(n19587), .Z(n38011) );
  NAND2_X1 U16243 ( .A1(n22931), .A2(n7160), .ZN(n38012) );
  BUF_X2 U16245 ( .I(n25487), .Z(n38013) );
  XOR2_X1 U16246 ( .A1(n23685), .A2(n14289), .Z(n16833) );
  NAND2_X2 U16251 ( .A1(n5181), .A2(n5183), .ZN(n14289) );
  XOR2_X1 U16252 ( .A1(n12690), .A2(n15844), .Z(n9400) );
  XOR2_X1 U16255 ( .A1(n9757), .A2(n27746), .Z(n12690) );
  NOR2_X2 U16257 ( .A1(n21521), .A2(n21587), .ZN(n8600) );
  NAND2_X2 U16258 ( .A1(n1081), .A2(n37508), .ZN(n9082) );
  AOI21_X2 U16262 ( .A1(n27686), .A2(n28193), .B(n37164), .ZN(n38014) );
  INV_X2 U16264 ( .I(n38015), .ZN(n34987) );
  XOR2_X1 U16265 ( .A1(n31485), .A2(n12084), .Z(n38015) );
  NAND2_X1 U16278 ( .A1(n11067), .A2(n37095), .ZN(n29372) );
  OAI22_X2 U16282 ( .A1(n29345), .A2(n39647), .B1(n12479), .B2(n19896), .ZN(
        n35465) );
  INV_X2 U16283 ( .I(n19846), .ZN(n35936) );
  NAND2_X2 U16284 ( .A1(n5768), .A2(n7770), .ZN(n24898) );
  NOR3_X2 U16287 ( .A1(n34071), .A2(n35297), .A3(n32797), .ZN(n27140) );
  XOR2_X1 U16290 ( .A1(n25), .A2(n25148), .Z(n33527) );
  XOR2_X1 U16291 ( .A1(n18366), .A2(n38016), .Z(n26995) );
  XOR2_X1 U16300 ( .A1(n26434), .A2(n31414), .Z(n38016) );
  OR2_X1 U16308 ( .A1(n35300), .A2(n32010), .Z(n24370) );
  OAI21_X2 U16309 ( .A1(n11133), .A2(n24119), .B(n11131), .ZN(n7529) );
  NOR2_X2 U16310 ( .A1(n35360), .A2(n38017), .ZN(n32608) );
  XOR2_X1 U16314 ( .A1(n20424), .A2(n38018), .Z(n33895) );
  XOR2_X1 U16317 ( .A1(n20730), .A2(n26222), .Z(n38018) );
  NAND2_X2 U16322 ( .A1(n18788), .A2(n19499), .ZN(n39232) );
  XNOR2_X1 U16324 ( .A1(n38208), .A2(n16618), .ZN(n39239) );
  XOR2_X1 U16329 ( .A1(n20586), .A2(n24052), .Z(n19188) );
  NAND2_X2 U16336 ( .A1(n39581), .A2(n39333), .ZN(n24052) );
  OAI21_X2 U16338 ( .A1(n13445), .A2(n37904), .B(n12307), .ZN(n9847) );
  XOR2_X1 U16339 ( .A1(n32895), .A2(n4900), .Z(n7140) );
  NOR2_X1 U16340 ( .A1(n21047), .A2(n23020), .ZN(n38019) );
  XOR2_X1 U16341 ( .A1(n33322), .A2(n29463), .Z(n5094) );
  OAI22_X2 U16348 ( .A1(n23593), .A2(n4148), .B1(n4149), .B2(n23594), .ZN(
        n33322) );
  OAI21_X2 U16350 ( .A1(n17863), .A2(n17862), .B(n10894), .ZN(n25113) );
  INV_X2 U16355 ( .I(n5063), .ZN(n38668) );
  NAND2_X1 U16356 ( .A1(n26918), .A2(n13392), .ZN(n33062) );
  NAND2_X2 U16357 ( .A1(n10461), .A2(n35427), .ZN(n27009) );
  XOR2_X1 U16358 ( .A1(n13439), .A2(n9246), .Z(n23802) );
  NAND2_X2 U16360 ( .A1(n33698), .A2(n23584), .ZN(n13439) );
  OAI21_X2 U16365 ( .A1(n23578), .A2(n6945), .B(n1138), .ZN(n21296) );
  NAND2_X2 U16366 ( .A1(n38576), .A2(n38020), .ZN(n36634) );
  OAI21_X2 U16369 ( .A1(n33101), .A2(n36556), .B(n34044), .ZN(n38020) );
  NAND2_X2 U16370 ( .A1(n1759), .A2(n33516), .ZN(n28066) );
  NOR2_X2 U16376 ( .A1(n37105), .A2(n36634), .ZN(n38916) );
  NAND2_X2 U16382 ( .A1(n16579), .A2(n12160), .ZN(n13516) );
  OAI21_X2 U16392 ( .A1(n28623), .A2(n33283), .B(n19161), .ZN(n33519) );
  NAND2_X2 U16393 ( .A1(n33283), .A2(n2147), .ZN(n19161) );
  AND2_X1 U16394 ( .A1(n35427), .A2(n9369), .Z(n27430) );
  BUF_X2 U16395 ( .I(n15037), .Z(n36549) );
  NOR3_X2 U16398 ( .A1(n33513), .A2(n39605), .A3(n24282), .ZN(n32542) );
  NAND2_X2 U16399 ( .A1(n29862), .A2(n9649), .ZN(n29908) );
  XOR2_X1 U16400 ( .A1(n24938), .A2(n25030), .Z(n38992) );
  NOR2_X2 U16401 ( .A1(n24607), .A2(n12846), .ZN(n25030) );
  NAND3_X2 U16403 ( .A1(n23511), .A2(n23510), .A3(n11245), .ZN(n15299) );
  NAND2_X2 U16405 ( .A1(n12156), .A2(n35427), .ZN(n11256) );
  OR2_X1 U16407 ( .A1(n30156), .A2(n14254), .Z(n31357) );
  XOR2_X1 U16408 ( .A1(n29100), .A2(n38384), .Z(n30156) );
  OR2_X1 U16412 ( .A1(n5282), .A2(n24515), .Z(n34143) );
  NAND2_X1 U16415 ( .A1(n38023), .A2(n1536), .ZN(n5292) );
  OAI22_X1 U16417 ( .A1(n1531), .A2(n25692), .B1(n8014), .B2(n12500), .ZN(
        n38023) );
  AOI22_X2 U16421 ( .A1(n8946), .A2(n33867), .B1(n27652), .B2(n13955), .ZN(
        n8944) );
  AOI21_X1 U16423 ( .A1(n28235), .A2(n28234), .B(n11283), .ZN(n38512) );
  XOR2_X1 U16424 ( .A1(n19862), .A2(n19902), .Z(n6923) );
  XOR2_X1 U16425 ( .A1(n27594), .A2(n27796), .Z(n27753) );
  NAND3_X2 U16427 ( .A1(n17151), .A2(n15275), .A3(n15277), .ZN(n27796) );
  XOR2_X1 U16435 ( .A1(n38026), .A2(n2176), .Z(n8526) );
  NAND2_X2 U16436 ( .A1(n36849), .A2(n32081), .ZN(n22488) );
  XOR2_X1 U16438 ( .A1(n9036), .A2(n29282), .Z(n13700) );
  NAND2_X2 U16439 ( .A1(n137), .A2(n6039), .ZN(n9036) );
  NOR2_X1 U16440 ( .A1(n36854), .A2(n28234), .ZN(n4415) );
  NOR2_X1 U16442 ( .A1(n2573), .A2(n4531), .ZN(n12379) );
  NAND2_X2 U16444 ( .A1(n4244), .A2(n38027), .ZN(n15716) );
  NAND2_X1 U16445 ( .A1(n33061), .A2(n18116), .ZN(n38027) );
  NAND2_X1 U16448 ( .A1(n39017), .A2(n15358), .ZN(n35709) );
  NAND2_X2 U16452 ( .A1(n14216), .A2(n7643), .ZN(n31486) );
  XOR2_X1 U16453 ( .A1(n31541), .A2(n4301), .Z(n22233) );
  XOR2_X1 U16456 ( .A1(n38028), .A2(n26204), .Z(n33067) );
  XNOR2_X1 U16463 ( .A1(n16610), .A2(n9576), .ZN(n26204) );
  NOR2_X2 U16465 ( .A1(n149), .A2(n4467), .ZN(n38029) );
  OAI21_X2 U16475 ( .A1(n31177), .A2(n31175), .B(n38030), .ZN(n39268) );
  AOI22_X2 U16482 ( .A1(n14645), .A2(n8735), .B1(n16590), .B2(n15872), .ZN(
        n38030) );
  XOR2_X1 U16483 ( .A1(n13569), .A2(n27470), .Z(n13568) );
  OR2_X1 U16484 ( .A1(n10375), .A2(n33431), .Z(n22834) );
  XOR2_X1 U16486 ( .A1(n22651), .A2(n12267), .Z(n22463) );
  OAI21_X2 U16488 ( .A1(n16624), .A2(n16623), .B(n22081), .ZN(n22651) );
  OAI22_X2 U16497 ( .A1(n1234), .A2(n14394), .B1(n26719), .B2(n735), .ZN(
        n11248) );
  XOR2_X1 U16499 ( .A1(n38427), .A2(n33576), .Z(n10686) );
  NAND2_X2 U16504 ( .A1(n16325), .A2(n14461), .ZN(n5509) );
  XOR2_X1 U16510 ( .A1(n28827), .A2(n29052), .Z(n8909) );
  NAND2_X2 U16512 ( .A1(n8910), .A2(n8911), .ZN(n28827) );
  XOR2_X1 U16513 ( .A1(n38031), .A2(n1700), .Z(Ciphertext[6]) );
  NOR2_X1 U16515 ( .A1(n9606), .A2(n9607), .ZN(n38031) );
  XOR2_X1 U16516 ( .A1(n10406), .A2(n10407), .Z(n11657) );
  OAI21_X2 U16517 ( .A1(n24355), .A2(n8359), .B(n19818), .ZN(n35666) );
  NOR2_X2 U16519 ( .A1(n39074), .A2(n32069), .ZN(n24355) );
  INV_X2 U16521 ( .I(n13761), .ZN(n29219) );
  NAND3_X2 U16522 ( .A1(n35502), .A2(n30655), .A3(n32267), .ZN(n13761) );
  NAND3_X2 U16524 ( .A1(n25360), .A2(n19971), .A3(n19311), .ZN(n39108) );
  NAND2_X1 U16525 ( .A1(n13663), .A2(n17248), .ZN(n39402) );
  INV_X4 U16526 ( .I(n24709), .ZN(n6491) );
  NAND2_X2 U16527 ( .A1(n12422), .A2(n12424), .ZN(n24709) );
  XOR2_X1 U16537 ( .A1(n21079), .A2(n38033), .Z(n19948) );
  XOR2_X1 U16541 ( .A1(n31692), .A2(n28853), .Z(n38033) );
  NOR2_X2 U16546 ( .A1(n27341), .A2(n32205), .ZN(n27133) );
  INV_X2 U16561 ( .I(n26888), .ZN(n27341) );
  NAND3_X2 U16564 ( .A1(n26698), .A2(n142), .A3(n26699), .ZN(n26888) );
  NAND3_X2 U16565 ( .A1(n36556), .A2(n19070), .A3(n17810), .ZN(n38034) );
  XOR2_X1 U16566 ( .A1(n38035), .A2(n19128), .Z(Ciphertext[20]) );
  NAND3_X1 U16567 ( .A1(n17955), .A2(n6841), .A3(n6842), .ZN(n38035) );
  XOR2_X1 U16568 ( .A1(n11794), .A2(n23869), .Z(n15114) );
  NOR2_X2 U16571 ( .A1(n38036), .A2(n24154), .ZN(n24698) );
  XOR2_X1 U16572 ( .A1(n13703), .A2(n13877), .Z(n39613) );
  OAI22_X2 U16574 ( .A1(n4089), .A2(n4253), .B1(n38572), .B2(n4254), .ZN(
        n13877) );
  XOR2_X1 U16576 ( .A1(n20294), .A2(n18153), .Z(n31752) );
  NOR2_X2 U16577 ( .A1(n23616), .A2(n38037), .ZN(n24038) );
  AOI21_X2 U16581 ( .A1(n36635), .A2(n39434), .B(n23614), .ZN(n38037) );
  XOR2_X1 U16587 ( .A1(n38038), .A2(n18993), .Z(Ciphertext[15]) );
  NOR2_X1 U16590 ( .A1(n14200), .A2(n14197), .ZN(n38038) );
  NAND2_X1 U16593 ( .A1(n26761), .A2(n26810), .ZN(n11515) );
  INV_X1 U16595 ( .I(n24974), .ZN(n35339) );
  XOR2_X1 U16596 ( .A1(n36748), .A2(n23609), .Z(n23677) );
  XOR2_X1 U16599 ( .A1(n30610), .A2(n30609), .Z(n5274) );
  XOR2_X1 U16602 ( .A1(n26321), .A2(n39667), .Z(n26630) );
  NAND2_X2 U16604 ( .A1(n38040), .A2(n38039), .ZN(n18303) );
  OAI21_X2 U16607 ( .A1(n13421), .A2(n21892), .B(n21893), .ZN(n38039) );
  OAI21_X2 U16613 ( .A1(n21896), .A2(n15528), .B(n21895), .ZN(n38040) );
  XOR2_X1 U16614 ( .A1(n10562), .A2(n27859), .Z(n10483) );
  XOR2_X1 U16615 ( .A1(n27779), .A2(n27778), .Z(n27859) );
  BUF_X2 U16618 ( .I(n38619), .Z(n38041) );
  INV_X4 U16620 ( .I(n26935), .ZN(n1093) );
  INV_X2 U16625 ( .I(n29070), .ZN(n7489) );
  XOR2_X1 U16643 ( .A1(n8634), .A2(n23950), .Z(n636) );
  XOR2_X1 U16645 ( .A1(n33322), .A2(n23680), .Z(n23950) );
  XOR2_X1 U16646 ( .A1(n25179), .A2(n25096), .Z(n31563) );
  NAND2_X2 U16647 ( .A1(n12832), .A2(n24085), .ZN(n25096) );
  NAND2_X2 U16648 ( .A1(n7892), .A2(n33437), .ZN(n9200) );
  NAND2_X2 U16649 ( .A1(n2684), .A2(n2685), .ZN(n23889) );
  NOR2_X2 U16651 ( .A1(n24802), .A2(n35901), .ZN(n15414) );
  XOR2_X1 U16656 ( .A1(n6130), .A2(n26026), .Z(n26399) );
  NOR2_X2 U16664 ( .A1(n33950), .A2(n25692), .ZN(n8222) );
  XOR2_X1 U16667 ( .A1(n32349), .A2(n38043), .Z(n9986) );
  INV_X2 U16668 ( .I(n25200), .ZN(n38043) );
  XOR2_X1 U16669 ( .A1(n25296), .A2(n24991), .Z(n25200) );
  NAND2_X2 U16676 ( .A1(n11614), .A2(n1433), .ZN(n13780) );
  XOR2_X1 U16681 ( .A1(n39378), .A2(n30849), .Z(n38048) );
  NAND2_X2 U16682 ( .A1(n17335), .A2(n2458), .ZN(n17333) );
  OR3_X2 U16687 ( .A1(n15515), .A2(n25480), .A3(n16933), .Z(n25529) );
  OAI22_X2 U16690 ( .A1(n17225), .A2(n1061), .B1(n1062), .B2(n20566), .ZN(
        n39240) );
  NAND3_X2 U16691 ( .A1(n29370), .A2(n39677), .A3(n4669), .ZN(n39208) );
  OAI21_X2 U16692 ( .A1(n11054), .A2(n37106), .B(n38044), .ZN(n8542) );
  XOR2_X1 U16694 ( .A1(n38045), .A2(n38711), .Z(n25544) );
  XOR2_X1 U16697 ( .A1(n5433), .A2(n38458), .Z(n38045) );
  XOR2_X1 U16699 ( .A1(n5803), .A2(n5804), .Z(n39353) );
  XOR2_X1 U16702 ( .A1(n38046), .A2(n19738), .Z(Ciphertext[92]) );
  NAND4_X2 U16703 ( .A1(n29714), .A2(n29716), .A3(n29713), .A4(n29715), .ZN(
        n38046) );
  NAND2_X2 U16706 ( .A1(n31960), .A2(n19911), .ZN(n15868) );
  XOR2_X1 U16710 ( .A1(n38048), .A2(n23410), .Z(n34473) );
  XOR2_X1 U16713 ( .A1(n8852), .A2(n18430), .Z(n29024) );
  NAND2_X2 U16716 ( .A1(n8854), .A2(n8853), .ZN(n18430) );
  XOR2_X1 U16718 ( .A1(n12840), .A2(n798), .Z(n19295) );
  NAND3_X2 U16719 ( .A1(n20177), .A2(n22819), .A3(n20176), .ZN(n38724) );
  AOI22_X2 U16725 ( .A1(n3309), .A2(n5591), .B1(n23412), .B2(n1636), .ZN(
        n38049) );
  OAI21_X2 U16726 ( .A1(n38782), .A2(n19941), .B(n16677), .ZN(n38050) );
  XOR2_X1 U16732 ( .A1(n26590), .A2(n19450), .Z(n13496) );
  INV_X2 U16735 ( .I(n26272), .ZN(n26687) );
  XOR2_X1 U16737 ( .A1(n29057), .A2(n18133), .Z(n19428) );
  NAND2_X2 U16738 ( .A1(n28338), .A2(n9442), .ZN(n18133) );
  XOR2_X1 U16739 ( .A1(n35065), .A2(n23982), .Z(n14386) );
  OAI22_X2 U16743 ( .A1(n10495), .A2(n10494), .B1(n5049), .B2(n1134), .ZN(
        n35065) );
  XOR2_X1 U16747 ( .A1(n26389), .A2(n26436), .Z(n26508) );
  NAND2_X2 U16749 ( .A1(n25926), .A2(n9226), .ZN(n26389) );
  XOR2_X1 U16750 ( .A1(n1661), .A2(n3953), .Z(n13842) );
  XOR2_X1 U16751 ( .A1(n22534), .A2(n22520), .Z(n22524) );
  XOR2_X1 U16753 ( .A1(n22628), .A2(n1662), .Z(n22534) );
  INV_X2 U16755 ( .I(n38052), .ZN(n15466) );
  XOR2_X1 U16760 ( .A1(Plaintext[168]), .A2(Key[168]), .Z(n38052) );
  NAND2_X2 U16762 ( .A1(n11337), .A2(n26935), .ZN(n11336) );
  NAND3_X2 U16764 ( .A1(n28491), .A2(n28490), .A3(n28489), .ZN(n28492) );
  BUF_X2 U16766 ( .I(n29344), .Z(n29458) );
  INV_X2 U16767 ( .I(n38053), .ZN(n17307) );
  NOR2_X2 U16770 ( .A1(n21460), .A2(n21459), .ZN(n38053) );
  OAI21_X2 U16776 ( .A1(n21539), .A2(n21542), .B(n9424), .ZN(n21459) );
  NOR2_X2 U16782 ( .A1(n12191), .A2(n5487), .ZN(n5490) );
  INV_X2 U16783 ( .I(n18681), .ZN(n12191) );
  NAND2_X2 U16784 ( .A1(n35006), .A2(n17201), .ZN(n18681) );
  XOR2_X1 U16787 ( .A1(n2627), .A2(n269), .Z(n3207) );
  NAND2_X2 U16790 ( .A1(n1834), .A2(n32184), .ZN(n2627) );
  NAND2_X2 U16791 ( .A1(n11225), .A2(n36483), .ZN(n27435) );
  INV_X1 U16794 ( .I(n19279), .ZN(n38626) );
  XOR2_X1 U16795 ( .A1(n12145), .A2(n39579), .Z(n36239) );
  NAND2_X2 U16796 ( .A1(n11279), .A2(n11280), .ZN(n35203) );
  AOI22_X2 U16801 ( .A1(n37225), .A2(n38055), .B1(n2012), .B2(n17960), .ZN(
        n2009) );
  INV_X2 U16804 ( .I(n1036), .ZN(n38055) );
  NAND2_X2 U16805 ( .A1(n38949), .A2(n39748), .ZN(n34350) );
  NOR2_X1 U16808 ( .A1(n15048), .A2(n11737), .ZN(n38765) );
  NAND2_X2 U16818 ( .A1(n38056), .A2(n27543), .ZN(n16853) );
  NAND2_X2 U16828 ( .A1(n38057), .A2(n13093), .ZN(n13414) );
  OAI21_X2 U16832 ( .A1(n32873), .A2(n32872), .B(n37883), .ZN(n38057) );
  NAND2_X2 U16833 ( .A1(n14833), .A2(n4424), .ZN(n2480) );
  XOR2_X1 U16838 ( .A1(n38352), .A2(n39698), .Z(n38058) );
  INV_X2 U16846 ( .I(n5282), .ZN(n24603) );
  XOR2_X1 U16849 ( .A1(n5625), .A2(n17884), .Z(n27496) );
  NOR2_X1 U16854 ( .A1(n22265), .A2(n22267), .ZN(n11684) );
  OAI21_X1 U16856 ( .A1(n36910), .A2(n9914), .B(n29224), .ZN(n13771) );
  INV_X1 U16857 ( .I(n29220), .ZN(n36910) );
  AND2_X1 U16863 ( .A1(n31357), .A2(n35870), .Z(n38236) );
  OAI21_X2 U16865 ( .A1(n38059), .A2(n34817), .B(n28212), .ZN(n39087) );
  NOR2_X2 U16869 ( .A1(n28213), .A2(n16950), .ZN(n38059) );
  INV_X2 U16880 ( .I(n8475), .ZN(n38799) );
  XOR2_X1 U16881 ( .A1(n27516), .A2(n19800), .Z(n31070) );
  NAND2_X2 U16883 ( .A1(n14058), .A2(n14057), .ZN(n27516) );
  OAI21_X2 U16884 ( .A1(n32343), .A2(n32344), .B(n11679), .ZN(n20190) );
  NOR2_X2 U16886 ( .A1(n6615), .A2(n38284), .ZN(n32343) );
  NAND3_X2 U16888 ( .A1(n6195), .A2(n32545), .A3(n6192), .ZN(n36386) );
  AOI21_X2 U16890 ( .A1(n29873), .A2(n29869), .B(n33297), .ZN(n38217) );
  NAND3_X2 U16893 ( .A1(n38757), .A2(n31170), .A3(n35547), .ZN(n30095) );
  INV_X2 U16896 ( .I(n13333), .ZN(n32555) );
  NOR3_X2 U16897 ( .A1(n30694), .A2(n25622), .A3(n33785), .ZN(n3010) );
  OR2_X1 U16903 ( .A1(n6932), .A2(n16619), .Z(n4949) );
  XOR2_X1 U16904 ( .A1(n6727), .A2(n25263), .Z(n25153) );
  NOR2_X1 U16909 ( .A1(n29627), .A2(n29617), .ZN(n38063) );
  XOR2_X1 U16911 ( .A1(n26437), .A2(n26009), .Z(n26528) );
  OR2_X2 U16914 ( .A1(n27875), .A2(n17378), .Z(n28199) );
  XOR2_X1 U16915 ( .A1(n16054), .A2(n6758), .Z(n29060) );
  AOI21_X2 U16919 ( .A1(n6789), .A2(n6788), .B(n38064), .ZN(n6786) );
  NOR3_X1 U16920 ( .A1(n5239), .A2(n5352), .A3(n34008), .ZN(n38064) );
  INV_X2 U16922 ( .I(n27588), .ZN(n27587) );
  NAND2_X2 U16923 ( .A1(n35332), .A2(n2722), .ZN(n27588) );
  NAND2_X2 U16930 ( .A1(n10231), .A2(n11616), .ZN(n26899) );
  INV_X2 U16938 ( .I(n38066), .ZN(n16174) );
  XNOR2_X1 U16941 ( .A1(n32431), .A2(n32432), .ZN(n38066) );
  NAND3_X1 U16947 ( .A1(n14375), .A2(n38168), .A3(n35855), .ZN(n18352) );
  XOR2_X1 U16950 ( .A1(n10233), .A2(n5584), .Z(n20960) );
  NAND3_X2 U16951 ( .A1(n9142), .A2(n29180), .A3(n7933), .ZN(n30117) );
  OR2_X1 U16952 ( .A1(n23468), .A2(n23467), .Z(n7534) );
  AND2_X1 U16954 ( .A1(n19782), .A2(n24465), .Z(n35873) );
  NAND2_X2 U16956 ( .A1(n38437), .A2(n26042), .ZN(n17178) );
  AND2_X1 U16957 ( .A1(n36810), .A2(n32471), .Z(n16299) );
  INV_X2 U16965 ( .I(n24827), .ZN(n11271) );
  NAND3_X2 U16968 ( .A1(n1877), .A2(n1875), .A3(n5432), .ZN(n24827) );
  XOR2_X1 U16979 ( .A1(n27480), .A2(n20167), .Z(n20166) );
  XOR2_X1 U16982 ( .A1(n27851), .A2(n5750), .Z(n27480) );
  XOR2_X1 U16985 ( .A1(n38067), .A2(n29295), .Z(Ciphertext[3]) );
  XOR2_X1 U16987 ( .A1(n28783), .A2(n12989), .Z(n29128) );
  NAND2_X2 U16990 ( .A1(n5397), .A2(n5398), .ZN(n28783) );
  NAND2_X2 U17001 ( .A1(n910), .A2(n2678), .ZN(n25977) );
  NOR2_X2 U17004 ( .A1(n19544), .A2(n7790), .ZN(n9025) );
  XOR2_X1 U17007 ( .A1(n14353), .A2(n17925), .Z(n14454) );
  INV_X1 U17012 ( .I(n38070), .ZN(n35360) );
  OAI21_X1 U17013 ( .A1(n34567), .A2(n34568), .B(n28735), .ZN(n38070) );
  INV_X2 U17015 ( .I(n12572), .ZN(n30211) );
  NAND3_X2 U17016 ( .A1(n39432), .A2(n7893), .A3(n39431), .ZN(n12572) );
  INV_X4 U17017 ( .I(n17685), .ZN(n937) );
  AOI22_X2 U17022 ( .A1(n17794), .A2(n29263), .B1(n37185), .B2(n16123), .ZN(
        n38071) );
  NAND2_X1 U17024 ( .A1(n38072), .A2(n10703), .ZN(n39551) );
  NOR2_X1 U17025 ( .A1(n39393), .A2(n39392), .ZN(n38072) );
  XOR2_X1 U17026 ( .A1(n23874), .A2(n19608), .Z(n23876) );
  INV_X2 U17029 ( .I(n24887), .ZN(n38073) );
  AND2_X1 U17033 ( .A1(n7044), .A2(n38073), .Z(n17863) );
  XOR2_X1 U17044 ( .A1(n22789), .A2(n22728), .Z(n22581) );
  NOR2_X2 U17048 ( .A1(n39190), .A2(n34433), .ZN(n34753) );
  AND2_X1 U17049 ( .A1(n19560), .A2(n24872), .Z(n30422) );
  NAND2_X2 U17050 ( .A1(n31161), .A2(n18148), .ZN(n19560) );
  NAND2_X2 U17053 ( .A1(n4246), .A2(n4247), .ZN(n38619) );
  XOR2_X1 U17058 ( .A1(n36617), .A2(n38076), .Z(n35544) );
  XNOR2_X1 U17070 ( .A1(n27845), .A2(n8875), .ZN(n2437) );
  NOR2_X2 U17074 ( .A1(n38247), .A2(n25820), .ZN(n31473) );
  NAND2_X2 U17075 ( .A1(n18686), .A2(n18685), .ZN(n5819) );
  AOI22_X2 U17078 ( .A1(n21943), .A2(n20923), .B1(n16128), .B2(n16052), .ZN(
        n18685) );
  INV_X4 U17081 ( .I(n3293), .ZN(n21583) );
  NAND2_X1 U17085 ( .A1(n31461), .A2(n8349), .ZN(n38077) );
  XOR2_X1 U17086 ( .A1(n8654), .A2(n37252), .Z(n9590) );
  XNOR2_X1 U17087 ( .A1(n39391), .A2(n8532), .ZN(n8654) );
  NOR2_X2 U17088 ( .A1(n35377), .A2(n34962), .ZN(n31945) );
  BUF_X2 U17089 ( .I(n27314), .Z(n38079) );
  XOR2_X1 U17090 ( .A1(n10636), .A2(n38080), .Z(n10733) );
  XOR2_X1 U17098 ( .A1(n12026), .A2(n12480), .Z(n38080) );
  INV_X2 U17104 ( .I(n38081), .ZN(n6640) );
  OAI21_X1 U17115 ( .A1(n12675), .A2(n10563), .B(n38959), .ZN(n9439) );
  NAND3_X2 U17117 ( .A1(n3583), .A2(n20472), .A3(n32927), .ZN(n39161) );
  OAI21_X2 U17122 ( .A1(n33437), .A2(n39083), .B(n30204), .ZN(n30206) );
  XOR2_X1 U17132 ( .A1(n15904), .A2(n38082), .Z(n32821) );
  XOR2_X1 U17135 ( .A1(n23809), .A2(n37224), .Z(n38082) );
  XOR2_X1 U17138 ( .A1(n11870), .A2(n11871), .Z(n13499) );
  BUF_X4 U17146 ( .I(n17095), .Z(n33335) );
  OAI21_X2 U17148 ( .A1(n10902), .A2(n31157), .B(n37524), .ZN(n26151) );
  XOR2_X1 U17152 ( .A1(n27787), .A2(n27632), .Z(n27527) );
  NAND2_X2 U17156 ( .A1(n27023), .A2(n27024), .ZN(n27787) );
  AOI21_X1 U17167 ( .A1(n39584), .A2(n9743), .B(n949), .ZN(n5162) );
  XOR2_X1 U17172 ( .A1(n24001), .A2(n33232), .Z(n33231) );
  OAI21_X2 U17175 ( .A1(n5591), .A2(n38085), .B(n23606), .ZN(n9331) );
  OR2_X1 U17180 ( .A1(n23308), .A2(n18850), .Z(n38085) );
  XOR2_X1 U17182 ( .A1(n10767), .A2(n12003), .Z(n3392) );
  XOR2_X1 U17186 ( .A1(n16096), .A2(n7464), .Z(n10767) );
  XOR2_X1 U17187 ( .A1(n29068), .A2(n38086), .Z(n21323) );
  XOR2_X1 U17191 ( .A1(n34178), .A2(n38087), .Z(n38086) );
  AND2_X1 U17195 ( .A1(n11150), .A2(n36708), .Z(n832) );
  NAND2_X2 U17196 ( .A1(n39290), .A2(n38088), .ZN(n3510) );
  NAND3_X1 U17198 ( .A1(n224), .A2(n34374), .A3(n9193), .ZN(n38088) );
  AND2_X1 U17213 ( .A1(n2597), .A2(n39699), .Z(n2595) );
  XOR2_X1 U17214 ( .A1(n10488), .A2(n22643), .Z(n10705) );
  AOI21_X2 U17215 ( .A1(n16027), .A2(n7771), .B(n347), .ZN(n22643) );
  AND2_X1 U17219 ( .A1(n28676), .A2(n28578), .Z(n9951) );
  OR2_X1 U17220 ( .A1(n9801), .A2(n11784), .Z(n13004) );
  XOR2_X1 U17222 ( .A1(n35105), .A2(n2196), .Z(n9801) );
  INV_X2 U17223 ( .I(n38089), .ZN(n18920) );
  XOR2_X1 U17227 ( .A1(n18922), .A2(n18921), .Z(n38089) );
  NAND2_X1 U17229 ( .A1(n38090), .A2(n19521), .ZN(n13913) );
  OAI21_X1 U17231 ( .A1(n34401), .A2(n14483), .B(n22901), .ZN(n38090) );
  INV_X2 U17234 ( .I(n14502), .ZN(n23201) );
  XOR2_X1 U17235 ( .A1(n10502), .A2(n10501), .Z(n14502) );
  XOR2_X1 U17240 ( .A1(n24033), .A2(n2220), .Z(n33578) );
  AOI22_X2 U17241 ( .A1(n3821), .A2(n33885), .B1(n21892), .B2(n21489), .ZN(
        n38091) );
  NOR2_X2 U17249 ( .A1(n32683), .A2(n11796), .ZN(n35434) );
  BUF_X4 U17251 ( .I(n5745), .Z(n5675) );
  NAND2_X2 U17253 ( .A1(n34632), .A2(n14506), .ZN(n15581) );
  NOR2_X2 U17255 ( .A1(n27484), .A2(n39296), .ZN(n11041) );
  NAND2_X2 U17256 ( .A1(n35576), .A2(n14502), .ZN(n3683) );
  INV_X2 U17257 ( .I(n14833), .ZN(n22128) );
  NAND2_X1 U17258 ( .A1(n30060), .A2(n30793), .ZN(n30062) );
  XOR2_X1 U17259 ( .A1(n4828), .A2(n31965), .Z(n26503) );
  OAI21_X2 U17264 ( .A1(n3519), .A2(n3518), .B(n3516), .ZN(n31965) );
  BUF_X2 U17266 ( .I(n3449), .Z(n38092) );
  NAND3_X2 U17267 ( .A1(n27200), .A2(n17298), .A3(n32961), .ZN(n38093) );
  NOR2_X2 U17270 ( .A1(n22927), .A2(n8141), .ZN(n20788) );
  AND2_X2 U17272 ( .A1(n8142), .A2(n22917), .Z(n8141) );
  NAND2_X2 U17273 ( .A1(n36527), .A2(n8507), .ZN(n38704) );
  INV_X2 U17274 ( .I(n21167), .ZN(n8445) );
  XOR2_X1 U17275 ( .A1(n38094), .A2(n22590), .Z(n22678) );
  XOR2_X1 U17276 ( .A1(n22529), .A2(n22528), .Z(n38094) );
  XOR2_X1 U17286 ( .A1(n7936), .A2(n38095), .Z(n3705) );
  XOR2_X1 U17290 ( .A1(n3703), .A2(n31547), .Z(n38095) );
  XOR2_X1 U17296 ( .A1(n21036), .A2(n38096), .Z(n11250) );
  XOR2_X1 U17297 ( .A1(n34531), .A2(n31320), .Z(n38096) );
  XOR2_X1 U17299 ( .A1(n3610), .A2(n15346), .Z(n9205) );
  NAND3_X2 U17305 ( .A1(n2588), .A2(n2589), .A3(n2590), .ZN(n3610) );
  NAND2_X1 U17306 ( .A1(n2765), .A2(n10463), .ZN(n4865) );
  NAND2_X2 U17308 ( .A1(n6099), .A2(n6098), .ZN(n2765) );
  XOR2_X1 U17310 ( .A1(n12741), .A2(n8940), .Z(n19374) );
  NAND2_X2 U17312 ( .A1(n11536), .A2(n11534), .ZN(n8940) );
  NAND2_X2 U17313 ( .A1(n17792), .A2(n21587), .ZN(n21520) );
  NAND2_X2 U17315 ( .A1(n38098), .A2(n6734), .ZN(n29555) );
  NAND2_X1 U17317 ( .A1(n20426), .A2(n32987), .ZN(n38098) );
  NAND2_X2 U17318 ( .A1(n3050), .A2(n27972), .ZN(n28948) );
  AND2_X1 U17326 ( .A1(n7901), .A2(n33644), .Z(n18354) );
  XOR2_X1 U17328 ( .A1(n22563), .A2(n16667), .Z(n7038) );
  NOR2_X2 U17331 ( .A1(n8947), .A2(n9485), .ZN(n8744) );
  INV_X2 U17332 ( .I(n38099), .ZN(n8947) );
  NAND2_X2 U17333 ( .A1(n8948), .A2(n22222), .ZN(n38099) );
  NAND3_X1 U17335 ( .A1(n7373), .A2(n18120), .A3(n30680), .ZN(n38101) );
  INV_X4 U17342 ( .I(n27064), .ZN(n1221) );
  NAND3_X1 U17345 ( .A1(n17365), .A2(n15308), .A3(n15209), .ZN(n15307) );
  NAND2_X2 U17349 ( .A1(n10883), .A2(n28685), .ZN(n11030) );
  NOR3_X2 U17352 ( .A1(n20578), .A2(n26841), .A3(n36392), .ZN(n36647) );
  AND2_X1 U17357 ( .A1(n39054), .A2(n17022), .Z(n38234) );
  XOR2_X1 U17360 ( .A1(n38103), .A2(n4397), .Z(n18853) );
  XOR2_X1 U17361 ( .A1(n5655), .A2(n6795), .Z(n38103) );
  XOR2_X1 U17365 ( .A1(n34513), .A2(n26262), .Z(n13171) );
  XOR2_X1 U17368 ( .A1(n13802), .A2(n8059), .Z(n27832) );
  NAND3_X2 U17369 ( .A1(n27040), .A2(n27039), .A3(n27041), .ZN(n13802) );
  AOI21_X2 U17372 ( .A1(n18901), .A2(n26825), .B(n38104), .ZN(n35036) );
  NOR2_X2 U17373 ( .A1(n26823), .A2(n26824), .ZN(n38104) );
  INV_X2 U17387 ( .I(n38106), .ZN(n10261) );
  NOR2_X1 U17388 ( .A1(n38106), .A2(n38105), .ZN(n6724) );
  NAND2_X2 U17389 ( .A1(n18686), .A2(n18685), .ZN(n38106) );
  XOR2_X1 U17396 ( .A1(n38107), .A2(n39259), .Z(n38554) );
  XOR2_X1 U17398 ( .A1(n27643), .A2(n37147), .Z(n38107) );
  NAND2_X1 U17399 ( .A1(n10210), .A2(n35869), .ZN(n3430) );
  INV_X2 U17406 ( .I(n38108), .ZN(n8604) );
  XNOR2_X1 U17408 ( .A1(n18663), .A2(n33831), .ZN(n38108) );
  OAI21_X2 U17409 ( .A1(n38338), .A2(n1110), .B(n25754), .ZN(n9305) );
  XOR2_X1 U17410 ( .A1(n25146), .A2(n25026), .Z(n25239) );
  NAND2_X2 U17412 ( .A1(n10876), .A2(n7495), .ZN(n23303) );
  XOR2_X1 U17414 ( .A1(n38344), .A2(n3151), .Z(n5558) );
  NAND3_X2 U17416 ( .A1(n13665), .A2(n18196), .A3(n37525), .ZN(n9912) );
  NOR2_X2 U17419 ( .A1(n22935), .A2(n8491), .ZN(n8386) );
  NAND2_X1 U17420 ( .A1(n6226), .A2(n36992), .ZN(n224) );
  NAND2_X1 U17425 ( .A1(n34068), .A2(n38114), .ZN(n31200) );
  XOR2_X1 U17429 ( .A1(n16765), .A2(n16766), .Z(n24164) );
  NOR2_X2 U17430 ( .A1(n28728), .A2(n28473), .ZN(n8092) );
  NAND2_X2 U17434 ( .A1(n27878), .A2(n4788), .ZN(n28728) );
  NAND2_X2 U17435 ( .A1(n37028), .A2(n37300), .ZN(n26236) );
  XOR2_X1 U17436 ( .A1(n22439), .A2(n22531), .Z(n22640) );
  NAND2_X2 U17439 ( .A1(n13614), .A2(n31476), .ZN(n22531) );
  INV_X2 U17445 ( .I(n8430), .ZN(n24789) );
  NAND2_X2 U17447 ( .A1(n39354), .A2(n32057), .ZN(n8430) );
  INV_X4 U17451 ( .I(n1755), .ZN(n34389) );
  XOR2_X1 U17453 ( .A1(n38110), .A2(n38109), .Z(n2778) );
  XOR2_X1 U17457 ( .A1(n2184), .A2(n2185), .Z(n38110) );
  BUF_X4 U17460 ( .I(n8205), .Z(n38609) );
  INV_X2 U17463 ( .I(n19930), .ZN(n1439) );
  XOR2_X1 U17471 ( .A1(n6848), .A2(n6796), .Z(n19930) );
  NAND2_X2 U17472 ( .A1(n30132), .A2(n18241), .ZN(n19098) );
  NAND3_X2 U17474 ( .A1(n26422), .A2(n3449), .A3(n37055), .ZN(n38394) );
  XOR2_X1 U17477 ( .A1(n36645), .A2(n6475), .Z(n32537) );
  XOR2_X1 U17478 ( .A1(n38111), .A2(n24015), .Z(n24317) );
  BUF_X4 U17485 ( .I(n12237), .Z(n38855) );
  NAND2_X2 U17490 ( .A1(n17989), .A2(n17499), .ZN(n34283) );
  NAND2_X2 U17491 ( .A1(n33359), .A2(n34283), .ZN(n38339) );
  INV_X2 U17492 ( .I(n27244), .ZN(n34606) );
  NAND3_X2 U17495 ( .A1(n15495), .A2(n20954), .A3(n23232), .ZN(n24079) );
  AOI21_X2 U17497 ( .A1(n20399), .A2(n1089), .B(n36549), .ZN(n36711) );
  NOR2_X1 U17501 ( .A1(n33289), .A2(n19857), .ZN(n8987) );
  NAND3_X2 U17502 ( .A1(n38112), .A2(n11501), .A3(n39786), .ZN(n17) );
  NAND2_X2 U17508 ( .A1(n33603), .A2(n11375), .ZN(n38112) );
  XOR2_X1 U17509 ( .A1(n16336), .A2(n16334), .Z(n33777) );
  NAND2_X2 U17510 ( .A1(n15733), .A2(n36473), .ZN(n16334) );
  AND2_X1 U17516 ( .A1(n23102), .A2(n9677), .Z(n3411) );
  OAI21_X2 U17519 ( .A1(n15459), .A2(n5051), .B(n38113), .ZN(n11241) );
  NOR2_X1 U17521 ( .A1(n38119), .A2(n23358), .ZN(n38114) );
  AOI21_X2 U17522 ( .A1(n28415), .A2(n34667), .B(n35199), .ZN(n38311) );
  NAND4_X2 U17523 ( .A1(n34192), .A2(n9364), .A3(n9357), .A4(n7595), .ZN(
        n18211) );
  NAND2_X2 U17526 ( .A1(n26125), .A2(n4190), .ZN(n39569) );
  NAND2_X1 U17527 ( .A1(n38116), .A2(n23487), .ZN(n23305) );
  OAI22_X1 U17533 ( .A1(n23488), .A2(n1632), .B1(n32017), .B2(n37774), .ZN(
        n38116) );
  XOR2_X1 U17534 ( .A1(n10616), .A2(n38117), .Z(n4059) );
  XOR2_X1 U17535 ( .A1(n18600), .A2(n25214), .Z(n38117) );
  XOR2_X1 U17536 ( .A1(n8546), .A2(n38118), .Z(n8544) );
  NOR2_X1 U17541 ( .A1(n33263), .A2(n37393), .ZN(n38432) );
  BUF_X4 U17544 ( .I(n29936), .Z(n16224) );
  INV_X4 U17547 ( .I(n4190), .ZN(n39454) );
  XOR2_X1 U17548 ( .A1(n27749), .A2(n37812), .Z(n38121) );
  XOR2_X1 U17550 ( .A1(n19642), .A2(n27738), .Z(n27502) );
  AOI22_X2 U17552 ( .A1(n7079), .A2(n2888), .B1(n25743), .B2(n33795), .ZN(
        n7080) );
  NAND2_X2 U17553 ( .A1(n18213), .A2(n18215), .ZN(n38122) );
  NAND3_X2 U17555 ( .A1(n38123), .A2(n17715), .A3(n30805), .ZN(n39104) );
  INV_X4 U17556 ( .I(n12306), .ZN(n36234) );
  OAI21_X2 U17557 ( .A1(n22969), .A2(n45), .B(n38124), .ZN(n23592) );
  OAI21_X1 U17559 ( .A1(n35994), .A2(n6009), .B(n13572), .ZN(n38124) );
  NAND2_X1 U17560 ( .A1(n34685), .A2(n25888), .ZN(n25850) );
  NAND2_X2 U17570 ( .A1(n7583), .A2(n33346), .ZN(n25489) );
  NAND2_X2 U17571 ( .A1(n38125), .A2(n34395), .ZN(n14956) );
  AOI21_X2 U17572 ( .A1(n37128), .A2(n7486), .B(n38126), .ZN(n38125) );
  NOR2_X2 U17575 ( .A1(n7486), .A2(n28073), .ZN(n38126) );
  NAND2_X2 U17581 ( .A1(n4584), .A2(n4581), .ZN(n10171) );
  NOR2_X1 U17585 ( .A1(n21840), .A2(n21903), .ZN(n21624) );
  OR2_X1 U17587 ( .A1(n17217), .A2(n856), .Z(n9061) );
  AND2_X1 U17592 ( .A1(n8849), .A2(n8850), .Z(n38127) );
  AOI21_X2 U17593 ( .A1(n24832), .A2(n24573), .B(n38128), .ZN(n16864) );
  OAI21_X2 U17594 ( .A1(n16208), .A2(n24832), .B(n24574), .ZN(n38128) );
  XNOR2_X1 U17595 ( .A1(n17310), .A2(n22552), .ZN(n6630) );
  OAI21_X2 U17596 ( .A1(n6582), .A2(n36946), .B(n22159), .ZN(n22552) );
  AOI21_X2 U17599 ( .A1(n38129), .A2(n19734), .B(n19962), .ZN(n2243) );
  NAND2_X1 U17600 ( .A1(n8229), .A2(n38429), .ZN(n39522) );
  NOR2_X2 U17601 ( .A1(n16733), .A2(n38130), .ZN(n16732) );
  NAND2_X2 U17602 ( .A1(n26870), .A2(n7975), .ZN(n27006) );
  XOR2_X1 U17605 ( .A1(n36778), .A2(n22580), .Z(n2471) );
  XOR2_X1 U17607 ( .A1(n20454), .A2(n27687), .Z(n27490) );
  XOR2_X1 U17608 ( .A1(n11399), .A2(n32505), .Z(n16425) );
  NAND2_X2 U17610 ( .A1(n19435), .A2(n20157), .ZN(n11526) );
  XOR2_X1 U17614 ( .A1(n27758), .A2(n27534), .Z(n3557) );
  NAND2_X2 U17620 ( .A1(n13400), .A2(n35790), .ZN(n27758) );
  XOR2_X1 U17622 ( .A1(n27667), .A2(n31061), .Z(n12304) );
  NAND2_X2 U17623 ( .A1(n15768), .A2(n37096), .ZN(n29361) );
  XOR2_X1 U17640 ( .A1(n22748), .A2(n22747), .Z(n5338) );
  XOR2_X1 U17642 ( .A1(n16804), .A2(n16805), .Z(n18186) );
  XOR2_X1 U17643 ( .A1(n27541), .A2(n34986), .Z(n16805) );
  OR2_X1 U17645 ( .A1(n25836), .A2(n19580), .Z(n18214) );
  AOI22_X2 U17647 ( .A1(n5164), .A2(n927), .B1(n26090), .B2(n37239), .ZN(
        n38131) );
  XOR2_X1 U17650 ( .A1(n1886), .A2(n1883), .Z(n10938) );
  NAND2_X2 U17652 ( .A1(n25975), .A2(n6056), .ZN(n15524) );
  NOR3_X2 U17654 ( .A1(n10882), .A2(n1548), .A3(n31780), .ZN(n32011) );
  NAND2_X2 U17656 ( .A1(n38132), .A2(n39622), .ZN(n25836) );
  XOR2_X1 U17657 ( .A1(n2782), .A2(n38181), .Z(n38133) );
  NAND2_X2 U17661 ( .A1(n24740), .A2(n24821), .ZN(n35785) );
  OAI21_X2 U17662 ( .A1(n14167), .A2(n24820), .B(n14166), .ZN(n24740) );
  BUF_X4 U17663 ( .I(n9920), .Z(n9321) );
  NAND2_X2 U17666 ( .A1(n28748), .A2(n9917), .ZN(n28623) );
  NAND2_X2 U17670 ( .A1(n8535), .A2(n8534), .ZN(n27633) );
  NAND2_X2 U17671 ( .A1(n23505), .A2(n20276), .ZN(n23596) );
  NOR2_X2 U17672 ( .A1(n23051), .A2(n4565), .ZN(n35932) );
  OR2_X1 U17675 ( .A1(n13717), .A2(n26001), .Z(n2657) );
  XOR2_X1 U17683 ( .A1(n38134), .A2(n30126), .Z(Ciphertext[166]) );
  NAND3_X2 U17685 ( .A1(n36005), .A2(n36420), .A3(n9261), .ZN(n38134) );
  BUF_X4 U17687 ( .I(n26459), .Z(n26909) );
  INV_X2 U17688 ( .I(n38135), .ZN(n39815) );
  XOR2_X1 U17689 ( .A1(n8567), .A2(n8565), .Z(n38135) );
  XOR2_X1 U17694 ( .A1(n38136), .A2(n1769), .Z(n32985) );
  BUF_X2 U17700 ( .I(n17890), .Z(n38137) );
  NOR2_X2 U17701 ( .A1(n31264), .A2(n37102), .ZN(n38138) );
  INV_X2 U17705 ( .I(n22510), .ZN(n22778) );
  NAND2_X2 U17713 ( .A1(n20256), .A2(n33655), .ZN(n22510) );
  AOI22_X1 U17718 ( .A1(n30098), .A2(n2489), .B1(n2484), .B2(n35175), .ZN(
        n36182) );
  NAND2_X2 U17719 ( .A1(n36736), .A2(n8730), .ZN(n38653) );
  XOR2_X1 U17722 ( .A1(n15305), .A2(n38139), .Z(n20883) );
  XOR2_X1 U17725 ( .A1(n15303), .A2(n15304), .Z(n38139) );
  XOR2_X1 U17726 ( .A1(n23973), .A2(n18175), .Z(n23937) );
  NAND2_X2 U17727 ( .A1(n39506), .A2(n32487), .ZN(n23973) );
  XOR2_X1 U17729 ( .A1(n35878), .A2(n22727), .Z(n13561) );
  INV_X1 U17734 ( .I(n38512), .ZN(n35374) );
  OAI21_X1 U17738 ( .A1(n33104), .A2(n12146), .B(n2091), .ZN(n36444) );
  INV_X2 U17739 ( .I(n17653), .ZN(n2848) );
  NAND2_X2 U17740 ( .A1(n32391), .A2(n5282), .ZN(n17891) );
  NOR3_X2 U17741 ( .A1(n35313), .A2(n31661), .A3(n36885), .ZN(n32054) );
  NAND3_X2 U17753 ( .A1(n20498), .A2(n29722), .A3(n17708), .ZN(n29714) );
  AND2_X1 U17754 ( .A1(n30184), .A2(n17996), .Z(n12301) );
  NAND2_X2 U17762 ( .A1(n23255), .A2(n33702), .ZN(n38175) );
  INV_X2 U17763 ( .I(n25813), .ZN(n1014) );
  OAI21_X2 U17765 ( .A1(n38775), .A2(n35580), .B(n38774), .ZN(n26650) );
  NOR2_X2 U17773 ( .A1(n15623), .A2(n3983), .ZN(n36224) );
  AOI22_X2 U17774 ( .A1(n26132), .A2(n1014), .B1(n6749), .B2(n25936), .ZN(
        n39625) );
  INV_X2 U17775 ( .I(n26459), .ZN(n26719) );
  NAND2_X2 U17782 ( .A1(n988), .A2(n27894), .ZN(n13955) );
  INV_X2 U17793 ( .I(n8412), .ZN(n27440) );
  AOI21_X2 U17796 ( .A1(n2868), .A2(n28224), .B(n28229), .ZN(n15571) );
  OAI22_X2 U17797 ( .A1(n33001), .A2(n32948), .B1(n36711), .B2(n38092), .ZN(
        n38402) );
  BUF_X4 U17801 ( .I(n38402), .Z(n32926) );
  NAND2_X2 U17804 ( .A1(n2740), .A2(n12443), .ZN(n12488) );
  NAND2_X2 U17805 ( .A1(n691), .A2(n29555), .ZN(n29547) );
  OR2_X1 U17806 ( .A1(n29437), .A2(n29438), .Z(n18495) );
  INV_X4 U17814 ( .I(n13366), .ZN(n28213) );
  OAI21_X1 U17815 ( .A1(n8307), .A2(n1198), .B(n38804), .ZN(n33161) );
  AOI22_X2 U17818 ( .A1(n12478), .A2(n7866), .B1(n1531), .B2(n25692), .ZN(
        n8223) );
  AOI22_X2 U17819 ( .A1(n8965), .A2(n38119), .B1(n8757), .B2(n23358), .ZN(
        n6517) );
  NAND2_X2 U17820 ( .A1(n8407), .A2(n25782), .ZN(n35786) );
  INV_X2 U17822 ( .I(n30257), .ZN(n30258) );
  INV_X2 U17828 ( .I(n23540), .ZN(n10495) );
  NAND2_X1 U17829 ( .A1(n38266), .A2(n36654), .ZN(n22825) );
  NAND2_X2 U17832 ( .A1(n945), .A2(n27233), .ZN(n7471) );
  AOI21_X2 U17833 ( .A1(n986), .A2(n20977), .B(n38443), .ZN(n8993) );
  NAND2_X2 U17835 ( .A1(n34740), .A2(n34739), .ZN(n34738) );
  NOR2_X2 U17836 ( .A1(n20010), .A2(n28279), .ZN(n30773) );
  AOI21_X2 U17837 ( .A1(n38404), .A2(n38702), .B(n2597), .ZN(n30550) );
  NOR3_X2 U17838 ( .A1(n310), .A2(n16461), .A3(n28200), .ZN(n35309) );
  NAND2_X2 U17840 ( .A1(n25692), .A2(n12478), .ZN(n12382) );
  NAND2_X2 U17847 ( .A1(n31486), .A2(n39768), .ZN(n38143) );
  OAI21_X1 U17848 ( .A1(n6204), .A2(n1407), .B(n31444), .ZN(n29194) );
  BUF_X4 U17857 ( .I(n28231), .Z(n19366) );
  INV_X2 U17858 ( .I(n29998), .ZN(n29949) );
  OAI22_X2 U17859 ( .A1(n30365), .A2(n1093), .B1(n38824), .B2(n38120), .ZN(
        n18023) );
  INV_X2 U17861 ( .I(n29781), .ZN(n1408) );
  NAND2_X1 U17863 ( .A1(n6831), .A2(n36375), .ZN(n38632) );
  NAND2_X2 U17866 ( .A1(n13151), .A2(n36791), .ZN(n13372) );
  OR2_X1 U17868 ( .A1(n5881), .A2(n5884), .Z(n38140) );
  INV_X1 U17870 ( .I(n25246), .ZN(n38895) );
  INV_X1 U17872 ( .I(n39793), .ZN(n25848) );
  NOR2_X1 U17876 ( .A1(n20157), .A2(n32977), .ZN(n30370) );
  NOR3_X1 U17882 ( .A1(n32977), .A2(n28049), .A3(n20157), .ZN(n10166) );
  NAND2_X1 U17884 ( .A1(n36391), .A2(n14601), .ZN(n12986) );
  INV_X1 U17893 ( .I(n29559), .ZN(n39003) );
  AOI21_X1 U17895 ( .A1(n27416), .A2(n19564), .B(n27110), .ZN(n27111) );
  NOR2_X1 U17896 ( .A1(n28131), .A2(n2868), .ZN(n15568) );
  CLKBUF_X4 U17900 ( .I(n20522), .Z(n33784) );
  NAND2_X1 U17902 ( .A1(n30241), .A2(n20525), .ZN(n31237) );
  NAND2_X1 U17903 ( .A1(n859), .A2(n26935), .ZN(n13777) );
  NAND2_X1 U17910 ( .A1(n29354), .A2(n29422), .ZN(n6865) );
  CLKBUF_X4 U17914 ( .I(n33961), .Z(n2782) );
  INV_X1 U17915 ( .I(n27802), .ZN(n1457) );
  NOR2_X1 U17917 ( .A1(n19475), .A2(n20160), .ZN(n38142) );
  INV_X1 U17918 ( .I(n29204), .ZN(n15601) );
  NAND2_X1 U17920 ( .A1(n25962), .A2(n16407), .ZN(n26027) );
  NAND3_X1 U17922 ( .A1(n27866), .A2(n19657), .A3(n9553), .ZN(n27685) );
  OR2_X1 U17932 ( .A1(n29869), .A2(n773), .Z(n5973) );
  NAND2_X1 U17933 ( .A1(n38506), .A2(n14030), .ZN(n38145) );
  NOR2_X1 U17934 ( .A1(n28142), .A2(n20184), .ZN(n20500) );
  CLKBUF_X4 U17935 ( .I(n28473), .Z(n5396) );
  CLKBUF_X4 U17936 ( .I(n17777), .Z(n11676) );
  NAND2_X1 U17945 ( .A1(n9802), .A2(n19580), .ZN(n30957) );
  NAND2_X1 U17948 ( .A1(n29701), .A2(n29700), .ZN(n16385) );
  OAI21_X1 U17951 ( .A1(n29699), .A2(n29700), .B(n29698), .ZN(n28513) );
  NAND2_X1 U17953 ( .A1(n30034), .A2(n30024), .ZN(n10942) );
  INV_X2 U17954 ( .I(n4879), .ZN(n29843) );
  NOR2_X1 U17955 ( .A1(n4879), .A2(n20793), .ZN(n3379) );
  OR2_X1 U17958 ( .A1(n39126), .A2(n32822), .Z(n5863) );
  NOR2_X1 U17961 ( .A1(n16154), .A2(n28143), .ZN(n7255) );
  AOI22_X1 U17962 ( .A1(n25420), .A2(n18031), .B1(n12381), .B2(n13166), .ZN(
        n38628) );
  INV_X1 U17967 ( .I(n21546), .ZN(n1692) );
  INV_X2 U17972 ( .I(n19696), .ZN(n19452) );
  BUF_X2 U17975 ( .I(n4382), .Z(n32385) );
  NOR2_X1 U17976 ( .A1(n39334), .A2(n28738), .ZN(n28743) );
  INV_X1 U17988 ( .I(n28286), .ZN(n28161) );
  NAND2_X1 U17992 ( .A1(n31143), .A2(n39731), .ZN(n38148) );
  NAND3_X1 U17993 ( .A1(n29712), .A2(n29719), .A3(n14337), .ZN(n29716) );
  OR2_X2 U17994 ( .A1(n9118), .A2(n26459), .Z(n26927) );
  AND2_X1 U17995 ( .A1(n33960), .A2(n15774), .Z(n33185) );
  CLKBUF_X1 U17997 ( .I(n7464), .Z(n34492) );
  NOR2_X1 U18000 ( .A1(n24169), .A2(n24396), .ZN(n23844) );
  NAND3_X1 U18001 ( .A1(n1142), .A2(n11307), .A3(n20782), .ZN(n23086) );
  NOR2_X1 U18002 ( .A1(n25942), .A2(n6579), .ZN(n9714) );
  OAI21_X1 U18004 ( .A1(n10800), .A2(n35690), .B(n10046), .ZN(n10799) );
  INV_X1 U18006 ( .I(n36571), .ZN(n34482) );
  INV_X2 U18007 ( .I(n26780), .ZN(n26948) );
  NOR2_X1 U18010 ( .A1(n28478), .A2(n1196), .ZN(n28479) );
  NAND2_X1 U18011 ( .A1(n1414), .A2(n1196), .ZN(n33229) );
  OAI21_X2 U18014 ( .A1(n20050), .A2(n20051), .B(n20049), .ZN(n38149) );
  OAI21_X1 U18026 ( .A1(n20050), .A2(n20051), .B(n20049), .ZN(n20210) );
  OR2_X1 U18044 ( .A1(n24536), .A2(n7705), .Z(n19532) );
  AND3_X1 U18053 ( .A1(n19398), .A2(n7705), .A3(n25683), .Z(n34025) );
  NAND2_X1 U18054 ( .A1(n29375), .A2(n37100), .ZN(n19244) );
  NAND2_X1 U18055 ( .A1(n29310), .A2(n29384), .ZN(n36994) );
  NAND2_X1 U18056 ( .A1(n35508), .A2(n36133), .ZN(n25534) );
  NOR2_X1 U18057 ( .A1(n32366), .A2(n1294), .ZN(n8214) );
  NAND2_X1 U18058 ( .A1(n11491), .A2(n11492), .ZN(n38150) );
  INV_X1 U18059 ( .I(n36523), .ZN(n36050) );
  INV_X1 U18063 ( .I(n7106), .ZN(n31425) );
  NAND3_X1 U18064 ( .A1(n7106), .A2(n12415), .A3(n26967), .ZN(n6797) );
  OR2_X1 U18066 ( .A1(n14387), .A2(n30217), .Z(n36739) );
  INV_X2 U18076 ( .I(n33963), .ZN(n10569) );
  NAND2_X1 U18079 ( .A1(n13370), .A2(n14856), .ZN(n13834) );
  OAI21_X1 U18080 ( .A1(n27927), .A2(n27926), .B(n36414), .ZN(n8910) );
  OR2_X1 U18081 ( .A1(n12371), .A2(n12372), .Z(n38151) );
  NAND2_X1 U18083 ( .A1(n11787), .A2(n11785), .ZN(n35029) );
  OAI21_X2 U18084 ( .A1(n27258), .A2(n27257), .B(n27256), .ZN(n38152) );
  OAI21_X1 U18085 ( .A1(n27258), .A2(n27257), .B(n27256), .ZN(n38153) );
  OAI21_X1 U18087 ( .A1(n27258), .A2(n27257), .B(n27256), .ZN(n27717) );
  NOR2_X2 U18089 ( .A1(n32697), .A2(n7588), .ZN(n27257) );
  CLKBUF_X4 U18093 ( .I(n26888), .Z(n27337) );
  AND2_X1 U18108 ( .A1(n2792), .A2(n29810), .Z(n14009) );
  NAND2_X2 U18111 ( .A1(n33563), .A2(n21164), .ZN(n38154) );
  INV_X1 U18114 ( .I(n18908), .ZN(n2113) );
  INV_X2 U18117 ( .I(n378), .ZN(n14793) );
  NAND2_X1 U18120 ( .A1(n378), .A2(n36922), .ZN(n36815) );
  NOR2_X1 U18121 ( .A1(n36922), .A2(n378), .ZN(n30644) );
  NAND2_X1 U18122 ( .A1(n378), .A2(n33293), .ZN(n7404) );
  OAI21_X1 U18124 ( .A1(n10338), .A2(n10524), .B(n8311), .ZN(n26270) );
  NOR2_X1 U18135 ( .A1(n27141), .A2(n10338), .ZN(n38494) );
  INV_X2 U18136 ( .I(n8000), .ZN(n10338) );
  OR3_X1 U18137 ( .A1(n8960), .A2(n27624), .A3(n16576), .Z(n7983) );
  NOR2_X1 U18138 ( .A1(n32186), .A2(n16576), .ZN(n28422) );
  OAI21_X1 U18139 ( .A1(n28328), .A2(n28327), .B(n39423), .ZN(n38970) );
  NOR2_X1 U18144 ( .A1(n39423), .A2(n39422), .ZN(n35548) );
  INV_X1 U18145 ( .I(n38461), .ZN(n5334) );
  NAND2_X1 U18148 ( .A1(n34386), .A2(n9823), .ZN(n38623) );
  INV_X1 U18162 ( .I(n15625), .ZN(n25277) );
  OR2_X2 U18165 ( .A1(n37079), .A2(n8395), .Z(n28043) );
  NOR2_X1 U18168 ( .A1(n27250), .A2(n33503), .ZN(n11854) );
  AOI21_X1 U18169 ( .A1(n13907), .A2(n310), .B(n13906), .ZN(n13905) );
  INV_X1 U18175 ( .I(n35705), .ZN(n1605) );
  NAND2_X1 U18182 ( .A1(n609), .A2(n35705), .ZN(n24451) );
  OR2_X1 U18185 ( .A1(n16459), .A2(n35705), .Z(n6933) );
  INV_X1 U18187 ( .I(n29336), .ZN(n38156) );
  AND2_X1 U18191 ( .A1(n32790), .A2(n14858), .Z(n29328) );
  CLKBUF_X12 U18197 ( .I(n29336), .Z(n32790) );
  OAI21_X1 U18198 ( .A1(n19669), .A2(n20691), .B(n27498), .ZN(n16856) );
  OAI21_X1 U18200 ( .A1(n6975), .A2(n27027), .B(n27251), .ZN(n33160) );
  NAND2_X1 U18202 ( .A1(n13088), .A2(n26988), .ZN(n6261) );
  NAND2_X1 U18207 ( .A1(n29800), .A2(n29799), .ZN(n5145) );
  NOR2_X1 U18208 ( .A1(n29800), .A2(n3614), .ZN(n39062) );
  NAND2_X1 U18214 ( .A1(n35273), .A2(n29616), .ZN(n29624) );
  NAND3_X2 U18216 ( .A1(n8031), .A2(n37728), .A3(n8030), .ZN(n10978) );
  CLKBUF_X4 U18219 ( .I(n833), .Z(n7284) );
  XNOR2_X1 U18220 ( .A1(n23832), .A2(n24050), .ZN(n17140) );
  XOR2_X1 U18231 ( .A1(n2805), .A2(n38157), .Z(n36380) );
  XOR2_X1 U18246 ( .A1(n23887), .A2(n678), .Z(n38157) );
  NOR2_X1 U18248 ( .A1(n28163), .A2(n5988), .ZN(n885) );
  BUF_X2 U18249 ( .I(n28163), .Z(n32705) );
  AOI21_X1 U18251 ( .A1(n28163), .A2(n16363), .B(n27979), .ZN(n35931) );
  CLKBUF_X1 U18252 ( .I(n30184), .Z(n31846) );
  AOI21_X1 U18256 ( .A1(n38683), .A2(n15317), .B(n26901), .ZN(n5589) );
  NAND3_X1 U18258 ( .A1(n26903), .A2(n26901), .A3(n11616), .ZN(n34843) );
  NAND2_X1 U18259 ( .A1(n34000), .A2(n1402), .ZN(n39312) );
  NOR2_X1 U18260 ( .A1(n39313), .A2(n34000), .ZN(n32335) );
  NAND2_X1 U18261 ( .A1(n8519), .A2(n22196), .ZN(n3435) );
  OAI21_X1 U18266 ( .A1(n5509), .A2(n13851), .B(n13322), .ZN(n13321) );
  NAND2_X1 U18270 ( .A1(n15963), .A2(n3988), .ZN(n35030) );
  AOI22_X1 U18273 ( .A1(n33139), .A2(n9627), .B1(n29333), .B2(n29340), .ZN(
        n31801) );
  INV_X2 U18279 ( .I(n12543), .ZN(n4950) );
  NOR2_X1 U18282 ( .A1(n26841), .A2(n36392), .ZN(n38798) );
  CLKBUF_X4 U18284 ( .I(n20595), .Z(n1548) );
  OAI22_X1 U18287 ( .A1(n19452), .A2(n1548), .B1(n16836), .B2(n16246), .ZN(
        n25402) );
  OAI21_X1 U18304 ( .A1(n1548), .A2(n953), .B(n16246), .ZN(n3877) );
  NAND2_X2 U18305 ( .A1(n32755), .A2(n38333), .ZN(n38158) );
  NOR2_X2 U18309 ( .A1(n4941), .A2(n30837), .ZN(n38159) );
  NAND2_X1 U18311 ( .A1(n32755), .A2(n38333), .ZN(n38964) );
  NAND2_X2 U18312 ( .A1(n32756), .A2(n32757), .ZN(n32755) );
  CLKBUF_X12 U18315 ( .I(n20883), .Z(n10346) );
  NOR2_X1 U18318 ( .A1(n13442), .A2(n35179), .ZN(n29566) );
  INV_X1 U18324 ( .I(n5031), .ZN(n26117) );
  NAND2_X1 U18329 ( .A1(n29889), .A2(n29888), .ZN(n11787) );
  NAND2_X1 U18330 ( .A1(n26905), .A2(n26564), .ZN(n15880) );
  NAND3_X1 U18335 ( .A1(n30858), .A2(n28444), .A3(n30857), .ZN(n27972) );
  NOR2_X1 U18339 ( .A1(n10746), .A2(n2456), .ZN(n9064) );
  NAND2_X1 U18340 ( .A1(n38871), .A2(n13890), .ZN(n38160) );
  AND2_X1 U18345 ( .A1(n26048), .A2(n26019), .Z(n26050) );
  NOR2_X1 U18357 ( .A1(n18281), .A2(n7905), .ZN(n28705) );
  NOR2_X1 U18360 ( .A1(n39019), .A2(n17286), .ZN(n29877) );
  NAND4_X1 U18362 ( .A1(n1560), .A2(n11601), .A3(n14874), .A4(n24754), .ZN(
        n11605) );
  OAI21_X1 U18363 ( .A1(n3631), .A2(n2121), .B(n38784), .ZN(n28923) );
  NAND2_X1 U18364 ( .A1(n9328), .A2(n9327), .ZN(n38162) );
  NAND2_X2 U18370 ( .A1(n27906), .A2(n9897), .ZN(n9327) );
  OR2_X2 U18372 ( .A1(n139), .A2(n32925), .Z(n38163) );
  OR2_X2 U18376 ( .A1(n139), .A2(n32925), .Z(n38164) );
  INV_X1 U18377 ( .I(n26591), .ZN(n15676) );
  NAND2_X1 U18378 ( .A1(n33200), .A2(n33199), .ZN(n27890) );
  NOR2_X1 U18380 ( .A1(n6892), .A2(n28609), .ZN(n28335) );
  OAI21_X1 U18381 ( .A1(n12238), .A2(n12611), .B(n28609), .ZN(n35574) );
  NAND3_X1 U18382 ( .A1(n178), .A2(n25670), .A3(n18164), .ZN(n10936) );
  NOR2_X1 U18383 ( .A1(n1066), .A2(n16559), .ZN(n35997) );
  INV_X1 U18385 ( .I(n9246), .ZN(n8045) );
  NAND2_X1 U18389 ( .A1(n12943), .A2(n9839), .ZN(n29365) );
  INV_X2 U18393 ( .I(n9839), .ZN(n13981) );
  AOI21_X2 U18399 ( .A1(n28623), .A2(n19161), .B(n977), .ZN(n13656) );
  INV_X2 U18400 ( .I(n28745), .ZN(n977) );
  INV_X1 U18404 ( .I(n36275), .ZN(n18190) );
  INV_X1 U18407 ( .I(n11939), .ZN(n31912) );
  OR3_X1 U18408 ( .A1(n968), .A2(n939), .A3(n3462), .Z(n30401) );
  CLKBUF_X4 U18413 ( .I(n28130), .Z(n2868) );
  INV_X1 U18418 ( .I(n39456), .ZN(n34479) );
  OAI21_X1 U18421 ( .A1(n21724), .A2(n4925), .B(n4924), .ZN(n21725) );
  INV_X1 U18425 ( .I(n12537), .ZN(n10058) );
  NOR2_X1 U18426 ( .A1(n11443), .A2(n27010), .ZN(n32490) );
  INV_X2 U18427 ( .I(n14557), .ZN(n30047) );
  CLKBUF_X4 U18428 ( .I(n14557), .Z(n36850) );
  AOI21_X2 U18437 ( .A1(n3798), .A2(n3799), .B(n33519), .ZN(n38165) );
  NAND2_X2 U18443 ( .A1(n977), .A2(n28746), .ZN(n3798) );
  INV_X2 U18454 ( .I(n29777), .ZN(n39313) );
  INV_X2 U18457 ( .I(n28398), .ZN(n16691) );
  NAND2_X1 U18460 ( .A1(n28398), .A2(n16303), .ZN(n16304) );
  NAND2_X1 U18463 ( .A1(n28398), .A2(n28755), .ZN(n27909) );
  OR2_X1 U18465 ( .A1(n16039), .A2(n15466), .Z(n21617) );
  NAND2_X1 U18466 ( .A1(n28422), .A2(n27624), .ZN(n31087) );
  INV_X1 U18469 ( .I(n16324), .ZN(n5290) );
  XNOR2_X1 U18470 ( .A1(n36254), .A2(n36255), .ZN(n38167) );
  NAND2_X1 U18474 ( .A1(n3944), .A2(n14448), .ZN(n38727) );
  NAND2_X1 U18475 ( .A1(n12488), .A2(n982), .ZN(n3981) );
  NAND2_X1 U18477 ( .A1(n12488), .A2(n2262), .ZN(n12487) );
  OAI21_X1 U18494 ( .A1(n33107), .A2(n33106), .B(n30953), .ZN(n18624) );
  CLKBUF_X12 U18496 ( .I(n2147), .Z(n30953) );
  NAND2_X1 U18498 ( .A1(n8314), .A2(n36385), .ZN(n1845) );
  OR2_X2 U18500 ( .A1(n26779), .A2(n20063), .Z(n26848) );
  NAND2_X1 U18501 ( .A1(n34857), .A2(n39140), .ZN(n39822) );
  NOR2_X1 U18502 ( .A1(n27963), .A2(n28050), .ZN(n10515) );
  NAND2_X1 U18503 ( .A1(n37754), .A2(n28279), .ZN(n27621) );
  INV_X1 U18504 ( .I(n12081), .ZN(n1397) );
  XOR2_X1 U18508 ( .A1(n38169), .A2(n38170), .Z(n34251) );
  XNOR2_X1 U18509 ( .A1(n27773), .A2(n19561), .ZN(n38169) );
  XOR2_X1 U18511 ( .A1(n9315), .A2(n15273), .Z(n38170) );
  NOR2_X1 U18512 ( .A1(n773), .A2(n1063), .ZN(n34858) );
  OR2_X1 U18520 ( .A1(n13758), .A2(n26219), .Z(n14862) );
  NAND2_X1 U18522 ( .A1(n27412), .A2(n36200), .ZN(n6353) );
  NOR2_X1 U18524 ( .A1(n21401), .A2(n21644), .ZN(n21720) );
  AOI21_X1 U18530 ( .A1(n21401), .A2(n32704), .B(n21909), .ZN(n13239) );
  NAND2_X1 U18534 ( .A1(n20120), .A2(n2752), .ZN(n38774) );
  BUF_X2 U18535 ( .I(n20120), .Z(n35580) );
  NAND2_X1 U18539 ( .A1(n15594), .A2(n20120), .ZN(n26748) );
  INV_X1 U18542 ( .I(n20120), .ZN(n8478) );
  AOI22_X1 U18545 ( .A1(n29796), .A2(n36096), .B1(n29798), .B2(n29797), .ZN(
        n36808) );
  AOI22_X1 U18548 ( .A1(n29784), .A2(n29783), .B1(n29798), .B2(n29789), .ZN(
        n39278) );
  OR3_X2 U18552 ( .A1(n30195), .A2(n35551), .A3(n4083), .Z(n35329) );
  NAND2_X1 U18555 ( .A1(n21759), .A2(n21545), .ZN(n21549) );
  OAI21_X1 U18556 ( .A1(n17997), .A2(n31846), .B(n2466), .ZN(n2465) );
  OR2_X2 U18560 ( .A1(n37896), .A2(n12519), .Z(n24401) );
  CLKBUF_X4 U18563 ( .I(n29452), .Z(n505) );
  INV_X2 U18565 ( .I(n29869), .ZN(n972) );
  AOI21_X1 U18576 ( .A1(n36225), .A2(n19476), .B(n11826), .ZN(n2769) );
  AOI21_X1 U18587 ( .A1(n1802), .A2(n21017), .B(n33945), .ZN(n38171) );
  AOI21_X1 U18589 ( .A1(n1802), .A2(n21017), .B(n33945), .ZN(n35317) );
  NOR2_X1 U18593 ( .A1(n37619), .A2(n12537), .ZN(n13403) );
  NAND2_X1 U18594 ( .A1(n35745), .A2(n15616), .ZN(n31146) );
  NAND3_X1 U18603 ( .A1(n17661), .A2(n27218), .A3(n15616), .ZN(n4948) );
  NOR2_X1 U18606 ( .A1(n4649), .A2(n1209), .ZN(n10084) );
  NOR2_X1 U18612 ( .A1(n22295), .A2(n5061), .ZN(n5127) );
  INV_X1 U18613 ( .I(n8988), .ZN(n38853) );
  INV_X1 U18617 ( .I(n12707), .ZN(n14128) );
  CLKBUF_X12 U18619 ( .I(n39528), .Z(n38951) );
  AOI21_X1 U18634 ( .A1(n37075), .A2(n8253), .B(n33662), .ZN(n2381) );
  AOI21_X1 U18635 ( .A1(n33082), .A2(n22907), .B(n22906), .ZN(n23391) );
  NAND2_X1 U18641 ( .A1(n6691), .A2(n14560), .ZN(n32042) );
  INV_X1 U18646 ( .I(n28484), .ZN(n28391) );
  NAND2_X1 U18652 ( .A1(n11089), .A2(n11087), .ZN(n38174) );
  INV_X1 U18654 ( .I(n11330), .ZN(n28609) );
  INV_X1 U18659 ( .I(n32623), .ZN(n3328) );
  NAND2_X1 U18661 ( .A1(n30244), .A2(n30245), .ZN(n30246) );
  NOR2_X1 U18668 ( .A1(n30245), .A2(n39187), .ZN(n10977) );
  NAND2_X1 U18669 ( .A1(n29815), .A2(n8677), .ZN(n29774) );
  NAND2_X1 U18670 ( .A1(n4520), .A2(n18601), .ZN(n4519) );
  INV_X2 U18671 ( .I(n5457), .ZN(n18601) );
  INV_X1 U18677 ( .I(n25700), .ZN(n31895) );
  NAND2_X1 U18681 ( .A1(n1944), .A2(n7454), .ZN(n28359) );
  NAND2_X1 U18684 ( .A1(n20830), .A2(n29458), .ZN(n20427) );
  OAI21_X1 U18685 ( .A1(n10648), .A2(n10988), .B(n17653), .ZN(n10645) );
  OR2_X2 U18687 ( .A1(n19543), .A2(n20778), .Z(n6349) );
  CLKBUF_X4 U18688 ( .I(n33086), .Z(n38337) );
  NAND2_X1 U18689 ( .A1(n28563), .A2(n1197), .ZN(n38856) );
  INV_X1 U18690 ( .I(n1197), .ZN(n38858) );
  AND2_X2 U18696 ( .A1(n2153), .A2(n33748), .Z(n14250) );
  NAND2_X2 U18698 ( .A1(n8145), .A2(n38651), .ZN(n23255) );
  INV_X2 U18702 ( .I(n17598), .ZN(n9553) );
  NOR2_X2 U18703 ( .A1(n33752), .A2(n6589), .ZN(n38176) );
  XOR2_X1 U18706 ( .A1(n9989), .A2(n26481), .Z(n38177) );
  XOR2_X1 U18715 ( .A1(n6630), .A2(n17513), .Z(n38179) );
  OR3_X2 U18718 ( .A1(n13300), .A2(n38749), .A3(n24515), .Z(n24777) );
  OR2_X2 U18720 ( .A1(n37245), .A2(n34977), .Z(n30412) );
  NAND2_X1 U18722 ( .A1(n8262), .A2(n7542), .ZN(n26647) );
  NAND2_X1 U18723 ( .A1(n1107), .A2(n25860), .ZN(n25708) );
  OAI21_X2 U18727 ( .A1(n4429), .A2(n4428), .B(n4076), .ZN(n38181) );
  NAND2_X1 U18728 ( .A1(n7497), .A2(n20351), .ZN(n22235) );
  OR2_X2 U18730 ( .A1(n4291), .A2(n8544), .Z(n23106) );
  NAND2_X1 U18734 ( .A1(n31234), .A2(n23349), .ZN(n2692) );
  NAND2_X1 U18738 ( .A1(n19332), .A2(n20995), .ZN(n26709) );
  INV_X1 U18742 ( .I(n2273), .ZN(n23317) );
  BUF_X2 U18743 ( .I(n29137), .Z(n30856) );
  NAND3_X1 U18751 ( .A1(n15327), .A2(n15328), .A3(n30057), .ZN(n32668) );
  INV_X1 U18753 ( .I(n29236), .ZN(n38945) );
  NAND2_X1 U18757 ( .A1(n39300), .A2(n20276), .ZN(n39299) );
  INV_X2 U18758 ( .I(n20276), .ZN(n23504) );
  NOR2_X1 U18777 ( .A1(n8190), .A2(n20276), .ZN(n8212) );
  NAND2_X1 U18794 ( .A1(n33455), .A2(n39477), .ZN(n26634) );
  INV_X1 U18796 ( .I(n16080), .ZN(n8305) );
  NAND2_X1 U18797 ( .A1(n3513), .A2(n34717), .ZN(n4033) );
  NOR2_X1 U18798 ( .A1(n1224), .A2(n34717), .ZN(n3514) );
  INV_X1 U18804 ( .I(n25558), .ZN(n38183) );
  NAND3_X1 U18813 ( .A1(n24763), .A2(n1269), .A3(n39098), .ZN(n24767) );
  AND2_X2 U18816 ( .A1(n199), .A2(n198), .Z(n38184) );
  OR2_X2 U18822 ( .A1(n15135), .A2(n2722), .Z(n27584) );
  NAND2_X1 U18825 ( .A1(n15135), .A2(n11020), .ZN(n36222) );
  NOR2_X1 U18829 ( .A1(n6218), .A2(n36539), .ZN(n8268) );
  NOR3_X1 U18837 ( .A1(n18907), .A2(n18402), .A3(n24203), .ZN(n34673) );
  NAND2_X1 U18841 ( .A1(n18907), .A2(n18402), .ZN(n39659) );
  NAND2_X1 U18855 ( .A1(n35985), .A2(n18907), .ZN(n16982) );
  CLKBUF_X12 U18858 ( .I(n13365), .Z(n7789) );
  INV_X2 U18859 ( .I(n21666), .ZN(n21834) );
  AOI21_X2 U18861 ( .A1(n2542), .A2(n25858), .B(n2541), .ZN(n12221) );
  INV_X2 U18863 ( .I(n13213), .ZN(n27251) );
  OAI21_X1 U18864 ( .A1(n24608), .A2(n19255), .B(n31161), .ZN(n36021) );
  OAI21_X1 U18872 ( .A1(n19255), .A2(n31161), .B(n9257), .ZN(n9256) );
  INV_X2 U18875 ( .I(n24232), .ZN(n24176) );
  OR2_X1 U18878 ( .A1(n37632), .A2(n12726), .Z(n11981) );
  OR2_X1 U18880 ( .A1(n15535), .A2(n12726), .Z(n280) );
  OAI22_X1 U18882 ( .A1(n34004), .A2(n39823), .B1(n31526), .B2(n17237), .ZN(
        n26843) );
  OAI21_X1 U18883 ( .A1(n29219), .A2(n31772), .B(n29222), .ZN(n12979) );
  XOR2_X1 U18891 ( .A1(n266), .A2(n17737), .Z(n38186) );
  OR2_X1 U18893 ( .A1(n38186), .A2(n29495), .Z(n20113) );
  OAI21_X1 U18900 ( .A1(n31179), .A2(n23237), .B(n23238), .ZN(n4288) );
  INV_X2 U18901 ( .I(n5554), .ZN(n8262) );
  NOR2_X1 U18902 ( .A1(n15579), .A2(n23461), .ZN(n31179) );
  INV_X2 U18903 ( .I(n15579), .ZN(n23462) );
  INV_X2 U18906 ( .I(n3649), .ZN(n25224) );
  NAND2_X1 U18907 ( .A1(n21476), .A2(n21587), .ZN(n21477) );
  NAND3_X1 U18912 ( .A1(n29677), .A2(n29667), .A3(n31538), .ZN(n29669) );
  NAND2_X1 U18913 ( .A1(n13804), .A2(n15768), .ZN(n13803) );
  INV_X1 U18915 ( .I(n11102), .ZN(n34894) );
  NAND2_X1 U18918 ( .A1(n34154), .A2(n7317), .ZN(n25807) );
  NOR2_X1 U18920 ( .A1(n22170), .A2(n21966), .ZN(n39173) );
  INV_X2 U18931 ( .I(n22170), .ZN(n20238) );
  INV_X2 U18939 ( .I(n38188), .ZN(n26918) );
  AOI21_X1 U18942 ( .A1(n5758), .A2(n5890), .B(n5757), .ZN(n38189) );
  AOI21_X1 U18943 ( .A1(n5758), .A2(n5890), .B(n5757), .ZN(n38190) );
  AOI21_X1 U18944 ( .A1(n5758), .A2(n5890), .B(n5757), .ZN(n5755) );
  NAND2_X1 U18945 ( .A1(n28725), .A2(n17801), .ZN(n5758) );
  XOR2_X1 U18947 ( .A1(n38813), .A2(n30612), .Z(n38191) );
  NAND2_X2 U18955 ( .A1(n38847), .A2(n8406), .ZN(n38192) );
  OAI21_X1 U18956 ( .A1(n28179), .A2(n14389), .B(n28181), .ZN(n32418) );
  NAND2_X2 U18961 ( .A1(n18605), .A2(n30585), .ZN(n38193) );
  BUF_X2 U18963 ( .I(n36150), .Z(n35684) );
  OR2_X2 U18969 ( .A1(n8889), .A2(n37815), .Z(n5111) );
  NOR2_X1 U18975 ( .A1(n4434), .A2(n27314), .ZN(n15917) );
  NOR2_X1 U18980 ( .A1(n18711), .A2(n31202), .ZN(n22138) );
  INV_X1 U18989 ( .I(n36509), .ZN(n27455) );
  OAI21_X2 U18991 ( .A1(n13445), .A2(n37904), .B(n12307), .ZN(n38194) );
  INV_X1 U18994 ( .I(n24106), .ZN(n24168) );
  NAND2_X2 U18995 ( .A1(n28305), .A2(n28304), .ZN(n38195) );
  NOR2_X1 U18997 ( .A1(n27097), .A2(n4771), .ZN(n38568) );
  NAND2_X1 U19000 ( .A1(n33950), .A2(n12478), .ZN(n12368) );
  OAI21_X1 U19005 ( .A1(n8608), .A2(n8607), .B(n25114), .ZN(n8606) );
  NAND3_X1 U19008 ( .A1(n30805), .A2(n14448), .A3(n28546), .ZN(n28470) );
  XOR2_X1 U19009 ( .A1(n3187), .A2(n3188), .Z(n38197) );
  NAND2_X2 U19010 ( .A1(n36535), .A2(n38841), .ZN(n38198) );
  NOR2_X2 U19011 ( .A1(n16911), .A2(n34581), .ZN(n38841) );
  NAND3_X1 U19012 ( .A1(n32960), .A2(n32962), .A3(n7424), .ZN(n30939) );
  OAI21_X1 U19014 ( .A1(n35508), .A2(n25484), .B(n611), .ZN(n25537) );
  OR2_X2 U19015 ( .A1(n3873), .A2(n30503), .Z(n11726) );
  INV_X2 U19018 ( .I(n24805), .ZN(n1026) );
  INV_X1 U19019 ( .I(n24805), .ZN(n38347) );
  INV_X1 U19020 ( .I(n11105), .ZN(n3100) );
  XOR2_X1 U19021 ( .A1(n5177), .A2(n5176), .Z(n38199) );
  NAND2_X2 U19022 ( .A1(n29472), .A2(n29469), .ZN(n38200) );
  OR2_X1 U19026 ( .A1(n38199), .A2(n20960), .Z(n15317) );
  INV_X1 U19039 ( .I(n31627), .ZN(n7714) );
  NAND2_X1 U19040 ( .A1(n11150), .A2(n138), .ZN(n39328) );
  NAND2_X1 U19041 ( .A1(n1108), .A2(n11150), .ZN(n15173) );
  NAND3_X2 U19043 ( .A1(n3399), .A2(n24907), .A3(n812), .ZN(n38201) );
  NAND3_X1 U19045 ( .A1(n3399), .A2(n24907), .A3(n812), .ZN(n25151) );
  XOR2_X1 U19046 ( .A1(n33722), .A2(n39115), .Z(n38202) );
  NAND2_X2 U19049 ( .A1(n31098), .A2(n3846), .ZN(n38203) );
  OAI21_X1 U19053 ( .A1(n35663), .A2(n5035), .B(n3923), .ZN(n38205) );
  NAND2_X1 U19054 ( .A1(n9250), .A2(n9248), .ZN(n38206) );
  INV_X2 U19055 ( .I(n17447), .ZN(n28212) );
  INV_X2 U19057 ( .I(n34479), .ZN(n33510) );
  INV_X1 U19059 ( .I(n2947), .ZN(n39203) );
  NOR2_X1 U19061 ( .A1(n495), .A2(n2947), .ZN(n459) );
  CLKBUF_X4 U19069 ( .I(n17833), .Z(n17792) );
  AOI21_X1 U19071 ( .A1(n32974), .A2(n25874), .B(n3575), .ZN(n36375) );
  NAND2_X1 U19072 ( .A1(n18866), .A2(n5258), .ZN(n7427) );
  INV_X2 U19073 ( .I(n5258), .ZN(n7426) );
  NAND2_X1 U19077 ( .A1(n30299), .A2(n15423), .ZN(n16213) );
  INV_X1 U19080 ( .I(n30299), .ZN(n23379) );
  NAND3_X2 U19086 ( .A1(n6195), .A2(n32545), .A3(n6192), .ZN(n38207) );
  INV_X2 U19098 ( .I(n16048), .ZN(n1039) );
  NAND2_X1 U19101 ( .A1(n30574), .A2(n16048), .ZN(n22987) );
  INV_X2 U19102 ( .I(n5211), .ZN(n9193) );
  AOI21_X2 U19104 ( .A1(n8238), .A2(n16575), .B(n34472), .ZN(n38208) );
  AOI21_X2 U19107 ( .A1(n2542), .A2(n25858), .B(n2541), .ZN(n38209) );
  AOI21_X1 U19108 ( .A1(n8238), .A2(n16575), .B(n34472), .ZN(n36842) );
  AOI21_X1 U19111 ( .A1(n38141), .A2(n29802), .B(n2792), .ZN(n5880) );
  INV_X1 U19113 ( .I(n4353), .ZN(n27318) );
  NAND2_X1 U19114 ( .A1(n4353), .A2(n13973), .ZN(n4345) );
  NAND3_X1 U19117 ( .A1(n35963), .A2(n31931), .A3(n39316), .ZN(n10841) );
  OAI22_X1 U19120 ( .A1(n12212), .A2(n35545), .B1(n10122), .B2(n31931), .ZN(
        n10078) );
  NAND2_X1 U19121 ( .A1(n35545), .A2(n31931), .ZN(n9350) );
  XNOR2_X1 U19126 ( .A1(n3292), .A2(n25065), .ZN(n38210) );
  INV_X2 U19133 ( .I(n8728), .ZN(n1388) );
  NAND2_X1 U19134 ( .A1(n8728), .A2(n29231), .ZN(n38944) );
  AOI21_X1 U19139 ( .A1(n35184), .A2(n7975), .B(n1480), .ZN(n2563) );
  CLKBUF_X12 U19140 ( .I(n20778), .Z(n9809) );
  INV_X2 U19141 ( .I(n10764), .ZN(n33815) );
  CLKBUF_X12 U19146 ( .I(n19930), .Z(n438) );
  NOR2_X1 U19149 ( .A1(n28546), .A2(n3944), .ZN(n17073) );
  INV_X2 U19150 ( .I(n3944), .ZN(n28643) );
  NAND2_X1 U19153 ( .A1(n28546), .A2(n3944), .ZN(n28647) );
  NOR2_X1 U19154 ( .A1(n9530), .A2(n25943), .ZN(n9529) );
  OAI21_X1 U19157 ( .A1(n22173), .A2(n5450), .B(n14833), .ZN(n14903) );
  NAND3_X1 U19161 ( .A1(n35901), .A2(n14064), .A3(n20128), .ZN(n17765) );
  NOR2_X1 U19165 ( .A1(n31433), .A2(n34279), .ZN(n35608) );
  NAND2_X1 U19168 ( .A1(n34279), .A2(n31433), .ZN(n39159) );
  OAI21_X2 U19175 ( .A1(n11735), .A2(n4463), .B(n4462), .ZN(n38212) );
  OAI21_X1 U19177 ( .A1(n7922), .A2(n5941), .B(n39417), .ZN(n36805) );
  NAND2_X2 U19178 ( .A1(n26648), .A2(n36953), .ZN(n38213) );
  NAND2_X2 U19182 ( .A1(n26641), .A2(n36911), .ZN(n36953) );
  INV_X2 U19183 ( .I(n939), .ZN(n920) );
  NAND2_X1 U19186 ( .A1(n9682), .A2(n4516), .ZN(n14985) );
  NAND2_X1 U19187 ( .A1(n39454), .A2(n4516), .ZN(n4511) );
  XOR2_X1 U19192 ( .A1(n36468), .A2(n14302), .Z(n38214) );
  INV_X1 U19194 ( .I(n25669), .ZN(n38963) );
  CLKBUF_X12 U19196 ( .I(n25669), .Z(n178) );
  XOR2_X1 U19197 ( .A1(n2215), .A2(n2214), .Z(n38215) );
  NAND3_X1 U19198 ( .A1(n999), .A2(n495), .A3(n27153), .ZN(n39707) );
  CLKBUF_X4 U19200 ( .I(n7654), .Z(n21804) );
  INV_X1 U19203 ( .I(n7654), .ZN(n21806) );
  INV_X1 U19204 ( .I(n28182), .ZN(n4457) );
  AND2_X1 U19206 ( .A1(n38199), .A2(n20960), .Z(n26752) );
  NOR2_X1 U19209 ( .A1(n27221), .A2(n5588), .ZN(n27224) );
  INV_X1 U19210 ( .I(n11569), .ZN(n25665) );
  OR3_X1 U19224 ( .A1(n17180), .A2(n25782), .A3(n8407), .Z(n25826) );
  NAND2_X1 U19225 ( .A1(n7096), .A2(n19326), .ZN(n27054) );
  INV_X1 U19233 ( .I(n19326), .ZN(n27343) );
  OAI21_X1 U19234 ( .A1(n27341), .A2(n27131), .B(n19326), .ZN(n4667) );
  INV_X1 U19237 ( .I(n6282), .ZN(n1104) );
  NAND2_X1 U19243 ( .A1(n32682), .A2(n36935), .ZN(n32681) );
  NOR2_X1 U19247 ( .A1(n11770), .A2(n2546), .ZN(n38218) );
  NOR2_X1 U19249 ( .A1(n11770), .A2(n2546), .ZN(n38219) );
  NOR2_X1 U19251 ( .A1(n11770), .A2(n2546), .ZN(n2443) );
  INV_X2 U19253 ( .I(n23472), .ZN(n23749) );
  AND2_X2 U19254 ( .A1(n39820), .A2(n14332), .Z(n25542) );
  CLKBUF_X12 U19255 ( .I(n5514), .Z(n31283) );
  INV_X1 U19261 ( .I(n5514), .ZN(n18816) );
  CLKBUF_X2 U19262 ( .I(n29678), .Z(n33128) );
  NOR2_X1 U19264 ( .A1(n36969), .A2(n33893), .ZN(n2922) );
  XOR2_X1 U19265 ( .A1(n1775), .A2(n16357), .Z(n38221) );
  NOR2_X1 U19268 ( .A1(n34008), .A2(n27985), .ZN(n28105) );
  NOR2_X1 U19269 ( .A1(n27484), .A2(n30758), .ZN(n31000) );
  NAND3_X1 U19277 ( .A1(n35115), .A2(n13753), .A3(n27484), .ZN(n4741) );
  INV_X1 U19278 ( .I(n25289), .ZN(n38511) );
  INV_X1 U19279 ( .I(n1234), .ZN(n26908) );
  NAND3_X2 U19280 ( .A1(n5344), .A2(n5342), .A3(n8048), .ZN(n38222) );
  XOR2_X1 U19281 ( .A1(n5731), .A2(n36339), .Z(n38223) );
  INV_X1 U19284 ( .I(n7990), .ZN(n7992) );
  XOR2_X1 U19293 ( .A1(n16696), .A2(n16698), .Z(n38224) );
  AOI21_X1 U19299 ( .A1(n27287), .A2(n1080), .B(n6010), .ZN(n38225) );
  AOI21_X1 U19300 ( .A1(n27287), .A2(n1080), .B(n6010), .ZN(n38226) );
  INV_X1 U19305 ( .I(n14869), .ZN(n38227) );
  NAND3_X2 U19306 ( .A1(n38516), .A2(n38525), .A3(n27242), .ZN(n38228) );
  NAND3_X2 U19307 ( .A1(n27238), .A2(n27237), .A3(n38690), .ZN(n38516) );
  NAND2_X1 U19309 ( .A1(n17685), .A2(n32675), .ZN(n21503) );
  NOR3_X1 U19311 ( .A1(n10242), .A2(n17685), .A3(n12077), .ZN(n12040) );
  CLKBUF_X12 U19312 ( .I(n29199), .Z(n30193) );
  INV_X1 U19319 ( .I(n29199), .ZN(n30229) );
  INV_X1 U19320 ( .I(n32043), .ZN(n12303) );
  AOI21_X1 U19322 ( .A1(n4008), .A2(n39098), .B(n5896), .ZN(n18326) );
  NOR2_X1 U19323 ( .A1(n35138), .A2(n692), .ZN(n2311) );
  AND2_X2 U19327 ( .A1(n22925), .A2(n18209), .Z(n22999) );
  INV_X1 U19336 ( .I(n35242), .ZN(n20041) );
  NOR2_X1 U19339 ( .A1(n1420), .A2(n38155), .ZN(n15963) );
  XOR2_X1 U19340 ( .A1(n38564), .A2(n3232), .Z(n38229) );
  INV_X1 U19341 ( .I(n8093), .ZN(n38230) );
  NOR2_X1 U19342 ( .A1(n28704), .A2(n38220), .ZN(n27897) );
  INV_X1 U19344 ( .I(n26558), .ZN(n35746) );
  NOR2_X1 U19350 ( .A1(n35254), .A2(n12198), .ZN(n30176) );
  INV_X1 U19351 ( .I(n28686), .ZN(n31045) );
  OAI21_X1 U19366 ( .A1(n1527), .A2(n38168), .B(n14375), .ZN(n3433) );
  INV_X2 U19368 ( .I(n5383), .ZN(n28608) );
  NAND2_X1 U19372 ( .A1(n5383), .A2(n36588), .ZN(n3637) );
  NAND2_X1 U19374 ( .A1(n7769), .A2(n10980), .ZN(n39076) );
  NOR2_X1 U19375 ( .A1(n16213), .A2(n23358), .ZN(n462) );
  NAND2_X1 U19378 ( .A1(n23379), .A2(n23358), .ZN(n23359) );
  NAND2_X1 U19379 ( .A1(n23358), .A2(n23250), .ZN(n31199) );
  NAND2_X2 U19381 ( .A1(n12660), .A2(n12661), .ZN(n10558) );
  NAND3_X2 U19384 ( .A1(n22048), .A2(n37199), .A3(n19089), .ZN(n12660) );
  INV_X2 U19386 ( .I(n38235), .ZN(n11363) );
  NOR2_X2 U19387 ( .A1(n25539), .A2(n39820), .ZN(n38235) );
  INV_X1 U19388 ( .I(n14282), .ZN(n38237) );
  INV_X2 U19389 ( .I(n38239), .ZN(n39810) );
  XOR2_X1 U19390 ( .A1(n7199), .A2(n7201), .Z(n38239) );
  XOR2_X1 U19391 ( .A1(n25172), .A2(n18428), .Z(n11369) );
  XOR2_X1 U19393 ( .A1(n26261), .A2(n31537), .Z(n9762) );
  XOR2_X1 U19398 ( .A1(n14353), .A2(n23710), .Z(n23887) );
  XOR2_X1 U19403 ( .A1(n35070), .A2(n38179), .Z(n17119) );
  NOR2_X1 U19405 ( .A1(n16948), .A2(n16949), .ZN(n17936) );
  XOR2_X1 U19406 ( .A1(n23666), .A2(n38240), .Z(n36272) );
  XOR2_X1 U19413 ( .A1(n23729), .A2(n12799), .Z(n38240) );
  AOI21_X1 U19414 ( .A1(n6581), .A2(n37589), .B(n14561), .ZN(n13206) );
  OAI21_X2 U19415 ( .A1(n11598), .A2(n21439), .B(n6690), .ZN(n33738) );
  AOI22_X2 U19416 ( .A1(n693), .A2(n21692), .B1(n21339), .B2(n21687), .ZN(
        n21439) );
  NAND2_X2 U19419 ( .A1(n21993), .A2(n21992), .ZN(n17310) );
  BUF_X2 U19422 ( .I(n39639), .Z(n38241) );
  OR2_X2 U19425 ( .A1(n18998), .A2(n8071), .Z(n22272) );
  AOI22_X1 U19427 ( .A1(n29599), .A2(n31667), .B1(n4786), .B2(n38420), .ZN(
        n33746) );
  XOR2_X1 U19430 ( .A1(n1618), .A2(n23686), .Z(n24033) );
  NAND2_X2 U19432 ( .A1(n34662), .A2(n37395), .ZN(n38242) );
  NOR2_X2 U19434 ( .A1(n38390), .A2(n7491), .ZN(n16013) );
  XOR2_X1 U19440 ( .A1(n36057), .A2(n38243), .Z(n14110) );
  XOR2_X1 U19442 ( .A1(n22454), .A2(n22766), .Z(n38243) );
  NAND2_X2 U19448 ( .A1(n38508), .A2(n35697), .ZN(n3015) );
  AND2_X1 U19451 ( .A1(n8604), .A2(n8395), .Z(n18628) );
  XOR2_X1 U19454 ( .A1(n5322), .A2(n6516), .Z(n24195) );
  BUF_X2 U19455 ( .I(n18425), .Z(n38248) );
  NAND2_X2 U19459 ( .A1(n22843), .A2(n2163), .ZN(n38249) );
  OAI21_X2 U19469 ( .A1(n13121), .A2(n19218), .B(n18162), .ZN(n32897) );
  XOR2_X1 U19473 ( .A1(n792), .A2(n3824), .Z(n3823) );
  XNOR2_X1 U19476 ( .A1(n3503), .A2(n18175), .ZN(n3824) );
  XOR2_X1 U19477 ( .A1(n14113), .A2(n38253), .Z(n7674) );
  XOR2_X1 U19478 ( .A1(n22603), .A2(n14112), .Z(n38253) );
  XOR2_X1 U19482 ( .A1(n27530), .A2(n38254), .Z(n27875) );
  XOR2_X1 U19483 ( .A1(n27527), .A2(n39465), .Z(n38254) );
  XOR2_X1 U19484 ( .A1(n18175), .A2(n32122), .Z(n23863) );
  AND2_X1 U19487 ( .A1(n740), .A2(n8556), .Z(n8652) );
  NAND2_X2 U19494 ( .A1(n36623), .A2(n5028), .ZN(n28730) );
  NAND2_X2 U19499 ( .A1(n31042), .A2(n38923), .ZN(n36623) );
  XOR2_X1 U19508 ( .A1(n4440), .A2(n16199), .Z(n4438) );
  XOR2_X1 U19511 ( .A1(n15346), .A2(n16226), .Z(n16199) );
  NAND2_X2 U19514 ( .A1(n39262), .A2(n27064), .ZN(n8372) );
  AND2_X1 U19517 ( .A1(n9118), .A2(n735), .Z(n6501) );
  XOR2_X1 U19519 ( .A1(n13369), .A2(n13367), .Z(n18156) );
  XOR2_X1 U19522 ( .A1(n8408), .A2(n8410), .Z(n32806) );
  OR2_X1 U19524 ( .A1(n38255), .A2(n30198), .Z(n2767) );
  NOR2_X2 U19525 ( .A1(n33861), .A2(n1755), .ZN(n30198) );
  INV_X1 U19528 ( .I(n29222), .ZN(n29224) );
  NAND2_X1 U19530 ( .A1(n29222), .A2(n6002), .ZN(n3415) );
  NOR2_X2 U19532 ( .A1(n38257), .A2(n38256), .ZN(n29222) );
  INV_X1 U19534 ( .I(n36694), .ZN(n38256) );
  OAI21_X1 U19541 ( .A1(n18278), .A2(n18039), .B(n38258), .ZN(n36862) );
  NAND2_X1 U19543 ( .A1(n29205), .A2(n18039), .ZN(n38258) );
  NAND2_X2 U19544 ( .A1(n10595), .A2(n34897), .ZN(n19326) );
  XOR2_X1 U19548 ( .A1(n26429), .A2(n12300), .Z(n12299) );
  XOR2_X1 U19549 ( .A1(n33027), .A2(n38619), .Z(n26429) );
  OAI21_X2 U19550 ( .A1(n11886), .A2(n29201), .B(n34983), .ZN(n29204) );
  NAND2_X2 U19551 ( .A1(n7745), .A2(n3945), .ZN(n3944) );
  XOR2_X1 U19553 ( .A1(n34491), .A2(n11814), .Z(n16500) );
  NOR2_X2 U19557 ( .A1(n7872), .A2(n28215), .ZN(n38443) );
  INV_X2 U19567 ( .I(n38259), .ZN(n20860) );
  OAI21_X1 U19569 ( .A1(n16577), .A2(n17708), .B(n38260), .ZN(n5778) );
  AOI22_X1 U19575 ( .A1(n5779), .A2(n20498), .B1(n29717), .B2(n29722), .ZN(
        n38260) );
  XOR2_X1 U19576 ( .A1(n22668), .A2(n38261), .Z(n649) );
  NAND2_X2 U19586 ( .A1(n17901), .A2(n17902), .ZN(n35241) );
  NOR2_X2 U19594 ( .A1(n14626), .A2(n16953), .ZN(n17901) );
  OAI21_X2 U19596 ( .A1(n8105), .A2(n26726), .B(n26725), .ZN(n27269) );
  XOR2_X1 U19599 ( .A1(n2005), .A2(n2002), .Z(n9649) );
  BUF_X2 U19601 ( .I(n20018), .Z(n38262) );
  XOR2_X1 U19603 ( .A1(n24017), .A2(n24016), .Z(n14719) );
  XOR2_X1 U19605 ( .A1(n24026), .A2(n38263), .Z(n39591) );
  XOR2_X1 U19607 ( .A1(n10722), .A2(n11180), .Z(n38263) );
  AOI21_X2 U19608 ( .A1(n36287), .A2(n34570), .B(n27103), .ZN(n27802) );
  NOR2_X1 U19610 ( .A1(n9489), .A2(n9487), .ZN(n5458) );
  XOR2_X1 U19612 ( .A1(n38264), .A2(n18316), .Z(n18315) );
  XOR2_X1 U19616 ( .A1(n18319), .A2(n30925), .Z(n38264) );
  XOR2_X1 U19617 ( .A1(n1262), .A2(n25086), .Z(n8240) );
  OAI22_X2 U19629 ( .A1(n14538), .A2(n15826), .B1(n20119), .B2(n1608), .ZN(
        n32637) );
  XOR2_X1 U19634 ( .A1(n27640), .A2(n38265), .Z(n39742) );
  INV_X1 U19638 ( .I(n29920), .ZN(n38265) );
  NAND2_X2 U19639 ( .A1(n14586), .A2(n38873), .ZN(n27640) );
  NAND2_X1 U19647 ( .A1(n19420), .A2(n8966), .ZN(n24500) );
  NOR2_X2 U19652 ( .A1(n38835), .A2(n32690), .ZN(n30696) );
  NAND2_X2 U19653 ( .A1(n9173), .A2(n35673), .ZN(n35187) );
  XOR2_X1 U19654 ( .A1(n23736), .A2(n23913), .Z(n12921) );
  XOR2_X1 U19659 ( .A1(n38267), .A2(n27465), .Z(Ciphertext[185]) );
  NAND2_X1 U19665 ( .A1(n27456), .A2(n37158), .ZN(n26641) );
  XOR2_X1 U19668 ( .A1(n26257), .A2(n13131), .Z(n17063) );
  XOR2_X1 U19676 ( .A1(n26381), .A2(n9870), .Z(n13131) );
  NAND2_X2 U19678 ( .A1(n2316), .A2(n25755), .ZN(n35138) );
  BUF_X2 U19679 ( .I(n32095), .Z(n38269) );
  NAND2_X2 U19681 ( .A1(n28256), .A2(n3989), .ZN(n28047) );
  XNOR2_X1 U19683 ( .A1(n10520), .A2(n6185), .ZN(n25222) );
  NAND2_X2 U19684 ( .A1(n38296), .A2(n38270), .ZN(n25813) );
  AOI22_X2 U19687 ( .A1(n12404), .A2(n1117), .B1(n19863), .B2(n25660), .ZN(
        n38270) );
  OAI21_X2 U19688 ( .A1(n37123), .A2(n9064), .B(n9063), .ZN(n29794) );
  XOR2_X1 U19689 ( .A1(n38271), .A2(n38969), .Z(n27919) );
  XOR2_X1 U19692 ( .A1(n33883), .A2(n27788), .Z(n38271) );
  NAND2_X2 U19698 ( .A1(n959), .A2(n626), .ZN(n33586) );
  NAND2_X2 U19699 ( .A1(n6054), .A2(n6053), .ZN(n23775) );
  AOI22_X2 U19700 ( .A1(n38274), .A2(n38272), .B1(n21527), .B2(n39627), .ZN(
        n39616) );
  NOR2_X2 U19701 ( .A1(n39627), .A2(n38273), .ZN(n38272) );
  INV_X2 U19704 ( .I(n35071), .ZN(n38274) );
  XOR2_X1 U19706 ( .A1(n29071), .A2(n28886), .Z(n28914) );
  NAND3_X2 U19710 ( .A1(n35415), .A2(n35414), .A3(n16632), .ZN(n11831) );
  XOR2_X1 U19712 ( .A1(n8183), .A2(n25252), .Z(n21253) );
  NAND2_X2 U19715 ( .A1(n12676), .A2(n35688), .ZN(n8183) );
  NAND2_X2 U19717 ( .A1(n4990), .A2(n30595), .ZN(n32748) );
  XOR2_X1 U19718 ( .A1(n35218), .A2(n8302), .Z(n36637) );
  NOR2_X2 U19719 ( .A1(n1333), .A2(n3003), .ZN(n22230) );
  INV_X2 U19722 ( .I(n31271), .ZN(n38839) );
  XOR2_X1 U19724 ( .A1(n5179), .A2(n36540), .Z(n31271) );
  NAND2_X2 U19725 ( .A1(n10128), .A2(n10126), .ZN(n38395) );
  XOR2_X1 U19728 ( .A1(n28971), .A2(n13639), .Z(n29123) );
  NAND2_X2 U19729 ( .A1(n28648), .A2(n18891), .ZN(n13639) );
  NAND2_X2 U19730 ( .A1(n34579), .A2(n38276), .ZN(n27023) );
  XOR2_X1 U19742 ( .A1(n6317), .A2(n6196), .Z(n20727) );
  NAND2_X2 U19743 ( .A1(n28416), .A2(n28417), .ZN(n6196) );
  NOR2_X2 U19744 ( .A1(n34685), .A2(n34350), .ZN(n25737) );
  XOR2_X1 U19745 ( .A1(n27807), .A2(n20846), .Z(n32647) );
  XOR2_X1 U19746 ( .A1(n33197), .A2(n25252), .Z(n25302) );
  NAND2_X1 U19753 ( .A1(n4516), .A2(n6904), .ZN(n12569) );
  NAND2_X2 U19757 ( .A1(n9540), .A2(n25559), .ZN(n4516) );
  NAND2_X2 U19759 ( .A1(n5675), .A2(n27274), .ZN(n27085) );
  NAND3_X2 U19760 ( .A1(n38277), .A2(n27151), .A3(n27148), .ZN(n27778) );
  AOI22_X2 U19761 ( .A1(n33910), .A2(n38278), .B1(n28401), .B2(n11490), .ZN(
        n11492) );
  NAND2_X2 U19765 ( .A1(n2937), .A2(n12537), .ZN(n38278) );
  AOI21_X2 U19767 ( .A1(n11591), .A2(n943), .B(n11590), .ZN(n13245) );
  INV_X2 U19768 ( .I(n38280), .ZN(n37054) );
  XOR2_X1 U19779 ( .A1(n3459), .A2(n3456), .Z(n38280) );
  NOR3_X1 U19782 ( .A1(n1429), .A2(n10907), .A3(n18871), .ZN(n32075) );
  XOR2_X1 U19783 ( .A1(n29050), .A2(n29125), .Z(n29158) );
  XOR2_X1 U19786 ( .A1(n38605), .A2(n21271), .Z(n36396) );
  XOR2_X1 U19791 ( .A1(n30502), .A2(n38890), .Z(n38781) );
  OAI22_X2 U19795 ( .A1(n924), .A2(n3388), .B1(n38214), .B2(n14458), .ZN(n8686) );
  OAI21_X2 U19806 ( .A1(n35295), .A2(n35296), .B(n32714), .ZN(n29438) );
  XOR2_X1 U19808 ( .A1(n22657), .A2(n22761), .Z(n22608) );
  NAND2_X2 U19816 ( .A1(n16548), .A2(n30212), .ZN(n38829) );
  NAND3_X2 U19819 ( .A1(n17648), .A2(n32598), .A3(n2632), .ZN(n39481) );
  NAND2_X2 U19823 ( .A1(n2633), .A2(n1633), .ZN(n17648) );
  NAND2_X2 U19825 ( .A1(n39503), .A2(n38281), .ZN(n27683) );
  AOI22_X1 U19826 ( .A1(n27017), .A2(n39424), .B1(n27224), .B2(n13278), .ZN(
        n38281) );
  NOR2_X2 U19827 ( .A1(n38283), .A2(n38282), .ZN(n22803) );
  INV_X1 U19828 ( .I(n14752), .ZN(n38284) );
  BUF_X2 U19829 ( .I(n24712), .Z(n38285) );
  AND2_X1 U19830 ( .A1(n20541), .A2(n33963), .Z(n38919) );
  NAND2_X2 U19831 ( .A1(n38286), .A2(n38354), .ZN(n16526) );
  XOR2_X1 U19835 ( .A1(n16552), .A2(n16554), .Z(n32750) );
  AOI21_X2 U19841 ( .A1(n37141), .A2(n32084), .B(n34643), .ZN(n16636) );
  NAND2_X2 U19848 ( .A1(n30311), .A2(n94), .ZN(n33944) );
  XOR2_X1 U19857 ( .A1(n6571), .A2(n11105), .Z(n26490) );
  NAND2_X2 U19858 ( .A1(n32380), .A2(n39777), .ZN(n11105) );
  XOR2_X1 U19861 ( .A1(n26567), .A2(n26334), .Z(n35721) );
  NAND2_X2 U19868 ( .A1(n9377), .A2(n31883), .ZN(n26567) );
  NOR2_X2 U19871 ( .A1(n33289), .A2(n35954), .ZN(n24219) );
  NOR2_X2 U19872 ( .A1(n22019), .A2(n2818), .ZN(n38287) );
  NAND2_X2 U19877 ( .A1(n38391), .A2(n38288), .ZN(n11120) );
  XOR2_X1 U19880 ( .A1(n38289), .A2(n1160), .Z(Ciphertext[22]) );
  NOR2_X1 U19887 ( .A1(n38348), .A2(n30577), .ZN(n38289) );
  NAND2_X2 U19889 ( .A1(n35158), .A2(n17420), .ZN(n27779) );
  OAI21_X2 U19891 ( .A1(n25838), .A2(n38982), .B(n25837), .ZN(n9989) );
  XOR2_X1 U19900 ( .A1(n33010), .A2(n38291), .Z(n23921) );
  INV_X2 U19904 ( .I(n24049), .ZN(n38291) );
  BUF_X2 U19906 ( .I(n388), .Z(n38292) );
  XOR2_X1 U19907 ( .A1(n38294), .A2(n20400), .Z(n18188) );
  XOR2_X1 U19909 ( .A1(n36628), .A2(n27648), .Z(n38294) );
  NAND2_X2 U19910 ( .A1(n35750), .A2(n34644), .ZN(n10032) );
  AOI22_X2 U19911 ( .A1(n18484), .A2(n2396), .B1(n24331), .B2(n24330), .ZN(
        n34263) );
  NOR2_X2 U19915 ( .A1(n12733), .A2(n24328), .ZN(n18484) );
  XOR2_X1 U19916 ( .A1(n38958), .A2(n38192), .Z(n38809) );
  NAND2_X2 U19917 ( .A1(n38847), .A2(n8406), .ZN(n7990) );
  XOR2_X1 U19918 ( .A1(n38295), .A2(n2351), .Z(n23202) );
  XOR2_X1 U19921 ( .A1(n14297), .A2(n2354), .Z(n38295) );
  OAI21_X2 U19924 ( .A1(n34099), .A2(n229), .B(n25662), .ZN(n38296) );
  XOR2_X1 U19925 ( .A1(n29039), .A2(n28920), .Z(n8678) );
  XOR2_X1 U19926 ( .A1(n9106), .A2(n12989), .Z(n28920) );
  XOR2_X1 U19927 ( .A1(n24019), .A2(n23676), .Z(n5255) );
  NAND2_X2 U19930 ( .A1(n38298), .A2(n38297), .ZN(n20255) );
  AOI22_X1 U19931 ( .A1(n32372), .A2(n12144), .B1(n17233), .B2(n14418), .ZN(
        n38297) );
  OAI21_X2 U19933 ( .A1(n21535), .A2(n21536), .B(n14501), .ZN(n38298) );
  XNOR2_X1 U19941 ( .A1(n26391), .A2(n19450), .ZN(n26449) );
  NAND3_X2 U19943 ( .A1(n38301), .A2(n37182), .A3(n9427), .ZN(n18994) );
  NAND2_X2 U19944 ( .A1(n28429), .A2(n12797), .ZN(n8729) );
  OAI21_X1 U19946 ( .A1(n37126), .A2(n4347), .B(n38308), .ZN(n8328) );
  XOR2_X1 U19948 ( .A1(n16109), .A2(n16110), .Z(n15865) );
  NAND2_X1 U19949 ( .A1(n22206), .A2(n19837), .ZN(n38932) );
  NAND2_X1 U19953 ( .A1(n38932), .A2(n38931), .ZN(n22211) );
  NOR2_X2 U19959 ( .A1(n12063), .A2(n6150), .ZN(n26334) );
  XOR2_X1 U19964 ( .A1(n23868), .A2(n675), .Z(n20485) );
  XOR2_X1 U19968 ( .A1(n36842), .A2(n19656), .Z(n23868) );
  NAND2_X2 U19972 ( .A1(n18170), .A2(n18171), .ZN(n20589) );
  XOR2_X1 U19973 ( .A1(n12215), .A2(n38309), .Z(n21116) );
  XOR2_X1 U19977 ( .A1(n31582), .A2(n28986), .Z(n38309) );
  OAI22_X2 U19978 ( .A1(n13427), .A2(n33849), .B1(n26811), .B2(n26810), .ZN(
        n12756) );
  INV_X2 U19985 ( .I(n38310), .ZN(n13427) );
  NOR2_X2 U19996 ( .A1(n12755), .A2(n13770), .ZN(n38310) );
  NAND2_X2 U19997 ( .A1(n17583), .A2(n5424), .ZN(n8423) );
  AND2_X1 U20002 ( .A1(n10940), .A2(n24408), .Z(n39271) );
  INV_X2 U20003 ( .I(n10520), .ZN(n25256) );
  NAND2_X2 U20004 ( .A1(n35664), .A2(n19559), .ZN(n23302) );
  INV_X1 U20009 ( .I(n2283), .ZN(n27520) );
  OR2_X1 U20023 ( .A1(n36371), .A2(n3644), .Z(n17998) );
  XOR2_X1 U20028 ( .A1(n18423), .A2(n18421), .Z(n34956) );
  NAND3_X2 U20029 ( .A1(n38312), .A2(n39324), .A3(n39325), .ZN(n35813) );
  XOR2_X1 U20031 ( .A1(n12520), .A2(n36389), .Z(n38486) );
  XNOR2_X1 U20033 ( .A1(n10683), .A2(n10684), .ZN(n38465) );
  NOR3_X2 U20034 ( .A1(n37108), .A2(n39303), .A3(n39752), .ZN(n35950) );
  XOR2_X1 U20035 ( .A1(n39804), .A2(n17310), .Z(n18239) );
  XOR2_X1 U20040 ( .A1(n26229), .A2(n38313), .Z(n38842) );
  XOR2_X1 U20041 ( .A1(n11298), .A2(n26525), .Z(n38313) );
  XOR2_X1 U20042 ( .A1(n38314), .A2(n20748), .Z(Ciphertext[165]) );
  NOR4_X2 U20046 ( .A1(n34706), .A2(n34707), .A3(n35625), .A4(n35624), .ZN(
        n38314) );
  NAND2_X2 U20049 ( .A1(n36099), .A2(n26113), .ZN(n39066) );
  NAND3_X2 U20050 ( .A1(n36678), .A2(n31004), .A3(n371), .ZN(n35665) );
  NAND2_X1 U20054 ( .A1(n1948), .A2(n15427), .ZN(n16146) );
  XOR2_X1 U20055 ( .A1(n38316), .A2(n38315), .Z(n31485) );
  XOR2_X1 U20057 ( .A1(n17189), .A2(n31576), .Z(n38315) );
  XOR2_X1 U20061 ( .A1(n1323), .A2(n31504), .Z(n38316) );
  AND2_X1 U20062 ( .A1(n5768), .A2(n38317), .Z(n12680) );
  XOR2_X1 U20063 ( .A1(n3976), .A2(n3975), .Z(n38742) );
  INV_X1 U20064 ( .I(n19783), .ZN(n38319) );
  INV_X1 U20066 ( .I(n14789), .ZN(n38320) );
  NAND3_X1 U20068 ( .A1(n11453), .A2(n38656), .A3(n19068), .ZN(n12746) );
  XOR2_X1 U20069 ( .A1(n38321), .A2(n23985), .Z(n23991) );
  XOR2_X1 U20070 ( .A1(n23984), .A2(n35235), .Z(n38321) );
  NAND2_X1 U20073 ( .A1(n3593), .A2(n38960), .ZN(n39016) );
  XOR2_X1 U20075 ( .A1(n38322), .A2(n11570), .Z(n32994) );
  XOR2_X1 U20077 ( .A1(n33924), .A2(n25197), .Z(n38322) );
  OAI22_X1 U20078 ( .A1(n21983), .A2(n3907), .B1(n3644), .B2(n38323), .ZN(
        n11440) );
  OR2_X1 U20080 ( .A1(n3907), .A2(n21982), .Z(n38323) );
  XOR2_X1 U20081 ( .A1(n38324), .A2(n19648), .Z(Ciphertext[99]) );
  NAND2_X1 U20085 ( .A1(n29736), .A2(n19369), .ZN(n38324) );
  XOR2_X1 U20086 ( .A1(n24074), .A2(n20973), .Z(n20550) );
  XOR2_X1 U20089 ( .A1(n23898), .A2(n23955), .Z(n24074) );
  NAND2_X2 U20092 ( .A1(n33161), .A2(n13755), .ZN(n38669) );
  XOR2_X1 U20093 ( .A1(n25234), .A2(n14214), .Z(n12997) );
  XOR2_X1 U20096 ( .A1(n38325), .A2(n19534), .Z(Ciphertext[113]) );
  NAND2_X1 U20098 ( .A1(n6441), .A2(n6438), .ZN(n38325) );
  XOR2_X1 U20099 ( .A1(n18335), .A2(n38326), .Z(n850) );
  XOR2_X1 U20105 ( .A1(n35202), .A2(n33735), .Z(n38326) );
  XOR2_X1 U20107 ( .A1(n29041), .A2(n31547), .Z(n28873) );
  OAI21_X2 U20116 ( .A1(n2335), .A2(n2334), .B(n33649), .ZN(n31547) );
  NAND2_X2 U20117 ( .A1(n31027), .A2(n30668), .ZN(n5424) );
  XOR2_X1 U20120 ( .A1(n18813), .A2(n7070), .Z(n39516) );
  BUF_X2 U20126 ( .I(n16123), .Z(n38328) );
  AND2_X1 U20132 ( .A1(n5514), .A2(n39011), .Z(n39110) );
  NAND3_X1 U20134 ( .A1(n24532), .A2(n6169), .A3(n957), .ZN(n38331) );
  NAND2_X2 U20135 ( .A1(n7487), .A2(n38332), .ZN(n24002) );
  AOI22_X2 U20136 ( .A1(n30460), .A2(n1644), .B1(n33080), .B2(n605), .ZN(
        n38332) );
  NAND2_X2 U20140 ( .A1(n27116), .A2(n7588), .ZN(n38333) );
  OR2_X1 U20150 ( .A1(n18619), .A2(n19949), .Z(n17586) );
  XOR2_X1 U20151 ( .A1(n26539), .A2(n26513), .Z(n5225) );
  XOR2_X1 U20155 ( .A1(n38619), .A2(n26161), .Z(n26513) );
  XNOR2_X1 U20159 ( .A1(n22551), .A2(n5463), .ZN(n39040) );
  XOR2_X1 U20164 ( .A1(n22586), .A2(n20392), .Z(n5463) );
  NOR2_X2 U20166 ( .A1(n14746), .A2(n20788), .ZN(n38334) );
  XOR2_X1 U20167 ( .A1(n25079), .A2(n38336), .Z(n39563) );
  NAND2_X2 U20168 ( .A1(n6574), .A2(n6837), .ZN(n25079) );
  NOR2_X1 U20169 ( .A1(n20739), .A2(n32043), .ZN(n28324) );
  INV_X1 U20179 ( .I(n39140), .ZN(n34524) );
  OAI21_X2 U20188 ( .A1(n36433), .A2(n36434), .B(n38642), .ZN(n39140) );
  AND3_X1 U20198 ( .A1(n3988), .A2(n28616), .A3(n6287), .Z(n5385) );
  AOI22_X2 U20201 ( .A1(n37181), .A2(n38338), .B1(n25627), .B2(n37748), .ZN(
        n31082) );
  NOR2_X2 U20204 ( .A1(n11476), .A2(n2272), .ZN(n38400) );
  AOI22_X2 U20207 ( .A1(n16206), .A2(n35326), .B1(n4871), .B2(n28548), .ZN(
        n35262) );
  NAND2_X2 U20212 ( .A1(n32651), .A2(n32637), .ZN(n16579) );
  NOR2_X1 U20215 ( .A1(n10913), .A2(n26978), .ZN(n34868) );
  NOR2_X2 U20223 ( .A1(n852), .A2(n17097), .ZN(n10913) );
  XOR2_X1 U20228 ( .A1(n39215), .A2(n10525), .Z(n34616) );
  NAND2_X2 U20230 ( .A1(n21245), .A2(n10472), .ZN(n19559) );
  INV_X2 U20240 ( .I(n19671), .ZN(n1299) );
  NAND2_X2 U20243 ( .A1(n13087), .A2(n39819), .ZN(n19671) );
  NAND2_X2 U20244 ( .A1(n4010), .A2(n10729), .ZN(n4301) );
  OAI22_X2 U20245 ( .A1(n7107), .A2(n33359), .B1(n7108), .B2(n38339), .ZN(
        n22659) );
  NAND2_X2 U20247 ( .A1(n38663), .A2(n39782), .ZN(n7512) );
  XOR2_X1 U20248 ( .A1(n10647), .A2(n4734), .Z(n11062) );
  NAND2_X2 U20249 ( .A1(n10646), .A2(n10645), .ZN(n10647) );
  NOR2_X2 U20253 ( .A1(n23072), .A2(n22919), .ZN(n36230) );
  NAND2_X2 U20255 ( .A1(n38634), .A2(n2850), .ZN(n17653) );
  NAND2_X2 U20262 ( .A1(n38340), .A2(n16763), .ZN(n21543) );
  XOR2_X1 U20264 ( .A1(n16627), .A2(n1558), .Z(n11570) );
  INV_X2 U20265 ( .I(n38341), .ZN(n21117) );
  NOR2_X2 U20267 ( .A1(n2654), .A2(n21982), .ZN(n38341) );
  NAND2_X2 U20268 ( .A1(n38342), .A2(n2941), .ZN(n18012) );
  XOR2_X1 U20278 ( .A1(n29029), .A2(n29030), .Z(n9768) );
  XOR2_X1 U20279 ( .A1(n15780), .A2(n29818), .Z(n29030) );
  XOR2_X1 U20296 ( .A1(n38343), .A2(n23876), .Z(n1923) );
  XOR2_X1 U20298 ( .A1(n13224), .A2(n36143), .Z(n38343) );
  XOR2_X1 U20300 ( .A1(n12014), .A2(n3150), .Z(n38344) );
  AND2_X2 U20303 ( .A1(n34134), .A2(n11657), .Z(n25364) );
  XOR2_X1 U20304 ( .A1(n17567), .A2(n35320), .Z(n21108) );
  NAND2_X2 U20305 ( .A1(n38469), .A2(n8320), .ZN(n17567) );
  XOR2_X1 U20306 ( .A1(n15517), .A2(n15516), .Z(n19928) );
  NAND2_X2 U20308 ( .A1(n8314), .A2(n1579), .ZN(n8317) );
  OAI21_X2 U20311 ( .A1(n28727), .A2(n8094), .B(n34525), .ZN(n8090) );
  INV_X2 U20316 ( .I(n39227), .ZN(n28727) );
  NAND3_X2 U20318 ( .A1(n27868), .A2(n27867), .A3(n18149), .ZN(n39227) );
  OAI21_X2 U20319 ( .A1(n1074), .A2(n12406), .B(n1200), .ZN(n38345) );
  NAND3_X2 U20320 ( .A1(n31695), .A2(n24957), .A3(n38346), .ZN(n26092) );
  NAND3_X1 U20321 ( .A1(n38338), .A2(n25756), .A3(n12675), .ZN(n38346) );
  INV_X2 U20324 ( .I(n26432), .ZN(n12934) );
  NOR2_X1 U20325 ( .A1(n20889), .A2(n35399), .ZN(n14777) );
  NAND2_X2 U20326 ( .A1(n21774), .A2(n21773), .ZN(n20889) );
  NAND2_X1 U20328 ( .A1(n25261), .A2(n11727), .ZN(n34411) );
  NAND2_X1 U20331 ( .A1(n11394), .A2(n11395), .ZN(n38348) );
  NAND2_X1 U20335 ( .A1(n38686), .A2(n33495), .ZN(n12704) );
  XOR2_X1 U20339 ( .A1(n23970), .A2(n23967), .Z(n23869) );
  NAND2_X2 U20340 ( .A1(n23301), .A2(n31052), .ZN(n23967) );
  OR2_X1 U20349 ( .A1(n33980), .A2(n28250), .Z(n28247) );
  XOR2_X1 U20351 ( .A1(n15995), .A2(n15994), .Z(n33980) );
  XOR2_X1 U20353 ( .A1(n23764), .A2(n38350), .Z(n37044) );
  INV_X2 U20359 ( .I(n23654), .ZN(n38350) );
  XOR2_X1 U20360 ( .A1(n38351), .A2(n6531), .Z(n6528) );
  XOR2_X1 U20361 ( .A1(n1620), .A2(n5699), .Z(n38351) );
  XOR2_X1 U20362 ( .A1(n29819), .A2(n29506), .Z(n38352) );
  OAI21_X2 U20364 ( .A1(n39034), .A2(n22863), .B(n9472), .ZN(n6213) );
  AND2_X2 U20366 ( .A1(n3839), .A2(n7696), .Z(n21461) );
  NAND2_X2 U20368 ( .A1(n16123), .A2(n14940), .ZN(n7207) );
  NOR2_X2 U20369 ( .A1(n961), .A2(n23401), .ZN(n38353) );
  OAI21_X2 U20371 ( .A1(n6744), .A2(n2898), .B(n37212), .ZN(n38354) );
  OAI21_X2 U20372 ( .A1(n3981), .A2(n9688), .B(n37006), .ZN(n2147) );
  XOR2_X1 U20374 ( .A1(n3652), .A2(n3650), .Z(n33446) );
  XOR2_X1 U20381 ( .A1(n9469), .A2(n9468), .Z(n39155) );
  OAI21_X2 U20382 ( .A1(n32937), .A2(n12146), .B(n38355), .ZN(n17806) );
  AOI21_X2 U20384 ( .A1(n36556), .A2(n19070), .B(n17810), .ZN(n38355) );
  NAND2_X1 U20386 ( .A1(n1211), .A2(n5402), .ZN(n6119) );
  NOR2_X2 U20388 ( .A1(n32325), .A2(n38356), .ZN(n18320) );
  NOR2_X2 U20394 ( .A1(n38359), .A2(n38358), .ZN(n38357) );
  INV_X2 U20395 ( .I(n25379), .ZN(n38358) );
  INV_X2 U20397 ( .I(n10674), .ZN(n38359) );
  XOR2_X1 U20400 ( .A1(n38361), .A2(n38360), .Z(n13759) );
  XOR2_X1 U20404 ( .A1(n26539), .A2(n15508), .Z(n38360) );
  XOR2_X1 U20406 ( .A1(n39743), .A2(n26419), .Z(n38361) );
  NAND2_X2 U20409 ( .A1(n14618), .A2(n19852), .ZN(n12227) );
  OR2_X2 U20419 ( .A1(n25355), .A2(n24896), .Z(n25389) );
  OAI22_X2 U20420 ( .A1(n3962), .A2(n37103), .B1(n3135), .B2(n1090), .ZN(
        n38435) );
  XOR2_X1 U20421 ( .A1(n6658), .A2(n31724), .Z(n32622) );
  INV_X2 U20424 ( .I(n5637), .ZN(n12231) );
  XOR2_X1 U20425 ( .A1(n28791), .A2(n6317), .Z(n5637) );
  XOR2_X1 U20428 ( .A1(n10401), .A2(n23945), .Z(n10400) );
  NAND3_X1 U20430 ( .A1(n33795), .A2(n2888), .A3(n3575), .ZN(n38633) );
  XOR2_X1 U20435 ( .A1(n33961), .A2(n20465), .Z(n7936) );
  NAND3_X2 U20437 ( .A1(n28521), .A2(n12947), .A3(n28520), .ZN(n20465) );
  NAND2_X1 U20439 ( .A1(n5671), .A2(n28285), .ZN(n34516) );
  XOR2_X1 U20440 ( .A1(n29049), .A2(n16355), .Z(n4393) );
  XOR2_X1 U20442 ( .A1(n1775), .A2(n16357), .Z(n16355) );
  XOR2_X1 U20445 ( .A1(n19608), .A2(n35196), .Z(n3929) );
  XOR2_X1 U20446 ( .A1(n19513), .A2(n29034), .Z(n15216) );
  AOI22_X2 U20447 ( .A1(n16474), .A2(n37311), .B1(n18836), .B2(n16475), .ZN(
        n19513) );
  XOR2_X1 U20448 ( .A1(n25046), .A2(n14563), .Z(n5033) );
  AOI21_X2 U20449 ( .A1(n6696), .A2(n1873), .B(n38364), .ZN(n39622) );
  XNOR2_X1 U20455 ( .A1(n5208), .A2(n29538), .ZN(n39720) );
  INV_X2 U20456 ( .I(n15922), .ZN(n38365) );
  NAND2_X1 U20462 ( .A1(n38367), .A2(n32472), .ZN(n38366) );
  NOR2_X1 U20463 ( .A1(n10272), .A2(n30716), .ZN(n38368) );
  BUF_X2 U20464 ( .I(n933), .Z(n38369) );
  XOR2_X1 U20465 ( .A1(n38371), .A2(n1370), .Z(Ciphertext[176]) );
  OAI21_X2 U20470 ( .A1(n13113), .A2(n13112), .B(n1771), .ZN(n23767) );
  NAND2_X2 U20472 ( .A1(n35690), .A2(n14206), .ZN(n1771) );
  XOR2_X1 U20476 ( .A1(n8324), .A2(n38430), .Z(n4894) );
  OAI21_X2 U20478 ( .A1(n19707), .A2(n1372), .B(n38372), .ZN(n22234) );
  NAND2_X2 U20483 ( .A1(n1372), .A2(n21755), .ZN(n38372) );
  OAI21_X2 U20485 ( .A1(n37143), .A2(n27163), .B(n27164), .ZN(n16997) );
  NOR2_X2 U20486 ( .A1(n15391), .A2(n38374), .ZN(n39200) );
  INV_X2 U20492 ( .I(n32107), .ZN(n7955) );
  OAI22_X2 U20495 ( .A1(n21553), .A2(n9886), .B1(n7954), .B2(n21719), .ZN(
        n32107) );
  XNOR2_X1 U20499 ( .A1(n21217), .A2(n20048), .ZN(n38763) );
  NAND2_X1 U20500 ( .A1(n22804), .A2(n14409), .ZN(n32676) );
  OAI21_X2 U20504 ( .A1(n8239), .A2(n13752), .B(n38376), .ZN(n10208) );
  BUF_X2 U20508 ( .I(n32623), .Z(n38377) );
  XOR2_X1 U20514 ( .A1(n32190), .A2(n18807), .Z(n2526) );
  NAND2_X2 U20515 ( .A1(n26113), .A2(n3642), .ZN(n17269) );
  NAND2_X2 U20522 ( .A1(n38476), .A2(n18349), .ZN(n26113) );
  OAI22_X2 U20528 ( .A1(n35902), .A2(n30671), .B1(n26966), .B2(n36234), .ZN(
        n27825) );
  NAND3_X2 U20531 ( .A1(n16621), .A2(n16634), .A3(n38378), .ZN(n22744) );
  NAND2_X2 U20532 ( .A1(n22136), .A2(n14196), .ZN(n38378) );
  NOR2_X2 U20533 ( .A1(n13601), .A2(n30304), .ZN(n13598) );
  NAND3_X2 U20534 ( .A1(n13600), .A2(n13599), .A3(n27874), .ZN(n30304) );
  NOR2_X2 U20535 ( .A1(n17869), .A2(n15868), .ZN(n22275) );
  OAI22_X1 U20536 ( .A1(n7515), .A2(n1121), .B1(n16210), .B2(n14283), .ZN(
        n24780) );
  NAND3_X2 U20537 ( .A1(n34167), .A2(n36159), .A3(n12326), .ZN(n34535) );
  NAND2_X2 U20542 ( .A1(n445), .A2(n5253), .ZN(n39038) );
  XOR2_X1 U20544 ( .A1(n7276), .A2(n38379), .Z(n22879) );
  XOR2_X1 U20548 ( .A1(n22745), .A2(n7275), .Z(n38379) );
  XOR2_X1 U20550 ( .A1(n6768), .A2(n39408), .Z(n39008) );
  OR2_X1 U20553 ( .A1(n36191), .A2(n34962), .Z(n38380) );
  XOR2_X1 U20556 ( .A1(n7288), .A2(n20460), .Z(n9787) );
  NAND2_X1 U20558 ( .A1(n5149), .A2(n20986), .ZN(n39174) );
  INV_X2 U20560 ( .I(n38381), .ZN(n36838) );
  NAND2_X2 U20566 ( .A1(n38450), .A2(n34930), .ZN(n38837) );
  AOI21_X2 U20570 ( .A1(n37255), .A2(n32682), .B(n38382), .ZN(n38717) );
  NOR3_X2 U20571 ( .A1(n7251), .A2(n36935), .A3(n9686), .ZN(n38382) );
  NOR2_X2 U20572 ( .A1(n38877), .A2(n27403), .ZN(n34036) );
  AND2_X1 U20575 ( .A1(n7485), .A2(n23577), .Z(n38726) );
  XOR2_X1 U20582 ( .A1(n38383), .A2(n13514), .Z(n14758) );
  XOR2_X1 U20583 ( .A1(n22518), .A2(n22519), .Z(n38383) );
  XOR2_X1 U20584 ( .A1(n29099), .A2(n12796), .Z(n38384) );
  NAND2_X1 U20585 ( .A1(n38751), .A2(n33384), .ZN(n2062) );
  BUF_X4 U20588 ( .I(n33993), .Z(n38448) );
  NAND2_X2 U20589 ( .A1(n13494), .A2(n14768), .ZN(n25179) );
  OAI21_X1 U20594 ( .A1(n33128), .A2(n29676), .B(n18042), .ZN(n29679) );
  XOR2_X1 U20595 ( .A1(n24014), .A2(n38385), .Z(n13654) );
  NAND2_X2 U20596 ( .A1(n38386), .A2(n16813), .ZN(n26571) );
  NOR3_X2 U20602 ( .A1(n38405), .A2(n38404), .A3(n34133), .ZN(n38387) );
  NOR2_X1 U20603 ( .A1(n5570), .A2(n921), .ZN(n9249) );
  INV_X2 U20607 ( .I(n5638), .ZN(n5570) );
  XOR2_X1 U20611 ( .A1(n1914), .A2(n1911), .Z(n5638) );
  NAND2_X2 U20612 ( .A1(n38388), .A2(n23041), .ZN(n23764) );
  NOR2_X2 U20613 ( .A1(n32060), .A2(n4707), .ZN(n38388) );
  OAI21_X2 U20617 ( .A1(n38493), .A2(n38494), .B(n21191), .ZN(n13213) );
  NOR2_X2 U20619 ( .A1(n23595), .A2(n23504), .ZN(n38929) );
  NOR2_X2 U20620 ( .A1(n24589), .A2(n31679), .ZN(n24538) );
  NAND2_X2 U20628 ( .A1(n5712), .A2(n5713), .ZN(n24589) );
  XOR2_X1 U20633 ( .A1(n9036), .A2(n33509), .Z(n29087) );
  MUX2_X1 U20634 ( .I0(n27897), .I1(n32002), .S(n31664), .Z(n27898) );
  NAND2_X2 U20636 ( .A1(n16706), .A2(n7190), .ZN(n31664) );
  XOR2_X1 U20638 ( .A1(n10939), .A2(n10239), .Z(n36406) );
  NAND2_X2 U20640 ( .A1(n9166), .A2(n11248), .ZN(n11818) );
  XOR2_X1 U20641 ( .A1(n26302), .A2(n26303), .Z(n26765) );
  XOR2_X1 U20642 ( .A1(n7475), .A2(n30094), .Z(n10100) );
  OAI22_X2 U20645 ( .A1(n35477), .A2(n36103), .B1(n23589), .B2(n2273), .ZN(
        n7475) );
  XOR2_X1 U20649 ( .A1(n26391), .A2(n38140), .Z(n7854) );
  NAND2_X2 U20650 ( .A1(n32897), .A2(n13118), .ZN(n26391) );
  NOR3_X1 U20653 ( .A1(n22940), .A2(n33969), .A3(n6646), .ZN(n38390) );
  XOR2_X1 U20654 ( .A1(n33863), .A2(n22508), .Z(n22765) );
  NOR2_X2 U20657 ( .A1(n14957), .A2(n667), .ZN(n22508) );
  XOR2_X1 U20663 ( .A1(n38392), .A2(n39049), .Z(n5211) );
  XOR2_X1 U20671 ( .A1(n39344), .A2(n5667), .Z(n38392) );
  NOR2_X2 U20674 ( .A1(n26092), .A2(n26093), .ZN(n25852) );
  NAND2_X2 U20675 ( .A1(n4595), .A2(n31165), .ZN(n26093) );
  NAND2_X2 U20676 ( .A1(n10216), .A2(n32366), .ZN(n23595) );
  NAND2_X2 U20681 ( .A1(n400), .A2(n15492), .ZN(n29231) );
  NAND2_X2 U20682 ( .A1(n25047), .A2(n36690), .ZN(n13843) );
  NAND2_X2 U20684 ( .A1(n25048), .A2(n3510), .ZN(n25047) );
  NAND2_X2 U20685 ( .A1(n23502), .A2(n32366), .ZN(n23374) );
  NAND2_X2 U20687 ( .A1(n12254), .A2(n12253), .ZN(n23502) );
  NAND2_X2 U20692 ( .A1(n38394), .A2(n39051), .ZN(n39050) );
  NAND2_X1 U20698 ( .A1(n36623), .A2(n3944), .ZN(n17715) );
  OAI21_X2 U20701 ( .A1(n10587), .A2(n9648), .B(n38396), .ZN(n28521) );
  AOI21_X2 U20702 ( .A1(n38529), .A2(n16295), .B(n37081), .ZN(n38396) );
  XOR2_X1 U20707 ( .A1(n18991), .A2(n32765), .Z(n14023) );
  NOR2_X2 U20708 ( .A1(n12504), .A2(n12503), .ZN(n18991) );
  NAND2_X2 U20714 ( .A1(n38398), .A2(n36277), .ZN(n26054) );
  XNOR2_X1 U20716 ( .A1(n1790), .A2(n24062), .ZN(n38975) );
  XOR2_X1 U20717 ( .A1(n23898), .A2(n23968), .Z(n23812) );
  NAND2_X2 U20721 ( .A1(n23224), .A2(n23223), .ZN(n23898) );
  INV_X2 U20724 ( .I(n17844), .ZN(n20839) );
  XOR2_X1 U20727 ( .A1(n32096), .A2(n18935), .Z(n17844) );
  OAI21_X2 U20733 ( .A1(n38400), .A2(n35880), .B(n23141), .ZN(n31908) );
  NAND3_X2 U20734 ( .A1(n36911), .A2(n39414), .A3(n27240), .ZN(n38525) );
  NAND2_X2 U20736 ( .A1(n38401), .A2(n16305), .ZN(n4391) );
  OAI21_X2 U20740 ( .A1(n21570), .A2(n21599), .B(n21870), .ZN(n38401) );
  XOR2_X1 U20757 ( .A1(n26595), .A2(n7018), .Z(n26491) );
  XOR2_X1 U20767 ( .A1(n4330), .A2(n32954), .Z(n867) );
  XOR2_X1 U20769 ( .A1(n29246), .A2(n38403), .Z(n12069) );
  XOR2_X1 U20773 ( .A1(n29832), .A2(n4905), .Z(n38403) );
  XOR2_X1 U20776 ( .A1(n29021), .A2(n29142), .Z(n10430) );
  NAND3_X2 U20779 ( .A1(n7849), .A2(n15602), .A3(n13422), .ZN(n29021) );
  NOR2_X2 U20780 ( .A1(n39366), .A2(n39365), .ZN(n39364) );
  INV_X2 U20781 ( .I(n38406), .ZN(n14179) );
  XNOR2_X1 U20784 ( .A1(n9435), .A2(n38567), .ZN(n38406) );
  NAND3_X2 U20785 ( .A1(n32833), .A2(n19391), .A3(n1417), .ZN(n1741) );
  NAND3_X2 U20788 ( .A1(n39736), .A2(n5924), .A3(n5923), .ZN(n17730) );
  AOI22_X2 U20792 ( .A1(n31603), .A2(n12081), .B1(n39280), .B2(n19544), .ZN(
        n3464) );
  AOI22_X2 U20793 ( .A1(n31764), .A2(n12156), .B1(n27226), .B2(n10461), .ZN(
        n5983) );
  NOR2_X2 U20796 ( .A1(n10051), .A2(n27184), .ZN(n27226) );
  OR2_X1 U20797 ( .A1(n25782), .A2(n26106), .Z(n11581) );
  OAI21_X2 U20800 ( .A1(n11442), .A2(n11589), .B(n11441), .ZN(n25782) );
  AOI22_X2 U20807 ( .A1(n3899), .A2(n28570), .B1(n3903), .B2(n33995), .ZN(
        n4002) );
  XOR2_X1 U20808 ( .A1(n24053), .A2(n23963), .Z(n23928) );
  NAND2_X2 U20814 ( .A1(n34421), .A2(n38859), .ZN(n24053) );
  NAND2_X2 U20816 ( .A1(n31719), .A2(n26122), .ZN(n38409) );
  XOR2_X1 U20820 ( .A1(n38410), .A2(n16268), .Z(n36463) );
  XOR2_X1 U20825 ( .A1(n36687), .A2(n6795), .Z(n38410) );
  XOR2_X1 U20827 ( .A1(n10226), .A2(n38411), .Z(n39511) );
  XOR2_X1 U20830 ( .A1(n27531), .A2(n27505), .Z(n38411) );
  XOR2_X1 U20832 ( .A1(n24064), .A2(n24002), .Z(n11267) );
  NAND2_X2 U20837 ( .A1(n23019), .A2(n23018), .ZN(n24064) );
  NOR2_X2 U20838 ( .A1(n196), .A2(n1688), .ZN(n13009) );
  OR2_X2 U20841 ( .A1(n38412), .A2(n10821), .Z(n10820) );
  AOI21_X1 U20843 ( .A1(n9466), .A2(n10875), .B(n20810), .ZN(n38412) );
  AOI21_X2 U20844 ( .A1(n2339), .A2(n8154), .B(n38413), .ZN(n38908) );
  NOR2_X1 U20847 ( .A1(n13371), .A2(n4748), .ZN(n38413) );
  NAND4_X2 U20862 ( .A1(n26913), .A2(n26914), .A3(n26915), .A4(n18749), .ZN(
        n27700) );
  NAND2_X2 U20868 ( .A1(n1891), .A2(n38414), .ZN(n18749) );
  INV_X2 U20870 ( .I(n38415), .ZN(n21644) );
  XNOR2_X1 U20872 ( .A1(n21399), .A2(Key[183]), .ZN(n38415) );
  INV_X2 U20877 ( .I(n9303), .ZN(n25753) );
  NAND2_X2 U20879 ( .A1(n25754), .A2(n25699), .ZN(n9303) );
  XOR2_X1 U20881 ( .A1(n14218), .A2(n13883), .Z(n12884) );
  XOR2_X1 U20885 ( .A1(n36566), .A2(n27767), .Z(n14218) );
  XOR2_X1 U20886 ( .A1(n9001), .A2(n17263), .Z(n26570) );
  NOR2_X2 U20891 ( .A1(n13387), .A2(n13388), .ZN(n9001) );
  XOR2_X1 U20897 ( .A1(n35257), .A2(n30063), .Z(n18736) );
  OAI21_X1 U20898 ( .A1(n3361), .A2(n3360), .B(n35646), .ZN(n35257) );
  INV_X2 U20899 ( .I(n29160), .ZN(n973) );
  NAND2_X2 U20900 ( .A1(n39364), .A2(n35351), .ZN(n29160) );
  AOI21_X2 U20902 ( .A1(n24175), .A2(n24328), .B(n6585), .ZN(n11373) );
  NAND2_X2 U20904 ( .A1(n38417), .A2(n14006), .ZN(n15373) );
  NAND3_X2 U20905 ( .A1(n1653), .A2(n6646), .A3(n38725), .ZN(n38417) );
  INV_X2 U20911 ( .I(n9108), .ZN(n1184) );
  XNOR2_X1 U20912 ( .A1(n25298), .A2(n25113), .ZN(n25144) );
  NOR2_X1 U20916 ( .A1(n38418), .A2(n2785), .ZN(n2784) );
  NOR2_X1 U20917 ( .A1(n2788), .A2(n33646), .ZN(n38418) );
  NAND2_X1 U20919 ( .A1(n3443), .A2(n7935), .ZN(n4058) );
  XOR2_X1 U20920 ( .A1(Plaintext[186]), .A2(Key[186]), .Z(n7935) );
  NAND2_X2 U20921 ( .A1(n33224), .A2(n38421), .ZN(n32831) );
  NOR2_X2 U20926 ( .A1(n38423), .A2(n38422), .ZN(n38421) );
  NOR2_X2 U20927 ( .A1(n24155), .A2(n9101), .ZN(n38423) );
  OAI21_X1 U20932 ( .A1(n21464), .A2(n21463), .B(n21645), .ZN(n9495) );
  OAI21_X2 U20933 ( .A1(n8264), .A2(n1570), .B(n30843), .ZN(n38424) );
  NAND2_X2 U20934 ( .A1(n20122), .A2(n39690), .ZN(n3575) );
  XOR2_X1 U20936 ( .A1(n19071), .A2(n23696), .Z(n6943) );
  BUF_X4 U20940 ( .I(n39648), .Z(n38561) );
  NAND3_X2 U20943 ( .A1(n38426), .A2(n25416), .A3(n38425), .ZN(n25509) );
  NAND2_X2 U20945 ( .A1(n9740), .A2(n38178), .ZN(n38426) );
  INV_X4 U20947 ( .I(n26029), .ZN(n16867) );
  NOR2_X2 U20948 ( .A1(n23120), .A2(n15947), .ZN(n31364) );
  NOR3_X2 U20949 ( .A1(n37074), .A2(n26799), .A3(n35282), .ZN(n38755) );
  NOR2_X2 U20956 ( .A1(n849), .A2(n4138), .ZN(n26799) );
  NAND3_X2 U20960 ( .A1(n36393), .A2(n23627), .A3(n36394), .ZN(n33672) );
  NAND2_X2 U20961 ( .A1(n2560), .A2(n2557), .ZN(n29617) );
  NAND2_X2 U20966 ( .A1(n23303), .A2(n11970), .ZN(n23489) );
  XOR2_X1 U20971 ( .A1(n34788), .A2(n24970), .Z(n38427) );
  INV_X2 U20972 ( .I(n38428), .ZN(n25307) );
  XNOR2_X1 U20976 ( .A1(n12592), .A2(n12594), .ZN(n38428) );
  NAND3_X1 U20977 ( .A1(n36737), .A2(n36739), .A3(n30211), .ZN(n38429) );
  OAI21_X2 U20979 ( .A1(n11714), .A2(n10013), .B(n24638), .ZN(n11713) );
  NAND2_X2 U20980 ( .A1(n35960), .A2(n3120), .ZN(n24638) );
  XOR2_X1 U20981 ( .A1(n1561), .A2(n25301), .Z(n8324) );
  XOR2_X1 U20986 ( .A1(n36138), .A2(n20333), .Z(n33505) );
  NAND2_X1 U20991 ( .A1(n3568), .A2(n25728), .ZN(n25729) );
  NOR2_X1 U20993 ( .A1(n14337), .A2(n29722), .ZN(n29709) );
  NAND2_X2 U20996 ( .A1(n1082), .A2(n38211), .ZN(n26807) );
  XOR2_X1 U21000 ( .A1(n10012), .A2(n25136), .Z(n25272) );
  XOR2_X1 U21003 ( .A1(n29045), .A2(n29040), .Z(n18813) );
  NOR2_X2 U21005 ( .A1(n21145), .A2(n20735), .ZN(n29040) );
  AOI21_X1 U21010 ( .A1(n28079), .A2(n987), .B(n883), .ZN(n7220) );
  NAND2_X2 U21011 ( .A1(n1252), .A2(n7986), .ZN(n39294) );
  XOR2_X1 U21029 ( .A1(n16833), .A2(n15974), .Z(n15973) );
  XOR2_X1 U21030 ( .A1(n38433), .A2(n34223), .Z(n8184) );
  XOR2_X1 U21035 ( .A1(n16019), .A2(n35728), .Z(n38433) );
  OR2_X1 U21039 ( .A1(n19135), .A2(n39050), .Z(n35617) );
  XOR2_X1 U21041 ( .A1(n20706), .A2(n38620), .Z(n2283) );
  XOR2_X1 U21047 ( .A1(n3035), .A2(n38434), .Z(n3974) );
  XOR2_X1 U21049 ( .A1(n14784), .A2(n26483), .Z(n38434) );
  INV_X2 U21052 ( .I(n4008), .ZN(n1120) );
  NAND2_X2 U21083 ( .A1(n32018), .A2(n36542), .ZN(n4008) );
  NOR2_X1 U21084 ( .A1(n17934), .A2(n10523), .ZN(n10524) );
  XOR2_X1 U21085 ( .A1(n17920), .A2(n17922), .Z(n17934) );
  XOR2_X1 U21089 ( .A1(n26391), .A2(n10225), .Z(n15288) );
  AOI22_X2 U21099 ( .A1(n21421), .A2(n10924), .B1(n21983), .B2(n37176), .ZN(
        n33736) );
  XOR2_X1 U21102 ( .A1(n13978), .A2(n16324), .Z(n13977) );
  NAND2_X2 U21112 ( .A1(n11529), .A2(n11530), .ZN(n16324) );
  NAND2_X2 U21113 ( .A1(n30795), .A2(n7978), .ZN(n30539) );
  NOR2_X2 U21114 ( .A1(n36626), .A2(n38436), .ZN(n39098) );
  AOI22_X2 U21115 ( .A1(n626), .A2(n10342), .B1(n11673), .B2(n3398), .ZN(
        n38436) );
  XOR2_X1 U21116 ( .A1(n27809), .A2(n27615), .Z(n8336) );
  XOR2_X1 U21117 ( .A1(n27542), .A2(n6033), .Z(n27809) );
  NAND2_X2 U21118 ( .A1(n39357), .A2(n4339), .ZN(n34195) );
  NAND2_X2 U21129 ( .A1(n38439), .A2(n38438), .ZN(n9539) );
  INV_X1 U21130 ( .I(n7982), .ZN(n38438) );
  XOR2_X1 U21131 ( .A1(n37338), .A2(n16162), .Z(n38440) );
  OR2_X2 U21133 ( .A1(n36868), .A2(n36355), .Z(n3574) );
  XOR2_X1 U21135 ( .A1(n19830), .A2(n20779), .Z(n9780) );
  INV_X1 U21137 ( .I(n23349), .ZN(n38441) );
  NOR2_X2 U21140 ( .A1(n10724), .A2(n38953), .ZN(n4248) );
  INV_X2 U21141 ( .I(n20691), .ZN(n39023) );
  NAND2_X2 U21143 ( .A1(n38618), .A2(n4014), .ZN(n20691) );
  OAI21_X2 U21145 ( .A1(n37203), .A2(n38463), .B(n38442), .ZN(n12741) );
  AOI22_X2 U21151 ( .A1(n10910), .A2(n34737), .B1(n10908), .B2(n28608), .ZN(
        n38442) );
  NAND3_X1 U21156 ( .A1(n11039), .A2(n13753), .A3(n35114), .ZN(n26844) );
  XOR2_X1 U21157 ( .A1(n13193), .A2(n6561), .Z(n31581) );
  NAND2_X2 U21158 ( .A1(n12822), .A2(n9968), .ZN(n13193) );
  OAI22_X2 U21159 ( .A1(n10458), .A2(n10457), .B1(n17502), .B2(n12522), .ZN(
        n31293) );
  AOI21_X2 U21170 ( .A1(n33264), .A2(n34598), .B(n38444), .ZN(n24661) );
  OAI22_X2 U21171 ( .A1(n7086), .A2(n15968), .B1(n14004), .B2(n24403), .ZN(
        n38444) );
  NAND2_X2 U21176 ( .A1(n35258), .A2(n36865), .ZN(n38638) );
  AOI22_X2 U21177 ( .A1(n25445), .A2(n32520), .B1(n33011), .B2(n33815), .ZN(
        n38672) );
  XOR2_X1 U21179 ( .A1(n3609), .A2(n5323), .Z(n23959) );
  NAND2_X2 U21182 ( .A1(n35864), .A2(n4251), .ZN(n3609) );
  INV_X2 U21184 ( .I(n38445), .ZN(n1230) );
  AND2_X1 U21185 ( .A1(n32043), .A2(n9958), .Z(n36995) );
  XOR2_X1 U21188 ( .A1(n18547), .A2(n12304), .Z(n32043) );
  XNOR2_X1 U21189 ( .A1(n12969), .A2(n15500), .ZN(n39245) );
  NAND2_X2 U21190 ( .A1(n33187), .A2(n38446), .ZN(n32898) );
  NAND2_X1 U21194 ( .A1(n367), .A2(n39176), .ZN(n4495) );
  AOI21_X2 U21196 ( .A1(n22262), .A2(n33738), .B(n33086), .ZN(n4339) );
  INV_X4 U21199 ( .I(n33748), .ZN(n33086) );
  AOI22_X2 U21200 ( .A1(n36578), .A2(n15099), .B1(n34048), .B2(n15096), .ZN(
        n33748) );
  OAI22_X2 U21202 ( .A1(n31147), .A2(n32012), .B1(n28614), .B2(n4002), .ZN(
        n5115) );
  XOR2_X1 U21203 ( .A1(n39282), .A2(n5114), .Z(n31329) );
  OR2_X1 U21204 ( .A1(n5112), .A2(n3675), .Z(n32449) );
  OR2_X2 U21207 ( .A1(n21722), .A2(n3507), .Z(n11852) );
  OAI22_X2 U21209 ( .A1(n28652), .A2(n35830), .B1(n28650), .B2(n30931), .ZN(
        n13027) );
  NAND3_X2 U21210 ( .A1(n14750), .A2(n14749), .A3(n22995), .ZN(n14748) );
  NAND2_X2 U21212 ( .A1(n6674), .A2(n20449), .ZN(n14750) );
  AOI22_X2 U21218 ( .A1(n11331), .A2(n4642), .B1(n11333), .B2(n13015), .ZN(
        n31367) );
  AOI22_X2 U21220 ( .A1(n39226), .A2(n579), .B1(n32684), .B2(n31721), .ZN(
        n5787) );
  NOR2_X2 U21222 ( .A1(n12675), .A2(n12931), .ZN(n579) );
  NAND3_X2 U21223 ( .A1(n26979), .A2(n17252), .A3(n17097), .ZN(n38450) );
  XOR2_X1 U21228 ( .A1(n28933), .A2(n28869), .Z(n36706) );
  XOR2_X1 U21231 ( .A1(n18785), .A2(n29070), .Z(n28933) );
  OAI21_X2 U21235 ( .A1(n23182), .A2(n32270), .B(n37137), .ZN(n23183) );
  NAND2_X2 U21239 ( .A1(n38451), .A2(n15583), .ZN(n31751) );
  NAND3_X2 U21243 ( .A1(n39585), .A2(n38834), .A3(n38328), .ZN(n38451) );
  OR2_X1 U21246 ( .A1(n24473), .A2(n7240), .Z(n38474) );
  NAND2_X2 U21252 ( .A1(n28066), .A2(n14500), .ZN(n5430) );
  AND2_X1 U21254 ( .A1(n20077), .A2(n32537), .Z(n22940) );
  CLKBUF_X4 U21255 ( .I(n26833), .Z(n38852) );
  INV_X4 U21263 ( .I(n38452), .ZN(n15573) );
  AND3_X2 U21265 ( .A1(n11648), .A2(n11649), .A3(n15446), .Z(n38452) );
  XOR2_X1 U21266 ( .A1(n34876), .A2(n36114), .Z(n38453) );
  XOR2_X1 U21269 ( .A1(n28949), .A2(n28950), .Z(n33434) );
  XOR2_X1 U21271 ( .A1(n38454), .A2(n19810), .Z(n26803) );
  XOR2_X1 U21273 ( .A1(n25986), .A2(n25985), .Z(n38454) );
  XOR2_X1 U21274 ( .A1(n32613), .A2(n11401), .Z(n38455) );
  AOI21_X2 U21279 ( .A1(n7978), .A2(n30795), .B(n26700), .ZN(n32262) );
  NAND2_X2 U21280 ( .A1(n39144), .A2(n38456), .ZN(n33258) );
  OAI21_X2 U21282 ( .A1(n39223), .A2(n39224), .B(n7986), .ZN(n38456) );
  NOR2_X2 U21287 ( .A1(n4427), .A2(n4062), .ZN(n25146) );
  XOR2_X1 U21290 ( .A1(n31227), .A2(n476), .Z(n4612) );
  XOR2_X1 U21292 ( .A1(n13649), .A2(n38457), .Z(n19658) );
  XOR2_X1 U21293 ( .A1(n23723), .A2(n23741), .Z(n38457) );
  XOR2_X1 U21294 ( .A1(n24992), .A2(n15186), .Z(n38458) );
  XOR2_X1 U21295 ( .A1(n39163), .A2(n23675), .Z(n34269) );
  NAND2_X2 U21299 ( .A1(n34884), .A2(n20984), .ZN(n23675) );
  NAND2_X1 U21303 ( .A1(n20619), .A2(n24470), .ZN(n36790) );
  NAND2_X2 U21304 ( .A1(n39643), .A2(n28392), .ZN(n6093) );
  NOR2_X2 U21305 ( .A1(n38460), .A2(n38459), .ZN(n19260) );
  AOI21_X2 U21307 ( .A1(n18997), .A2(n31583), .B(n29587), .ZN(n38459) );
  AOI21_X2 U21308 ( .A1(n20371), .A2(n29630), .B(n21264), .ZN(n38460) );
  XOR2_X1 U21309 ( .A1(n37874), .A2(n15682), .Z(n28845) );
  XNOR2_X1 U21310 ( .A1(n29048), .A2(n19843), .ZN(n38606) );
  NAND2_X2 U21311 ( .A1(n1904), .A2(n21287), .ZN(n6601) );
  OAI22_X2 U21312 ( .A1(n11861), .A2(n29946), .B1(n16510), .B2(n17240), .ZN(
        n1904) );
  XOR2_X1 U21315 ( .A1(n18001), .A2(n14173), .Z(n9943) );
  XOR2_X1 U21321 ( .A1(n27777), .A2(n38158), .Z(n5524) );
  XOR2_X1 U21342 ( .A1(n18160), .A2(n23707), .Z(n23997) );
  AOI21_X2 U21343 ( .A1(n9971), .A2(n1307), .B(n23442), .ZN(n18160) );
  AOI22_X2 U21347 ( .A1(n22977), .A2(n10828), .B1(n10470), .B2(n7266), .ZN(
        n10469) );
  NAND3_X2 U21350 ( .A1(n33669), .A2(n17532), .A3(n28163), .ZN(n31882) );
  NOR2_X1 U21355 ( .A1(n4713), .A2(n38513), .ZN(n15947) );
  AOI21_X1 U21356 ( .A1(n7789), .A2(n10702), .B(n29059), .ZN(n11777) );
  NAND2_X2 U21358 ( .A1(n2182), .A2(n36720), .ZN(n23373) );
  XOR2_X1 U21361 ( .A1(n38462), .A2(n1161), .Z(Ciphertext[171]) );
  OAI21_X1 U21366 ( .A1(n39079), .A2(n2506), .B(n2945), .ZN(n2203) );
  INV_X2 U21370 ( .I(n35813), .ZN(n24788) );
  OR2_X1 U21371 ( .A1(n12246), .A2(n31682), .Z(n12192) );
  XOR2_X1 U21372 ( .A1(n38464), .A2(n25090), .Z(n25159) );
  INV_X2 U21374 ( .I(n25133), .ZN(n38464) );
  NAND2_X2 U21379 ( .A1(n7064), .A2(n31290), .ZN(n25090) );
  XOR2_X1 U21380 ( .A1(n14719), .A2(n38465), .Z(n39277) );
  NAND2_X2 U21386 ( .A1(n38466), .A2(n13870), .ZN(n34644) );
  NOR2_X2 U21387 ( .A1(n31705), .A2(n11800), .ZN(n11695) );
  AOI22_X2 U21388 ( .A1(n1077), .A2(n9315), .B1(n20976), .B2(n10573), .ZN(
        n10579) );
  NAND2_X2 U21389 ( .A1(n1570), .A2(n257), .ZN(n12124) );
  XOR2_X1 U21392 ( .A1(n24711), .A2(n25192), .Z(n20554) );
  INV_X2 U21395 ( .I(n38467), .ZN(n8479) );
  NAND2_X2 U21396 ( .A1(n39131), .A2(n12133), .ZN(n11698) );
  NOR2_X2 U21405 ( .A1(n36964), .A2(n10708), .ZN(n35181) );
  XOR2_X1 U21408 ( .A1(n22635), .A2(n22633), .Z(n32847) );
  XOR2_X1 U21410 ( .A1(n22776), .A2(n22731), .Z(n22633) );
  NOR2_X1 U21411 ( .A1(n36786), .A2(n36787), .ZN(n39731) );
  AOI21_X2 U21419 ( .A1(n11424), .A2(n20336), .B(n11423), .ZN(n26278) );
  NAND3_X2 U21426 ( .A1(n20470), .A2(n39382), .A3(n27620), .ZN(n20662) );
  INV_X2 U21428 ( .I(n38470), .ZN(n28188) );
  NAND2_X1 U21429 ( .A1(n5101), .A2(n7542), .ZN(n36981) );
  AOI21_X2 U21437 ( .A1(n10521), .A2(n20064), .B(n10159), .ZN(n10520) );
  XOR2_X1 U21439 ( .A1(n18133), .A2(n38471), .Z(n38927) );
  XOR2_X1 U21440 ( .A1(n29113), .A2(n29983), .Z(n38471) );
  XOR2_X1 U21442 ( .A1(n29105), .A2(n16529), .Z(n12402) );
  NAND2_X1 U21443 ( .A1(n32649), .A2(n32648), .ZN(n39722) );
  NAND2_X2 U21444 ( .A1(n38474), .A2(n38472), .ZN(n10626) );
  NAND2_X2 U21447 ( .A1(n1081), .A2(n3851), .ZN(n3850) );
  OR2_X2 U21452 ( .A1(n28204), .A2(n21159), .Z(n9089) );
  XOR2_X1 U21457 ( .A1(n38205), .A2(n15219), .Z(n10412) );
  NOR2_X2 U21460 ( .A1(n38910), .A2(n3849), .ZN(n15219) );
  XOR2_X1 U21461 ( .A1(n5412), .A2(n33701), .Z(n5410) );
  NOR2_X2 U21463 ( .A1(n12447), .A2(n24174), .ZN(n39480) );
  NAND2_X2 U21465 ( .A1(n1607), .A2(n37954), .ZN(n12447) );
  NOR2_X2 U21467 ( .A1(n38475), .A2(n34042), .ZN(n12676) );
  XOR2_X1 U21471 ( .A1(n12973), .A2(n24058), .Z(n9548) );
  XOR2_X1 U21473 ( .A1(n2443), .A2(n1502), .Z(n2545) );
  OAI21_X2 U21479 ( .A1(n32712), .A2(n15284), .B(n12031), .ZN(n21140) );
  AOI21_X2 U21494 ( .A1(n8393), .A2(n2629), .B(n1742), .ZN(n35209) );
  AOI21_X2 U21498 ( .A1(n2865), .A2(n17269), .B(n930), .ZN(n1742) );
  NAND2_X2 U21500 ( .A1(n38478), .A2(n30850), .ZN(n24799) );
  XOR2_X1 U21504 ( .A1(n27760), .A2(n27413), .Z(n38624) );
  XOR2_X1 U21505 ( .A1(n27731), .A2(n7755), .Z(n27413) );
  NAND2_X2 U21507 ( .A1(n38479), .A2(n39592), .ZN(n2668) );
  XOR2_X1 U21509 ( .A1(n27778), .A2(n21093), .Z(n27515) );
  NAND2_X2 U21516 ( .A1(n10953), .A2(n36492), .ZN(n21093) );
  XOR2_X1 U21520 ( .A1(n29257), .A2(n29085), .Z(n17659) );
  XOR2_X1 U21522 ( .A1(n24030), .A2(n23883), .Z(n24001) );
  NOR2_X2 U21525 ( .A1(n1302), .A2(n1297), .ZN(n8390) );
  NAND2_X2 U21526 ( .A1(n23467), .A2(n16528), .ZN(n18989) );
  NOR2_X2 U21528 ( .A1(n38559), .A2(n6970), .ZN(n23467) );
  NAND2_X2 U21529 ( .A1(n14496), .A2(n20576), .ZN(n36969) );
  XOR2_X1 U21530 ( .A1(n20695), .A2(n24056), .Z(n39201) );
  XOR2_X1 U21531 ( .A1(n1613), .A2(n16138), .Z(n20695) );
  XOR2_X1 U21533 ( .A1(n39078), .A2(n17650), .Z(n19443) );
  OAI21_X2 U21541 ( .A1(n31470), .A2(n31471), .B(n10511), .ZN(n17650) );
  XOR2_X1 U21542 ( .A1(n38485), .A2(n22506), .Z(n2046) );
  XOR2_X1 U21557 ( .A1(n16912), .A2(n22701), .Z(n38485) );
  XOR2_X1 U21561 ( .A1(n20205), .A2(n24011), .Z(n23729) );
  NAND2_X2 U21564 ( .A1(n7482), .A2(n23422), .ZN(n20205) );
  XOR2_X1 U21566 ( .A1(n38510), .A2(n15857), .Z(n39285) );
  XOR2_X1 U21568 ( .A1(n38486), .A2(n7558), .Z(n12519) );
  XOR2_X1 U21569 ( .A1(n25031), .A2(n32433), .Z(n25167) );
  NAND2_X2 U21572 ( .A1(n17916), .A2(n4937), .ZN(n38493) );
  BUF_X2 U21573 ( .I(n17263), .Z(n38495) );
  NAND2_X1 U21578 ( .A1(n9836), .A2(n11777), .ZN(n39586) );
  OAI21_X2 U21581 ( .A1(n123), .A2(n683), .B(n38496), .ZN(n32763) );
  XOR2_X1 U21585 ( .A1(n3495), .A2(n38497), .Z(n8128) );
  XOR2_X1 U21592 ( .A1(n32346), .A2(n3493), .Z(n38497) );
  NAND2_X2 U21595 ( .A1(n9242), .A2(n36197), .ZN(n3983) );
  BUF_X1 U21596 ( .I(n6002), .Z(n35264) );
  INV_X2 U21598 ( .I(n38854), .ZN(n3899) );
  AOI22_X2 U21602 ( .A1(n2614), .A2(n17532), .B1(n33669), .B2(n2613), .ZN(
        n38596) );
  INV_X2 U21604 ( .I(n23550), .ZN(n38499) );
  AOI21_X2 U21616 ( .A1(n35191), .A2(n38499), .B(n37814), .ZN(n38615) );
  INV_X2 U21620 ( .I(n30981), .ZN(n27366) );
  NAND2_X2 U21621 ( .A1(n21101), .A2(n27363), .ZN(n30981) );
  XOR2_X1 U21622 ( .A1(n8059), .A2(n27862), .Z(n27642) );
  BUF_X2 U21625 ( .I(n26551), .Z(n38502) );
  OAI21_X2 U21626 ( .A1(n37249), .A2(n38503), .B(n9598), .ZN(n34463) );
  AND2_X1 U21627 ( .A1(n32080), .A2(n36463), .Z(n28288) );
  NOR2_X2 U21628 ( .A1(n33752), .A2(n6589), .ZN(n26481) );
  OAI21_X2 U21629 ( .A1(n4371), .A2(n4369), .B(n38504), .ZN(n28305) );
  XOR2_X1 U21634 ( .A1(n38624), .A2(n38505), .Z(n17777) );
  XOR2_X1 U21639 ( .A1(n12165), .A2(n27495), .Z(n38505) );
  INV_X2 U21650 ( .I(n24812), .ZN(n32651) );
  XOR2_X1 U21651 ( .A1(n10767), .A2(n13483), .Z(n13090) );
  XOR2_X1 U21654 ( .A1(n6384), .A2(n11753), .Z(n13483) );
  AOI22_X2 U21660 ( .A1(n28282), .A2(n28283), .B1(n36877), .B2(n16544), .ZN(
        n12787) );
  NAND2_X2 U21664 ( .A1(n33314), .A2(n38487), .ZN(n24121) );
  XOR2_X1 U21666 ( .A1(n27749), .A2(n38225), .Z(n3889) );
  XOR2_X1 U21674 ( .A1(n33645), .A2(n30170), .Z(n10492) );
  INV_X4 U21676 ( .I(n19255), .ZN(n31698) );
  NAND2_X2 U21677 ( .A1(n24455), .A2(n24456), .ZN(n19255) );
  NAND2_X2 U21678 ( .A1(n5264), .A2(n16859), .ZN(n27379) );
  AND2_X1 U21684 ( .A1(n585), .A2(n17871), .Z(n35075) );
  OAI22_X2 U21693 ( .A1(n15445), .A2(n25362), .B1(n15444), .B2(n19095), .ZN(
        n35003) );
  OAI21_X2 U21694 ( .A1(n28187), .A2(n14642), .B(n33002), .ZN(n38506) );
  NOR2_X2 U21696 ( .A1(n9969), .A2(n28191), .ZN(n28187) );
  NAND2_X2 U21697 ( .A1(n38506), .A2(n14030), .ZN(n13594) );
  NAND2_X2 U21698 ( .A1(n13492), .A2(n38947), .ZN(n38946) );
  XOR2_X1 U21700 ( .A1(n24961), .A2(n13634), .Z(n25262) );
  NAND2_X2 U21701 ( .A1(n62), .A2(n35022), .ZN(n13634) );
  XOR2_X1 U21702 ( .A1(n12749), .A2(n15265), .Z(n15261) );
  NAND2_X1 U21707 ( .A1(n3016), .A2(n24178), .ZN(n38508) );
  NAND3_X2 U21708 ( .A1(n18202), .A2(n28746), .A3(n18201), .ZN(n19408) );
  XOR2_X1 U21710 ( .A1(n19561), .A2(n35229), .Z(n4266) );
  XOR2_X1 U21711 ( .A1(n23688), .A2(n34435), .Z(n2695) );
  NOR2_X2 U21712 ( .A1(n38509), .A2(n35944), .ZN(n12910) );
  XOR2_X1 U21718 ( .A1(n25154), .A2(n38511), .Z(n38510) );
  XOR2_X1 U21720 ( .A1(n11756), .A2(n12233), .Z(n24610) );
  NAND3_X1 U21723 ( .A1(n15541), .A2(n37050), .A3(n826), .ZN(n12578) );
  CLKBUF_X2 U21725 ( .I(n22929), .Z(n39518) );
  NAND2_X2 U21729 ( .A1(n38549), .A2(n13454), .ZN(n8412) );
  NAND2_X2 U21731 ( .A1(n30302), .A2(n2029), .ZN(n26114) );
  NAND2_X2 U21740 ( .A1(n31964), .A2(n31963), .ZN(n2029) );
  BUF_X2 U21747 ( .I(n26530), .Z(n38514) );
  XOR2_X1 U21751 ( .A1(n15401), .A2(n38515), .Z(n27474) );
  NAND2_X2 U21755 ( .A1(n11855), .A2(n13211), .ZN(n15401) );
  XOR2_X1 U21757 ( .A1(n27542), .A2(n37101), .Z(n39515) );
  NAND2_X1 U21760 ( .A1(n16444), .A2(n25767), .ZN(n34595) );
  NAND2_X1 U21765 ( .A1(n28322), .A2(n14448), .ZN(n30380) );
  OAI21_X1 U21766 ( .A1(n25488), .A2(n32775), .B(n25487), .ZN(n32879) );
  XOR2_X1 U21767 ( .A1(n16696), .A2(n16698), .Z(n34561) );
  NAND3_X2 U21768 ( .A1(n38516), .A2(n38525), .A3(n27242), .ZN(n27528) );
  XOR2_X1 U21769 ( .A1(n38517), .A2(n38518), .Z(n28182) );
  XOR2_X1 U21770 ( .A1(n15844), .A2(n15785), .Z(n38517) );
  XOR2_X1 U21772 ( .A1(n27515), .A2(n763), .Z(n38518) );
  NAND2_X2 U21773 ( .A1(n12287), .A2(n24159), .ZN(n24903) );
  OAI21_X2 U21777 ( .A1(n30388), .A2(n25566), .B(n38520), .ZN(n14212) );
  OAI21_X2 U21779 ( .A1(n33897), .A2(n15459), .B(n10723), .ZN(n38520) );
  INV_X1 U21780 ( .I(n25170), .ZN(n1930) );
  BUF_X2 U21784 ( .I(n17101), .Z(n38523) );
  BUF_X2 U21786 ( .I(n23190), .Z(n38524) );
  NAND2_X2 U21787 ( .A1(n18632), .A2(n38526), .ZN(n17607) );
  NOR2_X2 U21792 ( .A1(n35314), .A2(n9135), .ZN(n38528) );
  NAND2_X2 U21798 ( .A1(n12074), .A2(n8696), .ZN(n32588) );
  INV_X2 U21801 ( .I(n14349), .ZN(n22323) );
  NAND2_X2 U21802 ( .A1(n21516), .A2(n16961), .ZN(n14349) );
  XOR2_X1 U21804 ( .A1(n11881), .A2(n38530), .Z(n11880) );
  BUF_X2 U21807 ( .I(n5859), .Z(n38531) );
  OAI22_X2 U21808 ( .A1(n14535), .A2(n17537), .B1(n17536), .B2(n37920), .ZN(
        n22411) );
  XOR2_X1 U21813 ( .A1(n29092), .A2(n29096), .Z(n29027) );
  NAND2_X2 U21814 ( .A1(n35583), .A2(n14929), .ZN(n29092) );
  XOR2_X1 U21816 ( .A1(n32608), .A2(n28851), .Z(n29073) );
  OAI21_X2 U21817 ( .A1(n12608), .A2(n12609), .B(n28524), .ZN(n28851) );
  XOR2_X1 U21818 ( .A1(n557), .A2(n34963), .Z(n11828) );
  INV_X2 U21819 ( .I(n39810), .ZN(n19082) );
  XOR2_X1 U21827 ( .A1(n4658), .A2(n35129), .Z(n33808) );
  AOI21_X2 U21828 ( .A1(n1966), .A2(n22148), .B(n1965), .ZN(n359) );
  XOR2_X1 U21833 ( .A1(n38532), .A2(n11922), .Z(n11350) );
  XOR2_X1 U21834 ( .A1(n9777), .A2(n5542), .Z(n38532) );
  XOR2_X1 U21835 ( .A1(n23835), .A2(n20486), .Z(n17492) );
  NOR2_X1 U21840 ( .A1(n32043), .A2(n36136), .ZN(n28028) );
  XOR2_X1 U21841 ( .A1(n23743), .A2(n18980), .Z(n1969) );
  NOR3_X2 U21842 ( .A1(n33793), .A2(n30334), .A3(n38533), .ZN(n33116) );
  NOR3_X2 U21847 ( .A1(n33629), .A2(n18281), .A3(n17735), .ZN(n38533) );
  XOR2_X1 U21856 ( .A1(n29294), .A2(n28957), .Z(n5782) );
  XOR2_X1 U21859 ( .A1(n16771), .A2(n29242), .Z(n28957) );
  NAND2_X1 U21864 ( .A1(n38535), .A2(n39001), .ZN(n38534) );
  INV_X2 U21866 ( .I(n12396), .ZN(n38535) );
  OAI21_X2 U21874 ( .A1(n38537), .A2(n3899), .B(n39020), .ZN(n3390) );
  INV_X2 U21876 ( .I(n33995), .ZN(n38537) );
  NAND2_X2 U21883 ( .A1(n38713), .A2(n36472), .ZN(n9802) );
  NAND2_X1 U21884 ( .A1(n214), .A2(n38538), .ZN(n2630) );
  NAND2_X1 U21886 ( .A1(n20418), .A2(n38981), .ZN(n38538) );
  OAI21_X1 U21888 ( .A1(n27403), .A2(n36865), .B(n994), .ZN(n33887) );
  INV_X4 U21890 ( .I(n13730), .ZN(n27403) );
  NAND3_X2 U21892 ( .A1(n33567), .A2(n26816), .A3(n16573), .ZN(n13730) );
  XOR2_X1 U21893 ( .A1(n18600), .A2(n38192), .Z(n16133) );
  XOR2_X1 U21898 ( .A1(n33582), .A2(n38539), .Z(n33601) );
  INV_X1 U21902 ( .I(n29043), .ZN(n38539) );
  NAND2_X2 U21906 ( .A1(n14286), .A2(n9714), .ZN(n5848) );
  NAND2_X2 U21911 ( .A1(n10323), .A2(n38540), .ZN(n22353) );
  OAI22_X1 U21918 ( .A1(n21867), .A2(n17948), .B1(n19549), .B2(n21868), .ZN(
        n38540) );
  OAI22_X2 U21920 ( .A1(n16887), .A2(n38541), .B1(n39526), .B2(n23056), .ZN(
        n35915) );
  OAI22_X2 U21922 ( .A1(n12710), .A2(n25862), .B1(n12712), .B2(n12711), .ZN(
        n26227) );
  NOR2_X2 U21926 ( .A1(n21181), .A2(n36846), .ZN(n27484) );
  OAI22_X1 U21927 ( .A1(n27332), .A2(n27333), .B1(n35115), .B2(n27331), .ZN(
        n27336) );
  XOR2_X1 U21928 ( .A1(n6427), .A2(n6430), .Z(n20080) );
  AOI22_X2 U21929 ( .A1(n7255), .A2(n39298), .B1(n37661), .B2(n9655), .ZN(
        n31785) );
  OAI21_X2 U21930 ( .A1(n5642), .A2(n14398), .B(n34774), .ZN(n33509) );
  NAND2_X2 U21933 ( .A1(n15713), .A2(n15716), .ZN(n39406) );
  NAND2_X2 U21948 ( .A1(n35301), .A2(n2953), .ZN(n23419) );
  XOR2_X1 U21949 ( .A1(n751), .A2(n38543), .Z(n851) );
  XOR2_X1 U21950 ( .A1(n26441), .A2(n29718), .Z(n38543) );
  NOR2_X2 U21953 ( .A1(n39618), .A2(n38544), .ZN(n18656) );
  NAND2_X2 U21961 ( .A1(n38547), .A2(n38545), .ZN(n38544) );
  XOR2_X1 U21963 ( .A1(n20392), .A2(n11974), .Z(n22452) );
  XOR2_X1 U21965 ( .A1(n35209), .A2(n14346), .Z(n5688) );
  NOR2_X2 U21966 ( .A1(n14226), .A2(n14224), .ZN(n14346) );
  NOR2_X2 U21968 ( .A1(n20566), .A2(n29346), .ZN(n39033) );
  INV_X2 U21971 ( .I(n13815), .ZN(n20566) );
  XOR2_X1 U21982 ( .A1(n9972), .A2(n11946), .Z(n13815) );
  NOR2_X2 U21985 ( .A1(n38551), .A2(n38550), .ZN(n14088) );
  INV_X2 U21986 ( .I(n12199), .ZN(n38551) );
  NAND2_X2 U21987 ( .A1(n38552), .A2(n26090), .ZN(n39158) );
  NAND2_X2 U21991 ( .A1(n4852), .A2(n25882), .ZN(n38552) );
  NOR2_X1 U21993 ( .A1(n32682), .A2(n9686), .ZN(n28625) );
  XOR2_X1 U21997 ( .A1(n38553), .A2(n30781), .Z(n31426) );
  XOR2_X1 U21998 ( .A1(n27709), .A2(n27718), .Z(n38553) );
  INV_X2 U22000 ( .I(n38554), .ZN(n27894) );
  NAND2_X1 U22002 ( .A1(n38611), .A2(n1627), .ZN(n14746) );
  NOR2_X2 U22007 ( .A1(n436), .A2(n39318), .ZN(n6405) );
  XOR2_X1 U22009 ( .A1(n38796), .A2(n12322), .Z(n10029) );
  XOR2_X1 U22010 ( .A1(n26288), .A2(n38753), .Z(n12322) );
  NAND2_X2 U22017 ( .A1(n25836), .A2(n19580), .ZN(n25808) );
  XOR2_X1 U22019 ( .A1(n24947), .A2(n24948), .Z(n24949) );
  XOR2_X1 U22021 ( .A1(n23902), .A2(n18160), .Z(n6987) );
  AOI21_X2 U22022 ( .A1(n4528), .A2(n1132), .B(n4526), .ZN(n23902) );
  XOR2_X1 U22023 ( .A1(n8324), .A2(n15011), .Z(n4869) );
  XNOR2_X1 U22035 ( .A1(n25221), .A2(n31579), .ZN(n38563) );
  BUF_X2 U22036 ( .I(n4108), .Z(n38555) );
  NAND2_X2 U22038 ( .A1(n38557), .A2(n22834), .ZN(n33257) );
  INV_X2 U22040 ( .I(n22829), .ZN(n38557) );
  NOR2_X2 U22047 ( .A1(n39096), .A2(n33431), .ZN(n22829) );
  INV_X4 U22051 ( .I(n38907), .ZN(n13973) );
  XOR2_X1 U22052 ( .A1(n28845), .A2(n38885), .Z(n34477) );
  XNOR2_X1 U22053 ( .A1(n38212), .A2(n1375), .ZN(n39335) );
  INV_X1 U22056 ( .I(n6591), .ZN(n37025) );
  XOR2_X1 U22062 ( .A1(n6593), .A2(n38558), .Z(n6591) );
  XOR2_X1 U22063 ( .A1(n9979), .A2(n24070), .Z(n208) );
  NAND2_X2 U22064 ( .A1(n18485), .A2(n39056), .ZN(n9979) );
  NOR2_X1 U22073 ( .A1(n29752), .A2(n29751), .ZN(n29758) );
  XOR2_X1 U22075 ( .A1(n7710), .A2(n29833), .Z(n7004) );
  AOI22_X2 U22078 ( .A1(n2125), .A2(n2124), .B1(n32385), .B2(n36722), .ZN(
        n19384) );
  NAND3_X1 U22079 ( .A1(n24098), .A2(n20517), .A3(n20041), .ZN(n6912) );
  XOR2_X1 U22082 ( .A1(n35842), .A2(n38562), .Z(n38966) );
  XOR2_X1 U22083 ( .A1(n25222), .A2(n38563), .Z(n38562) );
  XOR2_X1 U22084 ( .A1(n3232), .A2(n38564), .Z(n32599) );
  XOR2_X1 U22085 ( .A1(n22690), .A2(n32331), .Z(n38564) );
  NAND2_X2 U22086 ( .A1(n38565), .A2(n27102), .ZN(n36287) );
  XOR2_X1 U22087 ( .A1(n28951), .A2(n5862), .Z(n38567) );
  NOR2_X1 U22090 ( .A1(n36633), .A2(n30805), .ZN(n38924) );
  XOR2_X1 U22091 ( .A1(n25249), .A2(n17623), .Z(n38569) );
  NOR2_X2 U22094 ( .A1(n36850), .A2(n2160), .ZN(n12272) );
  INV_X1 U22097 ( .I(n29968), .ZN(n5678) );
  NAND2_X2 U22101 ( .A1(n34460), .A2(n39525), .ZN(n29968) );
  NAND2_X2 U22104 ( .A1(n38570), .A2(n31606), .ZN(n9917) );
  NOR2_X2 U22105 ( .A1(n32657), .A2(n33292), .ZN(n38570) );
  NOR2_X1 U22106 ( .A1(n25665), .A2(n20441), .ZN(n19336) );
  XOR2_X1 U22107 ( .A1(n11425), .A2(n3413), .Z(n20540) );
  NOR2_X2 U22111 ( .A1(n12456), .A2(n12458), .ZN(n11425) );
  OAI21_X2 U22112 ( .A1(n31530), .A2(n3112), .B(n3111), .ZN(n3110) );
  OAI21_X2 U22114 ( .A1(n38060), .A2(n18228), .B(n20671), .ZN(n38572) );
  XOR2_X1 U22117 ( .A1(n762), .A2(n2437), .Z(n2436) );
  XOR2_X1 U22119 ( .A1(n27546), .A2(n35998), .Z(n762) );
  NOR2_X2 U22120 ( .A1(n38573), .A2(n5738), .ZN(n31656) );
  NOR2_X2 U22134 ( .A1(n28712), .A2(n36414), .ZN(n38573) );
  NAND2_X1 U22142 ( .A1(n34254), .A2(n32468), .ZN(n39777) );
  NOR2_X2 U22144 ( .A1(n16682), .A2(n15867), .ZN(n3377) );
  XOR2_X1 U22148 ( .A1(n23997), .A2(n36233), .Z(n39665) );
  INV_X2 U22150 ( .I(n38575), .ZN(n34178) );
  XOR2_X1 U22152 ( .A1(n38575), .A2(n29054), .Z(n34091) );
  NAND2_X2 U22157 ( .A1(n36585), .A2(n15312), .ZN(n38575) );
  OAI21_X2 U22162 ( .A1(n36342), .A2(n33101), .B(n36341), .ZN(n38576) );
  NAND2_X1 U22163 ( .A1(n20793), .A2(n29769), .ZN(n29770) );
  NAND2_X2 U22164 ( .A1(n17373), .A2(n13389), .ZN(n17263) );
  NOR2_X2 U22165 ( .A1(n31393), .A2(n39453), .ZN(n33961) );
  AND2_X1 U22169 ( .A1(n7993), .A2(n14463), .Z(n14655) );
  OR2_X2 U22173 ( .A1(n38214), .A2(n14061), .Z(n16773) );
  NAND2_X2 U22177 ( .A1(n39464), .A2(n9608), .ZN(n23535) );
  OAI21_X1 U22178 ( .A1(n24764), .A2(n39098), .B(n7852), .ZN(n32221) );
  NAND2_X2 U22179 ( .A1(n32035), .A2(n25808), .ZN(n15298) );
  NAND2_X1 U22182 ( .A1(n10141), .A2(n24793), .ZN(n17106) );
  AOI22_X2 U22184 ( .A1(n38582), .A2(n36920), .B1(n7261), .B2(n5888), .ZN(
        n14874) );
  INV_X2 U22185 ( .I(n24579), .ZN(n38582) );
  NAND2_X2 U22190 ( .A1(n5137), .A2(n32091), .ZN(n24579) );
  NAND2_X2 U22191 ( .A1(n30173), .A2(n30172), .ZN(n4368) );
  NAND2_X2 U22192 ( .A1(n5139), .A2(n5138), .ZN(n18788) );
  NAND2_X2 U22195 ( .A1(n38583), .A2(n18915), .ZN(n23884) );
  OAI21_X2 U22206 ( .A1(n38499), .A2(n17521), .B(n36212), .ZN(n38583) );
  NOR2_X1 U22211 ( .A1(n21269), .A2(n33368), .ZN(n38864) );
  INV_X2 U22213 ( .I(n12924), .ZN(n33368) );
  XOR2_X1 U22215 ( .A1(n8888), .A2(n35142), .Z(n12924) );
  XOR2_X1 U22218 ( .A1(n26483), .A2(n12683), .Z(n38585) );
  INV_X2 U22222 ( .I(n38586), .ZN(n12049) );
  XNOR2_X1 U22228 ( .A1(n9768), .A2(n12039), .ZN(n38586) );
  XOR2_X1 U22229 ( .A1(n1065), .A2(n15617), .Z(n29056) );
  NAND2_X2 U22236 ( .A1(n13962), .A2(n13965), .ZN(n15617) );
  XOR2_X1 U22237 ( .A1(n22424), .A2(n22425), .Z(n22943) );
  XOR2_X1 U22238 ( .A1(n17838), .A2(n17839), .Z(n11622) );
  OAI21_X2 U22240 ( .A1(n31926), .A2(n31925), .B(n38587), .ZN(n7106) );
  XOR2_X1 U22243 ( .A1(n38588), .A2(n19825), .Z(Ciphertext[32]) );
  AOI22_X1 U22247 ( .A1(n13274), .A2(n15958), .B1(n13273), .B2(n13803), .ZN(
        n38588) );
  NOR2_X2 U22249 ( .A1(n38589), .A2(n29350), .ZN(n9839) );
  OAI22_X2 U22251 ( .A1(n4790), .A2(n5334), .B1(n5336), .B2(n1401), .ZN(n38589) );
  XOR2_X1 U22254 ( .A1(n28837), .A2(n11922), .Z(n3081) );
  XOR2_X1 U22256 ( .A1(n28925), .A2(n3082), .Z(n28837) );
  XOR2_X1 U22258 ( .A1(n29243), .A2(n38590), .Z(n37034) );
  XOR2_X1 U22260 ( .A1(n17243), .A2(n3665), .Z(n38590) );
  NAND3_X1 U22266 ( .A1(n1193), .A2(n5418), .A3(n31015), .ZN(n10361) );
  INV_X2 U22268 ( .I(n10980), .ZN(n38674) );
  XOR2_X1 U22279 ( .A1(n25324), .A2(n37110), .Z(n813) );
  NOR2_X1 U22281 ( .A1(n36422), .A2(n14439), .ZN(n22792) );
  NAND2_X1 U22284 ( .A1(n38592), .A2(n38591), .ZN(n18054) );
  NAND2_X2 U22286 ( .A1(n39361), .A2(n34220), .ZN(n10463) );
  NAND2_X2 U22293 ( .A1(n38593), .A2(n19109), .ZN(n29559) );
  NAND2_X1 U22296 ( .A1(n34804), .A2(n34806), .ZN(n38593) );
  OR2_X1 U22297 ( .A1(n38358), .A2(n25660), .Z(n25576) );
  NOR2_X1 U22301 ( .A1(n24608), .A2(n39704), .ZN(n7067) );
  NAND2_X2 U22309 ( .A1(n3794), .A2(n38596), .ZN(n11330) );
  INV_X1 U22315 ( .I(n34134), .ZN(n39021) );
  XNOR2_X1 U22318 ( .A1(n7076), .A2(n31289), .ZN(n34134) );
  INV_X2 U22319 ( .I(n38597), .ZN(n24404) );
  XOR2_X1 U22321 ( .A1(n13568), .A2(n3447), .Z(n3446) );
  XOR2_X1 U22322 ( .A1(n26197), .A2(n26225), .Z(n32839) );
  XOR2_X1 U22323 ( .A1(n15034), .A2(n38598), .Z(n15036) );
  XOR2_X1 U22324 ( .A1(n24641), .A2(n37231), .Z(n38598) );
  OAI21_X2 U22325 ( .A1(n38599), .A2(n1940), .B(n1939), .ZN(n1938) );
  NOR2_X1 U22347 ( .A1(n3690), .A2(n2502), .ZN(n38599) );
  AND2_X1 U22348 ( .A1(n22347), .A2(n22346), .Z(n10037) );
  NAND2_X2 U22351 ( .A1(n36753), .A2(n10630), .ZN(n22347) );
  INV_X2 U22353 ( .I(n32601), .ZN(n38600) );
  INV_X4 U22354 ( .I(n39663), .ZN(n2416) );
  XOR2_X1 U22366 ( .A1(n38602), .A2(n20257), .Z(n26921) );
  XOR2_X1 U22368 ( .A1(n20260), .A2(n32175), .Z(n38602) );
  XOR2_X1 U22371 ( .A1(n24039), .A2(n38603), .Z(n2168) );
  XOR2_X1 U22372 ( .A1(n36748), .A2(n36895), .Z(n38603) );
  XOR2_X1 U22373 ( .A1(n38988), .A2(n18491), .Z(n18525) );
  OR2_X1 U22374 ( .A1(n33483), .A2(n24192), .Z(n15258) );
  XOR2_X1 U22376 ( .A1(n15250), .A2(n7359), .Z(n33483) );
  AOI22_X2 U22381 ( .A1(n2520), .A2(n1890), .B1(n9201), .B2(n2519), .ZN(n2518)
         );
  XOR2_X1 U22383 ( .A1(n29158), .A2(n38606), .Z(n38605) );
  NAND2_X2 U22384 ( .A1(n28258), .A2(n27884), .ZN(n28171) );
  XOR2_X1 U22386 ( .A1(n27537), .A2(n34963), .Z(n27805) );
  NOR2_X2 U22391 ( .A1(n5769), .A2(n5770), .ZN(n34963) );
  XOR2_X1 U22393 ( .A1(n18785), .A2(n29104), .Z(n28603) );
  NAND3_X2 U22396 ( .A1(n28601), .A2(n34463), .A3(n34462), .ZN(n29104) );
  NAND2_X2 U22406 ( .A1(n27870), .A2(n19743), .ZN(n27871) );
  NAND2_X2 U22409 ( .A1(n14829), .A2(n14828), .ZN(n33307) );
  AOI21_X2 U22410 ( .A1(n21025), .A2(n16691), .B(n38607), .ZN(n21024) );
  NOR3_X2 U22413 ( .A1(n36814), .A2(n31924), .A3(n28299), .ZN(n38607) );
  NOR2_X2 U22414 ( .A1(n8090), .A2(n38608), .ZN(n11753) );
  INV_X2 U22416 ( .I(n26157), .ZN(n26394) );
  XOR2_X1 U22426 ( .A1(n38610), .A2(n39025), .Z(n33387) );
  NAND2_X1 U22428 ( .A1(n38408), .A2(n37088), .ZN(n31739) );
  AOI22_X2 U22431 ( .A1(n28513), .A2(n29702), .B1(n34793), .B2(n35858), .ZN(
        n29568) );
  XOR2_X1 U22435 ( .A1(n12865), .A2(n27480), .Z(n11237) );
  NAND2_X2 U22437 ( .A1(n5695), .A2(n16856), .ZN(n12865) );
  NOR2_X2 U22440 ( .A1(n38612), .A2(n556), .ZN(n27498) );
  AOI21_X2 U22442 ( .A1(n27205), .A2(n27206), .B(n27400), .ZN(n38612) );
  NAND2_X2 U22443 ( .A1(n38615), .A2(n38613), .ZN(n17745) );
  NAND2_X1 U22447 ( .A1(n38614), .A2(n23550), .ZN(n38613) );
  XOR2_X1 U22448 ( .A1(n24013), .A2(n38616), .Z(n39590) );
  XOR2_X1 U22455 ( .A1(n24012), .A2(n35640), .Z(n38616) );
  XOR2_X1 U22457 ( .A1(n31565), .A2(n31863), .Z(n11233) );
  NAND2_X2 U22461 ( .A1(n8213), .A2(n8211), .ZN(n24076) );
  AOI22_X2 U22464 ( .A1(n33667), .A2(n23505), .B1(n8214), .B2(n8190), .ZN(
        n8213) );
  INV_X2 U22468 ( .I(n21461), .ZN(n38617) );
  NOR2_X2 U22473 ( .A1(n38617), .A2(n21869), .ZN(n32114) );
  NAND2_X2 U22474 ( .A1(n56), .A2(n38621), .ZN(n34609) );
  NAND3_X2 U22476 ( .A1(n12704), .A2(n12705), .A3(n1115), .ZN(n38621) );
  XOR2_X1 U22478 ( .A1(n19632), .A2(n38622), .Z(n26931) );
  XOR2_X1 U22479 ( .A1(n26558), .A2(n26557), .Z(n38622) );
  NOR2_X2 U22481 ( .A1(n5311), .A2(n27407), .ZN(n5059) );
  XOR2_X1 U22486 ( .A1(n6066), .A2(n24959), .Z(n25257) );
  NOR2_X2 U22488 ( .A1(n38867), .A2(n30413), .ZN(n24959) );
  XOR2_X1 U22490 ( .A1(n23396), .A2(n37148), .Z(n7734) );
  XOR2_X1 U22492 ( .A1(n24023), .A2(n23764), .Z(n23396) );
  NAND2_X2 U22493 ( .A1(n34895), .A2(n11170), .ZN(n24712) );
  AOI21_X2 U22496 ( .A1(n1453), .A2(n2262), .B(n12443), .ZN(n4151) );
  XOR2_X1 U22497 ( .A1(n29167), .A2(n6719), .Z(n28909) );
  NOR2_X2 U22501 ( .A1(n35823), .A2(n16036), .ZN(n6719) );
  INV_X2 U22502 ( .I(n38627), .ZN(n35792) );
  NAND3_X2 U22503 ( .A1(n23160), .A2(n35684), .A3(n10436), .ZN(n38627) );
  NAND2_X2 U22505 ( .A1(n14794), .A2(n38628), .ZN(n378) );
  XOR2_X1 U22509 ( .A1(n27464), .A2(n27492), .Z(n27847) );
  NOR2_X2 U22511 ( .A1(n19803), .A2(n19802), .ZN(n27464) );
  NAND2_X2 U22513 ( .A1(n16535), .A2(n10209), .ZN(n17996) );
  NAND2_X2 U22516 ( .A1(n31425), .A2(n12556), .ZN(n4529) );
  OR2_X1 U22523 ( .A1(n6533), .A2(n36509), .Z(n27237) );
  NAND2_X2 U22524 ( .A1(n7800), .A2(n24240), .ZN(n24243) );
  XOR2_X1 U22527 ( .A1(n4086), .A2(n4085), .Z(n8452) );
  AND2_X1 U22528 ( .A1(n24898), .A2(n39505), .Z(n5030) );
  AOI22_X2 U22535 ( .A1(n10069), .A2(n20058), .B1(n14156), .B2(n6215), .ZN(
        n6214) );
  OAI21_X2 U22542 ( .A1(n33995), .A2(n38075), .B(n3903), .ZN(n6505) );
  NAND2_X1 U22546 ( .A1(n3373), .A2(n19098), .ZN(n3372) );
  OAI22_X2 U22548 ( .A1(n1079), .A2(n38638), .B1(n8453), .B2(n10946), .ZN(
        n15465) );
  XOR2_X1 U22550 ( .A1(n12971), .A2(n33334), .Z(n38639) );
  AOI22_X2 U22563 ( .A1(n22138), .A2(n22246), .B1(n22139), .B2(n35290), .ZN(
        n38640) );
  NAND2_X1 U22565 ( .A1(n19514), .A2(n25420), .ZN(n38642) );
  NAND2_X1 U22567 ( .A1(n38644), .A2(n34005), .ZN(n38643) );
  INV_X2 U22569 ( .I(n19821), .ZN(n38644) );
  NAND2_X2 U22570 ( .A1(n34683), .A2(n38645), .ZN(n22228) );
  AOI21_X2 U22573 ( .A1(n38647), .A2(n1351), .B(n38646), .ZN(n38645) );
  NOR2_X1 U22574 ( .A1(n17160), .A2(n1351), .ZN(n38646) );
  INV_X1 U22575 ( .I(n13348), .ZN(n38647) );
  XOR2_X1 U22579 ( .A1(n31352), .A2(n22605), .Z(n2030) );
  XOR2_X1 U22587 ( .A1(n38648), .A2(n11755), .Z(n36880) );
  NAND2_X2 U22588 ( .A1(n38780), .A2(n10949), .ZN(n11755) );
  XOR2_X1 U22602 ( .A1(n38649), .A2(n20674), .Z(n20677) );
  XOR2_X1 U22603 ( .A1(n21157), .A2(n10258), .Z(n38649) );
  NOR2_X2 U22604 ( .A1(n38650), .A2(n15969), .ZN(n23929) );
  INV_X2 U22612 ( .I(n33786), .ZN(n39300) );
  NAND2_X2 U22613 ( .A1(n13406), .A2(n13407), .ZN(n33786) );
  XOR2_X1 U22615 ( .A1(n1557), .A2(n25079), .Z(n25148) );
  NAND2_X1 U22617 ( .A1(n23342), .A2(n23343), .ZN(n23344) );
  NAND2_X2 U22620 ( .A1(n33894), .A2(n23624), .ZN(n23342) );
  XOR2_X1 U22621 ( .A1(n23982), .A2(n5290), .Z(n36079) );
  OR2_X1 U22622 ( .A1(n39265), .A2(n24868), .Z(n32268) );
  NAND2_X2 U22623 ( .A1(n4452), .A2(n4453), .ZN(n26098) );
  NAND2_X2 U22624 ( .A1(n20642), .A2(n28297), .ZN(n16096) );
  NAND3_X2 U22630 ( .A1(n20111), .A2(n27317), .A3(n27316), .ZN(n7549) );
  OAI21_X2 U22634 ( .A1(n8993), .A2(n38868), .B(n37828), .ZN(n32146) );
  XOR2_X1 U22635 ( .A1(n38654), .A2(n11210), .Z(n34218) );
  XOR2_X1 U22642 ( .A1(n27841), .A2(n27740), .Z(n38654) );
  AOI22_X2 U22644 ( .A1(n6314), .A2(n29453), .B1(n39647), .B2(n29378), .ZN(
        n39060) );
  XOR2_X1 U22648 ( .A1(n18930), .A2(n18705), .Z(n19478) );
  INV_X1 U22661 ( .I(n38843), .ZN(n17894) );
  OR2_X1 U22665 ( .A1(n38843), .A2(n34010), .Z(n17038) );
  XOR2_X1 U22666 ( .A1(n3320), .A2(n38655), .Z(n3885) );
  XOR2_X1 U22671 ( .A1(n33310), .A2(n38261), .Z(n38655) );
  NAND2_X2 U22672 ( .A1(n3964), .A2(n3966), .ZN(n29085) );
  NAND2_X2 U22676 ( .A1(n988), .A2(n10642), .ZN(n28276) );
  AOI21_X2 U22677 ( .A1(n14543), .A2(n28808), .B(n38657), .ZN(n16658) );
  XOR2_X1 U22680 ( .A1(n12401), .A2(n12400), .Z(n12399) );
  NOR2_X2 U22683 ( .A1(n27371), .A2(n31672), .ZN(n12374) );
  NAND2_X2 U22685 ( .A1(n27372), .A2(n27267), .ZN(n27371) );
  XOR2_X1 U22690 ( .A1(n24938), .A2(n25176), .Z(n25246) );
  NOR2_X2 U22694 ( .A1(n24815), .A2(n7321), .ZN(n25176) );
  XOR2_X1 U22695 ( .A1(n5731), .A2(n36339), .Z(n30465) );
  NAND2_X1 U22698 ( .A1(n39013), .A2(n36560), .ZN(n39131) );
  XOR2_X1 U22700 ( .A1(n10782), .A2(n27793), .Z(n8958) );
  XOR2_X1 U22702 ( .A1(n3163), .A2(n4734), .Z(n38659) );
  XOR2_X1 U22704 ( .A1(n28855), .A2(n28545), .Z(n12455) );
  XOR2_X1 U22707 ( .A1(n29067), .A2(n29819), .Z(n28855) );
  NAND2_X2 U22709 ( .A1(n10807), .A2(n37172), .ZN(n25827) );
  INV_X2 U22710 ( .I(n3496), .ZN(n33894) );
  NAND3_X2 U22715 ( .A1(n32909), .A2(n10437), .A3(n10438), .ZN(n3496) );
  XOR2_X1 U22719 ( .A1(n38660), .A2(n2159), .Z(n31107) );
  XOR2_X1 U22720 ( .A1(n3559), .A2(n27791), .Z(n38660) );
  XOR2_X1 U22721 ( .A1(n4412), .A2(n33039), .Z(n4409) );
  NAND2_X1 U22722 ( .A1(n23272), .A2(n18199), .ZN(n18198) );
  OR2_X1 U22726 ( .A1(n29199), .A2(n11348), .Z(n35869) );
  AOI22_X2 U22727 ( .A1(n25538), .A2(n13461), .B1(n39327), .B2(n12908), .ZN(
        n38663) );
  XOR2_X1 U22731 ( .A1(n38664), .A2(n18270), .Z(Ciphertext[16]) );
  NAND4_X2 U22733 ( .A1(n29233), .A2(n36232), .A3(n39306), .A4(n29234), .ZN(
        n38664) );
  XOR2_X1 U22738 ( .A1(n37129), .A2(n7549), .Z(n27817) );
  NOR2_X2 U22742 ( .A1(n14614), .A2(n6648), .ZN(n20112) );
  NOR2_X2 U22748 ( .A1(n32131), .A2(n7706), .ZN(n14614) );
  NAND3_X1 U22749 ( .A1(n5282), .A2(n24683), .A3(n13300), .ZN(n17893) );
  NAND2_X2 U22755 ( .A1(n8925), .A2(n33493), .ZN(n5282) );
  NAND3_X1 U22756 ( .A1(n20174), .A2(n20590), .A3(n19966), .ZN(n2356) );
  OR2_X1 U22757 ( .A1(n6515), .A2(n33599), .Z(n35150) );
  OAI21_X2 U22758 ( .A1(n38667), .A2(n34524), .B(n1020), .ZN(n3380) );
  NOR2_X2 U22759 ( .A1(n1104), .A2(n26055), .ZN(n38667) );
  XOR2_X1 U22762 ( .A1(n22509), .A2(n22510), .Z(n22661) );
  NAND3_X2 U22766 ( .A1(n24121), .A2(n17066), .A3(n35253), .ZN(n34693) );
  XOR2_X1 U22770 ( .A1(n6277), .A2(n38670), .Z(n24196) );
  XOR2_X1 U22772 ( .A1(n23711), .A2(n23865), .Z(n38670) );
  XOR2_X1 U22774 ( .A1(n9577), .A2(n7371), .Z(n26808) );
  XOR2_X1 U22778 ( .A1(n27613), .A2(n27614), .Z(n28157) );
  NAND2_X2 U22780 ( .A1(n24345), .A2(n5953), .ZN(n39413) );
  XOR2_X1 U22786 ( .A1(n26435), .A2(n26387), .Z(n26527) );
  NOR2_X2 U22788 ( .A1(n16525), .A2(n25821), .ZN(n26435) );
  AOI22_X2 U22790 ( .A1(n23297), .A2(n23462), .B1(n23298), .B2(n23460), .ZN(
        n23301) );
  NAND2_X1 U22801 ( .A1(n38727), .A2(n28546), .ZN(n19043) );
  AOI21_X2 U22802 ( .A1(n9375), .A2(n9380), .B(n38671), .ZN(n31883) );
  INV_X2 U22805 ( .I(n25532), .ZN(n38671) );
  NAND2_X2 U22809 ( .A1(n15085), .A2(n33440), .ZN(n25532) );
  XOR2_X1 U22812 ( .A1(n4081), .A2(n39119), .Z(n26651) );
  OAI22_X2 U22815 ( .A1(n4455), .A2(n4454), .B1(n32722), .B2(n25514), .ZN(
        n4453) );
  AOI22_X2 U22816 ( .A1(n30397), .A2(n21900), .B1(n21901), .B2(n275), .ZN(
        n15468) );
  NOR2_X2 U22817 ( .A1(n21840), .A2(n1348), .ZN(n21901) );
  BUF_X2 U22818 ( .I(n36371), .Z(n38673) );
  NAND2_X1 U22820 ( .A1(n29208), .A2(n15535), .ZN(n29205) );
  AOI21_X2 U22828 ( .A1(n38676), .A2(n23100), .B(n11659), .ZN(n13087) );
  NOR2_X2 U22830 ( .A1(n15330), .A2(n33082), .ZN(n38676) );
  NAND2_X2 U22835 ( .A1(n38677), .A2(n11260), .ZN(n24817) );
  NAND2_X1 U22844 ( .A1(n10219), .A2(n36872), .ZN(n38677) );
  XOR2_X1 U22848 ( .A1(n29088), .A2(n2392), .Z(n10185) );
  AND2_X1 U22849 ( .A1(n18827), .A2(n35648), .Z(n39806) );
  NAND3_X2 U22853 ( .A1(n5864), .A2(n5863), .A3(n38678), .ZN(n7023) );
  XOR2_X1 U22857 ( .A1(n14039), .A2(n38679), .Z(n30925) );
  NAND2_X2 U22868 ( .A1(n12046), .A2(n12045), .ZN(n14039) );
  AOI22_X2 U22869 ( .A1(n27344), .A2(n1225), .B1(n27342), .B2(n27343), .ZN(
        n27345) );
  OAI21_X2 U22878 ( .A1(n1029), .A2(n9825), .B(n17101), .ZN(n10654) );
  NAND2_X2 U22880 ( .A1(n24108), .A2(n24109), .ZN(n9825) );
  CLKBUF_X4 U22884 ( .I(n966), .Z(n39018) );
  OR2_X2 U22890 ( .A1(n2416), .A2(n39021), .Z(n36345) );
  NAND2_X2 U22896 ( .A1(n9835), .A2(n23475), .ZN(n19633) );
  NAND2_X1 U22900 ( .A1(n38223), .A2(n3937), .ZN(n9337) );
  XOR2_X1 U22908 ( .A1(n28967), .A2(n10328), .Z(n36746) );
  XOR2_X1 U22911 ( .A1(n26531), .A2(n32253), .Z(n12411) );
  OAI21_X2 U22919 ( .A1(n3244), .A2(n7699), .B(n39625), .ZN(n26531) );
  XOR2_X1 U22920 ( .A1(n36804), .A2(n38680), .Z(n12298) );
  XOR2_X1 U22930 ( .A1(n9184), .A2(n6688), .Z(n38680) );
  XOR2_X1 U22934 ( .A1(n18327), .A2(n38682), .Z(n39263) );
  XOR2_X1 U22945 ( .A1(n24702), .A2(n37121), .Z(n38682) );
  NAND2_X1 U22954 ( .A1(n38644), .A2(n11616), .ZN(n38683) );
  NAND2_X1 U22956 ( .A1(n1235), .A2(n38684), .ZN(n32725) );
  NAND2_X2 U22957 ( .A1(n12392), .A2(n23111), .ZN(n3119) );
  AOI21_X2 U22959 ( .A1(n38686), .A2(n38685), .B(n1115), .ZN(n34272) );
  INV_X2 U22963 ( .I(n34010), .ZN(n38685) );
  BUF_X2 U22971 ( .I(n35431), .Z(n38687) );
  NAND2_X2 U22972 ( .A1(n38689), .A2(n38688), .ZN(n26648) );
  XOR2_X1 U22973 ( .A1(n26262), .A2(n35212), .Z(n844) );
  OAI21_X2 U22976 ( .A1(n16239), .A2(n7888), .B(n25807), .ZN(n26262) );
  OAI21_X2 U22977 ( .A1(n16182), .A2(n6176), .B(n38691), .ZN(n15353) );
  NAND2_X2 U22983 ( .A1(n4160), .A2(n4161), .ZN(n6176) );
  NAND2_X2 U22984 ( .A1(n13233), .A2(n10346), .ZN(n29630) );
  XOR2_X1 U22985 ( .A1(n9894), .A2(n38692), .Z(n2052) );
  XOR2_X1 U22986 ( .A1(n11938), .A2(n36067), .Z(n38692) );
  AND2_X1 U22992 ( .A1(n36509), .A2(n36523), .Z(n32950) );
  INV_X2 U22994 ( .I(n18175), .ZN(n23757) );
  NAND2_X2 U23000 ( .A1(n38693), .A2(n36091), .ZN(n18175) );
  OR2_X1 U23009 ( .A1(n20818), .A2(n18389), .Z(n38693) );
  XOR2_X1 U23014 ( .A1(n17360), .A2(n17361), .Z(n36970) );
  NOR2_X2 U23015 ( .A1(n8641), .A2(n8640), .ZN(n39442) );
  NOR2_X2 U23022 ( .A1(n13308), .A2(n24301), .ZN(n38749) );
  AOI21_X2 U23028 ( .A1(n29781), .A2(n1402), .B(n481), .ZN(n2017) );
  NAND3_X1 U23029 ( .A1(n23518), .A2(n39001), .A3(n6373), .ZN(n38806) );
  AOI22_X2 U23031 ( .A1(n38800), .A2(n35288), .B1(n17778), .B2(n7902), .ZN(
        n39001) );
  OR2_X1 U23035 ( .A1(n20566), .A2(n29241), .Z(n38823) );
  AOI22_X2 U23037 ( .A1(n35369), .A2(n1186), .B1(n20621), .B2(n7486), .ZN(
        n20314) );
  BUF_X2 U23038 ( .I(n6056), .Z(n38694) );
  AND2_X1 U23039 ( .A1(n37188), .A2(n6136), .Z(n39530) );
  NAND2_X2 U23044 ( .A1(n6390), .A2(n6180), .ZN(n7961) );
  INV_X2 U23045 ( .I(n27314), .ZN(n27409) );
  OAI22_X2 U23046 ( .A1(n12714), .A2(n12713), .B1(n26766), .B2(n12078), .ZN(
        n27314) );
  NAND2_X2 U23048 ( .A1(n8253), .A2(n32191), .ZN(n27084) );
  NAND2_X2 U23050 ( .A1(n33098), .A2(n33097), .ZN(n8253) );
  AOI21_X2 U23059 ( .A1(n24155), .A2(n10220), .B(n2595), .ZN(n38695) );
  NAND2_X1 U23060 ( .A1(n25486), .A2(n18207), .ZN(n25305) );
  AOI22_X2 U23062 ( .A1(n38696), .A2(n24655), .B1(n24507), .B2(n33409), .ZN(
        n4729) );
  NOR2_X2 U23065 ( .A1(n19679), .A2(n37355), .ZN(n38696) );
  AND2_X1 U23066 ( .A1(n5383), .A2(n39435), .Z(n39473) );
  XOR2_X1 U23081 ( .A1(n38697), .A2(n19805), .Z(Ciphertext[76]) );
  NAND2_X2 U23085 ( .A1(n38698), .A2(n35762), .ZN(n29616) );
  XOR2_X1 U23089 ( .A1(n22659), .A2(n19128), .Z(n19127) );
  XNOR2_X1 U23094 ( .A1(n22702), .A2(n644), .ZN(n39039) );
  NAND3_X1 U23109 ( .A1(n9987), .A2(n5819), .A3(n21961), .ZN(n38699) );
  XOR2_X1 U23111 ( .A1(n31492), .A2(n39654), .Z(n11810) );
  NOR2_X1 U23113 ( .A1(n38701), .A2(n38700), .ZN(n39007) );
  INV_X1 U23116 ( .I(n5819), .ZN(n38701) );
  INV_X2 U23122 ( .I(n19142), .ZN(n38702) );
  NAND2_X2 U23130 ( .A1(n15811), .A2(n15814), .ZN(n17499) );
  INV_X1 U23132 ( .I(n5340), .ZN(n8703) );
  NOR2_X2 U23134 ( .A1(n12784), .A2(n28282), .ZN(n28167) );
  OR2_X1 U23138 ( .A1(n14212), .A2(n10986), .Z(n12552) );
  XOR2_X1 U23141 ( .A1(n27785), .A2(n20721), .Z(n32807) );
  OAI21_X1 U23144 ( .A1(n27282), .A2(n1227), .B(n38705), .ZN(n3718) );
  NAND2_X1 U23145 ( .A1(n27282), .A2(n3313), .ZN(n38705) );
  XOR2_X1 U23148 ( .A1(n3731), .A2(n18887), .Z(n38706) );
  XOR2_X1 U23153 ( .A1(n311), .A2(n10014), .Z(n11586) );
  NAND2_X2 U23155 ( .A1(n32883), .A2(n2182), .ZN(n9968) );
  NAND2_X2 U23158 ( .A1(n38708), .A2(n38707), .ZN(n29189) );
  NAND2_X2 U23165 ( .A1(n29187), .A2(n3631), .ZN(n38707) );
  NAND2_X2 U23181 ( .A1(n29188), .A2(n38709), .ZN(n38708) );
  NOR2_X1 U23182 ( .A1(n24091), .A2(n37066), .ZN(n39191) );
  XOR2_X1 U23184 ( .A1(n38820), .A2(n29816), .Z(n38710) );
  INV_X4 U23187 ( .I(n7445), .ZN(n24646) );
  NAND2_X2 U23189 ( .A1(n28087), .A2(n28086), .ZN(n33047) );
  XOR2_X1 U23193 ( .A1(n24997), .A2(n2653), .Z(n25210) );
  NAND2_X2 U23201 ( .A1(n16668), .A2(n14681), .ZN(n24997) );
  NAND2_X2 U23204 ( .A1(n15670), .A2(n26944), .ZN(n38715) );
  NAND2_X1 U23205 ( .A1(n19367), .A2(n12162), .ZN(n38716) );
  OAI21_X2 U23209 ( .A1(n36295), .A2(n13516), .B(n24616), .ZN(n34564) );
  OAI21_X2 U23210 ( .A1(n2331), .A2(n14278), .B(n38717), .ZN(n16017) );
  OAI22_X2 U23212 ( .A1(n22246), .A2(n38718), .B1(n35290), .B2(n9265), .ZN(
        n22036) );
  INV_X2 U23213 ( .I(n33713), .ZN(n38719) );
  NAND2_X2 U23215 ( .A1(n38721), .A2(n38720), .ZN(n23778) );
  NAND2_X1 U23226 ( .A1(n19633), .A2(n12011), .ZN(n38720) );
  OAI21_X2 U23227 ( .A1(n12008), .A2(n12009), .B(n34823), .ZN(n38721) );
  XOR2_X1 U23231 ( .A1(n29093), .A2(n1411), .Z(n28984) );
  INV_X2 U23234 ( .I(n31396), .ZN(n1411) );
  NOR2_X2 U23237 ( .A1(n34266), .A2(n18103), .ZN(n31396) );
  OAI21_X2 U23239 ( .A1(n2062), .A2(n17075), .B(n38722), .ZN(n39030) );
  AOI22_X2 U23240 ( .A1(n33113), .A2(n33115), .B1(n1984), .B2(n33114), .ZN(
        n38722) );
  XOR2_X1 U23249 ( .A1(n38723), .A2(n16975), .Z(n29768) );
  XOR2_X1 U23253 ( .A1(n20006), .A2(n489), .Z(n38723) );
  BUF_X2 U23256 ( .I(n34757), .Z(n38725) );
  INV_X4 U23259 ( .I(n24896), .ZN(n38782) );
  OR2_X1 U23269 ( .A1(n23489), .A2(n23602), .Z(n30631) );
  NOR2_X1 U23270 ( .A1(n5598), .A2(n21914), .ZN(n20832) );
  AND2_X1 U23272 ( .A1(n33316), .A2(n23444), .Z(n38893) );
  NAND2_X2 U23276 ( .A1(n38729), .A2(n38728), .ZN(n30372) );
  NAND2_X2 U23277 ( .A1(n38731), .A2(n38730), .ZN(n38729) );
  INV_X2 U23285 ( .I(n25542), .ZN(n38731) );
  BUF_X2 U23286 ( .I(n39820), .Z(n38732) );
  NAND3_X2 U23289 ( .A1(n38733), .A2(n36098), .A3(n36097), .ZN(n9310) );
  OAI21_X2 U23301 ( .A1(n37156), .A2(n7511), .B(n26564), .ZN(n38733) );
  XOR2_X1 U23303 ( .A1(n12534), .A2(n19359), .Z(n25152) );
  NAND3_X2 U23309 ( .A1(n5123), .A2(n5122), .A3(n31455), .ZN(n12534) );
  XOR2_X1 U23311 ( .A1(n38735), .A2(n26584), .Z(n11374) );
  XOR2_X1 U23312 ( .A1(n26365), .A2(n12667), .Z(n38735) );
  OAI21_X2 U23314 ( .A1(n20584), .A2(n31966), .B(n11518), .ZN(n14448) );
  NAND2_X2 U23315 ( .A1(n10469), .A2(n10471), .ZN(n11970) );
  OAI21_X2 U23316 ( .A1(n34618), .A2(n34619), .B(n9872), .ZN(n38737) );
  XOR2_X1 U23319 ( .A1(n35089), .A2(n36211), .Z(n34876) );
  INV_X1 U23320 ( .I(n38739), .ZN(n8210) );
  OAI21_X2 U23322 ( .A1(n31234), .A2(n31235), .B(n30274), .ZN(n13306) );
  NAND2_X2 U23323 ( .A1(n18330), .A2(n18331), .ZN(n11342) );
  OAI21_X2 U23326 ( .A1(n26220), .A2(n1494), .B(n38740), .ZN(n6376) );
  NOR2_X2 U23327 ( .A1(n34224), .A2(n37103), .ZN(n38740) );
  XOR2_X1 U23328 ( .A1(n27475), .A2(n38741), .Z(n34491) );
  INV_X2 U23335 ( .I(n8874), .ZN(n38741) );
  XOR2_X1 U23340 ( .A1(n26278), .A2(n35214), .Z(n11399) );
  NAND3_X2 U23341 ( .A1(n13184), .A2(n13182), .A3(n36801), .ZN(n20576) );
  INV_X2 U23343 ( .I(n38743), .ZN(n17390) );
  NOR2_X2 U23347 ( .A1(n38745), .A2(n38744), .ZN(n36408) );
  NOR2_X2 U23357 ( .A1(n10654), .A2(n2341), .ZN(n38745) );
  BUF_X2 U23366 ( .I(n20391), .Z(n38746) );
  NOR2_X2 U23368 ( .A1(n33036), .A2(n38747), .ZN(n12393) );
  NAND2_X2 U23376 ( .A1(n20405), .A2(n34389), .ZN(n6045) );
  BUF_X2 U23377 ( .I(n23550), .Z(n38748) );
  NOR2_X2 U23378 ( .A1(n31601), .A2(n30097), .ZN(n30087) );
  AOI21_X2 U23381 ( .A1(n3527), .A2(n19476), .B(n6044), .ZN(n31601) );
  XOR2_X1 U23383 ( .A1(n38750), .A2(n15331), .Z(n4016) );
  XOR2_X1 U23386 ( .A1(n3386), .A2(n20719), .Z(n38750) );
  XOR2_X1 U23387 ( .A1(n5603), .A2(n39028), .Z(n34757) );
  INV_X2 U23395 ( .I(n38751), .ZN(n1984) );
  NAND2_X2 U23397 ( .A1(n2416), .A2(n37086), .ZN(n38751) );
  NAND2_X2 U23398 ( .A1(n34326), .A2(n20084), .ZN(n29071) );
  OR2_X1 U23399 ( .A1(n1448), .A2(n28079), .Z(n7219) );
  OAI21_X2 U23408 ( .A1(n19006), .A2(n38754), .B(n23259), .ZN(n23910) );
  XOR2_X1 U23411 ( .A1(n25186), .A2(n25118), .Z(n11102) );
  NAND2_X2 U23414 ( .A1(n819), .A2(n24210), .ZN(n25118) );
  NAND2_X2 U23419 ( .A1(n21662), .A2(n21951), .ZN(n20367) );
  NAND2_X2 U23421 ( .A1(n32113), .A2(n17991), .ZN(n17989) );
  AOI21_X2 U23423 ( .A1(n23201), .A2(n38756), .B(n22850), .ZN(n2413) );
  NOR2_X1 U23425 ( .A1(n2350), .A2(n36369), .ZN(n38756) );
  XOR2_X1 U23426 ( .A1(n4354), .A2(n4355), .Z(n4356) );
  INV_X1 U23427 ( .I(n33883), .ZN(n27727) );
  XNOR2_X1 U23437 ( .A1(n27683), .A2(n27858), .ZN(n33883) );
  XOR2_X1 U23439 ( .A1(n38758), .A2(n34933), .Z(n18790) );
  XOR2_X1 U23443 ( .A1(n23549), .A2(n21045), .Z(n38758) );
  XOR2_X1 U23445 ( .A1(n23979), .A2(n23715), .Z(n23563) );
  XOR2_X1 U23446 ( .A1(n7498), .A2(n9911), .Z(n12631) );
  XOR2_X1 U23447 ( .A1(n11600), .A2(n20268), .Z(n20704) );
  XOR2_X1 U23448 ( .A1(n38759), .A2(n28787), .Z(n20453) );
  XOR2_X1 U23449 ( .A1(n2431), .A2(n29128), .Z(n38759) );
  XOR2_X1 U23450 ( .A1(n22561), .A2(n3528), .Z(n22758) );
  NOR2_X2 U23451 ( .A1(n637), .A2(n12155), .ZN(n22561) );
  OR2_X1 U23461 ( .A1(n29737), .A2(n19348), .Z(n19369) );
  NAND2_X2 U23463 ( .A1(n16057), .A2(n16056), .ZN(n24023) );
  XOR2_X1 U23467 ( .A1(n23786), .A2(n15777), .Z(n20602) );
  XOR2_X1 U23469 ( .A1(n11098), .A2(n23880), .Z(n15777) );
  OAI21_X2 U23471 ( .A1(n20863), .A2(n38302), .B(n14699), .ZN(n13351) );
  NAND3_X2 U23473 ( .A1(n31331), .A2(n31332), .A3(n15953), .ZN(n14365) );
  NAND2_X2 U23474 ( .A1(n39255), .A2(n38761), .ZN(n8163) );
  AOI22_X2 U23477 ( .A1(n24771), .A2(n24770), .B1(n24769), .B2(n11846), .ZN(
        n38761) );
  XOR2_X1 U23478 ( .A1(n38763), .A2(n6324), .Z(n39043) );
  OAI21_X2 U23481 ( .A1(n38765), .A2(n38764), .B(n27911), .ZN(n18480) );
  NAND2_X1 U23486 ( .A1(n22316), .A2(n3863), .ZN(n22270) );
  NAND2_X2 U23487 ( .A1(n2403), .A2(n5417), .ZN(n22316) );
  NAND2_X2 U23488 ( .A1(n32727), .A2(n32728), .ZN(n38766) );
  NAND2_X2 U23494 ( .A1(n37014), .A2(n23456), .ZN(n17995) );
  NAND2_X2 U23497 ( .A1(n18819), .A2(n32397), .ZN(n37014) );
  NOR2_X2 U23499 ( .A1(n24336), .A2(n24232), .ZN(n12250) );
  INV_X4 U23501 ( .I(n38768), .ZN(n22222) );
  OR2_X2 U23505 ( .A1(n33051), .A2(n21679), .Z(n38768) );
  NAND2_X2 U23508 ( .A1(n38769), .A2(n8058), .ZN(n23337) );
  NAND2_X2 U23512 ( .A1(n22705), .A2(n22926), .ZN(n38769) );
  NOR2_X2 U23513 ( .A1(n37106), .A2(n6822), .ZN(n34303) );
  XOR2_X1 U23514 ( .A1(n38770), .A2(n3571), .Z(n23827) );
  AOI22_X2 U23517 ( .A1(n23496), .A2(n5357), .B1(n23592), .B2(n34603), .ZN(
        n23594) );
  NAND2_X2 U23522 ( .A1(n29426), .A2(n29424), .ZN(n6314) );
  NAND2_X1 U23523 ( .A1(n5500), .A2(n38771), .ZN(n39775) );
  NAND2_X1 U23524 ( .A1(n7992), .A2(n4736), .ZN(n38771) );
  AND2_X1 U23529 ( .A1(n11831), .A2(n28484), .Z(n3019) );
  AOI22_X2 U23535 ( .A1(n34112), .A2(n14081), .B1(n18058), .B2(n25502), .ZN(
        n35453) );
  INV_X2 U23538 ( .I(n38772), .ZN(n3488) );
  OR2_X2 U23539 ( .A1(n1454), .A2(n18689), .Z(n28175) );
  XOR2_X1 U23548 ( .A1(n3320), .A2(n6365), .Z(n32293) );
  NAND2_X2 U23550 ( .A1(n27392), .A2(n35895), .ZN(n27393) );
  AOI21_X2 U23555 ( .A1(n38773), .A2(n14435), .B(n12954), .ZN(n15535) );
  NAND2_X2 U23559 ( .A1(n27661), .A2(n27557), .ZN(n10801) );
  NAND3_X2 U23561 ( .A1(n36250), .A2(n27431), .A3(n10755), .ZN(n27661) );
  NAND2_X2 U23562 ( .A1(n7619), .A2(n6615), .ZN(n38776) );
  INV_X2 U23575 ( .I(n39268), .ZN(n38777) );
  NAND2_X2 U23576 ( .A1(n36521), .A2(n36520), .ZN(n7096) );
  NAND3_X2 U23590 ( .A1(n20217), .A2(n26817), .A3(n26626), .ZN(n27095) );
  OAI21_X2 U23592 ( .A1(n38811), .A2(n36821), .B(n38848), .ZN(n31797) );
  XOR2_X1 U23595 ( .A1(n6825), .A2(n18428), .Z(n32734) );
  XOR2_X1 U23599 ( .A1(n25104), .A2(n17184), .Z(n18428) );
  NAND2_X2 U23602 ( .A1(n38778), .A2(n30726), .ZN(n12485) );
  OR2_X1 U23603 ( .A1(n25412), .A2(n25307), .Z(n38779) );
  NOR2_X2 U23620 ( .A1(n28643), .A2(n14448), .ZN(n28732) );
  NAND2_X1 U23621 ( .A1(n34111), .A2(n31185), .ZN(n38780) );
  NOR2_X2 U23628 ( .A1(n23119), .A2(n1145), .ZN(n23120) );
  NAND2_X1 U23632 ( .A1(n5570), .A2(n921), .ZN(n38785) );
  XOR2_X1 U23641 ( .A1(n18180), .A2(n26438), .Z(n26155) );
  NAND2_X2 U23647 ( .A1(n38786), .A2(n6105), .ZN(n36579) );
  OAI21_X2 U23648 ( .A1(n7293), .A2(n2625), .B(n7292), .ZN(n38786) );
  INV_X2 U23653 ( .I(n27102), .ZN(n38787) );
  NAND2_X2 U23654 ( .A1(n19030), .A2(n38787), .ZN(n27038) );
  AOI21_X1 U23655 ( .A1(n5471), .A2(n18816), .B(n39110), .ZN(n4449) );
  XOR2_X1 U23656 ( .A1(n2527), .A2(n2524), .Z(n5717) );
  INV_X2 U23658 ( .I(n9020), .ZN(n24136) );
  INV_X2 U23662 ( .I(n19233), .ZN(n38886) );
  XOR2_X1 U23665 ( .A1(n36760), .A2(n36759), .Z(n19233) );
  OAI21_X2 U23666 ( .A1(n944), .A2(n27269), .B(n38788), .ZN(n27374) );
  OAI21_X2 U23667 ( .A1(n36224), .A2(n28281), .B(n15622), .ZN(n38854) );
  XOR2_X1 U23669 ( .A1(n26413), .A2(n26412), .Z(n7374) );
  XOR2_X1 U23670 ( .A1(n26290), .A2(n39662), .Z(n26413) );
  NAND2_X2 U23671 ( .A1(n20988), .A2(n34693), .ZN(n24812) );
  XOR2_X1 U23675 ( .A1(n10706), .A2(n5486), .Z(n38791) );
  AOI22_X2 U23681 ( .A1(n34822), .A2(n22288), .B1(n22286), .B2(n22287), .ZN(
        n9486) );
  XOR2_X1 U23685 ( .A1(n21108), .A2(n28775), .Z(n19047) );
  NOR2_X2 U23686 ( .A1(n17849), .A2(n35272), .ZN(n19157) );
  NAND2_X2 U23690 ( .A1(n29401), .A2(n29402), .ZN(n35272) );
  NAND2_X2 U23692 ( .A1(n27298), .A2(n7757), .ZN(n27070) );
  XOR2_X1 U23696 ( .A1(n7737), .A2(n17579), .Z(n31633) );
  XOR2_X1 U23703 ( .A1(n27841), .A2(n38793), .Z(n9039) );
  XOR2_X1 U23704 ( .A1(n33398), .A2(n31620), .Z(n38793) );
  OAI22_X2 U23708 ( .A1(n38795), .A2(n38794), .B1(n18115), .B2(n1118), .ZN(
        n15525) );
  OAI21_X1 U23709 ( .A1(n9016), .A2(n10712), .B(n36595), .ZN(n3083) );
  XOR2_X1 U23710 ( .A1(n26450), .A2(n31154), .Z(n38796) );
  INV_X2 U23714 ( .I(n19425), .ZN(n38797) );
  XOR2_X1 U23715 ( .A1(n35241), .A2(n11755), .Z(n27636) );
  OR2_X1 U23723 ( .A1(n12334), .A2(n13082), .Z(n28074) );
  INV_X1 U23726 ( .I(n15019), .ZN(n21949) );
  NAND2_X2 U23727 ( .A1(n2555), .A2(n2554), .ZN(n29612) );
  NOR3_X2 U23735 ( .A1(n38238), .A2(n38798), .A3(n34061), .ZN(n32444) );
  XOR2_X1 U23743 ( .A1(n16096), .A2(n38799), .Z(n7766) );
  NOR2_X1 U23744 ( .A1(n14408), .A2(n30942), .ZN(n15142) );
  NAND2_X2 U23747 ( .A1(n14408), .A2(n1006), .ZN(n26661) );
  XOR2_X1 U23749 ( .A1(n3474), .A2(n3471), .Z(n17378) );
  INV_X2 U23753 ( .I(n38801), .ZN(n34123) );
  OAI22_X2 U23757 ( .A1(n9331), .A2(n23608), .B1(n32246), .B2(n98), .ZN(n24030) );
  XOR2_X1 U23758 ( .A1(n38802), .A2(n29506), .Z(Ciphertext[54]) );
  INV_X4 U23771 ( .I(n9333), .ZN(n9733) );
  NAND2_X2 U23772 ( .A1(n38803), .A2(n16231), .ZN(n9970) );
  OAI21_X2 U23773 ( .A1(n16016), .A2(n5980), .B(n5979), .ZN(n38803) );
  NOR2_X2 U23775 ( .A1(n38807), .A2(n46), .ZN(n10015) );
  AOI21_X2 U23779 ( .A1(n11363), .A2(n16825), .B(n38728), .ZN(n38807) );
  XOR2_X1 U23780 ( .A1(n28763), .A2(n36545), .Z(n21162) );
  NAND3_X1 U23785 ( .A1(n39206), .A2(n5311), .A3(n7606), .ZN(n16517) );
  XOR2_X1 U23788 ( .A1(n38808), .A2(n36284), .Z(n39608) );
  XOR2_X1 U23789 ( .A1(n39685), .A2(n37236), .Z(n38808) );
  XOR2_X1 U23791 ( .A1(n5323), .A2(n9518), .Z(n11215) );
  OR2_X1 U23792 ( .A1(n2416), .A2(n10665), .Z(n31619) );
  INV_X2 U23795 ( .I(n29439), .ZN(n1392) );
  AOI22_X1 U23796 ( .A1(n7154), .A2(n38848), .B1(n31986), .B2(n24792), .ZN(
        n9008) );
  XOR2_X1 U23799 ( .A1(n25253), .A2(n38809), .Z(n38815) );
  XOR2_X1 U23800 ( .A1(n7250), .A2(n25104), .Z(n25253) );
  INV_X2 U23801 ( .I(n38810), .ZN(n15549) );
  AOI21_X2 U23804 ( .A1(n26950), .A2(n13056), .B(n1236), .ZN(n38810) );
  OAI21_X2 U23809 ( .A1(n32640), .A2(n17897), .B(n20996), .ZN(n17896) );
  NOR2_X2 U23810 ( .A1(n19901), .A2(n37477), .ZN(n38811) );
  XOR2_X1 U23819 ( .A1(n35590), .A2(n39136), .Z(n11311) );
  NAND2_X2 U23823 ( .A1(n32282), .A2(n21959), .ZN(n39136) );
  XOR2_X1 U23825 ( .A1(n25251), .A2(n13763), .Z(n38814) );
  NOR2_X2 U23832 ( .A1(n26788), .A2(n1234), .ZN(n2362) );
  OAI21_X2 U23838 ( .A1(n19972), .A2(n1234), .B(n26909), .ZN(n26788) );
  OAI21_X2 U23844 ( .A1(n24429), .A2(n10815), .B(n38817), .ZN(n39253) );
  OAI21_X2 U23847 ( .A1(n18466), .A2(n14478), .B(n24373), .ZN(n38817) );
  NAND2_X2 U23849 ( .A1(n16224), .A2(n30047), .ZN(n11111) );
  NOR2_X2 U23850 ( .A1(n26682), .A2(n30500), .ZN(n32984) );
  OAI22_X2 U23851 ( .A1(n38819), .A2(n30550), .B1(n6715), .B2(n38404), .ZN(
        n35250) );
  AOI21_X2 U23856 ( .A1(n16141), .A2(n6715), .B(n10220), .ZN(n38819) );
  XOR2_X1 U23860 ( .A1(n2036), .A2(n38181), .Z(n38820) );
  NAND2_X2 U23863 ( .A1(n36016), .A2(n38821), .ZN(n7769) );
  AOI21_X2 U23865 ( .A1(n38823), .A2(n38822), .B(n1061), .ZN(n9869) );
  AOI21_X2 U23867 ( .A1(n3988), .A2(n28568), .B(n38826), .ZN(n19571) );
  NAND2_X2 U23868 ( .A1(n36124), .A2(n13378), .ZN(n38826) );
  XOR2_X1 U23876 ( .A1(n17342), .A2(n19825), .Z(n5610) );
  AOI22_X2 U23880 ( .A1(n17309), .A2(n32385), .B1(n11980), .B2(n38694), .ZN(
        n17342) );
  NAND3_X2 U23885 ( .A1(n27978), .A2(n27976), .A3(n37035), .ZN(n28616) );
  XOR2_X1 U23889 ( .A1(n12976), .A2(n38827), .Z(n24431) );
  XOR2_X1 U23891 ( .A1(n12798), .A2(n31466), .Z(n38827) );
  NAND2_X2 U23893 ( .A1(n38828), .A2(n17665), .ZN(n3840) );
  NAND3_X1 U23894 ( .A1(n12333), .A2(n9592), .A3(n35999), .ZN(n38828) );
  NOR2_X2 U23899 ( .A1(n20802), .A2(n25746), .ZN(n26026) );
  XOR2_X1 U23900 ( .A1(n542), .A2(n34391), .Z(n5993) );
  OAI21_X2 U23901 ( .A1(n35549), .A2(n35548), .B(n32983), .ZN(n542) );
  NAND3_X2 U23902 ( .A1(n11286), .A2(n34416), .A3(n11776), .ZN(n23903) );
  NAND3_X2 U23905 ( .A1(n38831), .A2(n36957), .A3(n5172), .ZN(n36509) );
  NAND3_X2 U23911 ( .A1(n18945), .A2(n34847), .A3(n18944), .ZN(n39772) );
  XOR2_X1 U23912 ( .A1(n1660), .A2(n22656), .Z(n13174) );
  NAND2_X2 U23914 ( .A1(n18124), .A2(n10366), .ZN(n31620) );
  AOI22_X2 U23916 ( .A1(n38833), .A2(n22326), .B1(n22249), .B2(n31383), .ZN(
        n13161) );
  INV_X2 U23919 ( .I(n13163), .ZN(n38833) );
  NOR2_X2 U23920 ( .A1(n30722), .A2(n37131), .ZN(n26744) );
  XOR2_X1 U23926 ( .A1(n28896), .A2(n28972), .Z(n16336) );
  BUF_X2 U23929 ( .I(n30232), .Z(n38834) );
  NAND2_X2 U23947 ( .A1(n33703), .A2(n36810), .ZN(n23400) );
  OAI21_X2 U23949 ( .A1(n7629), .A2(n7630), .B(n16058), .ZN(n24065) );
  BUF_X2 U23951 ( .I(n39030), .Z(n38835) );
  XOR2_X1 U23952 ( .A1(n12145), .A2(n26150), .Z(n7102) );
  INV_X2 U23956 ( .I(n22659), .ZN(n1669) );
  XNOR2_X1 U23967 ( .A1(Plaintext[93]), .A2(Key[93]), .ZN(n33147) );
  AOI21_X2 U23973 ( .A1(n2644), .A2(n21944), .B(n38836), .ZN(n4342) );
  NOR2_X2 U23982 ( .A1(n38837), .A2(n4982), .ZN(n5439) );
  INV_X2 U23990 ( .I(n22729), .ZN(n22628) );
  XOR2_X1 U23992 ( .A1(n22729), .A2(n38838), .Z(n509) );
  NOR2_X2 U23993 ( .A1(n32551), .A2(n20239), .ZN(n22729) );
  INV_X2 U23994 ( .I(n20352), .ZN(n38838) );
  NAND2_X1 U23995 ( .A1(n38840), .A2(n29210), .ZN(n29102) );
  NAND2_X1 U23998 ( .A1(n19765), .A2(n35870), .ZN(n38840) );
  XOR2_X1 U24002 ( .A1(n19571), .A2(n29254), .Z(n29094) );
  NOR2_X2 U24004 ( .A1(n19191), .A2(n34669), .ZN(n34371) );
  XOR2_X1 U24007 ( .A1(n8313), .A2(n17852), .Z(n18229) );
  NAND2_X2 U24010 ( .A1(n36535), .A2(n38841), .ZN(n6282) );
  NAND2_X2 U24011 ( .A1(n5928), .A2(n31424), .ZN(n29142) );
  XOR2_X1 U24012 ( .A1(n31599), .A2(n38021), .Z(n2476) );
  XOR2_X1 U24016 ( .A1(n38842), .A2(n1978), .Z(n11297) );
  XOR2_X1 U24017 ( .A1(n3157), .A2(n36529), .Z(n28117) );
  XOR2_X1 U24019 ( .A1(n33690), .A2(n3258), .Z(n36529) );
  NOR2_X2 U24021 ( .A1(n15159), .A2(n830), .ZN(n38843) );
  XOR2_X1 U24027 ( .A1(n38845), .A2(n37261), .Z(Ciphertext[110]) );
  OAI22_X1 U24030 ( .A1(n32466), .A2(n32467), .B1(n13606), .B2(n29812), .ZN(
        n38845) );
  OR2_X1 U24038 ( .A1(n37061), .A2(n33368), .Z(n20370) );
  XOR2_X1 U24045 ( .A1(n23952), .A2(n24002), .Z(n14220) );
  XOR2_X1 U24046 ( .A1(n38846), .A2(n22638), .Z(n12760) );
  XNOR2_X1 U24047 ( .A1(n22562), .A2(n22775), .ZN(n22638) );
  XOR2_X1 U24049 ( .A1(n34188), .A2(n37660), .Z(n38846) );
  NAND2_X2 U24054 ( .A1(n39182), .A2(n5494), .ZN(n38847) );
  NOR2_X2 U24056 ( .A1(n32745), .A2(n875), .ZN(n30365) );
  INV_X1 U24064 ( .I(n16053), .ZN(n22893) );
  NAND2_X1 U24066 ( .A1(n35246), .A2(n19594), .ZN(n16053) );
  XOR2_X1 U24068 ( .A1(n16526), .A2(n19527), .Z(n12297) );
  OAI21_X1 U24070 ( .A1(n37734), .A2(n30220), .B(n30158), .ZN(n2322) );
  XOR2_X1 U24072 ( .A1(n29057), .A2(n38962), .Z(n9131) );
  XOR2_X1 U24083 ( .A1(n12839), .A2(n30006), .Z(n10598) );
  NAND2_X2 U24084 ( .A1(n36949), .A2(n36951), .ZN(n12839) );
  NAND2_X2 U24086 ( .A1(n34010), .A2(n9526), .ZN(n19785) );
  XNOR2_X1 U24088 ( .A1(n13138), .A2(n18544), .ZN(n38849) );
  NOR2_X2 U24091 ( .A1(n6347), .A2(n22019), .ZN(n7355) );
  INV_X2 U24092 ( .I(n22574), .ZN(n35446) );
  BUF_X2 U24094 ( .I(n15439), .Z(n38850) );
  BUF_X2 U24099 ( .I(n15794), .Z(n38851) );
  XOR2_X1 U24107 ( .A1(n27830), .A2(n15776), .Z(n27635) );
  NAND2_X2 U24108 ( .A1(n26890), .A2(n34113), .ZN(n15776) );
  INV_X4 U24109 ( .I(n19998), .ZN(n997) );
  NAND2_X2 U24110 ( .A1(n3349), .A2(n19172), .ZN(n19998) );
  NOR2_X1 U24113 ( .A1(n13298), .A2(n34033), .ZN(n39436) );
  AND2_X1 U24117 ( .A1(n27137), .A2(n38853), .Z(n34660) );
  NAND2_X2 U24122 ( .A1(n34738), .A2(n9109), .ZN(n2431) );
  NAND2_X2 U24123 ( .A1(n31679), .A2(n35893), .ZN(n7846) );
  NAND2_X2 U24125 ( .A1(n3664), .A2(n28560), .ZN(n28563) );
  XOR2_X1 U24127 ( .A1(n2943), .A2(n16017), .Z(n16019) );
  NAND2_X2 U24138 ( .A1(n18625), .A2(n18624), .ZN(n2943) );
  NAND2_X1 U24142 ( .A1(n30548), .A2(n14845), .ZN(n38859) );
  NAND2_X1 U24143 ( .A1(n38614), .A2(n23423), .ZN(n14163) );
  NAND2_X2 U24144 ( .A1(n25635), .A2(n25634), .ZN(n13712) );
  XOR2_X1 U24146 ( .A1(n17727), .A2(n31214), .Z(n22438) );
  NAND2_X2 U24147 ( .A1(n3967), .A2(n3969), .ZN(n31214) );
  XOR2_X1 U24152 ( .A1(n12104), .A2(n12103), .Z(n31784) );
  INV_X2 U24161 ( .I(n10940), .ZN(n16590) );
  BUF_X2 U24163 ( .I(n14193), .Z(n38860) );
  NOR2_X2 U24168 ( .A1(n5156), .A2(n38861), .ZN(n5154) );
  INV_X2 U24171 ( .I(n25261), .ZN(n38862) );
  NOR2_X1 U24183 ( .A1(n37052), .A2(n11727), .ZN(n38863) );
  NOR2_X1 U24190 ( .A1(n12370), .A2(n5456), .ZN(n18670) );
  XOR2_X1 U24191 ( .A1(n27541), .A2(n27581), .Z(n32015) );
  NAND2_X2 U24193 ( .A1(n16997), .A2(n17829), .ZN(n27541) );
  OAI21_X2 U24195 ( .A1(n38865), .A2(n38864), .B(n21264), .ZN(n11001) );
  NOR2_X2 U24196 ( .A1(n32720), .A2(n29587), .ZN(n38865) );
  XOR2_X1 U24198 ( .A1(n11746), .A2(n11747), .Z(n19783) );
  AOI22_X2 U24204 ( .A1(n20791), .A2(n18920), .B1(n37468), .B2(n8735), .ZN(
        n24113) );
  XOR2_X1 U24207 ( .A1(n26489), .A2(n26553), .Z(n12300) );
  NAND2_X2 U24226 ( .A1(n7168), .A2(n7171), .ZN(n26489) );
  AOI21_X2 U24227 ( .A1(n32367), .A2(n32368), .B(n1567), .ZN(n38867) );
  OR2_X2 U24236 ( .A1(n32854), .A2(n11342), .Z(n30274) );
  NAND2_X2 U24243 ( .A1(n10996), .A2(n38869), .ZN(n22599) );
  XOR2_X1 U24246 ( .A1(n39742), .A2(n27169), .Z(n38870) );
  XOR2_X1 U24249 ( .A1(n38872), .A2(n34152), .Z(n34957) );
  XOR2_X1 U24254 ( .A1(n15529), .A2(n26601), .Z(n38872) );
  XNOR2_X1 U24257 ( .A1(n36386), .A2(n27534), .ZN(n479) );
  NAND2_X2 U24261 ( .A1(n31302), .A2(n36805), .ZN(n27534) );
  XOR2_X1 U24265 ( .A1(n5516), .A2(n709), .Z(n34200) );
  INV_X2 U24266 ( .I(n13311), .ZN(n36251) );
  NOR2_X2 U24267 ( .A1(n15289), .A2(n15290), .ZN(n13311) );
  NOR2_X1 U24283 ( .A1(n38874), .A2(n20053), .ZN(n1997) );
  INV_X2 U24289 ( .I(n15925), .ZN(n38874) );
  NAND2_X2 U24290 ( .A1(n24795), .A2(n35981), .ZN(n24597) );
  NAND2_X2 U24293 ( .A1(n14051), .A2(n14050), .ZN(n24795) );
  XOR2_X1 U24294 ( .A1(n6717), .A2(n15162), .Z(n38875) );
  XOR2_X1 U24295 ( .A1(n820), .A2(n38876), .Z(n13873) );
  XOR2_X1 U24308 ( .A1(n14350), .A2(n25260), .Z(n38876) );
  XOR2_X1 U24314 ( .A1(n26590), .A2(n26357), .Z(n26558) );
  OAI21_X2 U24315 ( .A1(n12895), .A2(n4801), .B(n25766), .ZN(n26590) );
  BUF_X2 U24318 ( .I(n19202), .Z(n38878) );
  AOI21_X2 U24319 ( .A1(n15943), .A2(n1119), .B(n38879), .ZN(n16581) );
  NOR3_X2 U24320 ( .A1(n38182), .A2(n3076), .A3(n30843), .ZN(n38879) );
  XOR2_X1 U24322 ( .A1(n23830), .A2(n38882), .Z(n5086) );
  XOR2_X1 U24323 ( .A1(n5959), .A2(n1612), .Z(n38882) );
  XOR2_X1 U24324 ( .A1(n23973), .A2(n9043), .Z(n23850) );
  MUX2_X1 U24334 ( .I0(n25931), .I1(n11888), .S(n38247), .Z(n15834) );
  XOR2_X1 U24340 ( .A1(n33511), .A2(n7288), .Z(n15810) );
  OR2_X1 U24341 ( .A1(n19424), .A2(n29900), .Z(n15358) );
  AND2_X1 U24342 ( .A1(n28079), .A2(n20860), .Z(n5022) );
  AOI21_X1 U24344 ( .A1(n8520), .A2(n38976), .B(n1687), .ZN(n7897) );
  XOR2_X1 U24345 ( .A1(n11308), .A2(n19221), .Z(n22650) );
  NAND2_X2 U24346 ( .A1(n7895), .A2(n11047), .ZN(n11308) );
  XOR2_X1 U24347 ( .A1(n28844), .A2(n2392), .Z(n38885) );
  NOR2_X2 U24348 ( .A1(n39687), .A2(n25450), .ZN(n26048) );
  OAI22_X2 U24349 ( .A1(n33459), .A2(n4957), .B1(n24172), .B2(n2268), .ZN(
        n24625) );
  NAND2_X2 U24352 ( .A1(n15559), .A2(n15558), .ZN(n20346) );
  XOR2_X1 U24353 ( .A1(n21036), .A2(n21149), .Z(n21035) );
  INV_X2 U24355 ( .I(n38887), .ZN(n39816) );
  XOR2_X1 U24359 ( .A1(n11119), .A2(n11118), .Z(n38887) );
  NOR2_X2 U24362 ( .A1(n1635), .A2(n30881), .ZN(n23256) );
  OAI22_X2 U24363 ( .A1(n3803), .A2(n20840), .B1(n34013), .B2(n13635), .ZN(
        n4143) );
  INV_X2 U24372 ( .I(n16265), .ZN(n30315) );
  OAI22_X2 U24376 ( .A1(n32663), .A2(n15926), .B1(n15929), .B2(n21694), .ZN(
        n16265) );
  INV_X2 U24377 ( .I(n33258), .ZN(n8006) );
  NAND3_X1 U24380 ( .A1(n3906), .A2(n962), .A3(n15911), .ZN(n12696) );
  OAI21_X2 U24382 ( .A1(n19564), .A2(n27180), .B(n33773), .ZN(n27110) );
  OR2_X1 U24387 ( .A1(n7843), .A2(n30800), .Z(n22199) );
  NAND3_X2 U24391 ( .A1(n20975), .A2(n4188), .A3(n17765), .ZN(n24924) );
  XOR2_X1 U24396 ( .A1(n38888), .A2(n3427), .Z(n3424) );
  XOR2_X1 U24404 ( .A1(n8183), .A2(n3426), .Z(n38888) );
  XOR2_X1 U24407 ( .A1(n38889), .A2(n25202), .Z(n320) );
  XOR2_X1 U24409 ( .A1(n38992), .A2(n25256), .Z(n38889) );
  NAND2_X1 U24410 ( .A1(n33879), .A2(n7901), .ZN(n31432) );
  NAND2_X2 U24421 ( .A1(n18599), .A2(n12416), .ZN(n33879) );
  XOR2_X1 U24422 ( .A1(n16556), .A2(n16558), .Z(n38901) );
  XOR2_X1 U24426 ( .A1(n5116), .A2(n23659), .Z(n38890) );
  NAND2_X2 U24427 ( .A1(n38891), .A2(n32789), .ZN(n34692) );
  NAND3_X2 U24428 ( .A1(n34940), .A2(n260), .A3(n34087), .ZN(n38891) );
  AOI22_X2 U24431 ( .A1(n38892), .A2(n23234), .B1(n20450), .B2(n23292), .ZN(
        n35301) );
  XOR2_X1 U24439 ( .A1(n25185), .A2(n38895), .Z(n1817) );
  OAI21_X2 U24442 ( .A1(n9367), .A2(n26929), .B(n38912), .ZN(n9369) );
  NAND2_X2 U24446 ( .A1(n27562), .A2(n27078), .ZN(n27731) );
  NAND2_X2 U24452 ( .A1(n33908), .A2(n14086), .ZN(n27562) );
  NAND2_X2 U24458 ( .A1(n34913), .A2(n27085), .ZN(n14058) );
  XOR2_X1 U24472 ( .A1(n18807), .A2(n23814), .Z(n19991) );
  NAND3_X2 U24473 ( .A1(n15604), .A2(n15603), .A3(n14576), .ZN(n18807) );
  NAND2_X2 U24475 ( .A1(n38897), .A2(n2404), .ZN(n22317) );
  OAI21_X2 U24485 ( .A1(n2628), .A2(n21924), .B(n38898), .ZN(n38897) );
  OAI22_X2 U24487 ( .A1(n35160), .A2(n16072), .B1(n16073), .B2(n34436), .ZN(
        n35648) );
  BUF_X2 U24488 ( .I(n6390), .Z(n38899) );
  XOR2_X1 U24497 ( .A1(n33083), .A2(n29887), .Z(n39141) );
  BUF_X2 U24503 ( .I(n14153), .Z(n38900) );
  XOR2_X1 U24505 ( .A1(n38902), .A2(n3701), .Z(n15794) );
  XOR2_X1 U24514 ( .A1(n39145), .A2(n10384), .Z(n38902) );
  NAND2_X2 U24528 ( .A1(n38904), .A2(n6048), .ZN(n22574) );
  NAND2_X2 U24536 ( .A1(n38921), .A2(n38920), .ZN(n38904) );
  XOR2_X1 U24542 ( .A1(n20152), .A2(n20151), .Z(n20153) );
  NAND2_X1 U24543 ( .A1(n39527), .A2(n32981), .ZN(n34131) );
  XOR2_X1 U24546 ( .A1(n6165), .A2(n30661), .Z(n32981) );
  XOR2_X1 U24547 ( .A1(n23936), .A2(n38905), .Z(n7558) );
  XOR2_X1 U24548 ( .A1(n25146), .A2(n38192), .Z(n32346) );
  AOI21_X1 U24551 ( .A1(n425), .A2(n15677), .B(n11734), .ZN(n25739) );
  INV_X2 U24556 ( .I(n34692), .ZN(n425) );
  NOR2_X2 U24560 ( .A1(n13607), .A2(n14600), .ZN(n10606) );
  INV_X2 U24562 ( .I(n7643), .ZN(n14600) );
  XOR2_X1 U24567 ( .A1(n17906), .A2(n17905), .Z(n7643) );
  NAND2_X2 U24569 ( .A1(n7625), .A2(n38908), .ZN(n38907) );
  NAND2_X2 U24570 ( .A1(n26063), .A2(n25941), .ZN(n38909) );
  AOI21_X2 U24571 ( .A1(n7454), .A2(n28494), .B(n35173), .ZN(n1944) );
  NOR2_X2 U24581 ( .A1(n9366), .A2(n7523), .ZN(n38912) );
  XOR2_X1 U24588 ( .A1(n28909), .A2(n38913), .Z(n31089) );
  XOR2_X1 U24590 ( .A1(n248), .A2(n17784), .Z(n38913) );
  XOR2_X1 U24594 ( .A1(n34752), .A2(n8844), .Z(n19226) );
  NAND2_X2 U24595 ( .A1(n3429), .A2(n12358), .ZN(n34813) );
  OAI21_X2 U24597 ( .A1(n23154), .A2(n22919), .B(n14738), .ZN(n33847) );
  NOR2_X2 U24598 ( .A1(n8173), .A2(n5957), .ZN(n24769) );
  OAI21_X2 U24600 ( .A1(n33598), .A2(n30339), .B(n28193), .ZN(n31098) );
  OAI22_X2 U24602 ( .A1(n36175), .A2(n3091), .B1(n26835), .B2(n16970), .ZN(
        n31014) );
  NAND3_X2 U24605 ( .A1(n23266), .A2(n23265), .A3(n23267), .ZN(n23905) );
  AOI21_X2 U24607 ( .A1(n17397), .A2(n7541), .B(n28681), .ZN(n28362) );
  INV_X2 U24617 ( .I(n13594), .ZN(n28681) );
  NOR2_X2 U24622 ( .A1(n2416), .A2(n37086), .ZN(n25366) );
  NAND2_X1 U24623 ( .A1(n28034), .A2(n36979), .ZN(n27956) );
  BUF_X2 U24628 ( .I(n34350), .Z(n38914) );
  NAND2_X2 U24632 ( .A1(n38915), .A2(n36767), .ZN(n34541) );
  NAND2_X2 U24633 ( .A1(n19785), .A2(n17894), .ZN(n38915) );
  NAND2_X2 U24644 ( .A1(n928), .A2(n38914), .ZN(n33109) );
  INV_X2 U24650 ( .I(n38916), .ZN(n24910) );
  NAND2_X1 U24651 ( .A1(n825), .A2(n25309), .ZN(n19968) );
  XOR2_X1 U24652 ( .A1(n25062), .A2(n25061), .Z(n25309) );
  INV_X1 U24653 ( .I(n39460), .ZN(n24073) );
  XOR2_X1 U24660 ( .A1(n26381), .A2(n26516), .Z(n21142) );
  NAND2_X2 U24662 ( .A1(n25655), .A2(n34486), .ZN(n26381) );
  XOR2_X1 U24665 ( .A1(n23623), .A2(n24012), .Z(n20777) );
  NAND2_X2 U24667 ( .A1(n18123), .A2(n18370), .ZN(n24012) );
  NOR2_X2 U24668 ( .A1(n32483), .A2(n38918), .ZN(n30504) );
  INV_X2 U24670 ( .I(n38922), .ZN(n34040) );
  NAND2_X2 U24672 ( .A1(n35443), .A2(n31986), .ZN(n38922) );
  NAND2_X2 U24676 ( .A1(n12279), .A2(n38925), .ZN(n24545) );
  NAND2_X1 U24681 ( .A1(n25943), .A2(n25345), .ZN(n3926) );
  OAI22_X2 U24685 ( .A1(n34083), .A2(n12599), .B1(n34487), .B2(n12601), .ZN(
        n25943) );
  NAND2_X2 U24690 ( .A1(n16250), .A2(n25989), .ZN(n26081) );
  NAND2_X2 U24692 ( .A1(n9479), .A2(n17173), .ZN(n16250) );
  AND2_X2 U24694 ( .A1(n14601), .A2(n35269), .Z(n30348) );
  AOI22_X2 U24697 ( .A1(n35137), .A2(n39317), .B1(n39406), .B2(n24879), .ZN(
        n24547) );
  XOR2_X1 U24705 ( .A1(n38927), .A2(n9436), .Z(n9435) );
  NAND3_X1 U24709 ( .A1(n36775), .A2(n19349), .A3(n38220), .ZN(n7480) );
  NOR2_X2 U24713 ( .A1(n35594), .A2(n38929), .ZN(n13075) );
  NOR2_X1 U24715 ( .A1(n25544), .A2(n15515), .ZN(n9816) );
  OAI21_X1 U24719 ( .A1(n25966), .A2(n18320), .B(n25962), .ZN(n38930) );
  NAND2_X2 U24724 ( .A1(n38933), .A2(n35448), .ZN(n5753) );
  NOR2_X2 U24728 ( .A1(n26), .A2(n22317), .ZN(n2028) );
  XOR2_X1 U24742 ( .A1(n26475), .A2(n34630), .Z(n14752) );
  XNOR2_X1 U24745 ( .A1(n29242), .A2(n9035), .ZN(n18526) );
  OAI22_X2 U24746 ( .A1(n4878), .A2(n28664), .B1(n15580), .B2(n12990), .ZN(
        n29242) );
  XOR2_X1 U24747 ( .A1(n11867), .A2(n20692), .Z(n35324) );
  XOR2_X1 U24759 ( .A1(n3161), .A2(n38934), .Z(n13039) );
  XOR2_X1 U24783 ( .A1(n3778), .A2(n3777), .Z(n38934) );
  NAND2_X2 U24788 ( .A1(n37080), .A2(n18990), .ZN(n19409) );
  NAND2_X2 U24790 ( .A1(n1444), .A2(n33955), .ZN(n28240) );
  INV_X4 U24791 ( .I(n38965), .ZN(n34001) );
  XOR2_X1 U24792 ( .A1(n29108), .A2(n38167), .Z(n9972) );
  XOR2_X1 U24795 ( .A1(n36255), .A2(n36254), .Z(n2142) );
  AOI22_X2 U24797 ( .A1(n12745), .A2(n9756), .B1(n12744), .B2(n7588), .ZN(
        n17349) );
  XOR2_X1 U24799 ( .A1(n5843), .A2(n38935), .Z(n39570) );
  XOR2_X1 U24800 ( .A1(n13935), .A2(n39609), .Z(n38935) );
  XOR2_X1 U24809 ( .A1(n20589), .A2(n4127), .Z(n27692) );
  NAND2_X2 U24813 ( .A1(n11089), .A2(n11087), .ZN(n4127) );
  XOR2_X1 U24826 ( .A1(n2170), .A2(n2168), .Z(n10559) );
  NAND2_X2 U24828 ( .A1(n39502), .A2(n38936), .ZN(n15792) );
  OAI21_X2 U24836 ( .A1(n10518), .A2(n10519), .B(n11891), .ZN(n38936) );
  INV_X2 U24837 ( .I(n20589), .ZN(n38937) );
  XOR2_X1 U24839 ( .A1(n8741), .A2(n33373), .Z(n17064) );
  XOR2_X1 U24841 ( .A1(n21077), .A2(n4856), .Z(n21074) );
  NAND2_X1 U24842 ( .A1(n3944), .A2(n5028), .ZN(n28644) );
  XOR2_X1 U24846 ( .A1(n523), .A2(n4393), .Z(n3526) );
  OAI21_X2 U24851 ( .A1(n38938), .A2(n14846), .B(n21406), .ZN(n22155) );
  NAND2_X2 U24852 ( .A1(n19210), .A2(n16177), .ZN(n38939) );
  XOR2_X1 U24853 ( .A1(n25154), .A2(n38940), .Z(n33058) );
  XOR2_X1 U24861 ( .A1(n36980), .A2(n33208), .Z(n38940) );
  XOR2_X1 U24865 ( .A1(Plaintext[155]), .A2(Key[155]), .Z(n39519) );
  NAND2_X1 U24869 ( .A1(n1265), .A2(n35893), .ZN(n38942) );
  XOR2_X1 U24870 ( .A1(n2436), .A2(n35425), .Z(n16631) );
  XOR2_X1 U24876 ( .A1(n4592), .A2(n9043), .Z(n23961) );
  NAND2_X2 U24880 ( .A1(n35285), .A2(n23648), .ZN(n4592) );
  INV_X4 U24883 ( .I(n25956), .ZN(n19740) );
  NAND2_X2 U24885 ( .A1(n34541), .A2(n11954), .ZN(n25956) );
  NAND2_X2 U24889 ( .A1(n14896), .A2(n14897), .ZN(n33996) );
  XOR2_X1 U24893 ( .A1(n38943), .A2(n19677), .Z(Ciphertext[163]) );
  OAI21_X1 U24894 ( .A1(n21006), .A2(n21005), .B(n30127), .ZN(n38943) );
  OAI21_X1 U24895 ( .A1(n8728), .A2(n38945), .B(n38944), .ZN(n29230) );
  AOI21_X2 U24897 ( .A1(n36979), .A2(n14376), .B(n38946), .ZN(n13323) );
  NAND2_X2 U24898 ( .A1(n28189), .A2(n16327), .ZN(n38947) );
  XOR2_X1 U24901 ( .A1(n10129), .A2(n27520), .Z(n13751) );
  NAND2_X2 U24904 ( .A1(n20245), .A2(n26806), .ZN(n32191) );
  OAI22_X1 U24905 ( .A1(n28736), .A2(n36935), .B1(n34861), .B2(n9686), .ZN(
        n28059) );
  NAND2_X2 U24907 ( .A1(n36209), .A2(n36640), .ZN(n35901) );
  NAND2_X2 U24910 ( .A1(n6800), .A2(n6799), .ZN(n39489) );
  NAND3_X2 U24911 ( .A1(n2417), .A2(n20881), .A3(n30694), .ZN(n38949) );
  XOR2_X1 U24918 ( .A1(n38209), .A2(n7481), .Z(n13324) );
  NAND2_X1 U24923 ( .A1(n29596), .A2(n29592), .ZN(n9865) );
  XOR2_X1 U24925 ( .A1(n25139), .A2(n25138), .Z(n25619) );
  NAND2_X2 U24931 ( .A1(n38952), .A2(n34967), .ZN(n4246) );
  NAND2_X2 U24935 ( .A1(n26081), .A2(n38953), .ZN(n38952) );
  NOR2_X1 U24936 ( .A1(n9135), .A2(n35314), .ZN(n15715) );
  XOR2_X1 U24943 ( .A1(n19374), .A2(n29151), .Z(n16193) );
  XOR2_X1 U24949 ( .A1(n38954), .A2(n14866), .Z(n30946) );
  XOR2_X1 U24950 ( .A1(n26508), .A2(n39596), .Z(n38954) );
  NOR2_X1 U24958 ( .A1(n19700), .A2(n19364), .ZN(n35297) );
  NAND2_X2 U24963 ( .A1(n5983), .A2(n31110), .ZN(n31535) );
  XOR2_X1 U24967 ( .A1(n22749), .A2(n22580), .Z(n22752) );
  NOR2_X2 U24976 ( .A1(n17637), .A2(n17634), .ZN(n22749) );
  AOI21_X2 U24977 ( .A1(n37104), .A2(n30859), .B(n26990), .ZN(n38955) );
  XOR2_X1 U24982 ( .A1(n5233), .A2(n37214), .Z(n39347) );
  NAND2_X2 U24986 ( .A1(n8977), .A2(n11924), .ZN(n19580) );
  INV_X2 U24988 ( .I(n20297), .ZN(n29346) );
  XOR2_X1 U24989 ( .A1(n13358), .A2(n13052), .Z(n20297) );
  OAI21_X2 U24990 ( .A1(n38956), .A2(n37239), .B(n424), .ZN(n6845) );
  INV_X2 U24992 ( .I(n27137), .ZN(n27350) );
  NAND2_X2 U24993 ( .A1(n39041), .A2(n34974), .ZN(n27137) );
  NAND2_X2 U24996 ( .A1(n3263), .A2(n14933), .ZN(n18070) );
  OR2_X1 U24998 ( .A1(n17197), .A2(n20056), .Z(n27929) );
  AOI21_X2 U25007 ( .A1(n1108), .A2(n952), .B(n17029), .ZN(n10530) );
  NAND3_X2 U25010 ( .A1(n3806), .A2(n3807), .A3(n32035), .ZN(n8972) );
  AOI22_X2 U25022 ( .A1(n5020), .A2(n28168), .B1(n28167), .B2(n7528), .ZN(
        n38957) );
  AOI22_X2 U25023 ( .A1(n8355), .A2(n14857), .B1(n12633), .B2(n12632), .ZN(
        n25252) );
  NAND2_X1 U25032 ( .A1(n9633), .A2(n38193), .ZN(n27114) );
  INV_X1 U25033 ( .I(n18526), .ZN(n31822) );
  AOI21_X2 U25036 ( .A1(n9599), .A2(n35888), .B(n4992), .ZN(n4991) );
  XOR2_X1 U25037 ( .A1(n7328), .A2(n25319), .Z(n36039) );
  BUF_X2 U25042 ( .I(n30494), .Z(n38960) );
  INV_X2 U25047 ( .I(n8423), .ZN(n35369) );
  NAND3_X2 U25050 ( .A1(n14116), .A2(n14115), .A3(n10032), .ZN(n27810) );
  AOI22_X2 U25055 ( .A1(n6097), .A2(n2835), .B1(n5327), .B2(n1519), .ZN(n26365) );
  XOR2_X1 U25065 ( .A1(n31617), .A2(n22203), .Z(n780) );
  NAND2_X2 U25069 ( .A1(n30603), .A2(n34252), .ZN(n30764) );
  NAND2_X2 U25072 ( .A1(n36187), .A2(n38961), .ZN(n11003) );
  NAND3_X1 U25091 ( .A1(n34103), .A2(n34411), .A3(n13943), .ZN(n38961) );
  XOR2_X1 U25092 ( .A1(n36497), .A2(n4540), .Z(n33848) );
  XOR2_X1 U25093 ( .A1(n34718), .A2(n38962), .Z(n660) );
  XOR2_X1 U25096 ( .A1(n1238), .A2(n26476), .Z(n26522) );
  NAND2_X2 U25097 ( .A1(n35992), .A2(n8133), .ZN(n26476) );
  NAND2_X2 U25109 ( .A1(n39002), .A2(n35839), .ZN(n18686) );
  OR2_X1 U25113 ( .A1(n25639), .A2(n38963), .Z(n39053) );
  NAND2_X2 U25114 ( .A1(n2798), .A2(n39401), .ZN(n10739) );
  OR2_X2 U25122 ( .A1(n20945), .A2(n10816), .Z(n13607) );
  XOR2_X1 U25125 ( .A1(n20618), .A2(n34856), .Z(n2209) );
  XOR2_X1 U25126 ( .A1(n36668), .A2(n29820), .Z(n17159) );
  INV_X2 U25131 ( .I(n38966), .ZN(n14081) );
  XOR2_X1 U25133 ( .A1(n8887), .A2(n29258), .Z(n35142) );
  XOR2_X1 U25136 ( .A1(n38968), .A2(n19217), .Z(n26545) );
  XOR2_X1 U25139 ( .A1(n27193), .A2(n27194), .Z(n38969) );
  OAI21_X2 U25142 ( .A1(n19379), .A2(n16774), .B(n38971), .ZN(n1919) );
  OAI21_X2 U25145 ( .A1(n19070), .A2(n8041), .B(n24257), .ZN(n23652) );
  NAND2_X2 U25146 ( .A1(n33104), .A2(n38972), .ZN(n24257) );
  INV_X2 U25158 ( .I(n18269), .ZN(n38972) );
  XOR2_X1 U25164 ( .A1(n38974), .A2(n13967), .Z(n33576) );
  XOR2_X1 U25173 ( .A1(n39582), .A2(n25238), .Z(n38974) );
  XOR2_X1 U25175 ( .A1(n26529), .A2(n26527), .Z(n5312) );
  XOR2_X1 U25177 ( .A1(n1986), .A2(n39529), .Z(n15853) );
  XOR2_X1 U25180 ( .A1(n1791), .A2(n38975), .Z(n39433) );
  NAND2_X2 U25182 ( .A1(n32524), .A2(n34301), .ZN(n7744) );
  AOI22_X2 U25196 ( .A1(n39283), .A2(n4781), .B1(n27306), .B2(n26791), .ZN(
        n32248) );
  XOR2_X1 U25198 ( .A1(n38977), .A2(n18700), .Z(Ciphertext[45]) );
  NOR2_X1 U25203 ( .A1(n19689), .A2(n29436), .ZN(n38977) );
  XOR2_X1 U25205 ( .A1(n27717), .A2(n37881), .Z(n10562) );
  NAND2_X2 U25208 ( .A1(n36343), .A2(n30373), .ZN(n24802) );
  NAND2_X2 U25209 ( .A1(n25954), .A2(n365), .ZN(n36008) );
  NAND2_X1 U25213 ( .A1(n22473), .A2(n34131), .ZN(n39199) );
  BUF_X2 U25217 ( .I(n26421), .Z(n38979) );
  AOI21_X2 U25219 ( .A1(n38980), .A2(n18877), .B(n12142), .ZN(n22292) );
  NAND2_X2 U25227 ( .A1(n36358), .A2(n15626), .ZN(n38980) );
  OR2_X1 U25237 ( .A1(n25861), .A2(n1107), .Z(n12710) );
  INV_X1 U25239 ( .I(n33997), .ZN(n38982) );
  NAND2_X2 U25240 ( .A1(n4150), .A2(n4151), .ZN(n28104) );
  NAND2_X2 U25242 ( .A1(n3914), .A2(n34939), .ZN(n7018) );
  NAND2_X2 U25247 ( .A1(n12171), .A2(n12170), .ZN(n14153) );
  NOR2_X2 U25249 ( .A1(n31876), .A2(n32869), .ZN(n1882) );
  NOR2_X2 U25251 ( .A1(n15890), .A2(n33792), .ZN(n39528) );
  NOR3_X2 U25254 ( .A1(n38600), .A2(n15176), .A3(n17511), .ZN(n35322) );
  XOR2_X1 U25256 ( .A1(n38985), .A2(n701), .Z(n12471) );
  XOR2_X1 U25258 ( .A1(n13652), .A2(n22520), .Z(n38985) );
  INV_X2 U25262 ( .I(n20570), .ZN(n38986) );
  AOI21_X2 U25264 ( .A1(n18484), .A2(n24228), .B(n38987), .ZN(n20229) );
  OAI21_X2 U25268 ( .A1(n30379), .A2(n2396), .B(n2400), .ZN(n38987) );
  XOR2_X1 U25269 ( .A1(n18493), .A2(n29119), .Z(n38988) );
  XOR2_X1 U25271 ( .A1(n6989), .A2(n26599), .Z(n26288) );
  XOR2_X1 U25280 ( .A1(n34653), .A2(n14374), .Z(n38989) );
  AOI22_X2 U25281 ( .A1(n24113), .A2(n18615), .B1(n24112), .B2(n24111), .ZN(
        n15281) );
  XOR2_X1 U25282 ( .A1(n38990), .A2(n1356), .Z(Ciphertext[95]) );
  NOR2_X2 U25287 ( .A1(n39101), .A2(n5949), .ZN(n38990) );
  XOR2_X1 U25289 ( .A1(n9930), .A2(n29092), .Z(n12562) );
  NAND2_X1 U25290 ( .A1(n33964), .A2(n17698), .ZN(n29694) );
  NAND2_X2 U25292 ( .A1(n33843), .A2(n15022), .ZN(n13879) );
  NAND2_X2 U25293 ( .A1(n5994), .A2(n34836), .ZN(n3963) );
  XOR2_X1 U25294 ( .A1(n38991), .A2(Key[151]), .Z(n39031) );
  XOR2_X1 U25300 ( .A1(n39024), .A2(n18452), .Z(n6449) );
  OAI21_X2 U25313 ( .A1(n18501), .A2(n23193), .B(n23192), .ZN(n39070) );
  OAI21_X2 U25320 ( .A1(n26619), .A2(n1236), .B(n14271), .ZN(n26618) );
  BUF_X2 U25326 ( .I(n25006), .Z(n38993) );
  XOR2_X1 U25329 ( .A1(n34902), .A2(n38994), .Z(n3404) );
  XOR2_X1 U25336 ( .A1(n990), .A2(n31602), .Z(n38994) );
  XOR2_X1 U25338 ( .A1(n7689), .A2(n39766), .Z(n13062) );
  NOR2_X2 U25344 ( .A1(n38995), .A2(n18538), .ZN(n23912) );
  NOR3_X1 U25347 ( .A1(n29813), .A2(n38141), .A3(n2792), .ZN(n6650) );
  XOR2_X1 U25358 ( .A1(n16019), .A2(n28947), .Z(n31031) );
  NAND2_X2 U25365 ( .A1(n38999), .A2(n38998), .ZN(n38997) );
  NAND2_X1 U25367 ( .A1(n28644), .A2(n28729), .ZN(n39000) );
  OAI21_X1 U25372 ( .A1(n20368), .A2(n21950), .B(n39658), .ZN(n21786) );
  NAND2_X1 U25375 ( .A1(n6405), .A2(n39423), .ZN(n28382) );
  NAND2_X2 U25376 ( .A1(n12751), .A2(n12752), .ZN(n39002) );
  OR2_X1 U25382 ( .A1(n29543), .A2(n39003), .Z(n7437) );
  OAI22_X2 U25385 ( .A1(n14744), .A2(n39004), .B1(n14743), .B2(n9797), .ZN(
        n23613) );
  NAND2_X2 U25388 ( .A1(n6254), .A2(n39005), .ZN(n6253) );
  OAI21_X2 U25391 ( .A1(n21001), .A2(n19486), .B(n39007), .ZN(n22284) );
  AOI22_X2 U25392 ( .A1(n24290), .A2(n7949), .B1(n1274), .B2(n8690), .ZN(
        n39538) );
  NOR2_X2 U25395 ( .A1(n13970), .A2(n232), .ZN(n24290) );
  INV_X4 U25398 ( .I(n39108), .ZN(n840) );
  XOR2_X1 U25403 ( .A1(n39008), .A2(n24057), .Z(n36066) );
  XOR2_X1 U25406 ( .A1(n14023), .A2(n8920), .Z(n24930) );
  AOI22_X2 U25409 ( .A1(n5921), .A2(n14337), .B1(n29719), .B2(n29720), .ZN(
        n29723) );
  NAND2_X2 U25411 ( .A1(n27343), .A2(n39009), .ZN(n34113) );
  NOR2_X2 U25420 ( .A1(n27344), .A2(n7620), .ZN(n39009) );
  NAND2_X2 U25432 ( .A1(n13875), .A2(n14277), .ZN(n36827) );
  INV_X2 U25439 ( .I(n39011), .ZN(n921) );
  XOR2_X1 U25441 ( .A1(n2547), .A2(n30578), .Z(n39011) );
  BUF_X2 U25447 ( .I(n36539), .Z(n39012) );
  XOR2_X1 U25453 ( .A1(n39665), .A2(n9243), .Z(n24318) );
  XOR2_X1 U25455 ( .A1(n32298), .A2(n27796), .Z(n32149) );
  AOI21_X2 U25456 ( .A1(n2377), .A2(n26871), .B(n36806), .ZN(n32298) );
  OAI21_X2 U25466 ( .A1(n30421), .A2(n24658), .B(n1121), .ZN(n39013) );
  NAND2_X2 U25468 ( .A1(n2796), .A2(n31657), .ZN(n36539) );
  NOR2_X2 U25471 ( .A1(n10030), .A2(n30675), .ZN(n197) );
  OR2_X1 U25472 ( .A1(n1109), .A2(n19153), .Z(n39800) );
  XOR2_X1 U25480 ( .A1(n20794), .A2(n32083), .Z(n20591) );
  OAI22_X2 U25483 ( .A1(n22127), .A2(n22255), .B1(n31481), .B2(n937), .ZN(
        n22731) );
  NAND2_X2 U25485 ( .A1(n24440), .A2(n19584), .ZN(n33457) );
  BUF_X2 U25486 ( .I(n18661), .Z(n39015) );
  NAND2_X2 U25489 ( .A1(n1949), .A2(n39016), .ZN(n15426) );
  AOI21_X2 U25493 ( .A1(n31913), .A2(n20157), .B(n39069), .ZN(n13727) );
  XOR2_X1 U25495 ( .A1(n13736), .A2(n16175), .Z(n10769) );
  OAI22_X2 U25497 ( .A1(n39248), .A2(n26111), .B1(n16860), .B2(n26112), .ZN(
        n14226) );
  BUF_X2 U25515 ( .I(n16803), .Z(n39019) );
  NOR2_X1 U25519 ( .A1(n16931), .A2(n32486), .ZN(n25641) );
  NAND2_X2 U25529 ( .A1(n39749), .A2(n32871), .ZN(n6590) );
  NAND2_X2 U25530 ( .A1(n14759), .A2(n15953), .ZN(n23117) );
  NAND2_X2 U25534 ( .A1(n32133), .A2(n18034), .ZN(n14759) );
  XOR2_X1 U25535 ( .A1(n33470), .A2(n38144), .Z(n16218) );
  NAND2_X2 U25539 ( .A1(n5377), .A2(n31273), .ZN(n33470) );
  NAND4_X2 U25544 ( .A1(n34292), .A2(n30062), .A3(n35095), .A4(n39022), .ZN(
        n39695) );
  NAND2_X2 U25545 ( .A1(n39023), .A2(n16848), .ZN(n27854) );
  NOR2_X2 U25546 ( .A1(n16211), .A2(n24545), .ZN(n24658) );
  XOR2_X1 U25557 ( .A1(n29001), .A2(n29000), .Z(n39024) );
  XOR2_X1 U25562 ( .A1(n27626), .A2(n11236), .Z(n18094) );
  XOR2_X1 U25567 ( .A1(n35270), .A2(n13289), .Z(n27626) );
  AOI21_X1 U25573 ( .A1(n34534), .A2(n29477), .B(n1396), .ZN(n12150) );
  INV_X2 U25574 ( .I(n29468), .ZN(n1396) );
  NOR2_X2 U25576 ( .A1(n23250), .A2(n30299), .ZN(n7631) );
  NAND2_X2 U25579 ( .A1(n33526), .A2(n32943), .ZN(n30299) );
  XOR2_X1 U25580 ( .A1(n12798), .A2(n24045), .Z(n16765) );
  XOR2_X1 U25584 ( .A1(n23697), .A2(n476), .Z(n24045) );
  AND2_X1 U25590 ( .A1(n36995), .A2(n28024), .Z(n20968) );
  NAND3_X1 U25593 ( .A1(n34482), .A2(n1101), .A3(n7110), .ZN(n17312) );
  NOR3_X2 U25598 ( .A1(n33081), .A2(n15651), .A3(n4893), .ZN(n39026) );
  XOR2_X1 U25601 ( .A1(n39027), .A2(n8119), .Z(n35143) );
  NAND2_X2 U25603 ( .A1(n12176), .A2(n11373), .ZN(n18110) );
  NAND2_X2 U25608 ( .A1(n30853), .A2(n35967), .ZN(n26627) );
  XOR2_X1 U25610 ( .A1(n22771), .A2(n13961), .Z(n39028) );
  XOR2_X1 U25611 ( .A1(n27804), .A2(n39029), .Z(n4362) );
  XOR2_X1 U25613 ( .A1(n1464), .A2(n35190), .Z(n39029) );
  INV_X2 U25616 ( .I(n7846), .ZN(n14523) );
  INV_X2 U25621 ( .I(n39031), .ZN(n35116) );
  OAI21_X2 U25626 ( .A1(n13351), .A2(n13350), .B(n5613), .ZN(n37016) );
  NAND2_X2 U25627 ( .A1(n34715), .A2(n32032), .ZN(n15558) );
  XOR2_X1 U25631 ( .A1(n16898), .A2(n22563), .Z(n22712) );
  NOR2_X2 U25633 ( .A1(n35668), .A2(n6557), .ZN(n16898) );
  NAND2_X1 U25634 ( .A1(n6949), .A2(n39152), .ZN(n22330) );
  INV_X2 U25637 ( .I(n39033), .ZN(n34064) );
  OAI21_X2 U25641 ( .A1(n34387), .A2(n4743), .B(n16263), .ZN(n10356) );
  AOI21_X2 U25642 ( .A1(n10352), .A2(n10351), .B(n39035), .ZN(n10349) );
  NOR2_X2 U25653 ( .A1(n30338), .A2(n28024), .ZN(n39035) );
  OAI21_X2 U25657 ( .A1(n35075), .A2(n34690), .B(n33077), .ZN(n24455) );
  NAND2_X2 U25659 ( .A1(n23766), .A2(n23765), .ZN(n13045) );
  NOR2_X1 U25663 ( .A1(n38728), .A2(n38732), .ZN(n34076) );
  NAND3_X2 U25665 ( .A1(n4038), .A2(n1217), .A3(n37076), .ZN(n39036) );
  XOR2_X1 U25667 ( .A1(n13914), .A2(n5003), .Z(n26625) );
  XOR2_X1 U25668 ( .A1(n15093), .A2(n2782), .Z(n39219) );
  BUF_X2 U25671 ( .I(n15737), .Z(n39037) );
  XOR2_X1 U25673 ( .A1(n39040), .A2(n39039), .Z(n39472) );
  NOR2_X2 U25675 ( .A1(n32016), .A2(n31018), .ZN(n39041) );
  INV_X4 U25684 ( .I(n27338), .ZN(n1225) );
  NAND2_X2 U25693 ( .A1(n81), .A2(n35772), .ZN(n27338) );
  OAI22_X2 U25695 ( .A1(n25491), .A2(n9594), .B1(n16113), .B2(n20924), .ZN(
        n33997) );
  XOR2_X1 U25697 ( .A1(n39447), .A2(n39042), .Z(n4291) );
  XOR2_X1 U25698 ( .A1(n22394), .A2(n22557), .Z(n39042) );
  INV_X2 U25702 ( .I(n39043), .ZN(n22925) );
  XOR2_X1 U25705 ( .A1(n25167), .A2(n30330), .Z(n39044) );
  NAND2_X2 U25706 ( .A1(n39046), .A2(n22926), .ZN(n39045) );
  NAND2_X2 U25708 ( .A1(n1235), .A2(n9618), .ZN(n14825) );
  NOR2_X2 U25715 ( .A1(n18055), .A2(n18056), .ZN(n20806) );
  INV_X4 U25716 ( .I(n8942), .ZN(n8707) );
  AND2_X1 U25718 ( .A1(n13492), .A2(n12909), .Z(n28035) );
  NAND2_X2 U25724 ( .A1(n6556), .A2(n14233), .ZN(n22563) );
  XOR2_X1 U25729 ( .A1(n24037), .A2(n18849), .Z(n39049) );
  OAI22_X2 U25734 ( .A1(n2491), .A2(n13588), .B1(n34892), .B2(n26727), .ZN(
        n39051) );
  INV_X2 U25735 ( .I(n39052), .ZN(n19410) );
  XNOR2_X1 U25736 ( .A1(n27646), .A2(n8424), .ZN(n39052) );
  AOI21_X2 U25741 ( .A1(n22999), .A2(n9797), .B(n37062), .ZN(n32614) );
  XOR2_X1 U25743 ( .A1(n37498), .A2(n25123), .Z(n13935) );
  OAI22_X2 U25746 ( .A1(n24744), .A2(n24547), .B1(n11751), .B2(n11642), .ZN(
        n25123) );
  AOI22_X2 U25747 ( .A1(n10698), .A2(n37674), .B1(n23052), .B2(n14556), .ZN(
        n33087) );
  XOR2_X1 U25761 ( .A1(n23781), .A2(n24073), .Z(n2107) );
  INV_X2 U25763 ( .I(n39054), .ZN(n30285) );
  NOR2_X2 U25764 ( .A1(n12360), .A2(n39055), .ZN(n32152) );
  NAND2_X1 U25769 ( .A1(n4525), .A2(n37088), .ZN(n39434) );
  XOR2_X1 U25772 ( .A1(n27707), .A2(n29394), .Z(n7651) );
  NAND2_X2 U25777 ( .A1(n20914), .A2(n32245), .ZN(n27707) );
  NAND2_X1 U25779 ( .A1(n2630), .A2(n32471), .ZN(n39056) );
  AND2_X1 U25780 ( .A1(n23682), .A2(n2394), .Z(n39057) );
  XOR2_X1 U25785 ( .A1(n12300), .A2(n33233), .Z(n39058) );
  NAND2_X1 U25787 ( .A1(n39059), .A2(n37341), .ZN(n13901) );
  AOI21_X2 U25789 ( .A1(n12802), .A2(n12804), .B(n12800), .ZN(n10054) );
  INV_X2 U25792 ( .I(n24761), .ZN(n39059) );
  XOR2_X1 U25793 ( .A1(n22629), .A2(n22652), .Z(n22787) );
  OAI22_X2 U25796 ( .A1(n22077), .A2(n20354), .B1(n20355), .B2(n22078), .ZN(
        n22629) );
  NAND2_X2 U25803 ( .A1(n13727), .A2(n13726), .ZN(n36935) );
  BUF_X2 U25809 ( .I(n26180), .Z(n39063) );
  NAND2_X2 U25813 ( .A1(n39730), .A2(n8208), .ZN(n27581) );
  INV_X1 U25822 ( .I(n3499), .ZN(n39115) );
  NOR3_X1 U25827 ( .A1(n39271), .A2(n24410), .A3(n37467), .ZN(n32818) );
  INV_X2 U25828 ( .I(n10559), .ZN(n39648) );
  NOR2_X2 U25839 ( .A1(n39480), .A2(n31443), .ZN(n39138) );
  AOI21_X2 U25843 ( .A1(n11513), .A2(n17047), .B(n39064), .ZN(n26353) );
  INV_X2 U25846 ( .I(n34279), .ZN(n39065) );
  INV_X2 U25849 ( .I(n27546), .ZN(n20829) );
  OAI22_X2 U25854 ( .A1(n3920), .A2(n27240), .B1(n3921), .B2(n35466), .ZN(
        n27546) );
  AOI22_X1 U25857 ( .A1(n24302), .A2(n24461), .B1(n14509), .B2(n19990), .ZN(
        n39796) );
  AOI21_X2 U25861 ( .A1(n39066), .A2(n17269), .B(n25925), .ZN(n18630) );
  AOI21_X2 U25866 ( .A1(n39068), .A2(n31603), .B(n9025), .ZN(n7893) );
  NOR2_X2 U25868 ( .A1(n10702), .A2(n30240), .ZN(n39068) );
  INV_X4 U25871 ( .I(n30211), .ZN(n39083) );
  NOR2_X1 U25874 ( .A1(n28119), .A2(n28049), .ZN(n39069) );
  OAI22_X1 U25876 ( .A1(n1126), .A2(n37267), .B1(n19864), .B2(n30279), .ZN(
        n31916) );
  XOR2_X1 U25877 ( .A1(n27710), .A2(n27781), .Z(n11730) );
  XOR2_X1 U25879 ( .A1(n23684), .A2(n23683), .Z(n39071) );
  NAND2_X2 U25882 ( .A1(n2628), .A2(n9316), .ZN(n3429) );
  NOR2_X2 U25890 ( .A1(n18657), .A2(n33899), .ZN(n2628) );
  NAND2_X2 U25895 ( .A1(n39072), .A2(n35729), .ZN(n27755) );
  MUX2_X1 U25907 ( .I0(n27119), .I1(n27118), .S(n32976), .Z(n39072) );
  NAND2_X2 U25913 ( .A1(n39501), .A2(n24673), .ZN(n18115) );
  OAI21_X2 U25915 ( .A1(n39165), .A2(n692), .B(n13971), .ZN(n17374) );
  NOR2_X2 U25917 ( .A1(n2798), .A2(n10143), .ZN(n8680) );
  BUF_X2 U25926 ( .I(n24470), .Z(n39074) );
  OAI22_X2 U25933 ( .A1(n18862), .A2(n26038), .B1(n18863), .B2(n25921), .ZN(
        n26511) );
  XOR2_X1 U25935 ( .A1(n36851), .A2(n8177), .Z(n8176) );
  XOR2_X1 U25938 ( .A1(n6746), .A2(n24075), .Z(n31655) );
  AND2_X1 U25942 ( .A1(n25490), .A2(n34427), .Z(n4715) );
  AOI22_X1 U25947 ( .A1(n5723), .A2(n36965), .B1(n35963), .B2(n31931), .ZN(
        n8052) );
  NAND2_X2 U25954 ( .A1(n33087), .A2(n8101), .ZN(n31931) );
  BUF_X4 U25955 ( .I(n36281), .Z(n39075) );
  INV_X1 U25958 ( .I(n39076), .ZN(n2898) );
  INV_X2 U25960 ( .I(n23918), .ZN(n36497) );
  XOR2_X1 U25968 ( .A1(n24034), .A2(n6560), .Z(n23918) );
  OAI21_X1 U25970 ( .A1(n20242), .A2(n21782), .B(n32123), .ZN(n21663) );
  OAI22_X2 U25981 ( .A1(n32202), .A2(n9798), .B1(n13451), .B2(n13450), .ZN(
        n23580) );
  OAI21_X2 U25985 ( .A1(n34081), .A2(n13320), .B(n35419), .ZN(n39077) );
  INV_X2 U25987 ( .I(n26361), .ZN(n39078) );
  NAND2_X2 U25988 ( .A1(n10510), .A2(n10509), .ZN(n26361) );
  NOR2_X1 U25992 ( .A1(n20242), .A2(n32123), .ZN(n20241) );
  OAI21_X1 U25993 ( .A1(n14438), .A2(n3700), .B(n3631), .ZN(n2859) );
  XOR2_X1 U25999 ( .A1(n39080), .A2(n29036), .Z(n2122) );
  XOR2_X1 U26000 ( .A1(n29095), .A2(n19309), .Z(n39080) );
  XOR2_X1 U26003 ( .A1(n22482), .A2(n39081), .Z(n130) );
  XOR2_X1 U26007 ( .A1(n22768), .A2(n33990), .Z(n39081) );
  XOR2_X1 U26008 ( .A1(n3649), .A2(n39082), .Z(n30330) );
  INV_X1 U26019 ( .I(n19953), .ZN(n39082) );
  AOI21_X2 U26039 ( .A1(n21505), .A2(n10345), .B(n32319), .ZN(n22254) );
  OAI21_X2 U26045 ( .A1(n31696), .A2(n30155), .B(n32777), .ZN(n18589) );
  OAI21_X2 U26049 ( .A1(n39107), .A2(n787), .B(n39084), .ZN(n11678) );
  OAI21_X2 U26050 ( .A1(n10018), .A2(n9841), .B(n20873), .ZN(n39084) );
  NOR2_X2 U26051 ( .A1(n35116), .A2(n37111), .ZN(n15019) );
  XOR2_X1 U26052 ( .A1(n27664), .A2(n27574), .Z(n27495) );
  NOR2_X2 U26055 ( .A1(n13721), .A2(n20149), .ZN(n27664) );
  AND2_X1 U26057 ( .A1(n22294), .A2(n22292), .Z(n22139) );
  XOR2_X1 U26058 ( .A1(n39086), .A2(n34152), .Z(n19459) );
  XOR2_X1 U26060 ( .A1(n36508), .A2(n21142), .Z(n39086) );
  NAND2_X2 U26067 ( .A1(n8350), .A2(n39087), .ZN(n28692) );
  NAND2_X2 U26069 ( .A1(n36404), .A2(n2625), .ZN(n31665) );
  XOR2_X1 U26071 ( .A1(n13115), .A2(n29038), .Z(n39088) );
  XOR2_X1 U26072 ( .A1(n1258), .A2(n14385), .Z(n25063) );
  XOR2_X1 U26073 ( .A1(n29096), .A2(n29063), .Z(n19600) );
  NAND3_X2 U26074 ( .A1(n14049), .A2(n6068), .A3(n6071), .ZN(n29096) );
  NAND2_X1 U26076 ( .A1(n13384), .A2(n38163), .ZN(n9263) );
  XOR2_X1 U26080 ( .A1(n2637), .A2(n39088), .Z(n29184) );
  XOR2_X1 U26081 ( .A1(n18620), .A2(n39089), .Z(n35164) );
  XOR2_X1 U26082 ( .A1(n23833), .A2(n18622), .Z(n39089) );
  NAND2_X2 U26084 ( .A1(n39498), .A2(n6541), .ZN(n25319) );
  XOR2_X1 U26087 ( .A1(n39090), .A2(n39310), .Z(n3804) );
  XOR2_X1 U26089 ( .A1(n23885), .A2(n1622), .Z(n39090) );
  NAND2_X1 U26095 ( .A1(n39091), .A2(n1451), .ZN(n19413) );
  OAI22_X1 U26096 ( .A1(n983), .A2(n28050), .B1(n14404), .B2(n28124), .ZN(
        n39091) );
  XOR2_X1 U26100 ( .A1(n18239), .A2(n22427), .Z(n34468) );
  NAND2_X2 U26104 ( .A1(n24624), .A2(n24734), .ZN(n25196) );
  NAND2_X2 U26107 ( .A1(n31712), .A2(n24769), .ZN(n8406) );
  AOI21_X2 U26113 ( .A1(n39092), .A2(n24083), .B(n24082), .ZN(n24735) );
  INV_X2 U26119 ( .I(n39094), .ZN(n19153) );
  XOR2_X1 U26121 ( .A1(n19154), .A2(n24633), .Z(n39094) );
  NAND2_X2 U26126 ( .A1(n39095), .A2(n2152), .ZN(n26263) );
  NAND2_X2 U26133 ( .A1(n39386), .A2(n26325), .ZN(n39095) );
  BUF_X2 U26134 ( .I(n10379), .Z(n39096) );
  INV_X2 U26136 ( .I(n39097), .ZN(n14638) );
  XOR2_X1 U26137 ( .A1(n10343), .A2(n28940), .Z(n39097) );
  XOR2_X1 U26139 ( .A1(n28978), .A2(n29081), .Z(n2004) );
  XOR2_X1 U26142 ( .A1(n29303), .A2(n14956), .Z(n29836) );
  OAI21_X2 U26144 ( .A1(n16920), .A2(n17007), .B(n28757), .ZN(n29303) );
  NAND2_X2 U26146 ( .A1(n959), .A2(n33712), .ZN(n18328) );
  NAND2_X2 U26147 ( .A1(n19965), .A2(n19964), .ZN(n25433) );
  AOI22_X2 U26148 ( .A1(n24363), .A2(n38984), .B1(n36082), .B2(n39099), .ZN(
        n24364) );
  XOR2_X1 U26150 ( .A1(n8277), .A2(n8276), .Z(n39100) );
  INV_X2 U26154 ( .I(n39073), .ZN(n23914) );
  NOR2_X2 U26158 ( .A1(n1270), .A2(n5282), .ZN(n24775) );
  XOR2_X1 U26164 ( .A1(n3885), .A2(n3886), .Z(n28204) );
  XOR2_X1 U26167 ( .A1(n13797), .A2(n39102), .Z(n29312) );
  XOR2_X1 U26168 ( .A1(n11346), .A2(n11922), .Z(n39102) );
  XOR2_X1 U26169 ( .A1(n23737), .A2(n14140), .Z(n39103) );
  XOR2_X1 U26174 ( .A1(n29058), .A2(n12244), .Z(n29304) );
  NAND2_X2 U26178 ( .A1(n28761), .A2(n19794), .ZN(n29058) );
  XOR2_X1 U26191 ( .A1(n10647), .A2(n10644), .Z(n11402) );
  OAI21_X2 U26195 ( .A1(n6293), .A2(n14915), .B(n14914), .ZN(n26055) );
  NAND2_X2 U26197 ( .A1(n34613), .A2(n5672), .ZN(n6293) );
  XOR2_X1 U26202 ( .A1(n39105), .A2(n1322), .Z(n34202) );
  XOR2_X1 U26203 ( .A1(n22588), .A2(n22531), .Z(n39105) );
  INV_X2 U26205 ( .I(n39106), .ZN(n26988) );
  XNOR2_X1 U26209 ( .A1(n13244), .A2(n7720), .ZN(n39106) );
  NOR2_X1 U26213 ( .A1(n23181), .A2(n22903), .ZN(n39107) );
  XOR2_X1 U26216 ( .A1(n26550), .A2(n26551), .Z(n26601) );
  OAI21_X2 U26218 ( .A1(n15552), .A2(n15551), .B(n25784), .ZN(n26551) );
  OAI22_X2 U26221 ( .A1(n4991), .A2(n3598), .B1(n39761), .B2(n34667), .ZN(
        n39189) );
  NAND2_X2 U26224 ( .A1(n4492), .A2(n39109), .ZN(n27690) );
  NAND3_X1 U26226 ( .A1(n27070), .A2(n36989), .A3(n27071), .ZN(n39109) );
  NAND2_X2 U26227 ( .A1(n6844), .A2(n6845), .ZN(n35654) );
  INV_X2 U26234 ( .I(n7023), .ZN(n10544) );
  OAI21_X2 U26235 ( .A1(n39150), .A2(n15986), .B(n27235), .ZN(n5994) );
  XOR2_X1 U26239 ( .A1(n27778), .A2(n27746), .Z(n27788) );
  OAI21_X2 U26245 ( .A1(n5461), .A2(n5462), .B(n39111), .ZN(n20392) );
  XOR2_X1 U26251 ( .A1(n27466), .A2(n32354), .Z(n20846) );
  NAND2_X2 U26254 ( .A1(n37163), .A2(n12814), .ZN(n5408) );
  INV_X2 U26260 ( .I(n39113), .ZN(n36361) );
  XOR2_X1 U26267 ( .A1(Plaintext[139]), .A2(Key[139]), .Z(n39113) );
  XOR2_X1 U26279 ( .A1(n15723), .A2(n39114), .Z(n32932) );
  XOR2_X1 U26282 ( .A1(n15721), .A2(n15722), .Z(n39114) );
  XOR2_X1 U26284 ( .A1(n33722), .A2(n39115), .Z(n15692) );
  XOR2_X1 U26285 ( .A1(n32135), .A2(n30169), .Z(n22627) );
  AOI22_X2 U26290 ( .A1(n4199), .A2(n35755), .B1(n4198), .B2(n31651), .ZN(
        n32135) );
  BUF_X4 U26300 ( .I(n13686), .Z(n39117) );
  NAND2_X2 U26307 ( .A1(n28245), .A2(n28244), .ZN(n28748) );
  XOR2_X1 U26314 ( .A1(n484), .A2(n343), .Z(n39118) );
  XOR2_X1 U26332 ( .A1(n4079), .A2(n4080), .Z(n39119) );
  OAI21_X2 U26333 ( .A1(n2017), .A2(n2016), .B(n2013), .ZN(n31538) );
  NAND3_X2 U26335 ( .A1(n10048), .A2(n14901), .A3(n11436), .ZN(n34421) );
  NAND2_X2 U26338 ( .A1(n8645), .A2(n8644), .ZN(n8875) );
  NAND2_X2 U26342 ( .A1(n12161), .A2(n39120), .ZN(n25263) );
  XOR2_X1 U26364 ( .A1(n39121), .A2(n18014), .Z(n18017) );
  XOR2_X1 U26371 ( .A1(n8240), .A2(n39544), .Z(n39121) );
  BUF_X2 U26372 ( .I(n30183), .Z(n39122) );
  INV_X2 U26374 ( .I(n39123), .ZN(n8205) );
  XNOR2_X1 U26384 ( .A1(n7115), .A2(n7112), .ZN(n39123) );
  NAND2_X1 U26385 ( .A1(n23247), .A2(n35232), .ZN(n13578) );
  OAI22_X2 U26388 ( .A1(n39124), .A2(n39714), .B1(n15633), .B2(n24910), .ZN(
        n24994) );
  INV_X2 U26402 ( .I(n13843), .ZN(n39124) );
  INV_X2 U26413 ( .I(n39125), .ZN(n22962) );
  NOR2_X2 U26419 ( .A1(n10047), .A2(n1046), .ZN(n39125) );
  NAND2_X1 U26425 ( .A1(n13105), .A2(n13104), .ZN(n39170) );
  NAND2_X1 U26427 ( .A1(n12694), .A2(n12505), .ZN(n39128) );
  XOR2_X1 U26434 ( .A1(n34414), .A2(n39130), .Z(n35395) );
  XOR2_X1 U26435 ( .A1(n2317), .A2(n25304), .Z(n39130) );
  XOR2_X1 U26440 ( .A1(n12999), .A2(n27773), .Z(n27751) );
  BUF_X2 U26441 ( .I(n30574), .Z(n39133) );
  NAND2_X2 U26449 ( .A1(n24779), .A2(n24545), .ZN(n24659) );
  OAI21_X2 U26455 ( .A1(n16069), .A2(n18479), .B(n16068), .ZN(n24779) );
  XOR2_X1 U26460 ( .A1(n39468), .A2(n25226), .Z(n15316) );
  NOR2_X2 U26462 ( .A1(n39134), .A2(n21196), .ZN(n29341) );
  AOI22_X2 U26463 ( .A1(n28510), .A2(n28509), .B1(n36414), .B2(n8218), .ZN(
        n8217) );
  XOR2_X1 U26476 ( .A1(n39135), .A2(n26262), .Z(n13853) );
  AND2_X1 U26480 ( .A1(n13278), .A2(n4272), .Z(n39532) );
  NOR2_X2 U26484 ( .A1(n8319), .A2(n24304), .ZN(n12686) );
  XOR2_X1 U26492 ( .A1(n39137), .A2(n6544), .Z(n4997) );
  XOR2_X1 U26499 ( .A1(n37149), .A2(n6546), .Z(n39137) );
  NAND2_X2 U26502 ( .A1(n39138), .A2(n34263), .ZN(n3760) );
  NAND2_X1 U26504 ( .A1(n39142), .A2(n31987), .ZN(n39139) );
  NAND2_X2 U26508 ( .A1(n21300), .A2(n33651), .ZN(n14387) );
  XOR2_X1 U26517 ( .A1(n11059), .A2(n39141), .Z(n31125) );
  XOR2_X1 U26519 ( .A1(n1506), .A2(n26511), .Z(n11059) );
  AND2_X1 U26521 ( .A1(n2001), .A2(n29956), .Z(n32539) );
  OR2_X1 U26525 ( .A1(n39140), .A2(n26055), .Z(n13168) );
  NOR2_X2 U26535 ( .A1(n20061), .A2(n39143), .ZN(n20059) );
  XOR2_X1 U26543 ( .A1(n3663), .A2(n35247), .Z(n35246) );
  XOR2_X1 U26546 ( .A1(n9719), .A2(n39136), .Z(n39145) );
  NOR2_X2 U26548 ( .A1(n10515), .A2(n10516), .ZN(n39502) );
  INV_X4 U26554 ( .I(n4576), .ZN(n7379) );
  OAI21_X2 U26555 ( .A1(n7934), .A2(n8498), .B(n35827), .ZN(n7253) );
  INV_X2 U26556 ( .I(n39148), .ZN(n7934) );
  NAND2_X2 U26560 ( .A1(n2717), .A2(n2716), .ZN(n39148) );
  XOR2_X1 U26561 ( .A1(n39149), .A2(n33954), .Z(n12673) );
  XOR2_X1 U26563 ( .A1(n20820), .A2(n16549), .Z(n39149) );
  XOR2_X1 U26566 ( .A1(n22599), .A2(n22656), .Z(n33177) );
  OAI21_X2 U26567 ( .A1(n8028), .A2(n1047), .B(n6032), .ZN(n22656) );
  XOR2_X1 U26570 ( .A1(n25247), .A2(n25175), .Z(n25185) );
  NOR3_X1 U26579 ( .A1(n12309), .A2(n18121), .A3(n13166), .ZN(n31745) );
  NAND2_X2 U26583 ( .A1(n29627), .A2(n29617), .ZN(n29611) );
  AOI22_X1 U26602 ( .A1(n6948), .A2(n9165), .B1(n10681), .B2(n4108), .ZN(
        n39152) );
  NAND2_X2 U26604 ( .A1(n1147), .A2(n5515), .ZN(n30594) );
  NAND2_X2 U26608 ( .A1(n23518), .A2(n19671), .ZN(n20817) );
  NAND2_X2 U26609 ( .A1(n6919), .A2(n37082), .ZN(n8039) );
  NAND2_X2 U26615 ( .A1(n39158), .A2(n19368), .ZN(n26599) );
  OR2_X1 U26618 ( .A1(n13686), .A2(n17034), .Z(n32527) );
  XOR2_X1 U26621 ( .A1(n39162), .A2(n17872), .Z(n7319) );
  XOR2_X1 U26623 ( .A1(n8884), .A2(n17874), .Z(n39162) );
  XOR2_X1 U26626 ( .A1(n26503), .A2(n26348), .Z(n11620) );
  INV_X4 U26627 ( .I(n7542), .ZN(n13294) );
  NAND2_X2 U26631 ( .A1(n2493), .A2(n39164), .ZN(n11247) );
  INV_X2 U26638 ( .I(n39166), .ZN(n253) );
  XOR2_X1 U26639 ( .A1(n10769), .A2(n10770), .Z(n39166) );
  XOR2_X1 U26643 ( .A1(n32685), .A2(n39167), .Z(n34427) );
  XOR2_X1 U26646 ( .A1(n25129), .A2(n25128), .Z(n39167) );
  XOR2_X1 U26651 ( .A1(n39168), .A2(n34955), .Z(n20958) );
  XOR2_X1 U26653 ( .A1(n22759), .A2(n20865), .Z(n39168) );
  XOR2_X1 U26654 ( .A1(n33870), .A2(n39169), .Z(n19266) );
  XOR2_X1 U26656 ( .A1(n14218), .A2(n1456), .Z(n39169) );
  XOR2_X1 U26657 ( .A1(n39170), .A2(n29221), .Z(Ciphertext[9]) );
  OAI21_X2 U26658 ( .A1(n1034), .A2(n305), .B(n38561), .ZN(n34711) );
  INV_X2 U26661 ( .I(n39171), .ZN(n9333) );
  NAND2_X2 U26663 ( .A1(n37219), .A2(n39204), .ZN(n4576) );
  AOI21_X2 U26667 ( .A1(n19270), .A2(n554), .B(n39173), .ZN(n19268) );
  XOR2_X1 U26673 ( .A1(n25010), .A2(n35339), .Z(n31281) );
  INV_X2 U26675 ( .I(n39175), .ZN(n7982) );
  XOR2_X1 U26680 ( .A1(Plaintext[41]), .A2(Key[41]), .Z(n39175) );
  AOI21_X2 U26693 ( .A1(n34195), .A2(n4337), .B(n4336), .ZN(n4493) );
  XOR2_X1 U26700 ( .A1(n15648), .A2(n9154), .Z(n39177) );
  XOR2_X1 U26708 ( .A1(n5381), .A2(n34722), .Z(n5382) );
  BUF_X2 U26712 ( .I(n10429), .Z(n9914) );
  NAND2_X2 U26713 ( .A1(n4888), .A2(n25473), .ZN(n35059) );
  XOR2_X1 U26717 ( .A1(n13483), .A2(n8602), .Z(n2161) );
  XOR2_X1 U26718 ( .A1(n16054), .A2(n28850), .Z(n8602) );
  NAND2_X2 U26723 ( .A1(n35420), .A2(n32411), .ZN(n28660) );
  OAI21_X2 U26730 ( .A1(n24346), .A2(n7834), .B(n1033), .ZN(n7800) );
  NAND2_X1 U26732 ( .A1(n3863), .A2(n22317), .ZN(n22319) );
  XOR2_X1 U26735 ( .A1(n36386), .A2(n27690), .Z(n3258) );
  OAI21_X2 U26742 ( .A1(n36099), .A2(n2534), .B(n910), .ZN(n2629) );
  NAND2_X2 U26747 ( .A1(n39180), .A2(n28403), .ZN(n31378) );
  NOR2_X1 U26748 ( .A1(n902), .A2(n35777), .ZN(n11094) );
  OAI21_X2 U26750 ( .A1(n39181), .A2(n21564), .B(n21562), .ZN(n35431) );
  INV_X1 U26754 ( .I(n21560), .ZN(n39181) );
  NAND2_X2 U26763 ( .A1(n17792), .A2(n19543), .ZN(n21560) );
  XOR2_X1 U26768 ( .A1(n29121), .A2(n3280), .Z(n11479) );
  AOI21_X2 U26771 ( .A1(n13807), .A2(n28614), .B(n13806), .ZN(n3280) );
  XOR2_X1 U26780 ( .A1(n36329), .A2(n15757), .Z(n878) );
  AOI22_X2 U26783 ( .A1(n6501), .A2(n26909), .B1(n1234), .B2(n26718), .ZN(
        n35794) );
  NOR2_X1 U26788 ( .A1(n26459), .A2(n20891), .ZN(n26718) );
  NAND2_X2 U26790 ( .A1(n2009), .A2(n12982), .ZN(n11372) );
  NAND2_X2 U26798 ( .A1(n39184), .A2(n31634), .ZN(n17791) );
  NOR2_X2 U26799 ( .A1(n18842), .A2(n37160), .ZN(n39184) );
  XOR2_X1 U26804 ( .A1(n39185), .A2(n3726), .Z(n36338) );
  XOR2_X1 U26807 ( .A1(n27673), .A2(n39186), .Z(n39185) );
  NOR2_X1 U26808 ( .A1(n13414), .A2(n12966), .ZN(n2012) );
  NAND2_X2 U26822 ( .A1(n18883), .A2(n36685), .ZN(n28590) );
  XOR2_X1 U26832 ( .A1(n6729), .A2(n6728), .Z(n11145) );
  OR2_X1 U26840 ( .A1(n28047), .A2(n39188), .Z(n34340) );
  NAND2_X2 U26849 ( .A1(n39189), .A2(n28592), .ZN(n28865) );
  AND2_X1 U26852 ( .A1(n4515), .A2(n32979), .Z(n39781) );
  XOR2_X1 U26854 ( .A1(n16755), .A2(n33182), .Z(n35080) );
  OR2_X1 U26856 ( .A1(n6945), .A2(n13370), .Z(n10432) );
  NOR2_X2 U26862 ( .A1(n18505), .A2(n22801), .ZN(n6945) );
  NAND3_X2 U26875 ( .A1(n24772), .A2(n24343), .A3(n3487), .ZN(n11601) );
  NAND2_X2 U26878 ( .A1(n25433), .A2(n7391), .ZN(n15991) );
  AOI21_X1 U26884 ( .A1(n14228), .A2(n951), .B(n39015), .ZN(n18464) );
  NAND2_X2 U26886 ( .A1(n10836), .A2(n11048), .ZN(n28051) );
  OAI21_X2 U26887 ( .A1(n6807), .A2(n19211), .B(n22262), .ZN(n32081) );
  XOR2_X1 U26891 ( .A1(n36305), .A2(n1969), .Z(n24276) );
  XOR2_X1 U26893 ( .A1(n39195), .A2(n24679), .Z(n10309) );
  XOR2_X1 U26894 ( .A1(n24676), .A2(n10199), .Z(n39195) );
  BUF_X4 U26895 ( .I(n985), .Z(n39235) );
  OAI21_X2 U26902 ( .A1(n32260), .A2(n23569), .B(n5792), .ZN(n5791) );
  OR3_X1 U26910 ( .A1(n21687), .A2(n7982), .A3(n21688), .Z(n7965) );
  XOR2_X1 U26913 ( .A1(n19112), .A2(n5802), .Z(n3141) );
  XOR2_X1 U26924 ( .A1(n20347), .A2(n25255), .Z(n33759) );
  NAND2_X2 U26925 ( .A1(n39197), .A2(n17062), .ZN(n15069) );
  NAND2_X2 U26927 ( .A1(n34268), .A2(n39415), .ZN(n39197) );
  NOR2_X2 U26929 ( .A1(n35917), .A2(n17388), .ZN(n39770) );
  XOR2_X1 U26930 ( .A1(n31348), .A2(n6456), .Z(n32534) );
  INV_X1 U26931 ( .I(n2947), .ZN(n999) );
  AOI21_X1 U26939 ( .A1(n39405), .A2(n39406), .B(n39317), .ZN(n15553) );
  NAND2_X2 U26946 ( .A1(n17806), .A2(n31650), .ZN(n39317) );
  OAI21_X1 U26954 ( .A1(n39261), .A2(n7387), .B(n34373), .ZN(n321) );
  AOI22_X2 U26955 ( .A1(n39199), .A2(n23013), .B1(n39198), .B2(n1318), .ZN(
        n23482) );
  OAI21_X2 U26956 ( .A1(n16678), .A2(n5702), .B(n33972), .ZN(n39198) );
  NOR2_X2 U26957 ( .A1(n32654), .A2(n31780), .ZN(n20683) );
  XOR2_X1 U26960 ( .A1(n26261), .A2(n26145), .Z(n26146) );
  NAND2_X2 U26961 ( .A1(n39200), .A2(n18309), .ZN(n1414) );
  AND3_X1 U26970 ( .A1(n28637), .A2(n39355), .A3(n33047), .Z(n39366) );
  XOR2_X1 U26972 ( .A1(n39201), .A2(n6780), .Z(n24280) );
  NAND2_X1 U26975 ( .A1(n29380), .A2(n14151), .ZN(n28901) );
  NAND2_X2 U26979 ( .A1(n1301), .A2(n35963), .ZN(n20998) );
  OAI21_X2 U26987 ( .A1(n39206), .A2(n39203), .B(n27154), .ZN(n3672) );
  NOR2_X2 U26989 ( .A1(n22456), .A2(n39205), .ZN(n39204) );
  XOR2_X1 U26993 ( .A1(n27496), .A2(n27654), .Z(n2042) );
  BUF_X2 U27000 ( .I(n27408), .Z(n39206) );
  XOR2_X1 U27005 ( .A1(n11740), .A2(n17657), .Z(n39207) );
  INV_X2 U27012 ( .I(n18998), .ZN(n9422) );
  NAND3_X2 U27014 ( .A1(n7964), .A2(n7963), .A3(n7965), .ZN(n18998) );
  XOR2_X1 U27018 ( .A1(n39208), .A2(n29371), .Z(Ciphertext[34]) );
  OR2_X1 U27021 ( .A1(n9604), .A2(n36361), .Z(n15626) );
  XOR2_X1 U27023 ( .A1(n1656), .A2(n22762), .Z(n6224) );
  INV_X2 U27026 ( .I(n22228), .ZN(n1331) );
  NOR2_X2 U27034 ( .A1(n20423), .A2(n5935), .ZN(n14921) );
  XOR2_X1 U27037 ( .A1(n22750), .A2(n3172), .Z(n2473) );
  XOR2_X1 U27041 ( .A1(n22492), .A2(n22491), .Z(n22750) );
  NAND2_X2 U27042 ( .A1(n13066), .A2(n13068), .ZN(n26357) );
  XOR2_X1 U27043 ( .A1(n33807), .A2(n39210), .Z(n34802) );
  XOR2_X1 U27044 ( .A1(n61), .A2(n39211), .Z(n39210) );
  INV_X2 U27050 ( .I(n31579), .ZN(n39211) );
  XOR2_X1 U27054 ( .A1(n39212), .A2(n15227), .Z(n17604) );
  XOR2_X1 U27055 ( .A1(n25200), .A2(n15226), .Z(n39212) );
  INV_X2 U27064 ( .I(n39213), .ZN(n34167) );
  NOR2_X2 U27077 ( .A1(n27399), .A2(n12327), .ZN(n39213) );
  OAI21_X2 U27078 ( .A1(n15249), .A2(n28111), .B(n15389), .ZN(n20200) );
  NOR2_X2 U27084 ( .A1(n8368), .A2(n4306), .ZN(n15249) );
  NAND2_X2 U27087 ( .A1(n12604), .A2(n19892), .ZN(n11868) );
  NAND2_X2 U27094 ( .A1(n2022), .A2(n3014), .ZN(n19892) );
  XOR2_X1 U27101 ( .A1(n17957), .A2(n29076), .Z(n5129) );
  XOR2_X1 U27102 ( .A1(n5130), .A2(n29082), .Z(n29076) );
  AOI22_X2 U27106 ( .A1(n11293), .A2(n37582), .B1(n11292), .B2(n7110), .ZN(
        n17890) );
  NAND2_X1 U27109 ( .A1(n17978), .A2(n28559), .ZN(n17977) );
  XOR2_X1 U27111 ( .A1(n38979), .A2(n26568), .Z(n39685) );
  XOR2_X1 U27118 ( .A1(n39217), .A2(n15421), .Z(n14608) );
  XOR2_X1 U27119 ( .A1(n36317), .A2(n27754), .Z(n39217) );
  XOR2_X1 U27120 ( .A1(n25243), .A2(n8163), .Z(n25032) );
  INV_X2 U27121 ( .I(n30619), .ZN(n29074) );
  XOR2_X1 U27122 ( .A1(n28874), .A2(n39220), .Z(n30619) );
  INV_X2 U27123 ( .I(n16309), .ZN(n39220) );
  XOR2_X1 U27124 ( .A1(n25217), .A2(n39221), .Z(n25062) );
  XOR2_X1 U27129 ( .A1(n25316), .A2(n19670), .Z(n39221) );
  XOR2_X1 U27130 ( .A1(n22443), .A2(n22527), .Z(n7510) );
  INV_X4 U27131 ( .I(n31955), .ZN(n27306) );
  NAND2_X1 U27137 ( .A1(n1086), .A2(n35332), .ZN(n15577) );
  NOR2_X2 U27138 ( .A1(n35038), .A2(n34057), .ZN(n31955) );
  AOI21_X2 U27142 ( .A1(n15941), .A2(n37014), .B(n1039), .ZN(n15949) );
  INV_X2 U27144 ( .I(n5363), .ZN(n39305) );
  NAND2_X2 U27149 ( .A1(n39646), .A2(n15999), .ZN(n5363) );
  NOR2_X2 U27155 ( .A1(n5798), .A2(n14472), .ZN(n39224) );
  NAND3_X2 U27160 ( .A1(n12893), .A2(n9146), .A3(n9145), .ZN(n10986) );
  XOR2_X1 U27168 ( .A1(n8300), .A2(n8298), .Z(n15873) );
  XOR2_X1 U27169 ( .A1(n23781), .A2(n23878), .Z(n6379) );
  NAND2_X2 U27175 ( .A1(n39225), .A2(n37217), .ZN(n39697) );
  NAND2_X2 U27177 ( .A1(n11511), .A2(n29), .ZN(n39225) );
  BUF_X2 U27178 ( .I(n25754), .Z(n39226) );
  OR2_X1 U27180 ( .A1(n9333), .A2(n37100), .Z(n5335) );
  XOR2_X1 U27195 ( .A1(n4612), .A2(n39228), .Z(n7115) );
  XOR2_X1 U27197 ( .A1(n39229), .A2(n38385), .Z(n39228) );
  INV_X2 U27204 ( .I(n17937), .ZN(n39229) );
  NOR2_X2 U27210 ( .A1(n39230), .A2(n8763), .ZN(n33563) );
  OR2_X1 U27215 ( .A1(n9839), .A2(n31307), .Z(n13839) );
  BUF_X2 U27221 ( .I(n36595), .Z(n39231) );
  INV_X2 U27223 ( .I(n39232), .ZN(n39817) );
  XOR2_X1 U27229 ( .A1(n7929), .A2(n28925), .Z(n39233) );
  XOR2_X1 U27232 ( .A1(n8301), .A2(n8396), .Z(n8395) );
  NAND2_X1 U27237 ( .A1(n26098), .A2(n10764), .ZN(n4990) );
  NOR2_X2 U27246 ( .A1(n39236), .A2(n33376), .ZN(n3071) );
  NAND2_X2 U27251 ( .A1(n14737), .A2(n14735), .ZN(n28594) );
  NAND2_X2 U27252 ( .A1(n38220), .A2(n31664), .ZN(n14735) );
  NAND2_X1 U27254 ( .A1(n36530), .A2(n12289), .ZN(n20421) );
  OAI21_X2 U27255 ( .A1(n39237), .A2(n35290), .B(n9265), .ZN(n18872) );
  OAI21_X2 U27266 ( .A1(n25845), .A2(n25844), .B(n39238), .ZN(n32106) );
  NAND3_X2 U27283 ( .A1(n25842), .A2(n25954), .A3(n37966), .ZN(n39238) );
  NAND2_X2 U27284 ( .A1(n30833), .A2(n253), .ZN(n24444) );
  XOR2_X1 U27289 ( .A1(n12586), .A2(n36803), .Z(n26919) );
  NOR2_X1 U27292 ( .A1(n36361), .A2(n35455), .ZN(n21780) );
  NAND2_X2 U27293 ( .A1(n35362), .A2(n6424), .ZN(n36226) );
  AOI22_X2 U27297 ( .A1(n29349), .A2(n1062), .B1(n29348), .B2(n39240), .ZN(
        n31307) );
  OR2_X1 U27298 ( .A1(n807), .A2(n24266), .Z(n11196) );
  NOR2_X1 U27307 ( .A1(n29421), .A2(n32946), .ZN(n12054) );
  INV_X2 U27311 ( .I(n39241), .ZN(n5836) );
  XOR2_X1 U27312 ( .A1(n8083), .A2(n35920), .Z(n39241) );
  BUF_X2 U27314 ( .I(n33738), .Z(n39242) );
  AOI21_X2 U27317 ( .A1(n7986), .A2(n6064), .B(n35962), .ZN(n36450) );
  NOR2_X1 U27321 ( .A1(n18601), .A2(n29338), .ZN(n18671) );
  NAND2_X2 U27327 ( .A1(n12060), .A2(n31810), .ZN(n14858) );
  OAI21_X2 U27329 ( .A1(n28287), .A2(n28288), .B(n28161), .ZN(n32077) );
  XOR2_X1 U27335 ( .A1(n31240), .A2(n37222), .Z(n16318) );
  XOR2_X1 U27351 ( .A1(n24056), .A2(n24057), .Z(n14821) );
  XOR2_X1 U27352 ( .A1(n10722), .A2(n23794), .Z(n24057) );
  OAI21_X2 U27353 ( .A1(n39244), .A2(n39243), .B(n3619), .ZN(n19294) );
  OAI21_X1 U27354 ( .A1(n9385), .A2(n24732), .B(n35250), .ZN(n3792) );
  OR2_X1 U27355 ( .A1(n26688), .A2(n26665), .Z(n18357) );
  NAND2_X2 U27368 ( .A1(n34311), .A2(n113), .ZN(n39484) );
  XOR2_X1 U27375 ( .A1(n5225), .A2(n5226), .Z(n20613) );
  NAND2_X2 U27379 ( .A1(n23389), .A2(n4525), .ZN(n23234) );
  XOR2_X1 U27383 ( .A1(n30838), .A2(n39246), .Z(n820) );
  XOR2_X1 U27396 ( .A1(n25216), .A2(n25258), .Z(n39246) );
  XOR2_X1 U27407 ( .A1(n6681), .A2(n34351), .Z(n31840) );
  XOR2_X1 U27408 ( .A1(n11201), .A2(n22645), .Z(n37023) );
  NAND2_X2 U27411 ( .A1(n12567), .A2(n22162), .ZN(n11201) );
  NOR2_X2 U27418 ( .A1(n3685), .A2(n2336), .ZN(n10065) );
  XOR2_X1 U27419 ( .A1(n17326), .A2(n39247), .Z(n29424) );
  OAI21_X2 U27422 ( .A1(n25727), .A2(n16264), .B(n39273), .ZN(n10723) );
  OAI21_X1 U27435 ( .A1(n31555), .A2(n26609), .B(n39825), .ZN(n34642) );
  XOR2_X1 U27439 ( .A1(n25243), .A2(n29838), .Z(n9325) );
  NAND3_X2 U27444 ( .A1(n24766), .A2(n24767), .A3(n24768), .ZN(n25243) );
  NOR2_X1 U27445 ( .A1(n13524), .A2(n30283), .ZN(n13523) );
  XOR2_X1 U27448 ( .A1(n27665), .A2(n27835), .Z(n18512) );
  INV_X1 U27451 ( .I(n35256), .ZN(n39449) );
  XOR2_X1 U27458 ( .A1(n10002), .A2(n27462), .Z(n27985) );
  INV_X2 U27463 ( .I(n18257), .ZN(n19716) );
  NAND2_X2 U27466 ( .A1(n9569), .A2(n9570), .ZN(n18257) );
  NAND2_X2 U27480 ( .A1(n17917), .A2(n22891), .ZN(n33163) );
  OAI22_X2 U27481 ( .A1(n7537), .A2(n22920), .B1(n19945), .B2(n22682), .ZN(
        n22891) );
  INV_X1 U27484 ( .I(n15459), .ZN(n39252) );
  NAND2_X2 U27489 ( .A1(n39253), .A2(n14895), .ZN(n31986) );
  XOR2_X1 U27492 ( .A1(n6571), .A2(n19816), .Z(n6572) );
  NOR2_X2 U27494 ( .A1(n4400), .A2(n4401), .ZN(n6571) );
  NAND2_X2 U27501 ( .A1(n17096), .A2(n19976), .ZN(n4139) );
  OAI21_X2 U27511 ( .A1(n19975), .A2(n17001), .B(n39242), .ZN(n17096) );
  XOR2_X1 U27512 ( .A1(n39254), .A2(n34145), .Z(n34351) );
  XOR2_X1 U27523 ( .A1(n37593), .A2(n33308), .Z(n39254) );
  NOR2_X2 U27525 ( .A1(n6282), .A2(n2349), .ZN(n25424) );
  NAND2_X2 U27526 ( .A1(n24536), .A2(n19418), .ZN(n25682) );
  OAI21_X2 U27527 ( .A1(n24772), .A2(n24686), .B(n5401), .ZN(n39256) );
  AOI21_X2 U27528 ( .A1(n20316), .A2(n38797), .B(n39257), .ZN(n16859) );
  XOR2_X1 U27536 ( .A1(n7018), .A2(n26596), .Z(n26261) );
  NAND2_X2 U27546 ( .A1(n33517), .A2(n35568), .ZN(n33030) );
  AOI22_X2 U27550 ( .A1(n3949), .A2(n24467), .B1(n24466), .B2(n1280), .ZN(
        n39354) );
  NOR2_X2 U27554 ( .A1(n19566), .A2(n37259), .ZN(n24466) );
  NOR2_X1 U27558 ( .A1(n15299), .A2(n388), .ZN(n4638) );
  OAI22_X2 U27564 ( .A1(n22851), .A2(n22859), .B1(n5436), .B2(n383), .ZN(n388)
         );
  INV_X4 U27567 ( .I(n33277), .ZN(n39416) );
  XOR2_X1 U27571 ( .A1(n17563), .A2(n638), .Z(n2398) );
  XOR2_X1 U27575 ( .A1(n35654), .A2(n26595), .Z(n26358) );
  NOR2_X2 U27578 ( .A1(n4460), .A2(n6178), .ZN(n26595) );
  NOR2_X2 U27580 ( .A1(n25661), .A2(n19153), .ZN(n25383) );
  NAND2_X2 U27583 ( .A1(n32929), .A2(n32928), .ZN(n39260) );
  XOR2_X1 U27585 ( .A1(n23712), .A2(n23893), .Z(n23734) );
  NAND3_X2 U27588 ( .A1(n23408), .A2(n23407), .A3(n23406), .ZN(n23893) );
  BUF_X2 U27591 ( .I(n12617), .Z(n39261) );
  INV_X2 U27594 ( .I(n33786), .ZN(n1133) );
  NOR2_X2 U27595 ( .A1(n36686), .A2(n31156), .ZN(n36187) );
  XOR2_X1 U27596 ( .A1(n12854), .A2(n12855), .Z(n7865) );
  AND2_X1 U27599 ( .A1(n24586), .A2(n10980), .Z(n39505) );
  NOR2_X2 U27608 ( .A1(n28626), .A2(n28625), .ZN(n14712) );
  INV_X2 U27624 ( .I(n39263), .ZN(n25498) );
  XOR2_X1 U27626 ( .A1(n10153), .A2(n39694), .Z(n12835) );
  XOR2_X1 U27629 ( .A1(n6177), .A2(n7481), .Z(n10153) );
  NAND2_X2 U27632 ( .A1(n4823), .A2(n14848), .ZN(n8493) );
  NAND2_X2 U27634 ( .A1(n8160), .A2(n24233), .ZN(n39370) );
  NAND2_X2 U27640 ( .A1(n3869), .A2(n1609), .ZN(n24233) );
  NOR2_X2 U27651 ( .A1(n13988), .A2(n7236), .ZN(n39264) );
  NOR2_X2 U27653 ( .A1(n2832), .A2(n30656), .ZN(n26591) );
  XOR2_X1 U27654 ( .A1(n3893), .A2(n39267), .Z(n3937) );
  XOR2_X1 U27659 ( .A1(n11570), .A2(n1556), .Z(n39267) );
  NAND2_X1 U27667 ( .A1(n14587), .A2(n21391), .ZN(n16289) );
  NAND2_X2 U27672 ( .A1(n4001), .A2(n25361), .ZN(n39269) );
  NOR2_X2 U27686 ( .A1(n1676), .A2(n17207), .ZN(n22136) );
  NAND3_X1 U27691 ( .A1(n33747), .A2(n6235), .A3(n23574), .ZN(n32927) );
  NAND3_X2 U27692 ( .A1(n7825), .A2(n30631), .A3(n30276), .ZN(n23970) );
  INV_X2 U27693 ( .I(n39270), .ZN(n34073) );
  XOR2_X1 U27694 ( .A1(n19015), .A2(n31849), .Z(n39270) );
  XOR2_X1 U27700 ( .A1(n208), .A2(n32441), .Z(n17776) );
  XOR2_X1 U27707 ( .A1(n25153), .A2(n21259), .Z(n5629) );
  AOI22_X2 U27713 ( .A1(n11159), .A2(n3803), .B1(n11160), .B2(n121), .ZN(
        n39492) );
  XOR2_X1 U27714 ( .A1(n34409), .A2(n27806), .Z(n34408) );
  XOR2_X1 U27725 ( .A1(n12411), .A2(n7726), .Z(n32375) );
  XOR2_X1 U27730 ( .A1(n39272), .A2(n27791), .Z(n3157) );
  XOR2_X1 U27734 ( .A1(n13448), .A2(n20659), .Z(n39272) );
  XOR2_X1 U27738 ( .A1(n13700), .A2(n2392), .Z(n33582) );
  INV_X2 U27741 ( .I(n11601), .ZN(n7350) );
  INV_X2 U27750 ( .I(n14193), .ZN(n15737) );
  NAND2_X2 U27752 ( .A1(n8845), .A2(n21211), .ZN(n24683) );
  NAND2_X2 U27759 ( .A1(n34577), .A2(n13717), .ZN(n8858) );
  NAND2_X2 U27761 ( .A1(n36693), .A2(n8863), .ZN(n13717) );
  OR2_X1 U27763 ( .A1(n33939), .A2(n13453), .Z(n8847) );
  NOR2_X1 U27768 ( .A1(n33516), .A2(n28272), .ZN(n8308) );
  NAND3_X2 U27771 ( .A1(n31358), .A2(n25467), .A3(n25469), .ZN(n17329) );
  INV_X1 U27773 ( .I(n13554), .ZN(n12387) );
  XOR2_X1 U27775 ( .A1(n15348), .A2(n30626), .Z(n15410) );
  XOR2_X1 U27782 ( .A1(n24417), .A2(n9113), .Z(n34347) );
  NAND3_X2 U27783 ( .A1(n9416), .A2(n24493), .A3(n9418), .ZN(n9113) );
  XOR2_X1 U27788 ( .A1(n27817), .A2(n14325), .Z(n27818) );
  OAI21_X2 U27806 ( .A1(n18272), .A2(n18271), .B(n6127), .ZN(n39275) );
  XOR2_X1 U27815 ( .A1(n28970), .A2(n34787), .Z(n2218) );
  INV_X2 U27818 ( .I(n39277), .ZN(n807) );
  XOR2_X1 U27825 ( .A1(n39278), .A2(n1711), .Z(Ciphertext[103]) );
  BUF_X2 U27826 ( .I(n17412), .Z(n39280) );
  NOR3_X2 U27829 ( .A1(n39281), .A2(n32054), .A3(n34942), .ZN(n16929) );
  XOR2_X1 U27832 ( .A1(n25262), .A2(n39600), .Z(n39282) );
  XOR2_X1 U27833 ( .A1(n19374), .A2(n35468), .Z(n3393) );
  INV_X2 U27837 ( .I(n39285), .ZN(n5042) );
  NAND2_X1 U27838 ( .A1(n39287), .A2(n39286), .ZN(n5070) );
  NOR2_X1 U27839 ( .A1(n9235), .A2(n20960), .ZN(n39286) );
  XOR2_X1 U27842 ( .A1(n35163), .A2(n39288), .Z(n16110) );
  XOR2_X1 U27849 ( .A1(n38385), .A2(n23957), .Z(n39288) );
  BUF_X2 U27850 ( .I(n6145), .Z(n39289) );
  AOI21_X2 U27853 ( .A1(n12227), .A2(n28023), .B(n27711), .ZN(n27908) );
  XOR2_X1 U27866 ( .A1(n35076), .A2(n5867), .Z(n10251) );
  XOR2_X1 U27874 ( .A1(n24047), .A2(n23969), .Z(n23936) );
  NAND3_X2 U27877 ( .A1(n31786), .A2(n1034), .A3(n24425), .ZN(n39290) );
  OAI22_X2 U27878 ( .A1(n39292), .A2(n39291), .B1(n2326), .B2(n1529), .ZN(
        n33027) );
  INV_X2 U27879 ( .I(n35333), .ZN(n39291) );
  INV_X2 U27882 ( .I(n26038), .ZN(n39292) );
  NAND2_X2 U27885 ( .A1(n39293), .A2(n30817), .ZN(n15439) );
  NOR2_X2 U27886 ( .A1(n14508), .A2(n15134), .ZN(n39293) );
  NAND2_X1 U27889 ( .A1(n39294), .A2(n24963), .ZN(n4756) );
  XOR2_X1 U27891 ( .A1(n19035), .A2(n16771), .Z(n29119) );
  NAND3_X2 U27893 ( .A1(n20878), .A2(n28410), .A3(n104), .ZN(n19035) );
  NAND3_X2 U27896 ( .A1(n23248), .A2(n12094), .A3(n23270), .ZN(n39533) );
  BUF_X2 U27908 ( .I(n3977), .Z(n39296) );
  XOR2_X1 U27914 ( .A1(n23961), .A2(n8904), .Z(n5179) );
  XOR2_X1 U27915 ( .A1(n14393), .A2(n19835), .Z(n19472) );
  NAND2_X2 U27917 ( .A1(n7080), .A2(n14253), .ZN(n14393) );
  OAI21_X2 U27920 ( .A1(n36703), .A2(n20500), .B(n2338), .ZN(n28344) );
  INV_X2 U27922 ( .I(n253), .ZN(n24440) );
  OAI21_X2 U27923 ( .A1(n39301), .A2(n1133), .B(n39299), .ZN(n23377) );
  NOR2_X2 U27924 ( .A1(n31157), .A2(n33952), .ZN(n39302) );
  INV_X2 U27925 ( .I(n21144), .ZN(n32712) );
  OAI22_X2 U27928 ( .A1(n1076), .A2(n20010), .B1(n36197), .B2(n35469), .ZN(
        n28281) );
  NAND2_X2 U27930 ( .A1(n39414), .A2(n8262), .ZN(n8261) );
  XOR2_X1 U27941 ( .A1(n18049), .A2(n18048), .Z(n20070) );
  INV_X2 U27942 ( .I(n3977), .ZN(n35115) );
  NAND2_X2 U27946 ( .A1(n35036), .A2(n4098), .ZN(n3977) );
  XOR2_X1 U27948 ( .A1(n28976), .A2(n28975), .Z(n29907) );
  BUF_X2 U27960 ( .I(n10482), .Z(n39303) );
  OAI21_X1 U27968 ( .A1(n33369), .A2(n27385), .B(n1471), .ZN(n27384) );
  NAND2_X2 U27971 ( .A1(n10693), .A2(n10689), .ZN(n24529) );
  NAND2_X2 U27972 ( .A1(n6027), .A2(n39304), .ZN(n27672) );
  AOI22_X2 U27975 ( .A1(n4610), .A2(n33336), .B1(n33369), .B2(n13222), .ZN(
        n39304) );
  XOR2_X1 U27981 ( .A1(n6905), .A2(n6906), .Z(n19982) );
  NAND3_X1 U27982 ( .A1(n31534), .A2(n29237), .A3(n14933), .ZN(n39306) );
  NAND2_X2 U28007 ( .A1(n39307), .A2(n13419), .ZN(n32282) );
  OAI21_X2 U28011 ( .A1(n3733), .A2(n7434), .B(n2840), .ZN(n39307) );
  NAND3_X1 U28019 ( .A1(n781), .A2(n20173), .A3(n19594), .ZN(n32283) );
  INV_X2 U28020 ( .I(n35246), .ZN(n781) );
  INV_X2 U28021 ( .I(n39308), .ZN(n29430) );
  OAI21_X2 U28023 ( .A1(n15089), .A2(n14873), .B(n36275), .ZN(n39308) );
  INV_X2 U28025 ( .I(n20619), .ZN(n24473) );
  NAND2_X1 U28029 ( .A1(n39309), .A2(n20619), .ZN(n4666) );
  XOR2_X1 U28031 ( .A1(n20615), .A2(n23864), .Z(n20619) );
  INV_X2 U28033 ( .I(n16816), .ZN(n39309) );
  XOR2_X1 U28040 ( .A1(n29111), .A2(n20727), .Z(n16584) );
  XOR2_X1 U28041 ( .A1(n8729), .A2(n29167), .Z(n29111) );
  OAI21_X2 U28051 ( .A1(n2731), .A2(n934), .B(n24674), .ZN(n31124) );
  OAI22_X2 U28057 ( .A1(n36665), .A2(n31827), .B1(n1103), .B2(n26129), .ZN(
        n5684) );
  NAND2_X2 U28058 ( .A1(n5277), .A2(n12778), .ZN(n25894) );
  XOR2_X1 U28066 ( .A1(n36206), .A2(n17288), .Z(n18830) );
  XOR2_X1 U28072 ( .A1(n39311), .A2(n3304), .Z(n13745) );
  XOR2_X1 U28073 ( .A1(n3301), .A2(n3303), .Z(n39311) );
  NAND2_X1 U28083 ( .A1(n7300), .A2(n39485), .ZN(n36526) );
  NOR2_X1 U28092 ( .A1(n19992), .A2(n39312), .ZN(n14432) );
  XOR2_X1 U28100 ( .A1(n23780), .A2(n39314), .Z(n39460) );
  AOI21_X2 U28101 ( .A1(n13627), .A2(n34920), .B(n13626), .ZN(n5498) );
  XOR2_X1 U28104 ( .A1(n25217), .A2(n39315), .Z(n25220) );
  XOR2_X1 U28106 ( .A1(n11267), .A2(n6051), .Z(n6389) );
  AOI21_X2 U28107 ( .A1(n4825), .A2(n9024), .B(n7635), .ZN(n39318) );
  BUF_X4 U28108 ( .I(n542), .Z(n39739) );
  AND2_X1 U28110 ( .A1(n892), .A2(n14405), .Z(n31696) );
  XOR2_X1 U28111 ( .A1(n16066), .A2(n27709), .Z(n6395) );
  XOR2_X1 U28112 ( .A1(n6033), .A2(n27787), .Z(n27709) );
  XOR2_X1 U28122 ( .A1(n22429), .A2(n18153), .Z(n6369) );
  XOR2_X1 U28123 ( .A1(n39319), .A2(n12853), .Z(n33326) );
  XOR2_X1 U28124 ( .A1(n21007), .A2(n33650), .Z(n39319) );
  OR3_X1 U28125 ( .A1(n39061), .A2(n25696), .A3(n20838), .Z(n2495) );
  INV_X2 U28126 ( .I(n23571), .ZN(n30524) );
  NOR2_X2 U28127 ( .A1(n28771), .A2(n9290), .ZN(n888) );
  OAI21_X2 U28134 ( .A1(n5910), .A2(n37164), .B(n34668), .ZN(n9328) );
  INV_X2 U28135 ( .I(n39323), .ZN(n18467) );
  XOR2_X1 U28136 ( .A1(Plaintext[6]), .A2(Key[6]), .Z(n39323) );
  NOR2_X2 U28149 ( .A1(n11595), .A2(n11635), .ZN(n11594) );
  NAND2_X1 U28156 ( .A1(n24266), .A2(n24309), .ZN(n39324) );
  NAND2_X1 U28171 ( .A1(n11194), .A2(n24448), .ZN(n39325) );
  XOR2_X1 U28181 ( .A1(n18180), .A2(n34148), .Z(n4918) );
  NAND2_X2 U28182 ( .A1(n9140), .A2(n12152), .ZN(n18180) );
  XOR2_X1 U28219 ( .A1(n12014), .A2(n34214), .Z(n26303) );
  XOR2_X1 U28223 ( .A1(n12455), .A2(n12453), .Z(n28550) );
  NAND2_X2 U28224 ( .A1(n3844), .A2(n3843), .ZN(n28473) );
  NAND2_X2 U28234 ( .A1(n8157), .A2(n9585), .ZN(n9035) );
  AOI22_X2 U28244 ( .A1(n34585), .A2(n38724), .B1(n8046), .B2(n1630), .ZN(
        n9246) );
  AND2_X2 U28256 ( .A1(n16080), .A2(n7500), .Z(n25427) );
  INV_X2 U28266 ( .I(n39326), .ZN(n28093) );
  INV_X2 U28281 ( .I(n36634), .ZN(n25053) );
  XOR2_X1 U28284 ( .A1(n27758), .A2(n27647), .Z(n27713) );
  OAI21_X2 U28296 ( .A1(n39329), .A2(n10974), .B(n26773), .ZN(n39542) );
  NOR2_X2 U28298 ( .A1(n26866), .A2(n1089), .ZN(n39329) );
  OAI21_X2 U28307 ( .A1(n39330), .A2(n21494), .B(n21493), .ZN(n22019) );
  OAI21_X2 U28308 ( .A1(n35043), .A2(n21804), .B(n35042), .ZN(n39330) );
  XOR2_X1 U28309 ( .A1(n27433), .A2(n34050), .Z(n34650) );
  XOR2_X1 U28314 ( .A1(n2515), .A2(n39331), .Z(n30597) );
  XOR2_X1 U28316 ( .A1(n26411), .A2(n37206), .Z(n39331) );
  XOR2_X1 U28317 ( .A1(n3665), .A2(n21056), .Z(n21055) );
  XOR2_X1 U28333 ( .A1(n16524), .A2(n23861), .Z(n24055) );
  NAND3_X2 U28334 ( .A1(n10123), .A2(n36903), .A3(n18499), .ZN(n35331) );
  NOR2_X1 U28337 ( .A1(n1186), .A2(n5424), .ZN(n39334) );
  XOR2_X1 U28351 ( .A1(n2041), .A2(n39335), .Z(n35957) );
  INV_X1 U28352 ( .I(n39535), .ZN(n28128) );
  AND2_X1 U28353 ( .A1(n39535), .A2(n28093), .Z(n8788) );
  INV_X1 U28358 ( .I(n39336), .ZN(n36152) );
  NOR2_X2 U28359 ( .A1(n34656), .A2(n3336), .ZN(n34995) );
  OAI21_X1 U28386 ( .A1(n39337), .A2(n29210), .B(n30193), .ZN(n16535) );
  NOR2_X1 U28388 ( .A1(n17238), .A2(n35210), .ZN(n39337) );
  AOI21_X2 U28400 ( .A1(n12199), .A2(n38548), .B(n37132), .ZN(n3659) );
  BUF_X2 U28407 ( .I(n4034), .Z(n39338) );
  INV_X2 U28408 ( .I(n39339), .ZN(n640) );
  XOR2_X1 U28409 ( .A1(n9687), .A2(n699), .Z(n39339) );
  XNOR2_X1 U28410 ( .A1(n23930), .A2(n24005), .ZN(n39378) );
  XOR2_X1 U28421 ( .A1(n18807), .A2(n19761), .Z(n10083) );
  NOR2_X1 U28445 ( .A1(n13926), .A2(n29566), .ZN(n39340) );
  XOR2_X1 U28463 ( .A1(n15973), .A2(n39341), .Z(n23934) );
  XOR2_X1 U28471 ( .A1(n15971), .A2(n15972), .Z(n39341) );
  BUF_X2 U28474 ( .I(n14408), .Z(n39342) );
  NOR2_X2 U28476 ( .A1(n39343), .A2(n10019), .ZN(n10193) );
  NOR2_X2 U28488 ( .A1(n38166), .A2(n39345), .ZN(n39379) );
  NOR2_X2 U28489 ( .A1(n29444), .A2(n29595), .ZN(n39345) );
  NAND2_X2 U28493 ( .A1(n39616), .A2(n21529), .ZN(n17861) );
  XOR2_X1 U28522 ( .A1(n39346), .A2(n13288), .Z(n13799) );
  XOR2_X1 U28523 ( .A1(n29257), .A2(n13287), .Z(n39346) );
  INV_X2 U28526 ( .I(n39347), .ZN(n5976) );
  BUF_X2 U28531 ( .I(n32608), .Z(n39348) );
  OAI22_X2 U28536 ( .A1(n17716), .A2(n8711), .B1(n10062), .B2(n26030), .ZN(
        n8708) );
  NAND2_X2 U28538 ( .A1(n16407), .A2(n16867), .ZN(n17716) );
  NAND2_X2 U28539 ( .A1(n39349), .A2(n34257), .ZN(n11729) );
  NOR2_X2 U28556 ( .A1(n4656), .A2(n20549), .ZN(n39349) );
  XOR2_X1 U28561 ( .A1(n26384), .A2(n34648), .Z(n19448) );
  OR2_X1 U28572 ( .A1(n33455), .A2(n18741), .Z(n13371) );
  XOR2_X1 U28575 ( .A1(n26577), .A2(n36864), .Z(n33455) );
  BUF_X2 U28576 ( .I(n4574), .Z(n39350) );
  NOR2_X2 U28577 ( .A1(n11364), .A2(n31383), .ZN(n39808) );
  BUF_X2 U28582 ( .I(n950), .Z(n39351) );
  NAND2_X2 U28583 ( .A1(n34846), .A2(n39352), .ZN(n10223) );
  NOR2_X1 U28584 ( .A1(n15509), .A2(n939), .ZN(n18278) );
  NOR2_X2 U28592 ( .A1(n31751), .A2(n19706), .ZN(n15509) );
  AND3_X1 U28600 ( .A1(n28109), .A2(n8368), .A3(n33955), .Z(n15391) );
  NAND2_X2 U28601 ( .A1(n32469), .A2(n26108), .ZN(n26107) );
  XOR2_X1 U28602 ( .A1(n25010), .A2(n25011), .Z(n18705) );
  XOR2_X1 U28606 ( .A1(n25080), .A2(n35722), .Z(n25010) );
  BUF_X2 U28612 ( .I(n6067), .Z(n39355) );
  BUF_X2 U28616 ( .I(n22129), .Z(n39356) );
  XOR2_X1 U28630 ( .A1(n18498), .A2(n39358), .Z(n8897) );
  XOR2_X1 U28631 ( .A1(n35318), .A2(n39359), .Z(n39358) );
  INV_X1 U28632 ( .I(n30120), .ZN(n39359) );
  NAND2_X2 U28634 ( .A1(n33438), .A2(n12080), .ZN(n22401) );
  NAND2_X2 U28638 ( .A1(n12776), .A2(n27099), .ZN(n13703) );
  XOR2_X1 U28640 ( .A1(n35445), .A2(n39360), .Z(n31207) );
  XOR2_X1 U28641 ( .A1(n660), .A2(n17988), .Z(n39360) );
  XOR2_X1 U28642 ( .A1(n27842), .A2(n1467), .Z(n27469) );
  NAND2_X1 U28645 ( .A1(n39126), .A2(n17114), .ZN(n10721) );
  NAND2_X1 U28648 ( .A1(n32294), .A2(n23610), .ZN(n33356) );
  XOR2_X1 U28652 ( .A1(n32765), .A2(n7990), .Z(n24561) );
  AOI22_X2 U28654 ( .A1(n10464), .A2(n919), .B1(n21836), .B2(n19620), .ZN(
        n39361) );
  INV_X2 U28655 ( .I(n39362), .ZN(n2393) );
  XOR2_X1 U28679 ( .A1(n26363), .A2(n26184), .Z(n17935) );
  XOR2_X1 U28684 ( .A1(n39621), .A2(n20892), .Z(n21301) );
  NOR2_X2 U28688 ( .A1(n39367), .A2(n10354), .ZN(n7243) );
  NOR2_X2 U28693 ( .A1(n30282), .A2(n24691), .ZN(n39367) );
  XOR2_X1 U28697 ( .A1(n22712), .A2(n22564), .Z(n5609) );
  NAND2_X2 U28699 ( .A1(n6293), .A2(n32580), .ZN(n7323) );
  OR2_X1 U28704 ( .A1(n33249), .A2(n20694), .Z(n21482) );
  XOR2_X1 U28711 ( .A1(n9007), .A2(n39369), .Z(n9338) );
  XOR2_X1 U28726 ( .A1(n34901), .A2(n9005), .Z(n39369) );
  OR2_X1 U28727 ( .A1(n12447), .A2(n24328), .Z(n20227) );
  NOR2_X2 U28741 ( .A1(n21666), .A2(n21435), .ZN(n21836) );
  NAND2_X2 U28747 ( .A1(n34406), .A2(n34407), .ZN(n34405) );
  NAND2_X2 U28763 ( .A1(n32763), .A2(n10914), .ZN(n33993) );
  NAND2_X2 U28772 ( .A1(n39370), .A2(n23694), .ZN(n423) );
  OAI21_X2 U28784 ( .A1(n5621), .A2(n34030), .B(n5380), .ZN(n33461) );
  NAND2_X2 U28786 ( .A1(n21478), .A2(n19388), .ZN(n3618) );
  AOI21_X2 U28788 ( .A1(n3620), .A2(n33240), .B(n39372), .ZN(n3619) );
  NOR2_X2 U28793 ( .A1(n39373), .A2(n39381), .ZN(n39372) );
  NAND2_X2 U28799 ( .A1(n33579), .A2(n37107), .ZN(n39381) );
  AND2_X1 U28800 ( .A1(n894), .A2(n39374), .Z(n36469) );
  NAND3_X1 U28801 ( .A1(n1404), .A2(n29596), .A3(n14417), .ZN(n39374) );
  NAND2_X2 U28811 ( .A1(n1006), .A2(n924), .ZN(n7596) );
  AOI21_X2 U28814 ( .A1(n39377), .A2(n39376), .B(n20357), .ZN(n13922) );
  NAND2_X2 U28815 ( .A1(n4388), .A2(n19778), .ZN(n39376) );
  OAI21_X2 U28819 ( .A1(n2410), .A2(n14417), .B(n39379), .ZN(n29475) );
  NAND2_X1 U28820 ( .A1(n24963), .A2(n1530), .ZN(n39380) );
  NAND2_X2 U28821 ( .A1(n28478), .A2(n1196), .ZN(n28370) );
  NAND2_X2 U28826 ( .A1(n3533), .A2(n3534), .ZN(n28478) );
  NAND2_X2 U28829 ( .A1(n24261), .A2(n39381), .ZN(n24263) );
  XOR2_X1 U28833 ( .A1(n39383), .A2(n15700), .Z(Ciphertext[169]) );
  AOI22_X1 U28842 ( .A1(n29015), .A2(n18424), .B1(n30139), .B2(n30146), .ZN(
        n39383) );
  AOI22_X2 U28852 ( .A1(n27348), .A2(n33146), .B1(n27351), .B2(n27350), .ZN(
        n10366) );
  NOR2_X1 U28853 ( .A1(n8798), .A2(n8988), .ZN(n27348) );
  XOR2_X1 U28857 ( .A1(n39384), .A2(n28782), .Z(n36514) );
  XOR2_X1 U28859 ( .A1(n28780), .A2(n32465), .Z(n39384) );
  NOR2_X2 U28860 ( .A1(n26737), .A2(n17024), .ZN(n17023) );
  XOR2_X1 U28863 ( .A1(n25237), .A2(n25179), .Z(n25188) );
  XOR2_X1 U28870 ( .A1(n39385), .A2(n36456), .Z(n34828) );
  XOR2_X1 U28885 ( .A1(n39651), .A2(n19025), .Z(n39385) );
  NAND2_X2 U28887 ( .A1(n31048), .A2(n12936), .ZN(n39583) );
  NOR3_X2 U28893 ( .A1(n8803), .A2(n8804), .A3(n24794), .ZN(n32019) );
  NAND2_X2 U28894 ( .A1(n11614), .A2(n8944), .ZN(n28505) );
  INV_X1 U28895 ( .I(n26325), .ZN(n1237) );
  NOR2_X2 U28896 ( .A1(n20851), .A2(n20852), .ZN(n26325) );
  NAND2_X2 U28897 ( .A1(n39387), .A2(n31180), .ZN(n16260) );
  OAI21_X2 U28907 ( .A1(n29383), .A2(n17444), .B(n29382), .ZN(n39387) );
  XOR2_X1 U28908 ( .A1(n13852), .A2(n8939), .Z(n17250) );
  NAND2_X2 U28913 ( .A1(n34781), .A2(n8934), .ZN(n8939) );
  NAND2_X2 U28914 ( .A1(n39388), .A2(n4028), .ZN(n28622) );
  OAI21_X2 U28928 ( .A1(n14378), .A2(n17711), .B(n24180), .ZN(n364) );
  NAND2_X2 U28937 ( .A1(n14378), .A2(n24142), .ZN(n24180) );
  XOR2_X1 U28945 ( .A1(n29296), .A2(n28610), .Z(n29140) );
  NAND2_X2 U28946 ( .A1(n20314), .A2(n28331), .ZN(n29296) );
  OAI21_X2 U28947 ( .A1(n1095), .A2(n1094), .B(n1787), .ZN(n26728) );
  XOR2_X1 U28948 ( .A1(n17569), .A2(n30409), .Z(n15118) );
  XOR2_X1 U28958 ( .A1(n22453), .A2(n9116), .Z(n17569) );
  NAND2_X2 U28974 ( .A1(n31795), .A2(n26887), .ZN(n27703) );
  XOR2_X1 U28989 ( .A1(n21268), .A2(n182), .Z(n24224) );
  NAND2_X2 U28990 ( .A1(n33209), .A2(n33328), .ZN(n1010) );
  NAND2_X2 U28997 ( .A1(n8659), .A2(n14237), .ZN(n39391) );
  AOI21_X2 U29001 ( .A1(n36777), .A2(n7905), .B(n39394), .ZN(n34751) );
  INV_X2 U29034 ( .I(n14735), .ZN(n39394) );
  OR2_X1 U29035 ( .A1(n24432), .A2(n19576), .Z(n20458) );
  XOR2_X1 U29044 ( .A1(n359), .A2(n22476), .Z(n22754) );
  XOR2_X1 U29055 ( .A1(n39395), .A2(n33320), .Z(Ciphertext[66]) );
  AOI22_X1 U29064 ( .A1(n31284), .A2(n29570), .B1(n13442), .B2(n20701), .ZN(
        n39395) );
  NAND2_X2 U29065 ( .A1(n39396), .A2(n16737), .ZN(n7317) );
  OAI21_X2 U29079 ( .A1(n14625), .A2(n16739), .B(n31780), .ZN(n39396) );
  BUF_X2 U29085 ( .I(n28114), .Z(n39399) );
  OR2_X2 U29089 ( .A1(n19821), .A2(n19423), .Z(n39824) );
  INV_X2 U29090 ( .I(n39400), .ZN(n14103) );
  NOR2_X2 U29093 ( .A1(n5427), .A2(n1198), .ZN(n39400) );
  XOR2_X1 U29094 ( .A1(n11479), .A2(n29002), .Z(n16601) );
  XOR2_X1 U29096 ( .A1(n28971), .A2(n28896), .Z(n29002) );
  XOR2_X1 U29097 ( .A1(n31215), .A2(n14802), .Z(n20171) );
  XOR2_X1 U29103 ( .A1(n26572), .A2(n39032), .Z(n14802) );
  AOI21_X2 U29108 ( .A1(n34484), .A2(n11421), .B(n35988), .ZN(n614) );
  OAI22_X2 U29116 ( .A1(n4808), .A2(n16686), .B1(n26824), .B2(n14488), .ZN(
        n35988) );
  INV_X2 U29117 ( .I(n39403), .ZN(n39811) );
  XOR2_X1 U29118 ( .A1(n11498), .A2(n7341), .Z(n39403) );
  NAND2_X2 U29120 ( .A1(n19914), .A2(n1006), .ZN(n14807) );
  INV_X2 U29121 ( .I(n39404), .ZN(n24140) );
  XNOR2_X1 U29124 ( .A1(n35481), .A2(n35480), .ZN(n39404) );
  INV_X2 U29125 ( .I(n24879), .ZN(n39405) );
  BUF_X2 U29126 ( .I(n9231), .Z(n39407) );
  AND2_X1 U29133 ( .A1(n15566), .A2(n34764), .Z(n9293) );
  XOR2_X1 U29136 ( .A1(n25232), .A2(n21154), .Z(n2662) );
  XOR2_X1 U29140 ( .A1(n28955), .A2(n39409), .Z(n33890) );
  XOR2_X1 U29142 ( .A1(n28951), .A2(n37254), .Z(n39409) );
  XOR2_X1 U29145 ( .A1(n32647), .A2(n39780), .Z(n28130) );
  INV_X1 U29147 ( .I(n27728), .ZN(n39410) );
  XOR2_X1 U29153 ( .A1(n17417), .A2(n27779), .Z(n27728) );
  OAI21_X2 U29167 ( .A1(n26053), .A2(n34153), .B(n33395), .ZN(n1760) );
  INV_X2 U29173 ( .I(n39411), .ZN(n21767) );
  XNOR2_X1 U29174 ( .A1(Plaintext[132]), .A2(Key[132]), .ZN(n39411) );
  NAND2_X2 U29175 ( .A1(n3744), .A2(n3745), .ZN(n23938) );
  XOR2_X1 U29183 ( .A1(n8894), .A2(n27758), .Z(n10539) );
  XOR2_X1 U29198 ( .A1(n36706), .A2(n15393), .Z(n17726) );
  XOR2_X1 U29199 ( .A1(n31535), .A2(n27470), .Z(n27715) );
  AOI22_X2 U29202 ( .A1(n33278), .A2(n33277), .B1(n33276), .B2(n1400), .ZN(
        n39734) );
  NOR2_X1 U29207 ( .A1(n22068), .A2(n32318), .ZN(n39801) );
  NAND3_X2 U29227 ( .A1(n17236), .A2(n28052), .A3(n10443), .ZN(n17234) );
  XOR2_X1 U29237 ( .A1(n7069), .A2(n27662), .Z(n7068) );
  NAND2_X2 U29239 ( .A1(n33563), .A2(n21164), .ZN(n27662) );
  NAND2_X2 U29241 ( .A1(n34866), .A2(n1436), .ZN(n39419) );
  NOR2_X2 U29251 ( .A1(n21114), .A2(n8840), .ZN(n24737) );
  AOI21_X2 U29255 ( .A1(n24217), .A2(n24218), .B(n20839), .ZN(n21114) );
  NAND2_X2 U29263 ( .A1(n28435), .A2(n8321), .ZN(n35320) );
  NOR2_X2 U29264 ( .A1(n3634), .A2(n31036), .ZN(n36595) );
  XOR2_X1 U29265 ( .A1(n28940), .A2(n29818), .Z(n29168) );
  NOR2_X2 U29266 ( .A1(n31608), .A2(n16503), .ZN(n28940) );
  NAND2_X1 U29269 ( .A1(n34476), .A2(n39421), .ZN(n30512) );
  AOI22_X1 U29271 ( .A1(n30070), .A2(n30076), .B1(n3815), .B2(n6687), .ZN(
        n39421) );
  NOR2_X1 U29272 ( .A1(n3927), .A2(n6405), .ZN(n39422) );
  OR2_X1 U29273 ( .A1(n39769), .A2(n29059), .Z(n39432) );
  OR2_X1 U29277 ( .A1(n2798), .A2(n39401), .Z(n16842) );
  XOR2_X1 U29279 ( .A1(n4438), .A2(n39427), .Z(n5975) );
  XOR2_X1 U29281 ( .A1(n28839), .A2(n28838), .Z(n2547) );
  XOR2_X1 U29282 ( .A1(n16357), .A2(n29828), .Z(n28839) );
  OAI21_X2 U29283 ( .A1(n2453), .A2(n2454), .B(n39428), .ZN(n14272) );
  AOI22_X2 U29284 ( .A1(n34073), .A2(n14390), .B1(n19823), .B2(n17464), .ZN(
        n23154) );
  XOR2_X1 U29285 ( .A1(n26555), .A2(n39429), .Z(n157) );
  XOR2_X1 U29290 ( .A1(n26194), .A2(n8002), .Z(n39429) );
  NAND3_X1 U29292 ( .A1(n13876), .A2(n876), .A3(n27970), .ZN(n13875) );
  OAI21_X2 U29293 ( .A1(n26353), .A2(n17786), .B(n20190), .ZN(n4272) );
  OAI21_X2 U29303 ( .A1(n27587), .A2(n27306), .B(n4781), .ZN(n27040) );
  OR2_X2 U29305 ( .A1(n8000), .A2(n21152), .Z(n8311) );
  XOR2_X1 U29307 ( .A1(n24575), .A2(n13190), .Z(n31075) );
  NOR2_X1 U29315 ( .A1(n32981), .A2(n36454), .ZN(n15033) );
  XOR2_X1 U29317 ( .A1(n39430), .A2(n33674), .Z(n8454) );
  XOR2_X1 U29323 ( .A1(n29836), .A2(n39490), .Z(n39430) );
  NAND2_X1 U29324 ( .A1(n2866), .A2(n12081), .ZN(n39431) );
  INV_X2 U29328 ( .I(n39433), .ZN(n8042) );
  NAND2_X2 U29329 ( .A1(n6601), .A2(n6599), .ZN(n2792) );
  NOR2_X2 U29337 ( .A1(n29559), .A2(n6252), .ZN(n29551) );
  NOR2_X1 U29342 ( .A1(n39435), .A2(n12527), .ZN(n10992) );
  NOR2_X1 U29343 ( .A1(n39436), .A2(n29012), .ZN(n36013) );
  NOR2_X2 U29345 ( .A1(n14833), .A2(n5450), .ZN(n21449) );
  NAND2_X2 U29348 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  XOR2_X1 U29352 ( .A1(n6596), .A2(n39437), .Z(n6657) );
  XOR2_X1 U29353 ( .A1(n25200), .A2(n37234), .Z(n39437) );
  XOR2_X1 U29359 ( .A1(n39438), .A2(n26309), .Z(n13528) );
  XOR2_X1 U29372 ( .A1(n12933), .A2(n12429), .Z(n39438) );
  NAND2_X2 U29376 ( .A1(n38881), .A2(n17960), .ZN(n17959) );
  XOR2_X1 U29379 ( .A1(n12181), .A2(n12180), .Z(n12179) );
  NAND2_X2 U29381 ( .A1(n6926), .A2(n32778), .ZN(n9668) );
  OAI22_X2 U29391 ( .A1(n39439), .A2(n36207), .B1(n36225), .B2(n16672), .ZN(
        n31453) );
  AOI22_X2 U29397 ( .A1(n34389), .A2(n30196), .B1(n1755), .B2(n33861), .ZN(
        n39439) );
  XOR2_X1 U29399 ( .A1(n382), .A2(n25252), .Z(n10616) );
  OAI22_X2 U29402 ( .A1(n24731), .A2(n11712), .B1(n24730), .B2(n39157), .ZN(
        n382) );
  OAI21_X2 U29404 ( .A1(n39441), .A2(n39440), .B(n14331), .ZN(n15953) );
  INV_X2 U29419 ( .I(n23200), .ZN(n39440) );
  NAND2_X2 U29426 ( .A1(n11183), .A2(n11185), .ZN(n23814) );
  INV_X2 U29434 ( .I(n39444), .ZN(n25434) );
  XNOR2_X1 U29437 ( .A1(n25220), .A2(n39657), .ZN(n39444) );
  XOR2_X1 U29439 ( .A1(Plaintext[80]), .A2(Key[80]), .Z(n39680) );
  XOR2_X1 U29447 ( .A1(n10301), .A2(n38213), .Z(n27601) );
  NAND2_X2 U29454 ( .A1(n26648), .A2(n36953), .ZN(n27689) );
  OAI21_X1 U29455 ( .A1(n29358), .A2(n7376), .B(n29372), .ZN(n13646) );
  OAI21_X2 U29467 ( .A1(n14311), .A2(n8089), .B(n39445), .ZN(n13766) );
  INV_X2 U29468 ( .I(n22133), .ZN(n39445) );
  OAI22_X2 U29488 ( .A1(n9252), .A2(n22131), .B1(n31573), .B2(n35780), .ZN(
        n22133) );
  INV_X2 U29497 ( .I(n39446), .ZN(n8197) );
  XNOR2_X1 U29502 ( .A1(n7037), .A2(n7040), .ZN(n39446) );
  XOR2_X1 U29503 ( .A1(n9187), .A2(n14902), .Z(n39447) );
  NOR2_X2 U29504 ( .A1(n18536), .A2(n18537), .ZN(n24857) );
  NOR2_X2 U29510 ( .A1(n1420), .A2(n9668), .ZN(n4531) );
  AND2_X1 U29513 ( .A1(n39449), .A2(n26863), .Z(n14732) );
  NOR2_X1 U29515 ( .A1(n4633), .A2(n34987), .ZN(n10634) );
  XOR2_X1 U29521 ( .A1(n39450), .A2(n34092), .Z(n10835) );
  XOR2_X1 U29526 ( .A1(n33505), .A2(n15405), .Z(n39450) );
  OAI21_X2 U29534 ( .A1(n14125), .A2(n39451), .B(n6295), .ZN(n2696) );
  AND2_X1 U29535 ( .A1(n5751), .A2(n14124), .Z(n39451) );
  NOR2_X2 U29536 ( .A1(n31948), .A2(n39452), .ZN(n32601) );
  NOR3_X1 U29542 ( .A1(n22792), .A2(n33925), .A3(n33544), .ZN(n39452) );
  XOR2_X1 U29547 ( .A1(n21227), .A2(n32383), .Z(n32382) );
  XOR2_X1 U29549 ( .A1(n11383), .A2(n3448), .Z(n21227) );
  NOR2_X1 U29550 ( .A1(n34286), .A2(n34285), .ZN(n39453) );
  NAND2_X2 U29559 ( .A1(n33987), .A2(n34526), .ZN(n6791) );
  INV_X1 U29563 ( .I(n26290), .ZN(n34009) );
  XNOR2_X1 U29569 ( .A1(n26381), .A2(n26290), .ZN(n32175) );
  NAND2_X2 U29572 ( .A1(n4189), .A2(n25891), .ZN(n26290) );
  OAI21_X1 U29580 ( .A1(n39602), .A2(n30989), .B(n33455), .ZN(n26578) );
  INV_X2 U29582 ( .I(n39455), .ZN(n2707) );
  XOR2_X1 U29589 ( .A1(n21035), .A2(n35626), .Z(n39456) );
  NAND3_X2 U29590 ( .A1(n17811), .A2(n19069), .A3(n33101), .ZN(n31650) );
  NAND2_X2 U29591 ( .A1(n39457), .A2(n6463), .ZN(n23707) );
  NAND2_X1 U29592 ( .A1(n18618), .A2(n34012), .ZN(n39457) );
  NAND3_X1 U29597 ( .A1(n23172), .A2(n39418), .A3(n38752), .ZN(n20176) );
  OAI21_X2 U29603 ( .A1(n39599), .A2(n6731), .B(n25637), .ZN(n39458) );
  XOR2_X1 U29604 ( .A1(n39459), .A2(n20270), .Z(n20394) );
  XOR2_X1 U29605 ( .A1(n39460), .A2(n24074), .Z(n39459) );
  NAND2_X2 U29609 ( .A1(n39461), .A2(n39338), .ZN(n7) );
  NAND2_X2 U29612 ( .A1(n27300), .A2(n4033), .ZN(n39461) );
  XOR2_X1 U29613 ( .A1(n27751), .A2(n39462), .Z(n19009) );
  XOR2_X1 U29614 ( .A1(n9013), .A2(n35464), .Z(n39462) );
  NAND3_X2 U29617 ( .A1(n4439), .A2(n13982), .A3(n23509), .ZN(n11669) );
  NOR2_X2 U29621 ( .A1(n3659), .A2(n30934), .ZN(n13155) );
  INV_X2 U29625 ( .I(n39463), .ZN(n37052) );
  XNOR2_X1 U29628 ( .A1(n6924), .A2(n6922), .ZN(n39463) );
  NAND2_X2 U29629 ( .A1(n39517), .A2(n26778), .ZN(n2947) );
  OAI21_X2 U29636 ( .A1(n22683), .A2(n8339), .B(n17568), .ZN(n39464) );
  XOR2_X1 U29638 ( .A1(n35218), .A2(n8402), .Z(n39465) );
  NAND2_X2 U29640 ( .A1(n39466), .A2(n9504), .ZN(n12289) );
  NAND2_X1 U29643 ( .A1(n9506), .A2(n19769), .ZN(n39466) );
  XOR2_X1 U29644 ( .A1(n24942), .A2(n5845), .Z(n15531) );
  AOI21_X2 U29645 ( .A1(n37208), .A2(n23225), .B(n15074), .ZN(n15073) );
  XOR2_X1 U29648 ( .A1(n16368), .A2(n17462), .Z(n9122) );
  NAND2_X2 U29665 ( .A1(n7725), .A2(n9178), .ZN(n39514) );
  OAI22_X2 U29672 ( .A1(n19134), .A2(n32228), .B1(n11295), .B2(n23124), .ZN(
        n14343) );
  INV_X2 U29680 ( .I(n20897), .ZN(n32228) );
  XOR2_X1 U29681 ( .A1(n11382), .A2(n32847), .Z(n20897) );
  NAND2_X2 U29686 ( .A1(n2193), .A2(n8570), .ZN(n9116) );
  NOR2_X2 U29687 ( .A1(n36507), .A2(n26372), .ZN(n27389) );
  INV_X2 U29691 ( .I(n35164), .ZN(n18619) );
  NAND2_X1 U29692 ( .A1(n39467), .A2(n24395), .ZN(n24181) );
  INV_X2 U29701 ( .I(n8760), .ZN(n39467) );
  NAND2_X2 U29703 ( .A1(n24716), .A2(n14534), .ZN(n25226) );
  NOR3_X1 U29705 ( .A1(n20418), .A2(n23399), .A3(n36810), .ZN(n23320) );
  XOR2_X1 U29706 ( .A1(n39809), .A2(n36190), .Z(n22968) );
  NOR3_X2 U29708 ( .A1(n840), .A2(n949), .A3(n9743), .ZN(n33433) );
  AOI21_X2 U29710 ( .A1(n34720), .A2(n37477), .B(n31796), .ZN(n39469) );
  OR2_X2 U29713 ( .A1(n5104), .A2(n39470), .Z(n34475) );
  OAI22_X1 U29714 ( .A1(n21519), .A2(n19397), .B1(n21520), .B2(n21521), .ZN(
        n39470) );
  XOR2_X1 U29725 ( .A1(n15776), .A2(n27703), .Z(n27500) );
  XOR2_X1 U29733 ( .A1(n39471), .A2(n1051), .Z(Ciphertext[161]) );
  AOI22_X1 U29741 ( .A1(n30107), .A2(n12204), .B1(n18483), .B2(n16180), .ZN(
        n39471) );
  XNOR2_X1 U29750 ( .A1(n26356), .A2(n9151), .ZN(n6477) );
  INV_X2 U29752 ( .I(n39472), .ZN(n17692) );
  XOR2_X1 U29754 ( .A1(n39474), .A2(n7180), .Z(n20649) );
  XOR2_X1 U29755 ( .A1(n28984), .A2(n7182), .Z(n39474) );
  NAND2_X2 U29761 ( .A1(n11889), .A2(n20859), .ZN(n36798) );
  XOR2_X1 U29763 ( .A1(n39475), .A2(n16601), .Z(n16599) );
  XOR2_X1 U29767 ( .A1(n33387), .A2(n14487), .Z(n39475) );
  NAND3_X2 U29769 ( .A1(n23248), .A2(n22852), .A3(n23270), .ZN(n15491) );
  XOR2_X1 U29772 ( .A1(n39476), .A2(n16679), .Z(n6165) );
  XOR2_X1 U29775 ( .A1(n2585), .A2(n34188), .Z(n39476) );
  NAND2_X2 U29778 ( .A1(n3120), .A2(n24637), .ZN(n24635) );
  OAI21_X2 U29796 ( .A1(n15496), .A2(n15497), .B(n24230), .ZN(n24637) );
  NAND2_X1 U29811 ( .A1(n36474), .A2(n29124), .ZN(n36473) );
  XOR2_X1 U29819 ( .A1(n30687), .A2(n13205), .Z(n36552) );
  INV_X4 U29823 ( .I(n7852), .ZN(n24691) );
  INV_X2 U29834 ( .I(n30989), .ZN(n39477) );
  BUF_X2 U29839 ( .I(n14379), .Z(n39478) );
  INV_X2 U29845 ( .I(n39479), .ZN(n39830) );
  XOR2_X1 U29846 ( .A1(n36127), .A2(n28320), .Z(n39479) );
  XOR2_X1 U29847 ( .A1(n9085), .A2(n26480), .Z(n26572) );
  AOI21_X2 U29851 ( .A1(n8709), .A2(n8711), .B(n8708), .ZN(n9085) );
  NAND2_X2 U29866 ( .A1(n32596), .A2(n39481), .ZN(n18300) );
  OR2_X2 U29869 ( .A1(n7631), .A2(n23380), .Z(n30364) );
  OAI21_X2 U29870 ( .A1(n39711), .A2(n20981), .B(n4716), .ZN(n14115) );
  NOR2_X2 U29872 ( .A1(n26152), .A2(n26153), .ZN(n27164) );
  XOR2_X1 U29874 ( .A1(n31807), .A2(n27178), .Z(n1859) );
  NAND2_X2 U29876 ( .A1(n27165), .A2(n21272), .ZN(n27387) );
  NAND2_X2 U29879 ( .A1(n26445), .A2(n26446), .ZN(n27165) );
  NAND2_X1 U29884 ( .A1(n39483), .A2(n39482), .ZN(n10556) );
  NAND2_X1 U29885 ( .A1(n12661), .A2(n12660), .ZN(n39483) );
  NAND2_X1 U29890 ( .A1(n5976), .A2(n5975), .ZN(n36304) );
  NAND2_X2 U29892 ( .A1(n1222), .A2(n27197), .ZN(n27354) );
  XOR2_X1 U29894 ( .A1(n39487), .A2(n22581), .Z(n1758) );
  XOR2_X1 U29895 ( .A1(n4720), .A2(n22492), .Z(n39487) );
  BUF_X2 U29897 ( .I(n2980), .Z(n39488) );
  NOR3_X2 U29903 ( .A1(n25499), .A2(n32365), .A3(n3735), .ZN(n19240) );
  NAND2_X2 U29912 ( .A1(n22327), .A2(n4108), .ZN(n13163) );
  NAND2_X2 U29916 ( .A1(n27144), .A2(n9593), .ZN(n19455) );
  OAI21_X2 U29927 ( .A1(n16708), .A2(n26684), .B(n16707), .ZN(n27144) );
  XOR2_X1 U29942 ( .A1(n39631), .A2(n29092), .Z(n39490) );
  NAND3_X2 U29960 ( .A1(n13616), .A2(n13615), .A3(n22056), .ZN(n22439) );
  XOR2_X1 U29972 ( .A1(n39493), .A2(n36513), .Z(Ciphertext[141]) );
  NOR2_X1 U29975 ( .A1(n36848), .A2(n32531), .ZN(n39493) );
  NOR2_X2 U29978 ( .A1(n18304), .A2(n35253), .ZN(n2057) );
  OAI21_X2 U29985 ( .A1(n37192), .A2(n39494), .B(n1223), .ZN(n34890) );
  NOR2_X1 U29989 ( .A1(n14327), .A2(n27389), .ZN(n39494) );
  BUF_X2 U29995 ( .I(n18959), .Z(n39495) );
  NAND2_X2 U29996 ( .A1(n5093), .A2(n9141), .ZN(n16107) );
  NAND2_X2 U29997 ( .A1(n5498), .A2(n5496), .ZN(n7432) );
  AND2_X1 U30005 ( .A1(n28236), .A2(n39488), .Z(n27990) );
  XOR2_X1 U30006 ( .A1(n35208), .A2(n39497), .Z(n32516) );
  INV_X2 U30009 ( .I(n29833), .ZN(n39497) );
  OAI22_X2 U30014 ( .A1(n28499), .A2(n27941), .B1(n4697), .B2(n28498), .ZN(
        n29833) );
  AOI21_X1 U30016 ( .A1(n11398), .A2(n11397), .B(n1379), .ZN(n30577) );
  NOR2_X1 U30017 ( .A1(n20321), .A2(n37084), .ZN(n34061) );
  AOI22_X2 U30019 ( .A1(n15292), .A2(n18293), .B1(n11900), .B2(n8495), .ZN(
        n4823) );
  NOR2_X2 U30022 ( .A1(n14783), .A2(n21930), .ZN(n15292) );
  XOR2_X1 U30023 ( .A1(n11739), .A2(n24077), .Z(n12798) );
  OAI21_X2 U30030 ( .A1(n4960), .A2(n21014), .B(n12746), .ZN(n24077) );
  NAND3_X1 U30034 ( .A1(n7852), .A2(n5896), .A3(n39098), .ZN(n34881) );
  NAND2_X1 U30035 ( .A1(n6539), .A2(n6540), .ZN(n39498) );
  NAND2_X1 U30039 ( .A1(n6353), .A2(n31875), .ZN(n39499) );
  BUF_X2 U30041 ( .I(n14817), .Z(n39500) );
  XOR2_X1 U30044 ( .A1(n22444), .A2(n22500), .Z(n22544) );
  NAND2_X2 U30045 ( .A1(n22347), .A2(n22346), .ZN(n22444) );
  XOR2_X1 U30049 ( .A1(n22648), .A2(n22715), .Z(n13961) );
  NAND2_X2 U30054 ( .A1(n33155), .A2(n16712), .ZN(n23794) );
  OAI21_X1 U30056 ( .A1(n30145), .A2(n30134), .B(n18424), .ZN(n30135) );
  NAND2_X2 U30058 ( .A1(n18588), .A2(n18241), .ZN(n18424) );
  XOR2_X1 U30059 ( .A1(n27647), .A2(n10301), .Z(n27820) );
  NAND2_X2 U30064 ( .A1(n34493), .A2(n16045), .ZN(n27647) );
  NAND2_X2 U30067 ( .A1(n30958), .A2(n12659), .ZN(n35919) );
  XOR2_X1 U30068 ( .A1(n25005), .A2(n16192), .Z(n16191) );
  NAND3_X1 U30071 ( .A1(n27334), .A2(n1218), .A3(n35115), .ZN(n26846) );
  NAND2_X1 U30072 ( .A1(n8650), .A2(n7607), .ZN(n2130) );
  NAND2_X2 U30078 ( .A1(n39509), .A2(n15834), .ZN(n334) );
  INV_X2 U30079 ( .I(n39511), .ZN(n4306) );
  XOR2_X1 U30080 ( .A1(n291), .A2(n4204), .Z(n39512) );
  NAND2_X1 U30084 ( .A1(n29532), .A2(n29525), .ZN(n29524) );
  NAND2_X2 U30085 ( .A1(n36469), .A2(n10259), .ZN(n29532) );
  NAND2_X2 U30087 ( .A1(n34982), .A2(n9535), .ZN(n34977) );
  NAND2_X2 U30088 ( .A1(n3193), .A2(n18696), .ZN(n28546) );
  OR3_X1 U30092 ( .A1(n23610), .A2(n1627), .A3(n37088), .Z(n35397) );
  XOR2_X1 U30093 ( .A1(n39516), .A2(n2727), .Z(n5514) );
  XOR2_X1 U30095 ( .A1(n36915), .A2(n33007), .Z(n26779) );
  XOR2_X1 U30097 ( .A1(n20753), .A2(n22642), .Z(n11377) );
  XOR2_X1 U30100 ( .A1(n17189), .A2(n22552), .Z(n22642) );
  OAI22_X2 U30105 ( .A1(n26955), .A2(n8415), .B1(n31982), .B2(n8103), .ZN(
        n39517) );
  NOR2_X2 U30106 ( .A1(n20376), .A2(n19017), .ZN(n20375) );
  NAND2_X2 U30111 ( .A1(n39771), .A2(n37180), .ZN(n19017) );
  INV_X2 U30112 ( .I(n39519), .ZN(n36728) );
  XOR2_X1 U30116 ( .A1(n34178), .A2(n38190), .Z(n15304) );
  XOR2_X1 U30122 ( .A1(n27645), .A2(n31233), .Z(n34544) );
  XOR2_X1 U30123 ( .A1(n19405), .A2(n12985), .Z(n39520) );
  AOI21_X2 U30126 ( .A1(n28543), .A2(n37956), .B(n11474), .ZN(n29067) );
  XOR2_X1 U30127 ( .A1(n38584), .A2(n26556), .Z(n26483) );
  NAND2_X2 U30135 ( .A1(n33557), .A2(n30199), .ZN(n30213) );
  XOR2_X1 U30139 ( .A1(n39522), .A2(n19908), .Z(Ciphertext[182]) );
  BUF_X2 U30143 ( .I(n16502), .Z(n39523) );
  AOI22_X2 U30146 ( .A1(n39524), .A2(n28450), .B1(n18972), .B2(n18971), .ZN(
        n27957) );
  NOR2_X2 U30147 ( .A1(n35830), .A2(n12543), .ZN(n39524) );
  OAI21_X2 U30148 ( .A1(n12276), .A2(n12275), .B(n30048), .ZN(n39525) );
  AOI22_X2 U30152 ( .A1(n5678), .A2(n13705), .B1(n31512), .B2(n29979), .ZN(
        n29982) );
  XOR2_X1 U30154 ( .A1(n6325), .A2(n37194), .Z(n7201) );
  XNOR2_X1 U30165 ( .A1(n12267), .A2(n22790), .ZN(n6325) );
  INV_X2 U30169 ( .I(n32981), .ZN(n4573) );
  NAND2_X1 U30172 ( .A1(n19097), .A2(n18081), .ZN(n29911) );
  XOR2_X1 U30175 ( .A1(n28999), .A2(n15565), .Z(n39529) );
  OAI21_X2 U30176 ( .A1(n39530), .A2(n32719), .B(n20764), .ZN(n13278) );
  XOR2_X1 U30178 ( .A1(n26572), .A2(n26229), .Z(n26577) );
  BUF_X2 U30182 ( .I(n20158), .Z(n39537) );
  INV_X2 U30183 ( .I(n33323), .ZN(n36867) );
  NAND3_X2 U30185 ( .A1(n14498), .A2(n19080), .A3(n18872), .ZN(n33323) );
  NAND2_X2 U30186 ( .A1(n39539), .A2(n33392), .ZN(n36301) );
  NAND2_X2 U30188 ( .A1(n24778), .A2(n39540), .ZN(n39539) );
  NAND2_X2 U30189 ( .A1(n19593), .A2(n13300), .ZN(n24778) );
  NOR2_X1 U30190 ( .A1(n23128), .A2(n13688), .ZN(n7504) );
  NAND2_X1 U30201 ( .A1(n3725), .A2(n2944), .ZN(n5107) );
  BUF_X2 U30202 ( .I(n19849), .Z(n39541) );
  NOR2_X2 U30204 ( .A1(n12509), .A2(n11240), .ZN(n11434) );
  XOR2_X1 U30205 ( .A1(n39543), .A2(n29854), .Z(Ciphertext[116]) );
  NAND2_X1 U30207 ( .A1(n19872), .A2(n30616), .ZN(n39543) );
  NOR2_X1 U30212 ( .A1(n6191), .A2(n4272), .ZN(n27017) );
  XOR2_X1 U30213 ( .A1(n5308), .A2(n25242), .Z(n39544) );
  XOR2_X1 U30214 ( .A1(n23931), .A2(n23841), .Z(n23985) );
  NAND2_X2 U30218 ( .A1(n23369), .A2(n23368), .ZN(n23841) );
  XOR2_X1 U30219 ( .A1(n233), .A2(n10309), .Z(n25380) );
  INV_X1 U30224 ( .I(n31488), .ZN(n39660) );
  NAND2_X2 U30227 ( .A1(n20108), .A2(n15884), .ZN(n32377) );
  INV_X2 U30228 ( .I(n4381), .ZN(n25975) );
  NAND2_X2 U30231 ( .A1(n2626), .A2(n18787), .ZN(n4381) );
  XOR2_X1 U30238 ( .A1(n14231), .A2(n19849), .Z(n11899) );
  NAND3_X2 U30240 ( .A1(n6409), .A2(n6408), .A3(n9500), .ZN(n19849) );
  AOI21_X2 U30242 ( .A1(n39545), .A2(n32977), .B(n10228), .ZN(n18571) );
  NAND2_X2 U30243 ( .A1(n345), .A2(n11526), .ZN(n39545) );
  AND2_X1 U30245 ( .A1(n4272), .A2(n39546), .Z(n20709) );
  XOR2_X1 U30249 ( .A1(n39547), .A2(n27726), .Z(n31442) );
  XOR2_X1 U30251 ( .A1(n32015), .A2(n27823), .Z(n39547) );
  OAI21_X2 U30252 ( .A1(n26236), .A2(n30883), .B(n14157), .ZN(n26035) );
  NAND2_X2 U30253 ( .A1(n31994), .A2(n39375), .ZN(n14157) );
  NAND2_X2 U30254 ( .A1(n7695), .A2(n8770), .ZN(n5126) );
  XOR2_X1 U30256 ( .A1(n39549), .A2(n8856), .Z(n32893) );
  XOR2_X1 U30263 ( .A1(n7358), .A2(n31541), .Z(n39549) );
  XOR2_X1 U30267 ( .A1(n25268), .A2(n25188), .Z(n39550) );
  XOR2_X1 U30268 ( .A1(Plaintext[120]), .A2(Key[120]), .Z(n33999) );
  OR2_X1 U30271 ( .A1(n26833), .A2(n30853), .Z(n32941) );
  XNOR2_X1 U30274 ( .A1(n22736), .A2(n22714), .ZN(n36195) );
  NAND2_X2 U30275 ( .A1(n39551), .A2(n39586), .ZN(n6002) );
  NAND2_X2 U30277 ( .A1(n22101), .A2(n38830), .ZN(n22098) );
  NAND2_X2 U30279 ( .A1(n27235), .A2(n27436), .ZN(n27150) );
  NOR2_X2 U30281 ( .A1(n20492), .A2(n20493), .ZN(n6435) );
  NOR2_X2 U30282 ( .A1(n13501), .A2(n33433), .ZN(n6844) );
  XOR2_X1 U30289 ( .A1(n39552), .A2(n7664), .Z(n10006) );
  XOR2_X1 U30291 ( .A1(n27683), .A2(n27632), .Z(n27782) );
  XOR2_X1 U30295 ( .A1(n27504), .A2(n19758), .Z(n27505) );
  NAND2_X2 U30296 ( .A1(n15058), .A2(n14084), .ZN(n27504) );
  XOR2_X1 U30299 ( .A1(n39553), .A2(n16532), .Z(n5603) );
  XOR2_X1 U30301 ( .A1(n16531), .A2(n17117), .Z(n39553) );
  NOR2_X1 U30304 ( .A1(n16946), .A2(n27320), .ZN(n39554) );
  XOR2_X1 U30307 ( .A1(n39556), .A2(n30179), .Z(Ciphertext[178]) );
  NAND3_X2 U30311 ( .A1(n34903), .A2(n5422), .A3(n17168), .ZN(n39556) );
  NOR2_X2 U30312 ( .A1(n24350), .A2(n24349), .ZN(n5957) );
  OAI21_X2 U30313 ( .A1(n20022), .A2(n20021), .B(n39557), .ZN(n27446) );
  XOR2_X1 U30318 ( .A1(n6196), .A2(n6930), .Z(n28985) );
  NAND2_X2 U30325 ( .A1(n11911), .A2(n9625), .ZN(n6930) );
  XOR2_X1 U30335 ( .A1(n14231), .A2(n30179), .Z(n25221) );
  AOI22_X2 U30339 ( .A1(n8296), .A2(n1122), .B1(n14266), .B2(n36228), .ZN(
        n14231) );
  XOR2_X1 U30342 ( .A1(n39558), .A2(n22590), .Z(n36038) );
  XOR2_X1 U30344 ( .A1(n7560), .A2(n39559), .Z(n39558) );
  XOR2_X1 U30345 ( .A1(n39560), .A2(n10365), .Z(n20087) );
  XOR2_X1 U30351 ( .A1(n28332), .A2(n28333), .Z(n39560) );
  NAND2_X2 U30353 ( .A1(n3535), .A2(n31319), .ZN(n35664) );
  XOR2_X1 U30355 ( .A1(n20213), .A2(n39561), .Z(n35711) );
  NAND2_X2 U30358 ( .A1(n15377), .A2(n15378), .ZN(n20213) );
  NAND2_X2 U30361 ( .A1(n39562), .A2(n11258), .ZN(n15030) );
  XOR2_X1 U30363 ( .A1(n39563), .A2(n518), .Z(n12293) );
  XOR2_X1 U30365 ( .A1(n26591), .A2(n26305), .Z(n26210) );
  NOR2_X2 U30368 ( .A1(n5881), .A2(n5884), .ZN(n26305) );
  XOR2_X1 U30369 ( .A1(n11350), .A2(n11349), .Z(n11348) );
  INV_X4 U30370 ( .I(n19279), .ZN(n32802) );
  NAND2_X2 U30371 ( .A1(n4538), .A2(n31376), .ZN(n6560) );
  AND2_X1 U30375 ( .A1(n4386), .A2(n11415), .Z(n3820) );
  NAND2_X2 U30381 ( .A1(n9746), .A2(n36700), .ZN(n14833) );
  NAND2_X1 U30385 ( .A1(n27185), .A2(n4964), .ZN(n39566) );
  XOR2_X1 U30387 ( .A1(n27845), .A2(n16613), .Z(n27763) );
  NAND2_X2 U30388 ( .A1(n39567), .A2(n3819), .ZN(n4378) );
  NOR2_X1 U30389 ( .A1(n25813), .A2(n25936), .ZN(n25937) );
  XOR2_X1 U30390 ( .A1(n27853), .A2(n35610), .Z(n27856) );
  NAND2_X2 U30393 ( .A1(n39568), .A2(n35492), .ZN(n25887) );
  NAND2_X2 U30394 ( .A1(n19759), .A2(n8131), .ZN(n5465) );
  NOR2_X2 U30397 ( .A1(n30342), .A2(n9889), .ZN(n17925) );
  INV_X2 U30401 ( .I(n39570), .ZN(n9893) );
  NOR2_X1 U30402 ( .A1(n980), .A2(n37804), .ZN(n18018) );
  BUF_X2 U30404 ( .I(n23969), .Z(n39575) );
  AOI22_X2 U30405 ( .A1(n26694), .A2(n19455), .B1(n3783), .B2(n21144), .ZN(
        n10998) );
  INV_X2 U30406 ( .I(n39577), .ZN(n17314) );
  XOR2_X1 U30408 ( .A1(n27857), .A2(n20032), .Z(n39577) );
  AOI21_X1 U30409 ( .A1(n30113), .A2(n30119), .B(n39578), .ZN(n30116) );
  XOR2_X1 U30413 ( .A1(n27757), .A2(n10707), .Z(n5484) );
  BUF_X2 U30415 ( .I(n12649), .Z(n39579) );
  XOR2_X1 U30417 ( .A1(n9119), .A2(n7623), .Z(n9118) );
  OAI22_X1 U30418 ( .A1(n28364), .A2(n1193), .B1(n28365), .B2(n33460), .ZN(
        n5150) );
  XOR2_X1 U30419 ( .A1(n39580), .A2(n36087), .Z(n15903) );
  XOR2_X1 U30420 ( .A1(n6291), .A2(n32090), .Z(n39580) );
  XOR2_X1 U30423 ( .A1(n20987), .A2(n35317), .Z(n39600) );
  NAND2_X2 U30424 ( .A1(n17093), .A2(n16842), .ZN(n39581) );
  NOR2_X1 U30426 ( .A1(n7099), .A2(n36435), .ZN(n4459) );
  AND2_X1 U30431 ( .A1(n13686), .A2(n36355), .Z(n10564) );
  BUF_X2 U30432 ( .I(n840), .Z(n39584) );
  NAND2_X2 U30433 ( .A1(n39587), .A2(n13264), .ZN(n24732) );
  NAND2_X2 U30435 ( .A1(n39589), .A2(n32408), .ZN(n3967) );
  OAI22_X2 U30436 ( .A1(n22220), .A2(n22223), .B1(n8792), .B2(n22222), .ZN(
        n39589) );
  OAI21_X2 U30437 ( .A1(n14082), .A2(n6592), .B(n19589), .ZN(n14273) );
  XOR2_X1 U30440 ( .A1(n39590), .A2(n13654), .Z(n205) );
  XOR2_X1 U30441 ( .A1(n39591), .A2(n17000), .Z(n19473) );
  XOR2_X1 U30443 ( .A1(n14191), .A2(n15978), .Z(n34611) );
  OR2_X1 U30444 ( .A1(n22084), .A2(n2257), .Z(n39592) );
  XOR2_X1 U30445 ( .A1(n26181), .A2(n26399), .Z(n6134) );
  XOR2_X1 U30448 ( .A1(n26585), .A2(n19847), .Z(n26181) );
  AOI22_X2 U30451 ( .A1(n39593), .A2(n28641), .B1(n28640), .B2(n15447), .ZN(
        n20452) );
  OAI22_X2 U30452 ( .A1(n15447), .A2(n28639), .B1(n4369), .B2(n28637), .ZN(
        n39593) );
  NOR3_X2 U30461 ( .A1(n7086), .A2(n13444), .A3(n20041), .ZN(n6914) );
  NAND2_X2 U30469 ( .A1(n32741), .A2(n16406), .ZN(n39681) );
  NAND2_X1 U30471 ( .A1(n336), .A2(n27422), .ZN(n33799) );
  NAND2_X1 U30473 ( .A1(n23518), .A2(n23517), .ZN(n19283) );
  NOR2_X2 U30476 ( .A1(n22842), .A2(n22841), .ZN(n23517) );
  NAND2_X1 U30477 ( .A1(n18850), .A2(n8660), .ZN(n23312) );
  NOR2_X2 U30478 ( .A1(n34001), .A2(n27363), .ZN(n16482) );
  NAND2_X2 U30480 ( .A1(n18023), .A2(n18024), .ZN(n27363) );
  BUF_X2 U30481 ( .I(n26729), .Z(n39595) );
  NAND2_X2 U30482 ( .A1(n6282), .A2(n2349), .ZN(n33539) );
  INV_X1 U30483 ( .I(n22552), .ZN(n39630) );
  XOR2_X1 U30484 ( .A1(n26509), .A2(n26587), .Z(n39596) );
  OAI21_X1 U30486 ( .A1(n26864), .A2(n26952), .B(n39737), .ZN(n32176) );
  INV_X2 U30493 ( .I(n39597), .ZN(n27200) );
  NOR2_X2 U30494 ( .A1(n17072), .A2(n7424), .ZN(n39597) );
  BUF_X2 U30496 ( .I(n1230), .Z(n39598) );
  NOR2_X1 U30501 ( .A1(n11415), .A2(n4356), .ZN(n33276) );
  NAND2_X1 U30503 ( .A1(n22939), .A2(n10247), .ZN(n39601) );
  NAND2_X1 U30504 ( .A1(n29946), .A2(n11861), .ZN(n29841) );
  XOR2_X1 U30507 ( .A1(n25183), .A2(n39604), .Z(n34911) );
  XOR2_X1 U30508 ( .A1(n39320), .A2(n37109), .Z(n39604) );
  XOR2_X1 U30509 ( .A1(n27805), .A2(n13568), .Z(n13608) );
  NAND2_X2 U30516 ( .A1(n17893), .A2(n17891), .ZN(n12846) );
  AOI21_X2 U30517 ( .A1(n34143), .A2(n24605), .B(n33392), .ZN(n24607) );
  NOR2_X2 U30518 ( .A1(n39606), .A2(n21852), .ZN(n21856) );
  OAI21_X2 U30519 ( .A1(n1355), .A2(n693), .B(n6234), .ZN(n39606) );
  BUF_X2 U30521 ( .I(n17861), .Z(n39607) );
  INV_X2 U30524 ( .I(n39608), .ZN(n34160) );
  XOR2_X1 U30525 ( .A1(n1556), .A2(n17445), .Z(n39609) );
  NOR2_X2 U30528 ( .A1(n11469), .A2(n39610), .ZN(n35793) );
  INV_X2 U30532 ( .I(n28491), .ZN(n39610) );
  NAND2_X2 U30533 ( .A1(n18910), .A2(n16619), .ZN(n28491) );
  XOR2_X1 U30538 ( .A1(n36961), .A2(n26474), .Z(n39612) );
  XOR2_X1 U30541 ( .A1(n39613), .A2(n12556), .Z(n4752) );
  XOR2_X1 U30543 ( .A1(n8952), .A2(n18577), .Z(n39614) );
  XOR2_X1 U30545 ( .A1(n26503), .A2(n39615), .Z(n412) );
  XOR2_X1 U30546 ( .A1(n26504), .A2(n36333), .Z(n39615) );
  AOI22_X2 U30551 ( .A1(n39617), .A2(n9543), .B1(n23042), .B2(n22833), .ZN(
        n7024) );
  INV_X2 U30554 ( .I(n13485), .ZN(n39617) );
  NAND2_X2 U30555 ( .A1(n38329), .A2(n33431), .ZN(n13485) );
  NAND2_X2 U30556 ( .A1(n32), .A2(n3913), .ZN(n3907) );
  NAND2_X2 U30557 ( .A1(n8699), .A2(n8294), .ZN(n10221) );
  NOR2_X2 U30564 ( .A1(n4173), .A2(n4172), .ZN(n39624) );
  OAI21_X2 U30567 ( .A1(n21713), .A2(n19542), .B(n21652), .ZN(n39619) );
  XOR2_X1 U30568 ( .A1(n24560), .A2(n24563), .Z(n39621) );
  OAI22_X2 U30571 ( .A1(n39546), .A2(n27221), .B1(n38488), .B2(n39424), .ZN(
        n27297) );
  XOR2_X1 U30575 ( .A1(n382), .A2(n25215), .Z(n8920) );
  NAND2_X2 U30578 ( .A1(n13386), .A2(n19682), .ZN(n24342) );
  XOR2_X1 U30584 ( .A1(n11451), .A2(n33809), .Z(n11449) );
  NAND2_X2 U30589 ( .A1(n39623), .A2(n7565), .ZN(n6944) );
  NAND3_X1 U30593 ( .A1(n24205), .A2(n37264), .A3(n24206), .ZN(n39623) );
  NAND2_X2 U30594 ( .A1(n39624), .A2(n34461), .ZN(n35500) );
  NOR2_X2 U30596 ( .A1(n30825), .A2(n37139), .ZN(n3993) );
  OAI21_X2 U30606 ( .A1(n2058), .A2(n7036), .B(n35647), .ZN(n5634) );
  NAND2_X2 U30607 ( .A1(n6786), .A2(n6790), .ZN(n28758) );
  AOI22_X2 U30608 ( .A1(n23011), .A2(n5702), .B1(n4931), .B2(n1318), .ZN(
        n16416) );
  XOR2_X1 U30611 ( .A1(n9923), .A2(n17494), .Z(n17698) );
  NAND2_X1 U30613 ( .A1(n8027), .A2(n39629), .ZN(n33667) );
  NAND2_X1 U30614 ( .A1(n33786), .A2(n32366), .ZN(n39629) );
  INV_X2 U30616 ( .I(n23970), .ZN(n15336) );
  AND2_X1 U30617 ( .A1(n33738), .A2(n2153), .Z(n21991) );
  XOR2_X1 U30618 ( .A1(n22464), .A2(n11974), .Z(n15671) );
  NAND2_X2 U30621 ( .A1(n38282), .A2(n12029), .ZN(n31049) );
  OR2_X1 U30622 ( .A1(n11764), .A2(n11763), .Z(n39633) );
  XOR2_X1 U30625 ( .A1(n10767), .A2(n39634), .Z(n34223) );
  OAI21_X2 U30626 ( .A1(n35819), .A2(n35820), .B(n39635), .ZN(n27914) );
  NAND2_X2 U30630 ( .A1(n28133), .A2(n28229), .ZN(n39635) );
  XOR2_X1 U30632 ( .A1(n12183), .A2(n36952), .Z(n7273) );
  XOR2_X1 U30633 ( .A1(n9943), .A2(n14062), .Z(n5891) );
  INV_X2 U30634 ( .I(n39638), .ZN(n11636) );
  INV_X2 U30637 ( .I(n39639), .ZN(n693) );
  XNOR2_X1 U30638 ( .A1(Plaintext[36]), .A2(Key[36]), .ZN(n39639) );
  NAND2_X1 U30639 ( .A1(n39642), .A2(n39640), .ZN(n26640) );
  NAND2_X1 U30644 ( .A1(n39641), .A2(n26764), .ZN(n39640) );
  INV_X1 U30653 ( .I(n26763), .ZN(n39641) );
  NAND2_X1 U30658 ( .A1(n13393), .A2(n26763), .ZN(n39642) );
  OAI22_X2 U30659 ( .A1(n19893), .A2(n8082), .B1(n16067), .B2(n28390), .ZN(
        n39643) );
  XOR2_X1 U30660 ( .A1(n39644), .A2(n16091), .Z(n287) );
  XOR2_X1 U30663 ( .A1(n37256), .A2(n35249), .Z(n39644) );
  AOI22_X2 U30665 ( .A1(n2434), .A2(n12080), .B1(n2435), .B2(n8749), .ZN(
        n31476) );
  XOR2_X1 U30667 ( .A1(Key[37]), .A2(Plaintext[37]), .Z(n35161) );
  OAI21_X2 U30668 ( .A1(n39645), .A2(n15739), .B(n33045), .ZN(n6089) );
  NOR2_X2 U30670 ( .A1(n31283), .A2(n921), .ZN(n3699) );
  NAND2_X2 U30673 ( .A1(n31205), .A2(n26023), .ZN(n25771) );
  NAND3_X1 U30677 ( .A1(n9553), .A2(n3511), .A3(n17197), .ZN(n33805) );
  INV_X2 U30679 ( .I(n32153), .ZN(n33599) );
  XOR2_X1 U30680 ( .A1(n30458), .A2(n30963), .Z(n32153) );
  OAI21_X2 U30681 ( .A1(n451), .A2(n450), .B(n38172), .ZN(n5344) );
  NAND2_X2 U30683 ( .A1(n20959), .A2(n39649), .ZN(n13917) );
  AOI22_X2 U30684 ( .A1(n15193), .A2(n20155), .B1(n16871), .B2(n39258), .ZN(
        n39649) );
  NAND2_X1 U30686 ( .A1(n30844), .A2(n38197), .ZN(n39821) );
  NAND2_X2 U30687 ( .A1(n38206), .A2(n18042), .ZN(n18908) );
  XOR2_X1 U30688 ( .A1(n34894), .A2(n4305), .Z(n31370) );
  AOI22_X1 U30691 ( .A1(n29577), .A2(n20437), .B1(n31899), .B2(n29575), .ZN(
        n17113) );
  NOR2_X2 U30692 ( .A1(n1222), .A2(n27197), .ZN(n3783) );
  XOR2_X1 U30694 ( .A1(n19024), .A2(n39652), .Z(n39651) );
  INV_X2 U30700 ( .I(n26498), .ZN(n39652) );
  AOI22_X2 U30701 ( .A1(n35274), .A2(n20357), .B1(n3833), .B2(n19778), .ZN(
        n36886) );
  NAND2_X2 U30702 ( .A1(n22304), .A2(n3835), .ZN(n35274) );
  NAND2_X2 U30705 ( .A1(n6228), .A2(n37215), .ZN(n6727) );
  INV_X2 U30706 ( .I(n39653), .ZN(n39814) );
  XOR2_X1 U30707 ( .A1(n10275), .A2(n10278), .Z(n39653) );
  INV_X1 U30708 ( .I(n27581), .ZN(n19396) );
  XOR2_X1 U30711 ( .A1(n27581), .A2(n27669), .Z(n27552) );
  XOR2_X1 U30712 ( .A1(n6757), .A2(n17455), .Z(n21098) );
  NAND2_X2 U30714 ( .A1(n25596), .A2(n35821), .ZN(n6757) );
  XOR2_X1 U30716 ( .A1(n27661), .A2(n27662), .Z(n27840) );
  NOR2_X1 U30717 ( .A1(n17121), .A2(n30194), .ZN(n17120) );
  XOR2_X1 U30721 ( .A1(n15592), .A2(n39655), .Z(n30966) );
  XOR2_X1 U30722 ( .A1(n5407), .A2(n25219), .Z(n39657) );
  NOR2_X2 U30725 ( .A1(n21738), .A2(n19335), .ZN(n22295) );
  OAI21_X2 U30726 ( .A1(n2057), .A2(n20989), .B(n24382), .ZN(n16184) );
  NOR2_X2 U30728 ( .A1(n33834), .A2(n18407), .ZN(n9412) );
  OR2_X2 U30729 ( .A1(n8653), .A2(n8517), .Z(n21899) );
  AOI21_X2 U30731 ( .A1(n22288), .A2(n1687), .B(n1328), .ZN(n5556) );
  XNOR2_X1 U30732 ( .A1(n31151), .A2(n33166), .ZN(n39663) );
  OR2_X1 U30733 ( .A1(n33347), .A2(n19410), .Z(n27934) );
  AND2_X2 U30737 ( .A1(n17424), .A2(n17425), .Z(n29461) );
  OR2_X1 U30739 ( .A1(n32899), .A2(n4880), .Z(n31786) );
  BUF_X2 U30741 ( .I(n13285), .Z(n39666) );
  XOR2_X1 U30743 ( .A1(n26318), .A2(n26317), .Z(n39667) );
  XOR2_X1 U30746 ( .A1(n26491), .A2(n2545), .Z(n32954) );
  OR2_X1 U30747 ( .A1(n35431), .A2(n21802), .Z(n39668) );
  OR2_X1 U30752 ( .A1(n1230), .A2(n14962), .Z(n26865) );
  NOR2_X2 U30753 ( .A1(n3562), .A2(n21869), .ZN(n21867) );
  NAND2_X2 U30754 ( .A1(n12529), .A2(n34340), .ZN(n5383) );
  INV_X2 U30756 ( .I(n39669), .ZN(n34116) );
  NOR2_X2 U30759 ( .A1(n14037), .A2(n18303), .ZN(n39669) );
  NAND2_X2 U30761 ( .A1(n12252), .A2(n155), .ZN(n26359) );
  INV_X2 U30765 ( .I(n27233), .ZN(n39671) );
  BUF_X2 U30770 ( .I(n21683), .Z(n39672) );
  XOR2_X1 U30771 ( .A1(n2512), .A2(n23841), .Z(n23866) );
  NOR2_X2 U30776 ( .A1(n13537), .A2(n39673), .ZN(n13536) );
  INV_X1 U30781 ( .I(n39674), .ZN(n39673) );
  NAND2_X1 U30785 ( .A1(n10414), .A2(n37051), .ZN(n39674) );
  XOR2_X1 U30786 ( .A1(n26435), .A2(n39675), .Z(n26201) );
  XOR2_X1 U30790 ( .A1(n34469), .A2(n20600), .Z(n39675) );
  AOI21_X2 U30797 ( .A1(n33753), .A2(n39248), .B(n39676), .ZN(n14504) );
  INV_X2 U30799 ( .I(n18661), .ZN(n39676) );
  BUF_X2 U30800 ( .I(n8219), .Z(n39678) );
  XOR2_X1 U30802 ( .A1(n39679), .A2(n26385), .Z(n18390) );
  XOR2_X1 U30803 ( .A1(n9984), .A2(n26176), .Z(n39679) );
  INV_X1 U30806 ( .I(n39488), .ZN(n2302) );
  XOR2_X1 U30807 ( .A1(n2134), .A2(n31794), .Z(n2980) );
  XOR2_X1 U30811 ( .A1(n31162), .A2(n13934), .Z(n29347) );
  XOR2_X1 U30813 ( .A1(n29142), .A2(n19866), .Z(n16091) );
  OAI21_X2 U30814 ( .A1(n36517), .A2(n17447), .B(n8788), .ZN(n12885) );
  XOR2_X1 U30817 ( .A1(n5316), .A2(n5315), .Z(n6145) );
  XOR2_X1 U30819 ( .A1(n27805), .A2(n12507), .Z(n19989) );
  NOR2_X1 U30820 ( .A1(n32204), .A2(n19163), .ZN(n34287) );
  XOR2_X1 U30821 ( .A1(n11290), .A2(n11288), .Z(n11481) );
  NOR3_X2 U30822 ( .A1(n19549), .A2(n39656), .A3(n16305), .ZN(n7315) );
  AND2_X2 U30823 ( .A1(n29968), .A2(n18896), .Z(n29973) );
  XOR2_X1 U30827 ( .A1(n12884), .A2(n39683), .Z(n3770) );
  XOR2_X1 U30828 ( .A1(n27753), .A2(n37195), .Z(n39683) );
  XOR2_X1 U30831 ( .A1(n3081), .A2(n3632), .Z(n18806) );
  XOR2_X1 U30832 ( .A1(n22639), .A2(n22640), .Z(n34289) );
  NOR2_X2 U30836 ( .A1(n6348), .A2(n39684), .ZN(n6347) );
  OAI22_X2 U30837 ( .A1(n21560), .A2(n19397), .B1(n21477), .B2(n8597), .ZN(
        n39684) );
  NOR2_X2 U30839 ( .A1(n11759), .A2(n36800), .ZN(n24673) );
  NAND2_X2 U30841 ( .A1(n21796), .A2(n7047), .ZN(n31202) );
  NOR2_X1 U30844 ( .A1(n24156), .A2(n37267), .ZN(n24303) );
  NAND3_X2 U30852 ( .A1(n28452), .A2(n35793), .A3(n4523), .ZN(n29121) );
  XOR2_X1 U30860 ( .A1(n15336), .A2(n31775), .Z(n13736) );
  NAND2_X1 U30861 ( .A1(n31812), .A2(n3978), .ZN(n39721) );
  OAI21_X2 U30864 ( .A1(n37981), .A2(n28639), .B(n39355), .ZN(n30757) );
  AOI21_X1 U30869 ( .A1(n6323), .A2(n29479), .B(n29478), .ZN(n6322) );
  XOR2_X1 U30870 ( .A1(n36544), .A2(n9989), .Z(n26183) );
  OAI22_X2 U30871 ( .A1(n20296), .A2(n1253), .B1(n20295), .B2(n25448), .ZN(
        n39687) );
  NAND2_X2 U30872 ( .A1(n20979), .A2(n10896), .ZN(n29644) );
  XOR2_X1 U30873 ( .A1(n5026), .A2(n39688), .Z(n6596) );
  XOR2_X1 U30874 ( .A1(n6598), .A2(n518), .Z(n39688) );
  AND2_X1 U30875 ( .A1(n19605), .A2(n28132), .Z(n28223) );
  BUF_X2 U30876 ( .I(n29659), .Z(n39689) );
  NAND2_X1 U30877 ( .A1(n35686), .A2(n24874), .ZN(n9211) );
  XOR2_X1 U30878 ( .A1(n38154), .A2(n20454), .Z(n10117) );
  NAND2_X1 U30879 ( .A1(n6946), .A2(n21995), .ZN(n6949) );
  AOI22_X2 U30880 ( .A1(n20121), .A2(n25688), .B1(n25393), .B2(n25689), .ZN(
        n39690) );
  XOR2_X1 U30881 ( .A1(n34469), .A2(n20213), .Z(n26569) );
  INV_X2 U30882 ( .I(n19443), .ZN(n39691) );
  NAND2_X1 U30883 ( .A1(n28017), .A2(n39692), .ZN(n31799) );
  XNOR2_X1 U30884 ( .A1(n23955), .A2(n37842), .ZN(n39728) );
  OR2_X1 U30885 ( .A1(n17692), .A2(n34013), .Z(n23023) );
  NAND3_X1 U30886 ( .A1(n22917), .A2(n23163), .A3(n36095), .ZN(n11877) );
  NAND2_X1 U30887 ( .A1(n9165), .A2(n22250), .ZN(n9711) );
  NAND2_X2 U30888 ( .A1(n7759), .A2(n9495), .ZN(n9165) );
  XOR2_X1 U30889 ( .A1(n39693), .A2(n22648), .Z(n487) );
  XOR2_X1 U30890 ( .A1(n291), .A2(n32309), .Z(n39694) );
  XOR2_X1 U30891 ( .A1(n39695), .A2(n30063), .Z(Ciphertext[144]) );
  NAND2_X2 U30892 ( .A1(n39697), .A2(n11507), .ZN(n11541) );
  BUF_X2 U30893 ( .I(n6196), .Z(n39698) );
  XOR2_X1 U30894 ( .A1(n28969), .A2(n17250), .Z(n10136) );
  XOR2_X1 U30895 ( .A1(n38147), .A2(n29104), .Z(n28969) );
  INV_X2 U30896 ( .I(n36380), .ZN(n39699) );
  AOI21_X1 U30897 ( .A1(n21873), .A2(n21874), .B(n21872), .ZN(n21879) );
  AOI21_X2 U30898 ( .A1(n39700), .A2(n37183), .B(n1546), .ZN(n7097) );
  OAI22_X2 U30899 ( .A1(n27085), .A2(n14261), .B1(n33979), .B2(n38211), .ZN(
        n11590) );
  NAND2_X2 U30900 ( .A1(n39701), .A2(n29948), .ZN(n29979) );
  NAND2_X1 U30901 ( .A1(n13085), .A2(n1904), .ZN(n39701) );
  AOI22_X2 U30902 ( .A1(n21020), .A2(n156), .B1(n39702), .B2(n9514), .ZN(n3904) );
  OR2_X1 U30903 ( .A1(n22796), .A2(n35213), .Z(n23030) );
  XOR2_X1 U30904 ( .A1(n130), .A2(n12205), .Z(n22796) );
  NOR2_X2 U30905 ( .A1(n23389), .A2(n4525), .ZN(n9639) );
  BUF_X2 U30906 ( .I(n24300), .Z(n39703) );
  BUF_X2 U30907 ( .I(n8430), .Z(n39704) );
  XOR2_X1 U30908 ( .A1(n26457), .A2(n4918), .Z(n35923) );
  AOI22_X2 U30909 ( .A1(n21766), .A2(n16945), .B1(n9759), .B2(n21499), .ZN(
        n39705) );
  XNOR2_X1 U30910 ( .A1(n22620), .A2(n22731), .ZN(n22429) );
  OAI21_X2 U30911 ( .A1(n5085), .A2(n37001), .B(n39707), .ZN(n11443) );
  XOR2_X1 U30912 ( .A1(n39708), .A2(n7553), .Z(n10737) );
  XOR2_X1 U30913 ( .A1(n291), .A2(n12838), .Z(n39708) );
  BUF_X2 U30914 ( .I(n18081), .Z(n39709) );
  XOR2_X1 U30915 ( .A1(n39710), .A2(n10920), .Z(n36373) );
  BUF_X2 U30916 ( .I(n34644), .Z(n39711) );
  XOR2_X1 U30917 ( .A1(n33601), .A2(n29033), .Z(n18288) );
  NAND2_X2 U30918 ( .A1(n31486), .A2(n39768), .ZN(n29747) );
  NAND2_X2 U30919 ( .A1(n39715), .A2(n31904), .ZN(n8375) );
  NAND2_X1 U30920 ( .A1(n25305), .A2(n1535), .ZN(n39715) );
  XOR2_X1 U30921 ( .A1(n10380), .A2(n33789), .Z(n10379) );
  XOR2_X1 U30922 ( .A1(n16607), .A2(n16605), .Z(n17313) );
  XOR2_X1 U30923 ( .A1(n8755), .A2(n29293), .Z(n29307) );
  NAND2_X1 U30924 ( .A1(n4880), .A2(n10559), .ZN(n34374) );
  XOR2_X1 U30925 ( .A1(n27598), .A2(n39717), .Z(n27603) );
  XOR2_X1 U30926 ( .A1(n27597), .A2(n27596), .Z(n39717) );
  XOR2_X1 U30927 ( .A1(n22541), .A2(n39718), .Z(n36812) );
  XOR2_X1 U30928 ( .A1(n31504), .A2(n39630), .Z(n39718) );
  XOR2_X1 U30929 ( .A1(n33452), .A2(n23988), .Z(n24043) );
  NOR2_X2 U30930 ( .A1(n23016), .A2(n23015), .ZN(n23988) );
  XOR2_X1 U30931 ( .A1(n25145), .A2(n39720), .Z(n39719) );
  OAI21_X1 U30932 ( .A1(n15028), .A2(n14529), .B(n31534), .ZN(n15027) );
  NOR2_X2 U30933 ( .A1(n32061), .A2(n23458), .ZN(n23297) );
  NAND2_X2 U30934 ( .A1(n39721), .A2(n4741), .ZN(n9757) );
  NAND2_X2 U30935 ( .A1(n39722), .A2(n15710), .ZN(n8728) );
  BUF_X2 U30936 ( .I(n33509), .Z(n39723) );
  XOR2_X1 U30937 ( .A1(n4302), .A2(n25085), .Z(n4305) );
  XOR2_X1 U30938 ( .A1(n39726), .A2(n29091), .Z(n29199) );
  XOR2_X1 U30939 ( .A1(n7936), .A2(n6675), .Z(n39726) );
  OAI21_X2 U30940 ( .A1(n34682), .A2(n13270), .B(n35258), .ZN(n33255) );
  XOR2_X1 U30941 ( .A1(n36000), .A2(n39727), .Z(n8760) );
  XOR2_X1 U30942 ( .A1(n23836), .A2(n39728), .Z(n39727) );
  NAND2_X2 U30943 ( .A1(n35926), .A2(n20825), .ZN(n12793) );
  NAND3_X2 U30944 ( .A1(n32159), .A2(n9330), .A3(n8013), .ZN(n8660) );
  AOI21_X2 U30945 ( .A1(n37106), .A2(n13495), .B(n24630), .ZN(n11082) );
  XOR2_X1 U30946 ( .A1(n23947), .A2(n24006), .Z(n15904) );
  XOR2_X1 U30947 ( .A1(n27818), .A2(n31996), .Z(n27884) );
  XOR2_X1 U30948 ( .A1(n8920), .A2(n21252), .Z(n8922) );
  NAND3_X2 U30949 ( .A1(n4938), .A2(n24389), .A3(n24388), .ZN(n19359) );
  AOI21_X1 U30950 ( .A1(n32196), .A2(n31340), .B(n26215), .ZN(n16814) );
  NAND2_X2 U30951 ( .A1(n12365), .A2(n14349), .ZN(n17976) );
  NAND2_X1 U30952 ( .A1(n39732), .A2(n21756), .ZN(n13521) );
  INV_X2 U30953 ( .I(n39733), .ZN(n39827) );
  XOR2_X1 U30954 ( .A1(n19727), .A2(n9707), .Z(n39733) );
  AOI21_X2 U30955 ( .A1(n39735), .A2(n13030), .B(n24727), .ZN(n25186) );
  XOR2_X1 U30956 ( .A1(n11416), .A2(n34181), .Z(n11415) );
  BUF_X2 U30957 ( .I(n30284), .Z(n39737) );
  NAND2_X2 U30958 ( .A1(n39738), .A2(n7179), .ZN(n16238) );
  AND2_X1 U30959 ( .A1(n28339), .A2(n28400), .Z(n13401) );
  NAND2_X2 U30960 ( .A1(n33585), .A2(n33138), .ZN(n23426) );
  NAND3_X2 U30961 ( .A1(n39740), .A2(n30391), .A3(n28863), .ZN(n29687) );
  XOR2_X1 U30962 ( .A1(n39741), .A2(n27701), .Z(n6644) );
  XOR2_X1 U30963 ( .A1(n10057), .A2(n19612), .Z(n39741) );
  XOR2_X1 U30964 ( .A1(n29088), .A2(n12707), .Z(n6635) );
  NAND2_X2 U30965 ( .A1(n35776), .A2(n33686), .ZN(n12707) );
  XOR2_X1 U30966 ( .A1(n38041), .A2(n13147), .Z(n39743) );
  NAND2_X2 U30967 ( .A1(n36186), .A2(n36082), .ZN(n30282) );
  NAND2_X2 U30968 ( .A1(n4143), .A2(n121), .ZN(n15559) );
  XOR2_X1 U30969 ( .A1(n30819), .A2(n17328), .Z(n39744) );
  BUF_X2 U30970 ( .I(n29996), .Z(n39745) );
  XNOR2_X1 U30971 ( .A1(n17398), .A2(n6142), .ZN(n39783) );
  NAND3_X1 U30972 ( .A1(n27934), .A2(n32977), .A3(n28118), .ZN(n28347) );
  OAI21_X2 U30973 ( .A1(n22036), .A2(n22037), .B(n20388), .ZN(n22509) );
  NAND2_X2 U30974 ( .A1(n13241), .A2(n39746), .ZN(n5061) );
  NOR2_X2 U30975 ( .A1(n39747), .A2(n22091), .ZN(n22014) );
  NOR3_X1 U30976 ( .A1(n9685), .A2(n1678), .A3(n22204), .ZN(n39747) );
  AOI22_X2 U30977 ( .A1(n25364), .A2(n33114), .B1(n25366), .B2(n2576), .ZN(
        n39748) );
  AND2_X1 U30978 ( .A1(n16095), .A2(n33304), .Z(n39749) );
  NAND2_X2 U30979 ( .A1(n1116), .A2(n32868), .ZN(n3451) );
  NAND2_X2 U30980 ( .A1(n21565), .A2(n13472), .ZN(n2166) );
  XOR2_X1 U30981 ( .A1(n39750), .A2(n11284), .Z(n17533) );
  XOR2_X1 U30982 ( .A1(n39751), .A2(n9196), .Z(n7741) );
  XOR2_X1 U30983 ( .A1(n9195), .A2(n27795), .Z(n39751) );
  OR3_X1 U30984 ( .A1(n14369), .A2(n6106), .A3(n21301), .Z(n25604) );
  BUF_X2 U30985 ( .I(n20267), .Z(n39752) );
  XOR2_X1 U30986 ( .A1(n35654), .A2(n2443), .Z(n2714) );
  INV_X2 U30987 ( .I(n39753), .ZN(n19016) );
  XOR2_X1 U30988 ( .A1(Plaintext[44]), .A2(Key[44]), .Z(n39753) );
  OAI21_X2 U30989 ( .A1(n39754), .A2(n12405), .B(n26794), .ZN(n27304) );
  NOR2_X2 U30990 ( .A1(n3041), .A2(n37589), .ZN(n14429) );
  OAI21_X2 U30991 ( .A1(n39755), .A2(n9170), .B(n27893), .ZN(n28704) );
  AOI21_X2 U30992 ( .A1(n9168), .A2(n37015), .B(n28419), .ZN(n39755) );
  OAI21_X2 U30993 ( .A1(n12352), .A2(n12214), .B(n39757), .ZN(n17884) );
  AOI22_X2 U30994 ( .A1(n12213), .A2(n27306), .B1(n27585), .B2(n26791), .ZN(
        n39757) );
  INV_X2 U30995 ( .I(n39759), .ZN(n3452) );
  XNOR2_X1 U30996 ( .A1(n22596), .A2(n22607), .ZN(n39759) );
  OAI22_X1 U30997 ( .A1(n1021), .A2(n2830), .B1(n15575), .B2(n17624), .ZN(
        n2833) );
  INV_X2 U30998 ( .I(n23912), .ZN(n39760) );
  INV_X2 U30999 ( .I(n28590), .ZN(n39761) );
  INV_X2 U31000 ( .I(n5859), .ZN(n31375) );
  NAND3_X2 U31001 ( .A1(n5858), .A2(n5857), .A3(n12578), .ZN(n5859) );
  XOR2_X1 U31002 ( .A1(n39762), .A2(n1809), .Z(n1805) );
  XOR2_X1 U31003 ( .A1(n31012), .A2(n1807), .Z(n39762) );
  XOR2_X1 U31004 ( .A1(n17623), .A2(n39763), .Z(n14953) );
  XOR2_X1 U31005 ( .A1(n5208), .A2(n25115), .Z(n39763) );
  XOR2_X1 U31006 ( .A1(n39764), .A2(n22511), .Z(n5340) );
  INV_X2 U31007 ( .I(n20335), .ZN(n39764) );
  OAI22_X2 U31008 ( .A1(n18392), .A2(n12260), .B1(n12257), .B2(n14451), .ZN(
        n13409) );
  XOR2_X1 U31009 ( .A1(n3290), .A2(n31125), .Z(n755) );
  XOR2_X1 U31010 ( .A1(n26397), .A2(n13064), .Z(n39766) );
  XOR2_X1 U31011 ( .A1(n28918), .A2(n28919), .Z(n29903) );
  INV_X2 U31012 ( .I(n21644), .ZN(n21909) );
  NAND2_X2 U31013 ( .A1(n23608), .A2(n1637), .ZN(n3744) );
  OAI21_X2 U31014 ( .A1(n19869), .A2(n18850), .B(n32013), .ZN(n23608) );
  XOR2_X1 U31015 ( .A1(n22640), .A2(n39767), .Z(n35343) );
  XOR2_X1 U31016 ( .A1(n12393), .A2(n35081), .Z(n39767) );
  XOR2_X1 U31017 ( .A1(n23902), .A2(n18849), .Z(n6564) );
  NAND2_X1 U31018 ( .A1(n29194), .A2(n29815), .ZN(n39768) );
  NOR2_X1 U31019 ( .A1(n19041), .A2(n29973), .ZN(n29963) );
  INV_X2 U31020 ( .I(n10959), .ZN(n11861) );
  INV_X1 U31021 ( .I(n26458), .ZN(n26318) );
  XOR2_X1 U31022 ( .A1(n26458), .A2(n17760), .Z(n17759) );
  XOR2_X1 U31023 ( .A1(n26365), .A2(n5031), .Z(n26458) );
  INV_X2 U31024 ( .I(n19728), .ZN(n19575) );
  NAND2_X2 U31025 ( .A1(n39770), .A2(n23466), .ZN(n2319) );
  OR2_X1 U31026 ( .A1(n21546), .A2(n21871), .Z(n11918) );
  XOR2_X1 U31027 ( .A1(n4561), .A2(n4562), .Z(n4564) );
  XOR2_X1 U31028 ( .A1(n39772), .A2(n19616), .Z(Ciphertext[85]) );
  NAND2_X2 U31029 ( .A1(n9884), .A2(n11001), .ZN(n29683) );
  AOI22_X2 U31030 ( .A1(n16367), .A2(n33349), .B1(n32616), .B2(n23556), .ZN(
        n11529) );
  NAND2_X2 U31031 ( .A1(n39773), .A2(n35159), .ZN(n26161) );
  XOR2_X1 U31032 ( .A1(n12818), .A2(n39774), .Z(n4086) );
  XOR2_X1 U31033 ( .A1(n7055), .A2(n27739), .Z(n39774) );
  XOR2_X1 U31034 ( .A1(n39775), .A2(n34136), .Z(n35435) );
  NAND2_X2 U31035 ( .A1(n37104), .A2(n33561), .ZN(n13854) );
  INV_X2 U31036 ( .I(n1414), .ZN(n4284) );
  XOR2_X1 U31037 ( .A1(n39776), .A2(n8747), .Z(n7459) );
  XOR2_X1 U31038 ( .A1(n2283), .A2(n31909), .Z(n39776) );
  OAI21_X2 U31039 ( .A1(n2915), .A2(n12449), .B(n12448), .ZN(n6177) );
  NAND2_X2 U31040 ( .A1(n24342), .A2(n24341), .ZN(n30464) );
  XOR2_X1 U31041 ( .A1(n18310), .A2(n16905), .Z(n34518) );
  XOR2_X1 U31042 ( .A1(n31401), .A2(n24941), .Z(n39778) );
  XOR2_X1 U31043 ( .A1(n22677), .A2(n22622), .Z(n22592) );
  XOR2_X1 U31044 ( .A1(n23971), .A2(n23974), .Z(n11118) );
  XOR2_X1 U31045 ( .A1(n18300), .A2(n23783), .Z(n23971) );
  XOR2_X1 U31046 ( .A1(n6369), .A2(n39779), .Z(n19680) );
  XOR2_X1 U31047 ( .A1(n22372), .A2(n6368), .Z(n39779) );
  INV_X2 U31048 ( .I(n257), .ZN(n8264) );
  NAND2_X2 U31049 ( .A1(n15223), .A2(n16430), .ZN(n257) );
  XOR2_X1 U31050 ( .A1(n17651), .A2(n22383), .Z(n8856) );
  OAI21_X2 U31051 ( .A1(n37179), .A2(n3699), .B(n2121), .ZN(n9250) );
  XOR2_X1 U31052 ( .A1(n25145), .A2(n25143), .Z(n13260) );
  XOR2_X1 U31053 ( .A1(n25097), .A2(n25211), .Z(n25145) );
  NAND2_X1 U31054 ( .A1(n34957), .A2(n26929), .ZN(n26635) );
  NOR2_X2 U31055 ( .A1(n39477), .A2(n31546), .ZN(n26929) );
  XOR2_X1 U31056 ( .A1(n27474), .A2(n15726), .Z(n39780) );
  NOR2_X2 U31057 ( .A1(n840), .A2(n11003), .ZN(n31917) );
  AND3_X1 U31058 ( .A1(n22326), .A2(n39489), .A3(n4108), .Z(n36085) );
  NOR2_X1 U31059 ( .A1(n21687), .A2(n21688), .ZN(n21691) );
  INV_X2 U31060 ( .I(n9964), .ZN(n21687) );
  XOR2_X1 U31061 ( .A1(Plaintext[38]), .A2(Key[38]), .Z(n9964) );
  XOR2_X1 U31062 ( .A1(n39783), .A2(n9430), .Z(n36113) );
  XOR2_X1 U31063 ( .A1(n8473), .A2(n31591), .Z(n8472) );
  NAND2_X2 U31064 ( .A1(n16657), .A2(n16658), .ZN(n8473) );
  NAND2_X2 U31065 ( .A1(n39784), .A2(n33730), .ZN(n7506) );
  NAND2_X2 U31066 ( .A1(n2974), .A2(n2977), .ZN(n39784) );
  NAND2_X2 U31067 ( .A1(n39785), .A2(n10657), .ZN(n22119) );
  XOR2_X1 U31068 ( .A1(n22731), .A2(n31562), .Z(n17413) );
  NOR2_X2 U31069 ( .A1(n8503), .A2(n8504), .ZN(n31562) );
  XOR2_X1 U31070 ( .A1(n10520), .A2(n30094), .Z(n642) );
  XOR2_X1 U31071 ( .A1(n39790), .A2(n17834), .Z(n17838) );
  XOR2_X1 U31072 ( .A1(n18600), .A2(n25250), .Z(n39790) );
  XOR2_X1 U31073 ( .A1(n39791), .A2(n14505), .Z(n779) );
  XOR2_X1 U31074 ( .A1(n1324), .A2(n39792), .Z(n39791) );
  INV_X2 U31075 ( .I(n8552), .ZN(n39792) );
  NOR3_X2 U31076 ( .A1(n16845), .A2(n14432), .A3(n29640), .ZN(n19318) );
  XOR2_X1 U31077 ( .A1(n32646), .A2(n1664), .Z(n9511) );
  NOR2_X2 U31078 ( .A1(n31966), .A2(n28109), .ZN(n39794) );
  INV_X1 U31079 ( .I(n28240), .ZN(n39795) );
  BUF_X2 U31080 ( .I(n7728), .Z(n39797) );
  XOR2_X1 U31081 ( .A1(n5279), .A2(n37197), .Z(n12283) );
  XOR2_X1 U31082 ( .A1(n22741), .A2(n1324), .Z(n5279) );
  NOR2_X2 U31083 ( .A1(n7391), .A2(n19813), .ZN(n15635) );
  INV_X2 U31084 ( .I(n39799), .ZN(n7391) );
  NOR2_X2 U31085 ( .A1(n733), .A2(n33948), .ZN(n39799) );
  OR2_X1 U31086 ( .A1(n35757), .A2(n7459), .Z(n8819) );
  XOR2_X1 U31087 ( .A1(n35542), .A2(n14608), .Z(n35757) );
  NAND2_X2 U31088 ( .A1(n10152), .A2(n20313), .ZN(n24162) );
  OAI22_X1 U31089 ( .A1(n2866), .A2(n39392), .B1(n19544), .B2(n29059), .ZN(
        n15492) );
  NOR2_X2 U31090 ( .A1(n7789), .A2(n30240), .ZN(n2866) );
  NAND2_X2 U31091 ( .A1(n20875), .A2(n39802), .ZN(n26089) );
  OAI21_X2 U31092 ( .A1(n10532), .A2(n17282), .B(n7236), .ZN(n39802) );
  OR2_X1 U31093 ( .A1(n35216), .A2(n32775), .Z(n18207) );
  NAND2_X2 U31094 ( .A1(n4083), .A2(n35551), .ZN(n16672) );
  OAI21_X2 U31095 ( .A1(n24187), .A2(n13167), .B(n10659), .ZN(n36664) );
  AOI22_X2 U31096 ( .A1(n1133), .A2(n7885), .B1(n7886), .B2(n23504), .ZN(n7884) );
  NAND2_X1 U31097 ( .A1(n27269), .A2(n35990), .ZN(n20377) );
  XOR2_X1 U31098 ( .A1(n39807), .A2(n33695), .Z(n20974) );
  XOR2_X1 U31099 ( .A1(n34489), .A2(n26513), .Z(n39807) );
  OAI22_X2 U31100 ( .A1(n39808), .A2(n34790), .B1(n8342), .B2(n21995), .ZN(
        n6893) );
  XOR2_X1 U31101 ( .A1(n17569), .A2(n38216), .Z(n39809) );
  INV_X2 U31102 ( .I(n7828), .ZN(n21239) );
  INV_X2 U31103 ( .I(n17564), .ZN(n23190) );
  INV_X1 U31104 ( .I(n38851), .ZN(n22964) );
  INV_X2 U31105 ( .I(n22853), .ZN(n14817) );
  OR2_X1 U31106 ( .A1(n4600), .A2(n31611), .Z(n39813) );
  AND2_X1 U31107 ( .A1(n18907), .A2(n18402), .Z(n39818) );
  BUF_X2 U31108 ( .I(n19223), .Z(n14082) );
  INV_X2 U31109 ( .I(n9751), .ZN(n36708) );
  XNOR2_X1 U31110 ( .A1(n30910), .A2(n13260), .ZN(n39820) );
  BUF_X2 U31111 ( .I(n6145), .Z(n5314) );
  OAI22_X2 U31112 ( .A1(n16073), .A2(n34436), .B1(n16072), .B2(n35160), .ZN(
        n35207) );
  AOI22_X2 U31113 ( .A1(n26097), .A2(n39351), .B1(n32748), .B2(n32747), .ZN(
        n35238) );
  XNOR2_X1 U31114 ( .A1(n15077), .A2(n15453), .ZN(n39823) );
  INV_X2 U31115 ( .I(n28125), .ZN(n10836) );
  OAI21_X2 U31116 ( .A1(n5160), .A2(n5158), .B(n31932), .ZN(n6067) );
  INV_X2 U31117 ( .I(n13927), .ZN(n18061) );
  INV_X2 U31118 ( .I(n3845), .ZN(n31888) );
  INV_X2 U31119 ( .I(n34325), .ZN(n777) );
  INV_X2 U31120 ( .I(n16803), .ZN(n967) );
  XNOR2_X1 U31121 ( .A1(n2996), .A2(n32092), .ZN(n39828) );
  INV_X2 U31122 ( .I(n29184), .ZN(n35551) );
endmodule


module SPEEDY_Top ( clk, Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFFSNQ_X1 \reg_in_reg[190]  ( .D(Plaintext[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[190]) );
  DFFSNQ_X1 \reg_in_reg[189]  ( .D(Plaintext[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[189]) );
  DFFSNQ_X1 \reg_in_reg[188]  ( .D(Plaintext[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[188]) );
  DFFSNQ_X1 \reg_in_reg[187]  ( .D(Plaintext[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[187]) );
  DFFSNQ_X1 \reg_in_reg[186]  ( .D(Plaintext[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[186]) );
  DFFSNQ_X1 \reg_in_reg[185]  ( .D(Plaintext[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[185]) );
  DFFSNQ_X1 \reg_in_reg[184]  ( .D(Plaintext[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[184]) );
  DFFSNQ_X1 \reg_in_reg[183]  ( .D(Plaintext[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[183]) );
  DFFSNQ_X1 \reg_in_reg[182]  ( .D(Plaintext[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[182]) );
  DFFSNQ_X1 \reg_in_reg[181]  ( .D(Plaintext[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[181]) );
  DFFSNQ_X1 \reg_in_reg[180]  ( .D(Plaintext[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[180]) );
  DFFSNQ_X1 \reg_in_reg[179]  ( .D(Plaintext[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[179]) );
  DFFSNQ_X1 \reg_in_reg[178]  ( .D(Plaintext[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[178]) );
  DFFSNQ_X1 \reg_in_reg[177]  ( .D(Plaintext[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[177]) );
  DFFSNQ_X1 \reg_in_reg[176]  ( .D(Plaintext[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[176]) );
  DFFSNQ_X1 \reg_in_reg[175]  ( .D(Plaintext[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[175]) );
  DFFSNQ_X1 \reg_in_reg[174]  ( .D(Plaintext[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[174]) );
  DFFSNQ_X1 \reg_in_reg[173]  ( .D(Plaintext[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[173]) );
  DFFSNQ_X1 \reg_in_reg[172]  ( .D(Plaintext[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[172]) );
  DFFSNQ_X1 \reg_in_reg[171]  ( .D(Plaintext[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[171]) );
  DFFSNQ_X1 \reg_in_reg[170]  ( .D(Plaintext[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[170]) );
  DFFSNQ_X1 \reg_in_reg[168]  ( .D(Plaintext[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[168]) );
  DFFSNQ_X1 \reg_in_reg[167]  ( .D(Plaintext[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[167]) );
  DFFSNQ_X1 \reg_in_reg[166]  ( .D(Plaintext[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[166]) );
  DFFSNQ_X1 \reg_in_reg[165]  ( .D(Plaintext[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[165]) );
  DFFSNQ_X1 \reg_in_reg[164]  ( .D(Plaintext[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[164]) );
  DFFSNQ_X1 \reg_in_reg[163]  ( .D(Plaintext[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[163]) );
  DFFSNQ_X1 \reg_in_reg[162]  ( .D(Plaintext[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[162]) );
  DFFSNQ_X1 \reg_in_reg[161]  ( .D(Plaintext[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[161]) );
  DFFSNQ_X1 \reg_in_reg[160]  ( .D(Plaintext[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[160]) );
  DFFSNQ_X1 \reg_in_reg[159]  ( .D(Plaintext[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[159]) );
  DFFSNQ_X1 \reg_in_reg[158]  ( .D(Plaintext[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[158]) );
  DFFSNQ_X1 \reg_in_reg[157]  ( .D(Plaintext[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[157]) );
  DFFSNQ_X1 \reg_in_reg[156]  ( .D(Plaintext[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[156]) );
  DFFSNQ_X1 \reg_in_reg[155]  ( .D(Plaintext[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[155]) );
  DFFSNQ_X1 \reg_in_reg[154]  ( .D(Plaintext[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[154]) );
  DFFSNQ_X1 \reg_in_reg[153]  ( .D(Plaintext[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[153]) );
  DFFSNQ_X1 \reg_in_reg[152]  ( .D(Plaintext[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[152]) );
  DFFSNQ_X1 \reg_in_reg[151]  ( .D(Plaintext[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[151]) );
  DFFSNQ_X1 \reg_in_reg[150]  ( .D(Plaintext[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[150]) );
  DFFSNQ_X1 \reg_in_reg[149]  ( .D(Plaintext[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[149]) );
  DFFSNQ_X1 \reg_in_reg[148]  ( .D(Plaintext[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[148]) );
  DFFSNQ_X1 \reg_in_reg[147]  ( .D(Plaintext[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[147]) );
  DFFSNQ_X1 \reg_in_reg[145]  ( .D(Plaintext[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[145]) );
  DFFSNQ_X1 \reg_in_reg[144]  ( .D(Plaintext[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[144]) );
  DFFSNQ_X1 \reg_in_reg[143]  ( .D(Plaintext[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[143]) );
  DFFSNQ_X1 \reg_in_reg[142]  ( .D(Plaintext[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[142]) );
  DFFSNQ_X1 \reg_in_reg[141]  ( .D(Plaintext[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[141]) );
  DFFSNQ_X1 \reg_in_reg[139]  ( .D(Plaintext[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[139]) );
  DFFSNQ_X1 \reg_in_reg[138]  ( .D(Plaintext[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[138]) );
  DFFSNQ_X1 \reg_in_reg[137]  ( .D(Plaintext[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[137]) );
  DFFSNQ_X1 \reg_in_reg[136]  ( .D(Plaintext[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[136]) );
  DFFSNQ_X1 \reg_in_reg[135]  ( .D(Plaintext[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[135]) );
  DFFSNQ_X1 \reg_in_reg[134]  ( .D(Plaintext[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[134]) );
  DFFSNQ_X1 \reg_in_reg[133]  ( .D(Plaintext[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[133]) );
  DFFSNQ_X1 \reg_in_reg[132]  ( .D(Plaintext[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[132]) );
  DFFSNQ_X1 \reg_in_reg[131]  ( .D(Plaintext[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[131]) );
  DFFSNQ_X1 \reg_in_reg[130]  ( .D(Plaintext[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[130]) );
  DFFSNQ_X1 \reg_in_reg[129]  ( .D(Plaintext[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[129]) );
  DFFSNQ_X1 \reg_in_reg[128]  ( .D(Plaintext[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[128]) );
  DFFSNQ_X1 \reg_in_reg[127]  ( .D(Plaintext[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[127]) );
  DFFSNQ_X1 \reg_in_reg[126]  ( .D(Plaintext[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[126]) );
  DFFSNQ_X1 \reg_in_reg[124]  ( .D(Plaintext[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[124]) );
  DFFSNQ_X1 \reg_in_reg[123]  ( .D(Plaintext[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[123]) );
  DFFSNQ_X1 \reg_in_reg[122]  ( .D(Plaintext[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[122]) );
  DFFSNQ_X1 \reg_in_reg[121]  ( .D(Plaintext[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[121]) );
  DFFSNQ_X1 \reg_in_reg[120]  ( .D(Plaintext[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[120]) );
  DFFSNQ_X1 \reg_in_reg[119]  ( .D(Plaintext[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[119]) );
  DFFSNQ_X1 \reg_in_reg[118]  ( .D(Plaintext[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[118]) );
  DFFSNQ_X1 \reg_in_reg[117]  ( .D(Plaintext[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[117]) );
  DFFSNQ_X1 \reg_in_reg[116]  ( .D(Plaintext[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[116]) );
  DFFSNQ_X1 \reg_in_reg[115]  ( .D(Plaintext[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[115]) );
  DFFSNQ_X1 \reg_in_reg[114]  ( .D(Plaintext[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[114]) );
  DFFSNQ_X1 \reg_in_reg[113]  ( .D(Plaintext[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[113]) );
  DFFSNQ_X1 \reg_in_reg[112]  ( .D(Plaintext[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[112]) );
  DFFSNQ_X1 \reg_in_reg[111]  ( .D(Plaintext[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[111]) );
  DFFSNQ_X1 \reg_in_reg[110]  ( .D(Plaintext[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[110]) );
  DFFSNQ_X1 \reg_in_reg[109]  ( .D(Plaintext[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[109]) );
  DFFSNQ_X1 \reg_in_reg[108]  ( .D(Plaintext[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[108]) );
  DFFSNQ_X1 \reg_in_reg[107]  ( .D(Plaintext[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[107]) );
  DFFSNQ_X1 \reg_in_reg[106]  ( .D(Plaintext[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[106]) );
  DFFSNQ_X1 \reg_in_reg[105]  ( .D(Plaintext[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[105]) );
  DFFSNQ_X1 \reg_in_reg[104]  ( .D(Plaintext[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[104]) );
  DFFSNQ_X1 \reg_in_reg[103]  ( .D(Plaintext[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[103]) );
  DFFSNQ_X1 \reg_in_reg[102]  ( .D(Plaintext[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[102]) );
  DFFSNQ_X1 \reg_in_reg[101]  ( .D(Plaintext[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[101]) );
  DFFSNQ_X1 \reg_in_reg[100]  ( .D(Plaintext[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[100]) );
  DFFSNQ_X1 \reg_in_reg[99]  ( .D(Plaintext[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[99]) );
  DFFSNQ_X1 \reg_in_reg[98]  ( .D(Plaintext[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[98]) );
  DFFSNQ_X1 \reg_in_reg[97]  ( .D(Plaintext[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[97]) );
  DFFSNQ_X1 \reg_in_reg[96]  ( .D(Plaintext[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[96]) );
  DFFSNQ_X1 \reg_in_reg[95]  ( .D(Plaintext[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[95]) );
  DFFSNQ_X1 \reg_in_reg[94]  ( .D(Plaintext[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[94]) );
  DFFSNQ_X1 \reg_in_reg[93]  ( .D(Plaintext[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[93]) );
  DFFSNQ_X1 \reg_in_reg[92]  ( .D(Plaintext[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[92]) );
  DFFSNQ_X1 \reg_in_reg[91]  ( .D(Plaintext[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[91]) );
  DFFSNQ_X1 \reg_in_reg[90]  ( .D(Plaintext[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[90]) );
  DFFSNQ_X1 \reg_in_reg[89]  ( .D(Plaintext[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[89]) );
  DFFSNQ_X1 \reg_in_reg[88]  ( .D(Plaintext[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[88]) );
  DFFSNQ_X1 \reg_in_reg[87]  ( .D(Plaintext[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[87]) );
  DFFSNQ_X1 \reg_in_reg[86]  ( .D(Plaintext[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[86]) );
  DFFSNQ_X1 \reg_in_reg[85]  ( .D(Plaintext[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[85]) );
  DFFSNQ_X1 \reg_in_reg[84]  ( .D(Plaintext[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[84]) );
  DFFSNQ_X1 \reg_in_reg[82]  ( .D(Plaintext[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[82]) );
  DFFSNQ_X1 \reg_in_reg[81]  ( .D(Plaintext[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[81]) );
  DFFSNQ_X1 \reg_in_reg[80]  ( .D(Plaintext[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[80]) );
  DFFSNQ_X1 \reg_in_reg[79]  ( .D(Plaintext[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[79]) );
  DFFSNQ_X1 \reg_in_reg[78]  ( .D(Plaintext[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[78]) );
  DFFSNQ_X1 \reg_in_reg[77]  ( .D(Plaintext[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[77]) );
  DFFSNQ_X1 \reg_in_reg[76]  ( .D(Plaintext[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[76]) );
  DFFSNQ_X1 \reg_in_reg[75]  ( .D(Plaintext[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[75]) );
  DFFSNQ_X1 \reg_in_reg[74]  ( .D(Plaintext[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[74]) );
  DFFSNQ_X1 \reg_in_reg[73]  ( .D(Plaintext[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[73]) );
  DFFSNQ_X1 \reg_in_reg[72]  ( .D(Plaintext[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[72]) );
  DFFSNQ_X1 \reg_in_reg[71]  ( .D(Plaintext[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[71]) );
  DFFSNQ_X1 \reg_in_reg[70]  ( .D(Plaintext[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[70]) );
  DFFSNQ_X1 \reg_in_reg[69]  ( .D(Plaintext[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[69]) );
  DFFSNQ_X1 \reg_in_reg[68]  ( .D(Plaintext[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[68]) );
  DFFSNQ_X1 \reg_in_reg[67]  ( .D(Plaintext[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[67]) );
  DFFSNQ_X1 \reg_in_reg[66]  ( .D(Plaintext[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[66]) );
  DFFSNQ_X1 \reg_in_reg[65]  ( .D(Plaintext[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[65]) );
  DFFSNQ_X1 \reg_in_reg[64]  ( .D(Plaintext[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[64]) );
  DFFSNQ_X1 \reg_in_reg[63]  ( .D(Plaintext[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[63]) );
  DFFSNQ_X1 \reg_in_reg[62]  ( .D(Plaintext[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[62]) );
  DFFSNQ_X1 \reg_in_reg[61]  ( .D(Plaintext[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[61]) );
  DFFSNQ_X1 \reg_in_reg[60]  ( .D(Plaintext[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[60]) );
  DFFSNQ_X1 \reg_in_reg[58]  ( .D(Plaintext[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[58]) );
  DFFSNQ_X1 \reg_in_reg[57]  ( .D(Plaintext[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[57]) );
  DFFSNQ_X1 \reg_in_reg[56]  ( .D(Plaintext[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[56]) );
  DFFSNQ_X1 \reg_in_reg[55]  ( .D(Plaintext[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[55]) );
  DFFSNQ_X1 \reg_in_reg[54]  ( .D(Plaintext[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[54]) );
  DFFSNQ_X1 \reg_in_reg[53]  ( .D(Plaintext[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[53]) );
  DFFSNQ_X1 \reg_in_reg[52]  ( .D(Plaintext[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[52]) );
  DFFSNQ_X1 \reg_in_reg[51]  ( .D(Plaintext[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[51]) );
  DFFSNQ_X1 \reg_in_reg[50]  ( .D(Plaintext[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[50]) );
  DFFSNQ_X1 \reg_in_reg[49]  ( .D(Plaintext[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[49]) );
  DFFSNQ_X1 \reg_in_reg[48]  ( .D(Plaintext[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[48]) );
  DFFSNQ_X1 \reg_in_reg[47]  ( .D(Plaintext[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[47]) );
  DFFSNQ_X1 \reg_in_reg[46]  ( .D(Plaintext[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[46]) );
  DFFSNQ_X1 \reg_in_reg[45]  ( .D(Plaintext[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[45]) );
  DFFSNQ_X1 \reg_in_reg[44]  ( .D(Plaintext[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[44]) );
  DFFSNQ_X1 \reg_in_reg[43]  ( .D(Plaintext[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[43]) );
  DFFSNQ_X1 \reg_in_reg[42]  ( .D(Plaintext[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[42]) );
  DFFSNQ_X1 \reg_in_reg[41]  ( .D(Plaintext[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[41]) );
  DFFSNQ_X1 \reg_in_reg[40]  ( .D(Plaintext[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[40]) );
  DFFSNQ_X1 \reg_in_reg[39]  ( .D(Plaintext[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[39]) );
  DFFSNQ_X1 \reg_in_reg[38]  ( .D(Plaintext[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[38]) );
  DFFSNQ_X1 \reg_in_reg[37]  ( .D(Plaintext[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[37]) );
  DFFSNQ_X1 \reg_in_reg[36]  ( .D(Plaintext[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[36]) );
  DFFSNQ_X1 \reg_in_reg[34]  ( .D(Plaintext[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[34]) );
  DFFSNQ_X1 \reg_in_reg[33]  ( .D(Plaintext[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[33]) );
  DFFSNQ_X1 \reg_in_reg[32]  ( .D(Plaintext[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[32]) );
  DFFSNQ_X1 \reg_in_reg[31]  ( .D(Plaintext[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[31]) );
  DFFSNQ_X1 \reg_in_reg[30]  ( .D(Plaintext[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[30]) );
  DFFSNQ_X1 \reg_in_reg[28]  ( .D(Plaintext[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[28]) );
  DFFSNQ_X1 \reg_in_reg[24]  ( .D(Plaintext[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[24]) );
  DFFSNQ_X1 \reg_in_reg[23]  ( .D(Plaintext[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[23]) );
  DFFSNQ_X1 \reg_in_reg[22]  ( .D(Plaintext[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[22]) );
  DFFSNQ_X1 \reg_in_reg[21]  ( .D(Plaintext[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[21]) );
  DFFSNQ_X1 \reg_in_reg[20]  ( .D(Plaintext[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[20]) );
  DFFSNQ_X1 \reg_in_reg[19]  ( .D(Plaintext[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[19]) );
  DFFSNQ_X1 \reg_in_reg[18]  ( .D(Plaintext[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[18]) );
  DFFSNQ_X1 \reg_in_reg[17]  ( .D(Plaintext[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[17]) );
  DFFSNQ_X1 \reg_in_reg[16]  ( .D(Plaintext[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[16]) );
  DFFSNQ_X1 \reg_in_reg[15]  ( .D(Plaintext[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[15]) );
  DFFSNQ_X1 \reg_in_reg[14]  ( .D(Plaintext[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[14]) );
  DFFSNQ_X1 \reg_in_reg[13]  ( .D(Plaintext[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[13]) );
  DFFSNQ_X1 \reg_in_reg[12]  ( .D(Plaintext[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[12]) );
  DFFSNQ_X1 \reg_in_reg[11]  ( .D(Plaintext[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[11]) );
  DFFSNQ_X1 \reg_in_reg[10]  ( .D(Plaintext[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[10]) );
  DFFSNQ_X1 \reg_in_reg[9]  ( .D(Plaintext[9]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[9]) );
  DFFSNQ_X1 \reg_in_reg[8]  ( .D(Plaintext[8]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[8]) );
  DFFSNQ_X1 \reg_in_reg[7]  ( .D(Plaintext[7]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[7]) );
  DFFSNQ_X1 \reg_in_reg[6]  ( .D(Plaintext[6]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[6]) );
  DFFSNQ_X1 \reg_in_reg[5]  ( .D(Plaintext[5]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[5]) );
  DFFSNQ_X1 \reg_in_reg[4]  ( .D(Plaintext[4]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[4]) );
  DFFSNQ_X1 \reg_in_reg[3]  ( .D(Plaintext[3]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[3]) );
  DFFSNQ_X1 \reg_in_reg[2]  ( .D(Plaintext[2]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[2]) );
  DFFSNQ_X1 \reg_in_reg[1]  ( .D(Plaintext[1]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[1]) );
  DFFSNQ_X1 \reg_in_reg[0]  ( .D(Plaintext[0]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[0]) );
  DFFSNQ_X1 \reg_key_reg[191]  ( .D(Key[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[191]) );
  DFFSNQ_X1 \reg_key_reg[190]  ( .D(Key[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[190]) );
  DFFSNQ_X1 \reg_key_reg[189]  ( .D(Key[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[189]) );
  DFFSNQ_X1 \reg_key_reg[188]  ( .D(Key[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[188]) );
  DFFSNQ_X1 \reg_key_reg[187]  ( .D(Key[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[187]) );
  DFFSNQ_X1 \reg_key_reg[186]  ( .D(Key[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[186]) );
  DFFSNQ_X1 \reg_key_reg[185]  ( .D(Key[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[185]) );
  DFFSNQ_X1 \reg_key_reg[184]  ( .D(Key[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[184]) );
  DFFSNQ_X1 \reg_key_reg[183]  ( .D(Key[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[183]) );
  DFFSNQ_X1 \reg_key_reg[182]  ( .D(Key[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[182]) );
  DFFSNQ_X1 \reg_key_reg[181]  ( .D(Key[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[181]) );
  DFFSNQ_X1 \reg_key_reg[180]  ( .D(Key[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[180]) );
  DFFSNQ_X1 \reg_key_reg[179]  ( .D(Key[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[179]) );
  DFFSNQ_X1 \reg_key_reg[178]  ( .D(Key[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[178]) );
  DFFSNQ_X1 \reg_key_reg[177]  ( .D(Key[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[177]) );
  DFFSNQ_X1 \reg_key_reg[176]  ( .D(Key[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[176]) );
  DFFSNQ_X1 \reg_key_reg[175]  ( .D(Key[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[175]) );
  DFFSNQ_X1 \reg_key_reg[174]  ( .D(Key[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[174]) );
  DFFSNQ_X1 \reg_key_reg[173]  ( .D(Key[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[173]) );
  DFFSNQ_X1 \reg_key_reg[172]  ( .D(Key[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[172]) );
  DFFSNQ_X1 \reg_key_reg[171]  ( .D(Key[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[171]) );
  DFFSNQ_X1 \reg_key_reg[170]  ( .D(Key[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[170]) );
  DFFSNQ_X1 \reg_key_reg[169]  ( .D(Key[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[169]) );
  DFFSNQ_X1 \reg_key_reg[168]  ( .D(Key[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[168]) );
  DFFSNQ_X1 \reg_key_reg[167]  ( .D(Key[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[167]) );
  DFFSNQ_X1 \reg_key_reg[166]  ( .D(Key[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[166]) );
  DFFSNQ_X1 \reg_key_reg[165]  ( .D(Key[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[165]) );
  DFFSNQ_X1 \reg_key_reg[164]  ( .D(Key[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[164]) );
  DFFSNQ_X1 \reg_key_reg[163]  ( .D(Key[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[163]) );
  DFFSNQ_X1 \reg_key_reg[162]  ( .D(Key[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[162]) );
  DFFSNQ_X1 \reg_key_reg[161]  ( .D(Key[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[161]) );
  DFFSNQ_X1 \reg_key_reg[160]  ( .D(Key[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[160]) );
  DFFSNQ_X1 \reg_key_reg[159]  ( .D(Key[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[159]) );
  DFFSNQ_X1 \reg_key_reg[158]  ( .D(Key[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[158]) );
  DFFSNQ_X1 \reg_key_reg[157]  ( .D(Key[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[157]) );
  DFFSNQ_X1 \reg_key_reg[156]  ( .D(Key[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[156]) );
  DFFSNQ_X1 \reg_key_reg[155]  ( .D(Key[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[155]) );
  DFFSNQ_X1 \reg_key_reg[154]  ( .D(Key[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[154]) );
  DFFSNQ_X1 \reg_key_reg[153]  ( .D(Key[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[153]) );
  DFFSNQ_X1 \reg_key_reg[152]  ( .D(Key[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[152]) );
  DFFSNQ_X1 \reg_key_reg[150]  ( .D(Key[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[150]) );
  DFFSNQ_X1 \reg_key_reg[149]  ( .D(Key[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[149]) );
  DFFSNQ_X1 \reg_key_reg[148]  ( .D(Key[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[148]) );
  DFFSNQ_X1 \reg_key_reg[147]  ( .D(Key[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[147]) );
  DFFSNQ_X1 \reg_key_reg[146]  ( .D(Key[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[146]) );
  DFFSNQ_X1 \reg_key_reg[145]  ( .D(Key[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[145]) );
  DFFSNQ_X1 \reg_key_reg[144]  ( .D(Key[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[144]) );
  DFFSNQ_X1 \reg_key_reg[143]  ( .D(Key[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[143]) );
  DFFSNQ_X1 \reg_key_reg[142]  ( .D(Key[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[142]) );
  DFFSNQ_X1 \reg_key_reg[141]  ( .D(Key[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[141]) );
  DFFSNQ_X1 \reg_key_reg[140]  ( .D(Key[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[140]) );
  DFFSNQ_X1 \reg_key_reg[139]  ( .D(Key[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[139]) );
  DFFSNQ_X1 \reg_key_reg[138]  ( .D(Key[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[138]) );
  DFFSNQ_X1 \reg_key_reg[137]  ( .D(Key[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[137]) );
  DFFSNQ_X1 \reg_key_reg[136]  ( .D(Key[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[136]) );
  DFFSNQ_X1 \reg_key_reg[135]  ( .D(Key[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[135]) );
  DFFSNQ_X1 \reg_key_reg[134]  ( .D(Key[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[134]) );
  DFFSNQ_X1 \reg_key_reg[133]  ( .D(Key[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[133]) );
  DFFSNQ_X1 \reg_key_reg[132]  ( .D(Key[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[132]) );
  DFFSNQ_X1 \reg_key_reg[131]  ( .D(Key[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[131]) );
  DFFSNQ_X1 \reg_key_reg[130]  ( .D(Key[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[130]) );
  DFFSNQ_X1 \reg_key_reg[129]  ( .D(Key[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[129]) );
  DFFSNQ_X1 \reg_key_reg[128]  ( .D(Key[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[128]) );
  DFFSNQ_X1 \reg_key_reg[127]  ( .D(Key[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[127]) );
  DFFSNQ_X1 \reg_key_reg[126]  ( .D(Key[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[126]) );
  DFFSNQ_X1 \reg_key_reg[125]  ( .D(Key[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[125]) );
  DFFSNQ_X1 \reg_key_reg[124]  ( .D(Key[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[124]) );
  DFFSNQ_X1 \reg_key_reg[123]  ( .D(Key[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[123]) );
  DFFSNQ_X1 \reg_key_reg[122]  ( .D(Key[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[122]) );
  DFFSNQ_X1 \reg_key_reg[121]  ( .D(Key[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[121]) );
  DFFSNQ_X1 \reg_key_reg[120]  ( .D(Key[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[120]) );
  DFFSNQ_X1 \reg_key_reg[119]  ( .D(Key[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[119]) );
  DFFSNQ_X1 \reg_key_reg[118]  ( .D(Key[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[118]) );
  DFFSNQ_X1 \reg_key_reg[117]  ( .D(Key[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[117]) );
  DFFSNQ_X1 \reg_key_reg[116]  ( .D(Key[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[116]) );
  DFFSNQ_X1 \reg_key_reg[115]  ( .D(Key[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[115]) );
  DFFSNQ_X1 \reg_key_reg[114]  ( .D(Key[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[114]) );
  DFFSNQ_X1 \reg_key_reg[113]  ( .D(Key[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[113]) );
  DFFSNQ_X1 \reg_key_reg[112]  ( .D(Key[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[112]) );
  DFFSNQ_X1 \reg_key_reg[111]  ( .D(Key[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[111]) );
  DFFSNQ_X1 \reg_key_reg[110]  ( .D(Key[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[110]) );
  DFFSNQ_X1 \reg_key_reg[109]  ( .D(Key[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[109]) );
  DFFSNQ_X1 \reg_key_reg[108]  ( .D(Key[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[108]) );
  DFFSNQ_X1 \reg_key_reg[107]  ( .D(Key[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[107]) );
  DFFSNQ_X1 \reg_key_reg[106]  ( .D(Key[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[106]) );
  DFFSNQ_X1 \reg_key_reg[105]  ( .D(Key[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[105]) );
  DFFSNQ_X1 \reg_key_reg[104]  ( .D(Key[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[104]) );
  DFFSNQ_X1 \reg_key_reg[103]  ( .D(Key[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[103]) );
  DFFSNQ_X1 \reg_key_reg[102]  ( .D(Key[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[102]) );
  DFFSNQ_X1 \reg_key_reg[101]  ( .D(Key[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[101]) );
  DFFSNQ_X1 \reg_key_reg[100]  ( .D(Key[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[100]) );
  DFFSNQ_X1 \reg_key_reg[99]  ( .D(Key[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[99]) );
  DFFSNQ_X1 \reg_key_reg[98]  ( .D(Key[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[98]) );
  DFFSNQ_X1 \reg_key_reg[97]  ( .D(Key[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[97]) );
  DFFSNQ_X1 \reg_key_reg[96]  ( .D(Key[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[96]) );
  DFFSNQ_X1 \reg_key_reg[95]  ( .D(Key[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[95]) );
  DFFSNQ_X1 \reg_key_reg[94]  ( .D(Key[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[94]) );
  DFFSNQ_X1 \reg_key_reg[93]  ( .D(Key[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[93]) );
  DFFSNQ_X1 \reg_key_reg[92]  ( .D(Key[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[92]) );
  DFFSNQ_X1 \reg_key_reg[91]  ( .D(Key[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[91]) );
  DFFSNQ_X1 \reg_key_reg[90]  ( .D(Key[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[90]) );
  DFFSNQ_X1 \reg_key_reg[89]  ( .D(Key[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[89]) );
  DFFSNQ_X1 \reg_key_reg[88]  ( .D(Key[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[88]) );
  DFFSNQ_X1 \reg_key_reg[87]  ( .D(Key[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[87]) );
  DFFSNQ_X1 \reg_key_reg[86]  ( .D(Key[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[86]) );
  DFFSNQ_X1 \reg_key_reg[85]  ( .D(Key[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[85]) );
  DFFSNQ_X1 \reg_key_reg[84]  ( .D(Key[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[84]) );
  DFFSNQ_X1 \reg_key_reg[83]  ( .D(Key[83]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[83]) );
  DFFSNQ_X1 \reg_key_reg[82]  ( .D(Key[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[82]) );
  DFFSNQ_X1 \reg_key_reg[81]  ( .D(Key[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[81]) );
  DFFSNQ_X1 \reg_key_reg[80]  ( .D(Key[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[80]) );
  DFFSNQ_X1 \reg_key_reg[79]  ( .D(Key[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[79]) );
  DFFSNQ_X1 \reg_key_reg[78]  ( .D(Key[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[78]) );
  DFFSNQ_X1 \reg_key_reg[77]  ( .D(Key[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[77]) );
  DFFSNQ_X1 \reg_key_reg[76]  ( .D(Key[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[76]) );
  DFFSNQ_X1 \reg_key_reg[75]  ( .D(Key[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[75]) );
  DFFSNQ_X1 \reg_key_reg[74]  ( .D(Key[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[74]) );
  DFFSNQ_X1 \reg_key_reg[73]  ( .D(Key[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[73]) );
  DFFSNQ_X1 \reg_key_reg[72]  ( .D(Key[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[72]) );
  DFFSNQ_X1 \reg_key_reg[71]  ( .D(Key[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[71]) );
  DFFSNQ_X1 \reg_key_reg[70]  ( .D(Key[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[70]) );
  DFFSNQ_X1 \reg_key_reg[69]  ( .D(Key[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[69]) );
  DFFSNQ_X1 \reg_key_reg[68]  ( .D(Key[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[68]) );
  DFFSNQ_X1 \reg_key_reg[67]  ( .D(Key[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[67]) );
  DFFSNQ_X1 \reg_key_reg[66]  ( .D(Key[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[66]) );
  DFFSNQ_X1 \reg_key_reg[65]  ( .D(Key[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[65]) );
  DFFSNQ_X1 \reg_key_reg[64]  ( .D(Key[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[64]) );
  DFFSNQ_X1 \reg_key_reg[63]  ( .D(Key[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[63]) );
  DFFSNQ_X1 \reg_key_reg[62]  ( .D(Key[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[62]) );
  DFFSNQ_X1 \reg_key_reg[61]  ( .D(Key[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[61]) );
  DFFSNQ_X1 \reg_key_reg[60]  ( .D(Key[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[60]) );
  DFFSNQ_X1 \reg_key_reg[59]  ( .D(Key[59]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[59]) );
  DFFSNQ_X1 \reg_key_reg[58]  ( .D(Key[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[58]) );
  DFFSNQ_X1 \reg_key_reg[57]  ( .D(Key[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[57]) );
  DFFSNQ_X1 \reg_key_reg[56]  ( .D(Key[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[56]) );
  DFFSNQ_X1 \reg_key_reg[55]  ( .D(Key[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[55]) );
  DFFSNQ_X1 \reg_key_reg[54]  ( .D(Key[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[54]) );
  DFFSNQ_X1 \reg_key_reg[53]  ( .D(Key[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[53]) );
  DFFSNQ_X1 \reg_key_reg[52]  ( .D(Key[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[52]) );
  DFFSNQ_X1 \reg_key_reg[51]  ( .D(Key[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[51]) );
  DFFSNQ_X1 \reg_key_reg[50]  ( .D(Key[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[50]) );
  DFFSNQ_X1 \reg_key_reg[49]  ( .D(Key[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[49]) );
  DFFSNQ_X1 \reg_key_reg[48]  ( .D(Key[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[48]) );
  DFFSNQ_X1 \reg_key_reg[47]  ( .D(Key[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[47]) );
  DFFSNQ_X1 \reg_key_reg[46]  ( .D(Key[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[46]) );
  DFFSNQ_X1 \reg_key_reg[45]  ( .D(Key[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[45]) );
  DFFSNQ_X1 \reg_key_reg[44]  ( .D(Key[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[44]) );
  DFFSNQ_X1 \reg_key_reg[43]  ( .D(Key[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[43]) );
  DFFSNQ_X1 \reg_key_reg[42]  ( .D(Key[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[42]) );
  DFFSNQ_X1 \reg_key_reg[41]  ( .D(Key[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[41]) );
  DFFSNQ_X1 \reg_key_reg[40]  ( .D(Key[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[40]) );
  DFFSNQ_X1 \reg_key_reg[39]  ( .D(Key[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[39]) );
  DFFSNQ_X1 \reg_key_reg[38]  ( .D(Key[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[38]) );
  DFFSNQ_X1 \reg_key_reg[36]  ( .D(Key[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[36]) );
  DFFSNQ_X1 \reg_key_reg[35]  ( .D(Key[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[35]) );
  DFFSNQ_X1 \reg_key_reg[34]  ( .D(Key[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[34]) );
  DFFSNQ_X1 \reg_key_reg[33]  ( .D(Key[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[33]) );
  DFFSNQ_X1 \reg_key_reg[32]  ( .D(Key[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[32]) );
  DFFSNQ_X1 \reg_key_reg[31]  ( .D(Key[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[31]) );
  DFFSNQ_X1 \reg_key_reg[30]  ( .D(Key[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[30]) );
  DFFSNQ_X1 \reg_key_reg[29]  ( .D(Key[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[29]) );
  DFFSNQ_X1 \reg_key_reg[28]  ( .D(Key[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[28]) );
  DFFSNQ_X1 \reg_key_reg[27]  ( .D(Key[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[27]) );
  DFFSNQ_X1 \reg_key_reg[26]  ( .D(Key[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[26]) );
  DFFSNQ_X1 \reg_key_reg[25]  ( .D(Key[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[25]) );
  DFFSNQ_X1 \reg_key_reg[24]  ( .D(Key[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[24]) );
  DFFSNQ_X1 \reg_key_reg[23]  ( .D(Key[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[23]) );
  DFFSNQ_X1 \reg_key_reg[22]  ( .D(Key[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[22]) );
  DFFSNQ_X1 \reg_key_reg[21]  ( .D(Key[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[21]) );
  DFFSNQ_X1 \reg_key_reg[20]  ( .D(Key[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[20]) );
  DFFSNQ_X1 \reg_key_reg[19]  ( .D(Key[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[19]) );
  DFFSNQ_X1 \reg_key_reg[18]  ( .D(Key[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[18]) );
  DFFSNQ_X1 \reg_key_reg[17]  ( .D(Key[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[17]) );
  DFFSNQ_X1 \reg_key_reg[16]  ( .D(Key[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[16]) );
  DFFSNQ_X1 \reg_key_reg[15]  ( .D(Key[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[15]) );
  DFFSNQ_X1 \reg_key_reg[14]  ( .D(Key[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[14]) );
  DFFSNQ_X1 \reg_key_reg[13]  ( .D(Key[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[13]) );
  DFFSNQ_X1 \reg_key_reg[12]  ( .D(Key[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[12]) );
  DFFSNQ_X1 \reg_key_reg[11]  ( .D(Key[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[11]) );
  DFFSNQ_X1 \reg_key_reg[10]  ( .D(Key[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[10]) );
  DFFSNQ_X1 \reg_key_reg[9]  ( .D(Key[9]), .CLK(clk), .SN(1'b1), .Q(reg_key[9]) );
  DFFSNQ_X1 \reg_key_reg[8]  ( .D(Key[8]), .CLK(clk), .SN(1'b1), .Q(reg_key[8]) );
  DFFSNQ_X1 \reg_key_reg[7]  ( .D(Key[7]), .CLK(clk), .SN(1'b1), .Q(reg_key[7]) );
  DFFSNQ_X1 \reg_key_reg[6]  ( .D(Key[6]), .CLK(clk), .SN(1'b1), .Q(reg_key[6]) );
  DFFSNQ_X1 \reg_key_reg[5]  ( .D(Key[5]), .CLK(clk), .SN(1'b1), .Q(reg_key[5]) );
  DFFSNQ_X1 \reg_key_reg[4]  ( .D(Key[4]), .CLK(clk), .SN(1'b1), .Q(reg_key[4]) );
  DFFSNQ_X1 \reg_key_reg[3]  ( .D(Key[3]), .CLK(clk), .SN(1'b1), .Q(reg_key[3]) );
  DFFSNQ_X1 \reg_key_reg[2]  ( .D(Key[2]), .CLK(clk), .SN(1'b1), .Q(reg_key[2]) );
  DFFSNQ_X1 \reg_key_reg[1]  ( .D(Key[1]), .CLK(clk), .SN(1'b1), .Q(reg_key[1]) );
  DFFSNQ_X1 \reg_key_reg[0]  ( .D(Key[0]), .CLK(clk), .SN(1'b1), .Q(reg_key[0]) );
  DFFSNQ_X1 \Ciphertext_reg[191]  ( .D(reg_out[191]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[191]) );
  DFFSNQ_X1 \Ciphertext_reg[188]  ( .D(reg_out[188]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[188]) );
  DFFSNQ_X1 \Ciphertext_reg[187]  ( .D(reg_out[187]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[187]) );
  DFFSNQ_X1 \Ciphertext_reg[184]  ( .D(reg_out[184]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[184]) );
  DFFSNQ_X1 \Ciphertext_reg[183]  ( .D(reg_out[183]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[183]) );
  DFFSNQ_X1 \Ciphertext_reg[181]  ( .D(reg_out[181]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[181]) );
  DFFSNQ_X1 \Ciphertext_reg[179]  ( .D(reg_out[179]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[179]) );
  DFFSNQ_X1 \Ciphertext_reg[178]  ( .D(reg_out[178]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[178]) );
  DFFSNQ_X1 \Ciphertext_reg[177]  ( .D(reg_out[177]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[177]) );
  DFFSNQ_X1 \Ciphertext_reg[176]  ( .D(reg_out[176]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[176]) );
  DFFSNQ_X1 \Ciphertext_reg[175]  ( .D(reg_out[175]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[175]) );
  DFFSNQ_X1 \Ciphertext_reg[173]  ( .D(reg_out[173]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[173]) );
  DFFSNQ_X1 \Ciphertext_reg[172]  ( .D(reg_out[172]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[172]) );
  DFFSNQ_X1 \Ciphertext_reg[170]  ( .D(reg_out[170]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[170]) );
  DFFSNQ_X1 \Ciphertext_reg[168]  ( .D(reg_out[168]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[168]) );
  DFFSNQ_X1 \Ciphertext_reg[167]  ( .D(reg_out[167]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[167]) );
  DFFSNQ_X1 \Ciphertext_reg[166]  ( .D(reg_out[166]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[166]) );
  DFFSNQ_X1 \Ciphertext_reg[163]  ( .D(reg_out[163]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[163]) );
  DFFSNQ_X1 \Ciphertext_reg[161]  ( .D(reg_out[161]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[161]) );
  DFFSNQ_X1 \Ciphertext_reg[158]  ( .D(reg_out[158]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[158]) );
  DFFSNQ_X1 \Ciphertext_reg[157]  ( .D(reg_out[157]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[157]) );
  DFFSNQ_X1 \Ciphertext_reg[156]  ( .D(reg_out[156]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[156]) );
  DFFSNQ_X1 \Ciphertext_reg[155]  ( .D(reg_out[155]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[155]) );
  DFFSNQ_X1 \Ciphertext_reg[151]  ( .D(reg_out[151]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[151]) );
  DFFSNQ_X1 \Ciphertext_reg[150]  ( .D(reg_out[150]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[150]) );
  DFFSNQ_X1 \Ciphertext_reg[149]  ( .D(reg_out[149]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[149]) );
  DFFSNQ_X1 \Ciphertext_reg[148]  ( .D(reg_out[148]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[148]) );
  DFFSNQ_X1 \Ciphertext_reg[147]  ( .D(reg_out[147]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[147]) );
  DFFSNQ_X1 \Ciphertext_reg[145]  ( .D(reg_out[145]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[145]) );
  DFFSNQ_X1 \Ciphertext_reg[144]  ( .D(reg_out[144]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[144]) );
  DFFSNQ_X1 \Ciphertext_reg[142]  ( .D(reg_out[142]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[142]) );
  DFFSNQ_X1 \Ciphertext_reg[141]  ( .D(reg_out[141]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[141]) );
  DFFSNQ_X1 \Ciphertext_reg[140]  ( .D(reg_out[140]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[140]) );
  DFFSNQ_X1 \Ciphertext_reg[139]  ( .D(reg_out[139]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[139]) );
  DFFSNQ_X1 \Ciphertext_reg[138]  ( .D(reg_out[138]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[138]) );
  DFFSNQ_X1 \Ciphertext_reg[135]  ( .D(reg_out[135]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[135]) );
  DFFSNQ_X1 \Ciphertext_reg[134]  ( .D(reg_out[134]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[134]) );
  DFFSNQ_X1 \Ciphertext_reg[129]  ( .D(reg_out[129]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[129]) );
  DFFSNQ_X1 \Ciphertext_reg[128]  ( .D(reg_out[128]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[128]) );
  DFFSNQ_X1 \Ciphertext_reg[127]  ( .D(reg_out[127]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[127]) );
  DFFSNQ_X1 \Ciphertext_reg[126]  ( .D(reg_out[126]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[126]) );
  DFFSNQ_X1 \Ciphertext_reg[123]  ( .D(reg_out[123]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[123]) );
  DFFSNQ_X1 \Ciphertext_reg[122]  ( .D(reg_out[122]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[122]) );
  DFFSNQ_X1 \Ciphertext_reg[121]  ( .D(reg_out[121]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[121]) );
  DFFSNQ_X1 \Ciphertext_reg[119]  ( .D(reg_out[119]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[119]) );
  DFFSNQ_X1 \Ciphertext_reg[118]  ( .D(reg_out[118]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[118]) );
  DFFSNQ_X1 \Ciphertext_reg[115]  ( .D(reg_out[115]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[115]) );
  DFFSNQ_X1 \Ciphertext_reg[113]  ( .D(reg_out[113]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[113]) );
  DFFSNQ_X1 \Ciphertext_reg[112]  ( .D(reg_out[112]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[112]) );
  DFFSNQ_X1 \Ciphertext_reg[110]  ( .D(reg_out[110]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[110]) );
  DFFSNQ_X1 \Ciphertext_reg[109]  ( .D(reg_out[109]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[109]) );
  DFFSNQ_X1 \Ciphertext_reg[108]  ( .D(reg_out[108]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[108]) );
  DFFSNQ_X1 \Ciphertext_reg[107]  ( .D(reg_out[107]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[107]) );
  DFFSNQ_X1 \Ciphertext_reg[106]  ( .D(reg_out[106]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[106]) );
  DFFSNQ_X1 \Ciphertext_reg[105]  ( .D(reg_out[105]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[105]) );
  DFFSNQ_X1 \Ciphertext_reg[104]  ( .D(reg_out[104]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[104]) );
  DFFSNQ_X1 \Ciphertext_reg[103]  ( .D(reg_out[103]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[103]) );
  DFFSNQ_X1 \Ciphertext_reg[102]  ( .D(reg_out[102]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[102]) );
  DFFSNQ_X1 \Ciphertext_reg[98]  ( .D(reg_out[98]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[98]) );
  DFFSNQ_X1 \Ciphertext_reg[96]  ( .D(reg_out[96]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[96]) );
  DFFSNQ_X1 \Ciphertext_reg[93]  ( .D(reg_out[93]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[93]) );
  DFFSNQ_X1 \Ciphertext_reg[92]  ( .D(reg_out[92]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[92]) );
  DFFSNQ_X1 \Ciphertext_reg[91]  ( .D(reg_out[91]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[91]) );
  DFFSNQ_X1 \Ciphertext_reg[90]  ( .D(reg_out[90]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[90]) );
  DFFSNQ_X1 \Ciphertext_reg[89]  ( .D(reg_out[89]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[89]) );
  DFFSNQ_X1 \Ciphertext_reg[86]  ( .D(reg_out[86]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[86]) );
  DFFSNQ_X1 \Ciphertext_reg[85]  ( .D(reg_out[85]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[85]) );
  DFFSNQ_X1 \Ciphertext_reg[84]  ( .D(reg_out[84]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[84]) );
  DFFSNQ_X1 \Ciphertext_reg[83]  ( .D(reg_out[83]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[83]) );
  DFFSNQ_X1 \Ciphertext_reg[82]  ( .D(reg_out[82]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[82]) );
  DFFSNQ_X1 \Ciphertext_reg[81]  ( .D(reg_out[81]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[81]) );
  DFFSNQ_X1 \Ciphertext_reg[80]  ( .D(reg_out[80]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[80]) );
  DFFSNQ_X1 \Ciphertext_reg[79]  ( .D(reg_out[79]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[79]) );
  DFFSNQ_X1 \Ciphertext_reg[78]  ( .D(reg_out[78]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[78]) );
  DFFSNQ_X1 \Ciphertext_reg[77]  ( .D(reg_out[77]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[77]) );
  DFFSNQ_X1 \Ciphertext_reg[76]  ( .D(reg_out[76]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[76]) );
  DFFSNQ_X1 \Ciphertext_reg[74]  ( .D(reg_out[74]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[74]) );
  DFFSNQ_X1 \Ciphertext_reg[73]  ( .D(reg_out[73]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[73]) );
  DFFSNQ_X1 \Ciphertext_reg[71]  ( .D(reg_out[71]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[71]) );
  DFFSNQ_X1 \Ciphertext_reg[70]  ( .D(reg_out[70]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[70]) );
  DFFSNQ_X1 \Ciphertext_reg[69]  ( .D(reg_out[69]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[69]) );
  DFFSNQ_X1 \Ciphertext_reg[68]  ( .D(reg_out[68]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[68]) );
  DFFSNQ_X1 \Ciphertext_reg[67]  ( .D(reg_out[67]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[67]) );
  DFFSNQ_X1 \Ciphertext_reg[66]  ( .D(reg_out[66]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[66]) );
  DFFSNQ_X1 \Ciphertext_reg[65]  ( .D(reg_out[65]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[65]) );
  DFFSNQ_X1 \Ciphertext_reg[64]  ( .D(reg_out[64]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[64]) );
  DFFSNQ_X1 \Ciphertext_reg[63]  ( .D(reg_out[63]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[63]) );
  DFFSNQ_X1 \Ciphertext_reg[62]  ( .D(reg_out[62]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[62]) );
  DFFSNQ_X1 \Ciphertext_reg[61]  ( .D(reg_out[61]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[61]) );
  DFFSNQ_X1 \Ciphertext_reg[60]  ( .D(reg_out[60]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[60]) );
  DFFSNQ_X1 \Ciphertext_reg[55]  ( .D(reg_out[55]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[55]) );
  DFFSNQ_X1 \Ciphertext_reg[53]  ( .D(reg_out[53]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[53]) );
  DFFSNQ_X1 \Ciphertext_reg[52]  ( .D(reg_out[52]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[52]) );
  DFFSNQ_X1 \Ciphertext_reg[51]  ( .D(reg_out[51]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[51]) );
  DFFSNQ_X1 \Ciphertext_reg[50]  ( .D(reg_out[50]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[50]) );
  DFFSNQ_X1 \Ciphertext_reg[48]  ( .D(reg_out[48]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[48]) );
  DFFSNQ_X1 \Ciphertext_reg[47]  ( .D(reg_out[47]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[47]) );
  DFFSNQ_X1 \Ciphertext_reg[46]  ( .D(reg_out[46]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[46]) );
  DFFSNQ_X1 \Ciphertext_reg[45]  ( .D(reg_out[45]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[45]) );
  DFFSNQ_X1 \Ciphertext_reg[44]  ( .D(reg_out[44]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[44]) );
  DFFSNQ_X1 \Ciphertext_reg[43]  ( .D(reg_out[43]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[43]) );
  DFFSNQ_X1 \Ciphertext_reg[42]  ( .D(reg_out[42]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[42]) );
  DFFSNQ_X1 \Ciphertext_reg[41]  ( .D(reg_out[41]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[41]) );
  DFFSNQ_X1 \Ciphertext_reg[40]  ( .D(reg_out[40]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[40]) );
  DFFSNQ_X1 \Ciphertext_reg[38]  ( .D(reg_out[38]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[38]) );
  DFFSNQ_X1 \Ciphertext_reg[37]  ( .D(reg_out[37]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[37]) );
  DFFSNQ_X1 \Ciphertext_reg[36]  ( .D(reg_out[36]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[36]) );
  DFFSNQ_X1 \Ciphertext_reg[35]  ( .D(reg_out[35]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[35]) );
  DFFSNQ_X1 \Ciphertext_reg[34]  ( .D(reg_out[34]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[34]) );
  DFFSNQ_X1 \Ciphertext_reg[31]  ( .D(reg_out[31]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[31]) );
  DFFSNQ_X1 \Ciphertext_reg[29]  ( .D(reg_out[29]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[29]) );
  DFFSNQ_X1 \Ciphertext_reg[27]  ( .D(reg_out[27]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[27]) );
  DFFSNQ_X1 \Ciphertext_reg[25]  ( .D(reg_out[25]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[25]) );
  DFFSNQ_X1 \Ciphertext_reg[24]  ( .D(reg_out[24]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[24]) );
  DFFSNQ_X1 \Ciphertext_reg[22]  ( .D(reg_out[22]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[22]) );
  DFFSNQ_X1 \Ciphertext_reg[19]  ( .D(reg_out[19]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[19]) );
  DFFSNQ_X1 \Ciphertext_reg[18]  ( .D(reg_out[18]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[18]) );
  DFFSNQ_X1 \Ciphertext_reg[17]  ( .D(reg_out[17]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[17]) );
  DFFSNQ_X1 \Ciphertext_reg[16]  ( .D(reg_out[16]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[16]) );
  DFFSNQ_X1 \Ciphertext_reg[15]  ( .D(reg_out[15]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[15]) );
  DFFSNQ_X1 \Ciphertext_reg[13]  ( .D(reg_out[13]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[13]) );
  DFFSNQ_X1 \Ciphertext_reg[12]  ( .D(reg_out[12]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[12]) );
  DFFSNQ_X1 \Ciphertext_reg[11]  ( .D(reg_out[11]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[11]) );
  DFFSNQ_X1 \Ciphertext_reg[7]  ( .D(reg_out[7]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[7]) );
  DFFSNQ_X1 \Ciphertext_reg[6]  ( .D(reg_out[6]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[6]) );
  DFFSNQ_X1 \Ciphertext_reg[5]  ( .D(reg_out[5]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[5]) );
  DFFSNQ_X1 \Ciphertext_reg[4]  ( .D(reg_out[4]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[4]) );
  DFFSNQ_X1 \Ciphertext_reg[2]  ( .D(reg_out[2]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[2]) );
  DFFSNQ_X1 \Ciphertext_reg[1]  ( .D(reg_out[1]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[1]) );
  DFFRNQ_X1 \Ciphertext_reg[160]  ( .D(reg_out[160]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[160]) );
  DFFRNQ_X1 \Ciphertext_reg[159]  ( .D(reg_out[159]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[159]) );
  DFFRNQ_X1 \Ciphertext_reg[10]  ( .D(reg_out[10]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[10]) );
  DFFRNQ_X1 \reg_in_reg[125]  ( .D(Plaintext[125]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[125]) );
  DFFRNQ_X1 \Ciphertext_reg[132]  ( .D(reg_out[132]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[132]) );
  DFFRNQ_X1 \Ciphertext_reg[49]  ( .D(reg_out[49]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[49]) );
  DFFRNQ_X1 \Ciphertext_reg[33]  ( .D(reg_out[33]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[33]) );
  DFFRNQ_X1 \Ciphertext_reg[3]  ( .D(reg_out[3]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[3]) );
  DFFRNQ_X1 \Ciphertext_reg[185]  ( .D(reg_out[185]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[185]) );
  DFFRNQ_X1 \reg_in_reg[25]  ( .D(Plaintext[25]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[25]) );
  DFFRNQ_X1 \Ciphertext_reg[99]  ( .D(reg_out[99]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[99]) );
  DFFRNQ_X1 \Ciphertext_reg[116]  ( .D(reg_out[116]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[116]) );
  DFFRNQ_X1 \Ciphertext_reg[32]  ( .D(reg_out[32]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[32]) );
  DFFRNQ_X1 \Ciphertext_reg[125]  ( .D(reg_out[125]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[125]) );
  DFFRNQ_X1 \Ciphertext_reg[94]  ( .D(reg_out[94]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[94]) );
  DFFRNQ_X1 \Ciphertext_reg[143]  ( .D(reg_out[143]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[143]) );
  DFFRNQ_X1 \Ciphertext_reg[75]  ( .D(reg_out[75]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[75]) );
  DFFRNQ_X1 \Ciphertext_reg[114]  ( .D(reg_out[114]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[114]) );
  DFFRNQ_X1 \Ciphertext_reg[186]  ( .D(reg_out[186]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[186]) );
  DFFRNQ_X1 \Ciphertext_reg[21]  ( .D(reg_out[21]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[21]) );
  DFFRNQ_X1 \Ciphertext_reg[154]  ( .D(reg_out[154]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[154]) );
  DFFRNQ_X1 \Ciphertext_reg[14]  ( .D(reg_out[14]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[14]) );
  DFFRNQ_X1 \reg_in_reg[140]  ( .D(Plaintext[140]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[140]) );
  DFFRNQ_X1 \Ciphertext_reg[20]  ( .D(reg_out[20]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[20]) );
  DFFRNQ_X1 \reg_in_reg[35]  ( .D(Plaintext[35]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[35]) );
  DFFRNQ_X1 \Ciphertext_reg[124]  ( .D(reg_out[124]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[124]) );
  DFFRNQ_X1 \Ciphertext_reg[136]  ( .D(reg_out[136]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[136]) );
  DFFRNQ_X1 \Ciphertext_reg[9]  ( .D(reg_out[9]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[9]) );
  DFFRNQ_X1 \Ciphertext_reg[28]  ( .D(reg_out[28]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[28]) );
  DFFRNQ_X1 \Ciphertext_reg[23]  ( .D(reg_out[23]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[23]) );
  DFFRNQ_X1 \Ciphertext_reg[111]  ( .D(reg_out[111]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[111]) );
  DFFRNQ_X1 \Ciphertext_reg[30]  ( .D(reg_out[30]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[30]) );
  DFFRNQ_X1 \Ciphertext_reg[101]  ( .D(reg_out[101]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[101]) );
  DFFRNQ_X1 \Ciphertext_reg[87]  ( .D(reg_out[87]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[87]) );
  DFFRNQ_X1 \reg_in_reg[169]  ( .D(Plaintext[169]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[169]) );
  DFFRNQ_X1 \Ciphertext_reg[117]  ( .D(reg_out[117]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[117]) );
  DFFRNQ_X1 \Ciphertext_reg[133]  ( .D(reg_out[133]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[133]) );
  DFFRNQ_X1 \Ciphertext_reg[146]  ( .D(reg_out[146]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[146]) );
  DFFSNQ_X1 \Ciphertext_reg[88]  ( .D(reg_out[88]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[88]) );
  DFFRNQ_X1 \Ciphertext_reg[72]  ( .D(reg_out[72]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[72]) );
  DFFRNQ_X1 \Ciphertext_reg[100]  ( .D(reg_out[100]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[100]) );
  DFFRNQ_X1 \Ciphertext_reg[130]  ( .D(reg_out[130]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[130]) );
  DFFRNQ_X1 \Ciphertext_reg[59]  ( .D(reg_out[59]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[59]) );
  DFFRNQ_X1 \Ciphertext_reg[0]  ( .D(reg_out[0]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[0]) );
  DFFRNQ_X1 \Ciphertext_reg[58]  ( .D(reg_out[58]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[58]) );
  DFFRNQ_X1 \Ciphertext_reg[26]  ( .D(reg_out[26]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[26]) );
  DFFRNQ_X1 \Ciphertext_reg[131]  ( .D(reg_out[131]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[131]) );
  DFFRNQ_X1 \Ciphertext_reg[189]  ( .D(reg_out[189]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[189]) );
  DFFRNQ_X1 \Ciphertext_reg[56]  ( .D(reg_out[56]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[56]) );
  DFFRNQ_X1 \Ciphertext_reg[54]  ( .D(reg_out[54]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[54]) );
  DFFRNQ_X1 \Ciphertext_reg[153]  ( .D(reg_out[153]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[153]) );
  DFFRNQ_X1 \Ciphertext_reg[174]  ( .D(reg_out[174]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[174]) );
  DFFRNQ_X1 \reg_in_reg[146]  ( .D(Plaintext[146]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[146]) );
  DFFRNQ_X1 \Ciphertext_reg[171]  ( .D(reg_out[171]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[171]) );
  DFFRNQ_X1 \Ciphertext_reg[180]  ( .D(reg_out[180]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[180]) );
  DFFRNQ_X1 \reg_key_reg[37]  ( .D(Key[37]), .CLK(clk), .RN(1'b1), .Q(
        reg_key[37]) );
  DFFRNQ_X1 \Ciphertext_reg[182]  ( .D(reg_out[182]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[182]) );
  DFFRNQ_X1 \reg_in_reg[83]  ( .D(Plaintext[83]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[83]) );
  DFFRNQ_X1 \Ciphertext_reg[152]  ( .D(reg_out[152]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[152]) );
  DFFRNQ_X1 \Ciphertext_reg[120]  ( .D(reg_out[120]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[120]) );
  DFFRNQ_X1 \Ciphertext_reg[137]  ( .D(reg_out[137]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[137]) );
  DFFSNQ_X1 \reg_in_reg[191]  ( .D(Plaintext[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[191]) );
  DFFRNQ_X1 \Ciphertext_reg[190]  ( .D(reg_out[190]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[190]) );
  DFFRNQ_X1 \Ciphertext_reg[97]  ( .D(reg_out[97]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[97]) );
  DFFRNQ_X1 \reg_in_reg[59]  ( .D(Plaintext[59]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[59]) );
  SPEEDY_Rounds7_0 SPEEDY_instance ( .Plaintext(reg_in), .Key(reg_key), 
        .Ciphertext(reg_out) );
  DFFRNQ_X1 \Ciphertext_reg[164]  ( .D(reg_out[164]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[164]) );
  DFFRNQ_X1 \Ciphertext_reg[162]  ( .D(reg_out[162]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[162]) );
  DFFSNQ_X1 \reg_in_reg[29]  ( .D(Plaintext[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[29]) );
  DFFRNQ_X1 \reg_in_reg[26]  ( .D(Plaintext[26]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[26]) );
  DFFRNQ_X1 \reg_key_reg[151]  ( .D(Key[151]), .CLK(clk), .RN(1'b1), .Q(
        reg_key[151]) );
  DFFRNQ_X1 \Ciphertext_reg[8]  ( .D(reg_out[8]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[8]) );
  DFFRNQ_X1 \Ciphertext_reg[95]  ( .D(reg_out[95]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[95]) );
  DFFSNQ_X1 \Ciphertext_reg[165]  ( .D(reg_out[165]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[165]) );
  DFFRNQ_X1 \Ciphertext_reg[169]  ( .D(reg_out[169]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[169]) );
  DFFSNQ_X1 \Ciphertext_reg[39]  ( .D(reg_out[39]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[39]) );
  DFFRNQ_X1 \reg_in_reg[27]  ( .D(Plaintext[27]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[27]) );
  DFFRNQ_X1 \Ciphertext_reg[57]  ( .D(reg_out[57]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[57]) );
endmodule

