module SPEEDY_Rounds6_0 ( Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31,
         n32, n34, n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n51, n52,
         n55, n58, n59, n60, n61, n62, n66, n68, n69, n70, n71, n72, n73, n75,
         n76, n77, n78, n79, n81, n82, n85, n87, n88, n89, n92, n95, n96, n97,
         n98, n100, n101, n102, n103, n104, n107, n108, n109, n111, n112, n113,
         n114, n115, n118, n119, n120, n121, n122, n123, n125, n126, n127,
         n128, n129, n131, n133, n135, n136, n137, n138, n139, n140, n141,
         n142, n144, n145, n146, n147, n148, n149, n151, n152, n153, n155,
         n156, n158, n159, n160, n161, n162, n164, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n185,
         n187, n188, n189, n190, n191, n194, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n223, n227, n231, n232, n233, n238, n239, n240, n244,
         n245, n246, n248, n249, n250, n257, n260, n261, n262, n263, n264,
         n266, n267, n268, n269, n270, n271, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n287, n288, n290, n291,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n307, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n343, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n376, n377, n379,
         n380, n381, n382, n383, n385, n386, n387, n388, n389, n391, n392,
         n394, n395, n396, n397, n398, n399, n400, n401, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n462, n463, n464,
         n465, n467, n468, n469, n470, n471, n472, n473, n474, n475, n477,
         n478, n479, n480, n481, n483, n484, n486, n488, n491, n492, n493,
         n494, n495, n496, n498, n499, n500, n501, n502, n504, n505, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n545, n546, n547, n548, n549, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n578, n579, n580, n581, n584, n585, n586, n587, n588, n589, n590,
         n593, n594, n595, n596, n597, n598, n599, n600, n602, n603, n605,
         n606, n607, n608, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n640, n641,
         n642, n644, n645, n646, n647, n648, n649, n650, n651, n652, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n692, n693, n695, n696, n697, n698, n699, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n718, n719, n720, n721, n722, n723, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n740, n741,
         n742, n743, n744, n746, n747, n749, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n775, n776, n777, n778, n779,
         n780, n781, n782, n784, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n804,
         n806, n807, n808, n809, n810, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n845, n847, n848, n849, n852, n853, n854,
         n855, n856, n857, n859, n860, n861, n862, n863, n864, n867, n868,
         n869, n870, n871, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n905, n906, n907, n908, n909, n910, n911, n912, n914, n915,
         n916, n918, n919, n920, n921, n923, n924, n925, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n965, n966, n967, n968, n969, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1032, n1033,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1065,
         n1066, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1095, n1096, n1097,
         n1098, n1099, n1100, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1152, n1153, n1154, n1155, n1156, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1208, n1210, n1211, n1212, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1235, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1272, n1273,
         n1275, n1276, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1299, n1300, n1301, n1302, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1351, n1352,
         n1353, n1355, n1357, n1358, n1359, n1361, n1362, n1363, n1364, n1365,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1526, n1527, n1528, n1530, n1531,
         n1532, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1556, n1557, n1558, n1559, n1561, n1562, n1563, n1564,
         n1566, n1568, n1569, n1570, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1604, n1605, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1653,
         n1654, n1655, n1656, n1658, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1718, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1852, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1938, n1939, n1940, n1941, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1987,
         n1988, n1990, n1991, n1992, n1993, n1995, n1996, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2015, n2016, n2017, n2018, n2020, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2064, n2066, n2067,
         n2068, n2069, n2070, n2071, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2124, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2183, n2184, n2185,
         n2186, n2187, n2188, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2198, n2199, n2202, n2203, n2204, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2238, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2338, n2339, n2341, n2342, n2344, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2435, n2436, n2437, n2438, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2520, n2521, n2522, n2523, n2524, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2580,
         n2581, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2648, n2649, n2650, n2651, n2652, n2653, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2673, n2674, n2675, n2677, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2701, n2702, n2703, n2704,
         n2706, n2708, n2709, n2710, n2711, n2713, n2714, n2715, n2717, n2718,
         n2720, n2721, n2722, n2724, n2725, n2726, n2727, n2728, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2821, n2823, n2824, n2826, n2827, n2828, n2829, n2830,
         n2831, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2857, n2858, n2859, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2951, n2952, n2953, n2955, n2956, n2957,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3016, n3018, n3022, n3024, n3025, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3093, n3094, n3095, n3096, n3097, n3098, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3109, n3110, n3111, n3112, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3152, n3153, n3155, n3156, n3157, n3158,
         n3159, n3160, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3280, n3281, n3282, n3283, n3284,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3365, n3366, n3367, n3368, n3369, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3469, n3470, n3471, n3472, n3473, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3532, n3533, n3534, n3535, n3536, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3561, n3562,
         n3563, n3564, n3565, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3578, n3579, n3580, n3581, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3620, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3645, n3646, n3647, n3648, n3650, n3651, n3652,
         n3653, n3655, n3656, n3657, n3658, n3660, n3661, n3662, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3688, n3689, n3690, n3691, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3791, n3792,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3804,
         n3805, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3826, n3827,
         n3828, n3829, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3898, n3899, n3900, n3901, n3903,
         n3904, n3906, n3907, n3908, n3909, n3910, n3912, n3913, n3914, n3916,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4120, n4121, n4122, n4123, n4124, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4221, n4222, n4224, n4225, n4226, n4227, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4272, n4273, n4274,
         n4276, n4277, n4278, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4311, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4326, n4327, n4328, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4495, n4496, n4497, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4520, n4521, n4522, n4523, n4524, n4525, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4536, n4537, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4556, n4557, n4558, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4600, n4601, n4602, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4624, n4625, n4626, n4627,
         n4628, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4686, n4687, n4688, n4689, n4691, n4692,
         n4694, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4777, n4778, n4779, n4780, n4781, n4782, n4784, n4785, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4832, n4833, n4834, n4835, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4848, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4906,
         n4907, n4908, n4909, n4910, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4936, n4937, n4938, n4939,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4953, n4954, n4956, n4957, n4958, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5006,
         n5007, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5017, n5018,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5068, n5070, n5071, n5072, n5073,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5119, n5120, n5121, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5427, n5428, n5429,
         n5432, n5433, n5434, n5436, n5437, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5563, n5564, n5565, n5566, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5581, n5582,
         n5583, n5584, n5585, n5586, n5588, n5589, n5590, n5591, n5593, n5594,
         n5595, n5596, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5658, n5659, n5660, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5719, n5720, n5722,
         n5723, n5724, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6319, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6742, n6743, n6744, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7018, n7019, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7097,
         n7098, n7099, n7100, n7101, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7132, n7133, n7135, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7310, n7311, n7312, n7313, n7314, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7524, n7525, n7526, n7527, n7528, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7556, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7881, n7882, n7883,
         n7884, n7885, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9143, n9144, n9145, n9146, n9147, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9208, n9209, n9210, n9211,
         n9212, n9213, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9293,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9325, n9326,
         n9327, n9328, n9329, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9342, n9343, n9345, n9346, n9348, n9349, n9350, n9351,
         n9354, n9355, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9490, n9491, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9512, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9984,
         n9985, n9986, n9989, n9990, n9991, n9992, n9993, n9994, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10031, n10032,
         n10033, n10034, n10035, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10103, n10104, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10122, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10151, n10152,
         n10154, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10538, n10539, n10540,
         n10541, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10627, n10628, n10629, n10630, n10632, n10633,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11103, n11104, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11199, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11324, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12526,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12546, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12592, n12593, n12594, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12619, n12620, n12621, n12622,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12852, n12853, n12854, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12887, n12888, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12973, n12974, n12975, n12976, n12977, n12979, n12980, n12981,
         n12982, n12983, n12984, n12986, n12987, n12988, n12991, n12993,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13202, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13254, n13255, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13286, n13287, n13288, n13289, n13291, n13292,
         n13294, n13295, n13296, n13297, n13298, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13341, n13342, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13436, n13437, n13438,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13449,
         n13450, n13453, n13454, n13457, n13458, n13459, n13460, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13633, n13634,
         n13635, n13636, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13646, n13647, n13648, n13649, n13650, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13690, n13691, n13692, n13693, n13695,
         n13696, n13697, n13698, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13977, n13978, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14097, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14188, n14189, n14190,
         n14191, n14192, n14194, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14273, n14274, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14744, n14745,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15316, n15317, n15318,
         n15319, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15559, n15560, n15562, n15563, n15564, n15565, n15566,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15604, n15605, n15606, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15625, n15626, n15627,
         n15628, n15629, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15739, n15740, n15741, n15742, n15744, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15757, n15758, n15759, n15760, n15761, n15762, n15764,
         n15765, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15890, n15891, n15892,
         n15893, n15894, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16041, n16042, n16043, n16045, n16046, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16080, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16154, n16155, n16156, n16157, n16158, n16159, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16276, n16277, n16278,
         n16280, n16281, n16283, n16284, n16285, n16286, n16287, n16288,
         n16290, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16339, n16340, n16341,
         n16342, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16593, n16595, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16712, n16713, n16714, n16715, n16716,
         n16717, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16789, n16790, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16806, n16807, n16808, n16809, n16810, n16811, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17148, n17150, n17151,
         n17152, n17153, n17154, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17291, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17463, n17464, n17465,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17551, n17552, n17553, n17554, n17555,
         n17556, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17705, n17706, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18116, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18714,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18869, n18870, n18871,
         n18872, n18873, n18874, n18876, n18877, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18907,
         n18908, n18909, n18911, n18912, n18913, n18914, n18916, n18917,
         n18918, n18919, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19035,
         n19036, n19037, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19056, n19057, n19059, n19060, n19061, n19062,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19213, n19214,
         n19215, n19217, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19359, n19360, n19361, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19395, n19396, n19397, n19398, n19399, n19400, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19451, n19452, n19456, n19457, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19490, n19491, n19492, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19518, n19519,
         n19520, n19521, n19522, n19523, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19645,
         n19646, n19647, n19648, n19649, n19650, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19758, n19759, n19760, n19761,
         n19762, n19764, n19765, n19766, n19767, n19768, n19769, n19772,
         n19773, n19774, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19920,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19941, n19942, n19943, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20013, n20014,
         n20015, n20016, n20017, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20058, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20109, n20111, n20112,
         n20113, n20114, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20199, n20200, n20201, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20319, n20320, n20321, n20322, n20323,
         n20324, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20501, n20502, n20503, n20504, n20505, n20507, n20508,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20525, n20526,
         n20527, n20528, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21023, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21070, n21071,
         n21072, n21073, n21074, n21075, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21389, n21390,
         n21391, n21392, n21393, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21781, n21782, n21783, n21784, n21785, n21786, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21844, n21845,
         n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853,
         n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861,
         n21862, n21863, n21864, n21865, n21866, n21868, n21869, n21870,
         n21871, n21872, n21873, n21874, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22052, n22053, n22054, n22055, n22056, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22070, n22071, n22072, n22074, n22075, n22076, n22077, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22095, n22096,
         n22097, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22155, n22156, n22157, n22158, n22159, n22161, n22162, n22163,
         n22164, n22165, n22166, n22168, n22169, n22170, n22172, n22173,
         n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181,
         n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22190,
         n22191, n22192, n22193, n22194, n22195, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22252, n22253, n22254, n22255, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22284, n22285,
         n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293,
         n22294, n22295, n22296, n22297, n22298, n22299, n22301, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22424, n22426, n22427, n22428, n22429,
         n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437,
         n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22446,
         n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454,
         n22455, n22456, n22458, n22459, n22461, n22462, n22463, n22464,
         n22465, n22466, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22482,
         n22483, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22521, n22522, n22523, n22524,
         n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
         n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
         n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
         n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
         n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
         n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572,
         n22573, n22574, n22575, n22576, n22578, n22579, n22580, n22581,
         n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589,
         n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597,
         n22598, n22600, n22601, n22602, n22603, n22604, n22605, n22606,
         n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614,
         n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622,
         n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630,
         n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638,
         n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646,
         n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654,
         n22655, n22656, n22657, n22658, n22659, n22661, n22663, n22664,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
         n22701, n22702, n22703, n22705, n22706, n22707, n22708, n22709,
         n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
         n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
         n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
         n22734, n22735, n22736, n22737, n22739, n22740, n22741, n22742,
         n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22779, n22780, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814, n22815, n22816, n22820, n22821,
         n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829,
         n22830, n22831, n22832, n22834, n22835, n22836, n22837, n22838,
         n22839, n22840, n22841, n22842, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22870, n22872, n22873, n22875, n22877,
         n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22886,
         n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894,
         n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902,
         n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910,
         n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918,
         n22919, n22920, n22921, n22922, n22923, n22926, n22927, n22928,
         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22952, n22953, n22954,
         n22955, n22956, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
         n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
         n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23005,
         n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013,
         n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
         n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
         n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037,
         n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045,
         n23046, n23047, n23048, n23049, n23050, n23052, n23053, n23054,
         n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062,
         n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070,
         n23071, n23072, n23073, n23074, n23076, n23077, n23079, n23080,
         n23081, n23082, n23085, n23086, n23087, n23088, n23089, n23090,
         n23091, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23112, n23113, n23114, n23115, n23116,
         n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124,
         n23125, n23126, n23127, n23128, n23129, n23131, n23132, n23133,
         n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
         n23142, n23143, n23145, n23146, n23147, n23148, n23149, n23150,
         n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158,
         n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166,
         n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174,
         n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182,
         n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190,
         n23191, n23193, n23194, n23195, n23196, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23241, n23242,
         n23243, n23244, n23245, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23334, n23335, n23336, n23337, n23338, n23339, n23340,
         n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348,
         n23349, n23350, n23353, n23354, n23355, n23356, n23357, n23358,
         n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366,
         n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374,
         n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382,
         n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390,
         n23391, n23392, n23393, n23394, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23410, n23411, n23413, n23414, n23416, n23417, n23418,
         n23419, n23420, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23458, n23460, n23461,
         n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
         n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477,
         n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
         n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
         n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
         n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
         n23544, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
         n23553, n23554, n23555, n23556, n23557, n23560, n23561, n23562,
         n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
         n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578,
         n23579, n23580, n23581, n23582, n23583, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23594, n23595, n23596,
         n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604,
         n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612,
         n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
         n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628,
         n23629, n23630, n23631, n23632, n23634, n23635, n23636, n23637,
         n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
         n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
         n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661,
         n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
         n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
         n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
         n23686, n23688, n23689, n23690, n23691, n23692, n23693, n23694,
         n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702,
         n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710,
         n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718,
         n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726,
         n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734,
         n23735, n23736, n23737, n23738, n23739, n23740, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23796, n23798, n23799, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23820,
         n23821, n23822, n23823, n23824, n23825, n23827, n23828, n23829,
         n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
         n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23846,
         n23847, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23871, n23872,
         n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23881,
         n23882, n23883, n23885, n23886, n23887, n23888, n23889, n23890,
         n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898,
         n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906,
         n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914,
         n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922,
         n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
         n23931, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23958, n23959, n23960, n23961, n23962, n23963, n23964,
         n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972,
         n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
         n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988,
         n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996,
         n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004,
         n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012,
         n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020,
         n24025, n24026, n24027, n24037, n24042, n24043, n24050, n24051,
         n24054, n24056, n24057, n24059, n24061, n24062, n24063, n24064,
         n24065, n24067, n24072, n24074, n24075, n24076, n24077, n24078,
         n24079, n24080, n24082, n24083, n24084, n24085, n24087, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24103, n24104, n24106, n24107,
         n24108, n24109, n24110, n24112, n24113, n24114, n24115, n24116,
         n24118, n24119, n24120, n24121, n24123, n24124, n24125, n24127,
         n24128, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
         n24137, n24138, n24139, n24140, n24141, n24143, n24144, n24146,
         n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
         n24155, n24158, n24159, n24160, n24161, n24162, n24163, n24164,
         n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
         n24174, n24177, n24178, n24179, n24180, n24181, n24182, n24183,
         n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
         n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
         n24200, n24202, n24203, n24204, n24205, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24217, n24218, n24219, n24220,
         n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24229,
         n24230, n24231, n24233, n24234, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24246, n24247, n24248,
         n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
         n24257, n24258, n24259, n24260, n24261, n24262, n24264, n24265,
         n24267, n24269, n24270, n24272, n24273, n24274, n24275, n24276,
         n24277, n24278, n24279, n24280, n24281, n24283, n24284, n24285,
         n24286, n24287, n24288, n24291, n24292, n24293, n24294, n24295,
         n24296, n24297, n24299, n24300, n24301, n24302, n24303, n24304,
         n24305, n24306, n24307, n24309, n24310, n24311, n24312, n24313,
         n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
         n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24349, n24350, n24351, n24352, n24353, n24354, n24356, n24357,
         n24360, n24361, n24362, n24364, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24383, n24384, n24385, n24386,
         n24387, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24418, n24420, n24421,
         n24422, n24423, n24424, n24426, n24427, n24428, n24429, n24430,
         n24431, n24433, n24434, n24435, n24439, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24451,
         n24452, n24453, n24454, n24456, n24457, n24458, n24459, n24460,
         n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468,
         n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476,
         n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
         n24485, n24486, n24487, n24488, n24490, n24491, n24492, n24493,
         n24494, n24495, n24496, n24498, n24499, n24500, n24501, n24502,
         n24503, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
         n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519,
         n24520, n24521, n24522, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24539, n24540, n24542, n24543, n24547, n24549, n24550, n24551,
         n24552, n24554, n24556, n24558, n24559, n24561, n24565, n24567,
         n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24581, n24582, n24583, n24584,
         n24585, n24586, n24587, n24588, n24589, n24591, n24592, n24594,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
         n24611, n24612, n24613, n24615, n24617, n24618, n24619, n24620,
         n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
         n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636,
         n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644,
         n24646, n24647, n24648, n24650, n24652, n24653, n24654, n24655,
         n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24664,
         n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672,
         n24673, n24674, n24675, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24691, n24692, n24694, n24697, n24698, n24699, n24700, n24701,
         n24702, n24703, n24704, n24706, n24707, n24709, n24710, n24711,
         n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
         n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
         n24728, n24729, n24730, n24733, n24734, n24735, n24736, n24737,
         n24738, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24763, n24764,
         n24765, n24767, n24768, n24769, n24770, n24771, n24772, n24773,
         n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781,
         n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789,
         n24790, n24791, n24792, n24794, n24795, n24796, n24797, n24798,
         n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806,
         n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814,
         n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
         n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
         n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
         n24839, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
         n24848, n24849, n24851, n24852, n24853, n24854, n24855, n24856,
         n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864,
         n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
         n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,
         n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888,
         n24889, n24890, n24891, n24892, n24893, n24895, n24896, n24897,
         n24898, n24899, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24935, n24936, n24937, n24938, n24940, n24941,
         n24942, n24943, n24944, n24946, n24947, n24948, n24949, n24950,
         n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958,
         n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966,
         n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974,
         n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982,
         n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990,
         n24991, n24992, n24993, n24994, n24995, n24996, n24998, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
         n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023,
         n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
         n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
         n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
         n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597;

  BUF_X1 U5 ( .A(n22354), .Z(n245) );
  XNOR2_X1 U8 ( .A(n21451), .B(n21450), .ZN(n22962) );
  XNOR2_X1 U10 ( .A(n21980), .B(n21745), .ZN(n21454) );
  OR2_X1 U16 ( .A1(n20230), .A2(n20498), .ZN(n170) );
  OR2_X1 U17 ( .A1(n20214), .A2(n20215), .ZN(n197) );
  INV_X1 U18 ( .A(n20464), .ZN(n20458) );
  INV_X1 U19 ( .A(n20618), .ZN(n7) );
  OR2_X1 U20 ( .A1(n3428), .A2(n20373), .ZN(n771) );
  INV_X1 U22 ( .A(n20216), .ZN(n100) );
  OR2_X1 U26 ( .A1(n19379), .A2(n19381), .ZN(n4007) );
  OR2_X1 U28 ( .A1(n19381), .A2(n19380), .ZN(n19204) );
  NAND2_X1 U30 ( .A1(n19039), .A2(n24582), .ZN(n194) );
  INV_X1 U36 ( .A(n16037), .ZN(n18516) );
  INV_X1 U40 ( .A(n365), .ZN(n46) );
  INV_X1 U41 ( .A(n17043), .ZN(n17373) );
  INV_X1 U49 ( .A(n3544), .ZN(n41) );
  OR2_X1 U50 ( .A1(n14926), .A2(n16028), .ZN(n161) );
  OR2_X1 U51 ( .A1(n15694), .A2(n16062), .ZN(n15600) );
  INV_X1 U52 ( .A(n16428), .ZN(n15958) );
  XNOR2_X1 U54 ( .A(n15096), .B(n12), .ZN(n15100) );
  INV_X1 U56 ( .A(n15358), .ZN(n75) );
  INV_X1 U57 ( .A(n15422), .ZN(n14442) );
  OR2_X1 U59 ( .A1(n14340), .A2(n25197), .ZN(n76) );
  OR2_X1 U60 ( .A1(n13921), .A2(n13653), .ZN(n96) );
  OR2_X1 U61 ( .A1(n13956), .A2(n13733), .ZN(n813) );
  AND2_X1 U62 ( .A1(n12704), .A2(n14078), .ZN(n13628) );
  AND3_X1 U63 ( .A1(n25435), .A2(n14235), .A3(n24402), .ZN(n182) );
  INV_X1 U66 ( .A(n14209), .ZN(n13811) );
  OR2_X1 U67 ( .A1(n13953), .A2(n24999), .ZN(n507) );
  OR2_X1 U69 ( .A1(n13209), .A2(n13208), .ZN(n136) );
  NAND2_X1 U70 ( .A1(n10395), .A2(n10394), .ZN(n508) );
  AND2_X1 U74 ( .A1(n13222), .A2(n13227), .ZN(n29) );
  AND2_X1 U76 ( .A1(n12454), .A2(n13061), .ZN(n4320) );
  INV_X1 U78 ( .A(n11892), .ZN(n12257) );
  INV_X1 U85 ( .A(n10630), .ZN(n44) );
  OAI21_X1 U86 ( .B1(n11338), .B2(n24082), .A(n10491), .ZN(n11935) );
  OAI211_X1 U90 ( .C1(n25), .C2(n9817), .A(n25046), .B(n24), .ZN(n655) );
  AND2_X1 U93 ( .A1(n25069), .A2(n9886), .ZN(n52) );
  INV_X1 U94 ( .A(n10148), .ZN(n10120) );
  XNOR2_X1 U96 ( .A(n8505), .B(n8504), .ZN(n8521) );
  CLKBUF_X1 U98 ( .A(Key[174]), .Z(n187) );
  NAND2_X1 U104 ( .A1(n7815), .A2(n9070), .ZN(n8507) );
  OR2_X1 U106 ( .A1(n248), .A2(n7232), .ZN(n3192) );
  OR2_X1 U107 ( .A1(n7099), .A2(n127), .ZN(n126) );
  OR2_X1 U108 ( .A1(n7522), .A2(n23), .ZN(n2949) );
  BUF_X1 U110 ( .A(n7057), .Z(n9068) );
  INV_X1 U111 ( .A(n7526), .ZN(n23) );
  MUX2_X1 U115 ( .A(n6107), .B(n6108), .S(n7033), .Z(n7526) );
  AND2_X1 U116 ( .A1(n4672), .A2(n7947), .ZN(n13) );
  OR2_X1 U118 ( .A1(n6945), .A2(n6944), .ZN(n70) );
  AND2_X1 U123 ( .A1(n23252), .A2(n3720), .ZN(n23254) );
  NOR2_X1 U124 ( .A1(n7284), .A2(n7776), .ZN(n7522) );
  NAND2_X1 U127 ( .A1(n17691), .A2(n17690), .ZN(n18004) );
  OR2_X1 U129 ( .A1(n13345), .A2(n12859), .ZN(n13349) );
  INV_X1 U130 ( .A(n22982), .ZN(n22530) );
  AND2_X1 U133 ( .A1(n16449), .A2(n223), .ZN(n131) );
  OR2_X1 U135 ( .A1(n7781), .A2(n7787), .ZN(n5266) );
  NOR2_X1 U137 ( .A1(n22987), .A2(n23379), .ZN(n22988) );
  OR2_X1 U139 ( .A1(n18994), .A2(n20319), .ZN(n615) );
  AND2_X1 U142 ( .A1(n23505), .A2(n3978), .ZN(n23513) );
  NOR2_X1 U145 ( .A1(n23937), .A2(n24948), .ZN(n104) );
  OR2_X1 U147 ( .A1(n22729), .A2(n22093), .ZN(n20893) );
  OR2_X1 U148 ( .A1(n23479), .A2(n23478), .ZN(n22736) );
  NAND2_X1 U156 ( .A1(n17620), .A2(n17623), .ZN(n16901) );
  MUX2_X2 U158 ( .A(n20254), .B(n20253), .S(n21844), .Z(n23860) );
  INV_X1 U162 ( .A(n10168), .ZN(n25) );
  OR2_X1 U163 ( .A1(n10168), .A2(n10169), .ZN(n24) );
  BUF_X1 U164 ( .A(n13453), .Z(n14302) );
  XNOR2_X2 U166 ( .A(n2633), .B(n2634), .ZN(n23014) );
  AND2_X2 U167 ( .A1(n2568), .A2(n2567), .ZN(n2569) );
  OAI21_X1 U170 ( .B1(n10028), .B2(n4787), .A(n9023), .ZN(n10941) );
  OR2_X1 U171 ( .A1(n20183), .A2(n20042), .ZN(n113) );
  XNOR2_X1 U172 ( .A(n11440), .B(n11640), .ZN(n12073) );
  INV_X1 U174 ( .A(n20913), .ZN(n347) );
  OAI22_X1 U178 ( .A1(n10793), .A2(n11196), .B1(n11199), .B2(n10789), .ZN(
        n10628) );
  OR2_X1 U180 ( .A1(n6819), .A2(n6895), .ZN(n190) );
  NAND2_X1 U181 ( .A1(n23393), .A2(n22026), .ZN(n23386) );
  NAND3_X1 U183 ( .A1(n24585), .A2(n16932), .A3(n17054), .ZN(n3593) );
  NAND2_X1 U187 ( .A1(n24589), .A2(n13386), .ZN(n1) );
  NAND2_X1 U188 ( .A1(n13644), .A2(n25011), .ZN(n3) );
  NAND2_X1 U190 ( .A1(n2801), .A2(n4), .ZN(n7829) );
  NAND2_X1 U193 ( .A1(n6), .A2(n5), .ZN(n20088) );
  NAND2_X1 U194 ( .A1(n20084), .A2(n24338), .ZN(n5) );
  NAND2_X1 U195 ( .A1(n8), .A2(n7), .ZN(n6) );
  NAND2_X1 U196 ( .A1(n20570), .A2(n20616), .ZN(n8) );
  NOR2_X1 U198 ( .A1(n25469), .A2(n9), .ZN(n1988) );
  NOR2_X1 U199 ( .A1(n19170), .A2(n19173), .ZN(n9) );
  XNOR2_X1 U202 ( .A(n18044), .B(n17590), .ZN(n10) );
  BUF_X1 U205 ( .A(n6849), .Z(n249) );
  XNOR2_X2 U208 ( .A(n14884), .B(n11), .ZN(n16595) );
  XNOR2_X1 U209 ( .A(n15176), .B(n12451), .ZN(n11) );
  OAI21_X1 U210 ( .B1(n24397), .B2(n23595), .A(n21944), .ZN(n21945) );
  NAND3_X1 U214 ( .A1(n5296), .A2(n10930), .A3(n10596), .ZN(n4213) );
  AOI22_X1 U215 ( .A1(n13813), .A2(n14209), .B1(n3340), .B2(n13422), .ZN(
        n12982) );
  NAND2_X1 U216 ( .A1(n13421), .A2(n1314), .ZN(n14209) );
  NAND2_X1 U218 ( .A1(n4259), .A2(n13), .ZN(n7949) );
  OR2_X2 U220 ( .A1(n2773), .A2(n7951), .ZN(n9149) );
  NAND2_X1 U221 ( .A1(n7035), .A2(n25424), .ZN(n6105) );
  NOR2_X1 U223 ( .A1(n3333), .A2(n3334), .ZN(n14) );
  AOI22_X1 U226 ( .A1(n8841), .A2(n15), .B1(n8842), .B2(n9729), .ZN(n10523) );
  OAI21_X1 U227 ( .B1(n9493), .B2(n426), .A(n9731), .ZN(n15) );
  NAND2_X1 U239 ( .A1(n9558), .A2(n4454), .ZN(n777) );
  NAND3_X1 U240 ( .A1(n13964), .A2(n13962), .A3(n13963), .ZN(n3801) );
  NOR2_X1 U244 ( .A1(n25246), .A2(n17419), .ZN(n17226) );
  NAND2_X1 U247 ( .A1(n3356), .A2(n25292), .ZN(n20) );
  OR2_X1 U248 ( .A1(n13010), .A2(n12919), .ZN(n21) );
  NAND3_X1 U249 ( .A1(n20519), .A2(n351), .A3(n22), .ZN(n73) );
  NAND2_X2 U252 ( .A1(n660), .A2(n9616), .ZN(n11205) );
  AOI22_X2 U257 ( .A1(n20222), .A2(n20272), .B1(n20515), .B2(n20221), .ZN(
        n21568) );
  NAND2_X1 U259 ( .A1(n17267), .A2(n15673), .ZN(n26) );
  NAND2_X1 U260 ( .A1(n16710), .A2(n17326), .ZN(n27) );
  NAND3_X1 U261 ( .A1(n10001), .A2(n10002), .A3(n10000), .ZN(n10004) );
  AOI21_X1 U263 ( .B1(n6782), .B2(n6781), .A(n6780), .ZN(n28) );
  NAND2_X1 U265 ( .A1(n12924), .A2(n29), .ZN(n12571) );
  NAND2_X2 U267 ( .A1(n608), .A2(n9204), .ZN(n10585) );
  XNOR2_X2 U269 ( .A(n5952), .B(Key[169]), .ZN(n6488) );
  NAND2_X1 U270 ( .A1(n12984), .A2(n780), .ZN(n779) );
  NAND3_X1 U272 ( .A1(n4296), .A2(n8026), .A3(n8025), .ZN(n9040) );
  INV_X1 U280 ( .A(n11598), .ZN(n31) );
  OR3_X1 U281 ( .A1(n7909), .A2(n7155), .A3(n7908), .ZN(n7156) );
  XNOR2_X1 U284 ( .A(n15443), .B(n15442), .ZN(n15545) );
  NOR2_X1 U285 ( .A1(n13028), .A2(n13023), .ZN(n11406) );
  NAND2_X1 U286 ( .A1(n34), .A2(n32), .ZN(n13854) );
  NAND2_X1 U287 ( .A1(n12549), .A2(n24220), .ZN(n32) );
  NAND3_X2 U291 ( .A1(n2424), .A2(n12575), .A3(n2423), .ZN(n13845) );
  AND2_X1 U294 ( .A1(n18902), .A2(n18772), .ZN(n762) );
  BUF_X1 U295 ( .A(n9269), .Z(n9947) );
  NAND2_X1 U296 ( .A1(n38), .A2(n24527), .ZN(n14044) );
  NAND2_X1 U298 ( .A1(n3559), .A2(n3558), .ZN(n38) );
  INV_X1 U301 ( .A(n18465), .ZN(n39) );
  AND3_X2 U302 ( .A1(n3251), .A2(n3250), .A3(n3252), .ZN(n11564) );
  NAND2_X1 U304 ( .A1(n42), .A2(n41), .ZN(n40) );
  NAND3_X2 U306 ( .A1(n2750), .A2(n6219), .A3(n2749), .ZN(n8341) );
  NAND2_X1 U312 ( .A1(n9064), .A2(n10050), .ZN(n9539) );
  OR2_X1 U313 ( .A1(n10751), .A2(n10904), .ZN(n10900) );
  OR2_X2 U316 ( .A1(n7244), .A2(n7243), .ZN(n8501) );
  OAI21_X1 U325 ( .B1(n2119), .B2(n6734), .A(n2118), .ZN(n6064) );
  OAI21_X1 U329 ( .B1(n16539), .B2(n17633), .A(n45), .ZN(n16792) );
  MUX2_X2 U331 ( .A(n22971), .B(n22970), .S(n22969), .Z(n23350) );
  XNOR2_X1 U332 ( .A(n47), .B(n2735), .ZN(Ciphertext[74]) );
  NAND3_X1 U333 ( .A1(n4605), .A2(n21955), .A3(n4607), .ZN(n47) );
  NAND2_X2 U335 ( .A1(n9415), .A2(n4655), .ZN(n10767) );
  NAND2_X1 U338 ( .A1(n2821), .A2(n13438), .ZN(n48) );
  OAI21_X1 U346 ( .B1(n52), .B2(n9887), .A(n51), .ZN(n9890) );
  NAND2_X1 U347 ( .A1(n9887), .A2(n9888), .ZN(n51) );
  INV_X1 U356 ( .A(n20291), .ZN(n55) );
  NAND2_X1 U357 ( .A1(n6301), .A2(n6488), .ZN(n6430) );
  NAND2_X1 U361 ( .A1(n17572), .A2(n17042), .ZN(n17043) );
  NAND2_X1 U363 ( .A1(n1148), .A2(n6977), .ZN(n6691) );
  NAND2_X1 U364 ( .A1(n1649), .A2(n10141), .ZN(n1648) );
  XNOR2_X2 U368 ( .A(n5913), .B(Key[18]), .ZN(n5916) );
  NAND2_X1 U369 ( .A1(n13236), .A2(n4499), .ZN(n12937) );
  NAND2_X1 U375 ( .A1(n2922), .A2(n9486), .ZN(n9487) );
  NAND3_X1 U376 ( .A1(n10181), .A2(n58), .A3(n10182), .ZN(n10183) );
  NAND2_X1 U377 ( .A1(n10179), .A2(n10178), .ZN(n58) );
  NAND3_X1 U380 ( .A1(n4846), .A2(n2259), .A3(n16355), .ZN(n2258) );
  NAND2_X1 U382 ( .A1(n13550), .A2(n14210), .ZN(n59) );
  NAND2_X1 U383 ( .A1(n6881), .A2(n6076), .ZN(n6643) );
  NAND2_X1 U384 ( .A1(n60), .A2(n942), .ZN(n941) );
  NAND2_X1 U385 ( .A1(n767), .A2(n6154), .ZN(n60) );
  NOR2_X2 U391 ( .A1(n13087), .A2(n13086), .ZN(n13712) );
  NAND2_X1 U392 ( .A1(n2938), .A2(n2941), .ZN(n13087) );
  OAI21_X1 U393 ( .B1(n3016), .B2(n20498), .A(n61), .ZN(n20270) );
  OAI21_X1 U398 ( .B1(n7228), .B2(n4812), .A(n7947), .ZN(n4811) );
  OR2_X1 U400 ( .A1(n15557), .A2(n25410), .ZN(n15750) );
  AOI22_X2 U404 ( .A1(n1570), .A2(n11038), .B1(n11040), .B2(n11039), .ZN(
        n11983) );
  NOR2_X1 U411 ( .A1(n23462), .A2(n22733), .ZN(n23020) );
  NAND2_X1 U412 ( .A1(n6052), .A2(n6051), .ZN(n6054) );
  NAND3_X1 U413 ( .A1(n16021), .A2(n287), .A3(n16846), .ZN(n16027) );
  NAND3_X1 U415 ( .A1(n7977), .A2(n3567), .A3(n3618), .ZN(n7516) );
  AND3_X2 U418 ( .A1(n1873), .A2(n3613), .A3(n3612), .ZN(n8807) );
  AOI22_X2 U419 ( .A1(n14025), .A2(n13877), .B1(n14334), .B2(n14333), .ZN(
        n13595) );
  NAND2_X1 U420 ( .A1(n66), .A2(n19032), .ZN(n4245) );
  NAND2_X1 U421 ( .A1(n19030), .A2(n19031), .ZN(n66) );
  INV_X1 U422 ( .A(n25215), .ZN(n370) );
  NAND2_X1 U423 ( .A1(n24569), .A2(n25215), .ZN(n5763) );
  AOI21_X2 U431 ( .B1(n7488), .B2(n7487), .A(n7486), .ZN(n9081) );
  XNOR2_X1 U432 ( .A(n68), .B(n2319), .ZN(Ciphertext[11]) );
  OAI211_X1 U433 ( .C1(n23082), .C2(n22578), .A(n23081), .B(n23080), .ZN(n68)
         );
  NAND2_X1 U436 ( .A1(n730), .A2(n3320), .ZN(n7758) );
  NAND2_X1 U438 ( .A1(n2387), .A2(n10884), .ZN(n3416) );
  NAND2_X1 U439 ( .A1(n2597), .A2(n22373), .ZN(n2596) );
  NAND2_X1 U442 ( .A1(n16717), .A2(n69), .ZN(n2823) );
  NAND3_X1 U443 ( .A1(n16715), .A2(n17598), .A3(n17596), .ZN(n69) );
  NAND2_X1 U445 ( .A1(n2996), .A2(n24458), .ZN(n14382) );
  NAND2_X1 U451 ( .A1(n1614), .A2(n1590), .ZN(n71) );
  NAND3_X1 U452 ( .A1(n73), .A2(n1438), .A3(n72), .ZN(n21675) );
  NAND2_X1 U453 ( .A1(n200), .A2(n20272), .ZN(n72) );
  AND2_X1 U455 ( .A1(n22889), .A2(n22093), .ZN(n21774) );
  NAND2_X1 U458 ( .A1(n13501), .A2(n13878), .ZN(n13511) );
  XNOR2_X1 U459 ( .A(n15506), .B(n75), .ZN(n15361) );
  NAND2_X1 U462 ( .A1(n17077), .A2(n17478), .ZN(n16897) );
  NAND3_X2 U466 ( .A1(n16374), .A2(n3775), .A3(n3774), .ZN(n18532) );
  NAND3_X1 U468 ( .A1(n616), .A2(n9071), .A3(n7430), .ZN(n775) );
  NAND2_X1 U469 ( .A1(n16210), .A2(n1496), .ZN(n17387) );
  NAND3_X1 U471 ( .A1(n6171), .A2(n6350), .A3(n6169), .ZN(n77) );
  NAND2_X1 U475 ( .A1(n22678), .A2(n23997), .ZN(n2618) );
  NAND2_X1 U478 ( .A1(n5208), .A2(n20193), .ZN(n5207) );
  NAND3_X1 U481 ( .A1(n10927), .A2(n10924), .A3(n10327), .ZN(n10328) );
  NAND3_X1 U483 ( .A1(n20388), .A2(n19345), .A3(n240), .ZN(n19023) );
  NAND2_X1 U484 ( .A1(n992), .A2(n78), .ZN(n15757) );
  NAND2_X1 U485 ( .A1(n16002), .A2(n16267), .ZN(n78) );
  BUF_X1 U487 ( .A(n5902), .Z(n6950) );
  AOI21_X2 U489 ( .B1(n17410), .B2(n15026), .A(n79), .ZN(n18326) );
  OAI21_X1 U490 ( .B1(n17410), .B2(n17257), .A(n15025), .ZN(n79) );
  XNOR2_X2 U493 ( .A(Key[61]), .B(Plaintext[61]), .ZN(n6963) );
  NAND2_X1 U496 ( .A1(n2767), .A2(n17013), .ZN(n4005) );
  NAND2_X1 U499 ( .A1(n131), .A2(n16236), .ZN(n16237) );
  MUX2_X1 U500 ( .A(n13073), .B(n12532), .S(n13067), .Z(n12475) );
  BUF_X1 U503 ( .A(n7147), .Z(n7699) );
  AND2_X2 U508 ( .A1(n6837), .A2(n467), .ZN(n7989) );
  NAND2_X1 U520 ( .A1(n81), .A2(n6540), .ZN(n6167) );
  NAND2_X1 U521 ( .A1(n5916), .A2(n6162), .ZN(n81) );
  NAND3_X2 U524 ( .A1(n13772), .A2(n82), .A3(n13771), .ZN(n14775) );
  INV_X1 U527 ( .A(n22736), .ZN(n23469) );
  NAND2_X1 U528 ( .A1(n25191), .A2(n12928), .ZN(n1971) );
  NAND3_X2 U529 ( .A1(n3039), .A2(n136), .A3(n13214), .ZN(n13988) );
  NAND3_X2 U531 ( .A1(n7493), .A2(n7491), .A3(n7492), .ZN(n3715) );
  BUF_X1 U535 ( .A(n22575), .Z(n23194) );
  XNOR2_X1 U538 ( .A(n85), .B(n1875), .ZN(Ciphertext[33]) );
  NOR2_X1 U539 ( .A1(n462), .A2(n22576), .ZN(n85) );
  INV_X1 U541 ( .A(n20572), .ZN(n87) );
  XNOR2_X2 U542 ( .A(n14681), .B(n14680), .ZN(n16109) );
  NAND2_X1 U545 ( .A1(n88), .A2(n16124), .ZN(n16127) );
  NAND2_X1 U546 ( .A1(n578), .A2(n381), .ZN(n88) );
  NAND3_X1 U548 ( .A1(n24103), .A2(n7897), .A3(n24861), .ZN(n5235) );
  AOI21_X2 U549 ( .B1(n89), .B2(n10852), .A(n2959), .ZN(n11703) );
  NAND2_X1 U550 ( .A1(n1167), .A2(n10847), .ZN(n89) );
  NAND2_X1 U551 ( .A1(n14028), .A2(n13877), .ZN(n13880) );
  NAND3_X2 U559 ( .A1(n5388), .A2(n1749), .A3(n1405), .ZN(n9188) );
  INV_X1 U560 ( .A(n17099), .ZN(n15869) );
  NAND2_X1 U561 ( .A1(n17120), .A2(n17119), .ZN(n17099) );
  NAND2_X1 U564 ( .A1(n24378), .A2(n20102), .ZN(n21035) );
  INV_X1 U573 ( .A(n11092), .ZN(n11090) );
  NAND2_X1 U574 ( .A1(n95), .A2(n11092), .ZN(n10764) );
  NAND3_X2 U575 ( .A1(n5362), .A2(n9535), .A3(n9534), .ZN(n11092) );
  XNOR2_X1 U577 ( .A(n8541), .B(n8540), .ZN(n9495) );
  OAI211_X2 U587 ( .C1(n15809), .C2(n15808), .A(n15807), .B(n15806), .ZN(
        n18289) );
  NAND3_X2 U588 ( .A1(n13381), .A2(n97), .A3(n96), .ZN(n14620) );
  NAND2_X1 U589 ( .A1(n13985), .A2(n13918), .ZN(n97) );
  NAND2_X1 U592 ( .A1(n25347), .A2(n20216), .ZN(n101) );
  NAND3_X2 U594 ( .A1(n15264), .A2(n3121), .A3(n15265), .ZN(n17342) );
  NAND2_X1 U596 ( .A1(n9487), .A2(n9488), .ZN(n102) );
  XNOR2_X2 U599 ( .A(n5779), .B(Key[91]), .ZN(n6712) );
  NAND2_X1 U600 ( .A1(n3407), .A2(n6277), .ZN(n791) );
  NAND2_X1 U601 ( .A1(n6517), .A2(n315), .ZN(n6277) );
  OAI21_X1 U602 ( .B1(n15783), .B2(n4678), .A(n2478), .ZN(n2891) );
  OAI21_X2 U604 ( .B1(n6387), .B2(n6386), .A(n6385), .ZN(n3979) );
  BUF_X1 U610 ( .A(n19250), .Z(n1551) );
  NAND3_X1 U612 ( .A1(n7718), .A2(n7715), .A3(n24577), .ZN(n7560) );
  NAND2_X1 U613 ( .A1(n23859), .A2(n23843), .ZN(n22982) );
  AOI22_X2 U616 ( .A1(n3191), .A2(n103), .B1(n10077), .B2(n10078), .ZN(n12053)
         );
  INV_X1 U617 ( .A(n11002), .ZN(n103) );
  NAND2_X1 U618 ( .A1(n5342), .A2(n5119), .ZN(n11002) );
  NAND2_X1 U619 ( .A1(n23924), .A2(n104), .ZN(n23915) );
  NAND2_X1 U631 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
  OAI211_X2 U634 ( .C1(n6750), .C2(n6749), .A(n6748), .B(n6747), .ZN(n7674) );
  INV_X1 U640 ( .A(n457), .ZN(n19325) );
  NAND2_X1 U641 ( .A1(n3748), .A2(n17872), .ZN(n457) );
  NAND2_X1 U646 ( .A1(n3302), .A2(n108), .ZN(n3301) );
  OR2_X1 U647 ( .A1(n14156), .A2(n5080), .ZN(n108) );
  XNOR2_X2 U649 ( .A(Key[63]), .B(Plaintext[63]), .ZN(n5800) );
  NAND2_X1 U651 ( .A1(n19244), .A2(n19615), .ZN(n109) );
  NAND3_X1 U654 ( .A1(n12652), .A2(n10360), .A3(n13177), .ZN(n10394) );
  NAND2_X1 U656 ( .A1(n15639), .A2(n16187), .ZN(n2051) );
  BUF_X2 U659 ( .A(n17845), .Z(n19464) );
  NAND3_X1 U660 ( .A1(n3549), .A2(n7500), .A3(n7991), .ZN(n2748) );
  AOI21_X2 U663 ( .B1(n15761), .B2(n3406), .A(n15760), .ZN(n17478) );
  NAND2_X1 U666 ( .A1(n11199), .A2(n10630), .ZN(n4047) );
  XNOR2_X1 U668 ( .A(n15072), .B(n15073), .ZN(n112) );
  NOR2_X1 U670 ( .A1(n16350), .A2(n24467), .ZN(n3333) );
  NAND2_X1 U671 ( .A1(n16597), .A2(n15822), .ZN(n16350) );
  NAND2_X1 U677 ( .A1(n5462), .A2(n16732), .ZN(n3306) );
  NAND2_X1 U679 ( .A1(n19398), .A2(n24326), .ZN(n114) );
  NAND2_X1 U680 ( .A1(n19399), .A2(n18899), .ZN(n115) );
  OAI21_X1 U685 ( .B1(n3655), .B2(n16876), .A(n17356), .ZN(n119) );
  NAND2_X1 U687 ( .A1(n16546), .A2(n17068), .ZN(n16733) );
  AND2_X1 U689 ( .A1(n14124), .A2(n3341), .ZN(n13815) );
  NAND2_X1 U690 ( .A1(n371), .A2(n16578), .ZN(n15538) );
  XNOR2_X1 U693 ( .A(n18466), .B(n16037), .ZN(n18401) );
  NAND3_X2 U694 ( .A1(n10920), .A2(n10921), .A3(n3182), .ZN(n12388) );
  NAND2_X1 U699 ( .A1(n122), .A2(n121), .ZN(n120) );
  INV_X1 U700 ( .A(n6802), .ZN(n121) );
  INV_X1 U701 ( .A(n24772), .ZN(n122) );
  OAI21_X1 U702 ( .B1(n12537), .B2(n14271), .A(n123), .ZN(n2774) );
  INV_X1 U703 ( .A(n13839), .ZN(n123) );
  NAND2_X1 U704 ( .A1(n9633), .A2(n9635), .ZN(n10039) );
  XNOR2_X2 U705 ( .A(n8870), .B(n8871), .ZN(n9635) );
  NOR2_X2 U706 ( .A1(n13007), .A2(n13008), .ZN(n13830) );
  INV_X1 U711 ( .A(n6826), .ZN(n6100) );
  NAND2_X1 U712 ( .A1(n6602), .A2(n7013), .ZN(n6826) );
  NAND3_X2 U714 ( .A1(n6227), .A2(n6228), .A3(n6229), .ZN(n7733) );
  NAND2_X1 U716 ( .A1(n14308), .A2(n14307), .ZN(n13956) );
  NAND2_X1 U718 ( .A1(n4249), .A2(n16002), .ZN(n994) );
  NAND2_X1 U719 ( .A1(n16004), .A2(n25009), .ZN(n4249) );
  OR2_X1 U723 ( .A1(n24470), .A2(n10935), .ZN(n10509) );
  BUF_X1 U724 ( .A(n16431), .Z(n17174) );
  OAI21_X1 U725 ( .B1(n7100), .B2(n126), .A(n125), .ZN(n7105) );
  NAND2_X1 U726 ( .A1(n7103), .A2(n127), .ZN(n125) );
  INV_X1 U727 ( .A(n7101), .ZN(n127) );
  OR2_X2 U729 ( .A1(n6131), .A2(n128), .ZN(n7615) );
  AOI21_X1 U730 ( .B1(n6129), .B2(n6260), .A(n6259), .ZN(n128) );
  NAND2_X1 U733 ( .A1(n6608), .A2(n6712), .ZN(n1925) );
  AND2_X2 U735 ( .A1(n727), .A2(n728), .ZN(n20319) );
  NAND2_X1 U737 ( .A1(n16126), .A2(n24458), .ZN(n129) );
  NAND2_X1 U743 ( .A1(n133), .A2(n24429), .ZN(n17156) );
  NAND2_X1 U745 ( .A1(n16046), .A2(n16045), .ZN(n133) );
  NAND2_X1 U747 ( .A1(n135), .A2(n24093), .ZN(n10375) );
  NAND3_X1 U751 ( .A1(n431), .A2(n7476), .A3(n7477), .ZN(n7425) );
  OR2_X1 U756 ( .A1(n1147), .A2(n6976), .ZN(n6388) );
  XNOR2_X2 U757 ( .A(n5829), .B(Key[134]), .ZN(n6358) );
  NAND2_X1 U759 ( .A1(n7185), .A2(n1862), .ZN(n7246) );
  NAND3_X2 U760 ( .A1(n2308), .A2(n2310), .A3(n2307), .ZN(n11749) );
  NAND2_X2 U763 ( .A1(n12732), .A2(n137), .ZN(n14510) );
  OR2_X2 U765 ( .A1(n16541), .A2(n16542), .ZN(n18659) );
  AOI22_X1 U767 ( .A1(n15945), .A2(n15943), .B1(n16443), .B2(n16440), .ZN(n138) );
  MUX2_X2 U768 ( .A(n9768), .B(n9767), .S(n11163), .Z(n12002) );
  OAI21_X1 U770 ( .B1(n17443), .B2(n17444), .A(n139), .ZN(n17448) );
  NAND2_X1 U772 ( .A1(n6904), .A2(n6902), .ZN(n6903) );
  NAND2_X2 U774 ( .A1(n4813), .A2(n4811), .ZN(n8867) );
  NAND2_X1 U777 ( .A1(n141), .A2(n140), .ZN(n23414) );
  OAI21_X1 U778 ( .B1(n23411), .B2(n24426), .A(n23420), .ZN(n140) );
  NAND2_X1 U779 ( .A1(n23413), .A2(n142), .ZN(n141) );
  NAND2_X1 U781 ( .A1(n7103), .A2(n6165), .ZN(n7098) );
  NAND2_X1 U782 ( .A1(n1611), .A2(n4819), .ZN(n2144) );
  NAND3_X1 U784 ( .A1(n4326), .A2(n11499), .A3(n11058), .ZN(n2152) );
  NAND2_X1 U790 ( .A1(n19380), .A2(n24335), .ZN(n19379) );
  OR2_X1 U791 ( .A1(n25035), .A2(n23411), .ZN(n3157) );
  XNOR2_X1 U796 ( .A(n144), .B(n4153), .ZN(Ciphertext[88]) );
  NAND2_X1 U797 ( .A1(n3156), .A2(n23414), .ZN(n144) );
  NAND3_X1 U798 ( .A1(n145), .A2(n2435), .A3(n10301), .ZN(n2433) );
  NAND2_X1 U799 ( .A1(n2386), .A2(n10302), .ZN(n145) );
  NAND2_X1 U800 ( .A1(n7133), .A2(n146), .ZN(n1848) );
  NAND2_X1 U801 ( .A1(n7132), .A2(n7598), .ZN(n146) );
  AOI21_X2 U802 ( .B1(n12590), .B2(n13350), .A(n2481), .ZN(n14064) );
  NAND3_X1 U805 ( .A1(n17236), .A2(n17237), .A3(n3872), .ZN(n17238) );
  NAND2_X1 U806 ( .A1(n9858), .A2(n238), .ZN(n9861) );
  XNOR2_X1 U810 ( .A(n147), .B(n8539), .ZN(n8540) );
  XNOR2_X1 U811 ( .A(n8891), .B(n8538), .ZN(n147) );
  NOR2_X2 U813 ( .A1(n12812), .A2(n12813), .ZN(n14325) );
  NAND2_X1 U814 ( .A1(n4962), .A2(n4963), .ZN(n12907) );
  OR2_X1 U817 ( .A1(n5992), .A2(n25045), .ZN(n7018) );
  OAI22_X2 U818 ( .A1(n16436), .A2(n16863), .B1(n16435), .B2(n17171), .ZN(
        n18335) );
  NOR2_X2 U829 ( .A1(n9439), .A2(n9438), .ZN(n12108) );
  XNOR2_X1 U830 ( .A(n149), .B(n4873), .ZN(n17606) );
  XNOR2_X1 U831 ( .A(n18183), .B(n18579), .ZN(n149) );
  BUF_X1 U832 ( .A(n9944), .Z(n9897) );
  BUF_X1 U834 ( .A(n5794), .Z(n6623) );
  OR2_X2 U837 ( .A1(n12887), .A2(n12888), .ZN(n14153) );
  INV_X1 U838 ( .A(n17027), .ZN(n17023) );
  NAND2_X1 U839 ( .A1(n17391), .A2(n17185), .ZN(n17027) );
  NAND2_X1 U848 ( .A1(n153), .A2(n152), .ZN(n151) );
  NAND2_X1 U849 ( .A1(n15828), .A2(n1846), .ZN(n152) );
  NAND2_X1 U850 ( .A1(n15829), .A2(n15638), .ZN(n153) );
  NAND2_X1 U855 ( .A1(n14130), .A2(n4844), .ZN(n13896) );
  NAND2_X2 U856 ( .A1(n1564), .A2(n3493), .ZN(n14130) );
  AND2_X2 U861 ( .A1(n10675), .A2(n10673), .ZN(n10985) );
  OAI211_X2 U862 ( .C1(n14058), .C2(n14057), .A(n2756), .B(n155), .ZN(n15119)
         );
  NAND2_X1 U863 ( .A1(n14056), .A2(n14058), .ZN(n155) );
  NAND2_X1 U864 ( .A1(n5863), .A2(n24592), .ZN(n6260) );
  NAND2_X1 U867 ( .A1(n3529), .A2(n3530), .ZN(n156) );
  NAND3_X1 U868 ( .A1(n7209), .A2(n7210), .A3(n2875), .ZN(n9769) );
  NAND2_X1 U869 ( .A1(n17181), .A2(n15907), .ZN(n15645) );
  XNOR2_X2 U874 ( .A(n14095), .B(n14094), .ZN(n16368) );
  NAND2_X1 U875 ( .A1(n158), .A2(n23058), .ZN(n22644) );
  INV_X1 U876 ( .A(n1322), .ZN(n158) );
  NAND2_X1 U877 ( .A1(n322), .A2(n23040), .ZN(n1322) );
  OR2_X2 U879 ( .A1(n5611), .A2(n5610), .ZN(n24012) );
  NOR2_X1 U881 ( .A1(n159), .A2(n23985), .ZN(n23986) );
  NAND2_X1 U882 ( .A1(n4476), .A2(n23984), .ZN(n159) );
  OAI21_X1 U883 ( .B1(n17067), .B2(n17069), .A(n369), .ZN(n723) );
  NAND2_X1 U886 ( .A1(n19646), .A2(n20343), .ZN(n19648) );
  NAND3_X1 U887 ( .A1(n160), .A2(n19104), .A3(n1706), .ZN(n20518) );
  NAND2_X1 U889 ( .A1(n15771), .A2(n161), .ZN(n15770) );
  NAND2_X1 U890 ( .A1(n162), .A2(n6307), .ZN(n7863) );
  NAND2_X1 U891 ( .A1(n909), .A2(n908), .ZN(n162) );
  NAND3_X2 U893 ( .A1(n15732), .A2(n15731), .A3(n468), .ZN(n18382) );
  NAND2_X1 U896 ( .A1(n24570), .A2(n17052), .ZN(n3434) );
  OAI211_X2 U898 ( .C1(n3921), .C2(n24257), .A(n3924), .B(n3920), .ZN(n7380)
         );
  NAND2_X2 U899 ( .A1(n4858), .A2(n3494), .ZN(n17131) );
  NAND2_X1 U900 ( .A1(n5162), .A2(n7237), .ZN(n4020) );
  AND2_X2 U906 ( .A1(n5197), .A2(n5199), .ZN(n10935) );
  XNOR2_X1 U907 ( .A(n15404), .B(n164), .ZN(n15406) );
  XNOR2_X1 U908 ( .A(n15402), .B(n15401), .ZN(n164) );
  NAND3_X1 U916 ( .A1(n3429), .A2(n1582), .A3(n1581), .ZN(n1580) );
  INV_X1 U920 ( .A(n22988), .ZN(n22992) );
  AND3_X2 U929 ( .A1(n1881), .A2(n2956), .A3(n20091), .ZN(n21182) );
  MUX2_X1 U932 ( .A(n5427), .B(n20498), .S(n19824), .Z(n19828) );
  NAND2_X1 U933 ( .A1(n20268), .A2(n1155), .ZN(n19824) );
  NAND2_X1 U935 ( .A1(n17211), .A2(n24529), .ZN(n16880) );
  NAND2_X1 U942 ( .A1(n20227), .A2(n20498), .ZN(n171) );
  NAND2_X1 U943 ( .A1(n172), .A2(n19082), .ZN(n20501) );
  NAND2_X1 U944 ( .A1(n5006), .A2(n5007), .ZN(n172) );
  NAND2_X1 U945 ( .A1(n17068), .A2(n1139), .ZN(n16732) );
  INV_X1 U949 ( .A(n20249), .ZN(n174) );
  NAND2_X1 U950 ( .A1(n19788), .A2(n20241), .ZN(n20248) );
  NAND2_X1 U953 ( .A1(n175), .A2(n5518), .ZN(n5517) );
  NAND2_X1 U954 ( .A1(n787), .A2(n1534), .ZN(n175) );
  NAND2_X1 U959 ( .A1(n13722), .A2(n391), .ZN(n4650) );
  AND2_X2 U967 ( .A1(n2147), .A2(n2146), .ZN(n7908) );
  NAND2_X1 U974 ( .A1(n20383), .A2(n20459), .ZN(n20464) );
  MUX2_X2 U977 ( .A(n19716), .B(n19715), .S(n19714), .Z(n21506) );
  OR2_X2 U978 ( .A1(n6626), .A2(n6627), .ZN(n7789) );
  NOR2_X2 U979 ( .A1(n11075), .A2(n11074), .ZN(n12196) );
  NAND2_X1 U981 ( .A1(n2682), .A2(n4765), .ZN(n178) );
  NAND2_X1 U982 ( .A1(n363), .A2(n19191), .ZN(n19566) );
  OAI21_X1 U983 ( .B1(n20312), .B2(n20125), .A(n179), .ZN(n19967) );
  NAND2_X1 U984 ( .A1(n20125), .A2(n20309), .ZN(n179) );
  XNOR2_X1 U989 ( .A(n180), .B(n20935), .ZN(Ciphertext[152]) );
  NAND4_X1 U990 ( .A1(n4954), .A2(n5732), .A3(n4953), .A4(n21833), .ZN(n180)
         );
  NAND3_X1 U991 ( .A1(n11148), .A2(n11147), .A3(n11143), .ZN(n10962) );
  XNOR2_X1 U992 ( .A(n181), .B(n8936), .ZN(n8939) );
  XNOR2_X1 U993 ( .A(n8937), .B(n9188), .ZN(n181) );
  NOR2_X2 U995 ( .A1(n19800), .A2(n19801), .ZN(n4227) );
  NAND2_X1 U996 ( .A1(n17729), .A2(n16888), .ZN(n17690) );
  NAND2_X1 U997 ( .A1(n9683), .A2(n4069), .ZN(n9686) );
  NOR2_X1 U998 ( .A1(n260), .A2(n10044), .ZN(n9683) );
  NAND2_X1 U999 ( .A1(n19519), .A2(n19522), .ZN(n19525) );
  INV_X1 U1000 ( .A(n7330), .ZN(n5704) );
  NAND2_X1 U1001 ( .A1(n3469), .A2(n7896), .ZN(n7330) );
  AND2_X2 U1003 ( .A1(n4726), .A2(n6197), .ZN(n2624) );
  AOI21_X1 U1005 ( .B1(n14231), .B2(n4560), .A(n182), .ZN(n4558) );
  NAND2_X1 U1010 ( .A1(n12428), .A2(n14315), .ZN(n183) );
  NAND2_X1 U1011 ( .A1(n12427), .A2(n14307), .ZN(n185) );
  OR2_X2 U1013 ( .A1(n7265), .A2(n7264), .ZN(n8899) );
  OR2_X1 U1015 ( .A1(n16809), .A2(n17081), .ZN(n16590) );
  OR2_X1 U1016 ( .A1(n19596), .A2(n18830), .ZN(n19254) );
  NAND2_X1 U1022 ( .A1(n1588), .A2(n22132), .ZN(n22343) );
  NAND2_X1 U1024 ( .A1(n3712), .A2(n16490), .ZN(n15761) );
  NAND2_X1 U1027 ( .A1(n23254), .A2(n189), .ZN(n188) );
  INV_X1 U1028 ( .A(n23256), .ZN(n189) );
  XNOR2_X2 U1031 ( .A(n14610), .B(n14609), .ZN(n16043) );
  OR3_X1 U1032 ( .A1(n9985), .A2(n9980), .A3(n9981), .ZN(n9739) );
  BUF_X1 U1034 ( .A(n6275), .Z(n6517) );
  NAND2_X1 U1039 ( .A1(n17284), .A2(n17293), .ZN(n17540) );
  NAND2_X2 U1040 ( .A1(n2934), .A2(n2935), .ZN(n17284) );
  AND3_X2 U1041 ( .A1(n2698), .A2(n2697), .A3(n2696), .ZN(n21084) );
  NAND3_X2 U1042 ( .A1(n4339), .A2(n22332), .A3(n22331), .ZN(n23165) );
  NAND2_X1 U1043 ( .A1(n12710), .A2(n12707), .ZN(n13074) );
  OAI21_X2 U1047 ( .B1(n1373), .B2(n1406), .A(n4252), .ZN(n11057) );
  NAND3_X1 U1048 ( .A1(n190), .A2(n6893), .A3(n6357), .ZN(n730) );
  NAND2_X1 U1054 ( .A1(n14075), .A2(n396), .ZN(n13851) );
  OAI21_X1 U1059 ( .B1(n19387), .B2(n24477), .A(n191), .ZN(n2706) );
  NAND2_X1 U1061 ( .A1(n10621), .A2(n10620), .ZN(n10622) );
  NAND2_X1 U1062 ( .A1(n232), .A2(n11212), .ZN(n10621) );
  NOR2_X2 U1066 ( .A1(n17200), .A2(n17201), .ZN(n18290) );
  NAND3_X1 U1069 ( .A1(n17572), .A2(n17042), .A3(n17573), .ZN(n15995) );
  NAND2_X2 U1071 ( .A1(n7455), .A2(n5161), .ZN(n9041) );
  NAND3_X1 U1075 ( .A1(n1861), .A2(n25366), .A3(n13345), .ZN(n12575) );
  MUX2_X2 U1082 ( .A(n10418), .B(n10417), .S(n10416), .Z(n11771) );
  NAND2_X1 U1087 ( .A1(n19404), .A2(n24929), .ZN(n19189) );
  NAND2_X1 U1088 ( .A1(n196), .A2(n194), .ZN(n19040) );
  OAI21_X1 U1090 ( .B1(n5233), .B2(n19036), .A(n19037), .ZN(n196) );
  AOI21_X2 U1091 ( .B1(n15998), .B2(n15997), .A(n15996), .ZN(n18312) );
  NAND3_X1 U1104 ( .A1(n197), .A2(n20508), .A3(n25223), .ZN(n4328) );
  NAND4_X2 U1105 ( .A1(n6691), .A2(n4828), .A3(n6689), .A4(n4829), .ZN(n7413)
         );
  XNOR2_X1 U1106 ( .A(Key[6]), .B(Plaintext[6]), .ZN(n6434) );
  OR2_X1 U1107 ( .A1(n11089), .A2(n11297), .ZN(n1058) );
  OR2_X1 U1108 ( .A1(n10451), .A2(n1499), .ZN(n3443) );
  OR2_X1 U1111 ( .A1(n13693), .A2(n13975), .ZN(n14508) );
  OR2_X1 U1114 ( .A1(n17343), .A2(n17241), .ZN(n1284) );
  INV_X1 U1116 ( .A(n19485), .ZN(n5280) );
  AND2_X1 U1119 ( .A1(n23748), .A2(n997), .ZN(n23744) );
  OR2_X1 U1120 ( .A1(n22633), .A2(n2040), .ZN(n509) );
  OR2_X1 U1121 ( .A1(n22634), .A2(n509), .ZN(n22640) );
  AND2_X1 U1122 ( .A1(n6426), .A2(n6467), .ZN(n198) );
  BUF_X1 U1123 ( .A(n6805), .Z(n8530) );
  AND2_X1 U1124 ( .A1(n7128), .A2(n7322), .ZN(n199) );
  AND2_X1 U1125 ( .A1(n20515), .A2(n20517), .ZN(n200) );
  OR2_X1 U1128 ( .A1(n10833), .A2(n9291), .ZN(n201) );
  OR2_X1 U1130 ( .A1(n10296), .A2(n5101), .ZN(n202) );
  OR2_X1 U1132 ( .A1(n10240), .A2(n10496), .ZN(n203) );
  AND3_X1 U1133 ( .A1(n11147), .A2(n11151), .A3(n714), .ZN(n204) );
  AND2_X2 U1135 ( .A1(n10569), .A2(n10568), .ZN(n13954) );
  OR2_X1 U1137 ( .A1(n14002), .A2(n14003), .ZN(n205) );
  OR3_X1 U1140 ( .A1(n17322), .A2(n17321), .A3(n17320), .ZN(n206) );
  OR2_X1 U1141 ( .A1(n17323), .A2(n17324), .ZN(n207) );
  OR3_X1 U1142 ( .A1(n17332), .A2(n17335), .A3(n376), .ZN(n208) );
  AND2_X1 U1145 ( .A1(n18764), .A2(n1475), .ZN(n209) );
  OR2_X1 U1149 ( .A1(n22456), .A2(n22270), .ZN(n211) );
  OR3_X1 U1151 ( .A1(n23839), .A2(n23857), .A3(n24469), .ZN(n212) );
  OR2_X2 U1153 ( .A1(n21871), .A2(n2921), .ZN(n23317) );
  XNOR2_X1 U1155 ( .A(n14561), .B(n14560), .ZN(n16149) );
  XNOR2_X2 U1166 ( .A(n13199), .B(n13198), .ZN(n16597) );
  XNOR2_X2 U1168 ( .A(n8496), .B(n8495), .ZN(n9798) );
  XNOR2_X2 U1169 ( .A(n14878), .B(n14877), .ZN(n15921) );
  XNOR2_X2 U1182 ( .A(n5896), .B(Key[53]), .ZN(n6560) );
  NOR2_X1 U1188 ( .A1(n15617), .A2(n15616), .ZN(n17062) );
  NOR2_X2 U1190 ( .A1(n14037), .A2(n3891), .ZN(n14846) );
  XNOR2_X1 U1198 ( .A(n8136), .B(n8135), .ZN(n9893) );
  AND2_X2 U1199 ( .A1(n3045), .A2(n3044), .ZN(n21591) );
  BUF_X1 U1211 ( .A(n11217), .Z(n232) );
  OAI21_X1 U1212 ( .B1(n5448), .B2(n10093), .A(n10092), .ZN(n11217) );
  NOR2_X1 U1216 ( .A1(n11928), .A2(n11927), .ZN(n14304) );
  XNOR2_X2 U1227 ( .A(n9093), .B(n9094), .ZN(n10060) );
  AND2_X2 U1229 ( .A1(n6092), .A2(n6093), .ZN(n5202) );
  OAI21_X2 U1233 ( .B1(n8384), .B2(n9327), .A(n8383), .ZN(n10931) );
  OAI211_X2 U1236 ( .C1(n7378), .C2(n7641), .A(n2787), .B(n7377), .ZN(n8517)
         );
  XNOR2_X1 U1244 ( .A(n8037), .B(n5157), .ZN(n9859) );
  XNOR2_X1 U1248 ( .A(n4385), .B(n17652), .ZN(n19485) );
  XNOR2_X2 U1256 ( .A(n11533), .B(n11532), .ZN(n12471) );
  XNOR2_X1 U1262 ( .A(n14412), .B(n14411), .ZN(n16428) );
  OR2_X1 U1264 ( .A1(n19596), .A2(n25001), .ZN(n808) );
  XNOR2_X1 U1272 ( .A(n8482), .B(n8481), .ZN(n9997) );
  OAI211_X2 U1273 ( .C1(n7645), .C2(n7736), .A(n7644), .B(n7643), .ZN(n8898)
         );
  XNOR2_X2 U1275 ( .A(Key[183]), .B(Plaintext[183]), .ZN(n6438) );
  AOI21_X2 U1279 ( .B1(n5814), .B2(n6242), .A(n5813), .ZN(n7577) );
  XNOR2_X1 U1281 ( .A(n6000), .B(Key[116]), .ZN(n6849) );
  XNOR2_X2 U1289 ( .A(n8750), .B(n8749), .ZN(n9762) );
  XNOR2_X2 U1297 ( .A(n4610), .B(n4611), .ZN(n3461) );
  BUF_X1 U1304 ( .A(n9255), .Z(n261) );
  OAI211_X1 U1305 ( .C1(n1183), .C2(n9934), .A(n1182), .B(n9933), .ZN(n10245)
         );
  XNOR2_X2 U1310 ( .A(n5943), .B(Key[182]), .ZN(n6174) );
  XNOR2_X1 U1314 ( .A(n21056), .B(n21057), .ZN(n22244) );
  NOR2_X1 U1316 ( .A1(n19510), .A2(n1419), .ZN(n20249) );
  INV_X1 U1319 ( .A(n19310), .ZN(n264) );
  NOR3_X1 U1322 ( .A1(n17576), .A2(n1638), .A3(n1637), .ZN(n17772) );
  INV_X1 U1327 ( .A(n17352), .ZN(n266) );
  INV_X1 U1328 ( .A(n16333), .ZN(n267) );
  INV_X1 U1332 ( .A(n10552), .ZN(n11160) );
  INV_X1 U1334 ( .A(n7591), .ZN(n268) );
  INV_X1 U1336 ( .A(n7965), .ZN(n270) );
  OR2_X1 U1337 ( .A1(n6174), .A2(n4866), .ZN(n6334) );
  INV_X1 U1338 ( .A(n5804), .ZN(n271) );
  CLKBUF_X1 U1340 ( .A(Key[83]), .Z(n2120) );
  CLKBUF_X1 U1341 ( .A(Key[11]), .Z(n1856) );
  CLKBUF_X1 U1343 ( .A(Key[124]), .Z(n765) );
  CLKBUF_X1 U1344 ( .A(Key[18]), .Z(n1833) );
  CLKBUF_X1 U1345 ( .A(Key[92]), .Z(n3183) );
  CLKBUF_X1 U1347 ( .A(Key[108]), .Z(n2834) );
  CLKBUF_X1 U1349 ( .A(Key[24]), .Z(n1865) );
  CLKBUF_X1 U1351 ( .A(Key[59]), .Z(n22886) );
  CLKBUF_X1 U1353 ( .A(Key[56]), .Z(n23679) );
  CLKBUF_X1 U1354 ( .A(Key[144]), .Z(n1952) );
  CLKBUF_X1 U1355 ( .A(Key[154]), .Z(n2744) );
  NOR2_X1 U1356 ( .A1(n24492), .A2(n23361), .ZN(n937) );
  INV_X1 U1357 ( .A(n22395), .ZN(n23292) );
  AND2_X1 U1359 ( .A1(n5223), .A2(n5222), .ZN(n23227) );
  OAI21_X1 U1360 ( .B1(n22503), .B2(n22504), .A(n22502), .ZN(n23442) );
  OAI211_X1 U1363 ( .C1(n22393), .C2(n22958), .A(n2857), .B(n1889), .ZN(n22395) );
  OAI21_X1 U1364 ( .B1(n22966), .B2(n334), .A(n833), .ZN(n22970) );
  OAI21_X1 U1365 ( .B1(n335), .B2(n810), .A(n809), .ZN(n21842) );
  OAI21_X1 U1370 ( .B1(n330), .B2(n25414), .A(n520), .ZN(n3642) );
  XNOR2_X1 U1371 ( .A(n20002), .B(n21083), .ZN(n22228) );
  XNOR2_X1 U1375 ( .A(n20731), .B(n20730), .ZN(n22323) );
  INV_X1 U1377 ( .A(n22449), .ZN(n274) );
  XNOR2_X1 U1378 ( .A(n3871), .B(n20252), .ZN(n22354) );
  OAI21_X1 U1386 ( .B1(n343), .B2(n20269), .A(n1154), .ZN(n19091) );
  OAI21_X1 U1387 ( .B1(n1256), .B2(n345), .A(n1255), .ZN(n20876) );
  OR2_X1 U1389 ( .A1(n20051), .A2(n2168), .ZN(n1072) );
  AND2_X1 U1390 ( .A1(n20338), .A2(n20666), .ZN(n19710) );
  INV_X1 U1393 ( .A(n19875), .ZN(n275) );
  AND2_X1 U1397 ( .A1(n348), .A2(n20479), .ZN(n1023) );
  INV_X1 U1398 ( .A(n20370), .ZN(n277) );
  OR2_X1 U1401 ( .A1(n4075), .A2(n18927), .ZN(n17942) );
  OR2_X1 U1403 ( .A1(n19613), .A2(n355), .ZN(n1805) );
  OR2_X1 U1404 ( .A1(n19360), .A2(n18817), .ZN(n1265) );
  AND2_X1 U1405 ( .A1(n19565), .A2(n19191), .ZN(n1051) );
  AND2_X1 U1406 ( .A1(n363), .A2(n19570), .ZN(n1049) );
  INV_X1 U1408 ( .A(n355), .ZN(n278) );
  XNOR2_X1 U1409 ( .A(n18282), .B(n3753), .ZN(n3773) );
  XNOR2_X1 U1410 ( .A(n18479), .B(n18480), .ZN(n19575) );
  INV_X1 U1412 ( .A(n19543), .ZN(n279) );
  XNOR2_X1 U1414 ( .A(n18321), .B(n18322), .ZN(n19568) );
  XNOR2_X1 U1417 ( .A(n17922), .B(n17923), .ZN(n4748) );
  XNOR2_X1 U1418 ( .A(n17819), .B(n444), .ZN(n17820) );
  XNOR2_X1 U1419 ( .A(n25390), .B(n450), .ZN(n17360) );
  AOI21_X1 U1424 ( .B1(n17143), .B2(n368), .A(n17146), .ZN(n474) );
  AOI22_X1 U1425 ( .A1(n16560), .A2(n17408), .B1(n17613), .B2(n17409), .ZN(
        n16563) );
  OAI211_X1 U1426 ( .C1(n366), .C2(n17473), .A(n17474), .B(n17475), .ZN(n515)
         );
  AND2_X1 U1428 ( .A1(n17044), .A2(n373), .ZN(n16767) );
  INV_X1 U1429 ( .A(n4004), .ZN(n281) );
  CLKBUF_X1 U1430 ( .A(n16527), .Z(n17453) );
  INV_X1 U1431 ( .A(n17173), .ZN(n282) );
  BUF_X1 U1432 ( .A(n16660), .Z(n17031) );
  INV_X1 U1433 ( .A(n1139), .ZN(n283) );
  INV_X1 U1435 ( .A(n17053), .ZN(n284) );
  INV_X1 U1437 ( .A(n17400), .ZN(n285) );
  NAND2_X1 U1440 ( .A1(n15835), .A2(n15836), .ZN(n16888) );
  BUF_X1 U1442 ( .A(n17065), .Z(n369) );
  INV_X1 U1449 ( .A(n17461), .ZN(n287) );
  INV_X1 U1451 ( .A(n15560), .ZN(n16023) );
  CLKBUF_X1 U1455 ( .A(n15710), .Z(n16438) );
  INV_X1 U1458 ( .A(n16334), .ZN(n290) );
  INV_X1 U1459 ( .A(n16042), .ZN(n291) );
  XNOR2_X1 U1463 ( .A(n14723), .B(n14722), .ZN(n15584) );
  INV_X1 U1464 ( .A(n16149), .ZN(n293) );
  XNOR2_X1 U1465 ( .A(n13499), .B(n13498), .ZN(n16332) );
  XNOR2_X1 U1466 ( .A(n14969), .B(n14968), .ZN(n16451) );
  XNOR2_X1 U1468 ( .A(n14979), .B(n14919), .ZN(n1091) );
  INV_X1 U1471 ( .A(n14997), .ZN(n295) );
  OAI21_X1 U1472 ( .B1(n14123), .B2(n14208), .A(n2214), .ZN(n14210) );
  AND2_X1 U1473 ( .A1(n394), .A2(n13951), .ZN(n749) );
  INV_X1 U1474 ( .A(n4844), .ZN(n14132) );
  INV_X1 U1475 ( .A(n14034), .ZN(n296) );
  INV_X1 U1476 ( .A(n14149), .ZN(n297) );
  INV_X1 U1477 ( .A(n14044), .ZN(n298) );
  INV_X1 U1478 ( .A(n13488), .ZN(n299) );
  NAND3_X1 U1480 ( .A1(n12422), .A2(n1086), .A3(n1087), .ZN(n13900) );
  INV_X1 U1483 ( .A(n13847), .ZN(n300) );
  OR2_X1 U1485 ( .A1(n12483), .A2(n12715), .ZN(n4057) );
  INV_X1 U1487 ( .A(n13328), .ZN(n301) );
  XNOR2_X1 U1488 ( .A(n12044), .B(n12043), .ZN(n2295) );
  OR2_X1 U1489 ( .A1(n13056), .A2(n13057), .ZN(n11438) );
  INV_X1 U1491 ( .A(n12784), .ZN(n302) );
  INV_X1 U1492 ( .A(n12796), .ZN(n303) );
  XNOR2_X1 U1493 ( .A(n12290), .B(n12289), .ZN(n13114) );
  INV_X1 U1496 ( .A(n4766), .ZN(n304) );
  XNOR2_X1 U1499 ( .A(n11977), .B(n11295), .ZN(n12114) );
  OR2_X1 U1504 ( .A1(n11101), .A2(n10914), .ZN(n10220) );
  NOR2_X1 U1506 ( .A1(n11342), .A2(n10632), .ZN(n10491) );
  AND2_X1 U1507 ( .A1(n10891), .A2(n10889), .ZN(n10438) );
  INV_X1 U1511 ( .A(n11122), .ZN(n305) );
  XNOR2_X1 U1518 ( .A(n7550), .B(n7549), .ZN(n9281) );
  INV_X1 U1519 ( .A(n1595), .ZN(n3292) );
  INV_X1 U1523 ( .A(n10061), .ZN(n309) );
  XNOR2_X1 U1524 ( .A(n9105), .B(n9104), .ZN(n9127) );
  INV_X1 U1526 ( .A(n8818), .ZN(n310) );
  OR2_X1 U1530 ( .A1(n8008), .A2(n8007), .ZN(n8970) );
  AND4_X1 U1531 ( .A1(n1195), .A2(n1190), .A3(n1191), .A4(n1193), .ZN(n1110)
         );
  BUF_X1 U1532 ( .A(n7108), .Z(n7532) );
  INV_X1 U1534 ( .A(n7609), .ZN(n311) );
  BUF_X1 U1535 ( .A(n7589), .Z(n7462) );
  CLKBUF_X1 U1536 ( .A(n7409), .Z(n7982) );
  INV_X1 U1540 ( .A(n7917), .ZN(n312) );
  INV_X1 U1543 ( .A(n1147), .ZN(n6687) );
  CLKBUF_X1 U1545 ( .A(n6066), .Z(n6688) );
  XNOR2_X1 U1548 ( .A(n5803), .B(Key[67]), .ZN(n5804) );
  CLKBUF_X1 U1549 ( .A(n6400), .Z(n6755) );
  CLKBUF_X1 U1550 ( .A(n6648), .Z(n7011) );
  INV_X1 U1552 ( .A(n6358), .ZN(n313) );
  CLKBUF_X1 U1555 ( .A(Key[109]), .Z(n925) );
  CLKBUF_X1 U1556 ( .A(Key[81]), .Z(n3062) );
  CLKBUF_X1 U1557 ( .A(Key[110]), .Z(n2049) );
  CLKBUF_X1 U1558 ( .A(Key[67]), .Z(n494) );
  CLKBUF_X1 U1559 ( .A(Key[126]), .Z(n1745) );
  CLKBUF_X1 U1560 ( .A(Key[123]), .Z(n21662) );
  CLKBUF_X1 U1562 ( .A(Key[177]), .Z(n20284) );
  CLKBUF_X1 U1563 ( .A(Key[170]), .Z(n1777) );
  CLKBUF_X1 U1565 ( .A(Key[31]), .Z(n2726) );
  CLKBUF_X1 U1568 ( .A(Key[128]), .Z(n2746) );
  CLKBUF_X1 U1569 ( .A(Key[125]), .Z(n2881) );
  CLKBUF_X1 U1570 ( .A(Key[88]), .Z(n891) );
  CLKBUF_X1 U1572 ( .A(Key[133]), .Z(n2826) );
  CLKBUF_X1 U1573 ( .A(Key[9]), .Z(n19392) );
  CLKBUF_X1 U1574 ( .A(Key[114]), .Z(n2211) );
  CLKBUF_X1 U1575 ( .A(Key[7]), .Z(n2222) );
  CLKBUF_X1 U1576 ( .A(Key[121]), .Z(n2145) );
  CLKBUF_X1 U1577 ( .A(Key[165]), .Z(n924) );
  CLKBUF_X1 U1578 ( .A(Key[21]), .Z(n17960) );
  CLKBUF_X1 U1579 ( .A(Key[160]), .Z(n1754) );
  CLKBUF_X1 U1580 ( .A(Key[135]), .Z(n3129) );
  CLKBUF_X1 U1582 ( .A(Key[129]), .Z(n876) );
  CLKBUF_X1 U1584 ( .A(Key[77]), .Z(n681) );
  CLKBUF_X1 U1585 ( .A(Key[118]), .Z(n3118) );
  CLKBUF_X1 U1586 ( .A(Key[104]), .Z(n3089) );
  CLKBUF_X1 U1587 ( .A(Key[130]), .Z(n2739) );
  CLKBUF_X1 U1588 ( .A(Key[70]), .Z(n663) );
  CLKBUF_X1 U1589 ( .A(Key[112]), .Z(n2126) );
  CLKBUF_X1 U1590 ( .A(Key[1]), .Z(n2805) );
  CLKBUF_X1 U1591 ( .A(Key[42]), .Z(n2761) );
  CLKBUF_X1 U1592 ( .A(Key[171]), .Z(n20690) );
  CLKBUF_X1 U1593 ( .A(Key[49]), .Z(n1827) );
  CLKBUF_X1 U1594 ( .A(Key[143]), .Z(n20609) );
  CLKBUF_X1 U1596 ( .A(Key[178]), .Z(n896) );
  CLKBUF_X1 U1598 ( .A(Key[39]), .Z(n2039) );
  CLKBUF_X1 U1599 ( .A(Key[17]), .Z(n1869) );
  CLKBUF_X1 U1602 ( .A(Key[52]), .Z(n1746) );
  CLKBUF_X1 U1603 ( .A(Key[22]), .Z(n1797) );
  CLKBUF_X1 U1604 ( .A(Key[95]), .Z(n14398) );
  CLKBUF_X1 U1606 ( .A(Key[147]), .Z(n1724) );
  CLKBUF_X1 U1610 ( .A(Key[16]), .Z(n853) );
  CLKBUF_X1 U1611 ( .A(Key[163]), .Z(n1757) );
  CLKBUF_X1 U1613 ( .A(Key[111]), .Z(n21204) );
  CLKBUF_X1 U1615 ( .A(Key[141]), .Z(n1804) );
  CLKBUF_X1 U1616 ( .A(Key[103]), .Z(n1951) );
  CLKBUF_X1 U1617 ( .A(Key[148]), .Z(n812) );
  CLKBUF_X1 U1618 ( .A(Key[120]), .Z(n3084) );
  CLKBUF_X1 U1619 ( .A(Key[127]), .Z(n1815) );
  CLKBUF_X1 U1620 ( .A(Key[76]), .Z(n2772) );
  CLKBUF_X1 U1622 ( .A(Key[71]), .Z(n2240) );
  CLKBUF_X1 U1623 ( .A(Key[85]), .Z(n2241) );
  CLKBUF_X1 U1624 ( .A(Key[69]), .Z(n860) );
  CLKBUF_X1 U1625 ( .A(Key[62]), .Z(n1863) );
  CLKBUF_X1 U1626 ( .A(Key[55]), .Z(n1739) );
  CLKBUF_X1 U1627 ( .A(Key[5]), .Z(n2991) );
  CLKBUF_X1 U1628 ( .A(Key[84]), .Z(n2193) );
  CLKBUF_X1 U1629 ( .A(Key[173]), .Z(n3158) );
  CLKBUF_X1 U1630 ( .A(Key[159]), .Z(n2044) );
  CLKBUF_X1 U1631 ( .A(Key[145]), .Z(n1792) );
  CLKBUF_X1 U1632 ( .A(Key[19]), .Z(n1835) );
  CLKBUF_X1 U1634 ( .A(Key[138]), .Z(n1801) );
  CLKBUF_X1 U1635 ( .A(Key[96]), .Z(n2717) );
  CLKBUF_X1 U1636 ( .A(Key[180]), .Z(n912) );
  CLKBUF_X1 U1637 ( .A(Key[47]), .Z(n889) );
  CLKBUF_X1 U1639 ( .A(Key[155]), .Z(n2989) );
  INV_X1 U1640 ( .A(n6521), .ZN(n315) );
  CLKBUF_X1 U1641 ( .A(Key[75]), .Z(n2882) );
  CLKBUF_X1 U1642 ( .A(Key[169]), .Z(n899) );
  CLKBUF_X1 U1644 ( .A(Key[162]), .Z(n921) );
  CLKBUF_X1 U1645 ( .A(Key[153]), .Z(n1891) );
  CLKBUF_X1 U1646 ( .A(Key[139]), .Z(n1810) );
  CLKBUF_X1 U1648 ( .A(Key[191]), .Z(n2847) );
  INV_X1 U1649 ( .A(n6243), .ZN(n316) );
  CLKBUF_X1 U1650 ( .A(Key[34]), .Z(n1789) );
  CLKBUF_X1 U1651 ( .A(Key[6]), .Z(n21623) );
  CLKBUF_X1 U1652 ( .A(Key[27]), .Z(n763) );
  CLKBUF_X1 U1653 ( .A(Key[188]), .Z(n3131) );
  CLKBUF_X1 U1654 ( .A(Key[10]), .Z(n20995) );
  CLKBUF_X1 U1655 ( .A(Key[181]), .Z(n1767) );
  CLKBUF_X1 U1658 ( .A(Key[80]), .Z(n2236) );
  CLKBUF_X1 U1659 ( .A(Key[86]), .Z(n3178) );
  CLKBUF_X1 U1660 ( .A(Key[72]), .Z(n1758) );
  CLKBUF_X1 U1661 ( .A(Key[73]), .Z(n881) );
  CLKBUF_X1 U1663 ( .A(Key[65]), .Z(n20046) );
  CLKBUF_X1 U1665 ( .A(Key[51]), .Z(n2087) );
  CLKBUF_X1 U1666 ( .A(Key[66]), .Z(n2990) );
  CLKBUF_X1 U1667 ( .A(Key[12]), .Z(n2208) );
  CLKBUF_X1 U1668 ( .A(Key[87]), .Z(n1826) );
  CLKBUF_X1 U1669 ( .A(Key[23]), .Z(n2190) );
  CLKBUF_X1 U1670 ( .A(Key[36]), .Z(n1364) );
  CLKBUF_X1 U1671 ( .A(Key[78]), .Z(n1924) );
  CLKBUF_X1 U1672 ( .A(Key[43]), .Z(n1768) );
  CLKBUF_X1 U1673 ( .A(Key[50]), .Z(n2005) );
  NOR2_X1 U1674 ( .A1(n23511), .A2(n23512), .ZN(n23522) );
  OAI211_X1 U1675 ( .C1(n23965), .C2(n23964), .A(n23963), .B(n878), .ZN(n3150)
         );
  OR2_X1 U1676 ( .A1(n23728), .A2(n23727), .ZN(n786) );
  OR2_X1 U1677 ( .A1(n22531), .A2(n22532), .ZN(n852) );
  OR2_X1 U1678 ( .A1(n23692), .A2(n23689), .ZN(n1145) );
  NOR2_X1 U1679 ( .A1(n23619), .A2(n23634), .ZN(n23652) );
  NOR2_X1 U1680 ( .A1(n23292), .A2(n23303), .ZN(n23298) );
  INV_X1 U1682 ( .A(n23311), .ZN(n4108) );
  AND2_X1 U1683 ( .A1(n23911), .A2(n23924), .ZN(n23941) );
  AND2_X1 U1687 ( .A1(n1683), .A2(n1686), .ZN(n23327) );
  BUF_X1 U1694 ( .A(n24010), .Z(n23982) );
  OAI21_X1 U1696 ( .B1(n21378), .B2(n25543), .A(n5048), .ZN(n22442) );
  INV_X1 U1699 ( .A(n23227), .ZN(n317) );
  INV_X1 U1701 ( .A(n23810), .ZN(n318) );
  AND3_X1 U1702 ( .A1(n5422), .A2(n5419), .A3(n1397), .ZN(n23361) );
  INV_X1 U1703 ( .A(n21863), .ZN(n23903) );
  OAI21_X1 U1705 ( .B1(n22497), .B2(n4719), .A(n2364), .ZN(n23443) );
  INV_X1 U1711 ( .A(n23442), .ZN(n321) );
  INV_X1 U1713 ( .A(n22698), .ZN(n322) );
  INV_X1 U1714 ( .A(n23972), .ZN(n878) );
  AND3_X1 U1716 ( .A1(n4781), .A2(n1691), .A3(n22729), .ZN(n23517) );
  OAI21_X1 U1719 ( .B1(n4591), .B2(n22408), .A(n24951), .ZN(n22414) );
  INV_X1 U1720 ( .A(n23543), .ZN(n323) );
  OAI21_X1 U1723 ( .B1(n20980), .B2(n20979), .A(n24902), .ZN(n1007) );
  AND2_X1 U1725 ( .A1(n22808), .A2(n4427), .ZN(n23993) );
  INV_X1 U1726 ( .A(n24879), .ZN(n324) );
  OR2_X1 U1728 ( .A1(n24951), .A2(n22565), .ZN(n650) );
  OR2_X1 U1729 ( .A1(n22953), .A2(n21878), .ZN(n1257) );
  OR2_X1 U1730 ( .A1(n22034), .A2(n24884), .ZN(n1258) );
  AND2_X1 U1731 ( .A1(n22667), .A2(n22670), .ZN(n919) );
  INV_X1 U1732 ( .A(n22219), .ZN(n22217) );
  OR2_X1 U1733 ( .A1(n4468), .A2(n4467), .ZN(n481) );
  INV_X1 U1734 ( .A(n3781), .ZN(n1686) );
  OR2_X1 U1736 ( .A1(n22322), .A2(n22456), .ZN(n22327) );
  NOR2_X1 U1737 ( .A1(n21802), .A2(n22198), .ZN(n23634) );
  INV_X1 U1738 ( .A(n22356), .ZN(n21348) );
  AND2_X1 U1741 ( .A1(n25082), .A2(n22361), .ZN(n1249) );
  OR2_X1 U1742 ( .A1(n21841), .A2(n22257), .ZN(n810) );
  OR2_X1 U1744 ( .A1(n22426), .A2(n2674), .ZN(n776) );
  XNOR2_X1 U1745 ( .A(n20783), .B(n20782), .ZN(n5084) );
  XNOR2_X1 U1746 ( .A(n20746), .B(n20745), .ZN(n22454) );
  OR2_X1 U1747 ( .A1(n21856), .A2(n22769), .ZN(n534) );
  OR2_X1 U1749 ( .A1(n21792), .A2(n3231), .ZN(n1163) );
  OR2_X1 U1751 ( .A1(n22261), .A2(n22398), .ZN(n22262) );
  INV_X1 U1752 ( .A(n2601), .ZN(n1146) );
  OR2_X1 U1753 ( .A1(n22056), .A2(n21836), .ZN(n1310) );
  CLKBUF_X1 U1757 ( .A(n21766), .Z(n22206) );
  INV_X1 U1758 ( .A(n22953), .ZN(n1293) );
  INV_X1 U1759 ( .A(n23574), .ZN(n325) );
  INV_X1 U1760 ( .A(n24971), .ZN(n326) );
  XNOR2_X1 U1761 ( .A(n21006), .B(n21007), .ZN(n22926) );
  AND2_X1 U1764 ( .A1(n4273), .A2(n22655), .ZN(n22811) );
  CLKBUF_X1 U1766 ( .A(n21265), .Z(n22614) );
  INV_X1 U1767 ( .A(n22888), .ZN(n327) );
  INV_X1 U1769 ( .A(n22228), .ZN(n328) );
  CLKBUF_X1 U1772 ( .A(n21759), .Z(n22197) );
  INV_X1 U1773 ( .A(n22323), .ZN(n329) );
  XNOR2_X1 U1774 ( .A(n20083), .B(n20082), .ZN(n22355) );
  INV_X1 U1777 ( .A(n23999), .ZN(n330) );
  XNOR2_X1 U1779 ( .A(n20988), .B(n20987), .ZN(n22715) );
  INV_X1 U1780 ( .A(n22657), .ZN(n331) );
  INV_X1 U1781 ( .A(n22257), .ZN(n332) );
  INV_X1 U1782 ( .A(n21934), .ZN(n333) );
  INV_X1 U1784 ( .A(n22968), .ZN(n334) );
  XNOR2_X1 U1785 ( .A(n21595), .B(n21594), .ZN(n22033) );
  XNOR2_X1 U1786 ( .A(n20642), .B(n20643), .ZN(n22333) );
  CLKBUF_X1 U1790 ( .A(n21209), .Z(n20634) );
  INV_X1 U1791 ( .A(n22252), .ZN(n335) );
  INV_X1 U1792 ( .A(n22222), .ZN(n336) );
  XNOR2_X1 U1793 ( .A(n21180), .B(n21179), .ZN(n22448) );
  INV_X1 U1794 ( .A(n22832), .ZN(n337) );
  INV_X1 U1795 ( .A(n22965), .ZN(n338) );
  XNOR2_X1 U1796 ( .A(n21621), .B(n21985), .ZN(n20957) );
  XNOR2_X1 U1797 ( .A(n21176), .B(n20594), .ZN(n21562) );
  XNOR2_X1 U1798 ( .A(n1153), .B(n20904), .ZN(n21496) );
  XNOR2_X1 U1799 ( .A(n21569), .B(n21402), .ZN(n21246) );
  XNOR2_X1 U1800 ( .A(n21688), .B(n596), .ZN(n21690) );
  NAND3_X1 U1802 ( .A1(n19048), .A2(n19050), .A3(n19049), .ZN(n20870) );
  XNOR2_X1 U1803 ( .A(n21687), .B(n21689), .ZN(n596) );
  OAI21_X1 U1814 ( .B1(n19706), .B2(n20614), .A(n19705), .ZN(n21975) );
  AND3_X1 U1815 ( .A1(n4183), .A2(n20266), .A3(n20265), .ZN(n4185) );
  MUX2_X1 U1820 ( .A(n21009), .B(n24581), .S(n20289), .Z(n20295) );
  OAI211_X1 U1824 ( .C1(n19939), .C2(n24077), .A(n3650), .B(n19339), .ZN(
        n21106) );
  OR2_X1 U1825 ( .A1(n20592), .A2(n20593), .ZN(n2362) );
  OAI21_X1 U1826 ( .B1(n636), .B2(n20527), .A(n20526), .ZN(n21013) );
  NOR2_X1 U1829 ( .A1(n20074), .A2(n19855), .ZN(n588) );
  NAND2_X1 U1831 ( .A1(n19938), .A2(n19939), .ZN(n2946) );
  AND2_X1 U1832 ( .A1(n20255), .A2(n19743), .ZN(n1256) );
  INV_X1 U1833 ( .A(n19511), .ZN(n754) );
  OR2_X1 U1834 ( .A1(n24076), .A2(n20616), .ZN(n19703) );
  AOI22_X1 U1835 ( .A1(n20478), .A2(n1024), .B1(n1023), .B2(n20480), .ZN(n1022) );
  INV_X1 U1836 ( .A(n20191), .ZN(n1242) );
  INV_X1 U1837 ( .A(n19743), .ZN(n2024) );
  INV_X1 U1840 ( .A(n19984), .ZN(n885) );
  AND2_X1 U1842 ( .A1(n20578), .A2(n20576), .ZN(n1205) );
  OR2_X1 U1843 ( .A1(n20165), .A2(n20395), .ZN(n2426) );
  OR2_X1 U1844 ( .A1(n1591), .A2(n17943), .ZN(n21031) );
  INV_X1 U1845 ( .A(n17943), .ZN(n21033) );
  INV_X1 U1847 ( .A(n20262), .ZN(n20409) );
  INV_X1 U1849 ( .A(n19887), .ZN(n339) );
  NAND2_X1 U1850 ( .A1(n1716), .A2(n1421), .ZN(n20094) );
  AND2_X1 U1851 ( .A1(n20523), .A2(n20522), .ZN(n21009) );
  NAND2_X1 U1853 ( .A1(n1980), .A2(n18394), .ZN(n20022) );
  OR2_X1 U1854 ( .A1(n19619), .A2(n19618), .ZN(n594) );
  INV_X1 U1856 ( .A(n20319), .ZN(n340) );
  NOR2_X1 U1857 ( .A1(n20142), .A2(n19975), .ZN(n19680) );
  BUF_X1 U1858 ( .A(n19774), .Z(n20384) );
  AND3_X1 U1859 ( .A1(n4916), .A2(n2983), .A3(n4915), .ZN(n17567) );
  NOR2_X1 U1860 ( .A1(n20497), .A2(n20498), .ZN(n20502) );
  NAND2_X1 U1865 ( .A1(n18547), .A2(n3055), .ZN(n20614) );
  INV_X1 U1867 ( .A(n20055), .ZN(n19928) );
  INV_X1 U1868 ( .A(n20317), .ZN(n341) );
  AOI21_X1 U1869 ( .B1(n19529), .B2(n1013), .A(n1011), .ZN(n1010) );
  AND2_X1 U1871 ( .A1(n3277), .A2(n3989), .ZN(n818) );
  NAND2_X1 U1873 ( .A1(n5646), .A2(n18827), .ZN(n20476) );
  INV_X1 U1876 ( .A(n20498), .ZN(n343) );
  INV_X1 U1880 ( .A(n20413), .ZN(n345) );
  INV_X1 U1883 ( .A(n20214), .ZN(n20199) );
  INV_X1 U1886 ( .A(n20909), .ZN(n346) );
  OAI21_X1 U1887 ( .B1(n1046), .B2(n1050), .A(n1048), .ZN(n20214) );
  INV_X1 U1891 ( .A(n20353), .ZN(n348) );
  OR2_X1 U1892 ( .A1(n17554), .A2(n19531), .ZN(n1015) );
  NAND2_X1 U1893 ( .A1(n19533), .A2(n19531), .ZN(n1016) );
  INV_X1 U1894 ( .A(n20367), .ZN(n349) );
  OR2_X1 U1895 ( .A1(n18443), .A2(n19164), .ZN(n1977) );
  AOI22_X1 U1896 ( .A1(n1001), .A2(n280), .B1(n19576), .B2(n25072), .ZN(n1000)
         );
  OAI21_X1 U1897 ( .B1(n19629), .B2(n4543), .A(n3379), .ZN(n19840) );
  OR2_X1 U1898 ( .A1(n1107), .A2(n264), .ZN(n1160) );
  INV_X1 U1899 ( .A(n20460), .ZN(n350) );
  INV_X1 U1900 ( .A(n20515), .ZN(n351) );
  NOR2_X1 U1901 ( .A1(n24982), .A2(n1002), .ZN(n1001) );
  INV_X1 U1902 ( .A(n19007), .ZN(n1005) );
  XNOR2_X1 U1903 ( .A(n4890), .B(n18384), .ZN(n18597) );
  AND2_X1 U1904 ( .A1(n1052), .A2(n5634), .ZN(n1050) );
  AND2_X1 U1905 ( .A1(n1051), .A2(n1047), .ZN(n1046) );
  AOI21_X1 U1906 ( .B1(n19269), .B2(n19534), .A(n4172), .ZN(n1012) );
  NAND2_X1 U1907 ( .A1(n1291), .A2(n19435), .ZN(n1290) );
  OR2_X1 U1908 ( .A1(n19435), .A2(n18833), .ZN(n1287) );
  BUF_X1 U1909 ( .A(n18772), .Z(n19125) );
  AND2_X1 U1912 ( .A1(n18788), .A2(n19397), .ZN(n18900) );
  NAND3_X1 U1913 ( .A1(n19060), .A2(n19059), .A3(n19007), .ZN(n19062) );
  AND2_X1 U1921 ( .A1(n4436), .A2(n1300), .ZN(n4435) );
  OR2_X1 U1922 ( .A1(n19311), .A2(n19309), .ZN(n696) );
  INV_X1 U1923 ( .A(n19186), .ZN(n19404) );
  INV_X1 U1924 ( .A(n19421), .ZN(n1306) );
  AND2_X1 U1925 ( .A1(n19419), .A2(n19420), .ZN(n1307) );
  AND2_X1 U1926 ( .A1(n988), .A2(n24982), .ZN(n1443) );
  XNOR2_X1 U1928 ( .A(n17647), .B(n17646), .ZN(n19490) );
  INV_X1 U1931 ( .A(n19487), .ZN(n352) );
  INV_X1 U1934 ( .A(n3773), .ZN(n353) );
  INV_X1 U1935 ( .A(n19575), .ZN(n354) );
  INV_X1 U1936 ( .A(n19238), .ZN(n355) );
  XNOR2_X1 U1938 ( .A(n17508), .B(n17507), .ZN(n19300) );
  INV_X1 U1939 ( .A(n19126), .ZN(n19543) );
  INV_X1 U1940 ( .A(n19418), .ZN(n19419) );
  INV_X1 U1941 ( .A(n19296), .ZN(n356) );
  INV_X1 U1942 ( .A(n19502), .ZN(n357) );
  XNOR2_X1 U1945 ( .A(n18427), .B(n18426), .ZN(n19162) );
  XNOR2_X1 U1947 ( .A(n16939), .B(n16938), .ZN(n19311) );
  INV_X1 U1948 ( .A(n19273), .ZN(n1053) );
  XNOR2_X1 U1949 ( .A(n18625), .B(n18624), .ZN(n19441) );
  INV_X1 U1950 ( .A(n19500), .ZN(n358) );
  INV_X1 U1954 ( .A(n19570), .ZN(n960) );
  XNOR2_X1 U1955 ( .A(n18462), .B(n18461), .ZN(n988) );
  OR2_X1 U1957 ( .A1(n19568), .A2(n19192), .ZN(n1047) );
  XNOR2_X1 U1960 ( .A(n4274), .B(n16626), .ZN(n19559) );
  INV_X1 U1962 ( .A(n18832), .ZN(n361) );
  XNOR2_X1 U1963 ( .A(n18273), .B(n18274), .ZN(n19126) );
  XNOR2_X1 U1964 ( .A(n18699), .B(n18698), .ZN(n19407) );
  XNOR2_X1 U1966 ( .A(n17308), .B(n17307), .ZN(n19329) );
  XNOR2_X1 U1969 ( .A(n18632), .B(n18631), .ZN(n19438) );
  XNOR2_X1 U1972 ( .A(n18379), .B(n18378), .ZN(n19428) );
  INV_X1 U1973 ( .A(n19568), .ZN(n362) );
  INV_X1 U1974 ( .A(n19192), .ZN(n363) );
  XNOR2_X1 U1975 ( .A(n17787), .B(n17786), .ZN(n19370) );
  XNOR2_X1 U1977 ( .A(n17874), .B(n3725), .ZN(n966) );
  XNOR2_X1 U1978 ( .A(n17638), .B(n17637), .ZN(n18051) );
  XNOR2_X1 U1980 ( .A(n18334), .B(n18407), .ZN(n17648) );
  XNOR2_X1 U1981 ( .A(n934), .B(n25411), .ZN(n18683) );
  AOI22_X1 U1982 ( .A1(n4267), .A2(n4266), .B1(n16610), .B2(n17054), .ZN(
        n17933) );
  XNOR2_X1 U1985 ( .A(n18674), .B(n18295), .ZN(n18387) );
  XNOR2_X1 U1992 ( .A(n17807), .B(n17913), .ZN(n18390) );
  OAI211_X1 U1993 ( .C1(n17030), .C2(n16662), .A(n4036), .B(n4035), .ZN(n17840) );
  OAI211_X1 U1998 ( .C1(n3601), .C2(n3603), .A(n3600), .B(n3599), .ZN(n18541)
         );
  AND2_X1 U2001 ( .A1(n3260), .A2(n16968), .ZN(n17662) );
  NAND2_X1 U2002 ( .A1(n15882), .A2(n935), .ZN(n934) );
  INV_X1 U2003 ( .A(n15610), .ZN(n1135) );
  AND2_X1 U2004 ( .A1(n2133), .A2(n2134), .ZN(n1253) );
  NAND2_X1 U2008 ( .A1(n16679), .A2(n5521), .ZN(n17807) );
  NAND3_X1 U2009 ( .A1(n1269), .A2(n15635), .A3(n15636), .ZN(n17875) );
  OAI211_X1 U2010 ( .C1(n2429), .C2(n17483), .A(n17480), .B(n2428), .ZN(n18365) );
  OAI21_X1 U2012 ( .B1(n17027), .B2(n3598), .A(n17026), .ZN(n18096) );
  AND2_X1 U2014 ( .A1(n17084), .A2(n16581), .ZN(n575) );
  OR2_X1 U2015 ( .A1(n17465), .A2(n25572), .ZN(n1313) );
  INV_X1 U2016 ( .A(n18310), .ZN(n364) );
  INV_X1 U2017 ( .A(n16615), .ZN(n469) );
  AOI21_X1 U2020 ( .B1(n16964), .B2(n16828), .A(n17441), .ZN(n16430) );
  AND2_X1 U2021 ( .A1(n2508), .A2(n2509), .ZN(n491) );
  NOR2_X1 U2022 ( .A1(n282), .A2(n17175), .ZN(n16523) );
  OAI211_X1 U2023 ( .C1(n16726), .C2(n16974), .A(n17335), .B(n16915), .ZN(
        n16605) );
  OAI21_X1 U2026 ( .B1(n24585), .B2(n16932), .A(n1270), .ZN(n1269) );
  INV_X1 U2027 ( .A(n16746), .ZN(n828) );
  OR2_X1 U2029 ( .A1(n16973), .A2(n17335), .ZN(n17337) );
  OR2_X1 U2030 ( .A1(n17482), .A2(n17481), .ZN(n2428) );
  OR2_X1 U2032 ( .A1(n15884), .A2(n15883), .ZN(n935) );
  OR2_X1 U2033 ( .A1(n17242), .A2(n17240), .ZN(n1283) );
  AND2_X1 U2034 ( .A1(n17193), .A2(n17031), .ZN(n572) );
  INV_X1 U2035 ( .A(n16731), .ZN(n17067) );
  AOI21_X1 U2038 ( .B1(n16929), .B2(n16932), .A(n17059), .ZN(n1270) );
  INV_X1 U2040 ( .A(n17284), .ZN(n17230) );
  OR2_X1 U2041 ( .A1(n17068), .A2(n1139), .ZN(n1138) );
  INV_X1 U2042 ( .A(n17302), .ZN(n470) );
  INV_X1 U2043 ( .A(n16539), .ZN(n365) );
  MUX2_X1 U2044 ( .A(n15163), .B(n15162), .S(n5447), .Z(n17379) );
  INV_X1 U2046 ( .A(n17293), .ZN(n16951) );
  INV_X1 U2048 ( .A(n16871), .ZN(n3602) );
  INV_X1 U2049 ( .A(n17629), .ZN(n366) );
  NOR2_X1 U2050 ( .A1(n17368), .A2(n24471), .ZN(n1546) );
  OR2_X1 U2051 ( .A1(n16795), .A2(n16551), .ZN(n16620) );
  NAND2_X1 U2059 ( .A1(n16245), .A2(n2202), .ZN(n17015) );
  AND3_X1 U2060 ( .A1(n1965), .A2(n16006), .A3(n1964), .ZN(n16846) );
  INV_X1 U2061 ( .A(n17413), .ZN(n16957) );
  INV_X1 U2062 ( .A(n25246), .ZN(n1230) );
  OAI21_X1 U2064 ( .B1(n4675), .B2(n4677), .A(n4676), .ZN(n17175) );
  AND2_X1 U2065 ( .A1(n25465), .A2(n17391), .ZN(n875) );
  INV_X1 U2066 ( .A(n17227), .ZN(n1231) );
  OR2_X1 U2067 ( .A1(n17227), .A2(n17419), .ZN(n1229) );
  INV_X1 U2068 ( .A(n15631), .ZN(n17060) );
  NAND2_X1 U2071 ( .A1(n16033), .A2(n1927), .ZN(n17464) );
  AOI22_X1 U2072 ( .A1(n16228), .A2(n16298), .B1(n16026), .B2(n16025), .ZN(
        n17461) );
  INV_X1 U2074 ( .A(n17141), .ZN(n368) );
  INV_X1 U2075 ( .A(n16261), .ZN(n17166) );
  NOR2_X1 U2080 ( .A1(n17622), .A2(n17624), .ZN(n17472) );
  INV_X1 U2083 ( .A(n17088), .ZN(n371) );
  AND2_X1 U2089 ( .A1(n4646), .A2(n4645), .ZN(n662) );
  OAI21_X1 U2091 ( .B1(n4985), .B2(n4984), .A(n4983), .ZN(n17288) );
  AND2_X1 U2092 ( .A1(n4197), .A2(n5212), .ZN(n1232) );
  NOR2_X1 U2093 ( .A1(n1382), .A2(n15866), .ZN(n4985) );
  NAND4_X1 U2094 ( .A1(n16088), .A2(n16104), .A3(n16087), .A4(n16086), .ZN(
        n16261) );
  AND2_X1 U2095 ( .A1(n15653), .A2(n16416), .ZN(n4984) );
  INV_X1 U2096 ( .A(n17573), .ZN(n373) );
  OAI211_X1 U2098 ( .C1(n16199), .C2(n3143), .A(n16201), .B(n3542), .ZN(n17386) );
  AND2_X1 U2099 ( .A1(n3122), .A2(n2212), .ZN(n16682) );
  INV_X1 U2101 ( .A(n16765), .ZN(n374) );
  INV_X1 U2103 ( .A(n17336), .ZN(n376) );
  OR2_X1 U2104 ( .A1(n15653), .A2(n15868), .ZN(n726) );
  OAI21_X1 U2105 ( .B1(n5414), .B2(n16194), .A(n3288), .ZN(n17622) );
  NOR2_X1 U2106 ( .A1(n1122), .A2(n16342), .ZN(n16347) );
  OR2_X1 U2107 ( .A1(n2251), .A2(n15537), .ZN(n516) );
  OR2_X1 U2108 ( .A1(n2607), .A2(n15564), .ZN(n1097) );
  NOR2_X1 U2109 ( .A1(n16404), .A2(n24062), .ZN(n3143) );
  AND2_X1 U2110 ( .A1(n15677), .A2(n15901), .ZN(n521) );
  NOR2_X1 U2112 ( .A1(n16392), .A2(n24537), .ZN(n15850) );
  BUF_X1 U2114 ( .A(n15545), .Z(n16475) );
  XNOR2_X1 U2115 ( .A(n2000), .B(n14597), .ZN(n16042) );
  INV_X1 U2116 ( .A(n15557), .ZN(n16010) );
  XNOR2_X1 U2117 ( .A(n14527), .B(n14526), .ZN(n16389) );
  INV_X1 U2118 ( .A(n24981), .ZN(n377) );
  XNOR2_X1 U2119 ( .A(n15140), .B(n1105), .ZN(n1103) );
  CLKBUF_X1 U2121 ( .A(n15640), .Z(n15907) );
  INV_X1 U2122 ( .A(n16109), .ZN(n379) );
  INV_X1 U2124 ( .A(n16423), .ZN(n707) );
  XNOR2_X1 U2125 ( .A(n13476), .B(n13475), .ZN(n16333) );
  XNOR2_X1 U2126 ( .A(n13939), .B(n13938), .ZN(n15970) );
  XNOR2_X1 U2129 ( .A(n15116), .B(n15115), .ZN(n16360) );
  XNOR2_X1 U2130 ( .A(n15469), .B(n15468), .ZN(n16473) );
  INV_X1 U2131 ( .A(n16067), .ZN(n380) );
  INV_X1 U2132 ( .A(n15646), .ZN(n16401) );
  XNOR2_X1 U2133 ( .A(n5192), .B(n14742), .ZN(n15583) );
  OR2_X1 U2138 ( .A1(n14926), .A2(n16029), .ZN(n2651) );
  XNOR2_X1 U2145 ( .A(n4399), .B(n15189), .ZN(n15198) );
  INV_X1 U2147 ( .A(n16176), .ZN(n15655) );
  INV_X1 U2148 ( .A(n16125), .ZN(n381) );
  CLKBUF_X1 U2149 ( .A(n13940), .Z(n15971) );
  XNOR2_X1 U2150 ( .A(n15014), .B(n15013), .ZN(n15560) );
  XNOR2_X1 U2153 ( .A(n14706), .B(n14707), .ZN(n16107) );
  INV_X1 U2154 ( .A(n15549), .ZN(n382) );
  INV_X1 U2156 ( .A(n15715), .ZN(n383) );
  XNOR2_X1 U2157 ( .A(n15086), .B(n15085), .ZN(n16290) );
  XNOR2_X1 U2158 ( .A(n15137), .B(n15136), .ZN(n16001) );
  XNOR2_X1 U2160 ( .A(n12909), .B(n14840), .ZN(n16349) );
  INV_X1 U2165 ( .A(n16449), .ZN(n385) );
  INV_X1 U2166 ( .A(n16381), .ZN(n386) );
  XNOR2_X1 U2167 ( .A(n14380), .B(n14379), .ZN(n16121) );
  INV_X1 U2168 ( .A(n15564), .ZN(n387) );
  INV_X1 U2169 ( .A(n16332), .ZN(n388) );
  XNOR2_X1 U2171 ( .A(n14657), .B(n14656), .ZN(n16129) );
  XNOR2_X1 U2172 ( .A(n14890), .B(n14894), .ZN(n796) );
  CLKBUF_X1 U2174 ( .A(n16219), .Z(n16458) );
  XNOR2_X1 U2177 ( .A(n14904), .B(n540), .ZN(n14905) );
  INV_X1 U2178 ( .A(n16219), .ZN(n389) );
  XNOR2_X1 U2179 ( .A(n12679), .B(n14845), .ZN(n15070) );
  XNOR2_X1 U2180 ( .A(n4859), .B(n1907), .ZN(n15405) );
  INV_X1 U2181 ( .A(n14788), .ZN(n1111) );
  INV_X1 U2182 ( .A(n3787), .ZN(n15188) );
  XNOR2_X1 U2183 ( .A(n15446), .B(n15109), .ZN(n540) );
  INV_X1 U2184 ( .A(n15177), .ZN(n5215) );
  XNOR2_X1 U2185 ( .A(n15293), .B(n1104), .ZN(n1102) );
  XNOR2_X1 U2190 ( .A(n15138), .B(n15483), .ZN(n1105) );
  NAND2_X1 U2191 ( .A1(n4558), .A2(n13690), .ZN(n15003) );
  NAND2_X1 U2194 ( .A1(n4330), .A2(n13483), .ZN(n15190) );
  XNOR2_X1 U2195 ( .A(n15386), .B(n1833), .ZN(n1104) );
  NAND2_X1 U2203 ( .A1(n2382), .A2(n2381), .ZN(n15463) );
  NAND4_X1 U2205 ( .A1(n14259), .A2(n14260), .A3(n14258), .A4(n14257), .ZN(
        n14958) );
  INV_X1 U2206 ( .A(n14043), .ZN(n985) );
  NAND3_X1 U2207 ( .A1(n2911), .A2(n13934), .A3(n2910), .ZN(n14997) );
  OR2_X1 U2209 ( .A1(n13667), .A2(n5753), .ZN(n13679) );
  NAND3_X1 U2210 ( .A1(n5332), .A2(n13567), .A3(n3983), .ZN(n15244) );
  NOR2_X1 U2214 ( .A1(n13895), .A2(n14130), .ZN(n620) );
  OAI21_X1 U2215 ( .B1(n13655), .B2(n13379), .A(n13989), .ZN(n13381) );
  AND2_X1 U2216 ( .A1(n14206), .A2(n14205), .ZN(n13551) );
  NOR2_X1 U2217 ( .A1(n14327), .A2(n13864), .ZN(n5246) );
  NOR2_X1 U2218 ( .A1(n13596), .A2(n13969), .ZN(n5520) );
  OR2_X1 U2219 ( .A1(n14328), .A2(n14041), .ZN(n12803) );
  OR2_X1 U2221 ( .A1(n10396), .A2(n508), .ZN(n967) );
  OR2_X1 U2223 ( .A1(n13995), .A2(n14235), .ZN(n795) );
  INV_X1 U2224 ( .A(n14076), .ZN(n13852) );
  OR2_X1 U2225 ( .A1(n13921), .A2(n13922), .ZN(n760) );
  AND2_X1 U2226 ( .A1(n24949), .A2(n13796), .ZN(n14180) );
  INV_X1 U2228 ( .A(n3959), .ZN(n13534) );
  OR2_X1 U2229 ( .A1(n14327), .A2(n14325), .ZN(n13863) );
  NOR2_X1 U2230 ( .A1(n14034), .A2(n14149), .ZN(n14151) );
  OR2_X1 U2231 ( .A1(n13851), .A2(n14078), .ZN(n13631) );
  OR2_X1 U2232 ( .A1(n13609), .A2(n14085), .ZN(n1060) );
  INV_X1 U2234 ( .A(n4116), .ZN(n14241) );
  NAND2_X1 U2235 ( .A1(n2317), .A2(n2316), .ZN(n14034) );
  INV_X1 U2236 ( .A(n13533), .ZN(n14088) );
  OR2_X1 U2237 ( .A1(n14022), .A2(n4510), .ZN(n13607) );
  INV_X1 U2238 ( .A(n13951), .ZN(n391) );
  NAND2_X1 U2239 ( .A1(n1017), .A2(n12890), .ZN(n14149) );
  OR2_X1 U2240 ( .A1(n14089), .A2(n13533), .ZN(n3959) );
  OAI21_X1 U2241 ( .B1(n12778), .B2(n12777), .A(n12776), .ZN(n13796) );
  AND2_X1 U2243 ( .A1(n612), .A2(n13502), .ZN(n13506) );
  AND2_X1 U2244 ( .A1(n13656), .A2(n13918), .ZN(n755) );
  INV_X1 U2245 ( .A(n13818), .ZN(n392) );
  NOR2_X1 U2248 ( .A1(n623), .A2(n12913), .ZN(n622) );
  NAND2_X1 U2249 ( .A1(n1081), .A2(n5022), .ZN(n4510) );
  AND4_X1 U2251 ( .A1(n13334), .A2(n13333), .A3(n13332), .A4(n13331), .ZN(
        n13682) );
  OAI211_X1 U2252 ( .C1(n1632), .C2(n13134), .A(n1631), .B(n1630), .ZN(n13552)
         );
  INV_X1 U2254 ( .A(n14049), .ZN(n13518) );
  INV_X1 U2255 ( .A(n14035), .ZN(n1028) );
  OR3_X1 U2256 ( .A1(n12119), .A2(n12118), .A3(n12117), .ZN(n1553) );
  AND2_X1 U2259 ( .A1(n5470), .A2(n4923), .ZN(n1127) );
  INV_X1 U2260 ( .A(n13503), .ZN(n612) );
  AND3_X1 U2261 ( .A1(n5310), .A2(n5309), .A3(n5314), .ZN(n14143) );
  INV_X1 U2262 ( .A(n14324), .ZN(n14041) );
  OR2_X1 U2263 ( .A1(n13128), .A2(n13127), .ZN(n14211) );
  OAI211_X2 U2266 ( .C1(n24487), .C2(n12558), .A(n12557), .B(n12556), .ZN(
        n14078) );
  OAI21_X1 U2267 ( .B1(n13021), .B2(n13020), .A(n13019), .ZN(n14225) );
  AND2_X1 U2268 ( .A1(n12828), .A2(n1508), .ZN(n13502) );
  INV_X1 U2270 ( .A(n13907), .ZN(n394) );
  AND3_X1 U2271 ( .A1(n4596), .A2(n4595), .A3(n25053), .ZN(n13681) );
  INV_X1 U2272 ( .A(n24999), .ZN(n395) );
  INV_X1 U2273 ( .A(n13419), .ZN(n1314) );
  OR2_X1 U2275 ( .A1(n12463), .A2(n12464), .ZN(n493) );
  AND2_X1 U2276 ( .A1(n1082), .A2(n12504), .ZN(n13537) );
  NAND3_X1 U2278 ( .A1(n12456), .A2(n12458), .A3(n12457), .ZN(n14049) );
  INV_X1 U2279 ( .A(n14269), .ZN(n397) );
  OAI21_X1 U2280 ( .B1(n3975), .B2(n3974), .A(n3972), .ZN(n14048) );
  AND2_X1 U2281 ( .A1(n12661), .A2(n13115), .ZN(n1267) );
  OR2_X1 U2282 ( .A1(n4587), .A2(n12995), .ZN(n1018) );
  OAI21_X1 U2283 ( .B1(n12937), .B2(n4493), .A(n1445), .ZN(n4491) );
  OR2_X1 U2285 ( .A1(n13220), .A2(n24513), .ZN(n780) );
  NOR2_X1 U2286 ( .A1(n12690), .A2(n12910), .ZN(n12598) );
  INV_X1 U2287 ( .A(n10200), .ZN(n499) );
  OR2_X1 U2288 ( .A1(n12179), .A2(n13093), .ZN(n597) );
  OR2_X1 U2289 ( .A1(n11328), .A2(n12993), .ZN(n1020) );
  BUF_X1 U2290 ( .A(n12868), .Z(n13119) );
  NOR2_X1 U2292 ( .A1(n12834), .A2(n13274), .ZN(n1201) );
  AND2_X1 U2294 ( .A1(n24346), .A2(n13272), .ZN(n4446) );
  INV_X1 U2295 ( .A(n12695), .ZN(n1200) );
  OR2_X1 U2296 ( .A1(n12792), .A2(n12995), .ZN(n12991) );
  AND2_X1 U2298 ( .A1(n12859), .A2(n12860), .ZN(n12863) );
  AOI21_X1 U2299 ( .B1(n1069), .B2(n12178), .A(n13092), .ZN(n4333) );
  OR2_X1 U2300 ( .A1(n12433), .A2(n13144), .ZN(n1915) );
  OR2_X1 U2301 ( .A1(n12738), .A2(n13162), .ZN(n3710) );
  AND2_X1 U2302 ( .A1(n12648), .A2(n12178), .ZN(n10200) );
  XNOR2_X1 U2306 ( .A(n12026), .B(n12027), .ZN(n13325) );
  INV_X1 U2307 ( .A(n12859), .ZN(n398) );
  CLKBUF_X1 U2309 ( .A(n12519), .Z(n12523) );
  BUF_X1 U2310 ( .A(n12520), .Z(n13040) );
  INV_X1 U2311 ( .A(n12454), .ZN(n13063) );
  XNOR2_X1 U2314 ( .A(n12361), .B(n12360), .ZN(n12861) );
  INV_X1 U2317 ( .A(n1324), .ZN(n10360) );
  INV_X1 U2318 ( .A(n12576), .ZN(n399) );
  XNOR2_X1 U2320 ( .A(n9971), .B(n9970), .ZN(n12178) );
  INV_X1 U2321 ( .A(n13335), .ZN(n400) );
  AND2_X1 U2322 ( .A1(n13027), .A2(n13028), .ZN(n563) );
  INV_X1 U2324 ( .A(n13050), .ZN(n401) );
  INV_X1 U2326 ( .A(n12725), .ZN(n403) );
  INV_X1 U2328 ( .A(n12600), .ZN(n404) );
  XNOR2_X1 U2329 ( .A(n12238), .B(n12237), .ZN(n13110) );
  XNOR2_X1 U2333 ( .A(n11364), .B(n11365), .ZN(n13213) );
  XNOR2_X1 U2335 ( .A(n12071), .B(n12070), .ZN(n13329) );
  INV_X1 U2336 ( .A(n13301), .ZN(n405) );
  XNOR2_X1 U2337 ( .A(n10708), .B(n10709), .ZN(n13130) );
  INV_X1 U2339 ( .A(n13124), .ZN(n406) );
  XNOR2_X1 U2340 ( .A(n11379), .B(n11378), .ZN(n12784) );
  XNOR2_X1 U2342 ( .A(n11443), .B(n11444), .ZN(n12796) );
  INV_X1 U2343 ( .A(n13267), .ZN(n407) );
  INV_X1 U2345 ( .A(n12795), .ZN(n408) );
  INV_X1 U2347 ( .A(n13056), .ZN(n409) );
  XNOR2_X1 U2352 ( .A(n4485), .B(n11744), .ZN(n13227) );
  XNOR2_X1 U2353 ( .A(n11810), .B(n11811), .ZN(n13235) );
  XNOR2_X1 U2354 ( .A(n12389), .B(n11247), .ZN(n11827) );
  INV_X1 U2355 ( .A(n11796), .ZN(n3648) );
  XNOR2_X1 U2356 ( .A(n9407), .B(n9406), .ZN(n9408) );
  XNOR2_X1 U2357 ( .A(n11414), .B(n12365), .ZN(n11356) );
  XNOR2_X1 U2358 ( .A(n11743), .B(n11745), .ZN(n4485) );
  XNOR2_X1 U2361 ( .A(n11464), .B(n2241), .ZN(n11315) );
  INV_X1 U2362 ( .A(n11253), .ZN(n11915) );
  XNOR2_X1 U2363 ( .A(n1177), .B(n11983), .ZN(n12088) );
  XNOR2_X1 U2366 ( .A(n4670), .B(n4668), .ZN(n11180) );
  MUX2_X1 U2370 ( .A(n11219), .B(n11218), .S(n233), .Z(n11568) );
  INV_X1 U2372 ( .A(n11845), .ZN(n12283) );
  AND3_X1 U2374 ( .A1(n10503), .A2(n3511), .A3(n3510), .ZN(n4670) );
  AOI22_X1 U2375 ( .A1(n10319), .A2(n10590), .B1(n10583), .B2(n10318), .ZN(
        n12248) );
  NAND3_X1 U2378 ( .A1(n10294), .A2(n10295), .A3(n202), .ZN(n11698) );
  AND3_X1 U2379 ( .A1(n9571), .A2(n9572), .A3(n4040), .ZN(n12402) );
  NAND4_X1 U2380 ( .A1(n1226), .A2(n1223), .A3(n1227), .A4(n1225), .ZN(n11253)
         );
  OAI211_X1 U2381 ( .C1(n10743), .C2(n10858), .A(n10742), .B(n10741), .ZN(
        n12066) );
  AND3_X1 U2382 ( .A1(n527), .A2(n526), .A3(n11050), .ZN(n12082) );
  NAND4_X1 U2383 ( .A1(n11174), .A2(n3384), .A3(n10383), .A4(n3385), .ZN(
        n11959) );
  AND2_X1 U2384 ( .A1(n531), .A2(n532), .ZN(n530) );
  OR2_X1 U2389 ( .A1(n11203), .A2(n11204), .ZN(n3011) );
  INV_X1 U2390 ( .A(n3443), .ZN(n10202) );
  NAND3_X1 U2391 ( .A1(n10928), .A2(n10929), .A3(n4691), .ZN(n12315) );
  AND2_X1 U2392 ( .A1(n10804), .A2(n10798), .ZN(n10806) );
  OAI21_X1 U2393 ( .B1(n10642), .B2(n11046), .A(n529), .ZN(n5671) );
  NOR2_X1 U2395 ( .A1(n10967), .A2(n10971), .ZN(n10818) );
  MUX2_X1 U2396 ( .A(n9210), .B(n9209), .S(n10587), .Z(n9216) );
  OR2_X1 U2397 ( .A1(n10805), .A2(n10799), .ZN(n735) );
  OR2_X1 U2398 ( .A1(n11082), .A2(n5559), .ZN(n1264) );
  OR2_X1 U2399 ( .A1(n11205), .A2(n11338), .ZN(n10821) );
  OR2_X1 U2400 ( .A1(n10527), .A2(n11529), .ZN(n525) );
  OR2_X1 U2402 ( .A1(n11091), .A2(n1057), .ZN(n1056) );
  INV_X1 U2403 ( .A(n10491), .ZN(n10233) );
  INV_X1 U2405 ( .A(n11212), .ZN(n3868) );
  NOR2_X1 U2406 ( .A1(n11099), .A2(n939), .ZN(n10782) );
  NOR2_X1 U2408 ( .A1(n10617), .A2(n10411), .ZN(n559) );
  INV_X1 U2409 ( .A(n11024), .ZN(n895) );
  INV_X1 U2410 ( .A(n11302), .ZN(n11300) );
  INV_X1 U2412 ( .A(n10887), .ZN(n10301) );
  INV_X1 U2413 ( .A(n939), .ZN(n10911) );
  CLKBUF_X1 U2414 ( .A(n11172), .Z(n1338) );
  INV_X1 U2415 ( .A(n232), .ZN(n10812) );
  INV_X1 U2416 ( .A(n10583), .ZN(n9443) );
  INV_X1 U2418 ( .A(n10798), .ZN(n10805) );
  INV_X1 U2419 ( .A(n4531), .ZN(n528) );
  INV_X1 U2420 ( .A(n11059), .ZN(n410) );
  NAND2_X1 U2424 ( .A1(n5535), .A2(n5534), .ZN(n10762) );
  INV_X1 U2426 ( .A(n9432), .ZN(n412) );
  INV_X1 U2427 ( .A(n10523), .ZN(n11024) );
  INV_X1 U2428 ( .A(n10277), .ZN(n413) );
  OR2_X1 U2430 ( .A1(n1181), .A2(n1963), .ZN(n10798) );
  INV_X1 U2431 ( .A(n11342), .ZN(n414) );
  OR2_X1 U2432 ( .A1(n9618), .A2(n9617), .ZN(n660) );
  INV_X1 U2434 ( .A(n11499), .ZN(n1218) );
  AND2_X1 U2435 ( .A1(n10778), .A2(n9502), .ZN(n1552) );
  INV_X1 U2436 ( .A(n10886), .ZN(n10541) );
  NAND2_X1 U2438 ( .A1(n9502), .A2(n10778), .ZN(n11099) );
  OAI21_X1 U2439 ( .B1(n9840), .B2(n10099), .A(n9839), .ZN(n10703) );
  INV_X1 U2440 ( .A(n11032), .ZN(n415) );
  AND2_X1 U2441 ( .A1(n9250), .A2(n1816), .ZN(n10855) );
  OR2_X1 U2444 ( .A1(n9201), .A2(n627), .ZN(n9582) );
  INV_X1 U2446 ( .A(n11039), .ZN(n416) );
  INV_X1 U2448 ( .A(n11163), .ZN(n417) );
  INV_X1 U2449 ( .A(n10889), .ZN(n418) );
  OAI211_X1 U2453 ( .C1(n3722), .C2(n5609), .A(n5608), .B(n3721), .ZN(n11121)
         );
  OR2_X1 U2454 ( .A1(n9128), .A2(n9129), .ZN(n11036) );
  OAI21_X1 U2455 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n10614) );
  AOI22_X1 U2458 ( .A1(n2140), .A2(n1796), .B1(n9501), .B2(n246), .ZN(n10778)
         );
  INV_X1 U2462 ( .A(n11298), .ZN(n419) );
  INV_X1 U2464 ( .A(n11130), .ZN(n420) );
  OAI22_X1 U2466 ( .A1(n5523), .A2(n24054), .B1(n9945), .B2(n1165), .ZN(n1181)
         );
  OAI21_X1 U2467 ( .B1(n10122), .B2(n9841), .A(n24087), .ZN(n2256) );
  OR2_X1 U2468 ( .A1(n9225), .A2(n9740), .ZN(n1168) );
  NOR2_X1 U2469 ( .A1(n2294), .A2(n1021), .ZN(n9693) );
  INV_X1 U2470 ( .A(n3305), .ZN(n699) );
  INV_X1 U2471 ( .A(n24085), .ZN(n2257) );
  OR2_X1 U2474 ( .A1(n9808), .A2(n9807), .ZN(n1318) );
  INV_X1 U2475 ( .A(n9417), .ZN(n9758) );
  NOR2_X1 U2477 ( .A1(n9872), .A2(n1021), .ZN(n1519) );
  AND2_X1 U2479 ( .A1(n9886), .A2(n9565), .ZN(n956) );
  AOI21_X1 U2480 ( .B1(n3292), .B2(n9281), .A(n9468), .ZN(n665) );
  AND2_X1 U2482 ( .A1(n8521), .A2(n9798), .ZN(n9314) );
  BUF_X1 U2483 ( .A(n8483), .Z(n9999) );
  OR2_X1 U2484 ( .A1(n24446), .A2(n4096), .ZN(n4097) );
  INV_X1 U2485 ( .A(n10108), .ZN(n9524) );
  INV_X1 U2487 ( .A(n9237), .ZN(n9697) );
  INV_X1 U2488 ( .A(n4254), .ZN(n1275) );
  OR2_X1 U2489 ( .A1(n9295), .A2(n9781), .ZN(n5025) );
  AND2_X1 U2490 ( .A1(n24535), .A2(n9990), .ZN(n9425) );
  NOR2_X1 U2491 ( .A1(n25005), .A2(n9418), .ZN(n9615) );
  INV_X1 U2492 ( .A(n9027), .ZN(n1021) );
  CLKBUF_X1 U2493 ( .A(n9297), .Z(n9780) );
  INV_X1 U2495 ( .A(n3292), .ZN(n1185) );
  BUF_X1 U2496 ( .A(n9398), .Z(n10136) );
  INV_X1 U2498 ( .A(n10251), .ZN(n10250) );
  NOR2_X1 U2499 ( .A1(n24087), .A2(n9843), .ZN(n2413) );
  OR2_X1 U2500 ( .A1(n10058), .A2(n4096), .ZN(n794) );
  CLKBUF_X1 U2501 ( .A(n9419), .Z(n9754) );
  INV_X1 U2505 ( .A(n8359), .ZN(n421) );
  INV_X1 U2507 ( .A(n24534), .ZN(n422) );
  XNOR2_X1 U2509 ( .A(n7454), .B(n7453), .ZN(n9962) );
  INV_X1 U2511 ( .A(n24505), .ZN(n424) );
  INV_X1 U2514 ( .A(n9779), .ZN(n425) );
  XNOR2_X1 U2515 ( .A(n8785), .B(n8784), .ZN(n9418) );
  INV_X1 U2516 ( .A(n9491), .ZN(n426) );
  INV_X1 U2517 ( .A(n9945), .ZN(n9942) );
  BUF_X1 U2518 ( .A(n8523), .Z(n9530) );
  BUF_X1 U2519 ( .A(n10071), .Z(n1330) );
  BUF_X1 U2520 ( .A(n9218), .Z(n10065) );
  XNOR2_X1 U2521 ( .A(n7042), .B(n7041), .ZN(n9918) );
  INV_X1 U2522 ( .A(n10109), .ZN(n4254) );
  XNOR2_X1 U2524 ( .A(n8816), .B(n8817), .ZN(n10018) );
  INV_X1 U2526 ( .A(n10071), .ZN(n427) );
  XNOR2_X1 U2528 ( .A(n8464), .B(n8463), .ZN(n9786) );
  XNOR2_X1 U2531 ( .A(n8944), .B(n8943), .ZN(n10046) );
  XNOR2_X1 U2532 ( .A(n8767), .B(n8768), .ZN(n9752) );
  XNOR2_X1 U2534 ( .A(n7497), .B(n7496), .ZN(n9964) );
  INV_X1 U2536 ( .A(n9837), .ZN(n428) );
  XNOR2_X1 U2537 ( .A(n8626), .B(n8625), .ZN(n10109) );
  INV_X1 U2540 ( .A(n9127), .ZN(n429) );
  XNOR2_X1 U2541 ( .A(n8559), .B(n2274), .ZN(n2276) );
  INV_X1 U2542 ( .A(n8951), .ZN(n5184) );
  XNOR2_X1 U2543 ( .A(n5344), .B(n8798), .ZN(n8198) );
  XNOR2_X1 U2545 ( .A(n8613), .B(n8280), .ZN(n9089) );
  XNOR2_X1 U2546 ( .A(n8980), .B(n1110), .ZN(n8778) );
  XNOR2_X1 U2548 ( .A(n8787), .B(n8450), .ZN(n9012) );
  OAI21_X1 U2557 ( .B1(n5116), .B2(n7952), .A(n2490), .ZN(n9159) );
  OAI21_X1 U2560 ( .B1(n3267), .B2(n7843), .A(n3265), .ZN(n8615) );
  NAND3_X1 U2561 ( .A1(n7745), .A2(n7746), .A3(n1972), .ZN(n9002) );
  OR2_X1 U2562 ( .A1(n4975), .A2(n7859), .ZN(n8789) );
  NAND2_X1 U2567 ( .A1(n7484), .A2(n4001), .ZN(n8795) );
  NOR2_X1 U2569 ( .A1(n7807), .A2(n7806), .ZN(n8450) );
  NAND3_X1 U2571 ( .A1(n7178), .A2(n7177), .A3(n7176), .ZN(n8917) );
  MUX2_X1 U2572 ( .A(n7446), .B(n7447), .S(n5607), .Z(n8492) );
  NAND3_X1 U2574 ( .A1(n2263), .A2(n7509), .A3(n2261), .ZN(n8769) );
  AND2_X1 U2575 ( .A1(n7158), .A2(n5345), .ZN(n7161) );
  NAND3_X1 U2577 ( .A1(n1848), .A2(n7137), .A3(n7138), .ZN(n8647) );
  NAND2_X1 U2579 ( .A1(n7729), .A2(n7728), .ZN(n8914) );
  AOI22_X1 U2581 ( .A1(n8024), .A2(n3258), .B1(n3259), .B2(n7532), .ZN(n3257)
         );
  OR2_X1 U2583 ( .A1(n3236), .A2(n2640), .ZN(n3235) );
  AND2_X1 U2584 ( .A1(n4145), .A2(n7953), .ZN(n842) );
  AND2_X1 U2585 ( .A1(n7282), .A2(n7281), .ZN(n533) );
  OAI21_X1 U2586 ( .B1(n806), .B2(n1345), .A(n2223), .ZN(n7487) );
  OAI21_X1 U2588 ( .B1(n3500), .B2(n7580), .A(n3498), .ZN(n8981) );
  AND2_X1 U2589 ( .A1(n7533), .A2(n7747), .ZN(n3258) );
  INV_X1 U2591 ( .A(n7349), .ZN(n1279) );
  OR2_X1 U2592 ( .A1(n7651), .A2(n7650), .ZN(n989) );
  OAI21_X1 U2593 ( .B1(n7322), .B2(n7890), .A(n311), .ZN(n1124) );
  INV_X1 U2594 ( .A(n941), .ZN(n7622) );
  OR2_X1 U2596 ( .A1(n2522), .A2(n8003), .ZN(n736) );
  AND2_X1 U2598 ( .A1(n7537), .A2(n7748), .ZN(n8011) );
  INV_X1 U2599 ( .A(n7444), .ZN(n7163) );
  OR2_X1 U2600 ( .A1(n7593), .A2(n7592), .ZN(n1190) );
  INV_X1 U2601 ( .A(n7754), .ZN(n7542) );
  OR2_X1 U2602 ( .A1(n7760), .A2(n7646), .ZN(n6194) );
  INV_X1 U2603 ( .A(n7683), .ZN(n7235) );
  INV_X1 U2605 ( .A(n512), .ZN(n7634) );
  INV_X1 U2607 ( .A(n1162), .ZN(n7676) );
  INV_X1 U2608 ( .A(n7074), .ZN(n7506) );
  OR3_X1 U2609 ( .A1(n7350), .A2(n5468), .A3(n7346), .ZN(n7253) );
  INV_X1 U2610 ( .A(n7078), .ZN(n3275) );
  NAND2_X1 U2611 ( .A1(n6581), .A2(n5604), .ZN(n7924) );
  INV_X1 U2612 ( .A(n7914), .ZN(n430) );
  CLKBUF_X1 U2614 ( .A(n6806), .Z(n7667) );
  CLKBUF_X1 U2615 ( .A(n7246), .Z(n7855) );
  OAI21_X1 U2616 ( .B1(n6443), .B2(n6296), .A(n6213), .ZN(n2640) );
  OR2_X1 U2617 ( .A1(n270), .A2(n7962), .ZN(n584) );
  INV_X1 U2618 ( .A(n7533), .ZN(n1975) );
  INV_X1 U2619 ( .A(n2624), .ZN(n7748) );
  AND2_X1 U2620 ( .A1(n2401), .A2(n2400), .ZN(n2402) );
  NOR2_X1 U2621 ( .A1(n1162), .A2(n1085), .ZN(n1084) );
  NAND2_X1 U2622 ( .A1(n3608), .A2(n6313), .ZN(n7861) );
  NAND2_X1 U2624 ( .A1(n764), .A2(n1174), .ZN(n7683) );
  NAND2_X1 U2626 ( .A1(n1433), .A2(n2899), .ZN(n7732) );
  INV_X1 U2627 ( .A(n7423), .ZN(n431) );
  NAND2_X1 U2628 ( .A1(n943), .A2(n944), .ZN(n942) );
  OAI211_X1 U2633 ( .C1(n5729), .C2(n6049), .A(n504), .B(n502), .ZN(n7108) );
  AND2_X1 U2636 ( .A1(n5890), .A2(n5889), .ZN(n7896) );
  INV_X1 U2637 ( .A(n7217), .ZN(n433) );
  INV_X1 U2638 ( .A(n7983), .ZN(n7827) );
  INV_X1 U2640 ( .A(n7224), .ZN(n434) );
  OAI21_X1 U2641 ( .B1(n5142), .B2(n5143), .A(n6273), .ZN(n7803) );
  AND2_X1 U2646 ( .A1(n5912), .A2(n5911), .ZN(n7347) );
  INV_X1 U2647 ( .A(n7915), .ZN(n435) );
  INV_X1 U2648 ( .A(n7664), .ZN(n436) );
  NAND2_X1 U2650 ( .A1(n6103), .A2(n6102), .ZN(n7768) );
  NAND2_X1 U2651 ( .A1(n1695), .A2(n568), .ZN(n1162) );
  INV_X1 U2653 ( .A(n6323), .ZN(n944) );
  OAI211_X1 U2654 ( .C1(n6412), .C2(n6051), .A(n6411), .B(n6410), .ZN(n7853)
         );
  AOI21_X1 U2658 ( .B1(n5088), .B2(n7024), .A(n2738), .ZN(n2737) );
  INV_X1 U2661 ( .A(n7962), .ZN(n437) );
  OAI21_X1 U2663 ( .B1(n709), .B2(n6553), .A(n708), .ZN(n1750) );
  AOI22_X1 U2664 ( .A1(n7005), .A2(n6835), .B1(n7004), .B2(n6836), .ZN(n467)
         );
  OR2_X1 U2665 ( .A1(n6177), .A2(n6178), .ZN(n7646) );
  INV_X1 U2667 ( .A(n1379), .ZN(n1085) );
  OR2_X1 U2668 ( .A1(n6463), .A2(n6464), .ZN(n773) );
  AND2_X1 U2669 ( .A1(n6274), .A2(n6324), .ZN(n6522) );
  OAI21_X1 U2670 ( .B1(n6906), .B2(n6905), .A(n6373), .ZN(n6475) );
  AND2_X1 U2671 ( .A1(n6519), .A2(n6275), .ZN(n6524) );
  AND2_X1 U2672 ( .A1(n6957), .A2(n6705), .ZN(n709) );
  AND2_X1 U2673 ( .A1(n6641), .A2(n6642), .ZN(n5635) );
  NAND2_X1 U2674 ( .A1(n6328), .A2(n5451), .ZN(n1079) );
  OAI21_X1 U2676 ( .B1(n669), .B2(n6674), .A(n668), .ZN(n6676) );
  INV_X1 U2677 ( .A(n6570), .ZN(n4754) );
  OR2_X1 U2678 ( .A1(n6588), .A2(n625), .ZN(n6226) );
  CLKBUF_X1 U2682 ( .A(n6187), .Z(n6347) );
  INV_X1 U2684 ( .A(n6999), .ZN(n947) );
  OR2_X1 U2687 ( .A1(n7035), .A2(n625), .ZN(n6591) );
  INV_X1 U2688 ( .A(n625), .ZN(n7033) );
  INV_X1 U2689 ( .A(n4324), .ZN(n708) );
  BUF_X1 U2690 ( .A(n6381), .Z(n7025) );
  INV_X1 U2691 ( .A(n6453), .ZN(n1106) );
  INV_X1 U2693 ( .A(n6683), .ZN(n6939) );
  INV_X1 U2696 ( .A(n6174), .ZN(n438) );
  INV_X1 U2697 ( .A(n6367), .ZN(n439) );
  BUF_X1 U2700 ( .A(n5887), .Z(n6679) );
  INV_X1 U2702 ( .A(n6324), .ZN(n440) );
  NOR2_X1 U2703 ( .A1(n6757), .A2(n6578), .ZN(n669) );
  INV_X1 U2705 ( .A(n1804), .ZN(n931) );
  INV_X1 U2706 ( .A(n5824), .ZN(n6372) );
  INV_X1 U2707 ( .A(n6496), .ZN(n441) );
  INV_X1 U2709 ( .A(n6578), .ZN(n5805) );
  INV_X1 U2710 ( .A(n23868), .ZN(n4189) );
  INV_X1 U2711 ( .A(n6381), .ZN(n442) );
  AOI21_X1 U2712 ( .B1(n6498), .B2(n6034), .A(n6434), .ZN(n2218) );
  AND3_X1 U2714 ( .A1(n6777), .A2(n6198), .A3(n6775), .ZN(n1295) );
  CLKBUF_X1 U2715 ( .A(Key[102]), .Z(n677) );
  CLKBUF_X1 U2717 ( .A(Key[140]), .Z(n3190) );
  CLKBUF_X1 U2721 ( .A(Key[64]), .Z(n2970) );
  CLKBUF_X1 U2722 ( .A(Key[53]), .Z(n2215) );
  INV_X1 U2723 ( .A(n2744), .ZN(n444) );
  CLKBUF_X1 U2725 ( .A(Key[30]), .Z(n3133) );
  XNOR2_X1 U2726 ( .A(Key[44]), .B(Plaintext[44]), .ZN(n6955) );
  INV_X1 U2727 ( .A(n1952), .ZN(n445) );
  CLKBUF_X1 U2728 ( .A(Key[57]), .Z(n887) );
  CLKBUF_X1 U2729 ( .A(Key[167]), .Z(n2743) );
  CLKBUF_X1 U2730 ( .A(Key[151]), .Z(n1874) );
  CLKBUF_X1 U2731 ( .A(Key[61]), .Z(n21046) );
  CLKBUF_X1 U2732 ( .A(Key[91]), .Z(n1935) );
  CLKBUF_X1 U2733 ( .A(Key[164]), .Z(n2137) );
  CLKBUF_X1 U2734 ( .A(Key[90]), .Z(n2034) );
  INV_X1 U2737 ( .A(n768), .ZN(n447) );
  INV_X1 U2740 ( .A(n7008), .ZN(n448) );
  CLKBUF_X1 U2741 ( .A(Key[187]), .Z(n888) );
  XNOR2_X1 U2743 ( .A(Plaintext[145]), .B(Key[145]), .ZN(n5824) );
  INV_X1 U2744 ( .A(n2834), .ZN(n449) );
  INV_X1 U2746 ( .A(n1833), .ZN(n450) );
  XNOR2_X1 U2749 ( .A(Key[187]), .B(Plaintext[187]), .ZN(n6195) );
  CLKBUF_X1 U2750 ( .A(Key[132]), .Z(n3155) );
  CLKBUF_X1 U2751 ( .A(Key[54]), .Z(n2795) );
  INV_X1 U2753 ( .A(n22886), .ZN(n451) );
  INV_X1 U2754 ( .A(n1865), .ZN(n452) );
  CLKBUF_X1 U2756 ( .A(Key[179]), .Z(n21964) );
  INV_X1 U2757 ( .A(n6050), .ZN(n453) );
  CLKBUF_X1 U2758 ( .A(Key[122]), .Z(n23476) );
  CLKBUF_X1 U2759 ( .A(Key[186]), .Z(n1726) );
  XNOR2_X1 U2760 ( .A(Key[85]), .B(Plaintext[85]), .ZN(n6243) );
  CLKBUF_X1 U2761 ( .A(Key[134]), .Z(n729) );
  CLKBUF_X1 U2762 ( .A(Key[8]), .Z(n3152) );
  INV_X1 U2763 ( .A(n7029), .ZN(n454) );
  CLKBUF_X1 U2764 ( .A(Key[26]), .Z(n3073) );
  INV_X1 U2765 ( .A(n765), .ZN(n455) );
  CLKBUF_X1 U2766 ( .A(Key[13]), .Z(n3125) );
  NAND2_X1 U2767 ( .A1(n19323), .A2(n456), .ZN(n19936) );
  NAND2_X1 U2768 ( .A1(n458), .A2(n457), .ZN(n456) );
  OAI211_X2 U2769 ( .C1(n13378), .C2(n13484), .A(n205), .B(n459), .ZN(n14805)
         );
  NAND2_X1 U2770 ( .A1(n13485), .A2(n652), .ZN(n459) );
  OR2_X1 U2772 ( .A1(n18959), .A2(n19470), .ZN(n18961) );
  NAND2_X1 U2773 ( .A1(n12272), .A2(n12864), .ZN(n13115) );
  AOI22_X1 U2775 ( .A1(n21919), .A2(n329), .B1(n22451), .B2(n22323), .ZN(
        n21920) );
  NAND2_X1 U2777 ( .A1(n1192), .A2(n1196), .ZN(n7237) );
  NOR2_X1 U2779 ( .A1(n5415), .A2(n22824), .ZN(n462) );
  OAI21_X1 U2780 ( .B1(n23948), .B2(n22826), .A(n463), .ZN(n23949) );
  OAI211_X2 U2782 ( .C1(n10894), .C2(n3119), .A(n465), .B(n464), .ZN(n12020)
         );
  NAND2_X1 U2783 ( .A1(n10892), .A2(n3119), .ZN(n464) );
  NAND2_X1 U2784 ( .A1(n10893), .A2(n11085), .ZN(n465) );
  NAND2_X1 U2786 ( .A1(n470), .A2(n469), .ZN(n468) );
  NAND2_X1 U2790 ( .A1(n7192), .A2(n8371), .ZN(n472) );
  NAND2_X1 U2791 ( .A1(n17142), .A2(n17141), .ZN(n473) );
  NAND2_X1 U2793 ( .A1(n3306), .A2(n16611), .ZN(n16614) );
  NAND3_X1 U2794 ( .A1(n7828), .A2(n7829), .A3(n7827), .ZN(n7830) );
  NAND2_X1 U2795 ( .A1(n1694), .A2(n12965), .ZN(n12968) );
  NAND2_X1 U2796 ( .A1(n477), .A2(n475), .ZN(n7717) );
  NAND2_X1 U2797 ( .A1(n8371), .A2(n24577), .ZN(n475) );
  NAND2_X1 U2799 ( .A1(n7715), .A2(n24878), .ZN(n477) );
  NAND3_X1 U2800 ( .A1(n16509), .A2(n16508), .A3(n25376), .ZN(n1812) );
  OAI211_X1 U2802 ( .C1(n16235), .C2(n257), .A(n478), .B(n385), .ZN(n14974) );
  NAND2_X1 U2803 ( .A1(n16235), .A2(n16450), .ZN(n478) );
  NAND2_X1 U2804 ( .A1(n480), .A2(n479), .ZN(n10769) );
  NAND3_X1 U2805 ( .A1(n10767), .A2(n10890), .A3(n4422), .ZN(n479) );
  NAND2_X1 U2806 ( .A1(n10768), .A2(n412), .ZN(n480) );
  MUX2_X1 U2807 ( .A(n23967), .B(n25017), .S(n23972), .Z(n23959) );
  OAI211_X2 U2810 ( .C1(n1604), .C2(n20369), .A(n484), .B(n483), .ZN(n21750)
         );
  NAND2_X1 U2811 ( .A1(n277), .A2(n24454), .ZN(n483) );
  NAND2_X1 U2812 ( .A1(n20370), .A2(n24531), .ZN(n484) );
  NAND2_X1 U2814 ( .A1(n17129), .A2(n17132), .ZN(n486) );
  XNOR2_X1 U2815 ( .A(n488), .B(n11348), .ZN(n11349) );
  XNOR2_X1 U2816 ( .A(n11347), .B(n11346), .ZN(n488) );
  NAND3_X1 U2817 ( .A1(n4013), .A2(n413), .A3(n10830), .ZN(n9646) );
  NAND3_X1 U2818 ( .A1(n4774), .A2(n17166), .A3(n25219), .ZN(n514) );
  NAND3_X1 U2822 ( .A1(n2485), .A2(n5624), .A3(n13353), .ZN(n2484) );
  NAND2_X1 U2823 ( .A1(n6718), .A2(n6712), .ZN(n6713) );
  NAND2_X1 U2824 ( .A1(n16193), .A2(n16191), .ZN(n15677) );
  NAND3_X1 U2829 ( .A1(n2728), .A2(n4554), .A3(n2727), .ZN(n492) );
  INV_X1 U2831 ( .A(Plaintext[65]), .ZN(n495) );
  NAND3_X1 U2832 ( .A1(n9454), .A2(n9564), .A3(n9885), .ZN(n2720) );
  OAI211_X1 U2833 ( .C1(n5269), .C2(n15921), .A(n496), .B(n389), .ZN(n15779)
         );
  NAND2_X1 U2834 ( .A1(n16464), .A2(n15921), .ZN(n496) );
  NAND2_X1 U2835 ( .A1(n13307), .A2(n11722), .ZN(n13309) );
  OR2_X1 U2838 ( .A1(n10201), .A2(n5323), .ZN(n498) );
  NAND3_X1 U2839 ( .A1(n1080), .A2(n4332), .A3(n499), .ZN(n1081) );
  AND2_X1 U2840 ( .A1(n6622), .A2(n6114), .ZN(n500) );
  NAND2_X1 U2842 ( .A1(n1609), .A2(n6114), .ZN(n505) );
  NAND2_X1 U2843 ( .A1(n1609), .A2(n500), .ZN(n504) );
  NAND2_X1 U2844 ( .A1(n505), .A2(n501), .ZN(n1610) );
  NAND2_X1 U2845 ( .A1(n6619), .A2(n316), .ZN(n501) );
  NAND3_X1 U2846 ( .A1(n6619), .A2(n6622), .A3(n316), .ZN(n502) );
  INV_X1 U2847 ( .A(n507), .ZN(n3302) );
  NOR2_X1 U2848 ( .A1(n508), .A2(n14158), .ZN(n13467) );
  NAND2_X1 U2849 ( .A1(n508), .A2(n14158), .ZN(n13776) );
  NOR2_X1 U2851 ( .A1(n5080), .A2(n24999), .ZN(n11022) );
  NAND2_X1 U2852 ( .A1(n5079), .A2(n507), .ZN(n13469) );
  OR2_X1 U2853 ( .A1(n22634), .A2(n22633), .ZN(n510) );
  NAND2_X1 U2854 ( .A1(n22636), .A2(n510), .ZN(n22641) );
  NAND2_X1 U2856 ( .A1(n512), .A2(n25253), .ZN(n7914) );
  NAND2_X1 U2857 ( .A1(n512), .A2(n7449), .ZN(n6486) );
  NAND2_X1 U2858 ( .A1(n3347), .A2(n511), .ZN(n7398) );
  AND2_X1 U2859 ( .A1(n512), .A2(n7918), .ZN(n511) );
  NAND2_X1 U2860 ( .A1(n430), .A2(n312), .ZN(n8075) );
  NAND3_X1 U2861 ( .A1(n3348), .A2(n512), .A3(n435), .ZN(n7159) );
  NAND3_X1 U2862 ( .A1(n2376), .A2(n2679), .A3(n22592), .ZN(n710) );
  OR2_X1 U2863 ( .A1(n25475), .A2(n8839), .ZN(n5277) );
  AOI21_X1 U2865 ( .B1(n20041), .B2(n20039), .A(n19862), .ZN(n513) );
  NAND2_X1 U2868 ( .A1(n515), .A2(n1841), .ZN(n18473) );
  NAND2_X1 U2869 ( .A1(n517), .A2(n516), .ZN(n17088) );
  OAI22_X1 U2870 ( .A1(n15536), .A2(n15788), .B1(n15535), .B2(n2253), .ZN(n517) );
  OR2_X1 U2871 ( .A1(n16231), .A2(n16232), .ZN(n15935) );
  OAI22_X1 U2872 ( .A1(n2814), .A2(n16739), .B1(n371), .B2(n16649), .ZN(n17090) );
  AOI22_X2 U2873 ( .A1(n5471), .A2(n12206), .B1(n5472), .B2(n3876), .ZN(n13460) );
  XNOR2_X1 U2874 ( .A(n12207), .B(n455), .ZN(n12208) );
  OAI21_X1 U2877 ( .B1(n19400), .B2(n18900), .A(n19163), .ZN(n519) );
  NAND2_X1 U2880 ( .A1(n23995), .A2(n25079), .ZN(n520) );
  OR2_X1 U2881 ( .A1(n10308), .A2(n4998), .ZN(n758) );
  NAND2_X1 U2882 ( .A1(n6341), .A2(n6187), .ZN(n6448) );
  NOR2_X1 U2883 ( .A1(n521), .A2(n15676), .ZN(n15678) );
  NAND2_X1 U2884 ( .A1(n523), .A2(n17449), .ZN(n522) );
  NAND2_X1 U2887 ( .A1(n2714), .A2(n10552), .ZN(n3196) );
  NAND3_X2 U2889 ( .A1(n10526), .A2(n525), .A3(n10525), .ZN(n12277) );
  NAND2_X1 U2890 ( .A1(n3556), .A2(n3555), .ZN(n16112) );
  NAND2_X1 U2892 ( .A1(n10013), .A2(n4531), .ZN(n526) );
  NAND2_X1 U2893 ( .A1(n10014), .A2(n528), .ZN(n527) );
  NAND2_X1 U2896 ( .A1(n11046), .A2(n11044), .ZN(n529) );
  INV_X1 U2897 ( .A(n10158), .ZN(n3305) );
  OR2_X1 U2898 ( .A1(n1100), .A2(n22359), .ZN(n972) );
  NOR2_X1 U2899 ( .A1(n5475), .A2(n20257), .ZN(n5473) );
  INV_X1 U2900 ( .A(n20255), .ZN(n20412) );
  NAND2_X1 U2901 ( .A1(n10242), .A2(n10497), .ZN(n531) );
  NAND2_X1 U2902 ( .A1(n10241), .A2(n2546), .ZN(n532) );
  NAND2_X1 U2903 ( .A1(n14075), .A2(n14076), .ZN(n13629) );
  OR2_X1 U2905 ( .A1(n25046), .A2(n8327), .ZN(n9591) );
  OR2_X1 U2906 ( .A1(n20422), .A2(n20419), .ZN(n1660) );
  NAND2_X1 U2907 ( .A1(n17160), .A2(n17163), .ZN(n16264) );
  NAND2_X1 U2910 ( .A1(n21293), .A2(n22771), .ZN(n535) );
  OAI21_X1 U2912 ( .B1(n23833), .B2(n23827), .A(n318), .ZN(n536) );
  NAND2_X1 U2913 ( .A1(n537), .A2(n11125), .ZN(n9243) );
  OAI22_X1 U2914 ( .A1(n305), .A2(n10460), .B1(n11124), .B2(n10850), .ZN(n537)
         );
  NAND2_X1 U2915 ( .A1(n16035), .A2(n16733), .ZN(n2096) );
  OAI21_X1 U2916 ( .B1(n13030), .B2(n302), .A(n538), .ZN(n12494) );
  NAND2_X1 U2917 ( .A1(n12786), .A2(n13023), .ZN(n538) );
  AOI22_X1 U2918 ( .A1(n3627), .A2(n3783), .B1(n3626), .B2(n17316), .ZN(n539)
         );
  INV_X1 U2919 ( .A(n542), .ZN(n541) );
  OAI21_X1 U2920 ( .B1(n11175), .B2(n10940), .A(n10939), .ZN(n542) );
  NAND2_X1 U2921 ( .A1(n543), .A2(n1375), .ZN(n11242) );
  NAND2_X1 U2923 ( .A1(n12624), .A2(n12878), .ZN(n5191) );
  NAND2_X1 U2924 ( .A1(n14182), .A2(n14178), .ZN(n13797) );
  INV_X1 U2925 ( .A(n13234), .ZN(n545) );
  NAND2_X1 U2926 ( .A1(n12936), .A2(n13234), .ZN(n546) );
  NAND2_X1 U2929 ( .A1(n18903), .A2(n353), .ZN(n548) );
  NAND2_X1 U2930 ( .A1(n18904), .A2(n3773), .ZN(n549) );
  OAI211_X1 U2935 ( .C1(n22624), .C2(n23058), .A(n553), .B(n552), .ZN(n22626)
         );
  NAND2_X1 U2936 ( .A1(n22643), .A2(n23059), .ZN(n552) );
  NAND2_X1 U2937 ( .A1(n23055), .A2(n22698), .ZN(n553) );
  NAND2_X1 U2938 ( .A1(n23301), .A2(n554), .ZN(n664) );
  AOI22_X1 U2939 ( .A1(n23298), .A2(n23297), .B1(n23300), .B2(n23299), .ZN(
        n554) );
  INV_X1 U2940 ( .A(n19422), .ZN(n1309) );
  NAND3_X1 U2941 ( .A1(n555), .A2(n4475), .A3(n4474), .ZN(n23977) );
  NAND2_X1 U2942 ( .A1(n23975), .A2(n23987), .ZN(n555) );
  INV_X1 U2944 ( .A(n557), .ZN(n556) );
  OAI21_X1 U2945 ( .B1(n9827), .B2(n10186), .A(n9586), .ZN(n557) );
  NAND2_X1 U2946 ( .A1(n561), .A2(n558), .ZN(n10345) );
  NAND2_X1 U2947 ( .A1(n560), .A2(n559), .ZN(n558) );
  INV_X1 U2948 ( .A(n10341), .ZN(n560) );
  NAND2_X1 U2949 ( .A1(n10342), .A2(n10411), .ZN(n561) );
  OR2_X1 U2951 ( .A1(n16106), .A2(n16108), .ZN(n15854) );
  INV_X1 U2952 ( .A(n13074), .ZN(n12708) );
  NAND2_X1 U2953 ( .A1(n4124), .A2(n562), .ZN(n4123) );
  NAND2_X1 U2954 ( .A1(n13029), .A2(n563), .ZN(n562) );
  NAND3_X2 U2955 ( .A1(n564), .A2(n15079), .A3(n15080), .ZN(n17424) );
  NAND2_X1 U2957 ( .A1(n13350), .A2(n12349), .ZN(n12330) );
  NAND3_X1 U2959 ( .A1(n424), .A2(n10089), .A3(n1348), .ZN(n9784) );
  XNOR2_X1 U2960 ( .A(n565), .B(n22875), .ZN(Ciphertext[9]) );
  OAI211_X1 U2961 ( .C1(n24350), .C2(n22578), .A(n1197), .B(n22873), .ZN(n565)
         );
  NAND2_X1 U2962 ( .A1(n4165), .A2(n2815), .ZN(n566) );
  NAND2_X1 U2963 ( .A1(n17090), .A2(n17091), .ZN(n567) );
  OR2_X1 U2964 ( .A1(n6742), .A2(n6104), .ZN(n568) );
  NAND2_X1 U2965 ( .A1(n7280), .A2(n8512), .ZN(n569) );
  OAI22_X1 U2966 ( .A1(n21930), .A2(n22465), .B1(n22462), .B2(n22459), .ZN(
        n570) );
  NAND2_X1 U2967 ( .A1(n17032), .A2(n571), .ZN(n18073) );
  NAND2_X1 U2968 ( .A1(n2111), .A2(n572), .ZN(n571) );
  NAND2_X1 U2970 ( .A1(n574), .A2(n573), .ZN(n2032) );
  INV_X1 U2971 ( .A(n24037), .ZN(n573) );
  NAND2_X1 U2972 ( .A1(n6921), .A2(n6920), .ZN(n574) );
  NAND2_X1 U2973 ( .A1(n25366), .A2(n25415), .ZN(n2422) );
  OAI21_X2 U2975 ( .B1(n16842), .B2(n17166), .A(n16841), .ZN(n18121) );
  NAND2_X1 U2977 ( .A1(n10858), .A2(n10860), .ZN(n10280) );
  NAND2_X1 U2978 ( .A1(n5064), .A2(n9250), .ZN(n10860) );
  OR2_X1 U2979 ( .A1(n10099), .A2(n10100), .ZN(n4302) );
  NAND2_X1 U2981 ( .A1(n19599), .A2(n19598), .ZN(n576) );
  NAND2_X1 U2983 ( .A1(n579), .A2(n25449), .ZN(n578) );
  INV_X1 U2984 ( .A(n16123), .ZN(n579) );
  OAI211_X1 U2985 ( .C1(n1231), .C2(n16957), .A(n1230), .B(n1229), .ZN(n1228)
         );
  NAND3_X1 U2986 ( .A1(n580), .A2(n1482), .A3(n2066), .ZN(n1722) );
  AND2_X1 U2988 ( .A1(n339), .A2(n19883), .ZN(n19916) );
  NAND2_X1 U2989 ( .A1(n1551), .A2(n4842), .ZN(n4841) );
  NAND2_X1 U2990 ( .A1(n7666), .A2(n7665), .ZN(n8534) );
  NAND2_X1 U2991 ( .A1(n581), .A2(n2121), .ZN(n16531) );
  NAND2_X1 U2992 ( .A1(n16526), .A2(n17451), .ZN(n581) );
  NAND2_X1 U2993 ( .A1(n2223), .A2(n584), .ZN(n7687) );
  NAND2_X1 U2994 ( .A1(n9675), .A2(n9674), .ZN(n1346) );
  AND2_X2 U2995 ( .A1(n586), .A2(n585), .ZN(n21985) );
  NAND2_X1 U2996 ( .A1(n20302), .A2(n20301), .ZN(n585) );
  NAND2_X1 U2997 ( .A1(n20300), .A2(n20299), .ZN(n586) );
  OAI21_X1 U2998 ( .B1(n12526), .B2(n25337), .A(n902), .ZN(n11452) );
  AOI21_X1 U3000 ( .B1(n20066), .B2(n20074), .A(n588), .ZN(n587) );
  INV_X1 U3002 ( .A(n15584), .ZN(n16105) );
  OR2_X1 U3003 ( .A1(n6195), .A2(n6444), .ZN(n640) );
  NAND2_X1 U3004 ( .A1(n589), .A2(n4044), .ZN(n15841) );
  NAND2_X1 U3005 ( .A1(n692), .A2(n4045), .ZN(n589) );
  OAI21_X1 U3006 ( .B1(n429), .B2(n10060), .A(n590), .ZN(n10067) );
  NAND2_X1 U3007 ( .A1(n10060), .A2(n10061), .ZN(n590) );
  OR2_X1 U3008 ( .A1(n17093), .A2(n24410), .ZN(n17687) );
  BUF_X2 U3009 ( .A(n6374), .Z(n6904) );
  NAND3_X1 U3010 ( .A1(n24468), .A2(n21840), .A3(n21822), .ZN(n21296) );
  NAND2_X1 U3014 ( .A1(n22403), .A2(n21885), .ZN(n593) );
  NAND2_X1 U3016 ( .A1(n6128), .A2(n6530), .ZN(n6129) );
  AOI21_X1 U3019 ( .B1(n907), .B2(n905), .A(n142), .ZN(n595) );
  NAND2_X1 U3020 ( .A1(n6257), .A2(n6256), .ZN(n2824) );
  NAND2_X1 U3022 ( .A1(n4906), .A2(n13094), .ZN(n598) );
  NAND2_X1 U3024 ( .A1(n11410), .A2(n11409), .ZN(n2117) );
  AND3_X2 U3025 ( .A1(n599), .A2(n13649), .A3(n13650), .ZN(n14104) );
  OAI211_X2 U3027 ( .C1(n20567), .C2(n20566), .A(n24530), .B(n600), .ZN(n21579) );
  NAND2_X1 U3028 ( .A1(n20565), .A2(n20564), .ZN(n600) );
  NAND2_X1 U3029 ( .A1(n20502), .A2(n20501), .ZN(n5424) );
  NAND2_X1 U3030 ( .A1(n605), .A2(n602), .ZN(n22854) );
  INV_X1 U3032 ( .A(n5421), .ZN(n603) );
  NAND2_X1 U3034 ( .A1(n22855), .A2(n24356), .ZN(n605) );
  INV_X1 U3035 ( .A(n14382), .ZN(n15620) );
  NAND3_X1 U3036 ( .A1(n10253), .A2(n10730), .A3(n606), .ZN(n10262) );
  OR2_X1 U3037 ( .A1(n10255), .A2(n10254), .ZN(n606) );
  NAND2_X1 U3038 ( .A1(n10254), .A2(n10129), .ZN(n10251) );
  AND2_X2 U3042 ( .A1(n2048), .A2(n1471), .ZN(n14327) );
  OAI21_X2 U3046 ( .B1(n16653), .B2(n16652), .A(n16651), .ZN(n18239) );
  NAND2_X1 U3047 ( .A1(n611), .A2(n610), .ZN(n9839) );
  NAND2_X1 U3048 ( .A1(n428), .A2(n8359), .ZN(n610) );
  NAND2_X1 U3049 ( .A1(n9838), .A2(n9837), .ZN(n611) );
  NAND2_X1 U3050 ( .A1(n10094), .A2(n9515), .ZN(n9838) );
  XNOR2_X2 U3052 ( .A(n17511), .B(n17512), .ZN(n19297) );
  NAND2_X1 U3053 ( .A1(n7887), .A2(n7883), .ZN(n3130) );
  NAND2_X1 U3054 ( .A1(n7882), .A2(n7585), .ZN(n7887) );
  NAND2_X1 U3057 ( .A1(n380), .A2(n16064), .ZN(n613) );
  AND2_X1 U3058 ( .A1(n22262), .A2(n1276), .ZN(n22135) );
  NAND2_X1 U3059 ( .A1(n615), .A2(n614), .ZN(n19715) );
  NAND2_X1 U3060 ( .A1(n20319), .A2(n19889), .ZN(n614) );
  NOR2_X1 U3061 ( .A1(n616), .A2(n7427), .ZN(n7199) );
  NAND2_X1 U3062 ( .A1(n7812), .A2(n9068), .ZN(n616) );
  INV_X1 U3063 ( .A(n617), .ZN(n16053) );
  NAND2_X1 U3064 ( .A1(n24352), .A2(n15706), .ZN(n617) );
  NOR2_X1 U3066 ( .A1(n14131), .A2(n620), .ZN(n14133) );
  NAND2_X1 U3067 ( .A1(n619), .A2(n618), .ZN(n12941) );
  NAND2_X1 U3068 ( .A1(n5751), .A2(n14132), .ZN(n618) );
  NOR2_X1 U3070 ( .A1(n1508), .A2(n12597), .ZN(n623) );
  NAND2_X1 U3071 ( .A1(n12912), .A2(n1508), .ZN(n624) );
  NAND2_X1 U3073 ( .A1(n25424), .A2(n625), .ZN(n7031) );
  NAND2_X1 U3074 ( .A1(n625), .A2(n6104), .ZN(n6005) );
  NAND3_X1 U3075 ( .A1(n6593), .A2(n6592), .A3(n626), .ZN(n6594) );
  NAND2_X1 U3076 ( .A1(n454), .A2(n7033), .ZN(n626) );
  NOR2_X1 U3077 ( .A1(n9398), .A2(n9365), .ZN(n627) );
  AND2_X1 U3078 ( .A1(n10136), .A2(n24026), .ZN(n9201) );
  NAND2_X1 U3079 ( .A1(n14853), .A2(n14852), .ZN(n628) );
  NAND2_X1 U3080 ( .A1(n21286), .A2(n629), .ZN(n21288) );
  OAI211_X1 U3081 ( .C1(n317), .C2(n23229), .A(n23218), .B(n630), .ZN(n629) );
  NAND2_X1 U3082 ( .A1(n317), .A2(n23220), .ZN(n630) );
  INV_X1 U3083 ( .A(n16311), .ZN(n16012) );
  NAND2_X1 U3084 ( .A1(n631), .A2(n16311), .ZN(n633) );
  OAI21_X1 U3085 ( .B1(n2173), .B2(n15198), .A(n632), .ZN(n631) );
  NAND2_X1 U3086 ( .A1(n15198), .A2(n16312), .ZN(n632) );
  NAND2_X1 U3089 ( .A1(n634), .A2(n633), .ZN(n635) );
  OAI21_X1 U3091 ( .B1(n17331), .B2(n635), .A(n17335), .ZN(n17339) );
  NOR2_X1 U3092 ( .A1(n19972), .A2(n636), .ZN(n19973) );
  OAI21_X1 U3093 ( .B1(n20530), .B2(n636), .A(n2852), .ZN(n18886) );
  INV_X1 U3094 ( .A(n20289), .ZN(n636) );
  NAND2_X1 U3095 ( .A1(n637), .A2(n6196), .ZN(n4726) );
  NAND2_X1 U3096 ( .A1(n6448), .A2(n637), .ZN(n4878) );
  NAND2_X1 U3097 ( .A1(n640), .A2(n6188), .ZN(n637) );
  XNOR2_X1 U3098 ( .A(n25390), .B(n447), .ZN(n18241) );
  XNOR2_X1 U3099 ( .A(n25390), .B(n452), .ZN(n16635) );
  XNOR2_X1 U3100 ( .A(n17873), .B(n445), .ZN(n17644) );
  XNOR2_X1 U3101 ( .A(n25390), .B(n449), .ZN(n18125) );
  NOR2_X1 U3102 ( .A1(n372), .A2(n17053), .ZN(n4298) );
  NAND2_X1 U3104 ( .A1(n9358), .A2(n9357), .ZN(n3324) );
  NAND2_X1 U3106 ( .A1(n24398), .A2(n24585), .ZN(n16609) );
  NAND2_X1 U3109 ( .A1(n25408), .A2(n12490), .ZN(n642) );
  NAND2_X1 U3111 ( .A1(n12534), .A2(n12535), .ZN(n12533) );
  NAND2_X1 U3112 ( .A1(n645), .A2(n376), .ZN(n644) );
  NAND2_X1 U3115 ( .A1(n994), .A2(n16266), .ZN(n646) );
  NAND2_X1 U3117 ( .A1(n10594), .A2(n10505), .ZN(n10930) );
  NAND3_X1 U3120 ( .A1(n10688), .A2(n10687), .A3(n10686), .ZN(n10689) );
  OR2_X1 U3121 ( .A1(n17299), .A2(n17297), .ZN(n16702) );
  OR2_X1 U3122 ( .A1(n22782), .A2(n24406), .ZN(n22365) );
  NAND3_X1 U3123 ( .A1(n1198), .A2(n22872), .A3(n22578), .ZN(n1197) );
  NAND3_X2 U3127 ( .A1(n15608), .A2(n879), .A3(n880), .ZN(n17068) );
  NAND2_X1 U3130 ( .A1(n16069), .A2(n4105), .ZN(n649) );
  NAND2_X1 U3131 ( .A1(n651), .A2(n650), .ZN(n21938) );
  NAND2_X1 U3132 ( .A1(n21935), .A2(n326), .ZN(n651) );
  XNOR2_X1 U3133 ( .A(n15222), .B(n15221), .ZN(n16192) );
  NOR2_X1 U3134 ( .A1(n13486), .A2(n24462), .ZN(n652) );
  NAND3_X1 U3135 ( .A1(n10547), .A2(n10705), .A3(n10702), .ZN(n10551) );
  AOI22_X1 U3139 ( .A1(n12866), .A2(n12865), .B1(n1513), .B2(n13114), .ZN(
        n4798) );
  NAND3_X1 U3140 ( .A1(n9456), .A2(n9455), .A3(n9887), .ZN(n957) );
  NAND2_X1 U3142 ( .A1(n657), .A2(n438), .ZN(n656) );
  NAND2_X1 U3143 ( .A1(n6439), .A2(n6438), .ZN(n657) );
  NAND2_X1 U3144 ( .A1(n6440), .A2(n6174), .ZN(n658) );
  NAND3_X2 U3145 ( .A1(n2943), .A2(n7649), .A3(n989), .ZN(n9043) );
  XNOR2_X1 U3146 ( .A(n659), .B(n5598), .ZN(Ciphertext[136]) );
  OAI211_X1 U3147 ( .C1(n23718), .C2(n3283), .A(n3280), .B(n23717), .ZN(n659)
         );
  NOR2_X2 U3148 ( .A1(n11252), .A2(n661), .ZN(n14294) );
  OAI22_X1 U3149 ( .A1(n12987), .A2(n13220), .B1(n4652), .B2(n12767), .ZN(n661) );
  NAND2_X1 U3150 ( .A1(n374), .A2(n662), .ZN(n17044) );
  NAND2_X1 U3151 ( .A1(n24903), .A2(n23303), .ZN(n23295) );
  XNOR2_X1 U3152 ( .A(n664), .B(n23302), .ZN(Ciphertext[57]) );
  NAND3_X1 U3153 ( .A1(n13506), .A2(n13507), .A3(n13505), .ZN(n13508) );
  NAND3_X1 U3154 ( .A1(n4597), .A2(n4600), .A3(n13437), .ZN(n2821) );
  XNOR2_X2 U3155 ( .A(n5822), .B(Key[146]), .ZN(n6377) );
  OAI211_X2 U3156 ( .C1(n17325), .C2(n17326), .A(n207), .B(n206), .ZN(n18447)
         );
  XNOR2_X1 U3157 ( .A(n11768), .B(n11764), .ZN(n667) );
  NAND2_X1 U3159 ( .A1(n6674), .A2(n6675), .ZN(n668) );
  NAND2_X1 U3160 ( .A1(n14584), .A2(n213), .ZN(n14585) );
  XNOR2_X1 U3162 ( .A(n18152), .B(n18147), .ZN(n670) );
  OAI211_X1 U3163 ( .C1(n1771), .C2(n13962), .A(n671), .B(n4293), .ZN(n1770)
         );
  NAND2_X1 U3164 ( .A1(n13962), .A2(n13963), .ZN(n671) );
  AND2_X2 U3165 ( .A1(n3744), .A2(n15768), .ZN(n16809) );
  NAND3_X1 U3166 ( .A1(n2003), .A2(n2002), .A3(n672), .ZN(n14976) );
  NOR2_X1 U3168 ( .A1(n16851), .A2(n1653), .ZN(n16847) );
  NAND3_X1 U3169 ( .A1(n674), .A2(n6494), .A3(n6489), .ZN(n6492) );
  NAND2_X1 U3170 ( .A1(n6487), .A2(n6488), .ZN(n674) );
  NAND3_X1 U3171 ( .A1(n675), .A2(n9884), .A3(n9563), .ZN(n9891) );
  NAND2_X1 U3172 ( .A1(n9883), .A2(n9882), .ZN(n675) );
  OAI211_X1 U3173 ( .C1(n7634), .C2(n7918), .A(n312), .B(n920), .ZN(n1280) );
  NAND2_X1 U3174 ( .A1(n7923), .A2(n5607), .ZN(n1088) );
  NAND2_X1 U3175 ( .A1(n12833), .A2(n5645), .ZN(n12850) );
  NAND2_X1 U3176 ( .A1(n9419), .A2(n9613), .ZN(n9972) );
  NAND2_X1 U3177 ( .A1(n1345), .A2(n270), .ZN(n2223) );
  AND2_X1 U3179 ( .A1(n2677), .A2(n710), .ZN(n5259) );
  NAND2_X1 U3180 ( .A1(n676), .A2(n13055), .ZN(n13059) );
  NOR2_X1 U3181 ( .A1(n409), .A2(n13057), .ZN(n676) );
  OR2_X1 U3182 ( .A1(n1248), .A2(n22359), .ZN(n782) );
  NAND2_X1 U3183 ( .A1(n2939), .A2(n401), .ZN(n2938) );
  NAND2_X1 U3184 ( .A1(n1962), .A2(n1961), .ZN(n1959) );
  OAI21_X1 U3185 ( .B1(n11085), .B2(n418), .A(n678), .ZN(n10894) );
  NAND2_X1 U3186 ( .A1(n11085), .A2(n10890), .ZN(n678) );
  XNOR2_X1 U3187 ( .A(n14827), .B(n15446), .ZN(n14430) );
  INV_X1 U3188 ( .A(n16572), .ZN(n17116) );
  OAI211_X1 U3189 ( .C1(n19070), .C2(n19612), .A(n19069), .B(n19068), .ZN(
        n1155) );
  NAND3_X1 U3192 ( .A1(n7841), .A2(n8370), .A3(n7843), .ZN(n7842) );
  NAND2_X1 U3194 ( .A1(n680), .A2(n4753), .ZN(n7578) );
  NAND2_X1 U3195 ( .A1(n4751), .A2(n4752), .ZN(n680) );
  NAND2_X1 U3196 ( .A1(n10684), .A2(n10363), .ZN(n3934) );
  NAND2_X1 U3197 ( .A1(n6405), .A2(n6404), .ZN(n1558) );
  NAND2_X1 U3199 ( .A1(n4806), .A2(n4807), .ZN(n693) );
  NAND2_X1 U3200 ( .A1(n2090), .A2(n16109), .ZN(n682) );
  NAND2_X1 U3201 ( .A1(n4689), .A2(n379), .ZN(n683) );
  OAI22_X1 U3204 ( .A1(n442), .A2(n249), .B1(n7021), .B2(n7026), .ZN(n6638) );
  NAND2_X1 U3205 ( .A1(n13548), .A2(n13551), .ZN(n684) );
  OAI21_X1 U3207 ( .B1(n707), .B2(n16170), .A(n706), .ZN(n15960) );
  NAND3_X1 U3208 ( .A1(n685), .A2(n12461), .A3(n12482), .ZN(n3454) );
  INV_X1 U3209 ( .A(n12709), .ZN(n685) );
  OAI22_X1 U3210 ( .A1(n16031), .A2(n24403), .B1(n16276), .B2(n16274), .ZN(
        n16032) );
  NAND2_X1 U3212 ( .A1(n3050), .A2(n4369), .ZN(n7421) );
  NAND2_X1 U3213 ( .A1(n16534), .A2(n16533), .ZN(n686) );
  NAND2_X1 U3216 ( .A1(n6380), .A2(n6379), .ZN(n4641) );
  XNOR2_X1 U3217 ( .A(n11796), .B(n12138), .ZN(n11469) );
  NAND2_X1 U3220 ( .A1(n16973), .A2(n17336), .ZN(n16726) );
  NAND2_X1 U3221 ( .A1(n25462), .A2(n25022), .ZN(n21146) );
  NAND2_X1 U3224 ( .A1(n19611), .A2(n2764), .ZN(n1590) );
  NAND2_X1 U3225 ( .A1(n13417), .A2(n24503), .ZN(n689) );
  NAND2_X1 U3226 ( .A1(n25278), .A2(n14099), .ZN(n690) );
  NAND3_X1 U3229 ( .A1(n693), .A2(n16686), .A3(n3723), .ZN(n17248) );
  NAND2_X1 U3230 ( .A1(n24339), .A2(n324), .ZN(n23389) );
  NAND2_X1 U3232 ( .A1(n731), .A2(n800), .ZN(n7214) );
  NAND3_X1 U3233 ( .A1(n3169), .A2(n14748), .A3(n16762), .ZN(n829) );
  AOI21_X1 U3235 ( .B1(n22848), .B2(n21709), .A(n22907), .ZN(n695) );
  OR2_X2 U3236 ( .A1(n722), .A2(n2449), .ZN(n12414) );
  NAND2_X1 U3238 ( .A1(n5633), .A2(n19191), .ZN(n5632) );
  NAND2_X1 U3239 ( .A1(n18923), .A2(n696), .ZN(n17011) );
  NAND2_X1 U3240 ( .A1(n14180), .A2(n14178), .ZN(n13771) );
  INV_X1 U3241 ( .A(n697), .ZN(n22269) );
  OAI22_X1 U3242 ( .A1(n22268), .A2(n22267), .B1(n22266), .B2(n25381), .ZN(
        n697) );
  NAND3_X1 U3245 ( .A1(n822), .A2(n821), .A3(n699), .ZN(n698) );
  NAND2_X1 U3247 ( .A1(n15314), .A2(n17342), .ZN(n16778) );
  NAND2_X1 U3249 ( .A1(n6037), .A2(n6503), .ZN(n703) );
  OAI21_X1 U3250 ( .B1(n13840), .B2(n397), .A(n704), .ZN(n13842) );
  NAND2_X1 U3251 ( .A1(n13840), .A2(n13837), .ZN(n704) );
  NAND3_X1 U3252 ( .A1(n13189), .A2(n3957), .A3(n13190), .ZN(n14108) );
  NAND3_X1 U3253 ( .A1(n9657), .A2(n9996), .A3(n9658), .ZN(n867) );
  OR2_X1 U3254 ( .A1(n16266), .A2(n16268), .ZN(n992) );
  AND2_X1 U3255 ( .A1(n14290), .A2(n13907), .ZN(n11454) );
  OR3_X1 U3256 ( .A1(n19393), .A2(n18788), .A3(n24407), .ZN(n18789) );
  OAI21_X1 U3257 ( .B1(n6329), .B2(n4621), .A(n6471), .ZN(n1078) );
  OAI21_X1 U3258 ( .B1(n406), .B2(n25430), .A(n705), .ZN(n12875) );
  NAND2_X1 U3259 ( .A1(n13352), .A2(n13353), .ZN(n705) );
  NAND2_X1 U3262 ( .A1(n6049), .A2(n6623), .ZN(n6624) );
  NAND2_X1 U3263 ( .A1(n1918), .A2(n11208), .ZN(n11211) );
  NAND2_X1 U3265 ( .A1(n6425), .A2(n198), .ZN(n2542) );
  NAND2_X1 U3267 ( .A1(n9979), .A2(n712), .ZN(n711) );
  INV_X1 U3268 ( .A(n713), .ZN(n712) );
  OAI21_X1 U3269 ( .B1(n9429), .B2(n9981), .A(n9980), .ZN(n713) );
  NAND3_X1 U3271 ( .A1(n10156), .A2(n25206), .A3(n10120), .ZN(n2254) );
  NAND3_X1 U3272 ( .A1(n5277), .A2(n25007), .A3(n5278), .ZN(n5272) );
  INV_X1 U3273 ( .A(n716), .ZN(Ciphertext[116]) );
  OAI211_X1 U3274 ( .C1(n21952), .C2(n21951), .A(n21949), .B(n21950), .ZN(n716) );
  NAND2_X1 U3275 ( .A1(n7212), .A2(n8530), .ZN(n800) );
  NAND3_X1 U3276 ( .A1(n346), .A2(n20486), .A3(n19634), .ZN(n19638) );
  NAND2_X1 U3277 ( .A1(n17255), .A2(n16561), .ZN(n17257) );
  NAND2_X1 U3279 ( .A1(n7720), .A2(n7719), .ZN(n8730) );
  NAND3_X1 U3280 ( .A1(n719), .A2(n1465), .A3(n718), .ZN(n23956) );
  NAND2_X1 U3281 ( .A1(n23953), .A2(n23969), .ZN(n718) );
  NAND2_X1 U3282 ( .A1(n23954), .A2(n23955), .ZN(n719) );
  OAI211_X2 U3283 ( .C1(n3971), .C2(n13162), .A(n3970), .B(n3969), .ZN(n1355)
         );
  NAND2_X1 U3284 ( .A1(n19190), .A2(n20511), .ZN(n837) );
  OR2_X2 U3286 ( .A1(n720), .A2(n4941), .ZN(n3725) );
  NAND2_X1 U3288 ( .A1(n721), .A2(n23011), .ZN(n23493) );
  NAND2_X1 U3289 ( .A1(n23480), .A2(n2710), .ZN(n721) );
  AOI21_X1 U3290 ( .B1(n10657), .B2(n10656), .A(n10661), .ZN(n722) );
  AOI21_X1 U3291 ( .B1(n10727), .B2(n10726), .A(n10868), .ZN(n1900) );
  NAND2_X1 U3292 ( .A1(n10286), .A2(n1658), .ZN(n10727) );
  XNOR2_X1 U3295 ( .A(n14979), .B(n14980), .ZN(n14981) );
  OAI211_X2 U3296 ( .C1(n13526), .C2(n13527), .A(n3329), .B(n3331), .ZN(n14979) );
  NAND2_X1 U3297 ( .A1(n12862), .A2(n725), .ZN(n13871) );
  NAND2_X1 U3298 ( .A1(n12858), .A2(n12863), .ZN(n725) );
  NAND2_X1 U3300 ( .A1(n13602), .A2(n14317), .ZN(n13603) );
  NAND2_X1 U3301 ( .A1(n17304), .A2(n17305), .ZN(n1244) );
  NAND2_X1 U3302 ( .A1(n14302), .A2(n14306), .ZN(n13889) );
  OAI21_X1 U3303 ( .B1(n6718), .B2(n24051), .A(n24500), .ZN(n6237) );
  NAND2_X1 U3305 ( .A1(n313), .A2(n6893), .ZN(n6816) );
  XNOR2_X2 U3306 ( .A(n5826), .B(Key[137]), .ZN(n6893) );
  NAND2_X1 U3307 ( .A1(n20317), .A2(n340), .ZN(n4960) );
  NAND2_X1 U3308 ( .A1(n17503), .A2(n17502), .ZN(n727) );
  INV_X1 U3309 ( .A(n2229), .ZN(n728) );
  NAND3_X1 U3313 ( .A1(n2325), .A2(n17227), .A3(n16954), .ZN(n4974) );
  NAND2_X1 U3314 ( .A1(n798), .A2(n7665), .ZN(n731) );
  NAND2_X1 U3316 ( .A1(n732), .A2(n19162), .ZN(n1979) );
  NAND2_X1 U3317 ( .A1(n3726), .A2(n19163), .ZN(n732) );
  NAND2_X1 U3318 ( .A1(n13212), .A2(n13211), .ZN(n13005) );
  NAND2_X1 U3319 ( .A1(n733), .A2(n16734), .ZN(n16735) );
  NAND2_X1 U3320 ( .A1(n16733), .A2(n16732), .ZN(n733) );
  NAND2_X1 U3321 ( .A1(n6904), .A2(n6089), .ZN(n6090) );
  NAND3_X1 U3323 ( .A1(n1058), .A2(n2878), .A3(n11302), .ZN(n734) );
  OAI21_X1 U3324 ( .B1(n10650), .B2(n10651), .A(n735), .ZN(n10652) );
  NAND3_X2 U3325 ( .A1(n737), .A2(n736), .A3(n8004), .ZN(n8965) );
  NAND2_X1 U3326 ( .A1(n7756), .A2(n7755), .ZN(n737) );
  NAND4_X1 U3331 ( .A1(n741), .A2(n14367), .A3(n14366), .A4(n740), .ZN(n14368)
         );
  NAND2_X1 U3332 ( .A1(n14363), .A2(n5526), .ZN(n740) );
  NAND2_X1 U3333 ( .A1(n14365), .A2(n14364), .ZN(n741) );
  NAND2_X1 U3334 ( .A1(n19395), .A2(n19162), .ZN(n18790) );
  NAND3_X1 U3338 ( .A1(n4215), .A2(n21366), .A3(n21365), .ZN(Ciphertext[160])
         );
  NAND2_X1 U3339 ( .A1(n16347), .A2(n25441), .ZN(n2702) );
  NAND2_X1 U3340 ( .A1(n744), .A2(n743), .ZN(n1832) );
  AOI21_X1 U3341 ( .B1(n24080), .B2(n15822), .A(n16597), .ZN(n743) );
  NAND2_X1 U3342 ( .A1(n16595), .A2(n24467), .ZN(n744) );
  NAND3_X1 U3343 ( .A1(n10134), .A2(n10141), .A3(n10138), .ZN(n9370) );
  INV_X1 U3346 ( .A(n16398), .ZN(n746) );
  NAND2_X1 U3348 ( .A1(n3937), .A2(n22461), .ZN(n747) );
  NAND2_X1 U3349 ( .A1(n24253), .A2(n24592), .ZN(n6015) );
  OR2_X1 U3352 ( .A1(n16546), .A2(n17068), .ZN(n1071) );
  NAND2_X1 U3353 ( .A1(n24973), .A2(n749), .ZN(n2303) );
  NAND3_X2 U3355 ( .A1(n751), .A2(n16617), .A3(n752), .ZN(n18431) );
  NAND2_X1 U3356 ( .A1(n3377), .A2(n469), .ZN(n752) );
  OAI21_X1 U3357 ( .B1(n19817), .B2(n754), .A(n753), .ZN(n19512) );
  NAND2_X1 U3358 ( .A1(n19817), .A2(n1344), .ZN(n753) );
  NAND2_X1 U3360 ( .A1(n757), .A2(n756), .ZN(n15718) );
  NAND2_X1 U3361 ( .A1(n24981), .A2(n15951), .ZN(n756) );
  NAND3_X1 U3362 ( .A1(n10307), .A2(n759), .A3(n758), .ZN(n11776) );
  OAI21_X1 U3363 ( .B1(n10305), .B2(n10306), .A(n4998), .ZN(n759) );
  NAND2_X1 U3366 ( .A1(n762), .A2(n19543), .ZN(n3665) );
  NAND2_X1 U3367 ( .A1(n2879), .A2(n7010), .ZN(n764) );
  NAND2_X1 U3369 ( .A1(n766), .A2(n437), .ZN(n1192) );
  NAND2_X1 U3370 ( .A1(n7235), .A2(n7961), .ZN(n766) );
  NAND3_X1 U3372 ( .A1(n6153), .A2(n6277), .A3(n440), .ZN(n767) );
  NAND2_X1 U3374 ( .A1(n1160), .A2(n1161), .ZN(n1159) );
  NAND2_X1 U3375 ( .A1(n5744), .A2(n1689), .ZN(n11133) );
  NOR2_X1 U3376 ( .A1(n420), .A2(n10838), .ZN(n5744) );
  NAND2_X1 U3377 ( .A1(n12597), .A2(n12824), .ZN(n12690) );
  NAND2_X1 U3378 ( .A1(n770), .A2(n769), .ZN(n14080) );
  NAND2_X1 U3380 ( .A1(n14076), .A2(n396), .ZN(n770) );
  NAND3_X1 U3381 ( .A1(n771), .A2(n20370), .A3(n349), .ZN(n3430) );
  NAND2_X1 U3382 ( .A1(n6556), .A2(n6697), .ZN(n1961) );
  NAND2_X1 U3383 ( .A1(n19581), .A2(n19579), .ZN(n18880) );
  OAI22_X1 U3385 ( .A1(n3211), .A2(n3212), .B1(n3210), .B2(n22972), .ZN(n772)
         );
  AOI21_X2 U3386 ( .B1(n19440), .B2(n3986), .A(n19439), .ZN(n20588) );
  NAND2_X1 U3388 ( .A1(n3116), .A2(n3072), .ZN(n9254) );
  AOI22_X1 U3391 ( .A1(n4513), .A2(n23645), .B1(n24320), .B2(n23652), .ZN(
        n22153) );
  NOR2_X1 U3396 ( .A1(n1201), .A2(n1200), .ZN(n4447) );
  NOR2_X1 U3397 ( .A1(n5472), .A2(n4923), .ZN(n898) );
  XNOR2_X1 U3398 ( .A(n15342), .B(n15238), .ZN(n15239) );
  NAND2_X1 U3401 ( .A1(n7431), .A2(n775), .ZN(n8339) );
  NAND2_X1 U3404 ( .A1(n7057), .A2(n9067), .ZN(n3249) );
  NAND3_X2 U3405 ( .A1(n3171), .A2(n2078), .A3(n6340), .ZN(n9067) );
  AOI21_X1 U3406 ( .B1(n777), .B2(n9560), .A(n9559), .ZN(n9561) );
  NAND2_X1 U3407 ( .A1(n1365), .A2(n16073), .ZN(n16074) );
  NAND2_X1 U3408 ( .A1(n778), .A2(n14178), .ZN(n4593) );
  NAND2_X1 U3409 ( .A1(n14181), .A2(n13796), .ZN(n778) );
  NAND4_X1 U3412 ( .A1(n23872), .A2(n3077), .A3(n3078), .A4(n23871), .ZN(
        n23874) );
  XNOR2_X1 U3413 ( .A(n781), .B(n21080), .ZN(n21082) );
  XNOR2_X1 U3414 ( .A(n21081), .B(n21429), .ZN(n781) );
  NAND2_X1 U3415 ( .A1(n7211), .A2(n7662), .ZN(n6548) );
  NAND2_X1 U3416 ( .A1(n9589), .A2(n9588), .ZN(n3551) );
  NAND2_X1 U3419 ( .A1(n14320), .A2(n13871), .ZN(n14459) );
  NAND2_X1 U3421 ( .A1(n22671), .A2(n22784), .ZN(n22672) );
  NAND3_X1 U3428 ( .A1(n23587), .A2(n23588), .A3(n23586), .ZN(n23590) );
  NAND2_X1 U3429 ( .A1(n10117), .A2(n784), .ZN(n9532) );
  NAND2_X1 U3430 ( .A1(n9530), .A2(n9531), .ZN(n784) );
  INV_X1 U3432 ( .A(n17734), .ZN(n4934) );
  NAND2_X1 U3433 ( .A1(n1086), .A2(n1087), .ZN(n12423) );
  NAND2_X1 U3434 ( .A1(n13177), .A2(n12506), .ZN(n13174) );
  OAI211_X2 U3435 ( .C1(n3656), .C2(n20165), .A(n19950), .B(n19949), .ZN(
        n21713) );
  OR2_X1 U3438 ( .A1(n10065), .A2(n10064), .ZN(n787) );
  OAI21_X1 U3439 ( .B1(n4083), .B2(n5158), .A(n4082), .ZN(n788) );
  NOR2_X2 U3440 ( .A1(n19020), .A2(n789), .ZN(n21639) );
  OAI22_X1 U3441 ( .A1(n20532), .A2(n20536), .B1(n19019), .B2(n20447), .ZN(
        n789) );
  XNOR2_X1 U3443 ( .A(n4687), .B(n4688), .ZN(n801) );
  NAND4_X1 U3444 ( .A1(n3425), .A2(n3426), .A3(n13964), .A4(n3427), .ZN(n790)
         );
  NAND3_X1 U3446 ( .A1(n6464), .A2(n6459), .A3(n6455), .ZN(n2078) );
  NAND2_X1 U3447 ( .A1(n3815), .A2(n16603), .ZN(n3816) );
  NAND2_X1 U3448 ( .A1(n2028), .A2(n2027), .ZN(n4511) );
  XNOR2_X1 U3450 ( .A(n792), .B(n23183), .ZN(Ciphertext[29]) );
  OAI22_X1 U3451 ( .A1(n23180), .A2(n23179), .B1(n23182), .B2(n23181), .ZN(
        n792) );
  NAND2_X1 U3452 ( .A1(n1145), .A2(n23688), .ZN(n1144) );
  INV_X1 U3453 ( .A(n933), .ZN(n7710) );
  NAND2_X1 U3454 ( .A1(n7865), .A2(n7862), .ZN(n933) );
  NAND3_X1 U3455 ( .A1(n10729), .A2(n10482), .A3(n10481), .ZN(n1178) );
  NAND3_X1 U3456 ( .A1(n6938), .A2(n6281), .A3(n793), .ZN(n5911) );
  OR2_X1 U3457 ( .A1(n6944), .A2(n5910), .ZN(n793) );
  NAND2_X1 U3458 ( .A1(n5910), .A2(n5887), .ZN(n6938) );
  XNOR2_X2 U3461 ( .A(n796), .B(n838), .ZN(n16274) );
  OR2_X1 U3462 ( .A1(n16334), .A2(n25092), .ZN(n981) );
  NAND2_X1 U3463 ( .A1(n14021), .A2(n14022), .ZN(n13540) );
  NAND2_X1 U3464 ( .A1(n22762), .A2(n23294), .ZN(n22761) );
  NAND2_X1 U3467 ( .A1(n4336), .A2(n13067), .ZN(n4340) );
  XNOR2_X1 U3471 ( .A(n17678), .B(n17679), .ZN(n797) );
  OAI21_X1 U3473 ( .B1(n8528), .B2(n269), .A(n799), .ZN(n798) );
  NAND2_X1 U3474 ( .A1(n7211), .A2(n8531), .ZN(n799) );
  NAND2_X1 U3476 ( .A1(n7933), .A2(n7932), .ZN(n2165) );
  NAND2_X1 U3477 ( .A1(n7163), .A2(n7923), .ZN(n7933) );
  NAND3_X2 U3478 ( .A1(n8352), .A2(n3708), .A3(n8351), .ZN(n8952) );
  AOI21_X1 U3480 ( .B1(n3764), .B2(n3765), .A(n16406), .ZN(n802) );
  NAND2_X1 U3481 ( .A1(n949), .A2(n6097), .ZN(n8005) );
  INV_X1 U3483 ( .A(n16997), .ZN(n17000) );
  NAND2_X1 U3484 ( .A1(n17574), .A2(n17368), .ZN(n16997) );
  XNOR2_X1 U3487 ( .A(n804), .B(n14470), .ZN(n14471) );
  XNOR2_X1 U3488 ( .A(n14469), .B(n14675), .ZN(n804) );
  INV_X1 U3490 ( .A(n7682), .ZN(n806) );
  NOR2_X1 U3495 ( .A1(n808), .A2(n19255), .ZN(n19073) );
  NAND2_X1 U3496 ( .A1(n21841), .A2(n22255), .ZN(n809) );
  AOI22_X2 U3497 ( .A1(n14007), .A2(n14006), .B1(n14005), .B2(n14004), .ZN(
        n14980) );
  NAND2_X1 U3500 ( .A1(n16902), .A2(n16539), .ZN(n17473) );
  NAND2_X1 U3501 ( .A1(n1116), .A2(n1118), .ZN(n5906) );
  NAND3_X1 U3502 ( .A1(n13462), .A2(n814), .A3(n813), .ZN(n14676) );
  NAND2_X1 U3503 ( .A1(n4921), .A2(n13959), .ZN(n814) );
  NAND2_X1 U3504 ( .A1(n17012), .A2(n4004), .ZN(n3516) );
  INV_X1 U3505 ( .A(n7920), .ZN(n1282) );
  NAND2_X1 U3507 ( .A1(n20912), .A2(n815), .ZN(n21736) );
  NAND3_X1 U3508 ( .A1(n817), .A2(n347), .A3(n816), .ZN(n815) );
  NAND2_X1 U3509 ( .A1(n20911), .A2(n346), .ZN(n816) );
  NAND2_X1 U3510 ( .A1(n20910), .A2(n20909), .ZN(n817) );
  NAND2_X1 U3511 ( .A1(n21888), .A2(n22265), .ZN(n22266) );
  NAND3_X1 U3513 ( .A1(n819), .A2(n4188), .A3(n4187), .ZN(Ciphertext[166]) );
  OAI21_X1 U3514 ( .B1(n4193), .B2(n4192), .A(n23868), .ZN(n819) );
  XNOR2_X1 U3515 ( .A(n820), .B(n19946), .ZN(n19966) );
  XNOR2_X1 U3516 ( .A(n19955), .B(n24899), .ZN(n820) );
  NOR2_X2 U3517 ( .A1(n1312), .A2(n20037), .ZN(n23857) );
  NAND2_X1 U3519 ( .A1(n14507), .A2(n24556), .ZN(n13977) );
  NAND2_X1 U3520 ( .A1(n9850), .A2(n9849), .ZN(n821) );
  NAND2_X1 U3521 ( .A1(n9384), .A2(n9592), .ZN(n822) );
  INV_X1 U3522 ( .A(n17486), .ZN(n17093) );
  NAND2_X1 U3524 ( .A1(n14327), .A2(n14328), .ZN(n14329) );
  NAND3_X1 U3525 ( .A1(n1589), .A2(n4235), .A3(n4237), .ZN(n4229) );
  NAND2_X1 U3526 ( .A1(n4230), .A2(n23200), .ZN(n1589) );
  INV_X1 U3528 ( .A(n2632), .ZN(n12829) );
  NAND2_X1 U3529 ( .A1(n13265), .A2(n2632), .ZN(n2631) );
  NAND2_X1 U3530 ( .A1(n4653), .A2(n17641), .ZN(n19917) );
  XNOR2_X1 U3531 ( .A(n823), .B(n18492), .ZN(n18494) );
  XNOR2_X1 U3532 ( .A(n18490), .B(n18491), .ZN(n823) );
  OAI211_X1 U3533 ( .C1(n22537), .C2(n23265), .A(n825), .B(n824), .ZN(n22538)
         );
  NAND2_X1 U3534 ( .A1(n22535), .A2(n23265), .ZN(n824) );
  NAND2_X1 U3535 ( .A1(n22536), .A2(n23281), .ZN(n825) );
  NAND2_X1 U3536 ( .A1(n829), .A2(n826), .ZN(n18251) );
  NAND2_X1 U3537 ( .A1(n828), .A2(n827), .ZN(n826) );
  INV_X1 U3538 ( .A(n17248), .ZN(n827) );
  AOI22_X1 U3539 ( .A1(n6558), .A2(n830), .B1(n6415), .B2(n6560), .ZN(n6417)
         );
  NAND2_X1 U3540 ( .A1(n6693), .A2(n6695), .ZN(n830) );
  XNOR2_X1 U3541 ( .A(n831), .B(n20505), .ZN(n20521) );
  XNOR2_X1 U3542 ( .A(n20504), .B(n21600), .ZN(n831) );
  NAND3_X1 U3543 ( .A1(n212), .A2(n4903), .A3(n832), .ZN(n2760) );
  NAND2_X1 U3544 ( .A1(n22530), .A2(n23860), .ZN(n832) );
  NAND2_X1 U3546 ( .A1(n22966), .A2(n24411), .ZN(n833) );
  OAI22_X1 U3547 ( .A1(n834), .A2(n14063), .B1(n13847), .B2(n13845), .ZN(
        n13849) );
  NOR2_X1 U3548 ( .A1(n13844), .A2(n13843), .ZN(n834) );
  AOI22_X2 U3549 ( .A1(n13310), .A2(n13309), .B1(n13312), .B2(n13311), .ZN(
        n13924) );
  NAND3_X1 U3552 ( .A1(n6051), .A2(n6746), .A3(n453), .ZN(n6747) );
  XNOR2_X2 U3553 ( .A(n5831), .B(Key[142]), .ZN(n6795) );
  NAND2_X1 U3554 ( .A1(n1774), .A2(n12665), .ZN(n1773) );
  NOR2_X2 U3555 ( .A1(n837), .A2(n19193), .ZN(n21514) );
  XNOR2_X1 U3557 ( .A(n14891), .B(n14893), .ZN(n838) );
  NAND3_X1 U3558 ( .A1(n22461), .A2(n22462), .A3(n3845), .ZN(n4339) );
  NAND3_X1 U3559 ( .A1(n13185), .A2(n24640), .A3(n12740), .ZN(n13105) );
  NAND2_X1 U3560 ( .A1(n5451), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U3561 ( .A1(n1599), .A2(n1793), .ZN(n20376) );
  NAND2_X1 U3562 ( .A1(n6776), .A2(n6292), .ZN(n6481) );
  AND2_X2 U3563 ( .A1(n10674), .A2(n1453), .ZN(n11163) );
  NOR2_X1 U3565 ( .A1(n1294), .A2(n1295), .ZN(n839) );
  NAND2_X1 U3566 ( .A1(n19686), .A2(n20149), .ZN(n19687) );
  NAND2_X1 U3567 ( .A1(n23690), .A2(n2305), .ZN(n22998) );
  NAND3_X2 U3569 ( .A1(n4619), .A2(n6316), .A3(n6317), .ZN(n7865) );
  OAI21_X1 U3570 ( .B1(n22109), .B2(n22929), .A(n22108), .ZN(n840) );
  NAND2_X1 U3571 ( .A1(n1530), .A2(n841), .ZN(n8088) );
  NAND2_X1 U3572 ( .A1(n3352), .A2(n842), .ZN(n841) );
  XNOR2_X1 U3573 ( .A(n843), .B(n23564), .ZN(Ciphertext[112]) );
  OAI211_X1 U3574 ( .C1(n23563), .C2(n23562), .A(n23560), .B(n23561), .ZN(n843) );
  NAND2_X1 U3576 ( .A1(n12633), .A2(n12206), .ZN(n5470) );
  OAI21_X2 U3580 ( .B1(n25036), .B2(n14083), .A(n12574), .ZN(n14857) );
  NAND3_X1 U3581 ( .A1(n13206), .A2(n1335), .A3(n13207), .ZN(n1725) );
  OAI22_X1 U3583 ( .A1(n845), .A2(n20186), .B1(n20043), .B2(n20191), .ZN(
        n20044) );
  NAND2_X1 U3584 ( .A1(n20041), .A2(n20042), .ZN(n845) );
  NAND2_X1 U3585 ( .A1(n2346), .A2(n19592), .ZN(n19589) );
  NAND2_X1 U3588 ( .A1(n9929), .A2(n9934), .ZN(n847) );
  NAND2_X1 U3589 ( .A1(n7838), .A2(n25217), .ZN(n848) );
  NAND2_X1 U3592 ( .A1(n16250), .A2(n16018), .ZN(n849) );
  NOR2_X1 U3595 ( .A1(n22533), .A2(n852), .ZN(n22534) );
  AOI21_X1 U3596 ( .B1(n18718), .B2(n19497), .A(n19499), .ZN(n18723) );
  XNOR2_X1 U3597 ( .A(n854), .B(n20812), .ZN(n20814) );
  XNOR2_X1 U3598 ( .A(n20811), .B(n24896), .ZN(n854) );
  NAND2_X1 U3601 ( .A1(n14010), .A2(n14254), .ZN(n855) );
  NAND2_X1 U3602 ( .A1(n14255), .A2(n14252), .ZN(n856) );
  NAND2_X1 U3606 ( .A1(n10219), .A2(n857), .ZN(n11616) );
  NAND2_X1 U3607 ( .A1(n10220), .A2(n10782), .ZN(n857) );
  INV_X1 U3609 ( .A(n8697), .ZN(n5553) );
  XNOR2_X1 U3610 ( .A(n9106), .B(n8959), .ZN(n8697) );
  XNOR2_X1 U3611 ( .A(n11943), .B(n11944), .ZN(n3473) );
  NAND3_X1 U3614 ( .A1(n5187), .A2(n5188), .A3(n20255), .ZN(n5186) );
  NAND3_X1 U3617 ( .A1(n5366), .A2(n281), .A3(n5367), .ZN(n5599) );
  NAND3_X1 U3619 ( .A1(n22506), .A2(n23443), .A3(n321), .ZN(n23444) );
  OAI211_X1 U3621 ( .C1(n1175), .C2(n6776), .A(n6290), .B(n6775), .ZN(n6199)
         );
  OAI21_X1 U3622 ( .B1(n20226), .B2(n3016), .A(n862), .ZN(n20271) );
  NAND2_X1 U3623 ( .A1(n3016), .A2(n20268), .ZN(n862) );
  NAND2_X1 U3624 ( .A1(n6894), .A2(n313), .ZN(n2914) );
  OAI21_X1 U3625 ( .B1(n13013), .B2(n13245), .A(n863), .ZN(n12563) );
  NAND2_X1 U3626 ( .A1(n13245), .A2(n25199), .ZN(n863) );
  OR2_X1 U3627 ( .A1(n19786), .A2(n19987), .ZN(n19753) );
  NOR2_X1 U3628 ( .A1(n21382), .A2(n22323), .ZN(n22322) );
  OR2_X1 U3629 ( .A1(n13132), .A2(n25033), .ZN(n1844) );
  OAI21_X1 U3630 ( .B1(n10570), .B2(n416), .A(n864), .ZN(n10576) );
  NAND2_X1 U3631 ( .A1(n10570), .A2(n10571), .ZN(n864) );
  XNOR2_X2 U3632 ( .A(n1884), .B(n14404), .ZN(n16170) );
  INV_X1 U3633 ( .A(n21909), .ZN(n22275) );
  NAND2_X1 U3634 ( .A1(n21910), .A2(n22138), .ZN(n21909) );
  INV_X1 U3635 ( .A(n1095), .ZN(n15709) );
  XNOR2_X1 U3637 ( .A(n868), .B(n14414), .ZN(n14422) );
  XNOR2_X1 U3638 ( .A(n14960), .B(n14413), .ZN(n868) );
  NAND3_X1 U3639 ( .A1(n6338), .A2(n6510), .A3(n6337), .ZN(n3171) );
  NAND2_X1 U3641 ( .A1(n4499), .A2(n13298), .ZN(n1818) );
  NAND2_X1 U3642 ( .A1(n3557), .A2(n13200), .ZN(n870) );
  NAND2_X1 U3643 ( .A1(n22952), .A2(n871), .ZN(n1889) );
  NOR2_X1 U3644 ( .A1(n24884), .A2(n22954), .ZN(n871) );
  NAND2_X1 U3646 ( .A1(n6359), .A2(n6360), .ZN(n873) );
  NAND2_X1 U3647 ( .A1(n25041), .A2(n22836), .ZN(n22895) );
  NAND2_X2 U3649 ( .A1(n874), .A2(n4796), .ZN(n13868) );
  NAND2_X1 U3650 ( .A1(n4333), .A2(n4332), .ZN(n874) );
  NOR2_X1 U3651 ( .A1(n5481), .A2(n19532), .ZN(n5475) );
  AOI21_X1 U3652 ( .B1(n17388), .B2(n17387), .A(n875), .ZN(n17393) );
  AOI22_X1 U3654 ( .A1(n877), .A2(n23531), .B1(n23008), .B2(n23505), .ZN(
        n22930) );
  NAND2_X1 U3655 ( .A1(n23013), .A2(n24313), .ZN(n877) );
  NAND2_X1 U3656 ( .A1(n21356), .A2(n23828), .ZN(n21357) );
  NAND2_X1 U3657 ( .A1(n8528), .A2(n269), .ZN(n4994) );
  NAND3_X1 U3660 ( .A1(n24589), .A2(n13646), .A3(n13824), .ZN(n13650) );
  NAND2_X1 U3662 ( .A1(n16509), .A2(n15605), .ZN(n880) );
  NAND2_X1 U3664 ( .A1(n9601), .A2(n9602), .ZN(n9607) );
  NAND2_X1 U3665 ( .A1(n6916), .A2(n6912), .ZN(n5845) );
  AND3_X1 U3666 ( .A1(n3350), .A2(n13991), .A3(n3349), .ZN(n1112) );
  INV_X1 U3667 ( .A(n17122), .ZN(n2580) );
  OAI211_X1 U3668 ( .C1(n10414), .C2(n10617), .A(n10413), .B(n977), .ZN(n11237) );
  NAND2_X1 U3669 ( .A1(n882), .A2(n1975), .ZN(n8026) );
  NAND2_X1 U3670 ( .A1(n1840), .A2(n8023), .ZN(n882) );
  NAND2_X1 U3671 ( .A1(n7882), .A2(n7883), .ZN(n7885) );
  OR2_X2 U3672 ( .A1(n5850), .A2(n5849), .ZN(n7883) );
  NAND2_X1 U3674 ( .A1(n19515), .A2(n19984), .ZN(n883) );
  NAND2_X1 U3675 ( .A1(n19516), .A2(n885), .ZN(n884) );
  XNOR2_X1 U3677 ( .A(n1111), .B(n1359), .ZN(n14370) );
  NAND2_X1 U3678 ( .A1(n7322), .A2(n7323), .ZN(n2733) );
  AND2_X2 U3679 ( .A1(n6009), .A2(n6008), .ZN(n7322) );
  XNOR2_X2 U3680 ( .A(Key[74]), .B(Plaintext[74]), .ZN(n5774) );
  AND2_X1 U3681 ( .A1(n16572), .A2(n890), .ZN(n16802) );
  INV_X1 U3682 ( .A(n17122), .ZN(n890) );
  NAND2_X1 U3685 ( .A1(n2753), .A2(n22240), .ZN(n22062) );
  NAND2_X1 U3686 ( .A1(n1243), .A2(n1246), .ZN(n892) );
  NAND2_X1 U3687 ( .A1(n24480), .A2(n11143), .ZN(n10304) );
  NAND2_X1 U3691 ( .A1(n13322), .A2(n13318), .ZN(n893) );
  OAI21_X1 U3692 ( .B1(n11525), .B2(n895), .A(n894), .ZN(n10581) );
  NAND2_X1 U3693 ( .A1(n11525), .A2(n25060), .ZN(n894) );
  AOI22_X1 U3694 ( .A1(n17454), .A2(n17455), .B1(n17456), .B2(n17457), .ZN(
        n17458) );
  OAI21_X1 U3696 ( .B1(n6371), .B2(n6658), .A(n6370), .ZN(n897) );
  NAND2_X1 U3698 ( .A1(n19821), .A2(n19788), .ZN(n19819) );
  NAND2_X1 U3699 ( .A1(n1680), .A2(n2853), .ZN(n23579) );
  OR2_X1 U3700 ( .A1(n25401), .A2(n6488), .ZN(n5953) );
  NOR2_X1 U3701 ( .A1(n1127), .A2(n898), .ZN(n14308) );
  NOR2_X1 U3702 ( .A1(n900), .A2(n10788), .ZN(n4051) );
  NOR2_X1 U3703 ( .A1(n1824), .A2(n10793), .ZN(n900) );
  XNOR2_X2 U3704 ( .A(n5817), .B(Key[126]), .ZN(n6367) );
  OAI21_X1 U3706 ( .B1(n16475), .B2(n16474), .A(n901), .ZN(n15460) );
  NAND2_X1 U3707 ( .A1(n16475), .A2(n15546), .ZN(n901) );
  XNOR2_X1 U3708 ( .A(n18308), .B(n934), .ZN(n17926) );
  NAND2_X1 U3709 ( .A1(n11438), .A2(n25337), .ZN(n902) );
  NAND2_X1 U3710 ( .A1(n20560), .A2(n20094), .ZN(n19727) );
  AOI21_X2 U3711 ( .B1(n19726), .B2(n19719), .A(n19725), .ZN(n20560) );
  XNOR2_X1 U3712 ( .A(n903), .B(n21696), .ZN(n21698) );
  XNOR2_X1 U3713 ( .A(n21695), .B(n21694), .ZN(n903) );
  NAND3_X1 U3714 ( .A1(n14416), .A2(n14278), .A3(n24958), .ZN(n13444) );
  NAND3_X1 U3715 ( .A1(n2514), .A2(n14946), .A3(n13801), .ZN(n13802) );
  NAND2_X1 U3716 ( .A1(n906), .A2(n23411), .ZN(n905) );
  INV_X1 U3717 ( .A(n23410), .ZN(n906) );
  NAND2_X1 U3718 ( .A1(n23418), .A2(n24947), .ZN(n907) );
  NAND3_X1 U3719 ( .A1(n3544), .A2(n16406), .A3(n24062), .ZN(n5212) );
  NAND2_X1 U3720 ( .A1(n6488), .A2(n6781), .ZN(n908) );
  NAND2_X1 U3721 ( .A1(n6305), .A2(n6304), .ZN(n909) );
  NAND2_X1 U3722 ( .A1(n910), .A2(n24007), .ZN(n3485) );
  NAND2_X1 U3723 ( .A1(n3486), .A2(n24005), .ZN(n910) );
  XNOR2_X1 U3724 ( .A(n911), .B(n14903), .ZN(n14906) );
  XNOR2_X1 U3725 ( .A(n14901), .B(n15112), .ZN(n911) );
  NAND3_X1 U3728 ( .A1(n914), .A2(n5029), .A3(n5032), .ZN(Ciphertext[14]) );
  NAND2_X1 U3729 ( .A1(n5028), .A2(n5031), .ZN(n914) );
  NAND2_X1 U3730 ( .A1(n915), .A2(n13988), .ZN(n13990) );
  INV_X1 U3731 ( .A(n13987), .ZN(n915) );
  NAND2_X1 U3732 ( .A1(n5416), .A2(n13247), .ZN(n13987) );
  NAND2_X1 U3733 ( .A1(n7328), .A2(n7897), .ZN(n7332) );
  NAND2_X1 U3734 ( .A1(n24952), .A2(n23112), .ZN(n5035) );
  XNOR2_X1 U3735 ( .A(n916), .B(n449), .ZN(Ciphertext[180]) );
  NAND2_X1 U3736 ( .A1(n23950), .A2(n23951), .ZN(n916) );
  OR2_X1 U3737 ( .A1(n6987), .A2(n6244), .ZN(n6247) );
  OAI211_X2 U3740 ( .C1(n5595), .C2(n7187), .A(n918), .B(n7645), .ZN(n8909) );
  NAND2_X1 U3741 ( .A1(n5593), .A2(n5595), .ZN(n918) );
  AOI21_X1 U3742 ( .B1(n22468), .B2(n22675), .A(n919), .ZN(n22470) );
  NAND2_X1 U3743 ( .A1(n7918), .A2(n435), .ZN(n920) );
  OR3_X1 U3744 ( .A1(n20290), .A2(n21008), .A3(n20523), .ZN(n2852) );
  NAND3_X2 U3746 ( .A1(n21933), .A2(n21932), .A3(n21931), .ZN(n23201) );
  NAND2_X1 U3747 ( .A1(n1299), .A2(n18914), .ZN(n18916) );
  OR2_X1 U3748 ( .A1(n19185), .A2(n19548), .ZN(n1710) );
  OR2_X1 U3750 ( .A1(n3822), .A2(n17613), .ZN(n16562) );
  NAND2_X1 U3751 ( .A1(n17408), .A2(n16561), .ZN(n3822) );
  NAND4_X2 U3752 ( .A1(n5984), .A2(n5985), .A3(n5983), .A4(n5982), .ZN(n7604)
         );
  AND2_X1 U3753 ( .A1(n17173), .A2(n927), .ZN(n16435) );
  NAND2_X1 U3754 ( .A1(n17175), .A2(n16434), .ZN(n927) );
  AOI21_X1 U3755 ( .B1(n17174), .B2(n282), .A(n17175), .ZN(n4413) );
  NAND2_X1 U3756 ( .A1(n22961), .A2(n24343), .ZN(n932) );
  XNOR2_X1 U3757 ( .A(n928), .B(n931), .ZN(Ciphertext[69]) );
  NAND3_X1 U3758 ( .A1(n929), .A2(n3014), .A3(n22995), .ZN(n928) );
  NAND3_X1 U3759 ( .A1(n930), .A2(n932), .A3(n23340), .ZN(n929) );
  OR2_X1 U3760 ( .A1(n23354), .A2(n23349), .ZN(n930) );
  INV_X1 U3761 ( .A(n932), .ZN(n22996) );
  AOI21_X1 U3762 ( .B1(n933), .B2(n7868), .A(n3570), .ZN(n7711) );
  XNOR2_X1 U3763 ( .A(n18310), .B(n934), .ZN(n16000) );
  XNOR2_X1 U3764 ( .A(n934), .B(n1777), .ZN(n17883) );
  XNOR2_X1 U3765 ( .A(n18285), .B(n934), .ZN(n18286) );
  NAND2_X1 U3766 ( .A1(n936), .A2(n24585), .ZN(n17056) );
  INV_X1 U3767 ( .A(n16932), .ZN(n936) );
  NOR2_X1 U3768 ( .A1(n24398), .A2(n16932), .ZN(n16610) );
  NAND2_X1 U3769 ( .A1(n23350), .A2(n23349), .ZN(n938) );
  NAND2_X1 U3770 ( .A1(n937), .A2(n23350), .ZN(n3014) );
  OAI21_X1 U3771 ( .B1(n24343), .B2(n24400), .A(n938), .ZN(n23037) );
  AOI22_X1 U3772 ( .A1(n22979), .A2(n22996), .B1(n23363), .B2(n938), .ZN(
        n22980) );
  NAND2_X1 U3774 ( .A1(n24753), .A2(n939), .ZN(n11096) );
  XNOR2_X1 U3776 ( .A(n13642), .B(n13641), .ZN(n940) );
  NAND2_X1 U3777 ( .A1(n24960), .A2(n25500), .ZN(n15811) );
  OAI21_X1 U3778 ( .B1(n3544), .B2(n24960), .A(n15646), .ZN(n16199) );
  NAND2_X1 U3779 ( .A1(n941), .A2(n7382), .ZN(n7303) );
  NAND3_X1 U3780 ( .A1(n7386), .A2(n7618), .A3(n941), .ZN(n7203) );
  NAND2_X1 U3781 ( .A1(n7383), .A2(n941), .ZN(n7389) );
  AOI21_X1 U3782 ( .B1(n7616), .B2(n941), .A(n7615), .ZN(n7624) );
  INV_X1 U3783 ( .A(n6156), .ZN(n943) );
  NAND2_X1 U3784 ( .A1(n8005), .A2(n7754), .ZN(n8003) );
  NAND3_X1 U3785 ( .A1(n945), .A2(n6074), .A3(n6073), .ZN(n7754) );
  NAND2_X1 U3786 ( .A1(n6657), .A2(n946), .ZN(n945) );
  NAND2_X1 U3787 ( .A1(n6658), .A2(n947), .ZN(n946) );
  NAND2_X1 U3788 ( .A1(n950), .A2(n448), .ZN(n949) );
  NAND2_X1 U3789 ( .A1(n6834), .A2(n7009), .ZN(n950) );
  NAND3_X1 U3792 ( .A1(n18967), .A2(n19300), .A3(n3653), .ZN(n951) );
  INV_X1 U3793 ( .A(n19297), .ZN(n3653) );
  NAND3_X1 U3794 ( .A1(n18856), .A2(n18970), .A3(n18928), .ZN(n952) );
  NAND2_X1 U3796 ( .A1(n9475), .A2(n9476), .ZN(n953) );
  AOI21_X1 U3797 ( .B1(n9473), .B2(n9864), .A(n9860), .ZN(n954) );
  AND2_X1 U3798 ( .A1(n10886), .A2(n10887), .ZN(n9477) );
  NAND2_X1 U3799 ( .A1(n9456), .A2(n956), .ZN(n955) );
  NAND2_X1 U3800 ( .A1(n961), .A2(n959), .ZN(n958) );
  NAND3_X1 U3801 ( .A1(n362), .A2(n19192), .A3(n960), .ZN(n959) );
  NAND2_X1 U3802 ( .A1(n19571), .A2(n19570), .ZN(n961) );
  AOI21_X1 U3803 ( .B1(n19567), .B2(n19566), .A(n19565), .ZN(n962) );
  NAND3_X1 U3804 ( .A1(n17230), .A2(n2285), .A3(n16951), .ZN(n14589) );
  NAND3_X1 U3805 ( .A1(n1656), .A2(n1655), .A3(n24537), .ZN(n963) );
  OAI21_X1 U3806 ( .B1(n16917), .B2(n17335), .A(n16915), .ZN(n16919) );
  XNOR2_X1 U3809 ( .A(n966), .B(n18436), .ZN(n18441) );
  INV_X1 U3810 ( .A(n966), .ZN(n4808) );
  INV_X1 U3811 ( .A(n17874), .ZN(n4942) );
  NAND2_X1 U3812 ( .A1(n967), .A2(n4356), .ZN(n4355) );
  NAND3_X1 U3813 ( .A1(n967), .A2(n14159), .A3(n5080), .ZN(n3085) );
  AOI22_X2 U3814 ( .A1(n1235), .A2(n15868), .B1(n15867), .B2(n16141), .ZN(
        n17119) );
  AND2_X2 U3815 ( .A1(n969), .A2(n968), .ZN(n17120) );
  NAND2_X1 U3816 ( .A1(n15855), .A2(n24928), .ZN(n968) );
  NAND3_X1 U3818 ( .A1(n23828), .A2(n23827), .A3(n318), .ZN(n21349) );
  AND2_X1 U3819 ( .A1(n4219), .A2(n1099), .ZN(n971) );
  NAND2_X1 U3820 ( .A1(n303), .A2(n12795), .ZN(n973) );
  OAI21_X1 U3822 ( .B1(n12799), .B2(n12798), .A(n12797), .ZN(n974) );
  INV_X1 U3823 ( .A(n1646), .ZN(n975) );
  AOI21_X2 U3824 ( .B1(n976), .B2(n12802), .A(n12801), .ZN(n14328) );
  NAND2_X1 U3826 ( .A1(n978), .A2(n10611), .ZN(n977) );
  NAND2_X1 U3827 ( .A1(n10614), .A2(n10486), .ZN(n10611) );
  NAND2_X1 U3828 ( .A1(n979), .A2(n980), .ZN(n978) );
  NAND2_X1 U3829 ( .A1(n10412), .A2(n10411), .ZN(n979) );
  NAND2_X1 U3830 ( .A1(n10486), .A2(n10411), .ZN(n980) );
  OAI211_X1 U3831 ( .C1(n388), .C2(n16334), .A(n981), .B(n15755), .ZN(n5317)
         );
  NAND2_X1 U3833 ( .A1(n21031), .A2(n21038), .ZN(n2248) );
  OR2_X1 U3835 ( .A1(n298), .A2(n13863), .ZN(n984) );
  NAND2_X1 U3836 ( .A1(n986), .A2(n16342), .ZN(n17620) );
  NAND2_X1 U3837 ( .A1(n987), .A2(n4926), .ZN(n986) );
  NOR2_X1 U3839 ( .A1(n19575), .A2(n988), .ZN(n1098) );
  MUX2_X1 U3840 ( .A(n988), .B(n24982), .S(n19575), .Z(n1004) );
  NAND2_X1 U3841 ( .A1(n7390), .A2(n7647), .ZN(n7649) );
  INV_X1 U3842 ( .A(n7646), .ZN(n7390) );
  AND2_X1 U3843 ( .A1(n12817), .A2(n14088), .ZN(n990) );
  NAND2_X1 U3844 ( .A1(n4510), .A2(n14085), .ZN(n12817) );
  NAND2_X1 U3845 ( .A1(n13537), .A2(n13536), .ZN(n14085) );
  NAND2_X1 U3848 ( .A1(n15757), .A2(n16001), .ZN(n995) );
  XNOR2_X2 U3849 ( .A(n15144), .B(n15145), .ZN(n16266) );
  AOI21_X1 U3852 ( .B1(n3856), .B2(n22253), .A(n332), .ZN(n996) );
  AOI21_X1 U3854 ( .B1(n22254), .B2(n24468), .A(n24362), .ZN(n998) );
  NAND2_X1 U3856 ( .A1(n20354), .A2(n20352), .ZN(n999) );
  NAND2_X1 U3857 ( .A1(n20003), .A2(n20479), .ZN(n20352) );
  INV_X1 U3858 ( .A(n19057), .ZN(n19060) );
  INV_X1 U3859 ( .A(n19578), .ZN(n1002) );
  NAND2_X1 U3861 ( .A1(n1005), .A2(n1004), .ZN(n1003) );
  AND2_X1 U3862 ( .A1(n23645), .A2(n23640), .ZN(n23653) );
  OAI211_X1 U3863 ( .C1(n22116), .C2(n22072), .A(n22169), .B(n22115), .ZN(
        n1006) );
  OAI211_X1 U3864 ( .C1(n20353), .C2(n20480), .A(n1008), .B(n20003), .ZN(n1992) );
  NAND4_X2 U3866 ( .A1(n4717), .A2(n4716), .A3(n3388), .A4(n3389), .ZN(n20479)
         );
  INV_X1 U3867 ( .A(n20479), .ZN(n2168) );
  INV_X1 U3868 ( .A(n1012), .ZN(n1011) );
  INV_X1 U3869 ( .A(n19269), .ZN(n1013) );
  NAND3_X1 U3870 ( .A1(n1019), .A2(n12991), .A3(n1018), .ZN(n1017) );
  NAND2_X1 U3871 ( .A1(n2608), .A2(n1020), .ZN(n1019) );
  NAND2_X1 U3873 ( .A1(n9872), .A2(n1021), .ZN(n9879) );
  NAND3_X1 U3874 ( .A1(n4993), .A2(n2294), .A3(n1021), .ZN(n9032) );
  MUX2_X1 U3875 ( .A(n9872), .B(n24549), .S(n9027), .Z(n9549) );
  INV_X1 U3877 ( .A(n20003), .ZN(n20477) );
  NOR2_X1 U3878 ( .A1(n20003), .A2(n20479), .ZN(n1024) );
  NAND2_X1 U3880 ( .A1(n1028), .A2(n1027), .ZN(n1026) );
  AND2_X1 U3882 ( .A1(n18834), .A2(n24478), .ZN(n2695) );
  NAND2_X1 U3883 ( .A1(n19438), .A2(n24478), .ZN(n18835) );
  NAND2_X1 U3884 ( .A1(n18642), .A2(n1029), .ZN(n18643) );
  AND2_X1 U3885 ( .A1(n24478), .A2(n25422), .ZN(n1029) );
  INV_X1 U3887 ( .A(n18651), .ZN(n1030) );
  NAND2_X1 U3888 ( .A1(n19081), .A2(n24478), .ZN(n18651) );
  NAND2_X1 U3891 ( .A1(n17629), .A2(n16539), .ZN(n1032) );
  INV_X1 U3892 ( .A(n2566), .ZN(n1033) );
  XNOR2_X1 U3893 ( .A(n18633), .B(n5120), .ZN(n18634) );
  NAND3_X1 U3895 ( .A1(n17629), .A2(n2561), .A3(n17633), .ZN(n1036) );
  NAND2_X1 U3896 ( .A1(n1038), .A2(n434), .ZN(n1037) );
  NAND2_X1 U3897 ( .A1(n1039), .A2(n7078), .ZN(n1038) );
  NAND2_X1 U3898 ( .A1(n7674), .A2(n25251), .ZN(n1039) );
  NAND2_X1 U3899 ( .A1(n1041), .A2(n6869), .ZN(n1040) );
  NAND2_X1 U3900 ( .A1(n7506), .A2(n1379), .ZN(n6869) );
  NAND2_X1 U3901 ( .A1(n7510), .A2(n7509), .ZN(n1041) );
  NAND2_X1 U3902 ( .A1(n1162), .A2(n7224), .ZN(n7509) );
  OR2_X2 U3903 ( .A1(n6868), .A2(n6867), .ZN(n7224) );
  NAND2_X1 U3904 ( .A1(n7078), .A2(n7674), .ZN(n7510) );
  NAND2_X1 U3905 ( .A1(n3274), .A2(n3273), .ZN(n7078) );
  NAND2_X1 U3906 ( .A1(n1043), .A2(n1042), .ZN(n1045) );
  NAND2_X1 U3907 ( .A1(n297), .A2(n14153), .ZN(n1042) );
  NAND2_X1 U3908 ( .A1(n14154), .A2(n13805), .ZN(n1043) );
  NAND3_X2 U3909 ( .A1(n1045), .A2(n14152), .A3(n1044), .ZN(n15055) );
  NAND2_X1 U3910 ( .A1(n14151), .A2(n14150), .ZN(n1044) );
  NAND2_X1 U3911 ( .A1(n1049), .A2(n19568), .ZN(n1048) );
  INV_X1 U3912 ( .A(n19191), .ZN(n5634) );
  XNOR2_X2 U3913 ( .A(n18307), .B(n18306), .ZN(n19191) );
  NAND2_X1 U3914 ( .A1(n19568), .A2(n1053), .ZN(n1052) );
  INV_X1 U3915 ( .A(n11297), .ZN(n11091) );
  NAND2_X1 U3916 ( .A1(n9528), .A2(n2855), .ZN(n11297) );
  NAND2_X1 U3918 ( .A1(n1055), .A2(n11302), .ZN(n1054) );
  INV_X1 U3919 ( .A(n11297), .ZN(n1055) );
  NAND2_X1 U3920 ( .A1(n10762), .A2(n11298), .ZN(n1057) );
  AOI22_X2 U3921 ( .A1(n10896), .A2(n1059), .B1(n10898), .B2(n10897), .ZN(
        n11627) );
  INV_X1 U3922 ( .A(n1055), .ZN(n1059) );
  NAND2_X1 U3923 ( .A1(n391), .A2(n11454), .ZN(n2301) );
  NAND2_X1 U3924 ( .A1(n14088), .A2(n4510), .ZN(n1062) );
  INV_X1 U3925 ( .A(n25372), .ZN(n21648) );
  XNOR2_X1 U3926 ( .A(n21650), .B(n1063), .ZN(n21651) );
  XNOR2_X1 U3927 ( .A(n25372), .B(n24319), .ZN(n1063) );
  OAI22_X1 U3929 ( .A1(n22941), .A2(n337), .B1(n22832), .B2(n22940), .ZN(n1066) );
  NAND2_X1 U3931 ( .A1(n25063), .A2(n1066), .ZN(n1065) );
  NAND2_X1 U3932 ( .A1(n22830), .A2(n22832), .ZN(n1068) );
  NOR2_X1 U3933 ( .A1(n23398), .A2(n23420), .ZN(n22868) );
  NAND2_X1 U3934 ( .A1(n13097), .A2(n1069), .ZN(n1080) );
  NAND2_X1 U3936 ( .A1(n13094), .A2(n3492), .ZN(n1069) );
  NAND3_X1 U3937 ( .A1(n16612), .A2(n16730), .A3(n283), .ZN(n1070) );
  NAND2_X1 U3938 ( .A1(n5761), .A2(n1071), .ZN(n16613) );
  NAND2_X1 U3939 ( .A1(n1073), .A2(n1072), .ZN(n20053) );
  NAND2_X1 U3940 ( .A1(n20480), .A2(n20476), .ZN(n20051) );
  NAND2_X1 U3941 ( .A1(n20048), .A2(n2168), .ZN(n1073) );
  NAND2_X1 U3942 ( .A1(n1075), .A2(n23311), .ZN(n5660) );
  NAND2_X1 U3943 ( .A1(n5662), .A2(n5664), .ZN(n1074) );
  OAI22_X1 U3946 ( .A1(n21891), .A2(n24881), .B1(n4109), .B2(n22974), .ZN(
        n1076) );
  NOR2_X1 U3947 ( .A1(n7590), .A2(n7591), .ZN(n1194) );
  OAI21_X2 U3948 ( .B1(n5452), .B2(n1079), .A(n1077), .ZN(n7591) );
  NAND2_X1 U3949 ( .A1(n1078), .A2(n1698), .ZN(n1077) );
  NAND2_X1 U3950 ( .A1(n6315), .A2(n6467), .ZN(n6328) );
  NAND3_X1 U3951 ( .A1(n13119), .A2(n13113), .A3(n12503), .ZN(n1082) );
  NAND2_X1 U3952 ( .A1(n7508), .A2(n1083), .ZN(n2263) );
  NAND2_X1 U3953 ( .A1(n1084), .A2(n7506), .ZN(n1083) );
  INV_X1 U3954 ( .A(n13900), .ZN(n13958) );
  NAND2_X1 U3955 ( .A1(n12659), .A2(n12503), .ZN(n1087) );
  NAND2_X1 U3956 ( .A1(n12291), .A2(n3328), .ZN(n1086) );
  NAND2_X1 U3957 ( .A1(n13958), .A2(n13903), .ZN(n13459) );
  AOI21_X1 U3958 ( .B1(n7262), .B2(n1088), .A(n7261), .ZN(n7265) );
  XNOR2_X1 U3959 ( .A(n1089), .B(n8263), .ZN(n8267) );
  INV_X1 U3960 ( .A(n8851), .ZN(n1089) );
  XNOR2_X1 U3961 ( .A(n1090), .B(n8851), .ZN(n8838) );
  INV_X1 U3962 ( .A(n8835), .ZN(n1090) );
  XNOR2_X1 U3963 ( .A(n1091), .B(n15338), .ZN(n14652) );
  XNOR2_X1 U3964 ( .A(n1091), .B(n15485), .ZN(n15492) );
  XNOR2_X1 U3965 ( .A(n1091), .B(n15239), .ZN(n15243) );
  OAI21_X1 U3968 ( .B1(n9953), .B2(n9955), .A(n9949), .ZN(n1093) );
  NAND2_X1 U3970 ( .A1(n16439), .A2(n1095), .ZN(n16446) );
  OAI22_X1 U3971 ( .A1(n1097), .A2(n16492), .B1(n16490), .B2(n387), .ZN(n1096)
         );
  NAND3_X1 U3973 ( .A1(n21839), .A2(n22361), .A3(n245), .ZN(n1099) );
  NAND2_X1 U3974 ( .A1(n24608), .A2(n22356), .ZN(n1100) );
  NAND2_X1 U3977 ( .A1(n6189), .A2(n1106), .ZN(n4881) );
  NAND2_X1 U3978 ( .A1(n6195), .A2(n6445), .ZN(n6453) );
  NAND2_X1 U3979 ( .A1(n19315), .A2(n19312), .ZN(n1107) );
  NAND2_X1 U3980 ( .A1(n17563), .A2(n1107), .ZN(n17565) );
  NOR2_X1 U3981 ( .A1(n1109), .A2(n19984), .ZN(n1108) );
  NOR2_X2 U3982 ( .A1(n1159), .A2(n18926), .ZN(n19984) );
  INV_X1 U3983 ( .A(n24464), .ZN(n1109) );
  XNOR2_X1 U3984 ( .A(n1110), .B(n8615), .ZN(n8071) );
  XNOR2_X1 U3985 ( .A(n9034), .B(n1110), .ZN(n9037) );
  XNOR2_X1 U3986 ( .A(n8491), .B(n1110), .ZN(n7980) );
  XNOR2_X1 U3987 ( .A(n8537), .B(n1110), .ZN(n7594) );
  NAND2_X1 U3988 ( .A1(n16474), .A2(n16473), .ZN(n15688) );
  NAND3_X1 U3989 ( .A1(n16469), .A2(n15546), .A3(n16471), .ZN(n1113) );
  NAND3_X1 U3990 ( .A1(n16472), .A2(n16473), .A3(n16474), .ZN(n1114) );
  MUX2_X1 U3991 ( .A(n16578), .B(n17086), .S(n16649), .Z(n15875) );
  NAND2_X1 U3992 ( .A1(n15795), .A2(n16069), .ZN(n1115) );
  NAND2_X1 U3994 ( .A1(n1119), .A2(n6255), .ZN(n1116) );
  NAND2_X1 U3995 ( .A1(n5905), .A2(n25437), .ZN(n1118) );
  AOI21_X1 U3996 ( .B1(n6254), .B2(n1119), .A(n6528), .ZN(n6258) );
  NAND2_X1 U3997 ( .A1(n6948), .A2(n6529), .ZN(n1119) );
  OAI22_X1 U3998 ( .A1(n19565), .A2(n19273), .B1(n19192), .B2(n19570), .ZN(
        n19274) );
  XNOR2_X2 U3999 ( .A(n18330), .B(n18329), .ZN(n19570) );
  NAND2_X1 U4000 ( .A1(n19274), .A2(n18907), .ZN(n1120) );
  NAND2_X1 U4001 ( .A1(n363), .A2(n19570), .ZN(n18907) );
  NAND2_X1 U4002 ( .A1(n18794), .A2(n18793), .ZN(n1121) );
  INV_X1 U4004 ( .A(n15667), .ZN(n1123) );
  NOR2_X1 U4005 ( .A1(n3947), .A2(n25092), .ZN(n16335) );
  AND2_X1 U4006 ( .A1(n267), .A2(n16332), .ZN(n16339) );
  OAI21_X2 U4008 ( .B1(n12426), .B2(n13150), .A(n1125), .ZN(n14307) );
  NAND2_X1 U4009 ( .A1(n1126), .A2(n13129), .ZN(n1125) );
  OAI21_X1 U4010 ( .B1(n13148), .B2(n13130), .A(n13131), .ZN(n1126) );
  NAND3_X1 U4011 ( .A1(n1128), .A2(n7139), .A3(n7896), .ZN(n7143) );
  NAND2_X1 U4012 ( .A1(n1130), .A2(n3469), .ZN(n1128) );
  INV_X1 U4013 ( .A(n3469), .ZN(n7902) );
  NAND2_X2 U4014 ( .A1(n1129), .A2(n1398), .ZN(n3469) );
  NAND2_X1 U4015 ( .A1(n5876), .A2(n5875), .ZN(n1129) );
  INV_X1 U4016 ( .A(n7327), .ZN(n1130) );
  NAND3_X1 U4018 ( .A1(n1138), .A2(n17067), .A3(n17066), .ZN(n1133) );
  NAND2_X1 U4019 ( .A1(n17069), .A2(n1139), .ZN(n16734) );
  NAND3_X1 U4020 ( .A1(n15609), .A2(n1136), .A3(n1134), .ZN(n18262) );
  NAND2_X1 U4021 ( .A1(n1135), .A2(n283), .ZN(n1134) );
  NAND2_X1 U4022 ( .A1(n16730), .A2(n1137), .ZN(n1136) );
  AND2_X1 U4023 ( .A1(n1139), .A2(n16546), .ZN(n1137) );
  XNOR2_X1 U4024 ( .A(n1140), .B(n23693), .ZN(Ciphertext[129]) );
  NAND3_X1 U4025 ( .A1(n1143), .A2(n1142), .A3(n1141), .ZN(n1140) );
  NAND2_X1 U4026 ( .A1(n23691), .A2(n25026), .ZN(n1141) );
  NAND2_X1 U4027 ( .A1(n25405), .A2(n23686), .ZN(n1142) );
  NOR2_X1 U4028 ( .A1(n23670), .A2(n25026), .ZN(n23686) );
  NAND2_X1 U4029 ( .A1(n1144), .A2(n23670), .ZN(n1143) );
  NAND3_X1 U4030 ( .A1(n4702), .A2(n4703), .A3(n4700), .ZN(Ciphertext[130]) );
  NAND2_X1 U4031 ( .A1(n22200), .A2(n1146), .ZN(n22179) );
  NAND2_X1 U4032 ( .A1(n325), .A2(n1146), .ZN(n4362) );
  OAI21_X1 U4033 ( .B1(n325), .B2(n1146), .A(n22200), .ZN(n21804) );
  NAND2_X1 U4035 ( .A1(n6976), .A2(n1147), .ZN(n6692) );
  NAND2_X1 U4037 ( .A1(n6686), .A2(n1147), .ZN(n6390) );
  INV_X1 U4039 ( .A(n6690), .ZN(n1149) );
  NAND2_X1 U4040 ( .A1(n1150), .A2(n4110), .ZN(n1613) );
  NAND2_X1 U4042 ( .A1(n4175), .A2(n20384), .ZN(n1152) );
  NAND2_X1 U4043 ( .A1(n1613), .A2(n4176), .ZN(n21743) );
  OAI21_X2 U4044 ( .B1(n19882), .B2(n20554), .A(n19881), .ZN(n1153) );
  XNOR2_X1 U4045 ( .A(n1153), .B(n21985), .ZN(n20818) );
  XNOR2_X1 U4046 ( .A(n1153), .B(n452), .ZN(n20991) );
  XNOR2_X1 U4047 ( .A(n1153), .B(n1758), .ZN(n21462) );
  NOR2_X1 U4049 ( .A1(n23652), .A2(n23649), .ZN(n22151) );
  NAND2_X1 U4050 ( .A1(n20856), .A2(n2601), .ZN(n1156) );
  NAND2_X1 U4051 ( .A1(n21802), .A2(n22200), .ZN(n1158) );
  NAND2_X1 U4052 ( .A1(n18922), .A2(n264), .ZN(n1161) );
  NAND2_X1 U4053 ( .A1(n14044), .A2(n5246), .ZN(n1930) );
  NAND2_X1 U4054 ( .A1(n20111), .A2(n19916), .ZN(n5123) );
  NOR2_X2 U4055 ( .A1(n17714), .A2(n17713), .ZN(n19883) );
  NAND3_X1 U4056 ( .A1(n1162), .A2(n7078), .A3(n25251), .ZN(n7075) );
  MUX2_X2 U4057 ( .A(n7226), .B(n7227), .S(n7676), .Z(n8491) );
  NAND2_X1 U4059 ( .A1(n24083), .A2(n9944), .ZN(n1165) );
  MUX2_X1 U4061 ( .A(n10848), .B(n10850), .S(n11122), .Z(n1166) );
  NAND2_X1 U4063 ( .A1(n3546), .A2(n1479), .ZN(n10848) );
  INV_X1 U4064 ( .A(n11124), .ZN(n1167) );
  NAND2_X1 U4066 ( .A1(n10721), .A2(n11124), .ZN(n1170) );
  OAI211_X1 U4067 ( .C1(n7008), .C2(n7009), .A(n1173), .B(n7006), .ZN(n1174)
         );
  NAND2_X1 U4068 ( .A1(n7009), .A2(n7004), .ZN(n1173) );
  NAND2_X1 U4069 ( .A1(n283), .A2(n17068), .ZN(n16611) );
  NAND3_X1 U4070 ( .A1(n283), .A2(n17068), .A3(n16612), .ZN(n5307) );
  INV_X1 U4071 ( .A(n6198), .ZN(n1175) );
  NOR2_X1 U4073 ( .A1(n25480), .A2(n1176), .ZN(n5964) );
  AOI21_X1 U4074 ( .B1(n6923), .B2(n6922), .A(n1176), .ZN(n6928) );
  INV_X1 U4075 ( .A(n6776), .ZN(n1176) );
  XNOR2_X1 U4076 ( .A(n1177), .B(n21662), .ZN(n10431) );
  XNOR2_X1 U4077 ( .A(n1177), .B(n21553), .ZN(n9406) );
  XNOR2_X1 U4078 ( .A(n11735), .B(n1177), .ZN(n10638) );
  XNOR2_X1 U4079 ( .A(n11564), .B(n1177), .ZN(n11537) );
  NAND3_X2 U4080 ( .A1(n9404), .A2(n9405), .A3(n1178), .ZN(n1177) );
  NOR2_X2 U4081 ( .A1(n19840), .A2(n1179), .ZN(n3198) );
  OAI22_X1 U4082 ( .A1(n3203), .A2(n19390), .B1(n24909), .B2(n3202), .ZN(n1179) );
  AND2_X1 U4083 ( .A1(n3198), .A2(n19839), .ZN(n19842) );
  NAND2_X1 U4085 ( .A1(n411), .A2(n10798), .ZN(n1180) );
  NAND2_X1 U4086 ( .A1(n10651), .A2(n10245), .ZN(n10243) );
  NAND2_X1 U4087 ( .A1(n9932), .A2(n25217), .ZN(n1182) );
  AOI22_X1 U4088 ( .A1(n9345), .A2(n9928), .B1(n9926), .B2(n9925), .ZN(n1183)
         );
  AOI21_X2 U4089 ( .B1(n1186), .B2(n1185), .A(n1184), .ZN(n10651) );
  NAND2_X1 U4090 ( .A1(n1602), .A2(n4166), .ZN(n1184) );
  OAI21_X2 U4091 ( .B1(n17730), .B2(n1189), .A(n1187), .ZN(n18370) );
  MUX2_X1 U4092 ( .A(n17731), .B(n1188), .S(n25472), .Z(n1187) );
  NAND2_X1 U4093 ( .A1(n17733), .A2(n17486), .ZN(n1188) );
  MUX2_X1 U4094 ( .A(n17728), .B(n17729), .S(n17486), .Z(n1189) );
  NOR2_X2 U4095 ( .A1(n15841), .A2(n15840), .ZN(n17486) );
  NAND2_X1 U4096 ( .A1(n1194), .A2(n7588), .ZN(n1191) );
  NAND3_X1 U4097 ( .A1(n1839), .A2(n7590), .A3(n7462), .ZN(n1193) );
  NAND2_X1 U4098 ( .A1(n7588), .A2(n7590), .ZN(n7593) );
  NAND3_X1 U4099 ( .A1(n2035), .A2(n7591), .A3(n7464), .ZN(n1195) );
  NAND2_X1 U4100 ( .A1(n7236), .A2(n7962), .ZN(n1196) );
  NAND2_X1 U4101 ( .A1(n25024), .A2(n23064), .ZN(n1198) );
  NAND2_X1 U4102 ( .A1(n1199), .A2(n10951), .ZN(n10957) );
  NAND2_X1 U4103 ( .A1(n2754), .A2(n10950), .ZN(n1199) );
  NAND2_X1 U4104 ( .A1(n10698), .A2(n25074), .ZN(n10950) );
  NAND2_X1 U4105 ( .A1(n13275), .A2(n1201), .ZN(n13276) );
  NOR2_X1 U4107 ( .A1(n367), .A2(n4004), .ZN(n3655) );
  OR2_X1 U4109 ( .A1(n16272), .A2(n4516), .ZN(n1202) );
  NAND2_X1 U4110 ( .A1(n296), .A2(n1028), .ZN(n1204) );
  NAND3_X1 U4111 ( .A1(n296), .A2(n1028), .A3(n14153), .ZN(n14152) );
  NOR2_X1 U4113 ( .A1(n13512), .A2(n14031), .ZN(n1203) );
  AND2_X1 U4114 ( .A1(n20193), .A2(n20576), .ZN(n1206) );
  NAND2_X1 U4116 ( .A1(n3198), .A2(n20576), .ZN(n20438) );
  NAND2_X1 U4118 ( .A1(n1208), .A2(n15811), .ZN(n15812) );
  NAND2_X1 U4119 ( .A1(n16404), .A2(n16401), .ZN(n1208) );
  OR2_X1 U4121 ( .A1(n9523), .A2(n1210), .ZN(n3028) );
  INV_X1 U4122 ( .A(n9843), .ZN(n1210) );
  OR2_X1 U4123 ( .A1(n1211), .A2(n19103), .ZN(n18021) );
  NOR2_X1 U4124 ( .A1(n19360), .A2(n24312), .ZN(n1211) );
  INV_X1 U4126 ( .A(n18817), .ZN(n1212) );
  NAND2_X1 U4127 ( .A1(n16404), .A2(n15646), .ZN(n1214) );
  NAND2_X1 U4129 ( .A1(n9803), .A2(n11053), .ZN(n1216) );
  NAND2_X1 U4130 ( .A1(n1218), .A2(n11058), .ZN(n1217) );
  NAND2_X1 U4131 ( .A1(n1523), .A2(n11499), .ZN(n1219) );
  NAND2_X1 U4132 ( .A1(n9802), .A2(n11499), .ZN(n1220) );
  NAND2_X1 U4133 ( .A1(n24499), .A2(n12459), .ZN(n12653) );
  OAI21_X1 U4135 ( .B1(n13177), .B2(n13176), .A(n12506), .ZN(n10362) );
  INV_X1 U4137 ( .A(n11205), .ZN(n1224) );
  NAND2_X1 U4138 ( .A1(n4152), .A2(n10819), .ZN(n1226) );
  NAND3_X1 U4140 ( .A1(n25025), .A2(n11342), .A3(n1224), .ZN(n1223) );
  NAND2_X1 U4141 ( .A1(n10232), .A2(n414), .ZN(n1227) );
  NAND2_X1 U4143 ( .A1(n1233), .A2(n1228), .ZN(n18146) );
  NAND2_X1 U4144 ( .A1(n14353), .A2(n25246), .ZN(n1233) );
  NAND2_X1 U4145 ( .A1(n15865), .A2(n15866), .ZN(n1235) );
  XNOR2_X2 U4147 ( .A(n21315), .B(n21314), .ZN(n22222) );
  INV_X1 U4148 ( .A(n22221), .ZN(n1238) );
  XNOR2_X2 U4149 ( .A(n21330), .B(n21329), .ZN(n22221) );
  NAND2_X1 U4150 ( .A1(n1239), .A2(n10558), .ZN(n10337) );
  INV_X1 U4151 ( .A(n25250), .ZN(n1239) );
  NAND3_X1 U4152 ( .A1(n1239), .A2(n10559), .A3(n10655), .ZN(n4540) );
  NAND2_X1 U4153 ( .A1(n1240), .A2(n10314), .ZN(n10316) );
  NAND2_X1 U4154 ( .A1(n10558), .A2(n25250), .ZN(n1240) );
  NOR2_X1 U4155 ( .A1(n19862), .A2(n1242), .ZN(n19865) );
  OAI21_X1 U4156 ( .B1(n20038), .B2(n20191), .A(n1241), .ZN(n20040) );
  NAND2_X1 U4157 ( .A1(n20038), .A2(n20039), .ZN(n1241) );
  NOR2_X1 U4158 ( .A1(n20185), .A2(n1242), .ZN(n20187) );
  NAND2_X1 U4159 ( .A1(n1244), .A2(n17598), .ZN(n1243) );
  NAND3_X1 U4160 ( .A1(n3316), .A2(n4574), .A3(n1483), .ZN(n1245) );
  NAND2_X1 U4161 ( .A1(n17596), .A2(n24543), .ZN(n1246) );
  NOR2_X1 U4162 ( .A1(n14180), .A2(n1247), .ZN(n14183) );
  INV_X1 U4163 ( .A(n14181), .ZN(n1247) );
  INV_X1 U4164 ( .A(n21839), .ZN(n22358) );
  NOR2_X1 U4165 ( .A1(n22361), .A2(n22358), .ZN(n1248) );
  AND2_X1 U4166 ( .A1(n21782), .A2(n22361), .ZN(n22359) );
  INV_X1 U4167 ( .A(n21838), .ZN(n21782) );
  NAND2_X1 U4170 ( .A1(n24172), .A2(n19459), .ZN(n1251) );
  NAND2_X1 U4171 ( .A1(n15938), .A2(n16247), .ZN(n2359) );
  NAND2_X1 U4172 ( .A1(n16018), .A2(n15938), .ZN(n15568) );
  NAND2_X1 U4173 ( .A1(n17058), .A2(n17057), .ZN(n1252) );
  NAND2_X1 U4174 ( .A1(n1254), .A2(n7893), .ZN(n7455) );
  NAND2_X1 U4175 ( .A1(n1254), .A2(n7889), .ZN(n7325) );
  OAI21_X1 U4176 ( .B1(n20410), .B2(n20411), .A(n345), .ZN(n1255) );
  NAND2_X1 U4177 ( .A1(n20872), .A2(n20412), .ZN(n20873) );
  MUX2_X1 U4178 ( .A(n25421), .B(n20411), .S(n20262), .Z(n20872) );
  MUX2_X1 U4179 ( .A(n22952), .B(n22033), .S(n22954), .Z(n1259) );
  XNOR2_X2 U4180 ( .A(n21605), .B(n21604), .ZN(n22954) );
  AND2_X1 U4182 ( .A1(n15804), .A2(n1261), .ZN(n4337) );
  NOR2_X1 U4183 ( .A1(n15856), .A2(n1261), .ZN(n15858) );
  MUX2_X1 U4185 ( .A(n15856), .B(n16117), .S(n1261), .Z(n4338) );
  MUX2_X1 U4186 ( .A(n15614), .B(n15613), .S(n1261), .Z(n15617) );
  XNOR2_X2 U4188 ( .A(n14481), .B(n14480), .ZN(n1261) );
  INV_X1 U4190 ( .A(n1263), .ZN(n1262) );
  NAND2_X1 U4193 ( .A1(n3119), .A2(n10767), .ZN(n11082) );
  NAND2_X1 U4194 ( .A1(n1503), .A2(n1504), .ZN(n20383) );
  NAND2_X1 U4195 ( .A1(n3943), .A2(n1506), .ZN(n1503) );
  NAND2_X1 U4196 ( .A1(n1266), .A2(n1265), .ZN(n3943) );
  NAND2_X1 U4197 ( .A1(n1268), .A2(n12503), .ZN(n5402) );
  XNOR2_X1 U4200 ( .A(n18258), .B(n25000), .ZN(n18619) );
  NAND2_X1 U4202 ( .A1(n9524), .A2(n9774), .ZN(n1272) );
  NAND2_X1 U4203 ( .A1(n25393), .A2(n9772), .ZN(n1273) );
  INV_X1 U4206 ( .A(n22268), .ZN(n1276) );
  NAND2_X1 U4209 ( .A1(n7914), .A2(n7917), .ZN(n1281) );
  NAND2_X1 U4210 ( .A1(n7634), .A2(n7449), .ZN(n7920) );
  INV_X1 U4211 ( .A(n17237), .ZN(n1285) );
  OAI211_X1 U4212 ( .C1(n16859), .C2(n17236), .A(n1284), .B(n1283), .ZN(n16860) );
  NAND2_X1 U4213 ( .A1(n17341), .A2(n3872), .ZN(n1286) );
  INV_X1 U4214 ( .A(n17346), .ZN(n17236) );
  NAND2_X2 U4215 ( .A1(n1763), .A2(n15365), .ZN(n17346) );
  AND3_X2 U4216 ( .A1(n15309), .A2(n1812), .A3(n15310), .ZN(n17241) );
  INV_X1 U4217 ( .A(n1289), .ZN(n1288) );
  AOI21_X1 U4218 ( .B1(n18835), .B2(n19437), .A(n25422), .ZN(n1289) );
  NAND2_X1 U4219 ( .A1(n361), .A2(n18834), .ZN(n19437) );
  AND2_X1 U4220 ( .A1(n19441), .A2(n25422), .ZN(n1291) );
  INV_X1 U4221 ( .A(n19441), .ZN(n19245) );
  AND2_X1 U4222 ( .A1(n24922), .A2(n24885), .ZN(n22956) );
  NOR2_X1 U4223 ( .A1(n22958), .A2(n1292), .ZN(n21879) );
  NAND2_X1 U4224 ( .A1(n24884), .A2(n1293), .ZN(n1292) );
  NOR2_X1 U4225 ( .A1(n6481), .A2(n6198), .ZN(n1294) );
  INV_X1 U4227 ( .A(n9418), .ZN(n9973) );
  NAND2_X1 U4228 ( .A1(n25005), .A2(n9418), .ZN(n9417) );
  NAND2_X1 U4229 ( .A1(n1296), .A2(n1712), .ZN(n19726) );
  NAND2_X1 U4230 ( .A1(n1714), .A2(n19404), .ZN(n1296) );
  OR2_X1 U4232 ( .A1(n6244), .A2(n1297), .ZN(n6641) );
  NAND2_X1 U4233 ( .A1(n6987), .A2(n6640), .ZN(n1297) );
  INV_X1 U4235 ( .A(n19261), .ZN(n1299) );
  NOR2_X1 U4236 ( .A1(n19264), .A2(n1300), .ZN(n17558) );
  AOI21_X1 U4237 ( .B1(n1299), .B2(n19264), .A(n1300), .ZN(n18918) );
  INV_X1 U4238 ( .A(n18914), .ZN(n1300) );
  NAND2_X1 U4239 ( .A1(n1304), .A2(n1301), .ZN(n21282) );
  NAND2_X1 U4240 ( .A1(n22578), .A2(n1302), .ZN(n1301) );
  NAND2_X1 U4241 ( .A1(n23064), .A2(n23077), .ZN(n1302) );
  NAND2_X1 U4244 ( .A1(n1309), .A2(n18586), .ZN(n1308) );
  AOI21_X1 U4245 ( .B1(n1311), .B2(n1310), .A(n328), .ZN(n1312) );
  INV_X1 U4246 ( .A(n21794), .ZN(n1311) );
  NAND3_X2 U4247 ( .A1(n2811), .A2(n16501), .A3(n1313), .ZN(n18331) );
  NAND2_X1 U4250 ( .A1(n12979), .A2(n25053), .ZN(n1315) );
  INV_X1 U4252 ( .A(n9808), .ZN(n9339) );
  AND2_X1 U4253 ( .A1(n10284), .A2(n11113), .ZN(n10285) );
  NAND2_X1 U4254 ( .A1(n10870), .A2(n10873), .ZN(n10284) );
  NAND2_X1 U4255 ( .A1(n9337), .A2(n9529), .ZN(n1317) );
  NAND3_X1 U4256 ( .A1(n6274), .A2(n6324), .A3(n315), .ZN(n1320) );
  NAND2_X1 U4258 ( .A1(n6518), .A2(n6517), .ZN(n1321) );
  NAND3_X1 U4259 ( .A1(n1322), .A2(n23053), .A3(n23052), .ZN(n23054) );
  INV_X1 U4260 ( .A(n23571), .ZN(n1323) );
  INV_X2 U4261 ( .A(n18596), .ZN(n19760) );
  XNOR2_X1 U4262 ( .A(n11237), .B(n11568), .ZN(n11880) );
  AND2_X1 U4263 ( .A1(n5440), .A2(n13868), .ZN(n13600) );
  XNOR2_X1 U4264 ( .A(n10320), .B(n1325), .ZN(n1324) );
  XOR2_X1 U4265 ( .A(n11536), .B(n10310), .Z(n1325) );
  OR2_X1 U4266 ( .A1(n10772), .A2(n415), .ZN(n11033) );
  INV_X1 U4269 ( .A(n24397), .ZN(n1328) );
  OAI211_X1 U4270 ( .C1(n12931), .C2(n12930), .A(n4457), .B(n12929), .ZN(n1331) );
  OR2_X1 U4271 ( .A1(n8752), .A2(n2159), .ZN(n1332) );
  XNOR2_X1 U4272 ( .A(n14426), .B(n14425), .ZN(n16423) );
  XNOR2_X1 U4273 ( .A(n8717), .B(n8718), .ZN(n10071) );
  OAI211_X1 U4274 ( .C1(n12931), .C2(n12930), .A(n4457), .B(n12929), .ZN(
        n14129) );
  XOR2_X1 U4276 ( .A(n18266), .B(n18265), .Z(n1334) );
  XOR2_X1 U4277 ( .A(n11364), .B(n11365), .Z(n1335) );
  XNOR2_X1 U4278 ( .A(n3141), .B(n21748), .ZN(n1336) );
  XOR2_X1 U4279 ( .A(n8088), .B(n9169), .Z(n1337) );
  OR2_X1 U4280 ( .A1(n17293), .A2(n17233), .ZN(n1339) );
  XNOR2_X1 U4282 ( .A(n3141), .B(n21748), .ZN(n22245) );
  NAND2_X1 U4287 ( .A1(n14236), .A2(n14235), .ZN(n1342) );
  NAND2_X1 U4288 ( .A1(n14234), .A2(n14233), .ZN(n1343) );
  XOR2_X1 U4292 ( .A(n11243), .B(n11741), .Z(n12322) );
  INV_X1 U4293 ( .A(n15715), .ZN(n16474) );
  OAI21_X1 U4294 ( .B1(n15820), .B2(n15819), .A(n16426), .ZN(n15835) );
  OAI211_X2 U4295 ( .C1(n11008), .C2(n4088), .A(n4495), .B(n1921), .ZN(n12295)
         );
  AND2_X1 U4296 ( .A1(n19320), .A2(n19319), .ZN(n1344) );
  NAND2_X1 U4297 ( .A1(n10093), .A2(n9676), .ZN(n1347) );
  XNOR2_X1 U4298 ( .A(n2276), .B(n1903), .ZN(n1348) );
  XNOR2_X1 U4299 ( .A(n1903), .B(n2276), .ZN(n9779) );
  NAND3_X1 U4300 ( .A1(n1727), .A2(n2926), .A3(n5231), .ZN(n1349) );
  NOR2_X1 U4302 ( .A1(n13523), .A2(n13522), .ZN(n1351) );
  XNOR2_X1 U4303 ( .A(n20750), .B(n20749), .ZN(n1352) );
  XNOR2_X1 U4304 ( .A(n11650), .B(n11649), .ZN(n1353) );
  NAND3_X1 U4306 ( .A1(n1727), .A2(n2926), .A3(n5231), .ZN(n23157) );
  NOR2_X1 U4307 ( .A1(n13523), .A2(n13522), .ZN(n15005) );
  XNOR2_X1 U4308 ( .A(n18527), .B(n18526), .ZN(n19238) );
  XNOR2_X1 U4309 ( .A(n20750), .B(n20749), .ZN(n22270) );
  XNOR2_X1 U4310 ( .A(n11650), .B(n11649), .ZN(n13159) );
  XOR2_X1 U4311 ( .A(n14763), .B(n15106), .Z(n14767) );
  XOR2_X1 U4312 ( .A(n14858), .B(n14857), .Z(n15160) );
  AOI21_X2 U4314 ( .B1(n15759), .B2(n5666), .A(n5668), .ZN(n16539) );
  OAI21_X1 U4315 ( .B1(n1871), .B2(n9691), .A(n9690), .ZN(n10961) );
  INV_X1 U4316 ( .A(n11158), .ZN(n1358) );
  NOR2_X1 U4320 ( .A1(n13799), .A2(n13798), .ZN(n1359) );
  XOR2_X1 U4322 ( .A(n18379), .B(n18378), .Z(n1361) );
  NOR2_X1 U4323 ( .A1(n13799), .A2(n13798), .ZN(n14982) );
  XNOR2_X1 U4324 ( .A(n8939), .B(n2276), .ZN(n9255) );
  MUX2_X1 U4325 ( .A(n22706), .B(n23278), .S(n23265), .Z(n22707) );
  INV_X1 U4326 ( .A(n23265), .ZN(n23274) );
  AND2_X1 U4327 ( .A1(n13035), .A2(n13036), .ZN(n1362) );
  OAI21_X2 U4329 ( .B1(n12923), .B2(n12924), .A(n12922), .ZN(n14127) );
  XOR2_X1 U4330 ( .A(n8427), .B(n8846), .Z(n8628) );
  XNOR2_X2 U4332 ( .A(n5894), .B(Key[50]), .ZN(n6699) );
  AOI22_X1 U4333 ( .A1(n16015), .A2(n16345), .B1(n16014), .B2(n24539), .ZN(
        n17463) );
  INV_X1 U4335 ( .A(n16106), .ZN(n4689) );
  AOI21_X1 U4336 ( .B1(n15592), .B2(n15591), .A(n15590), .ZN(n17065) );
  OAI21_X2 U4337 ( .B1(n6711), .B2(n7998), .A(n6710), .ZN(n8846) );
  INV_X1 U4342 ( .A(n7628), .ZN(n7913) );
  OR2_X1 U4343 ( .A1(n9433), .A2(n10037), .ZN(n9714) );
  XNOR2_X1 U4344 ( .A(n310), .B(n8506), .ZN(n8084) );
  INV_X1 U4345 ( .A(n10169), .ZN(n2207) );
  INV_X1 U4347 ( .A(n12040), .ZN(n12213) );
  INV_X1 U4348 ( .A(n10934), .ZN(n2311) );
  XNOR2_X1 U4349 ( .A(n3899), .B(n12355), .ZN(n11194) );
  INV_X1 U4350 ( .A(n11268), .ZN(n3899) );
  OR2_X1 U4351 ( .A1(n10811), .A2(n10812), .ZN(n5629) );
  OR2_X1 U4352 ( .A1(n11298), .A2(n10762), .ZN(n10763) );
  INV_X1 U4353 ( .A(n25027), .ZN(n3512) );
  OR2_X1 U4354 ( .A1(n12773), .A2(n12774), .ZN(n13069) );
  NOR2_X1 U4355 ( .A1(n13071), .A2(n12470), .ZN(n1544) );
  INV_X1 U4356 ( .A(n12856), .ZN(n4196) );
  INV_X1 U4357 ( .A(n13347), .ZN(n3766) );
  XNOR2_X1 U4358 ( .A(n11076), .B(n11582), .ZN(n12046) );
  XNOR2_X1 U4360 ( .A(n12131), .B(n3206), .ZN(n3204) );
  XNOR2_X1 U4361 ( .A(n12127), .B(n2834), .ZN(n3206) );
  XNOR2_X1 U4362 ( .A(n4996), .B(n4995), .ZN(n11328) );
  XNOR2_X1 U4363 ( .A(n11321), .B(n11320), .ZN(n4995) );
  NOR2_X1 U4364 ( .A1(n12951), .A2(n2295), .ZN(n12604) );
  AND2_X1 U4365 ( .A1(n24346), .A2(n404), .ZN(n3813) );
  XNOR2_X1 U4367 ( .A(n3862), .B(n3861), .ZN(n11722) );
  XNOR2_X1 U4368 ( .A(n11880), .B(n11700), .ZN(n3861) );
  XNOR2_X1 U4369 ( .A(n11699), .B(n11702), .ZN(n3862) );
  INV_X1 U4371 ( .A(n3341), .ZN(n14206) );
  INV_X1 U4372 ( .A(n13386), .ZN(n13646) );
  OR2_X1 U4373 ( .A1(n13277), .A2(n24346), .ZN(n4387) );
  INV_X1 U4374 ( .A(n13864), .ZN(n5230) );
  MUX2_X1 U4375 ( .A(n13401), .B(n13400), .S(n14225), .Z(n13402) );
  INV_X1 U4376 ( .A(n15802), .ZN(n16075) );
  INV_X1 U4377 ( .A(n16394), .ZN(n16167) );
  AND2_X1 U4378 ( .A1(n15198), .A2(n3554), .ZN(n3553) );
  XNOR2_X1 U4379 ( .A(n2862), .B(n14555), .ZN(n16151) );
  INV_X1 U4380 ( .A(n16312), .ZN(n16309) );
  OR2_X1 U4381 ( .A1(n4869), .A2(n15647), .ZN(n4575) );
  INV_X1 U4382 ( .A(n15640), .ZN(n3380) );
  INV_X1 U4383 ( .A(n17183), .ZN(n16204) );
  XNOR2_X1 U4384 ( .A(n4967), .B(n4965), .ZN(n16422) );
  XNOR2_X1 U4385 ( .A(n14428), .B(n4966), .ZN(n4965) );
  NOR2_X1 U4386 ( .A1(n24981), .A2(n5039), .ZN(n5038) );
  AND2_X1 U4387 ( .A1(n16481), .A2(n16480), .ZN(n5039) );
  AOI22_X1 U4388 ( .A1(n16495), .A2(n16494), .B1(n16493), .B2(n16492), .ZN(
        n16516) );
  OAI211_X1 U4389 ( .C1(n16104), .C2(n16105), .A(n3409), .B(n3408), .ZN(n17524) );
  OR2_X1 U4390 ( .A1(n16103), .A2(n3410), .ZN(n3409) );
  INV_X1 U4391 ( .A(n17524), .ZN(n16863) );
  OR2_X1 U4392 ( .A1(n16798), .A2(n5375), .ZN(n5240) );
  XNOR2_X1 U4393 ( .A(n17814), .B(n18562), .ZN(n17815) );
  INV_X1 U4394 ( .A(n1653), .ZN(n17144) );
  NAND3_X1 U4395 ( .A1(n16468), .A2(n4725), .A3(n4724), .ZN(n16984) );
  OR2_X1 U4397 ( .A1(n15796), .A2(n382), .ZN(n4858) );
  INV_X1 U4398 ( .A(n17515), .ZN(n18258) );
  OR2_X1 U4399 ( .A1(n19520), .A2(n19284), .ZN(n4433) );
  XNOR2_X1 U4401 ( .A(n1386), .B(n17092), .ZN(n4214) );
  NAND2_X1 U4403 ( .A1(n18840), .A2(n19322), .ZN(n3584) );
  OR2_X1 U4404 ( .A1(n18961), .A2(n19467), .ZN(n3579) );
  INV_X1 U4405 ( .A(n17567), .ZN(n19714) );
  OR2_X1 U4406 ( .A1(n20203), .A2(n20204), .ZN(n1664) );
  XNOR2_X1 U4407 ( .A(n3823), .B(n21043), .ZN(n21229) );
  XNOR2_X1 U4408 ( .A(n21266), .B(n24485), .ZN(n3746) );
  OR2_X1 U4410 ( .A1(n20368), .A2(n24454), .ZN(n20303) );
  XNOR2_X1 U4411 ( .A(n19161), .B(n19160), .ZN(n22255) );
  OR2_X1 U4412 ( .A1(n6034), .A2(n441), .ZN(n6171) );
  INV_X1 U4414 ( .A(n7782), .ZN(n7174) );
  AND2_X1 U4415 ( .A1(n2974), .A2(n2973), .ZN(n6613) );
  INV_X1 U4416 ( .A(n7991), .ZN(n7357) );
  INV_X1 U4418 ( .A(n8132), .ZN(n8845) );
  INV_X1 U4419 ( .A(n8428), .ZN(n4335) );
  XNOR2_X1 U4420 ( .A(n8476), .B(n2191), .ZN(n4395) );
  NAND2_X1 U4422 ( .A1(n1693), .A2(n1692), .ZN(n7234) );
  AND2_X1 U4423 ( .A1(n7004), .A2(n448), .ZN(n5148) );
  OR2_X1 U4424 ( .A1(n7892), .A2(n7322), .ZN(n3082) );
  XNOR2_X1 U4425 ( .A(n8730), .B(n8468), .ZN(n8797) );
  OR2_X1 U4427 ( .A1(n9220), .A2(n9705), .ZN(n3721) );
  NAND2_X1 U4428 ( .A1(n7532), .A2(n7533), .ZN(n1972) );
  INV_X1 U4429 ( .A(n8476), .ZN(n4401) );
  OR2_X1 U4430 ( .A1(n9127), .A2(n10063), .ZN(n9220) );
  NOR2_X1 U4431 ( .A1(n1517), .A2(n24549), .ZN(n9876) );
  INV_X1 U4432 ( .A(n10138), .ZN(n1649) );
  OR2_X1 U4433 ( .A1(n10099), .A2(n9515), .ZN(n10097) );
  OAI21_X1 U4434 ( .B1(n2267), .B2(n9615), .A(n1412), .ZN(n3546) );
  OR2_X1 U4435 ( .A1(n9754), .A2(n9613), .ZN(n1412) );
  AND2_X1 U4436 ( .A1(n10161), .A2(n24984), .ZN(n9382) );
  BUF_X1 U4437 ( .A(n9515), .Z(n10098) );
  XNOR2_X1 U4440 ( .A(n8806), .B(n1831), .ZN(n2491) );
  NOR2_X1 U4441 ( .A1(n4254), .A2(n25393), .ZN(n3865) );
  AND2_X1 U4443 ( .A1(n13049), .A2(n13048), .ZN(n1545) );
  AND2_X1 U4444 ( .A1(n2524), .A2(n2523), .ZN(n10312) );
  INV_X1 U4445 ( .A(n3375), .ZN(n11307) );
  AND2_X1 U4446 ( .A1(n11012), .A2(n11045), .ZN(n10415) );
  INV_X1 U4447 ( .A(n2295), .ZN(n13327) );
  OR2_X1 U4448 ( .A1(n13076), .A2(n3704), .ZN(n13080) );
  INV_X1 U4449 ( .A(n3492), .ZN(n4405) );
  OR2_X1 U4450 ( .A1(n10711), .A2(n13132), .ZN(n13158) );
  XNOR2_X1 U4451 ( .A(n11546), .B(n11547), .ZN(n12773) );
  INV_X1 U4452 ( .A(n11981), .ZN(n4931) );
  INV_X1 U4453 ( .A(n12934), .ZN(n5361) );
  OAI211_X1 U4456 ( .C1(n13104), .C2(n13103), .A(n12658), .B(n12657), .ZN(
        n12668) );
  INV_X1 U4457 ( .A(n3958), .ZN(n12654) );
  XNOR2_X1 U4458 ( .A(n11760), .B(n4134), .ZN(n13223) );
  OR2_X1 U4459 ( .A1(n3460), .A2(n3492), .ZN(n5325) );
  XNOR2_X1 U4460 ( .A(n11268), .B(n3900), .ZN(n11626) );
  NOR2_X1 U4461 ( .A1(n12583), .A2(n24554), .ZN(n12624) );
  OR2_X1 U4462 ( .A1(n13122), .A2(n5626), .ZN(n2516) );
  OR2_X1 U4463 ( .A1(n12873), .A2(n13123), .ZN(n2515) );
  OR2_X1 U4465 ( .A1(n12452), .A2(n304), .ZN(n3523) );
  OR2_X1 U4466 ( .A1(n12453), .A2(n4766), .ZN(n3524) );
  OR2_X1 U4467 ( .A1(n13025), .A2(n13030), .ZN(n1634) );
  NOR2_X1 U4469 ( .A1(n4790), .A2(n4789), .ZN(n4788) );
  AND2_X1 U4470 ( .A1(n4791), .A2(n3858), .ZN(n3860) );
  OR2_X1 U4472 ( .A1(n5359), .A2(n4499), .ZN(n2715) );
  AND2_X1 U4473 ( .A1(n12610), .A2(n1971), .ZN(n1970) );
  OR2_X1 U4474 ( .A1(n12606), .A2(n12683), .ZN(n2840) );
  OAI21_X1 U4475 ( .B1(n12965), .B2(n3813), .A(n13273), .ZN(n2158) );
  INV_X1 U4476 ( .A(n14167), .ZN(n14164) );
  OR2_X1 U4478 ( .A1(n4529), .A2(n12634), .ZN(n2721) );
  AOI21_X1 U4479 ( .B1(n14067), .B2(n13845), .A(n13627), .ZN(n12592) );
  INV_X1 U4480 ( .A(n15556), .ZN(n2173) );
  AND3_X1 U4481 ( .A1(n14327), .A2(n14044), .A3(n13864), .ZN(n2225) );
  NOR2_X1 U4482 ( .A1(n4870), .A2(n24062), .ZN(n4869) );
  OR2_X1 U4484 ( .A1(n16206), .A2(n15640), .ZN(n16207) );
  AND2_X1 U4485 ( .A1(n16324), .A2(n2610), .ZN(n16194) );
  AOI22_X1 U4486 ( .A1(n388), .A2(n290), .B1(n1123), .B2(n16331), .ZN(n16185)
         );
  XNOR2_X1 U4487 ( .A(n15237), .B(n15236), .ZN(n15674) );
  OAI21_X1 U4488 ( .B1(n386), .B2(n15992), .A(n15991), .ZN(n4646) );
  INV_X1 U4489 ( .A(n15839), .ZN(n16175) );
  XNOR2_X1 U4490 ( .A(n5757), .B(n13424), .ZN(n15915) );
  XNOR2_X1 U4491 ( .A(n4712), .B(n3694), .ZN(n16418) );
  INV_X1 U4492 ( .A(n16246), .ZN(n16253) );
  AND2_X1 U4493 ( .A1(n25484), .A2(n15764), .ZN(n15940) );
  INV_X1 U4496 ( .A(n16418), .ZN(n16413) );
  INV_X1 U4497 ( .A(n15842), .ZN(n2996) );
  XNOR2_X1 U4499 ( .A(n14592), .B(n1383), .ZN(n4205) );
  XNOR2_X1 U4500 ( .A(n4095), .B(n14593), .ZN(n4204) );
  INV_X1 U4501 ( .A(n2253), .ZN(n2251) );
  OAI21_X1 U4503 ( .B1(n16274), .B2(n16029), .A(n2280), .ZN(n16034) );
  AOI22_X1 U4504 ( .A1(n16133), .A2(n16075), .B1(n16132), .B2(n16131), .ZN(
        n16431) );
  OR2_X1 U4505 ( .A1(n15983), .A2(n16163), .ZN(n3008) );
  NAND3_X1 U4507 ( .A1(n16146), .A2(n2541), .A3(n16098), .ZN(n16434) );
  AOI22_X1 U4508 ( .A1(n16838), .A2(n16261), .B1(n16533), .B2(n17165), .ZN(
        n16378) );
  XNOR2_X1 U4509 ( .A(n17811), .B(n17969), .ZN(n18248) );
  INV_X1 U4511 ( .A(n17815), .ZN(n18287) );
  INV_X1 U4512 ( .A(n19278), .ZN(n5573) );
  XNOR2_X1 U4513 ( .A(n17639), .B(n18051), .ZN(n18734) );
  XNOR2_X1 U4514 ( .A(n18578), .B(n18577), .ZN(n18998) );
  AND2_X1 U4515 ( .A1(n18998), .A2(n19418), .ZN(n19002) );
  INV_X1 U4516 ( .A(n19488), .ZN(n19346) );
  AND2_X1 U4517 ( .A1(n18734), .A2(n19476), .ZN(n5685) );
  XNOR2_X1 U4518 ( .A(n18354), .B(n18353), .ZN(n18385) );
  INV_X1 U4519 ( .A(n18998), .ZN(n19421) );
  OR2_X1 U4520 ( .A1(n19413), .A2(n25469), .ZN(n19409) );
  XNOR2_X1 U4521 ( .A(n2692), .B(n17777), .ZN(n2029) );
  XNOR2_X1 U4522 ( .A(n18681), .B(n18682), .ZN(n19408) );
  XNOR2_X1 U4524 ( .A(n18123), .B(n23191), .ZN(n18438) );
  OR2_X1 U4526 ( .A1(n18907), .A2(n19568), .ZN(n2512) );
  XNOR2_X1 U4527 ( .A(n4268), .B(n18363), .ZN(n4274) );
  INV_X1 U4528 ( .A(n18520), .ZN(n16600) );
  XNOR2_X1 U4529 ( .A(n4808), .B(n17375), .ZN(n17376) );
  OR2_X1 U4530 ( .A1(n25423), .A2(n19436), .ZN(n5007) );
  AND2_X1 U4531 ( .A1(n357), .A2(n19500), .ZN(n18986) );
  XNOR2_X1 U4532 ( .A(n18175), .B(n18174), .ZN(n19520) );
  AND2_X1 U4533 ( .A1(n5572), .A2(n2626), .ZN(n20258) );
  AND2_X1 U4534 ( .A1(n19540), .A2(n19126), .ZN(n2626) );
  OR2_X1 U4535 ( .A1(n2132), .A2(n24477), .ZN(n4542) );
  XNOR2_X1 U4536 ( .A(n21164), .B(n21165), .ZN(n1605) );
  XNOR2_X1 U4537 ( .A(n4908), .B(n21532), .ZN(n17951) );
  INV_X1 U4538 ( .A(n21481), .ZN(n4908) );
  AOI21_X1 U4539 ( .B1(n22609), .B2(n22813), .A(n4272), .ZN(n22610) );
  NOR2_X1 U4540 ( .A1(n22495), .A2(n22494), .ZN(n4719) );
  OR2_X1 U4541 ( .A1(n21822), .A2(n22257), .ZN(n2987) );
  INV_X1 U4542 ( .A(n22255), .ZN(n4373) );
  OAI21_X1 U4543 ( .B1(n3741), .B2(n22811), .A(n22813), .ZN(n3740) );
  XNOR2_X1 U4544 ( .A(n20697), .B(n5286), .ZN(n20465) );
  OR2_X1 U4546 ( .A1(n6688), .A2(n4830), .ZN(n4829) );
  INV_X1 U4547 ( .A(n6648), .ZN(n7006) );
  XNOR2_X1 U4548 ( .A(Plaintext[122]), .B(Key[122]), .ZN(n6648) );
  OR2_X1 U4549 ( .A1(n6396), .A2(n6732), .ZN(n4178) );
  NAND2_X1 U4550 ( .A1(n6607), .A2(n6606), .ZN(n1926) );
  OR2_X1 U4552 ( .A1(n6528), .A2(n6529), .ZN(n4681) );
  OR2_X1 U4553 ( .A1(n6165), .A2(n7101), .ZN(n6545) );
  OR2_X1 U4554 ( .A1(n8022), .A2(n8021), .ZN(n1840) );
  OAI21_X1 U4555 ( .B1(n6094), .B2(n7006), .A(n7005), .ZN(n2879) );
  AND2_X1 U4556 ( .A1(n442), .A2(n7026), .ZN(n5089) );
  INV_X1 U4558 ( .A(n5924), .ZN(n3922) );
  AND2_X1 U4559 ( .A1(n7776), .A2(n7767), .ZN(n1786) );
  INV_X1 U4561 ( .A(n6805), .ZN(n7665) );
  INV_X1 U4562 ( .A(n8782), .ZN(n8537) );
  OR2_X1 U4563 ( .A1(n7456), .A2(n311), .ZN(n5161) );
  INV_X1 U4564 ( .A(n7257), .ZN(n7341) );
  NAND2_X1 U4565 ( .A1(n6537), .A2(n4744), .ZN(n7664) );
  INV_X1 U4566 ( .A(n8336), .ZN(n8172) );
  OR2_X1 U4567 ( .A1(n4136), .A2(n4002), .ZN(n4001) );
  NAND2_X1 U4568 ( .A1(n4883), .A2(n7068), .ZN(n2560) );
  OAI21_X1 U4569 ( .B1(n7221), .B2(n7064), .A(n431), .ZN(n4883) );
  NAND2_X1 U4570 ( .A1(n5636), .A2(n5635), .ZN(n7629) );
  NAND3_X1 U4571 ( .A1(n4377), .A2(n7538), .A3(n7539), .ZN(n9007) );
  XNOR2_X1 U4572 ( .A(n8150), .B(n5504), .ZN(n8157) );
  XNOR2_X1 U4573 ( .A(n4395), .B(n8342), .ZN(n8343) );
  XNOR2_X1 U4574 ( .A(n8612), .B(n8981), .ZN(n8889) );
  XNOR2_X1 U4575 ( .A(n7119), .B(n7120), .ZN(n9955) );
  INV_X1 U4576 ( .A(n9012), .ZN(n8665) );
  XNOR2_X1 U4577 ( .A(n8451), .B(n8454), .ZN(n1906) );
  INV_X1 U4578 ( .A(n9335), .ZN(n9334) );
  XNOR2_X1 U4579 ( .A(n8183), .B(n3507), .ZN(n3506) );
  AND2_X1 U4581 ( .A1(n25207), .A2(n10149), .ZN(n2740) );
  XNOR2_X1 U4582 ( .A(n8336), .B(n1528), .ZN(n8070) );
  INV_X1 U4584 ( .A(n9829), .ZN(n10178) );
  INV_X1 U4585 ( .A(n10614), .ZN(n10488) );
  INV_X1 U4586 ( .A(n9244), .ZN(n9866) );
  XNOR2_X1 U4587 ( .A(n9079), .B(n9078), .ZN(n10050) );
  XNOR2_X1 U4588 ( .A(n2446), .B(n8087), .ZN(n9692) );
  OR2_X1 U4589 ( .A1(n9454), .A2(n8157), .ZN(n9566) );
  OR2_X1 U4590 ( .A1(n9219), .A2(n10060), .ZN(n5608) );
  INV_X1 U4591 ( .A(n9515), .ZN(n4300) );
  AND2_X1 U4592 ( .A1(n10100), .A2(n9837), .ZN(n9327) );
  NOR2_X1 U4593 ( .A1(n10406), .A2(n10405), .ZN(n10992) );
  INV_X1 U4594 ( .A(n11036), .ZN(n5392) );
  INV_X1 U4596 ( .A(n10935), .ZN(n10508) );
  NAND3_X1 U4597 ( .A1(n1671), .A2(n1670), .A3(n1668), .ZN(n4422) );
  OR2_X1 U4598 ( .A1(n9436), .A2(n9435), .ZN(n1670) );
  NAND2_X1 U4599 ( .A1(n1669), .A2(n9434), .ZN(n1668) );
  INV_X1 U4600 ( .A(n9382), .ZN(n5105) );
  OR2_X1 U4601 ( .A1(n10172), .A2(n25), .ZN(n4212) );
  OR2_X1 U4602 ( .A1(n9815), .A2(n2207), .ZN(n2548) );
  AND3_X1 U4603 ( .A1(n10753), .A2(n2866), .A3(n2865), .ZN(n10760) );
  NAND2_X1 U4604 ( .A1(n2268), .A2(n9976), .ZN(n10416) );
  AND2_X1 U4605 ( .A1(n25499), .A2(n12942), .ZN(n2918) );
  OR2_X1 U4606 ( .A1(n3387), .A2(n10590), .ZN(n10591) );
  INV_X1 U4607 ( .A(n11704), .ZN(n3812) );
  XNOR2_X1 U4608 ( .A(n1388), .B(n12340), .ZN(n13353) );
  OAI21_X1 U4609 ( .B1(n4462), .B2(n420), .A(n4464), .ZN(n4461) );
  INV_X1 U4610 ( .A(n12613), .ZN(n3859) );
  OR2_X1 U4611 ( .A1(n10623), .A2(n11212), .ZN(n10624) );
  XNOR2_X1 U4612 ( .A(n11820), .B(n11819), .ZN(n13301) );
  INV_X1 U4613 ( .A(n405), .ZN(n4493) );
  AND2_X1 U4614 ( .A1(n13245), .A2(n13014), .ZN(n13018) );
  NOR2_X1 U4615 ( .A1(n25198), .A2(n13014), .ZN(n13016) );
  XNOR2_X1 U4616 ( .A(n11661), .B(n3208), .ZN(n11248) );
  AND2_X1 U4617 ( .A1(n13228), .A2(n11328), .ZN(n2291) );
  AND3_X1 U4618 ( .A1(n12612), .A2(n3859), .A3(n13303), .ZN(n4790) );
  OR2_X1 U4619 ( .A1(n13018), .A2(n13017), .ZN(n3558) );
  BUF_X1 U4620 ( .A(n13037), .Z(n13044) );
  OR2_X1 U4621 ( .A1(n13076), .A2(n12713), .ZN(n2192) );
  INV_X1 U4622 ( .A(n24573), .ZN(n3590) );
  AND3_X1 U4624 ( .A1(n25494), .A2(n13051), .A3(n4094), .ZN(n13086) );
  INV_X1 U4625 ( .A(n13998), .ZN(n13993) );
  INV_X1 U4626 ( .A(n12897), .ZN(n4861) );
  INV_X1 U4627 ( .A(n25248), .ZN(n2437) );
  XNOR2_X1 U4628 ( .A(n10198), .B(n10197), .ZN(n3492) );
  OAI21_X1 U4629 ( .B1(n12483), .B2(n12711), .A(n4060), .ZN(n4059) );
  AND2_X1 U4630 ( .A1(n13989), .A2(n13918), .ZN(n13984) );
  OR2_X1 U4631 ( .A1(n4729), .A2(n3766), .ZN(n2423) );
  OR2_X1 U4632 ( .A1(n12899), .A2(n13279), .ZN(n11867) );
  INV_X1 U4633 ( .A(n4241), .ZN(n12946) );
  XNOR2_X1 U4634 ( .A(n11835), .B(n11834), .ZN(n12902) );
  OR3_X1 U4635 ( .A1(n13222), .A2(n24965), .A3(n13227), .ZN(n4484) );
  INV_X1 U4636 ( .A(n14150), .ZN(n5102) );
  INV_X1 U4637 ( .A(n12767), .ZN(n2493) );
  INV_X1 U4638 ( .A(n13216), .ZN(n12986) );
  AOI22_X1 U4639 ( .A1(n13009), .A2(n11754), .B1(n13221), .B2(n12885), .ZN(
        n13010) );
  OR2_X1 U4642 ( .A1(n2608), .A2(n2837), .ZN(n12567) );
  AND2_X1 U4643 ( .A1(n13796), .A2(n13792), .ZN(n13579) );
  AND2_X1 U4644 ( .A1(n3788), .A2(n3786), .ZN(n3787) );
  OAI211_X1 U4645 ( .C1(n14268), .C2(n123), .A(n14267), .B(n3789), .ZN(n3788)
         );
  AND2_X1 U4646 ( .A1(n13884), .A2(n13597), .ZN(n13596) );
  OR2_X1 U4647 ( .A1(n12918), .A2(n24490), .ZN(n12570) );
  INV_X1 U4648 ( .A(n14048), .ZN(n14050) );
  OAI21_X1 U4649 ( .B1(n12426), .B2(n12666), .A(n10787), .ZN(n13953) );
  OR2_X1 U4650 ( .A1(n12437), .A2(n13138), .ZN(n2929) );
  OAI21_X1 U4651 ( .B1(n5013), .B2(n25061), .A(n13162), .ZN(n5012) );
  OR2_X1 U4652 ( .A1(n13164), .A2(n13163), .ZN(n4867) );
  AND2_X1 U4653 ( .A1(n4868), .A2(n14112), .ZN(n13581) );
  AND2_X1 U4654 ( .A1(n13485), .A2(n12669), .ZN(n13262) );
  OR2_X1 U4655 ( .A1(n14944), .A2(n25458), .ZN(n14144) );
  INV_X1 U4656 ( .A(n14826), .ZN(n15111) );
  INV_X1 U4657 ( .A(n13597), .ZN(n13724) );
  OR2_X1 U4658 ( .A1(n1578), .A2(n12555), .ZN(n12556) );
  AND2_X1 U4659 ( .A1(n5140), .A2(n4634), .ZN(n12072) );
  AND2_X1 U4660 ( .A1(n13325), .A2(n13323), .ZN(n5140) );
  INV_X1 U4661 ( .A(n14325), .ZN(n14330) );
  INV_X1 U4663 ( .A(n14221), .ZN(n4019) );
  INV_X1 U4664 ( .A(n13829), .ZN(n14119) );
  INV_X1 U4665 ( .A(n13966), .ZN(n13883) );
  INV_X1 U4666 ( .A(n13997), .ZN(n14235) );
  INV_X1 U4667 ( .A(n13682), .ZN(n14233) );
  AND2_X1 U4668 ( .A1(n14204), .A2(n3341), .ZN(n13814) );
  AND2_X1 U4669 ( .A1(n13446), .A2(n13445), .ZN(n2863) );
  OAI21_X1 U4670 ( .B1(n13819), .B2(n13385), .A(n13646), .ZN(n2658) );
  AND2_X1 U4671 ( .A1(n1790), .A2(n16051), .ZN(n15540) );
  OR2_X1 U4672 ( .A1(n13440), .A2(n14101), .ZN(n4598) );
  XNOR2_X1 U4673 ( .A(n14391), .B(n15452), .ZN(n15093) );
  XNOR2_X1 U4674 ( .A(n14358), .B(n14357), .ZN(n15842) );
  XNOR2_X1 U4675 ( .A(n13450), .B(n3787), .ZN(n3471) );
  XNOR2_X1 U4676 ( .A(n15177), .B(n5216), .ZN(n14964) );
  OR2_X1 U4677 ( .A1(n13676), .A2(n5221), .ZN(n13489) );
  OAI21_X1 U4678 ( .B1(n13484), .B2(n13487), .A(n3071), .ZN(n4415) );
  INV_X1 U4679 ( .A(n16368), .ZN(n15814) );
  OR2_X1 U4680 ( .A1(n15940), .A2(n2605), .ZN(n2604) );
  INV_X1 U4681 ( .A(n4765), .ZN(n14201) );
  AOI22_X1 U4683 ( .A1(n1621), .A2(n16285), .B1(n15747), .B2(n24539), .ZN(
        n17623) );
  INV_X1 U4684 ( .A(n5376), .ZN(n16622) );
  OAI21_X1 U4685 ( .B1(n16481), .B2(n15953), .A(n15696), .ZN(n5495) );
  OAI21_X1 U4686 ( .B1(n25238), .B2(n15695), .A(n16483), .ZN(n5493) );
  AND2_X1 U4687 ( .A1(n17276), .A2(n17254), .ZN(n17247) );
  AND2_X1 U4688 ( .A1(n16368), .A2(n17183), .ZN(n17181) );
  OR2_X1 U4690 ( .A1(n2549), .A2(n17442), .ZN(n16961) );
  OR2_X1 U4691 ( .A1(n17356), .A2(n17351), .ZN(n5366) );
  AND2_X1 U4692 ( .A1(n24942), .A2(n17450), .ZN(n17152) );
  INV_X1 U4693 ( .A(n3604), .ZN(n3598) );
  OAI21_X1 U4694 ( .B1(n16411), .B2(n3061), .A(n3060), .ZN(n16421) );
  INV_X1 U4695 ( .A(n17050), .ZN(n2613) );
  AND2_X1 U4697 ( .A1(n16323), .A2(n25447), .ZN(n15258) );
  AND2_X1 U4698 ( .A1(n4541), .A2(n15604), .ZN(n15693) );
  OAI22_X1 U4699 ( .A1(n4482), .A2(n17356), .B1(n16316), .B2(n367), .ZN(n16318) );
  NAND3_X1 U4700 ( .A1(n16758), .A2(n16757), .A3(n2324), .ZN(n17931) );
  OR2_X1 U4701 ( .A1(n15602), .A2(n16060), .ZN(n1673) );
  INV_X1 U4702 ( .A(n18646), .ZN(n18552) );
  NOR2_X1 U4703 ( .A1(n16671), .A2(n2530), .ZN(n2937) );
  OR2_X1 U4705 ( .A1(n16978), .A2(n17336), .ZN(n4246) );
  OR2_X1 U4706 ( .A1(n16431), .A2(n16434), .ZN(n16522) );
  NOR2_X1 U4707 ( .A1(n5522), .A2(n17572), .ZN(n3004) );
  AND2_X1 U4708 ( .A1(n1616), .A2(n1615), .ZN(n16719) );
  OR2_X1 U4709 ( .A1(n17025), .A2(n17389), .ZN(n1852) );
  OR2_X1 U4710 ( .A1(n4566), .A2(n17602), .ZN(n4565) );
  AOI21_X1 U4711 ( .B1(n4564), .B2(n4563), .A(n2968), .ZN(n4562) );
  OAI21_X1 U4712 ( .B1(n3956), .B2(n25215), .A(n3948), .ZN(n18254) );
  AOI21_X1 U4714 ( .B1(n3458), .B2(n3457), .A(n3391), .ZN(n3390) );
  AND2_X1 U4715 ( .A1(n25226), .A2(n25245), .ZN(n3391) );
  INV_X1 U4717 ( .A(n18123), .ZN(n18437) );
  INV_X1 U4718 ( .A(n19077), .ZN(n18862) );
  OR3_X1 U4719 ( .A1(n25245), .A2(n17131), .A3(n25226), .ZN(n15806) );
  OR2_X1 U4720 ( .A1(n17418), .A2(n17419), .ZN(n2054) );
  NAND2_X1 U4721 ( .A1(n2183), .A2(n2110), .ZN(n17811) );
  AND2_X1 U4722 ( .A1(n17198), .A2(n17395), .ZN(n2112) );
  XNOR2_X1 U4723 ( .A(n18397), .B(n17520), .ZN(n18627) );
  OAI21_X1 U4724 ( .B1(n17461), .B2(n288), .A(n17464), .ZN(n5158) );
  XNOR2_X1 U4725 ( .A(n3703), .B(n18187), .ZN(n18291) );
  AOI22_X1 U4726 ( .A1(n3930), .A2(n16985), .B1(n3929), .B2(n17144), .ZN(n3928) );
  OR2_X1 U4727 ( .A1(n3432), .A2(n17053), .ZN(n3431) );
  OR2_X1 U4728 ( .A1(n16895), .A2(n2372), .ZN(n2373) );
  AOI21_X1 U4729 ( .B1(n5386), .B2(n17479), .A(n2181), .ZN(n2374) );
  INV_X1 U4730 ( .A(n16513), .ZN(n16618) );
  OR2_X1 U4731 ( .A1(n16703), .A2(n16705), .ZN(n16617) );
  XNOR2_X1 U4732 ( .A(n24536), .B(n17757), .ZN(n18363) );
  NAND2_X1 U4733 ( .A1(n4304), .A2(n16908), .ZN(n2583) );
  NAND3_X1 U4734 ( .A1(n16182), .A2(n16181), .A3(n5017), .ZN(n17863) );
  AND2_X1 U4735 ( .A1(n16984), .A2(n16985), .ZN(n2161) );
  AND2_X1 U4736 ( .A1(n17122), .A2(n17114), .ZN(n16801) );
  AND2_X1 U4737 ( .A1(n25422), .A2(n19436), .ZN(n3985) );
  NOR2_X1 U4738 ( .A1(n1427), .A2(n5573), .ZN(n5569) );
  INV_X1 U4739 ( .A(n20192), .ZN(n5208) );
  XNOR2_X1 U4740 ( .A(n21160), .B(n21750), .ZN(n21163) );
  XNOR2_X1 U4741 ( .A(n21266), .B(n21160), .ZN(n21611) );
  OAI211_X1 U4742 ( .C1(n20220), .C2(n20510), .A(n1809), .B(n1808), .ZN(n21495) );
  INV_X1 U4743 ( .A(n19710), .ZN(n4713) );
  OAI22_X1 U4748 ( .A1(n5499), .A2(n25345), .B1(n2606), .B2(n20214), .ZN(
        n20513) );
  NAND2_X1 U4750 ( .A1(n20207), .A2(n4264), .ZN(n4263) );
  AND2_X1 U4751 ( .A1(n20206), .A2(n4265), .ZN(n4264) );
  OR2_X1 U4753 ( .A1(n20548), .A2(n20124), .ZN(n4569) );
  INV_X1 U4754 ( .A(n22721), .ZN(n2711) );
  INV_X1 U4755 ( .A(n20336), .ZN(n19708) );
  INV_X1 U4756 ( .A(n20459), .ZN(n4489) );
  OAI22_X1 U4757 ( .A1(n20128), .A2(n20130), .B1(n20130), .B2(n20129), .ZN(
        n5491) );
  AND2_X1 U4758 ( .A1(n21523), .A2(n2563), .ZN(n20926) );
  INV_X1 U4759 ( .A(n3115), .ZN(n2563) );
  NOR2_X1 U4761 ( .A1(n19984), .A2(n19983), .ZN(n2098) );
  OR2_X1 U4762 ( .A1(n20117), .A2(n20116), .ZN(n2873) );
  OR2_X1 U4763 ( .A1(n20114), .A2(n20111), .ZN(n2874) );
  XNOR2_X1 U4764 ( .A(n21599), .B(n21520), .ZN(n21192) );
  XNOR2_X1 U4765 ( .A(n21550), .B(n21981), .ZN(n21209) );
  NOR2_X1 U4766 ( .A1(n25383), .A2(n2431), .ZN(n20375) );
  OR2_X1 U4767 ( .A1(n20374), .A2(n2432), .ZN(n2431) );
  OR2_X1 U4768 ( .A1(n19682), .A2(n20302), .ZN(n2135) );
  NAND3_X1 U4770 ( .A1(n19986), .A2(n19987), .A3(n21068), .ZN(n3963) );
  XNOR2_X1 U4772 ( .A(n22006), .B(n25400), .ZN(n4396) );
  XNOR2_X1 U4773 ( .A(n2465), .B(n25483), .ZN(n20745) );
  XNOR2_X1 U4774 ( .A(n21699), .B(n23183), .ZN(n2465) );
  INV_X1 U4775 ( .A(n329), .ZN(n5224) );
  XNOR2_X1 U4776 ( .A(n20972), .B(n20678), .ZN(n4100) );
  NOR2_X1 U4777 ( .A1(n22209), .A2(n22064), .ZN(n22092) );
  XNOR2_X1 U4778 ( .A(n21724), .B(n21723), .ZN(n2633) );
  XNOR2_X1 U4781 ( .A(n21737), .B(n21734), .ZN(n4687) );
  OR2_X1 U4782 ( .A1(n23016), .A2(n23014), .ZN(n22914) );
  XNOR2_X1 U4783 ( .A(n20918), .B(n1628), .ZN(n2315) );
  INV_X1 U4784 ( .A(n21538), .ZN(n1628) );
  INV_X1 U4785 ( .A(n22227), .ZN(n3231) );
  OR2_X1 U4786 ( .A1(n22228), .A2(n22231), .ZN(n3230) );
  XNOR2_X1 U4787 ( .A(n20324), .B(n3746), .ZN(n4169) );
  OR2_X1 U4788 ( .A1(n22770), .A2(n5378), .ZN(n5377) );
  INV_X1 U4789 ( .A(n22812), .ZN(n4469) );
  OR2_X1 U4790 ( .A1(n5712), .A2(n21856), .ZN(n22772) );
  NAND4_X1 U4794 ( .A1(n23202), .A2(n22569), .A3(n24889), .A4(n22561), .ZN(
        n4237) );
  AND2_X1 U4795 ( .A1(n23805), .A2(n24895), .ZN(n2591) );
  INV_X1 U4797 ( .A(n3856), .ZN(n19625) );
  INV_X1 U4798 ( .A(n23843), .ZN(n23862) );
  INV_X1 U4799 ( .A(n6733), .ZN(n2119) );
  XNOR2_X1 U4800 ( .A(n5847), .B(Key[161]), .ZN(n6770) );
  OR2_X1 U4801 ( .A1(n6297), .A2(n6438), .ZN(n5946) );
  AOI21_X1 U4802 ( .B1(n6703), .B2(n24405), .A(n6959), .ZN(n4324) );
  INV_X1 U4803 ( .A(n8021), .ZN(n7531) );
  OR2_X1 U4804 ( .A1(n6162), .A2(n6265), .ZN(n2534) );
  OR2_X1 U4805 ( .A1(n5910), .A2(n5887), .ZN(n4503) );
  OAI21_X1 U4807 ( .B1(n6771), .B2(n24037), .A(n6770), .ZN(n6772) );
  INV_X1 U4808 ( .A(n4672), .ZN(n7945) );
  OR2_X1 U4809 ( .A1(n7858), .A2(n7857), .ZN(n4976) );
  INV_X1 U4810 ( .A(n7413), .ZN(n4827) );
  NOR2_X1 U4811 ( .A1(n5824), .A2(n6473), .ZN(n6899) );
  OAI21_X1 U4812 ( .B1(n5975), .B2(n6987), .A(n5974), .ZN(n5978) );
  AND2_X1 U4813 ( .A1(n5798), .A2(n5799), .ZN(n7481) );
  OR2_X1 U4814 ( .A1(n7861), .A2(n7862), .ZN(n3571) );
  INV_X1 U4815 ( .A(n7781), .ZN(n7419) );
  AND3_X1 U4816 ( .A1(n3588), .A2(n3344), .A3(n7531), .ZN(n3587) );
  AND2_X1 U4817 ( .A1(n4708), .A2(n4711), .ZN(n4707) );
  AND3_X1 U4818 ( .A1(n7930), .A2(n7931), .A3(n7929), .ZN(n4545) );
  INV_X1 U4819 ( .A(n2402), .ZN(n8024) );
  OR2_X1 U4820 ( .A1(n6768), .A2(n6767), .ZN(n2976) );
  INV_X1 U4821 ( .A(n7335), .ZN(n7592) );
  OR2_X1 U4823 ( .A1(n6494), .A2(n6493), .ZN(n1575) );
  OAI211_X1 U4825 ( .C1(n1468), .C2(n4376), .A(n7079), .B(n4375), .ZN(n8452)
         );
  OR2_X1 U4826 ( .A1(n6040), .A2(n6165), .ZN(n6041) );
  INV_X1 U4827 ( .A(n8960), .ZN(n8908) );
  OAI211_X1 U4828 ( .C1(n6752), .C2(n6674), .A(n6578), .B(n1807), .ZN(n2495)
         );
  OR2_X1 U4829 ( .A1(n6400), .A2(n6757), .ZN(n1807) );
  INV_X1 U4830 ( .A(n6572), .ZN(n6058) );
  OR2_X1 U4831 ( .A1(n6059), .A2(n6967), .ZN(n3838) );
  AND2_X1 U4832 ( .A1(n2355), .A2(n1175), .ZN(n2349) );
  INV_X1 U4833 ( .A(n6314), .ZN(n5452) );
  OR2_X1 U4834 ( .A1(n6233), .A2(n6715), .ZN(n6110) );
  XNOR2_X1 U4835 ( .A(n8721), .B(n2272), .ZN(n8756) );
  INV_X1 U4836 ( .A(n8755), .ZN(n2272) );
  OAI21_X1 U4837 ( .B1(n7045), .B2(n7174), .A(n3496), .ZN(n8812) );
  OAI21_X1 U4838 ( .B1(n5606), .B2(n5605), .A(n5607), .ZN(n5603) );
  AND2_X1 U4839 ( .A1(n7157), .A2(n7156), .ZN(n5345) );
  INV_X1 U4840 ( .A(n7364), .ZN(n7911) );
  INV_X1 U4841 ( .A(n7629), .ZN(n7910) );
  INV_X1 U4842 ( .A(n3979), .ZN(n8371) );
  OR2_X1 U4843 ( .A1(n6413), .A2(n7721), .ZN(n1879) );
  OR2_X1 U4844 ( .A1(n7115), .A2(n7761), .ZN(n5691) );
  INV_X1 U4845 ( .A(n2145), .ZN(n5690) );
  INV_X1 U4847 ( .A(n6549), .ZN(n7671) );
  AND2_X1 U4848 ( .A1(n3680), .A2(n7541), .ZN(n3679) );
  XNOR2_X1 U4849 ( .A(n8796), .B(n8795), .ZN(n9137) );
  XNOR2_X1 U4850 ( .A(n9007), .B(n2560), .ZN(n9115) );
  INV_X1 U4851 ( .A(n7553), .ZN(n2323) );
  OAI22_X1 U4852 ( .A1(n7043), .A2(n3730), .B1(n9355), .B2(n7044), .ZN(n4481)
         );
  OR2_X1 U4854 ( .A1(n7073), .A2(n437), .ZN(n3814) );
  XNOR2_X1 U4855 ( .A(n4802), .B(n8691), .ZN(n8994) );
  OR2_X1 U4856 ( .A1(n7909), .A2(n7364), .ZN(n4825) );
  XNOR2_X1 U4857 ( .A(n8237), .B(n3715), .ZN(n4913) );
  XNOR2_X1 U4858 ( .A(n4378), .B(n8639), .ZN(n9111) );
  INV_X1 U4859 ( .A(n10186), .ZN(n9520) );
  OAI21_X1 U4860 ( .B1(n9717), .B2(n9716), .A(n9715), .ZN(n10533) );
  AND2_X1 U4861 ( .A1(n9713), .A2(n10037), .ZN(n1669) );
  INV_X1 U4863 ( .A(n9702), .ZN(n4656) );
  AND2_X1 U4864 ( .A1(n3762), .A2(n10571), .ZN(n3758) );
  AND2_X1 U4865 ( .A1(n10942), .A2(n5392), .ZN(n3761) );
  INV_X1 U4866 ( .A(n9355), .ZN(n3730) );
  AND2_X1 U4867 ( .A1(n10848), .A2(n10850), .ZN(n5077) );
  INV_X1 U4868 ( .A(n11121), .ZN(n10460) );
  AND2_X1 U4869 ( .A1(n10682), .A2(n11004), .ZN(n11006) );
  AND2_X1 U4870 ( .A1(n9673), .A2(n5279), .ZN(n1532) );
  INV_X1 U4871 ( .A(n9795), .ZN(n5279) );
  INV_X1 U4873 ( .A(n11190), .ZN(n10480) );
  OAI21_X1 U4874 ( .B1(n1519), .B2(n2294), .A(n4993), .ZN(n1518) );
  OAI21_X1 U4875 ( .B1(n9693), .B2(n9876), .A(n9692), .ZN(n1520) );
  OR2_X1 U4876 ( .A1(n9664), .A2(n9985), .ZN(n2011) );
  INV_X1 U4877 ( .A(n9737), .ZN(n9982) );
  OR2_X1 U4880 ( .A1(n8526), .A2(n9334), .ZN(n2046) );
  AND2_X1 U4881 ( .A1(n9838), .A2(n428), .ZN(n9517) );
  INV_X1 U4882 ( .A(n10482), .ZN(n10457) );
  INV_X1 U4883 ( .A(n12147), .ZN(n12282) );
  OR2_X1 U4885 ( .A1(n10489), .A2(n10617), .ZN(n5062) );
  OR2_X1 U4887 ( .A1(n2148), .A2(n10985), .ZN(n11164) );
  OR2_X1 U4889 ( .A1(n10283), .A2(n10190), .ZN(n2226) );
  AND2_X1 U4890 ( .A1(n5393), .A2(n5392), .ZN(n5391) );
  OR2_X1 U4891 ( .A1(n10620), .A2(n233), .ZN(n3724) );
  AND2_X1 U4892 ( .A1(n2849), .A2(n10218), .ZN(n10219) );
  XNOR2_X1 U4893 ( .A(n2917), .B(n12023), .ZN(n12181) );
  AND2_X1 U4894 ( .A1(n11122), .A2(n10722), .ZN(n10723) );
  OR2_X1 U4895 ( .A1(n10936), .A2(n10935), .ZN(n2307) );
  OR2_X1 U4896 ( .A1(n5296), .A2(n2311), .ZN(n2310) );
  OR2_X1 U4897 ( .A1(n10549), .A2(n10699), .ZN(n4758) );
  OR2_X1 U4899 ( .A1(n2584), .A2(n10596), .ZN(n10600) );
  OR2_X1 U4900 ( .A1(n301), .A2(n2295), .ZN(n5312) );
  XNOR2_X1 U4901 ( .A(n11567), .B(n11566), .ZN(n12520) );
  INV_X1 U4902 ( .A(n12396), .ZN(n3269) );
  OR2_X1 U4903 ( .A1(n3573), .A2(n11069), .ZN(n10348) );
  INV_X1 U4904 ( .A(n11295), .ZN(n3448) );
  XNOR2_X1 U4905 ( .A(n11385), .B(n11653), .ZN(n11848) );
  NAND2_X1 U4906 ( .A1(n10659), .A2(n10660), .ZN(n2450) );
  INV_X1 U4907 ( .A(n12167), .ZN(n11486) );
  XNOR2_X1 U4908 ( .A(n12381), .B(n12048), .ZN(n11812) );
  OR2_X1 U4909 ( .A1(n11050), .A2(n11051), .ZN(n3144) );
  INV_X1 U4910 ( .A(n11787), .ZN(n12081) );
  OR2_X1 U4911 ( .A1(n10293), .A2(n11129), .ZN(n10295) );
  XNOR2_X1 U4912 ( .A(n4670), .B(n23476), .ZN(n11225) );
  AND2_X1 U4913 ( .A1(n14141), .A2(n14143), .ZN(n2178) );
  INV_X1 U4914 ( .A(n403), .ZN(n3974) );
  AOI21_X1 U4915 ( .B1(n13178), .B2(n24499), .A(n3968), .ZN(n3975) );
  OR2_X1 U4916 ( .A1(n12469), .A2(n12470), .ZN(n4336) );
  INV_X1 U4917 ( .A(n12470), .ZN(n13066) );
  OR2_X1 U4918 ( .A1(n13234), .A2(n13298), .ZN(n2544) );
  AND2_X1 U4919 ( .A1(n14124), .A2(n14208), .ZN(n13813) );
  INV_X1 U4920 ( .A(n13843), .ZN(n14067) );
  OR2_X1 U4921 ( .A1(n14294), .A2(n13907), .ZN(n11369) );
  OR2_X1 U4922 ( .A1(n13568), .A2(n13569), .ZN(n2603) );
  NOR2_X1 U4923 ( .A1(n14017), .A2(n2573), .ZN(n14020) );
  AND2_X1 U4924 ( .A1(n14089), .A2(n13533), .ZN(n2573) );
  INV_X1 U4925 ( .A(n13901), .ZN(n13959) );
  INV_X1 U4927 ( .A(n14301), .ZN(n3966) );
  OAI211_X1 U4928 ( .C1(n13591), .C2(n13864), .A(n2417), .B(n5150), .ZN(n14698) );
  OR2_X1 U4929 ( .A1(n12803), .A2(n298), .ZN(n2417) );
  AND2_X1 U4931 ( .A1(n14321), .A2(n3401), .ZN(n13500) );
  XNOR2_X1 U4932 ( .A(n15005), .B(n1907), .ZN(n13524) );
  INV_X1 U4933 ( .A(n15476), .ZN(n1907) );
  OR2_X1 U4934 ( .A1(n13807), .A2(n3717), .ZN(n13515) );
  OR2_X1 U4935 ( .A1(n4452), .A2(n14165), .ZN(n4451) );
  OAI211_X1 U4936 ( .C1(n4763), .C2(n14166), .A(n14170), .B(n4762), .ZN(n14697) );
  OR2_X1 U4937 ( .A1(n14171), .A2(n14172), .ZN(n4762) );
  AND2_X1 U4938 ( .A1(n14268), .A2(n14269), .ZN(n12542) );
  OR2_X1 U4939 ( .A1(n14226), .A2(n14225), .ZN(n1747) );
  NOR2_X1 U4941 ( .A1(n14000), .A2(n12669), .ZN(n14004) );
  AND2_X1 U4943 ( .A1(n14102), .A2(n14216), .ZN(n4876) );
  INV_X1 U4944 ( .A(n14102), .ZN(n4877) );
  AND2_X1 U4945 ( .A1(n2570), .A2(n3888), .ZN(n14202) );
  OR2_X1 U4946 ( .A1(n3338), .A2(n12639), .ZN(n4765) );
  OR2_X1 U4947 ( .A1(n13701), .A2(n13923), .ZN(n13707) );
  AND2_X1 U4948 ( .A1(n13995), .A2(n25435), .ZN(n14236) );
  OAI21_X1 U4949 ( .B1(n3808), .B2(n3807), .A(n13712), .ZN(n11681) );
  INV_X1 U4952 ( .A(n2242), .ZN(n3233) );
  OR2_X1 U4954 ( .A1(n14334), .A2(n14336), .ZN(n3059) );
  XNOR2_X1 U4955 ( .A(n13906), .B(n5251), .ZN(n15411) );
  INV_X1 U4956 ( .A(n14940), .ZN(n4557) );
  OAI21_X1 U4957 ( .B1(n24152), .B2(n14306), .A(n12120), .ZN(n12176) );
  NAND2_X1 U4958 ( .A1(n13525), .A2(n13864), .ZN(n2507) );
  AND2_X1 U4959 ( .A1(n3777), .A2(n3776), .ZN(n14437) );
  XNOR2_X1 U4960 ( .A(n15111), .B(n15112), .ZN(n15114) );
  AND2_X1 U4961 ( .A1(n4382), .A2(n4383), .ZN(n13263) );
  OR2_X1 U4963 ( .A1(n4016), .A2(n2457), .ZN(n4015) );
  XNOR2_X1 U4964 ( .A(n4637), .B(n4635), .ZN(n4897) );
  INV_X1 U4965 ( .A(n2375), .ZN(n16050) );
  INV_X1 U4966 ( .A(n14915), .ZN(n4095) );
  NOR2_X1 U4967 ( .A1(n11806), .A2(n13966), .ZN(n13470) );
  OR2_X1 U4968 ( .A1(n13968), .A2(n13969), .ZN(n3802) );
  OR2_X1 U4969 ( .A1(n4019), .A2(n14219), .ZN(n13831) );
  AOI21_X1 U4970 ( .B1(n2170), .B2(n2172), .A(n1868), .ZN(n1867) );
  OAI211_X1 U4971 ( .C1(n14107), .C2(n14112), .A(n14109), .B(n13582), .ZN(
        n3983) );
  XNOR2_X1 U4972 ( .A(n15071), .B(n14594), .ZN(n14389) );
  OR2_X1 U4973 ( .A1(n14144), .A2(n3887), .ZN(n3678) );
  XNOR2_X1 U4974 ( .A(n14902), .B(n14936), .ZN(n4966) );
  OAI21_X1 U4975 ( .B1(n3756), .B2(n13843), .A(n300), .ZN(n3755) );
  AOI22_X1 U4976 ( .A1(n13597), .A2(n13966), .B1(n11806), .B2(n13969), .ZN(
        n13598) );
  OAI211_X1 U4977 ( .C1(n14123), .C2(n13814), .A(n13548), .B(n14122), .ZN(
        n2382) );
  XNOR2_X1 U4978 ( .A(n15062), .B(n15133), .ZN(n15462) );
  XNOR2_X1 U4979 ( .A(n15119), .B(n14775), .ZN(n15461) );
  AOI21_X1 U4980 ( .B1(n13477), .B2(n14141), .A(n14140), .ZN(n5297) );
  INV_X1 U4981 ( .A(n14141), .ZN(n5299) );
  INV_X1 U4982 ( .A(n16095), .ZN(n1762) );
  XNOR2_X1 U4984 ( .A(n13441), .B(n4582), .ZN(n4581) );
  OR2_X1 U4985 ( .A1(n16410), .A2(n16414), .ZN(n3061) );
  OR2_X1 U4986 ( .A1(n15583), .A2(n16100), .ZN(n5245) );
  AND2_X1 U4987 ( .A1(n17275), .A2(n17273), .ZN(n2511) );
  OR2_X1 U4989 ( .A1(n16225), .A2(n24506), .ZN(n5383) );
  OR2_X1 U4990 ( .A1(n2587), .A2(n16796), .ZN(n5243) );
  AND2_X1 U4991 ( .A1(n15953), .A2(n16480), .ZN(n4773) );
  AND2_X1 U4993 ( .A1(n17326), .A2(n17265), .ZN(n17266) );
  OR2_X1 U4994 ( .A1(n16324), .A2(n16323), .ZN(n15899) );
  INV_X1 U4995 ( .A(n17015), .ZN(n17214) );
  OR2_X1 U4996 ( .A1(n17324), .A2(n17326), .ZN(n3991) );
  INV_X1 U4997 ( .A(n16892), .ZN(n16893) );
  INV_X1 U5000 ( .A(n15612), .ZN(n15856) );
  INV_X1 U5001 ( .A(n15611), .ZN(n16117) );
  OR2_X1 U5002 ( .A1(n16118), .A2(n15804), .ZN(n2518) );
  AND2_X1 U5003 ( .A1(n17435), .A2(n17434), .ZN(n16429) );
  AND2_X1 U5004 ( .A1(n17421), .A2(n17381), .ZN(n17426) );
  OR2_X1 U5005 ( .A1(n17185), .A2(n25465), .ZN(n17025) );
  OR2_X1 U5006 ( .A1(n17123), .A2(n4664), .ZN(n4663) );
  INV_X1 U5007 ( .A(n1896), .ZN(n4664) );
  NOR2_X1 U5009 ( .A1(n17282), .A2(n17254), .ZN(n4941) );
  INV_X1 U5010 ( .A(n5018), .ZN(n16662) );
  OR2_X1 U5012 ( .A1(n3955), .A2(n370), .ZN(n3953) );
  NAND3_X1 U5013 ( .A1(n2265), .A2(n16953), .A3(n2264), .ZN(n17791) );
  INV_X1 U5014 ( .A(n17532), .ZN(n18293) );
  AND2_X1 U5015 ( .A1(n17618), .A2(n17617), .ZN(n18018) );
  OR2_X1 U5016 ( .A1(n17457), .A2(n5073), .ZN(n17459) );
  XNOR2_X1 U5017 ( .A(n17724), .B(n17725), .ZN(n18812) );
  OAI21_X1 U5018 ( .B1(n3602), .B2(n17391), .A(n17388), .ZN(n3601) );
  NOR2_X1 U5019 ( .A1(n17186), .A2(n3317), .ZN(n3603) );
  XNOR2_X1 U5020 ( .A(n24888), .B(n18275), .ZN(n18475) );
  INV_X1 U5021 ( .A(n19445), .ZN(n19449) );
  OR2_X1 U5022 ( .A1(n16740), .A2(n17084), .ZN(n4614) );
  OR2_X1 U5024 ( .A1(n16557), .A2(n17211), .ZN(n16259) );
  XNOR2_X1 U5026 ( .A(n17709), .B(n18466), .ZN(n17882) );
  AND2_X1 U5027 ( .A1(n17312), .A2(n17305), .ZN(n3626) );
  INV_X1 U5028 ( .A(n18812), .ZN(n19390) );
  AND2_X1 U5029 ( .A1(n17524), .A2(n17171), .ZN(n16823) );
  XNOR2_X1 U5030 ( .A(n3706), .B(n18660), .ZN(n2692) );
  AND2_X1 U5031 ( .A1(n17575), .A2(n17574), .ZN(n1637) );
  AOI21_X1 U5032 ( .B1(n1640), .B2(n1639), .A(n17574), .ZN(n1638) );
  XNOR2_X1 U5033 ( .A(n17970), .B(n17811), .ZN(n18463) );
  INV_X1 U5035 ( .A(n18128), .ZN(n18371) );
  INV_X1 U5037 ( .A(n18448), .ZN(n3197) );
  OR2_X1 U5038 ( .A1(n19088), .A2(n19419), .ZN(n19089) );
  OR2_X1 U5039 ( .A1(n16630), .A2(n16629), .ZN(n16631) );
  XNOR2_X1 U5040 ( .A(n18257), .B(n18256), .ZN(n19278) );
  INV_X1 U5041 ( .A(n19470), .ZN(n3748) );
  XNOR2_X1 U5042 ( .A(n2283), .B(n18388), .ZN(n18458) );
  OR2_X1 U5043 ( .A1(n16734), .A2(n17067), .ZN(n5674) );
  XNOR2_X1 U5044 ( .A(n18227), .B(n18293), .ZN(n17679) );
  XNOR2_X1 U5045 ( .A(n17112), .B(n17113), .ZN(n17496) );
  OR2_X1 U5046 ( .A1(n16845), .A2(n2064), .ZN(n5136) );
  XNOR2_X1 U5047 ( .A(n18559), .B(n23151), .ZN(n2334) );
  XNOR2_X1 U5048 ( .A(n17673), .B(n2332), .ZN(n19488) );
  INV_X1 U5049 ( .A(n20386), .ZN(n19345) );
  NOR2_X1 U5051 ( .A1(n19361), .A2(n19210), .ZN(n4853) );
  OR2_X1 U5052 ( .A1(n18998), .A2(n19420), .ZN(n19088) );
  OAI21_X1 U5053 ( .B1(n19426), .B2(n19760), .A(n2663), .ZN(n19761) );
  INV_X1 U5054 ( .A(n19302), .ZN(n18766) );
  AND2_X1 U5055 ( .A1(n19413), .A2(n19408), .ZN(n1890) );
  AND2_X1 U5056 ( .A1(n2216), .A2(n19376), .ZN(n2410) );
  BUF_X1 U5057 ( .A(n19021), .Z(n17762) );
  OR2_X1 U5058 ( .A1(n19460), .A2(n18976), .ZN(n18978) );
  OR2_X1 U5059 ( .A1(n20536), .A2(n20145), .ZN(n20146) );
  OR2_X1 U5060 ( .A1(n18851), .A2(n19479), .ZN(n4403) );
  OR2_X1 U5061 ( .A1(n17554), .A2(n19272), .ZN(n4916) );
  OR2_X1 U5062 ( .A1(n19539), .A2(n3773), .ZN(n3751) );
  OR2_X1 U5063 ( .A1(n19520), .A2(n19522), .ZN(n18206) );
  AND2_X1 U5064 ( .A1(n19568), .A2(n19570), .ZN(n3995) );
  OAI21_X1 U5065 ( .B1(n19570), .B2(n19191), .A(n19192), .ZN(n3996) );
  OAI21_X1 U5066 ( .B1(n19106), .B2(n19105), .A(n2464), .ZN(n2462) );
  INV_X1 U5067 ( .A(n19799), .ZN(n1522) );
  INV_X1 U5068 ( .A(n19128), .ZN(n18767) );
  INV_X1 U5069 ( .A(n18790), .ZN(n19400) );
  INV_X1 U5070 ( .A(n19522), .ZN(n18895) );
  INV_X1 U5072 ( .A(n19304), .ZN(n18947) );
  AND2_X1 U5074 ( .A1(n19531), .A2(n24329), .ZN(n19535) );
  AND2_X1 U5075 ( .A1(n19579), .A2(n19580), .ZN(n2069) );
  XNOR2_X1 U5076 ( .A(n18066), .B(n18065), .ZN(n19077) );
  INV_X1 U5077 ( .A(n19311), .ZN(n5371) );
  XNOR2_X1 U5078 ( .A(n17008), .B(n17007), .ZN(n19312) );
  XNOR2_X1 U5079 ( .A(n5302), .B(n5305), .ZN(n5301) );
  XNOR2_X1 U5080 ( .A(n17033), .B(n3534), .ZN(n17034) );
  AND2_X1 U5081 ( .A1(n20598), .A2(n20599), .ZN(n19740) );
  OR2_X1 U5082 ( .A1(n25223), .A2(n20215), .ZN(n2606) );
  XNOR2_X1 U5083 ( .A(n2569), .B(n25222), .ZN(n21494) );
  XNOR2_X1 U5084 ( .A(n21501), .B(n21500), .ZN(n21502) );
  INV_X1 U5085 ( .A(n20533), .ZN(n20539) );
  INV_X1 U5088 ( .A(n18729), .ZN(n19228) );
  AND2_X1 U5089 ( .A1(n20111), .A2(n20109), .ZN(n3326) );
  AND2_X1 U5091 ( .A1(n19658), .A2(n3240), .ZN(n3241) );
  OR2_X1 U5093 ( .A1(n18783), .A2(n19407), .ZN(n5670) );
  OR2_X1 U5094 ( .A1(n20016), .A2(n20137), .ZN(n19994) );
  INV_X1 U5095 ( .A(n19917), .ZN(n20117) );
  AND2_X1 U5096 ( .A1(n18994), .A2(n20319), .ZN(n19691) );
  OR2_X1 U5098 ( .A1(n5189), .A2(n2024), .ZN(n5185) );
  AND2_X1 U5099 ( .A1(n20960), .A2(n20451), .ZN(n1614) );
  XNOR2_X1 U5100 ( .A(n21573), .B(n21721), .ZN(n21217) );
  OAI21_X1 U5101 ( .B1(n22465), .B2(n22462), .A(n22464), .ZN(n3906) );
  INV_X1 U5102 ( .A(n24042), .ZN(n2679) );
  OR2_X1 U5103 ( .A1(n20446), .A2(n20447), .ZN(n3075) );
  OR2_X1 U5105 ( .A1(n22421), .A2(n2674), .ZN(n2671) );
  OR2_X1 U5106 ( .A1(n22887), .A2(n22728), .ZN(n3836) );
  XNOR2_X1 U5107 ( .A(n21608), .B(n20826), .ZN(n20881) );
  OR2_X1 U5108 ( .A1(n22241), .A2(n22242), .ZN(n2753) );
  AOI21_X2 U5109 ( .B1(n2356), .B2(n19156), .A(n2358), .ZN(n21266) );
  INV_X1 U5110 ( .A(n20697), .ZN(n21325) );
  NOR2_X1 U5111 ( .A1(n22656), .A2(n25241), .ZN(n3741) );
  INV_X1 U5112 ( .A(n1605), .ZN(n2393) );
  NOR2_X1 U5113 ( .A1(n22592), .A2(n1605), .ZN(n22590) );
  AND2_X1 U5114 ( .A1(n25066), .A2(n2393), .ZN(n21188) );
  OAI21_X1 U5116 ( .B1(n2828), .B2(n21368), .A(n5539), .ZN(n22511) );
  AND2_X1 U5117 ( .A1(n25471), .A2(n22590), .ZN(n22318) );
  OR2_X1 U5118 ( .A1(n24971), .A2(n1593), .ZN(n21936) );
  NOR2_X1 U5119 ( .A1(n21883), .A2(n22401), .ZN(n22263) );
  AND2_X1 U5120 ( .A1(n22335), .A2(n22338), .ZN(n4442) );
  AND2_X1 U5121 ( .A1(n22268), .A2(n22396), .ZN(n3781) );
  NOR2_X1 U5122 ( .A1(n4098), .A2(n22975), .ZN(n4372) );
  NOR2_X1 U5124 ( .A1(n22198), .A2(n23574), .ZN(n23573) );
  OR2_X1 U5125 ( .A1(n22166), .A2(n22072), .ZN(n1679) );
  AND2_X1 U5126 ( .A1(n22911), .A2(n23464), .ZN(n2691) );
  INV_X1 U5127 ( .A(n22072), .ZN(n4064) );
  OR2_X1 U5128 ( .A1(n22092), .A2(n22156), .ZN(n22067) );
  XNOR2_X1 U5129 ( .A(n20835), .B(n20834), .ZN(n23575) );
  INV_X1 U5132 ( .A(n21903), .ZN(n2477) );
  OR2_X1 U5133 ( .A1(n24895), .A2(n23002), .ZN(n21902) );
  INV_X1 U5134 ( .A(n24895), .ZN(n4533) );
  OAI21_X1 U5135 ( .B1(n4473), .B2(n22812), .A(n4471), .ZN(n22826) );
  OR2_X1 U5136 ( .A1(n22658), .A2(n4469), .ZN(n4471) );
  OR2_X1 U5137 ( .A1(n23480), .A2(n23481), .ZN(n2539) );
  OR2_X1 U5138 ( .A1(n23053), .A2(n23048), .ZN(n3909) );
  NAND2_X1 U5139 ( .A1(n23042), .A2(n3913), .ZN(n3912) );
  AND2_X1 U5140 ( .A1(n23049), .A2(n23048), .ZN(n3913) );
  OR2_X1 U5141 ( .A1(n21930), .A2(n22464), .ZN(n21931) );
  AND2_X1 U5142 ( .A1(n5084), .A2(n22400), .ZN(n21915) );
  INV_X1 U5143 ( .A(n4236), .ZN(n4233) );
  INV_X1 U5144 ( .A(Key[58]), .ZN(n4236) );
  NOR2_X1 U5145 ( .A1(n21924), .A2(n2376), .ZN(n21925) );
  AOI22_X1 U5146 ( .A1(n1440), .A2(n22326), .B1(n21918), .B2(n5224), .ZN(n5223) );
  OAI22_X1 U5147 ( .A1(n22284), .A2(n2904), .B1(n22563), .B2(n22285), .ZN(
        n22287) );
  INV_X1 U5148 ( .A(n22563), .ZN(n2904) );
  NOR2_X1 U5149 ( .A1(n25550), .A2(n23277), .ZN(n22536) );
  INV_X1 U5150 ( .A(n23317), .ZN(n23318) );
  OAI21_X1 U5151 ( .B1(n22863), .B2(n22862), .A(n23462), .ZN(n1799) );
  OR2_X1 U5152 ( .A1(n22858), .A2(n22857), .ZN(n3264) );
  OAI21_X1 U5153 ( .B1(n23443), .B2(n22527), .A(n5348), .ZN(n22529) );
  OR2_X1 U5154 ( .A1(n23443), .A2(n1370), .ZN(n4033) );
  INV_X1 U5155 ( .A(n2710), .ZN(n23491) );
  AOI21_X1 U5156 ( .B1(n2313), .B2(n22206), .A(n22209), .ZN(n5226) );
  AOI21_X1 U5157 ( .B1(n22156), .B2(n22159), .A(n22092), .ZN(n5227) );
  INV_X1 U5158 ( .A(n22208), .ZN(n2313) );
  NOR2_X1 U5159 ( .A1(n22058), .A2(n22228), .ZN(n4398) );
  INV_X1 U5160 ( .A(n3227), .ZN(n3226) );
  AND2_X1 U5161 ( .A1(n23853), .A2(n24469), .ZN(n3737) );
  OR2_X1 U5162 ( .A1(n3641), .A2(n23998), .ZN(n3640) );
  NOR2_X1 U5164 ( .A1(n22810), .A2(n22813), .ZN(n4468) );
  OR2_X1 U5165 ( .A1(n24012), .A2(n24006), .ZN(n3486) );
  OR2_X1 U5166 ( .A1(n6752), .A2(n6675), .ZN(n6753) );
  OR2_X1 U5167 ( .A1(n6758), .A2(n6757), .ZN(n3276) );
  AND2_X1 U5169 ( .A1(n6776), .A2(n6198), .ZN(n4078) );
  OR2_X1 U5170 ( .A1(n6679), .A2(n6944), .ZN(n2843) );
  INV_X1 U5171 ( .A(n4866), .ZN(n6335) );
  OR2_X1 U5172 ( .A1(n6530), .A2(n6531), .ZN(n4746) );
  AOI21_X1 U5173 ( .B1(n6516), .B2(n6515), .A(n6514), .ZN(n6806) );
  NOR2_X1 U5175 ( .A1(n7952), .A2(n7423), .ZN(n4483) );
  AND2_X1 U5176 ( .A1(n1698), .A2(n4621), .ZN(n2160) );
  INV_X1 U5177 ( .A(n4621), .ZN(n6425) );
  AND2_X1 U5179 ( .A1(n6712), .A2(n24501), .ZN(n3445) );
  OR2_X1 U5180 ( .A1(n7255), .A2(n7600), .ZN(n1902) );
  AND2_X1 U5181 ( .A1(n6682), .A2(n6685), .ZN(n4826) );
  NAND2_X1 U5182 ( .A1(n2279), .A2(n2278), .ZN(n7864) );
  NAND3_X1 U5183 ( .A1(n6293), .A2(n6481), .A3(n6198), .ZN(n2278) );
  OR2_X1 U5184 ( .A1(n6489), .A2(n6493), .ZN(n6781) );
  INV_X1 U5185 ( .A(n7732), .ZN(n7640) );
  OR2_X1 U5186 ( .A1(n4621), .A2(n6470), .ZN(n6203) );
  OAI21_X1 U5187 ( .B1(n25404), .B2(n1698), .A(n5966), .ZN(n1696) );
  AOI21_X1 U5188 ( .B1(n2351), .B2(n2350), .A(n5964), .ZN(n7461) );
  INV_X1 U5189 ( .A(n2352), .ZN(n2351) );
  OR2_X1 U5190 ( .A1(n6692), .A2(n6977), .ZN(n4828) );
  AND2_X1 U5191 ( .A1(n7532), .A2(n5738), .ZN(n2196) );
  INV_X1 U5192 ( .A(n2534), .ZN(n7100) );
  OAI211_X1 U5193 ( .C1(n7103), .C2(n6539), .A(n2532), .B(n6543), .ZN(n7104)
         );
  OR2_X1 U5195 ( .A1(n7975), .A2(n7976), .ZN(n7517) );
  INV_X1 U5197 ( .A(n7234), .ZN(n7682) );
  AND2_X1 U5198 ( .A1(n6733), .A2(n6395), .ZN(n2900) );
  INV_X1 U5200 ( .A(n7525), .ZN(n1677) );
  OR2_X1 U5201 ( .A1(n7768), .A2(n7526), .ZN(n4247) );
  AND2_X1 U5202 ( .A1(n5574), .A2(n3444), .ZN(n1641) );
  INV_X1 U5203 ( .A(n1558), .ZN(n1559) );
  OR2_X1 U5204 ( .A1(n25253), .A2(n7449), .ZN(n7636) );
  AND2_X1 U5206 ( .A1(n6301), .A2(n6784), .ZN(n1561) );
  INV_X1 U5207 ( .A(n9066), .ZN(n7427) );
  NOR2_X1 U5208 ( .A1(n7217), .A2(n8316), .ZN(n7698) );
  INV_X1 U5209 ( .A(n7595), .ZN(n7135) );
  OR2_X1 U5210 ( .A1(n6805), .A2(n8527), .ZN(n6549) );
  INV_X1 U5212 ( .A(n7860), .ZN(n4537) );
  OR2_X1 U5214 ( .A1(n6403), .A2(n6752), .ZN(n1735) );
  OR2_X1 U5215 ( .A1(n6630), .A2(n6407), .ZN(n6412) );
  INV_X1 U5216 ( .A(n7474), .ZN(n5413) );
  INV_X1 U5217 ( .A(n7615), .ZN(n7385) );
  OR2_X1 U5218 ( .A1(n7896), .A2(n3469), .ZN(n2846) );
  INV_X1 U5220 ( .A(n8457), .ZN(n8764) );
  INV_X1 U5221 ( .A(n4400), .ZN(n7971) );
  INV_X1 U5222 ( .A(n7349), .ZN(n8508) );
  AND2_X1 U5223 ( .A1(n4259), .A2(n7657), .ZN(n7228) );
  AND2_X1 U5224 ( .A1(n5651), .A2(n6772), .ZN(n2836) );
  AND2_X1 U5225 ( .A1(n6312), .A2(n6311), .ZN(n3608) );
  AND2_X1 U5226 ( .A1(n7862), .A2(n7864), .ZN(n7553) );
  INV_X1 U5227 ( .A(n8005), .ZN(n7543) );
  AOI21_X1 U5228 ( .B1(n6171), .B2(n6170), .A(n6350), .ZN(n5068) );
  AND2_X1 U5229 ( .A1(n6191), .A2(n7761), .ZN(n7391) );
  INV_X1 U5230 ( .A(n5202), .ZN(n3268) );
  NOR2_X1 U5231 ( .A1(n8005), .A2(n7292), .ZN(n2520) );
  OR2_X1 U5232 ( .A1(n9066), .A2(n9067), .ZN(n7428) );
  NOR2_X1 U5233 ( .A1(n7588), .A2(n7335), .ZN(n7338) );
  INV_X1 U5234 ( .A(n7943), .ZN(n6931) );
  OR2_X1 U5235 ( .A1(n7489), .A2(n7943), .ZN(n6929) );
  INV_X1 U5236 ( .A(n8316), .ZN(n8314) );
  INV_X1 U5237 ( .A(n7255), .ZN(n7598) );
  INV_X1 U5238 ( .A(n7537), .ZN(n8013) );
  OR2_X1 U5239 ( .A1(n6582), .A2(n6755), .ZN(n5604) );
  INV_X1 U5240 ( .A(n5607), .ZN(n5460) );
  OR2_X1 U5241 ( .A1(n6243), .A2(n6114), .ZN(n6720) );
  OR2_X1 U5242 ( .A1(n6824), .A2(n6829), .ZN(n4122) );
  AND2_X1 U5243 ( .A1(n7475), .A2(n7474), .ZN(n7221) );
  INV_X1 U5244 ( .A(n1345), .ZN(n3488) );
  OR2_X1 U5245 ( .A1(n7961), .A2(n7683), .ZN(n7485) );
  OR2_X1 U5246 ( .A1(n7942), .A2(n4672), .ZN(n3677) );
  AND2_X1 U5247 ( .A1(n7861), .A2(n7707), .ZN(n7271) );
  INV_X1 U5248 ( .A(n7861), .ZN(n7868) );
  NAND2_X1 U5250 ( .A1(n1839), .A2(n7462), .ZN(n5552) );
  AND2_X1 U5251 ( .A1(n268), .A2(n5970), .ZN(n5549) );
  OR2_X1 U5252 ( .A1(n7908), .A2(n7364), .ZN(n5390) );
  AND2_X1 U5254 ( .A1(n25252), .A2(n7768), .ZN(n7525) );
  INV_X1 U5255 ( .A(n7322), .ZN(n7891) );
  OR2_X1 U5256 ( .A1(n4839), .A2(n442), .ZN(n3142) );
  INV_X1 U5257 ( .A(n7578), .ZN(n7576) );
  AND2_X1 U5259 ( .A1(n7141), .A2(n7902), .ZN(n2780) );
  NAND3_X1 U5260 ( .A1(n5265), .A2(n5268), .A3(n5263), .ZN(n8477) );
  AND2_X1 U5261 ( .A1(n7734), .A2(n7642), .ZN(n7730) );
  OR2_X1 U5262 ( .A1(n6950), .A2(n25437), .ZN(n4757) );
  AOI21_X1 U5263 ( .B1(n3923), .B2(n6553), .A(n3922), .ZN(n3921) );
  OR2_X1 U5264 ( .A1(n6137), .A2(n6705), .ZN(n3924) );
  OR2_X1 U5265 ( .A1(n440), .A2(n6524), .ZN(n6154) );
  OR2_X1 U5266 ( .A1(n6963), .A2(n6570), .ZN(n6571) );
  OR2_X1 U5267 ( .A1(n6688), .A2(n6686), .ZN(n6567) );
  OR2_X1 U5268 ( .A1(n1985), .A2(n7965), .ZN(n7236) );
  OR2_X1 U5269 ( .A1(n7070), .A2(n7962), .ZN(n1984) );
  AND2_X1 U5270 ( .A1(n5713), .A2(n7433), .ZN(n2858) );
  OR2_X1 U5271 ( .A1(n7175), .A2(n7782), .ZN(n7176) );
  AOI21_X1 U5272 ( .B1(n4705), .B2(n3344), .A(n3587), .ZN(n4710) );
  OR2_X1 U5274 ( .A1(n3979), .A2(n8367), .ZN(n7558) );
  INV_X1 U5275 ( .A(n8616), .ZN(n8400) );
  AND2_X1 U5276 ( .A1(n7740), .A2(n7811), .ZN(n4803) );
  OR2_X1 U5277 ( .A1(n9469), .A2(n1595), .ZN(n1594) );
  INV_X1 U5278 ( .A(n9959), .ZN(n2876) );
  AND2_X2 U5279 ( .A1(n2275), .A2(n4785), .ZN(n8721) );
  OR2_X1 U5280 ( .A1(n4784), .A2(n7661), .ZN(n2275) );
  XNOR2_X1 U5281 ( .A(n8806), .B(n8492), .ZN(n8714) );
  OR2_X1 U5282 ( .A1(n7345), .A2(n7600), .ZN(n1999) );
  INV_X1 U5283 ( .A(n8501), .ZN(n8973) );
  INV_X1 U5284 ( .A(n2058), .ZN(n5328) );
  INV_X1 U5285 ( .A(n8798), .ZN(n5343) );
  XNOR2_X1 U5286 ( .A(n2560), .B(n8923), .ZN(n7083) );
  XNOR2_X1 U5287 ( .A(n8416), .B(n8415), .ZN(n10157) );
  AND2_X1 U5288 ( .A1(n9843), .A2(n10149), .ZN(n9844) );
  INV_X1 U5289 ( .A(n9211), .ZN(n7437) );
  INV_X1 U5291 ( .A(n25232), .ZN(n5621) );
  AND2_X1 U5292 ( .A1(n10951), .A2(n25074), .ZN(n5106) );
  INV_X1 U5293 ( .A(n10703), .ZN(n5107) );
  AND2_X1 U5294 ( .A1(n9435), .A2(n9635), .ZN(n1939) );
  XNOR2_X1 U5295 ( .A(n8130), .B(n8129), .ZN(n9944) );
  AND2_X1 U5296 ( .A1(n24083), .A2(n9899), .ZN(n9289) );
  OR2_X1 U5297 ( .A1(n10168), .A2(n10166), .ZN(n2091) );
  INV_X1 U5298 ( .A(n10811), .ZN(n5628) );
  INV_X1 U5299 ( .A(n10314), .ZN(n10165) );
  AND2_X1 U5300 ( .A1(n11215), .A2(n10669), .ZN(n5085) );
  AND2_X1 U5301 ( .A1(n10942), .A2(n11039), .ZN(n2870) );
  AND2_X1 U5302 ( .A1(n9872), .A2(n2294), .ZN(n2293) );
  AOI21_X1 U5303 ( .B1(n9883), .B2(n25069), .A(n9563), .ZN(n5066) );
  INV_X1 U5305 ( .A(n11046), .ZN(n10641) );
  INV_X1 U5306 ( .A(n10757), .ZN(n2867) );
  NAND2_X1 U5307 ( .A1(n9342), .A2(n1464), .ZN(n1658) );
  OR2_X1 U5308 ( .A1(n9668), .A2(n9999), .ZN(n9311) );
  OR2_X1 U5309 ( .A1(n10054), .A2(n10052), .ZN(n1871) );
  AND2_X1 U5311 ( .A1(n10989), .A2(n10406), .ZN(n10996) );
  OR2_X1 U5312 ( .A1(n25229), .A2(n10737), .ZN(n10283) );
  INV_X1 U5313 ( .A(n10858), .ZN(n10859) );
  NOR2_X1 U5314 ( .A1(n8178), .A2(n8179), .ZN(n10994) );
  AND2_X1 U5315 ( .A1(n10406), .A2(n10990), .ZN(n8146) );
  OR2_X1 U5316 ( .A1(n3467), .A2(n11101), .ZN(n2849) );
  INV_X1 U5317 ( .A(n10891), .ZN(n2185) );
  OR3_X1 U5318 ( .A1(n10830), .A2(n10831), .A3(n10836), .ZN(n4778) );
  OR2_X1 U5319 ( .A1(n25217), .A2(n9603), .ZN(n2928) );
  INV_X1 U5320 ( .A(n12261), .ZN(n12218) );
  NOR2_X1 U5321 ( .A1(n4251), .A2(n11059), .ZN(n4392) );
  AND2_X1 U5322 ( .A1(n11052), .A2(n11058), .ZN(n4391) );
  INV_X1 U5323 ( .A(n10627), .ZN(n11563) );
  OR2_X1 U5324 ( .A1(n10924), .A2(n10993), .ZN(n4929) );
  OR2_X1 U5325 ( .A1(n10185), .A2(n9520), .ZN(n5534) );
  INV_X1 U5326 ( .A(n10558), .ZN(n10556) );
  INV_X1 U5327 ( .A(n4521), .ZN(n9810) );
  NAND4_X1 U5328 ( .A1(n2152), .A2(n11056), .A3(n3163), .A4(n1389), .ZN(n4759)
         );
  INV_X1 U5329 ( .A(n10504), .ZN(n4671) );
  INV_X1 U5330 ( .A(n10951), .ZN(n10955) );
  INV_X1 U5331 ( .A(n11152), .ZN(n11147) );
  AND3_X1 U5332 ( .A1(n10447), .A2(n10448), .A3(n10446), .ZN(n11412) );
  AOI21_X1 U5333 ( .B1(n11300), .B2(n419), .A(n11299), .ZN(n11306) );
  INV_X1 U5334 ( .A(n11146), .ZN(n2060) );
  NOR2_X1 U5335 ( .A1(n25249), .A2(n10714), .ZN(n11131) );
  INV_X1 U5337 ( .A(n10398), .ZN(n10661) );
  INV_X1 U5338 ( .A(n2243), .ZN(n10830) );
  INV_X1 U5339 ( .A(n10941), .ZN(n10944) );
  OAI21_X1 U5340 ( .B1(n9919), .B2(n9355), .A(n3967), .ZN(n9136) );
  AND2_X1 U5341 ( .A1(n9135), .A2(n9912), .ZN(n2810) );
  AND2_X1 U5342 ( .A1(n9461), .A2(n9463), .ZN(n3967) );
  INV_X1 U5343 ( .A(n11113), .ZN(n11110) );
  INV_X1 U5345 ( .A(n12221), .ZN(n5180) );
  INV_X1 U5346 ( .A(n11044), .ZN(n4532) );
  INV_X1 U5347 ( .A(n11012), .ZN(n2681) );
  NOR2_X1 U5348 ( .A1(n11024), .A2(n8934), .ZN(n3771) );
  AND2_X1 U5349 ( .A1(n10858), .A2(n25230), .ZN(n5727) );
  INV_X1 U5350 ( .A(n12134), .ZN(n12109) );
  INV_X1 U5351 ( .A(n11628), .ZN(n12356) );
  INV_X1 U5352 ( .A(n5340), .ZN(n10261) );
  OAI21_X1 U5353 ( .B1(n10148), .B2(n5357), .A(n5355), .ZN(n10867) );
  INV_X1 U5354 ( .A(n1658), .ZN(n10875) );
  INV_X1 U5356 ( .A(n5448), .ZN(n2498) );
  OR2_X1 U5357 ( .A1(n11070), .A2(n25203), .ZN(n3573) );
  INV_X1 U5358 ( .A(n11412), .ZN(n12168) );
  INV_X1 U5359 ( .A(n1499), .ZN(n10759) );
  NOR2_X1 U5360 ( .A1(n10753), .A2(n1499), .ZN(n3750) );
  INV_X1 U5361 ( .A(n3324), .ZN(n10291) );
  XNOR2_X1 U5362 ( .A(n12261), .B(n3158), .ZN(n12220) );
  OR2_X1 U5363 ( .A1(n4937), .A2(n10734), .ZN(n2830) );
  XNOR2_X1 U5364 ( .A(n3418), .B(n12180), .ZN(n12182) );
  XNOR2_X1 U5365 ( .A(n12306), .B(n3133), .ZN(n3418) );
  XNOR2_X1 U5366 ( .A(n11913), .B(n11914), .ZN(n2271) );
  XNOR2_X1 U5367 ( .A(n12128), .B(n12355), .ZN(n3207) );
  INV_X1 U5368 ( .A(n2739), .ZN(n4107) );
  XNOR2_X1 U5369 ( .A(n11268), .B(n3901), .ZN(n12266) );
  INV_X1 U5370 ( .A(n12315), .ZN(n5181) );
  OR2_X1 U5371 ( .A1(n10940), .A2(n24591), .ZN(n3252) );
  XNOR2_X1 U5372 ( .A(n25396), .B(n5514), .ZN(n11571) );
  INV_X1 U5373 ( .A(n11542), .ZN(n1699) );
  INV_X1 U5374 ( .A(n4759), .ZN(n11706) );
  NAND2_X1 U5376 ( .A1(n11081), .A2(n4421), .ZN(n10222) );
  OR2_X1 U5377 ( .A1(n10767), .A2(n4422), .ZN(n4421) );
  INV_X1 U5378 ( .A(n13153), .ZN(n1632) );
  INV_X1 U5379 ( .A(n11424), .ZN(n10490) );
  AND2_X1 U5380 ( .A1(n2628), .A2(n11342), .ZN(n10493) );
  OR2_X1 U5381 ( .A1(n10425), .A2(n10596), .ZN(n4211) );
  INV_X1 U5382 ( .A(n1543), .ZN(n1538) );
  INV_X1 U5383 ( .A(n1544), .ZN(n1537) );
  INV_X1 U5385 ( .A(n11199), .ZN(n10229) );
  XNOR2_X1 U5386 ( .A(n11401), .B(n2602), .ZN(n11665) );
  AND2_X1 U5388 ( .A1(n24930), .A2(n3688), .ZN(n11596) );
  NOR2_X1 U5389 ( .A1(n414), .A2(n4711), .ZN(n11934) );
  INV_X1 U5391 ( .A(n12219), .ZN(n5182) );
  AOI22_X1 U5392 ( .A1(n9241), .A2(n11124), .B1(n10846), .B2(n305), .ZN(n9242)
         );
  AND2_X1 U5393 ( .A1(n2680), .A2(n11012), .ZN(n10013) );
  OR2_X1 U5394 ( .A1(n13347), .A2(n12636), .ZN(n12858) );
  AND2_X1 U5395 ( .A1(n13169), .A2(n13167), .ZN(n12721) );
  INV_X1 U5397 ( .A(n302), .ZN(n1636) );
  INV_X1 U5402 ( .A(n24512), .ZN(n13215) );
  OR2_X1 U5403 ( .A1(n13040), .A2(n12800), .ZN(n4639) );
  OR2_X1 U5405 ( .A1(n12685), .A2(n5311), .ZN(n5314) );
  OR2_X1 U5406 ( .A1(n12684), .A2(n24422), .ZN(n5309) );
  NOR2_X1 U5407 ( .A1(n3689), .A2(n24373), .ZN(n13172) );
  INV_X1 U5408 ( .A(n12669), .ZN(n3563) );
  AND2_X1 U5409 ( .A1(n14333), .A2(n14339), .ZN(n13878) );
  OR2_X1 U5410 ( .A1(n13146), .A2(n13145), .ZN(n5543) );
  OR2_X1 U5411 ( .A1(n5412), .A2(n12858), .ZN(n3339) );
  INV_X1 U5412 ( .A(n13109), .ZN(n4529) );
  INV_X1 U5413 ( .A(n13485), .ZN(n14005) );
  INV_X1 U5414 ( .A(n14362), .ZN(n3698) );
  AND2_X1 U5415 ( .A1(n13569), .A2(n13394), .ZN(n3808) );
  NOR2_X1 U5416 ( .A1(n11601), .A2(n11600), .ZN(n3807) );
  AND2_X1 U5417 ( .A1(n13323), .A2(n2295), .ZN(n12848) );
  INV_X1 U5419 ( .A(n14107), .ZN(n13566) );
  INV_X1 U5420 ( .A(n13265), .ZN(n5644) );
  INV_X1 U5421 ( .A(n14129), .ZN(n13893) );
  AND2_X1 U5422 ( .A1(n13868), .A2(n14317), .ZN(n3501) );
  INV_X1 U5423 ( .A(n13647), .ZN(n13819) );
  INV_X1 U5424 ( .A(n14328), .ZN(n2505) );
  AND2_X1 U5425 ( .A1(n12633), .A2(n4923), .ZN(n5471) );
  OR2_X1 U5426 ( .A1(n13953), .A2(n14158), .ZN(n4356) );
  INV_X1 U5427 ( .A(n14211), .ZN(n13437) );
  AOI22_X1 U5429 ( .A1(n12876), .A2(n13357), .B1(n13359), .B2(n24554), .ZN(
        n2889) );
  AND2_X1 U5431 ( .A1(n14035), .A2(n14034), .ZN(n13806) );
  OAI21_X1 U5433 ( .B1(n12507), .B2(n12506), .A(n3633), .ZN(n3632) );
  OR2_X1 U5434 ( .A1(n14022), .A2(n13533), .ZN(n13609) );
  AND2_X1 U5435 ( .A1(n12018), .A2(n1527), .ZN(n1526) );
  NOR2_X1 U5437 ( .A1(n14172), .A2(n14165), .ZN(n3383) );
  NOR2_X1 U5439 ( .A1(n14000), .A2(n12668), .ZN(n13676) );
  INV_X1 U5440 ( .A(n14165), .ZN(n13741) );
  INV_X1 U5442 ( .A(n14190), .ZN(n14142) );
  INV_X1 U5443 ( .A(n12536), .ZN(n13759) );
  AND2_X1 U5444 ( .A1(n14274), .A2(n14268), .ZN(n13764) );
  AOI21_X1 U5445 ( .B1(n13733), .B2(n13732), .A(n13731), .ZN(n14594) );
  AND2_X1 U5446 ( .A1(n14106), .A2(n14108), .ZN(n1933) );
  AND3_X1 U5447 ( .A1(n13792), .A2(n13796), .A3(n13578), .ZN(n4331) );
  OR2_X1 U5448 ( .A1(n14302), .A2(n14301), .ZN(n13454) );
  AND2_X1 U5449 ( .A1(n14153), .A2(n3717), .ZN(n3716) );
  INV_X1 U5450 ( .A(n14089), .ZN(n14018) );
  OR2_X1 U5451 ( .A1(n13824), .A2(n13560), .ZN(n13389) );
  INV_X1 U5453 ( .A(n13048), .ZN(n12489) );
  INV_X1 U5454 ( .A(n4059), .ZN(n4058) );
  OR2_X1 U5456 ( .A1(n12843), .A2(n12946), .ZN(n2770) );
  OR2_X1 U5457 ( .A1(n12844), .A2(n12845), .ZN(n2769) );
  AND2_X1 U5458 ( .A1(n14294), .A2(n14290), .ZN(n13722) );
  NOR2_X1 U5459 ( .A1(n13895), .A2(n4844), .ZN(n4043) );
  AND2_X1 U5460 ( .A1(n399), .A2(n13338), .ZN(n12959) );
  INV_X1 U5461 ( .A(n14124), .ZN(n14123) );
  INV_X1 U5462 ( .A(n13422), .ZN(n2378) );
  INV_X1 U5463 ( .A(n14205), .ZN(n2379) );
  OR2_X1 U5465 ( .A1(n14219), .A2(n14222), .ZN(n13022) );
  OR2_X1 U5466 ( .A1(n13863), .A2(n13864), .ZN(n12814) );
  OAI211_X1 U5468 ( .C1(n5485), .C2(n5487), .A(n5483), .B(n5482), .ZN(n14966)
         );
  OAI21_X1 U5469 ( .B1(n15216), .B2(n15215), .A(n16641), .ZN(n16945) );
  OR2_X1 U5473 ( .A1(n16422), .A2(n16427), .ZN(n16171) );
  OAI21_X1 U5474 ( .B1(n13724), .B2(n11806), .A(n1771), .ZN(n13727) );
  AND2_X1 U5475 ( .A1(n14078), .A2(n14077), .ZN(n2122) );
  AND2_X1 U5476 ( .A1(n16443), .A2(n16442), .ZN(n2809) );
  OR2_X1 U5477 ( .A1(n16038), .A2(n16043), .ZN(n3578) );
  XNOR2_X1 U5478 ( .A(n14830), .B(n1371), .ZN(n15564) );
  INV_X1 U5479 ( .A(n14500), .ZN(n14806) );
  OR2_X1 U5480 ( .A1(n386), .A2(n25210), .ZN(n4026) );
  XNOR2_X1 U5481 ( .A(n15435), .B(n15434), .ZN(n15470) );
  OR2_X1 U5482 ( .A1(n15714), .A2(n16470), .ZN(n4972) );
  INV_X1 U5483 ( .A(n24539), .ZN(n4927) );
  OR2_X1 U5484 ( .A1(n15977), .A2(n16394), .ZN(n1656) );
  INV_X1 U5485 ( .A(n16225), .ZN(n16301) );
  OR2_X1 U5486 ( .A1(n15686), .A2(n16437), .ZN(n2637) );
  OR2_X1 U5487 ( .A1(n16076), .A2(n14664), .ZN(n3636) );
  INV_X1 U5488 ( .A(n16207), .ZN(n4914) );
  AND2_X1 U5490 ( .A1(n17421), .A2(n16945), .ZN(n2234) );
  NOR2_X1 U5491 ( .A1(n2375), .A2(n4897), .ZN(n15691) );
  NOR2_X1 U5492 ( .A1(n16048), .A2(n15605), .ZN(n15604) );
  XNOR2_X1 U5493 ( .A(n3471), .B(n14962), .ZN(n2407) );
  INV_X1 U5494 ( .A(n15953), .ZN(n15717) );
  XNOR2_X1 U5495 ( .A(n5009), .B(n15352), .ZN(n15353) );
  OR2_X1 U5496 ( .A1(n17085), .A2(n17088), .ZN(n3103) );
  INV_X1 U5497 ( .A(n4985), .ZN(n4981) );
  INV_X1 U5498 ( .A(n15314), .ZN(n17343) );
  XNOR2_X1 U5501 ( .A(n2969), .B(n1907), .ZN(n14693) );
  AND2_X1 U5502 ( .A1(n16595), .A2(n24587), .ZN(n15824) );
  AND2_X1 U5503 ( .A1(n5447), .A2(n5667), .ZN(n5668) );
  OAI211_X1 U5504 ( .C1(n5447), .C2(n16001), .A(n15758), .B(n3658), .ZN(n5666)
         );
  OAI21_X1 U5505 ( .B1(n16185), .B2(n15915), .A(n5317), .ZN(n1516) );
  OR2_X1 U5506 ( .A1(n16355), .A2(n16360), .ZN(n4496) );
  OR2_X1 U5507 ( .A1(n16770), .A2(n17039), .ZN(n17363) );
  INV_X1 U5509 ( .A(n15937), .ZN(n5168) );
  NOR2_X1 U5510 ( .A1(n15695), .A2(n15953), .ZN(n16482) );
  XNOR2_X1 U5511 ( .A(n14262), .B(n14263), .ZN(n15837) );
  AND2_X1 U5512 ( .A1(n4046), .A2(n15837), .ZN(n15839) );
  AND2_X1 U5514 ( .A1(n16551), .A2(n5376), .ZN(n15739) );
  OR2_X1 U5516 ( .A1(n14787), .A2(n24163), .ZN(n3067) );
  XNOR2_X1 U5517 ( .A(n14822), .B(n14821), .ZN(n16230) );
  INV_X1 U5518 ( .A(n17320), .ZN(n2287) );
  AND2_X1 U5519 ( .A1(n16769), .A2(n17364), .ZN(n2530) );
  OAI21_X1 U5520 ( .B1(n24586), .B2(n4807), .A(n4806), .ZN(n16687) );
  OR2_X1 U5521 ( .A1(n4353), .A2(n15594), .ZN(n4938) );
  OR2_X1 U5522 ( .A1(n3702), .A2(n16438), .ZN(n2202) );
  AND2_X1 U5523 ( .A1(n16241), .A2(n16437), .ZN(n3702) );
  INV_X1 U5524 ( .A(n17212), .ZN(n5512) );
  INV_X1 U5525 ( .A(n15470), .ZN(n16472) );
  INV_X1 U5528 ( .A(n17728), .ZN(n1704) );
  OR2_X1 U5529 ( .A1(n17690), .A2(n17485), .ZN(n1701) );
  AND2_X1 U5531 ( .A1(n14585), .A2(n1676), .ZN(n1675) );
  INV_X1 U5532 ( .A(n17433), .ZN(n3000) );
  AND2_X1 U5533 ( .A1(n17312), .A2(n17316), .ZN(n16716) );
  OR2_X1 U5534 ( .A1(n17596), .A2(n24543), .ZN(n4564) );
  OR2_X1 U5535 ( .A1(n17364), .A2(n25058), .ZN(n3951) );
  OR2_X1 U5536 ( .A1(n16064), .A2(n16067), .ZN(n4105) );
  NOR2_X1 U5537 ( .A1(n25245), .A2(n17132), .ZN(n3457) );
  OR2_X1 U5538 ( .A1(n15668), .A2(n290), .ZN(n2286) );
  OR2_X1 U5539 ( .A1(n17319), .A2(n16607), .ZN(n16923) );
  OAI21_X1 U5540 ( .B1(n13547), .B2(n267), .A(n13546), .ZN(n17225) );
  INV_X1 U5541 ( .A(n17225), .ZN(n16956) );
  INV_X1 U5542 ( .A(n17387), .ZN(n3604) );
  NAND3_X1 U5543 ( .A1(n382), .A2(n25446), .A3(n15550), .ZN(n5596) );
  AOI22_X1 U5544 ( .A1(n16828), .A2(n16962), .B1(n1612), .B2(n24444), .ZN(
        n17128) );
  OR2_X1 U5545 ( .A1(n15266), .A2(n24429), .ZN(n3121) );
  OAI21_X1 U5547 ( .B1(n15940), .B2(n24163), .A(n24162), .ZN(n2344) );
  INV_X1 U5548 ( .A(n16927), .ZN(n17322) );
  INV_X1 U5549 ( .A(n16971), .ZN(n17332) );
  OR2_X1 U5550 ( .A1(n25409), .A2(n15584), .ZN(n3503) );
  AND2_X1 U5551 ( .A1(n17316), .A2(n24543), .ZN(n3627) );
  AND2_X1 U5552 ( .A1(n17320), .A2(n16927), .ZN(n17267) );
  AND2_X1 U5553 ( .A1(n17371), .A2(n17042), .ZN(n16766) );
  OR2_X1 U5554 ( .A1(n17414), .A2(n17225), .ZN(n5705) );
  INV_X1 U5555 ( .A(n16486), .ZN(n16518) );
  AND2_X1 U5556 ( .A1(n16851), .A2(n17138), .ZN(n3930) );
  AND2_X1 U5557 ( .A1(n17145), .A2(n16984), .ZN(n3929) );
  INV_X1 U5558 ( .A(n3778), .ZN(n14864) );
  OR2_X1 U5559 ( .A1(n17608), .A2(n17409), .ZN(n16743) );
  OR2_X1 U5560 ( .A1(n16311), .A2(n16312), .ZN(n1817) );
  OR2_X1 U5561 ( .A1(n16298), .A2(n4957), .ZN(n4956) );
  INV_X1 U5562 ( .A(n17131), .ZN(n16655) );
  AND3_X1 U5563 ( .A1(n17081), .A2(n17078), .A3(n17478), .ZN(n2181) );
  NOR2_X1 U5566 ( .A1(n16353), .A2(n16595), .ZN(n3334) );
  INV_X1 U5567 ( .A(n17114), .ZN(n4304) );
  INV_X1 U5568 ( .A(n17520), .ZN(n18311) );
  INV_X1 U5569 ( .A(n16921), .ZN(n17596) );
  AND2_X1 U5570 ( .A1(n17068), .A2(n16731), .ZN(n4286) );
  INV_X1 U5571 ( .A(n16769), .ZN(n3685) );
  NOR2_X1 U5572 ( .A1(n1451), .A2(n1498), .ZN(n1497) );
  AND2_X1 U5573 ( .A1(n15970), .A2(n16186), .ZN(n3223) );
  INV_X1 U5574 ( .A(n17624), .ZN(n4284) );
  INV_X1 U5575 ( .A(n17622), .ZN(n4285) );
  AND2_X1 U5576 ( .A1(n16112), .A2(n17524), .ZN(n17527) );
  AOI21_X1 U5578 ( .B1(n17314), .B2(n16921), .A(n2968), .ZN(n3782) );
  OR2_X1 U5580 ( .A1(n16440), .A2(n16442), .ZN(n15947) );
  XNOR2_X1 U5581 ( .A(n18375), .B(n16866), .ZN(n16867) );
  INV_X1 U5582 ( .A(n16846), .ZN(n16499) );
  OR2_X1 U5583 ( .A1(n16034), .A2(n15573), .ZN(n1927) );
  INV_X1 U5584 ( .A(n17410), .ZN(n17609) );
  INV_X1 U5585 ( .A(n16561), .ZN(n17407) );
  OR2_X1 U5586 ( .A1(n16961), .A2(n17445), .ZN(n3260) );
  NAND2_X1 U5587 ( .A1(n15845), .A2(n2992), .ZN(n17122) );
  XNOR2_X1 U5589 ( .A(n18157), .B(n24886), .ZN(n18159) );
  INV_X1 U5590 ( .A(n4114), .ZN(n2216) );
  OR2_X1 U5591 ( .A1(n19312), .A2(n19310), .ZN(n18843) );
  XNOR2_X1 U5592 ( .A(n4269), .B(n18429), .ZN(n4268) );
  INV_X1 U5593 ( .A(n18694), .ZN(n4269) );
  INV_X1 U5594 ( .A(n19413), .ZN(n3491) );
  BUF_X1 U5595 ( .A(n16910), .Z(n17907) );
  XNOR2_X1 U5596 ( .A(n2001), .B(n18128), .ZN(n18464) );
  INV_X1 U5597 ( .A(n18129), .ZN(n2001) );
  INV_X1 U5598 ( .A(n18172), .ZN(n4971) );
  INV_X1 U5599 ( .A(n19255), .ZN(n18870) );
  XNOR2_X1 U5600 ( .A(n18520), .B(n18519), .ZN(n19064) );
  AND2_X1 U5601 ( .A1(n19238), .A2(n18883), .ZN(n19067) );
  AND2_X1 U5602 ( .A1(n19331), .A2(n4291), .ZN(n5213) );
  INV_X1 U5603 ( .A(n20586), .ZN(n19951) );
  AND2_X1 U5604 ( .A1(n280), .A2(n19575), .ZN(n5155) );
  INV_X1 U5606 ( .A(n19064), .ZN(n2298) );
  AND2_X1 U5607 ( .A1(n19065), .A2(n25012), .ZN(n2328) );
  AND2_X1 U5608 ( .A1(n25012), .A2(n19064), .ZN(n19616) );
  AND2_X1 U5611 ( .A1(n17945), .A2(n4291), .ZN(n4288) );
  OR2_X1 U5612 ( .A1(n19202), .A2(n3412), .ZN(n19839) );
  NAND2_X1 U5613 ( .A1(n276), .A2(n24463), .ZN(n5132) );
  OR2_X1 U5615 ( .A1(n17872), .A2(n18959), .ZN(n3583) );
  AOI21_X1 U5616 ( .B1(n20554), .B2(n20555), .A(n2594), .ZN(n20559) );
  INV_X1 U5617 ( .A(n1590), .ZN(n2688) );
  OAI211_X1 U5618 ( .C1(n19080), .C2(n5134), .A(n19251), .B(n1501), .ZN(n5427)
         );
  AOI22_X1 U5619 ( .A1(n19079), .A2(n19592), .B1(n2346), .B2(n1502), .ZN(n1501) );
  AND2_X1 U5620 ( .A1(n18808), .A2(n19078), .ZN(n1502) );
  OR2_X1 U5621 ( .A1(n19532), .A2(n19272), .ZN(n5652) );
  NAND2_X1 U5622 ( .A1(n4857), .A2(n1505), .ZN(n1504) );
  OR2_X1 U5624 ( .A1(n19009), .A2(n19170), .ZN(n3820) );
  INV_X1 U5625 ( .A(n20149), .ZN(n20147) );
  OR2_X1 U5626 ( .A1(n19087), .A2(n24584), .ZN(n3668) );
  INV_X1 U5627 ( .A(n5427), .ZN(n20497) );
  AND2_X1 U5628 ( .A1(n20268), .A2(n20501), .ZN(n20225) );
  OAI21_X1 U5629 ( .B1(n18720), .B2(n18721), .A(n357), .ZN(n18722) );
  INV_X1 U5630 ( .A(n5475), .ZN(n5474) );
  INV_X1 U5631 ( .A(n5569), .ZN(n5568) );
  INV_X1 U5632 ( .A(n20576), .ZN(n19841) );
  OR2_X1 U5633 ( .A1(n24583), .A2(n4291), .ZN(n4287) );
  INV_X1 U5634 ( .A(n20345), .ZN(n1557) );
  OR2_X1 U5636 ( .A1(n100), .A2(n20507), .ZN(n5499) );
  INV_X1 U5637 ( .A(n20614), .ZN(n2330) );
  INV_X1 U5638 ( .A(n20617), .ZN(n20570) );
  INV_X1 U5639 ( .A(n20616), .ZN(n20569) );
  NOR2_X1 U5640 ( .A1(n5590), .A2(n20414), .ZN(n5733) );
  INV_X1 U5641 ( .A(n21533), .ZN(n4164) );
  OAI21_X1 U5643 ( .B1(n18828), .B2(n19002), .A(n4195), .ZN(n4194) );
  OR2_X1 U5644 ( .A1(n19777), .A2(n20173), .ZN(n20234) );
  OR2_X1 U5645 ( .A1(n19255), .A2(n25001), .ZN(n3388) );
  INV_X1 U5646 ( .A(n20269), .ZN(n20224) );
  INV_X1 U5647 ( .A(n20414), .ZN(n5591) );
  OR2_X1 U5648 ( .A1(n19112), .A2(n2642), .ZN(n18867) );
  OR2_X1 U5649 ( .A1(n19252), .A2(n19078), .ZN(n2804) );
  AND2_X1 U5650 ( .A1(n7), .A2(n20614), .ZN(n20572) );
  INV_X1 U5652 ( .A(n20145), .ZN(n20447) );
  OR2_X1 U5653 ( .A1(n20149), .A2(n19018), .ZN(n20532) );
  OR2_X1 U5654 ( .A1(n19168), .A2(n19002), .ZN(n2927) );
  OR2_X1 U5655 ( .A1(n25422), .A2(n19246), .ZN(n3987) );
  INV_X1 U5656 ( .A(n20335), .ZN(n20666) );
  OR2_X1 U5657 ( .A1(n20142), .A2(n19979), .ZN(n2074) );
  OR2_X1 U5658 ( .A1(n5007), .A2(n19441), .ZN(n2693) );
  OAI211_X1 U5659 ( .C1(n20114), .C2(n19887), .A(n19886), .B(n19885), .ZN(
        n20904) );
  INV_X1 U5660 ( .A(n18978), .ZN(n17892) );
  INV_X1 U5661 ( .A(n1591), .ZN(n19893) );
  INV_X1 U5662 ( .A(n20518), .ZN(n20276) );
  INV_X1 U5663 ( .A(n20437), .ZN(n20583) );
  INV_X1 U5664 ( .A(n20193), .ZN(n20577) );
  OR2_X1 U5665 ( .A1(n25205), .A2(n20231), .ZN(n19803) );
  AND2_X1 U5666 ( .A1(n2594), .A2(n20557), .ZN(n19880) );
  AOI21_X1 U5667 ( .B1(n352), .B2(n19345), .A(n19344), .ZN(n19348) );
  INV_X1 U5668 ( .A(n19383), .ZN(n4008) );
  OR2_X1 U5669 ( .A1(n19168), .A2(n19421), .ZN(n4578) );
  INV_X1 U5670 ( .A(n19423), .ZN(n4579) );
  OR2_X1 U5671 ( .A1(n18818), .A2(n19211), .ZN(n4851) );
  NOR2_X1 U5672 ( .A1(n24275), .A2(n20913), .ZN(n20362) );
  AND2_X1 U5673 ( .A1(n5132), .A2(n5131), .ZN(n5130) );
  INV_X1 U5674 ( .A(n20019), .ZN(n4728) );
  INV_X1 U5675 ( .A(n19703), .ZN(n20623) );
  INV_X1 U5676 ( .A(n19849), .ZN(n19852) );
  INV_X1 U5677 ( .A(n19661), .ZN(n19657) );
  NOR2_X1 U5678 ( .A1(n20555), .A2(n20554), .ZN(n2369) );
  INV_X1 U5679 ( .A(n20089), .ZN(n2370) );
  AND2_X1 U5680 ( .A1(n20330), .A2(n3480), .ZN(n20090) );
  AND2_X1 U5681 ( .A1(n4616), .A2(n4066), .ZN(n20009) );
  AND2_X1 U5682 ( .A1(n5686), .A2(n5685), .ZN(n17895) );
  OR2_X1 U5683 ( .A1(n20071), .A2(n3240), .ZN(n19661) );
  AND2_X1 U5684 ( .A1(n20518), .A2(n20516), .ZN(n19799) );
  INV_X1 U5685 ( .A(n19979), .ZN(n20296) );
  INV_X1 U5686 ( .A(n20142), .ZN(n20297) );
  NAND2_X1 U5687 ( .A1(n3239), .A2(n18846), .ZN(n19658) );
  OR2_X1 U5688 ( .A1(n19406), .A2(n19407), .ZN(n18782) );
  OR2_X1 U5689 ( .A1(n25489), .A2(n19397), .ZN(n4809) );
  NOR2_X1 U5690 ( .A1(n19510), .A2(n1419), .ZN(n3195) );
  INV_X1 U5691 ( .A(n20419), .ZN(n4509) );
  INV_X1 U5692 ( .A(n20174), .ZN(n20589) );
  NOR2_X1 U5693 ( .A1(n20576), .A2(n20578), .ZN(n20432) );
  NAND2_X1 U5694 ( .A1(n19843), .A2(n19839), .ZN(n20437) );
  OR2_X1 U5695 ( .A1(n5207), .A2(n20194), .ZN(n5206) );
  INV_X1 U5696 ( .A(n20411), .ZN(n20263) );
  NAND2_X1 U5698 ( .A1(n18974), .A2(n19478), .ZN(n4402) );
  INV_X1 U5699 ( .A(n19658), .ZN(n20069) );
  INV_X1 U5700 ( .A(n3428), .ZN(n2432) );
  OAI21_X1 U5701 ( .B1(n1601), .B2(n1600), .A(n24454), .ZN(n1599) );
  AND2_X1 U5702 ( .A1(n20370), .A2(n20374), .ZN(n1601) );
  OR2_X1 U5703 ( .A1(n19173), .A2(n19407), .ZN(n18826) );
  OAI22_X1 U5704 ( .A1(n20280), .A2(n20279), .B1(n20343), .B2(n20345), .ZN(
        n2699) );
  OAI21_X1 U5705 ( .B1(n20298), .B2(n19979), .A(n4615), .ZN(n20302) );
  OR2_X1 U5706 ( .A1(n19785), .A2(n24464), .ZN(n19750) );
  OR2_X1 U5708 ( .A1(n20022), .A2(n18395), .ZN(n19729) );
  OR2_X1 U5709 ( .A1(n18728), .A2(n2578), .ZN(n2854) );
  AND2_X1 U5710 ( .A1(n19490), .A2(n240), .ZN(n2578) );
  OR2_X1 U5711 ( .A1(n18717), .A2(n18990), .ZN(n2304) );
  AOI21_X1 U5712 ( .B1(n20562), .B2(n20094), .A(n25221), .ZN(n2469) );
  OR2_X1 U5713 ( .A1(n20560), .A2(n20094), .ZN(n2470) );
  INV_X1 U5714 ( .A(n20126), .ZN(n20312) );
  AND2_X1 U5715 ( .A1(n20345), .A2(n3671), .ZN(n4460) );
  OR2_X1 U5717 ( .A1(n20230), .A2(n343), .ZN(n5425) );
  INV_X1 U5718 ( .A(n19586), .ZN(n2068) );
  NOR2_X1 U5719 ( .A1(n4480), .A2(n19592), .ZN(n4479) );
  NOR2_X2 U5720 ( .A1(n19604), .A2(n19603), .ZN(n20960) );
  OR2_X1 U5723 ( .A1(n20411), .A2(n4184), .ZN(n4183) );
  OR2_X1 U5724 ( .A1(n20591), .A2(n20588), .ZN(n2724) );
  XNOR2_X1 U5726 ( .A(n21967), .B(n21735), .ZN(n4688) );
  AOI22_X1 U5727 ( .A1(n17849), .A2(n20117), .B1(n3326), .B2(n25388), .ZN(
        n3325) );
  NOR2_X1 U5729 ( .A1(n22355), .A2(n22356), .ZN(n4221) );
  INV_X1 U5730 ( .A(n19888), .ZN(n4174) );
  XNOR2_X1 U5731 ( .A(n21640), .B(n21596), .ZN(n20831) );
  INV_X1 U5733 ( .A(n22803), .ZN(n22585) );
  AND2_X1 U5735 ( .A1(n22452), .A2(n21918), .ZN(n5584) );
  NOR2_X1 U5736 ( .A1(n22779), .A2(n22782), .ZN(n22780) );
  INV_X1 U5737 ( .A(n23196), .ZN(n4113) );
  INV_X1 U5738 ( .A(n22333), .ZN(n21368) );
  OR2_X1 U5739 ( .A1(n22977), .A2(n22389), .ZN(n3210) );
  AOI21_X1 U5740 ( .B1(n1766), .B2(n1765), .A(n22941), .ZN(n22942) );
  NAND2_X1 U5741 ( .A1(n24932), .A2(n22829), .ZN(n4608) );
  INV_X1 U5742 ( .A(n4633), .ZN(n22436) );
  NOR2_X1 U5743 ( .A1(n22959), .A2(n24885), .ZN(n22858) );
  AND2_X1 U5744 ( .A1(n24397), .A2(n23592), .ZN(n21946) );
  INV_X1 U5745 ( .A(n22159), .ZN(n2312) );
  INV_X1 U5746 ( .A(n21829), .ZN(n1728) );
  NOR2_X1 U5747 ( .A1(n21825), .A2(n22252), .ZN(n22521) );
  NOR2_X1 U5751 ( .A1(n331), .A2(n25241), .ZN(n22609) );
  INV_X1 U5752 ( .A(n4273), .ZN(n4168) );
  NAND2_X1 U5753 ( .A1(n22363), .A2(n25241), .ZN(n2528) );
  OAI21_X1 U5754 ( .B1(n22806), .B2(n22807), .A(n24992), .ZN(n4427) );
  INV_X1 U5755 ( .A(n24325), .ZN(n4630) );
  AND2_X1 U5756 ( .A1(n24381), .A2(n23714), .ZN(n3282) );
  OR2_X1 U5760 ( .A1(n22450), .A2(n274), .ZN(n5260) );
  INV_X1 U5761 ( .A(n23104), .ZN(n23123) );
  OR2_X1 U5763 ( .A1(n21379), .A2(n274), .ZN(n5048) );
  OR2_X1 U5764 ( .A1(n23165), .A2(n23178), .ZN(n22553) );
  AOI22_X1 U5765 ( .A1(n22324), .A2(n22325), .B1(n22452), .B2(n22456), .ZN(
        n3682) );
  OR2_X1 U5766 ( .A1(n23190), .A2(n23200), .ZN(n3037) );
  INV_X1 U5768 ( .A(n22561), .ZN(n22573) );
  INV_X1 U5769 ( .A(n3720), .ZN(n2869) );
  OR2_X1 U5770 ( .A1(n3720), .A2(n23252), .ZN(n3719) );
  NAND2_X1 U5771 ( .A1(n23252), .A2(n23253), .ZN(n4243) );
  AND2_X1 U5773 ( .A1(n3623), .A2(n22508), .ZN(n2861) );
  AOI21_X1 U5775 ( .B1(n25081), .B2(n1500), .A(n24309), .ZN(n2921) );
  OR2_X1 U5776 ( .A1(n21886), .A2(n3781), .ZN(n1684) );
  OR2_X1 U5777 ( .A1(n1685), .A2(n3781), .ZN(n1682) );
  OR2_X1 U5778 ( .A1(n4372), .A2(n22972), .ZN(n22978) );
  OR2_X1 U5779 ( .A1(n22744), .A2(n4606), .ZN(n4605) );
  OR2_X1 U5781 ( .A1(n22430), .A2(n23368), .ZN(n3528) );
  INV_X1 U5782 ( .A(n22026), .ZN(n23392) );
  AND2_X1 U5783 ( .A1(n23449), .A2(n22528), .ZN(n4311) );
  INV_X1 U5784 ( .A(n23480), .ZN(n23492) );
  OR2_X1 U5785 ( .A1(n23480), .A2(n2710), .ZN(n23485) );
  INV_X1 U5787 ( .A(n4949), .ZN(n23516) );
  INV_X1 U5788 ( .A(n23531), .ZN(n5701) );
  AND2_X1 U5789 ( .A1(n23592), .A2(n23596), .ZN(n5437) );
  AND3_X1 U5791 ( .A1(n22727), .A2(n20893), .A3(n20892), .ZN(n20895) );
  NOR2_X1 U5792 ( .A1(n23645), .A2(n23634), .ZN(n23629) );
  NOR2_X1 U5793 ( .A1(n23665), .A2(n5507), .ZN(n23669) );
  INV_X1 U5794 ( .A(n23727), .ZN(n3283) );
  AND2_X1 U5796 ( .A1(n24362), .A2(n4374), .ZN(n23752) );
  AND2_X1 U5797 ( .A1(n23767), .A2(n25051), .ZN(n2982) );
  AND2_X1 U5798 ( .A1(n23769), .A2(n25051), .ZN(n2783) );
  OR2_X1 U5799 ( .A1(n23789), .A2(n24307), .ZN(n4954) );
  AND2_X1 U5800 ( .A1(n22043), .A2(n23805), .ZN(n3495) );
  OR2_X1 U5801 ( .A1(n24392), .A2(n3201), .ZN(n23789) );
  AND2_X1 U5802 ( .A1(n3456), .A2(n3070), .ZN(n21346) );
  OR2_X1 U5803 ( .A1(n22214), .A2(n21341), .ZN(n3070) );
  OR2_X1 U5804 ( .A1(n21352), .A2(n21362), .ZN(n4216) );
  INV_X1 U5805 ( .A(n25391), .ZN(n23831) );
  AND2_X1 U5806 ( .A1(n24428), .A2(n4186), .ZN(n4192) );
  AND2_X1 U5807 ( .A1(n25399), .A2(n23860), .ZN(n4186) );
  OR2_X1 U5808 ( .A1(n23861), .A2(n23860), .ZN(n4190) );
  INV_X1 U5810 ( .A(n24006), .ZN(n4478) );
  OR2_X1 U5811 ( .A1(n4478), .A2(n24440), .ZN(n4475) );
  OR2_X1 U5812 ( .A1(n23988), .A2(n23983), .ZN(n23989) );
  OR2_X1 U5813 ( .A1(n23993), .A2(n24006), .ZN(n23979) );
  INV_X1 U5814 ( .A(n24019), .ZN(n24008) );
  NOR2_X1 U5815 ( .A1(n22775), .A2(n22774), .ZN(n5610) );
  AOI21_X1 U5816 ( .B1(n2538), .B2(n23499), .A(n2535), .ZN(n23012) );
  OR2_X1 U5817 ( .A1(n23058), .A2(n22699), .ZN(n3914) );
  NOR2_X1 U5818 ( .A1(n1422), .A2(n23200), .ZN(n4234) );
  OAI21_X1 U5819 ( .B1(n23218), .B2(n23219), .A(n2084), .ZN(n22652) );
  AND2_X1 U5820 ( .A1(n22296), .A2(n23245), .ZN(n3586) );
  OAI21_X1 U5821 ( .B1(n22851), .B2(n2961), .A(n2960), .ZN(n22867) );
  OR2_X1 U5822 ( .A1(n4032), .A2(n924), .ZN(n4029) );
  AND4_X1 U5823 ( .A1(n3441), .A2(n22085), .A3(n22084), .A4(n22083), .ZN(
        Ciphertext[133]) );
  INV_X1 U5824 ( .A(n1815), .ZN(n2588) );
  NOR2_X1 U5825 ( .A1(n24895), .A2(n22043), .ZN(n2590) );
  AND2_X1 U5826 ( .A1(n2475), .A2(n2473), .ZN(n21905) );
  OR2_X1 U5827 ( .A1(n23866), .A2(n24428), .ZN(n4816) );
  AOI21_X1 U5828 ( .B1(n22828), .B2(n25076), .A(n3840), .ZN(n3843) );
  INV_X1 U5829 ( .A(n20975), .ZN(n5131) );
  INV_X1 U5830 ( .A(n17107), .ZN(n4684) );
  XOR2_X1 U5831 ( .A(n14828), .B(n14829), .Z(n1371) );
  INV_X1 U5832 ( .A(n23723), .ZN(n5284) );
  INV_X1 U5833 ( .A(n22354), .ZN(n21844) );
  INV_X1 U5834 ( .A(n16578), .ZN(n2814) );
  INV_X1 U5835 ( .A(n6560), .ZN(n6934) );
  NAND3_X1 U5836 ( .A1(n24474), .A2(n7657), .A3(n7947), .ZN(n1372) );
  INV_X1 U5837 ( .A(n7589), .ZN(n7588) );
  AND3_X1 U5838 ( .A1(n5948), .A2(n5947), .A3(n5949), .ZN(n7589) );
  OR2_X1 U5839 ( .A1(n9805), .A2(n9804), .ZN(n1373) );
  OR2_X1 U5840 ( .A1(n12546), .A2(n12903), .ZN(n1374) );
  INV_X1 U5841 ( .A(n4897), .ZN(n4541) );
  INV_X1 U5842 ( .A(n10746), .ZN(n4341) );
  AND2_X1 U5843 ( .A1(n10811), .A2(n1448), .ZN(n1375) );
  XNOR2_X1 U5845 ( .A(n17992), .B(n17991), .ZN(n2540) );
  XNOR2_X1 U5846 ( .A(n9573), .B(n3360), .ZN(n13092) );
  INV_X1 U5847 ( .A(n13092), .ZN(n12871) );
  AND2_X1 U5848 ( .A1(n12767), .A2(n13216), .ZN(n1376) );
  OR2_X1 U5849 ( .A1(n25198), .A2(n13011), .ZN(n1377) );
  INV_X1 U5850 ( .A(n7382), .ZN(n1895) );
  OR3_X1 U5851 ( .A1(n22941), .A2(n22829), .A3(n22832), .ZN(n1378) );
  INV_X1 U5852 ( .A(n7573), .ZN(n3366) );
  INV_X1 U5853 ( .A(n4880), .ZN(n7651) );
  OR2_X1 U5854 ( .A1(n6719), .A2(n6718), .ZN(n1379) );
  INV_X1 U5856 ( .A(n7580), .ZN(n4136) );
  INV_X1 U5857 ( .A(n23120), .ZN(n5036) );
  INV_X1 U5858 ( .A(n20395), .ZN(n3656) );
  AND2_X1 U5859 ( .A1(n4136), .A2(n7575), .ZN(n1380) );
  INV_X1 U5860 ( .A(n13969), .ZN(n4293) );
  INV_X1 U5861 ( .A(n1535), .ZN(n16615) );
  BUF_X1 U5862 ( .A(n12178), .Z(n13097) );
  INV_X1 U5863 ( .A(n22809), .ZN(n22812) );
  AND2_X1 U5864 ( .A1(n16409), .A2(n14472), .ZN(n1382) );
  INV_X1 U5865 ( .A(n23799), .ZN(n23002) );
  XOR2_X1 U5866 ( .A(n15120), .B(n1951), .Z(n1383) );
  XOR2_X1 U5867 ( .A(n11847), .B(n11846), .Z(n1384) );
  XOR2_X1 U5868 ( .A(n9084), .B(n9083), .Z(n1385) );
  INV_X1 U5869 ( .A(n19613), .ZN(n1806) );
  INV_X1 U5870 ( .A(n13996), .ZN(n13995) );
  INV_X1 U5871 ( .A(n17391), .ZN(n3317) );
  XOR2_X1 U5872 ( .A(n18269), .B(n1835), .Z(n1386) );
  XOR2_X1 U5874 ( .A(n12337), .B(n12336), .Z(n1388) );
  INV_X1 U5875 ( .A(n20588), .ZN(n5093) );
  INV_X1 U5877 ( .A(n22464), .ZN(n3908) );
  INV_X1 U5879 ( .A(n7767), .ZN(n3013) );
  INV_X1 U5880 ( .A(n22387), .ZN(n4109) );
  INV_X1 U5881 ( .A(n8934), .ZN(n10922) );
  INV_X1 U5882 ( .A(n14112), .ZN(n5333) );
  INV_X1 U5883 ( .A(n14850), .ZN(n14416) );
  INV_X1 U5884 ( .A(n17351), .ZN(n17013) );
  OR3_X1 U5885 ( .A1(n11059), .A2(n11058), .A3(n11057), .ZN(n1389) );
  INV_X1 U5888 ( .A(n3671), .ZN(n20279) );
  INV_X1 U5889 ( .A(n22317), .ZN(n2376) );
  INV_X1 U5892 ( .A(n12737), .ZN(n5112) );
  OR3_X1 U5893 ( .A1(n22926), .A2(n25070), .A3(n22188), .ZN(n1390) );
  INV_X1 U5894 ( .A(n6498), .ZN(n6271) );
  INV_X1 U5895 ( .A(n16991), .ZN(n2064) );
  OR2_X1 U5896 ( .A1(n25445), .A2(n13437), .ZN(n1391) );
  AND2_X1 U5898 ( .A1(n16002), .A2(n24366), .ZN(n1392) );
  INV_X1 U5899 ( .A(n19490), .ZN(n5454) );
  OR3_X1 U5900 ( .A1(n405), .A2(n545), .A3(n4499), .ZN(n1393) );
  OR2_X1 U5901 ( .A1(n16817), .A2(n24410), .ZN(n1394) );
  OR2_X1 U5903 ( .A1(n14330), .A2(n14329), .ZN(n1395) );
  OR3_X1 U5904 ( .A1(n22107), .A2(n25070), .A3(n22927), .ZN(n1396) );
  OR3_X1 U5905 ( .A1(n22933), .A2(n22932), .A3(n25004), .ZN(n1397) );
  INV_X1 U5906 ( .A(n22973), .ZN(n3213) );
  INV_X1 U5907 ( .A(n13329), .ZN(n4634) );
  NAND3_X1 U5908 ( .A1(n6690), .A2(n24579), .A3(n6976), .ZN(n1398) );
  OR2_X1 U5909 ( .A1(n9625), .A2(n9681), .ZN(n1399) );
  INV_X1 U5910 ( .A(n22838), .ZN(n2326) );
  INV_X1 U5911 ( .A(n20549), .ZN(n20124) );
  XNOR2_X1 U5912 ( .A(n8201), .B(n8202), .ZN(n10149) );
  INV_X1 U5913 ( .A(n10149), .ZN(n9841) );
  OAI21_X1 U5914 ( .B1(n3709), .B2(n1392), .A(n4515), .ZN(n16607) );
  INV_X1 U5916 ( .A(n13871), .ZN(n3401) );
  INV_X1 U5917 ( .A(n16221), .ZN(n16461) );
  OR2_X1 U5918 ( .A1(n10680), .A2(n4737), .ZN(n1401) );
  OR2_X1 U5919 ( .A1(n7081), .A2(n7943), .ZN(n1402) );
  XNOR2_X1 U5920 ( .A(n18145), .B(n4214), .ZN(n2464) );
  INV_X1 U5921 ( .A(n2464), .ZN(n3412) );
  OR2_X1 U5922 ( .A1(n4069), .A2(n10047), .ZN(n1403) );
  INV_X1 U5923 ( .A(n8477), .ZN(n2191) );
  INV_X1 U5924 ( .A(n12607), .ZN(n13266) );
  XNOR2_X1 U5925 ( .A(n12001), .B(n12000), .ZN(n12607) );
  INV_X1 U5926 ( .A(n7733), .ZN(n5432) );
  XNOR2_X1 U5927 ( .A(n8438), .B(n8437), .ZN(n10079) );
  INV_X1 U5928 ( .A(n16096), .ZN(n4418) );
  OAI211_X1 U5929 ( .C1(n19376), .C2(n19222), .A(n5441), .B(n5442), .ZN(n20140) );
  OAI211_X1 U5930 ( .C1(n4543), .C2(n19022), .A(n4542), .B(n19629), .ZN(n19975) );
  INV_X1 U5931 ( .A(n19975), .ZN(n20298) );
  INV_X1 U5932 ( .A(n17572), .ZN(n3371) );
  INV_X1 U5933 ( .A(n9281), .ZN(n9963) );
  XNOR2_X1 U5934 ( .A(n4182), .B(n12271), .ZN(n12865) );
  XNOR2_X1 U5935 ( .A(n18712), .B(n18711), .ZN(n22257) );
  AND3_X1 U5937 ( .A1(n19112), .A2(n19233), .A3(n19608), .ZN(n1404) );
  OR2_X1 U5938 ( .A1(n7912), .A2(n7364), .ZN(n1405) );
  INV_X1 U5939 ( .A(n9964), .ZN(n3290) );
  INV_X1 U5940 ( .A(n20422), .ZN(n1662) );
  AND2_X1 U5941 ( .A1(n9806), .A2(n9807), .ZN(n1406) );
  OR3_X1 U5942 ( .A1(n14003), .A2(n13486), .A3(n14000), .ZN(n1407) );
  INV_X1 U5943 ( .A(n12861), .ZN(n5412) );
  INV_X1 U5944 ( .A(n6848), .ZN(n4643) );
  XOR2_X1 U5945 ( .A(n18557), .B(n18043), .Z(n1408) );
  XNOR2_X1 U5946 ( .A(n8248), .B(n8247), .ZN(n10177) );
  XNOR2_X1 U5947 ( .A(n21518), .B(n21519), .ZN(n22946) );
  XNOR2_X1 U5948 ( .A(n14673), .B(n14674), .ZN(n16108) );
  INV_X1 U5949 ( .A(n16108), .ZN(n2090) );
  XNOR2_X1 U5951 ( .A(n10530), .B(n10529), .ZN(n13165) );
  XOR2_X1 U5952 ( .A(n18489), .B(n5286), .Z(n1410) );
  XOR2_X1 U5953 ( .A(n14897), .B(n21944), .Z(n1411) );
  INV_X1 U5955 ( .A(n6955), .ZN(n3926) );
  XNOR2_X1 U5957 ( .A(n17793), .B(n17794), .ZN(n19365) );
  INV_X1 U5958 ( .A(n20517), .ZN(n3522) );
  INV_X1 U5959 ( .A(n17276), .ZN(n17274) );
  INV_X1 U5960 ( .A(n18597), .ZN(n19179) );
  AND3_X1 U5961 ( .A1(n7855), .A2(n24072), .A3(n7721), .ZN(n1413) );
  NAND3_X1 U5962 ( .A1(n4838), .A2(n3142), .A3(n6003), .ZN(n7893) );
  XOR2_X1 U5963 ( .A(n8588), .B(n1776), .Z(n1414) );
  OR2_X1 U5964 ( .A1(n15625), .A2(n16147), .ZN(n1415) );
  INV_X1 U5965 ( .A(n11529), .ZN(n11026) );
  INV_X1 U5966 ( .A(n7862), .ZN(n4536) );
  OR3_X1 U5967 ( .A1(n17421), .A2(n17425), .A3(n17424), .ZN(n1416) );
  OR2_X1 U5968 ( .A1(n21852), .A2(n22656), .ZN(n1417) );
  INV_X1 U5969 ( .A(n24572), .ZN(n4225) );
  INV_X1 U5971 ( .A(n20042), .ZN(n19862) );
  AND2_X1 U5972 ( .A1(n10993), .A2(n10990), .ZN(n1418) );
  XNOR2_X1 U5973 ( .A(n20709), .B(n20710), .ZN(n22562) );
  XNOR2_X1 U5974 ( .A(n18084), .B(n5135), .ZN(n18808) );
  AND2_X1 U5975 ( .A1(n19301), .A2(n19300), .ZN(n1419) );
  INV_X1 U5976 ( .A(n20597), .ZN(n5044) );
  OR2_X1 U5977 ( .A1(n20480), .A2(n20478), .ZN(n1420) );
  XNOR2_X1 U5978 ( .A(n14648), .B(n14647), .ZN(n16073) );
  OR2_X1 U5979 ( .A1(n5572), .A2(n19277), .ZN(n1421) );
  OR2_X1 U5980 ( .A1(n24889), .A2(n23201), .ZN(n1422) );
  OR2_X1 U5981 ( .A1(n19587), .A2(n24483), .ZN(n1423) );
  INV_X1 U5982 ( .A(n16434), .ZN(n17170) );
  AND2_X1 U5983 ( .A1(n20593), .A2(n20590), .ZN(n1424) );
  OR2_X1 U5984 ( .A1(n19013), .A2(n19436), .ZN(n1425) );
  OR2_X1 U5985 ( .A1(n19584), .A2(n19105), .ZN(n1426) );
  OR2_X1 U5986 ( .A1(n19277), .A2(n19126), .ZN(n1427) );
  NAND2_X1 U5987 ( .A1(n1642), .A2(n5574), .ZN(n7731) );
  INV_X1 U5988 ( .A(n7731), .ZN(n5595) );
  AND2_X1 U5989 ( .A1(n22656), .A2(n22606), .ZN(n1428) );
  OR2_X1 U5990 ( .A1(n19408), .A2(n19413), .ZN(n1429) );
  AND2_X1 U5991 ( .A1(n10596), .A2(n10935), .ZN(n1430) );
  AND2_X1 U5992 ( .A1(n22901), .A2(n22847), .ZN(n1431) );
  AND2_X1 U5993 ( .A1(n20019), .A2(n18985), .ZN(n1432) );
  INV_X1 U5994 ( .A(n2321), .ZN(n14090) );
  OAI211_X1 U5995 ( .C1(n12501), .C2(n13148), .A(n2575), .B(n2574), .ZN(n2321)
         );
  AND3_X1 U5996 ( .A1(n6241), .A2(n6242), .A3(n6240), .ZN(n1433) );
  AND2_X1 U5997 ( .A1(n16359), .A2(n16355), .ZN(n1434) );
  OR3_X1 U5998 ( .A1(n22505), .A2(n25063), .A3(n22722), .ZN(n1435) );
  OR2_X1 U5999 ( .A1(n19396), .A2(n19397), .ZN(n1436) );
  OR3_X1 U6000 ( .A1(n25572), .A2(n16846), .A3(n5052), .ZN(n1437) );
  OR3_X1 U6001 ( .A1(n20518), .A2(n20517), .A3(n20516), .ZN(n1438) );
  INV_X1 U6002 ( .A(n10571), .ZN(n3760) );
  INV_X1 U6003 ( .A(n22528), .ZN(n3242) );
  AND2_X1 U6004 ( .A1(n12471), .A2(n12773), .ZN(n1439) );
  INV_X1 U6005 ( .A(n7890), .ZN(n7606) );
  OR2_X1 U6006 ( .A1(n24311), .A2(n22323), .ZN(n1440) );
  INV_X1 U6007 ( .A(n13235), .ZN(n12546) );
  AND2_X1 U6008 ( .A1(n6729), .A2(n6732), .ZN(n1441) );
  OR2_X1 U6009 ( .A1(n23690), .A2(n23689), .ZN(n1442) );
  INV_X1 U6010 ( .A(n20136), .ZN(n1954) );
  INV_X1 U6011 ( .A(n23595), .ZN(n23591) );
  OR2_X1 U6012 ( .A1(n15670), .A2(n15915), .ZN(n1444) );
  BUF_X1 U6013 ( .A(n5888), .Z(n6940) );
  INV_X1 U6015 ( .A(n11116), .ZN(n11111) );
  OR2_X1 U6016 ( .A1(n14509), .A2(n14440), .ZN(n1446) );
  AND2_X1 U6017 ( .A1(n11159), .A2(n11158), .ZN(n1447) );
  OR2_X1 U6018 ( .A1(n10670), .A2(n11214), .ZN(n1448) );
  AND2_X1 U6019 ( .A1(n20126), .A2(n20124), .ZN(n1449) );
  NOR2_X1 U6020 ( .A1(n24588), .A2(n14303), .ZN(n1450) );
  AND2_X1 U6021 ( .A1(n17180), .A2(n17181), .ZN(n1451) );
  OR2_X1 U6022 ( .A1(n20437), .A2(n24940), .ZN(n1452) );
  AND2_X1 U6024 ( .A1(n9765), .A2(n9766), .ZN(n1453) );
  INV_X1 U6025 ( .A(n17305), .ZN(n3783) );
  INV_X1 U6026 ( .A(n21828), .ZN(n3201) );
  AND2_X1 U6027 ( .A1(n7588), .A2(n5971), .ZN(n1454) );
  OR2_X1 U6028 ( .A1(n3480), .A2(n20328), .ZN(n1455) );
  OR2_X1 U6029 ( .A1(n13316), .A2(n12945), .ZN(n1456) );
  AND2_X1 U6030 ( .A1(n331), .A2(n22656), .ZN(n1457) );
  INV_X1 U6032 ( .A(n12928), .ZN(n5672) );
  INV_X1 U6033 ( .A(n23714), .ZN(n23716) );
  OR2_X1 U6034 ( .A1(n13552), .A2(n24376), .ZN(n1459) );
  XNOR2_X1 U6036 ( .A(n7356), .B(n7355), .ZN(n10125) );
  INV_X1 U6037 ( .A(n10125), .ZN(n5057) );
  AND2_X1 U6038 ( .A1(n9695), .A2(n9699), .ZN(n1460) );
  XOR2_X1 U6039 ( .A(n21743), .B(n860), .Z(n1461) );
  NOR2_X1 U6040 ( .A1(n23730), .A2(n24991), .ZN(n1462) );
  INV_X1 U6041 ( .A(n11178), .ZN(n3386) );
  AND2_X1 U6042 ( .A1(n8318), .A2(n8319), .ZN(n1463) );
  OR2_X1 U6043 ( .A1(n25064), .A2(n1577), .ZN(n1464) );
  INV_X1 U6044 ( .A(n14306), .ZN(n1527) );
  INV_X1 U6045 ( .A(n20272), .ZN(n20520) );
  OR2_X1 U6047 ( .A1(n23969), .A2(n23972), .ZN(n1465) );
  NOR2_X1 U6049 ( .A1(n22159), .A2(n22158), .ZN(n1467) );
  INV_X1 U6050 ( .A(n19381), .ZN(n19377) );
  AND2_X1 U6051 ( .A1(n13088), .A2(n13394), .ZN(n14359) );
  AND2_X1 U6052 ( .A1(n7506), .A2(n1379), .ZN(n1468) );
  OR2_X1 U6053 ( .A1(n20073), .A2(n20072), .ZN(n1469) );
  INV_X1 U6055 ( .A(n17379), .ZN(n5406) );
  OR2_X1 U6056 ( .A1(n12793), .A2(n12792), .ZN(n1471) );
  OR2_X1 U6057 ( .A1(n15937), .A2(n24387), .ZN(n1472) );
  AND2_X1 U6058 ( .A1(n17298), .A2(n1535), .ZN(n1473) );
  INV_X1 U6059 ( .A(n12540), .ZN(n13220) );
  INV_X1 U6060 ( .A(n11755), .ZN(n12885) );
  INV_X1 U6061 ( .A(n7590), .ZN(n2035) );
  AND2_X1 U6062 ( .A1(n14462), .A2(n3501), .ZN(n1474) );
  INV_X1 U6063 ( .A(n7211), .ZN(n7666) );
  NAND2_X1 U6064 ( .A1(n4179), .A2(n13173), .ZN(n14107) );
  NAND3_X1 U6065 ( .A1(n19272), .A2(n19530), .A3(n1013), .ZN(n1475) );
  INV_X1 U6066 ( .A(n4754), .ZN(n4752) );
  INV_X1 U6067 ( .A(n17872), .ZN(n18945) );
  BUF_X1 U6068 ( .A(n17872), .Z(n19471) );
  INV_X1 U6069 ( .A(n22459), .ZN(n22463) );
  OR2_X1 U6070 ( .A1(n25058), .A2(n17362), .ZN(n1476) );
  NOR2_X1 U6071 ( .A1(n25075), .A2(n22655), .ZN(n1477) );
  OR2_X1 U6072 ( .A1(n22928), .A2(n24379), .ZN(n1478) );
  INV_X1 U6073 ( .A(n17970), .ZN(n5300) );
  INV_X1 U6074 ( .A(n2556), .ZN(n5487) );
  OR2_X1 U6075 ( .A1(n9236), .A2(n9416), .ZN(n1479) );
  NAND2_X1 U6076 ( .A1(n22490), .A2(n25055), .ZN(n1480) );
  OR2_X1 U6077 ( .A1(n11121), .A2(n11123), .ZN(n1481) );
  NAND2_X1 U6078 ( .A1(n22254), .A2(n21822), .ZN(n1482) );
  OR2_X1 U6079 ( .A1(n15646), .A2(n25500), .ZN(n1483) );
  OR2_X1 U6080 ( .A1(n20343), .A2(n20277), .ZN(n1484) );
  OR2_X1 U6081 ( .A1(n7782), .A2(n7418), .ZN(n1485) );
  OR2_X1 U6083 ( .A1(n20190), .A2(n20191), .ZN(n1487) );
  BUF_X1 U6084 ( .A(n15674), .Z(n16328) );
  AND2_X1 U6085 ( .A1(n24954), .A2(n23993), .ZN(n1488) );
  INV_X1 U6086 ( .A(n14143), .ZN(n5641) );
  INV_X1 U6087 ( .A(n8527), .ZN(n7087) );
  INV_X1 U6088 ( .A(n13549), .ZN(n14204) );
  INV_X1 U6089 ( .A(n13569), .ZN(n13589) );
  AND2_X1 U6091 ( .A1(n19964), .A2(n349), .ZN(n1489) );
  INV_X1 U6092 ( .A(n10548), .ZN(n10702) );
  BUF_X1 U6093 ( .A(n12663), .Z(n13152) );
  INV_X1 U6094 ( .A(n13968), .ZN(n1771) );
  INV_X1 U6095 ( .A(n23327), .ZN(n5659) );
  INV_X1 U6096 ( .A(n20400), .ZN(n20417) );
  AND2_X1 U6097 ( .A1(n7693), .A2(n7694), .ZN(n1490) );
  OR2_X1 U6098 ( .A1(n24498), .A2(n5131), .ZN(n1491) );
  INV_X1 U6099 ( .A(n20091), .ZN(n2368) );
  NAND2_X1 U6100 ( .A1(n16990), .A2(n17039), .ZN(n1492) );
  AND2_X1 U6101 ( .A1(n20368), .A2(n20373), .ZN(n3767) );
  INV_X1 U6102 ( .A(n14319), .ZN(n4794) );
  OR2_X1 U6103 ( .A1(n18912), .A2(n19138), .ZN(n1493) );
  INV_X1 U6104 ( .A(n924), .ZN(n4034) );
  AND2_X1 U6105 ( .A1(n5353), .A2(n5354), .ZN(n1494) );
  OR2_X1 U6106 ( .A1(n11342), .A2(n3344), .ZN(n1495) );
  INV_X1 U6107 ( .A(n21964), .ZN(n2319) );
  INV_X1 U6108 ( .A(n21046), .ZN(n4023) );
  INV_X1 U6109 ( .A(n2137), .ZN(n4668) );
  INV_X1 U6110 ( .A(n925), .ZN(n5433) );
  INV_X1 U6111 ( .A(n3155), .ZN(n3901) );
  INV_X1 U6112 ( .A(n888), .ZN(n1528) );
  INV_X1 U6113 ( .A(n4711), .ZN(n3344) );
  INV_X1 U6114 ( .A(n22089), .ZN(n5286) );
  INV_X1 U6115 ( .A(n853), .ZN(n4153) );
  INV_X1 U6116 ( .A(n1831), .ZN(n4761) );
  INV_X1 U6117 ( .A(n677), .ZN(n5514) );
  INV_X1 U6118 ( .A(n2034), .ZN(n3900) );
  INV_X1 U6119 ( .A(n763), .ZN(n2964) );
  INV_X1 U6120 ( .A(n3152), .ZN(n5251) );
  INV_X1 U6121 ( .A(n1935), .ZN(n4589) );
  INV_X1 U6122 ( .A(n2970), .ZN(n5598) );
  INV_X1 U6123 ( .A(n2743), .ZN(n3208) );
  INV_X1 U6124 ( .A(Key[41]), .ZN(n3696) );
  NAND2_X1 U6125 ( .A1(n1497), .A2(n1496), .ZN(n17184) );
  OAI21_X1 U6126 ( .B1(n16208), .B2(n16209), .A(n16207), .ZN(n1496) );
  NOR2_X1 U6127 ( .A1(n17182), .A2(n17183), .ZN(n1498) );
  NAND2_X1 U6128 ( .A1(n10753), .A2(n1499), .ZN(n4506) );
  NAND2_X1 U6129 ( .A1(n4505), .A2(n1499), .ZN(n4507) );
  NAND2_X1 U6130 ( .A1(n10452), .A2(n1499), .ZN(n10290) );
  AND2_X1 U6131 ( .A1(n10455), .A2(n1499), .ZN(n2385) );
  NAND2_X1 U6132 ( .A1(n23334), .A2(n24341), .ZN(n1500) );
  XNOR2_X2 U6133 ( .A(n21396), .B(n21397), .ZN(n23334) );
  NAND2_X1 U6135 ( .A1(n4052), .A2(n18862), .ZN(n19080) );
  NAND2_X1 U6137 ( .A1(n19361), .A2(n24447), .ZN(n1506) );
  AND2_X1 U6138 ( .A1(n25392), .A2(n24312), .ZN(n1505) );
  INV_X1 U6140 ( .A(n4442), .ZN(n1507) );
  NAND2_X1 U6141 ( .A1(n12827), .A2(n25466), .ZN(n1508) );
  NAND2_X1 U6142 ( .A1(n14457), .A2(n4794), .ZN(n14460) );
  OR2_X1 U6143 ( .A1(n1509), .A2(n25398), .ZN(n5698) );
  INV_X1 U6144 ( .A(n6523), .ZN(n1509) );
  AND2_X1 U6145 ( .A1(n16350), .A2(n1511), .ZN(n16598) );
  OAI21_X1 U6146 ( .B1(n24890), .B2(n16595), .A(n24080), .ZN(n1510) );
  NAND3_X1 U6147 ( .A1(n15885), .A2(n15890), .A3(n24587), .ZN(n1511) );
  NOR2_X1 U6148 ( .A1(n24587), .A2(n16597), .ZN(n1512) );
  NAND2_X1 U6149 ( .A1(n1513), .A2(n13116), .ZN(n2097) );
  NOR2_X1 U6150 ( .A1(n3328), .A2(n12272), .ZN(n1513) );
  NOR2_X1 U6151 ( .A1(n22800), .A2(n1514), .ZN(n22659) );
  NOR2_X1 U6152 ( .A1(n12942), .A2(n1515), .ZN(n11921) );
  NAND2_X1 U6153 ( .A1(n1515), .A2(n13317), .ZN(n13321) );
  INV_X1 U6154 ( .A(n4241), .ZN(n1515) );
  NAND2_X1 U6156 ( .A1(n1516), .A2(n2562), .ZN(n5316) );
  NAND2_X1 U6157 ( .A1(n1516), .A2(n16901), .ZN(n17474) );
  INV_X1 U6158 ( .A(n9694), .ZN(n1517) );
  INV_X1 U6159 ( .A(n2294), .ZN(n9875) );
  NAND2_X1 U6160 ( .A1(n1520), .A2(n1518), .ZN(n10534) );
  NAND2_X1 U6162 ( .A1(n19117), .A2(n1522), .ZN(n1521) );
  INV_X1 U6163 ( .A(n11057), .ZN(n1523) );
  NAND2_X1 U6164 ( .A1(n1524), .A2(n11059), .ZN(n10697) );
  NOR2_X1 U6165 ( .A1(n1218), .A2(n11057), .ZN(n1524) );
  AND2_X1 U6167 ( .A1(n24588), .A2(n14301), .ZN(n12018) );
  NAND2_X1 U6169 ( .A1(n3352), .A2(n4144), .ZN(n1530) );
  NAND2_X1 U6170 ( .A1(n1531), .A2(n431), .ZN(n3352) );
  NAND4_X1 U6172 ( .A1(n5273), .A2(n1532), .A3(n5274), .A4(n5271), .ZN(n10477)
         );
  NAND2_X1 U6173 ( .A1(n9127), .A2(n10064), .ZN(n1534) );
  OR2_X1 U6174 ( .A1(n1535), .A2(n17296), .ZN(n16513) );
  NOR2_X1 U6175 ( .A1(n1535), .A2(n17299), .ZN(n16706) );
  OR2_X1 U6176 ( .A1(n4508), .A2(n1535), .ZN(n16703) );
  NAND3_X1 U6177 ( .A1(n1541), .A2(n13643), .A3(n1536), .ZN(n13648) );
  NAND3_X1 U6178 ( .A1(n1538), .A2(n13079), .A3(n1537), .ZN(n1536) );
  NAND3_X1 U6179 ( .A1(n1540), .A2(n13079), .A3(n1539), .ZN(n13818) );
  NAND2_X1 U6180 ( .A1(n1543), .A2(n4340), .ZN(n1540) );
  NAND2_X1 U6181 ( .A1(n1542), .A2(n13079), .ZN(n1541) );
  INV_X1 U6182 ( .A(n4340), .ZN(n1542) );
  NAND2_X1 U6183 ( .A1(n13069), .A2(n13070), .ZN(n1543) );
  NOR2_X1 U6184 ( .A1(n3423), .A2(n1545), .ZN(n3422) );
  XNOR2_X2 U6185 ( .A(n4316), .B(n11617), .ZN(n13048) );
  XNOR2_X2 U6186 ( .A(n11605), .B(n11606), .ZN(n13049) );
  NAND2_X1 U6187 ( .A1(n1546), .A2(n17042), .ZN(n3372) );
  AOI21_X1 U6188 ( .B1(n17572), .B2(n1546), .A(n3004), .ZN(n3003) );
  XNOR2_X2 U6189 ( .A(Plaintext[29]), .B(Key[29]), .ZN(n6531) );
  MUX2_X1 U6190 ( .A(n18881), .B(n18880), .S(n2464), .Z(n1547) );
  NAND2_X1 U6192 ( .A1(n2069), .A2(n3412), .ZN(n1548) );
  NAND2_X1 U6193 ( .A1(n17224), .A2(n1549), .ZN(n2324) );
  AND2_X1 U6194 ( .A1(n25433), .A2(n17225), .ZN(n1549) );
  NAND2_X1 U6197 ( .A1(n6434), .A2(n6498), .ZN(n6168) );
  AND2_X1 U6198 ( .A1(n20909), .A2(n20491), .ZN(n1550) );
  XNOR2_X2 U6199 ( .A(n7654), .B(n7655), .ZN(n9599) );
  OR2_X1 U6200 ( .A1(n3353), .A2(n13829), .ZN(n13556) );
  OR2_X1 U6201 ( .A1(n4545), .A2(n7932), .ZN(n2164) );
  AND2_X1 U6202 ( .A1(n7924), .A2(n7932), .ZN(n5606) );
  AND2_X1 U6203 ( .A1(n4380), .A2(n4379), .ZN(n1554) );
  OR2_X1 U6204 ( .A1(n6789), .A2(n6905), .ZN(n5247) );
  INV_X1 U6205 ( .A(n7007), .ZN(n7005) );
  INV_X1 U6206 ( .A(n14242), .ZN(n13633) );
  INV_X1 U6208 ( .A(n4436), .ZN(n19265) );
  INV_X1 U6209 ( .A(n16397), .ZN(n3630) );
  INV_X1 U6210 ( .A(n7803), .ZN(n7795) );
  NOR2_X1 U6211 ( .A1(n441), .A2(n6271), .ZN(n5143) );
  OR2_X1 U6212 ( .A1(n5707), .A2(n25433), .ZN(n4572) );
  AND2_X1 U6213 ( .A1(n25450), .A2(n1363), .ZN(n21928) );
  INV_X1 U6215 ( .A(n16220), .ZN(n5269) );
  OR2_X1 U6217 ( .A1(n16901), .A2(n16902), .ZN(n2247) );
  XNOR2_X1 U6218 ( .A(n18285), .B(n18685), .ZN(n18372) );
  INV_X1 U6219 ( .A(n15746), .ZN(n1654) );
  OR2_X1 U6220 ( .A1(n24540), .A2(n25441), .ZN(n4926) );
  OAI211_X1 U6221 ( .C1(n9857), .C2(n9864), .A(n25464), .B(n4622), .ZN(n10517)
         );
  INV_X1 U6223 ( .A(n2404), .ZN(n7085) );
  AND2_X1 U6224 ( .A1(n7013), .A2(n6827), .ZN(n1876) );
  OR2_X1 U6225 ( .A1(n23281), .A2(n24349), .ZN(n5529) );
  OR2_X1 U6226 ( .A1(n24411), .A2(n22962), .ZN(n22964) );
  INV_X1 U6227 ( .A(n22967), .ZN(n21476) );
  OR2_X1 U6228 ( .A1(n2587), .A2(n16550), .ZN(n2508) );
  INV_X1 U6229 ( .A(n16550), .ZN(n16794) );
  OR2_X1 U6230 ( .A1(n16550), .A2(n16796), .ZN(n16619) );
  OR2_X1 U6231 ( .A1(n12648), .A2(n12178), .ZN(n5321) );
  AND2_X1 U6232 ( .A1(n24549), .A2(n9692), .ZN(n9028) );
  OR2_X1 U6233 ( .A1(n24549), .A2(n9027), .ZN(n3117) );
  XNOR2_X1 U6234 ( .A(n1813), .B(n8789), .ZN(n8549) );
  INV_X1 U6235 ( .A(n8366), .ZN(n1813) );
  XNOR2_X1 U6236 ( .A(n21215), .B(n20223), .ZN(n3871) );
  INV_X1 U6238 ( .A(n24547), .ZN(n4334) );
  OR2_X1 U6239 ( .A1(n6444), .A2(n6445), .ZN(n6021) );
  OR2_X1 U6240 ( .A1(n23069), .A2(n23064), .ZN(n4990) );
  OR2_X1 U6241 ( .A1(n12652), .A2(n403), .ZN(n3935) );
  OR2_X1 U6243 ( .A1(n25477), .A2(n20597), .ZN(n5365) );
  XNOR2_X1 U6244 ( .A(n11309), .B(n3647), .ZN(n12792) );
  OAI21_X1 U6245 ( .B1(n7893), .B2(n7604), .A(n7606), .ZN(n7326) );
  NOR2_X1 U6246 ( .A1(n9782), .A2(n9781), .ZN(n9676) );
  AND2_X1 U6247 ( .A1(n2718), .A2(n15811), .ZN(n3316) );
  INV_X1 U6248 ( .A(n13888), .ZN(n13945) );
  OAI21_X1 U6249 ( .B1(n9064), .B2(n10050), .A(n9866), .ZN(n9869) );
  AOI21_X1 U6250 ( .B1(n9064), .B2(n9244), .A(n24446), .ZN(n3489) );
  AND2_X1 U6251 ( .A1(n9064), .A2(n24092), .ZN(n10054) );
  AND2_X1 U6253 ( .A1(n3195), .A2(n19939), .ZN(n19817) );
  AND2_X1 U6254 ( .A1(n19302), .A2(n19133), .ZN(n3568) );
  NOR2_X1 U6255 ( .A1(n388), .A2(n15667), .ZN(n15917) );
  OR2_X1 U6256 ( .A1(n14510), .A2(n13974), .ZN(n3777) );
  INV_X1 U6257 ( .A(n13974), .ZN(n14436) );
  NOR2_X1 U6258 ( .A1(n13161), .A2(n12454), .ZN(n5013) );
  AND2_X1 U6259 ( .A1(n23869), .A2(n23905), .ZN(n23888) );
  NOR2_X1 U6260 ( .A1(n25414), .A2(n25079), .ZN(n2616) );
  AND2_X1 U6262 ( .A1(n25001), .A2(n19598), .ZN(n4715) );
  OR2_X1 U6264 ( .A1(n6775), .A2(n6292), .ZN(n6293) );
  OR2_X1 U6265 ( .A1(n6775), .A2(n6777), .ZN(n2353) );
  NOR2_X1 U6266 ( .A1(n10464), .A2(n10720), .ZN(n4500) );
  AOI22_X1 U6267 ( .A1(n7827), .A2(n7985), .B1(n7984), .B2(n7046), .ZN(n7513)
         );
  AND2_X1 U6268 ( .A1(n7985), .A2(n7983), .ZN(n1690) );
  OR2_X1 U6269 ( .A1(n7827), .A2(n7985), .ZN(n2082) );
  INV_X1 U6270 ( .A(n21140), .ZN(n22779) );
  INV_X1 U6271 ( .A(n18290), .ZN(n17637) );
  OR2_X1 U6272 ( .A1(n3472), .A2(n10125), .ZN(n9379) );
  XNOR2_X1 U6273 ( .A(n15267), .B(n15160), .ZN(n3669) );
  AND2_X1 U6275 ( .A1(n24321), .A2(n23303), .ZN(n23300) );
  OR2_X1 U6276 ( .A1(n24321), .A2(n23303), .ZN(n3623) );
  OR2_X1 U6277 ( .A1(n20255), .A2(n25421), .ZN(n5189) );
  NOR2_X1 U6278 ( .A1(n18895), .A2(n19526), .ZN(n19720) );
  OAI22_X1 U6279 ( .A1(n5003), .A2(n18795), .B1(n19526), .B2(n5496), .ZN(
        n19528) );
  INV_X1 U6280 ( .A(n19526), .ZN(n19283) );
  OR2_X1 U6282 ( .A1(n22868), .A2(n23411), .ZN(n2961) );
  AND2_X1 U6283 ( .A1(n24421), .A2(n19290), .ZN(n3094) );
  INV_X1 U6284 ( .A(n12792), .ZN(n4680) );
  AND2_X1 U6285 ( .A1(n13228), .A2(n12792), .ZN(n13229) );
  AND2_X1 U6286 ( .A1(n12792), .A2(n12995), .ZN(n2837) );
  OR2_X1 U6287 ( .A1(n7008), .A2(n7004), .ZN(n6833) );
  XNOR2_X1 U6288 ( .A(n24413), .B(n8981), .ZN(n8183) );
  OR2_X1 U6289 ( .A1(n22162), .A2(n22221), .ZN(n21830) );
  OAI21_X1 U6290 ( .B1(n18994), .B2(n20316), .A(n20319), .ZN(n2179) );
  AND2_X1 U6291 ( .A1(n12993), .A2(n4587), .ZN(n13230) );
  OR2_X1 U6292 ( .A1(n12791), .A2(n12993), .ZN(n5041) );
  OR2_X1 U6293 ( .A1(n9449), .A2(n9907), .ZN(n9936) );
  AND2_X1 U6294 ( .A1(n23273), .A2(n25550), .ZN(n22535) );
  AND2_X1 U6296 ( .A1(n22409), .A2(n22407), .ZN(n22133) );
  OR2_X1 U6297 ( .A1(n22562), .A2(n22407), .ZN(n1588) );
  OR2_X1 U6298 ( .A1(n16109), .A2(n16108), .ZN(n2020) );
  INV_X1 U6299 ( .A(n12272), .ZN(n13113) );
  OR2_X1 U6300 ( .A1(n6795), .A2(n6076), .ZN(n3894) );
  OR2_X1 U6301 ( .A1(n23555), .A2(n23546), .ZN(n5397) );
  INV_X1 U6302 ( .A(n16452), .ZN(n16235) );
  NOR2_X1 U6303 ( .A1(n12785), .A2(n13027), .ZN(n1635) );
  INV_X1 U6304 ( .A(n12785), .ZN(n13029) );
  OAI21_X1 U6305 ( .B1(n20963), .B2(n24354), .A(n20962), .ZN(n21452) );
  INV_X1 U6306 ( .A(n16192), .ZN(n16196) );
  XNOR2_X1 U6307 ( .A(n15218), .B(n14955), .ZN(n2862) );
  AND2_X1 U6312 ( .A1(n16266), .A2(n25009), .ZN(n5667) );
  OAI22_X1 U6313 ( .A1(n3287), .A2(n12824), .B1(n13288), .B2(n13289), .ZN(
        n13297) );
  XNOR2_X1 U6314 ( .A(n15430), .B(n15523), .ZN(n15106) );
  OR2_X1 U6315 ( .A1(n16356), .A2(n16290), .ZN(n4846) );
  OAI21_X1 U6316 ( .B1(n3517), .B2(n367), .A(n3514), .ZN(n3706) );
  AOI22_X1 U6317 ( .A1(n17356), .A2(n17351), .B1(n17012), .B2(n25491), .ZN(
        n3517) );
  XNOR2_X1 U6318 ( .A(n21601), .B(n21675), .ZN(n21023) );
  AND2_X1 U6319 ( .A1(n19366), .A2(n19370), .ZN(n19098) );
  NOR2_X1 U6321 ( .A1(n12459), .A2(n12724), .ZN(n3968) );
  NOR2_X1 U6323 ( .A1(n8021), .A2(n7278), .ZN(n3259) );
  INV_X1 U6324 ( .A(n24415), .ZN(n4350) );
  OAI211_X1 U6326 ( .C1(n13119), .C2(n12660), .A(n2571), .B(n12865), .ZN(
        n12422) );
  INV_X1 U6327 ( .A(n9989), .ZN(n9747) );
  INV_X1 U6329 ( .A(n18982), .ZN(n20137) );
  OR2_X1 U6330 ( .A1(n3822), .A2(n17607), .ZN(n16941) );
  OR2_X1 U6332 ( .A1(n22099), .A2(n22729), .ZN(n2981) );
  INV_X1 U6333 ( .A(n22729), .ZN(n3837) );
  INV_X1 U6334 ( .A(n19300), .ZN(n18970) );
  INV_X1 U6335 ( .A(n2607), .ZN(n16229) );
  AND2_X1 U6336 ( .A1(n16492), .A2(n24387), .ZN(n5169) );
  OR2_X1 U6337 ( .A1(n10007), .A2(n9484), .ZN(n9722) );
  OR2_X1 U6338 ( .A1(n6814), .A2(n6815), .ZN(n2800) );
  NAND2_X1 U6339 ( .A1(n18763), .A2(n4172), .ZN(n1556) );
  NAND3_X1 U6340 ( .A1(n1733), .A2(n20343), .A3(n1557), .ZN(n19650) );
  NAND2_X1 U6341 ( .A1(n1558), .A2(n4752), .ZN(n1862) );
  NAND2_X1 U6342 ( .A1(n4752), .A2(n1559), .ZN(n6406) );
  OAI21_X1 U6344 ( .B1(n8146), .B2(n10927), .A(n1562), .ZN(n10408) );
  NAND2_X1 U6345 ( .A1(n10407), .A2(n10927), .ZN(n1562) );
  NAND3_X1 U6346 ( .A1(n13349), .A2(n13346), .A3(n12861), .ZN(n2023) );
  NAND2_X1 U6347 ( .A1(n6937), .A2(n1563), .ZN(n6562) );
  NAND2_X1 U6348 ( .A1(n6559), .A2(n6934), .ZN(n1563) );
  INV_X1 U6349 ( .A(n12611), .ZN(n13304) );
  NAND2_X1 U6352 ( .A1(n13304), .A2(n12555), .ZN(n1566) );
  INV_X1 U6354 ( .A(n12555), .ZN(n13303) );
  XNOR2_X1 U6355 ( .A(n1568), .B(n3093), .ZN(n11336) );
  XNOR2_X1 U6356 ( .A(n1568), .B(n2881), .ZN(n12010) );
  XNOR2_X1 U6357 ( .A(n1568), .B(n14398), .ZN(n10706) );
  XNOR2_X1 U6358 ( .A(n1568), .B(n2782), .ZN(n11483) );
  XNOR2_X1 U6359 ( .A(n1568), .B(n12314), .ZN(n11614) );
  XNOR2_X1 U6360 ( .A(n1568), .B(n12391), .ZN(n12392) );
  OAI21_X1 U6361 ( .B1(n11038), .B2(n10942), .A(n1569), .ZN(n11040) );
  NAND2_X1 U6362 ( .A1(n10941), .A2(n11036), .ZN(n1569) );
  NAND2_X1 U6363 ( .A1(n11037), .A2(n11036), .ZN(n1570) );
  NAND2_X1 U6364 ( .A1(n10571), .A2(n10941), .ZN(n11037) );
  NAND2_X1 U6366 ( .A1(n12689), .A2(n12946), .ZN(n1572) );
  NAND2_X1 U6367 ( .A1(n7634), .A2(n1573), .ZN(n7160) );
  NAND2_X1 U6368 ( .A1(n1574), .A2(n25253), .ZN(n1573) );
  NAND2_X1 U6369 ( .A1(n7915), .A2(n7917), .ZN(n1574) );
  NAND3_X1 U6370 ( .A1(n1575), .A2(n6491), .A3(n6492), .ZN(n7915) );
  INV_X1 U6371 ( .A(Plaintext[59]), .ZN(n1576) );
  INV_X1 U6373 ( .A(n10166), .ZN(n1577) );
  NOR2_X1 U6374 ( .A1(n12555), .A2(n25248), .ZN(n13306) );
  NAND2_X1 U6375 ( .A1(n12914), .A2(n12613), .ZN(n1578) );
  NAND2_X1 U6376 ( .A1(n1579), .A2(n14264), .ZN(n5693) );
  AND2_X2 U6377 ( .A1(n1583), .A2(n1580), .ZN(n21115) );
  NAND2_X1 U6378 ( .A1(n25383), .A2(n2432), .ZN(n1581) );
  NAND2_X1 U6379 ( .A1(n19963), .A2(n20369), .ZN(n1582) );
  AOI21_X1 U6380 ( .B1(n3767), .B2(n24558), .A(n1489), .ZN(n1583) );
  AND2_X1 U6381 ( .A1(n17472), .A2(n17629), .ZN(n1842) );
  NAND2_X1 U6383 ( .A1(n22133), .A2(n1586), .ZN(n1585) );
  NAND2_X1 U6384 ( .A1(n22566), .A2(n22563), .ZN(n1586) );
  NAND2_X1 U6385 ( .A1(n22343), .A2(n22406), .ZN(n1587) );
  NAND4_X1 U6386 ( .A1(n4235), .A2(n1589), .A3(n4233), .A4(n4237), .ZN(n4232)
         );
  NAND2_X1 U6387 ( .A1(n1590), .A2(n20448), .ZN(n20449) );
  NOR2_X1 U6388 ( .A1(n1590), .A2(n20451), .ZN(n20158) );
  NAND2_X1 U6390 ( .A1(n1591), .A2(n20100), .ZN(n17946) );
  AND2_X1 U6391 ( .A1(n1591), .A2(n20103), .ZN(n2358) );
  NOR2_X1 U6392 ( .A1(n1591), .A2(n20101), .ZN(n19915) );
  NAND2_X1 U6393 ( .A1(n21033), .A2(n1591), .ZN(n20105) );
  OAI21_X1 U6394 ( .B1(n21033), .B2(n1591), .A(n20101), .ZN(n19156) );
  OAI21_X1 U6395 ( .B1(n7645), .B2(n5595), .A(n1592), .ZN(n7569) );
  NAND3_X1 U6396 ( .A1(n25151), .A2(n24578), .A3(n7640), .ZN(n1592) );
  NAND2_X1 U6397 ( .A1(n4018), .A2(n6237), .ZN(n1643) );
  INV_X1 U6398 ( .A(n22409), .ZN(n1593) );
  OR2_X1 U6399 ( .A1(n22341), .A2(n24971), .ZN(n22568) );
  AOI22_X2 U6400 ( .A1(n22343), .A2(n22412), .B1(n22342), .B2(n326), .ZN(
        n23166) );
  NOR2_X1 U6401 ( .A1(n9964), .A2(n1595), .ZN(n9965) );
  AOI21_X1 U6403 ( .B1(n9469), .B2(n1595), .A(n9964), .ZN(n8142) );
  MUX2_X1 U6405 ( .A(n9964), .B(n9203), .S(n3292), .Z(n9204) );
  AOI21_X1 U6406 ( .B1(n1597), .B2(n7854), .A(n1596), .ZN(n1598) );
  OR2_X1 U6407 ( .A1(n7722), .A2(n7721), .ZN(n1597) );
  OAI21_X2 U6408 ( .B1(n1598), .B2(n1413), .A(n7724), .ZN(n8478) );
  NOR2_X1 U6409 ( .A1(n20370), .A2(n20369), .ZN(n1600) );
  MUX2_X1 U6412 ( .A(n20368), .B(n20370), .S(n3428), .Z(n1604) );
  AND2_X1 U6414 ( .A1(n22592), .A2(n1605), .ZN(n21189) );
  NAND2_X1 U6415 ( .A1(n25066), .A2(n1605), .ZN(n22450) );
  NOR2_X1 U6416 ( .A1(n25066), .A2(n1605), .ZN(n21923) );
  INV_X1 U6417 ( .A(n7735), .ZN(n7641) );
  NAND2_X1 U6418 ( .A1(n1607), .A2(n7735), .ZN(n7644) );
  NAND2_X1 U6419 ( .A1(n1608), .A2(n7732), .ZN(n1607) );
  NAND2_X1 U6420 ( .A1(n7731), .A2(n7733), .ZN(n1608) );
  INV_X1 U6421 ( .A(n5796), .ZN(n6049) );
  INV_X1 U6422 ( .A(n5796), .ZN(n1609) );
  NAND2_X1 U6423 ( .A1(n1610), .A2(n6728), .ZN(n1642) );
  INV_X1 U6424 ( .A(n16830), .ZN(n1611) );
  NAND2_X1 U6426 ( .A1(n2688), .A2(n1614), .ZN(n2687) );
  NOR2_X1 U6427 ( .A1(n16714), .A2(n17312), .ZN(n1616) );
  NAND2_X1 U6428 ( .A1(n16715), .A2(n17304), .ZN(n1615) );
  INV_X1 U6429 ( .A(n17304), .ZN(n17597) );
  OAI211_X2 U6430 ( .C1(n18815), .C2(n19384), .A(n18814), .B(n1617), .ZN(
        n20491) );
  NAND2_X1 U6431 ( .A1(n19633), .A2(n1617), .ZN(n19636) );
  NAND2_X1 U6432 ( .A1(n18813), .A2(n24909), .ZN(n1617) );
  AND2_X1 U6433 ( .A1(n1619), .A2(n23649), .ZN(n23606) );
  NAND2_X1 U6434 ( .A1(n23638), .A2(n1618), .ZN(n23641) );
  AND3_X1 U6435 ( .A1(n23640), .A2(n23639), .A3(n1619), .ZN(n1618) );
  NAND3_X1 U6436 ( .A1(n23638), .A2(n23640), .A3(n1619), .ZN(n23631) );
  NAND2_X1 U6437 ( .A1(n1622), .A2(n1620), .ZN(n16348) );
  NAND2_X1 U6438 ( .A1(n1621), .A2(n16345), .ZN(n1620) );
  NOR2_X1 U6439 ( .A1(n1654), .A2(n16342), .ZN(n1621) );
  NAND2_X1 U6440 ( .A1(n16346), .A2(n16281), .ZN(n1622) );
  AOI21_X1 U6442 ( .B1(n1624), .B2(n16764), .A(n17274), .ZN(n1623) );
  NAND2_X1 U6443 ( .A1(n17248), .A2(n17273), .ZN(n16764) );
  AOI21_X1 U6445 ( .B1(n16762), .B2(n17252), .A(n1626), .ZN(n1625) );
  INV_X1 U6446 ( .A(n17275), .ZN(n1626) );
  NAND2_X1 U6447 ( .A1(n24300), .A2(n17272), .ZN(n16762) );
  AND2_X1 U6448 ( .A1(n22158), .A2(n2315), .ZN(n22211) );
  OR2_X1 U6449 ( .A1(n2315), .A2(n22158), .ZN(n22065) );
  NAND2_X1 U6450 ( .A1(n1467), .A2(n2315), .ZN(n22161) );
  OAI22_X2 U6451 ( .A1(n21771), .A2(n21770), .B1(n21769), .B2(n1627), .ZN(
        n23596) );
  INV_X1 U6452 ( .A(n2315), .ZN(n1627) );
  AND2_X1 U6453 ( .A1(n18982), .A2(n1629), .ZN(n5566) );
  NAND2_X1 U6454 ( .A1(n19992), .A2(n25378), .ZN(n19993) );
  NAND2_X1 U6456 ( .A1(n1432), .A2(n25378), .ZN(n5563) );
  NAND2_X1 U6457 ( .A1(n13131), .A2(n13151), .ZN(n13153) );
  NAND3_X1 U6458 ( .A1(n13131), .A2(n1774), .A3(n13152), .ZN(n1630) );
  NAND2_X1 U6459 ( .A1(n13133), .A2(n13132), .ZN(n1631) );
  NAND2_X1 U6460 ( .A1(n24376), .A2(n13552), .ZN(n4600) );
  NAND2_X1 U6461 ( .A1(n14268), .A2(n14267), .ZN(n13623) );
  NAND2_X1 U6462 ( .A1(n1636), .A2(n1635), .ZN(n1633) );
  NAND2_X1 U6463 ( .A1(n3371), .A2(n17571), .ZN(n1639) );
  NAND2_X1 U6464 ( .A1(n3374), .A2(n17572), .ZN(n1640) );
  NAND4_X1 U6465 ( .A1(n1641), .A2(n1643), .A3(n7733), .A4(n1642), .ZN(n7567)
         );
  NAND2_X1 U6466 ( .A1(n1645), .A2(n1644), .ZN(n22522) );
  OR2_X1 U6467 ( .A1(n24362), .A2(n21841), .ZN(n1644) );
  NAND2_X1 U6468 ( .A1(n21822), .A2(n21841), .ZN(n1645) );
  XNOR2_X2 U6469 ( .A(n19054), .B(n19053), .ZN(n21841) );
  NAND3_X1 U6470 ( .A1(n21798), .A2(n21796), .A3(n21797), .ZN(n23772) );
  NAND2_X1 U6471 ( .A1(n1646), .A2(n12800), .ZN(n12481) );
  NAND2_X1 U6472 ( .A1(n1646), .A2(n12797), .ZN(n4618) );
  NAND2_X1 U6473 ( .A1(n1648), .A2(n1647), .ZN(n9583) );
  NAND2_X1 U6474 ( .A1(n10136), .A2(n10138), .ZN(n1647) );
  NAND3_X1 U6475 ( .A1(n9367), .A2(n9366), .A3(n1649), .ZN(n9371) );
  MUX2_X1 U6476 ( .A(n5742), .B(n9400), .S(n10138), .Z(n9401) );
  OAI21_X1 U6477 ( .B1(n9201), .B2(n10146), .A(n1649), .ZN(n9202) );
  NAND2_X1 U6478 ( .A1(n17145), .A2(n1653), .ZN(n16848) );
  AOI21_X1 U6480 ( .B1(n16496), .B2(n1653), .A(n16847), .ZN(n16497) );
  NAND2_X1 U6482 ( .A1(n15977), .A2(n15849), .ZN(n1655) );
  NAND2_X1 U6483 ( .A1(n10284), .A2(n1658), .ZN(n3532) );
  NAND2_X1 U6485 ( .A1(n1658), .A2(n11113), .ZN(n11114) );
  INV_X1 U6487 ( .A(n20430), .ZN(n20209) );
  NAND2_X1 U6488 ( .A1(n20400), .A2(n1663), .ZN(n1661) );
  NOR2_X1 U6489 ( .A1(n20415), .A2(n20419), .ZN(n1663) );
  NAND2_X1 U6490 ( .A1(n1666), .A2(n20597), .ZN(n1665) );
  NAND2_X1 U6491 ( .A1(n19846), .A2(n20599), .ZN(n1666) );
  INV_X1 U6492 ( .A(n25477), .ZN(n1667) );
  NAND2_X1 U6493 ( .A1(n9718), .A2(n9635), .ZN(n9436) );
  NAND2_X1 U6494 ( .A1(n1672), .A2(n9634), .ZN(n1671) );
  OAI21_X1 U6495 ( .B1(n9434), .B2(n9710), .A(n9714), .ZN(n1672) );
  NAND3_X1 U6497 ( .A1(n16095), .A2(n15625), .A3(n16147), .ZN(n1676) );
  XNOR2_X2 U6498 ( .A(n14567), .B(n14566), .ZN(n16095) );
  NAND2_X1 U6499 ( .A1(n1677), .A2(n4247), .ZN(n7528) );
  NAND2_X1 U6500 ( .A1(n22113), .A2(n1678), .ZN(n1680) );
  NOR2_X1 U6501 ( .A1(n22072), .A2(n22917), .ZN(n1678) );
  NOR2_X1 U6504 ( .A1(n1681), .A2(n12768), .ZN(n12769) );
  OAI21_X1 U6505 ( .B1(n1681), .B2(n4651), .A(n13218), .ZN(n4547) );
  NAND2_X1 U6506 ( .A1(n13215), .A2(n12767), .ZN(n1681) );
  OR2_X1 U6508 ( .A1(n21887), .A2(n22263), .ZN(n1685) );
  NAND2_X1 U6509 ( .A1(n1685), .A2(n21886), .ZN(n1683) );
  AND2_X1 U6510 ( .A1(n382), .A2(n16067), .ZN(n16065) );
  AOI21_X1 U6511 ( .B1(n380), .B2(n16064), .A(n16060), .ZN(n15796) );
  INV_X1 U6512 ( .A(n11128), .ZN(n1689) );
  NAND3_X1 U6516 ( .A1(n10839), .A2(n11129), .A3(n1689), .ZN(n10716) );
  NAND3_X1 U6517 ( .A1(n10840), .A2(n420), .A3(n1689), .ZN(n10843) );
  NAND2_X1 U6518 ( .A1(n1690), .A2(n7048), .ZN(n6852) );
  OR2_X1 U6519 ( .A1(n21774), .A2(n1691), .ZN(n2513) );
  NAND2_X1 U6520 ( .A1(n327), .A2(n22728), .ZN(n1691) );
  NAND2_X1 U6521 ( .A1(n7034), .A2(n454), .ZN(n1692) );
  NAND2_X1 U6522 ( .A1(n2270), .A2(n7035), .ZN(n1693) );
  MUX2_X1 U6523 ( .A(n1345), .B(n270), .S(n7682), .Z(n7071) );
  INV_X1 U6524 ( .A(n12964), .ZN(n1694) );
  NAND2_X1 U6525 ( .A1(n6740), .A2(n6739), .ZN(n1695) );
  OAI21_X1 U6526 ( .B1(n434), .B2(n7674), .A(n7676), .ZN(n7673) );
  INV_X1 U6527 ( .A(n1696), .ZN(n1697) );
  XNOR2_X2 U6528 ( .A(n5969), .B(Key[179]), .ZN(n1698) );
  NAND2_X1 U6529 ( .A1(n5966), .A2(n1698), .ZN(n6468) );
  NAND2_X1 U6530 ( .A1(n1697), .A2(n5449), .ZN(n5450) );
  NOR2_X1 U6531 ( .A1(n6469), .A2(n1698), .ZN(n7692) );
  XNOR2_X1 U6532 ( .A(n11661), .B(n1699), .ZN(n10707) );
  XNOR2_X1 U6533 ( .A(n11750), .B(n1700), .ZN(n11752) );
  INV_X1 U6534 ( .A(n11661), .ZN(n1700) );
  XNOR2_X1 U6535 ( .A(n25493), .B(n18157), .ZN(n18305) );
  NAND2_X1 U6536 ( .A1(n15834), .A2(n25472), .ZN(n1702) );
  NAND3_X1 U6537 ( .A1(n1704), .A2(n17729), .A3(n17485), .ZN(n1703) );
  NAND3_X1 U6538 ( .A1(n17735), .A2(n24410), .A3(n17093), .ZN(n1705) );
  OAI211_X1 U6539 ( .C1(n19361), .C2(n25392), .A(n1707), .B(n19211), .ZN(n1706) );
  NAND2_X1 U6540 ( .A1(n25392), .A2(n19359), .ZN(n1707) );
  NAND3_X1 U6541 ( .A1(n15779), .A2(n15778), .A3(n15777), .ZN(n17075) );
  INV_X1 U6542 ( .A(n17075), .ZN(n17077) );
  OR2_X1 U6543 ( .A1(n7460), .A2(n268), .ZN(n1904) );
  OAI21_X1 U6547 ( .B1(n19549), .B2(n1710), .A(n19403), .ZN(n2722) );
  INV_X1 U6548 ( .A(n19548), .ZN(n1711) );
  NAND2_X1 U6549 ( .A1(n19552), .A2(n1713), .ZN(n1712) );
  AND2_X1 U6550 ( .A1(n19185), .A2(n25057), .ZN(n1713) );
  NAND2_X1 U6551 ( .A1(n19552), .A2(n19185), .ZN(n1714) );
  NOR2_X1 U6552 ( .A1(n25057), .A2(n1715), .ZN(n19725) );
  NAND2_X1 U6553 ( .A1(n19546), .A2(n19186), .ZN(n1715) );
  NAND2_X1 U6557 ( .A1(n16038), .A2(n2253), .ZN(n1718) );
  NAND2_X1 U6560 ( .A1(n10573), .A2(n11037), .ZN(n10575) );
  NAND2_X1 U6561 ( .A1(n1721), .A2(n1720), .ZN(n18941) );
  NAND2_X1 U6562 ( .A1(n18937), .A2(n19327), .ZN(n1720) );
  NAND2_X1 U6563 ( .A1(n18936), .A2(n19328), .ZN(n1721) );
  NAND2_X2 U6564 ( .A1(n1722), .A2(n21296), .ZN(n23828) );
  XNOR2_X2 U6565 ( .A(n1723), .B(n7436), .ZN(n3472) );
  XNOR2_X1 U6566 ( .A(n7552), .B(n7435), .ZN(n1723) );
  XNOR2_X1 U6567 ( .A(n11517), .B(n11516), .ZN(n11533) );
  OAI21_X1 U6568 ( .B1(n12550), .B2(n13001), .A(n1725), .ZN(n12553) );
  XNOR2_X1 U6571 ( .A(n4386), .B(n8702), .ZN(n9737) );
  NOR2_X1 U6572 ( .A1(n20264), .A2(n20262), .ZN(n19741) );
  INV_X1 U6573 ( .A(n7863), .ZN(n3570) );
  XNOR2_X1 U6574 ( .A(n25436), .B(n14952), .ZN(n14915) );
  NOR2_X1 U6576 ( .A1(n18756), .A2(n5239), .ZN(n5238) );
  OR2_X1 U6577 ( .A1(n21385), .A2(n21918), .ZN(n1727) );
  NAND3_X2 U6578 ( .A1(n5288), .A2(n9373), .A3(n5740), .ZN(n10756) );
  MUX2_X1 U6579 ( .A(n20515), .B(n20514), .S(n20517), .Z(n20275) );
  NAND2_X1 U6580 ( .A1(n19267), .A2(n19266), .ZN(n1729) );
  NAND2_X1 U6581 ( .A1(n19268), .A2(n18917), .ZN(n1730) );
  OAI21_X1 U6582 ( .B1(n24399), .B2(n17559), .A(n1731), .ZN(n18759) );
  NAND2_X1 U6583 ( .A1(n19264), .A2(n19261), .ZN(n1731) );
  OAI21_X1 U6585 ( .B1(n20343), .B2(n24414), .A(n1732), .ZN(n20278) );
  NAND2_X1 U6586 ( .A1(n1733), .A2(n20346), .ZN(n1732) );
  INV_X1 U6587 ( .A(n20277), .ZN(n1733) );
  NAND3_X1 U6588 ( .A1(n6403), .A2(n6401), .A3(n5805), .ZN(n1734) );
  OAI21_X1 U6589 ( .B1(n7563), .B2(n7853), .A(n24072), .ZN(n1737) );
  NAND3_X1 U6590 ( .A1(n24977), .A2(n23416), .A3(n25035), .ZN(n1738) );
  NAND3_X1 U6591 ( .A1(n22563), .A2(n22562), .A3(n22409), .ZN(n20714) );
  NAND3_X2 U6592 ( .A1(n16816), .A2(n16815), .A3(n1394), .ZN(n18149) );
  AOI21_X1 U6593 ( .B1(n16112), .B2(n17170), .A(n17171), .ZN(n16134) );
  NOR2_X2 U6595 ( .A1(n20283), .A2(n2138), .ZN(n20475) );
  NOR2_X1 U6596 ( .A1(n17437), .A2(n1782), .ZN(n1781) );
  NAND2_X1 U6599 ( .A1(n1741), .A2(n7826), .ZN(n6855) );
  OAI21_X1 U6600 ( .B1(n7828), .B2(n7048), .A(n7825), .ZN(n1741) );
  NAND2_X1 U6601 ( .A1(n14508), .A2(n14509), .ZN(n14512) );
  NAND2_X1 U6602 ( .A1(n13693), .A2(n24556), .ZN(n14509) );
  NAND3_X1 U6604 ( .A1(n14124), .A2(n14206), .A3(n14204), .ZN(n3850) );
  NAND2_X1 U6605 ( .A1(n24574), .A2(n10284), .ZN(n9580) );
  NAND2_X1 U6606 ( .A1(n2930), .A2(n2931), .ZN(n5912) );
  NAND3_X1 U6608 ( .A1(n4116), .A2(n14240), .A3(n13200), .ZN(n4117) );
  NAND2_X1 U6609 ( .A1(n7216), .A2(n1743), .ZN(n1742) );
  INV_X1 U6610 ( .A(n2404), .ZN(n1743) );
  NAND2_X1 U6611 ( .A1(n7215), .A2(n2404), .ZN(n1744) );
  NAND2_X1 U6612 ( .A1(n6504), .A2(n6501), .ZN(n6437) );
  AOI22_X1 U6614 ( .A1(n3366), .A2(n7575), .B1(n7573), .B2(n7574), .ZN(n3500)
         );
  NAND2_X1 U6615 ( .A1(n14220), .A2(n14225), .ZN(n1748) );
  AND2_X1 U6616 ( .A1(n4884), .A2(n19237), .ZN(n19610) );
  NAND2_X1 U6617 ( .A1(n5387), .A2(n7913), .ZN(n1749) );
  OAI21_X1 U6618 ( .B1(n9187), .B2(n9397), .A(n10141), .ZN(n1751) );
  XNOR2_X1 U6619 ( .A(n1752), .B(n23063), .ZN(Ciphertext[5]) );
  NAND2_X1 U6620 ( .A1(n1834), .A2(n23061), .ZN(n1752) );
  NAND2_X1 U6621 ( .A1(n1753), .A2(n24043), .ZN(n22594) );
  NAND2_X1 U6622 ( .A1(n5046), .A2(n2393), .ZN(n1753) );
  OR2_X1 U6624 ( .A1(n13211), .A2(n13207), .ZN(n13006) );
  NAND2_X1 U6625 ( .A1(n5651), .A2(n6772), .ZN(n5650) );
  NOR2_X1 U6626 ( .A1(n19910), .A2(n19911), .ZN(n1755) );
  XNOR2_X2 U6627 ( .A(n6035), .B(Key[7]), .ZN(n6351) );
  XNOR2_X1 U6628 ( .A(n17813), .B(n17812), .ZN(n1759) );
  NAND2_X1 U6629 ( .A1(n1761), .A2(n1760), .ZN(n4420) );
  NAND2_X1 U6630 ( .A1(n15864), .A2(n16095), .ZN(n1760) );
  NAND2_X1 U6631 ( .A1(n16151), .A2(n16149), .ZN(n15864) );
  NAND2_X1 U6632 ( .A1(n1415), .A2(n1762), .ZN(n1761) );
  NAND3_X1 U6633 ( .A1(n6752), .A2(n6578), .A3(n6751), .ZN(n6402) );
  OAI21_X1 U6634 ( .B1(n4772), .B2(n4773), .A(n15952), .ZN(n1763) );
  NAND2_X1 U6635 ( .A1(n3413), .A2(n3414), .ZN(n1764) );
  NAND2_X1 U6636 ( .A1(n22939), .A2(n24932), .ZN(n1765) );
  NAND2_X1 U6637 ( .A1(n22027), .A2(n22938), .ZN(n1766) );
  INV_X1 U6639 ( .A(n23869), .ZN(n23889) );
  NAND3_X1 U6641 ( .A1(n3268), .A2(n2522), .A3(n7758), .ZN(n1769) );
  NAND3_X1 U6642 ( .A1(n13157), .A2(n13151), .A3(n25033), .ZN(n13154) );
  OR2_X2 U6644 ( .A1(n13659), .A2(n13660), .ZN(n12669) );
  NAND2_X1 U6645 ( .A1(n1773), .A2(n1772), .ZN(n13659) );
  NAND2_X1 U6646 ( .A1(n12664), .A2(n13148), .ZN(n1772) );
  INV_X1 U6647 ( .A(n13148), .ZN(n1774) );
  XNOR2_X2 U6648 ( .A(n5879), .B(Key[32]), .ZN(n5903) );
  NAND2_X1 U6649 ( .A1(n1941), .A2(n10763), .ZN(n10896) );
  NAND2_X1 U6650 ( .A1(n18739), .A2(n18977), .ZN(n17888) );
  NAND2_X2 U6651 ( .A1(n20106), .A2(n2010), .ZN(n21469) );
  INV_X1 U6652 ( .A(n10713), .ZN(n10840) );
  OAI211_X1 U6653 ( .C1(n13217), .C2(n12986), .A(n4945), .B(n13218), .ZN(
        n12765) );
  NAND2_X1 U6654 ( .A1(n13902), .A2(n4524), .ZN(n13957) );
  NAND2_X1 U6655 ( .A1(n6474), .A2(n6789), .ZN(n6476) );
  XNOR2_X2 U6656 ( .A(n5979), .B(Key[121]), .ZN(n7004) );
  OR2_X1 U6657 ( .A1(n9064), .A2(n10050), .ZN(n3998) );
  XNOR2_X2 U6658 ( .A(n5965), .B(Key[177]), .ZN(n4621) );
  OR2_X1 U6660 ( .A1(n15637), .A2(n16397), .ZN(n2420) );
  NAND2_X1 U6661 ( .A1(n1779), .A2(n1778), .ZN(n7888) );
  NAND2_X1 U6662 ( .A1(n7885), .A2(n7884), .ZN(n1778) );
  NAND2_X1 U6664 ( .A1(n1612), .A2(n1780), .ZN(n17444) );
  NAND2_X1 U6665 ( .A1(n17436), .A2(n1781), .ZN(n1780) );
  NAND3_X1 U6666 ( .A1(n17434), .A2(n17435), .A3(n17433), .ZN(n1782) );
  NAND2_X1 U6669 ( .A1(n1784), .A2(n13067), .ZN(n1783) );
  NAND2_X1 U6670 ( .A1(n12472), .A2(n12471), .ZN(n1784) );
  XNOR2_X2 U6671 ( .A(Key[99]), .B(Plaintext[99]), .ZN(n7029) );
  OAI21_X1 U6673 ( .B1(n1460), .B2(n9697), .A(n1785), .ZN(n9701) );
  NAND2_X1 U6674 ( .A1(n9698), .A2(n9697), .ZN(n1785) );
  NAND2_X1 U6675 ( .A1(n7288), .A2(n1786), .ZN(n7287) );
  INV_X1 U6676 ( .A(n7510), .ZN(n2262) );
  OAI21_X1 U6677 ( .B1(n1788), .B2(n13096), .A(n1787), .ZN(n13100) );
  NAND2_X1 U6678 ( .A1(n13096), .A2(n13095), .ZN(n1787) );
  NAND2_X1 U6679 ( .A1(n13097), .A2(n12871), .ZN(n1788) );
  INV_X1 U6680 ( .A(n8221), .ZN(n7811) );
  MUX2_X1 U6681 ( .A(n8220), .B(n7812), .S(n8221), .Z(n7815) );
  NOR2_X1 U6682 ( .A1(n15706), .A2(n4897), .ZN(n1790) );
  OAI21_X1 U6683 ( .B1(n15824), .B2(n24080), .A(n2336), .ZN(n1791) );
  INV_X1 U6684 ( .A(n9884), .ZN(n5739) );
  INV_X1 U6685 ( .A(n19774), .ZN(n20461) );
  OR2_X1 U6686 ( .A1(n15803), .A2(n17134), .ZN(n15807) );
  NAND2_X1 U6687 ( .A1(n20372), .A2(n19962), .ZN(n1793) );
  XNOR2_X1 U6688 ( .A(n15021), .B(n15020), .ZN(n4957) );
  NAND2_X1 U6689 ( .A1(n19760), .A2(n18385), .ZN(n1982) );
  INV_X1 U6691 ( .A(n16095), .ZN(n16097) );
  INV_X1 U6692 ( .A(n9769), .ZN(n10681) );
  XNOR2_X1 U6693 ( .A(n12167), .B(n12295), .ZN(n11946) );
  XNOR2_X1 U6694 ( .A(n3471), .B(n14598), .ZN(n2000) );
  OR3_X1 U6695 ( .A1(n11169), .A2(n11171), .A3(n8660), .ZN(n3384) );
  NAND2_X1 U6696 ( .A1(n3982), .A2(n16528), .ZN(n16529) );
  NAND2_X1 U6697 ( .A1(n1795), .A2(n1794), .ZN(n10001) );
  NAND2_X1 U6698 ( .A1(n246), .A2(n9998), .ZN(n1794) );
  NAND2_X1 U6699 ( .A1(n25453), .A2(n1796), .ZN(n1795) );
  INV_X1 U6700 ( .A(n9997), .ZN(n1796) );
  AOI21_X1 U6702 ( .B1(n6134), .B2(n6164), .A(n6162), .ZN(n1798) );
  NAND2_X1 U6703 ( .A1(n16219), .A2(n16220), .ZN(n16216) );
  OR2_X1 U6704 ( .A1(n9832), .A2(n9829), .ZN(n9827) );
  NAND2_X1 U6705 ( .A1(n6156), .A2(n6523), .ZN(n6278) );
  NAND2_X1 U6707 ( .A1(n9564), .A2(n9565), .ZN(n9884) );
  XNOR2_X1 U6709 ( .A(n4670), .B(n3512), .ZN(n11690) );
  NAND2_X1 U6710 ( .A1(n350), .A2(n3657), .ZN(n20462) );
  NAND3_X1 U6712 ( .A1(n2326), .A2(n22893), .A3(n22835), .ZN(n1802) );
  NAND2_X1 U6713 ( .A1(n5766), .A2(n25438), .ZN(n1803) );
  INV_X1 U6714 ( .A(n6997), .ZN(n3109) );
  OAI211_X1 U6716 ( .C1(n19239), .C2(n278), .A(n3919), .B(n1805), .ZN(n3918)
         );
  INV_X1 U6718 ( .A(n20218), .ZN(n1809) );
  OAI21_X1 U6719 ( .B1(n4684), .B2(n17130), .A(n1811), .ZN(n16789) );
  NAND2_X1 U6720 ( .A1(n4684), .A2(n25227), .ZN(n1811) );
  XNOR2_X2 U6721 ( .A(n5871), .B(Key[42]), .ZN(n5924) );
  NAND2_X1 U6722 ( .A1(n2892), .A2(n5105), .ZN(n10934) );
  AND2_X1 U6723 ( .A1(n7604), .A2(n7323), .ZN(n2552) );
  NAND2_X1 U6724 ( .A1(n13216), .A2(n13217), .ZN(n12539) );
  AND2_X2 U6725 ( .A1(n5297), .A2(n5298), .ZN(n15446) );
  INV_X1 U6726 ( .A(n16171), .ZN(n15820) );
  NAND2_X1 U6727 ( .A1(n6487), .A2(n6301), .ZN(n6302) );
  NAND2_X1 U6729 ( .A1(n3064), .A2(n3066), .ZN(n12529) );
  AND3_X2 U6730 ( .A1(n14887), .A2(n14888), .A3(n15925), .ZN(n17608) );
  OAI21_X1 U6731 ( .B1(n348), .B2(n4065), .A(n20476), .ZN(n5244) );
  NOR2_X1 U6732 ( .A1(n16539), .A2(n2247), .ZN(n2246) );
  XNOR2_X2 U6733 ( .A(n11318), .B(n11317), .ZN(n12993) );
  NAND2_X1 U6734 ( .A1(n25246), .A2(n17413), .ZN(n17418) );
  NAND2_X1 U6735 ( .A1(n7792), .A2(n7793), .ZN(n8366) );
  NAND2_X1 U6736 ( .A1(n2160), .A2(n6326), .ZN(n6327) );
  NAND2_X1 U6738 ( .A1(n9753), .A2(n9613), .ZN(n1814) );
  NAND2_X1 U6739 ( .A1(n10855), .A2(n25230), .ZN(n10282) );
  NAND2_X1 U6740 ( .A1(n5065), .A2(n5066), .ZN(n1816) );
  NAND2_X1 U6741 ( .A1(n16310), .A2(n1817), .ZN(n16313) );
  AND3_X1 U6742 ( .A1(n250), .A2(n6848), .A3(n7025), .ZN(n2738) );
  OR2_X1 U6743 ( .A1(n15846), .A2(n16154), .ZN(n2992) );
  NAND2_X1 U6744 ( .A1(n1818), .A2(n2544), .ZN(n2543) );
  XNOR2_X1 U6745 ( .A(n3931), .B(n5513), .ZN(n16440) );
  INV_X1 U6746 ( .A(n17130), .ZN(n3458) );
  NAND2_X1 U6747 ( .A1(n13891), .A2(n1819), .ZN(n15523) );
  NAND2_X1 U6748 ( .A1(n1820), .A2(n13728), .ZN(n1819) );
  NAND2_X1 U6749 ( .A1(n13889), .A2(n13944), .ZN(n1820) );
  OR2_X1 U6751 ( .A1(n15929), .A2(n15725), .ZN(n15730) );
  INV_X1 U6752 ( .A(n13394), .ZN(n2629) );
  OR2_X1 U6753 ( .A1(n6556), .A2(n6414), .ZN(n6935) );
  INV_X1 U6754 ( .A(n13807), .ZN(n14035) );
  INV_X1 U6755 ( .A(n9681), .ZN(n4069) );
  INV_X1 U6756 ( .A(n15583), .ZN(n5100) );
  XNOR2_X1 U6757 ( .A(n2077), .B(n11906), .ZN(n5749) );
  INV_X1 U6758 ( .A(n24542), .ZN(n17598) );
  XNOR2_X1 U6759 ( .A(n3233), .B(n15191), .ZN(n15155) );
  XNOR2_X1 U6761 ( .A(n12214), .B(n11990), .ZN(n1821) );
  NAND3_X2 U6762 ( .A1(n5527), .A2(n5525), .A3(n13588), .ZN(n15230) );
  NAND2_X1 U6763 ( .A1(n1823), .A2(n1436), .ZN(n1822) );
  INV_X1 U6764 ( .A(n18901), .ZN(n1823) );
  NAND2_X1 U6765 ( .A1(n11201), .A2(n10630), .ZN(n1824) );
  NAND3_X1 U6766 ( .A1(n6949), .A2(n6255), .A3(n5903), .ZN(n5528) );
  NAND2_X1 U6767 ( .A1(n1825), .A2(n377), .ZN(n5546) );
  NOR2_X1 U6768 ( .A1(n15695), .A2(n25238), .ZN(n1825) );
  NAND2_X1 U6769 ( .A1(n1441), .A2(n6731), .ZN(n1922) );
  NAND2_X1 U6770 ( .A1(n6734), .A2(n6238), .ZN(n6731) );
  NAND2_X1 U6772 ( .A1(n20909), .A2(n20491), .ZN(n20483) );
  NAND3_X1 U6773 ( .A1(n16262), .A2(n16261), .A3(n25219), .ZN(n16263) );
  NAND2_X1 U6774 ( .A1(n353), .A2(n19125), .ZN(n5571) );
  XOR2_X1 U6775 ( .A(n18281), .B(n18280), .Z(n3753) );
  INV_X1 U6776 ( .A(n13302), .ZN(n1828) );
  NAND2_X1 U6777 ( .A1(n9664), .A2(n9985), .ZN(n9742) );
  NAND2_X1 U6778 ( .A1(n2668), .A2(n2669), .ZN(n2238) );
  NAND3_X2 U6779 ( .A1(n4889), .A2(n1402), .A3(n1372), .ZN(n8787) );
  OAI21_X1 U6780 ( .B1(n25223), .B2(n25347), .A(n1996), .ZN(n19816) );
  AOI22_X1 U6781 ( .A1(n1830), .A2(n6468), .B1(n5451), .B2(n6467), .ZN(n7690)
         );
  NAND2_X1 U6782 ( .A1(n25404), .A2(n6425), .ZN(n1830) );
  OR2_X1 U6783 ( .A1(n23062), .A2(n322), .ZN(n1834) );
  INV_X1 U6784 ( .A(n10100), .ZN(n9836) );
  OAI21_X1 U6785 ( .B1(n17003), .B2(n17051), .A(n3643), .ZN(n3646) );
  XNOR2_X1 U6789 ( .A(n10601), .B(n3565), .ZN(n10602) );
  INV_X1 U6790 ( .A(n5971), .ZN(n1839) );
  NAND2_X1 U6791 ( .A1(n1842), .A2(n17473), .ZN(n1841) );
  INV_X1 U6792 ( .A(n4503), .ZN(n5884) );
  NAND2_X1 U6793 ( .A1(n1844), .A2(n1843), .ZN(n12501) );
  NAND2_X1 U6794 ( .A1(n25033), .A2(n13130), .ZN(n1843) );
  OAI21_X1 U6795 ( .B1(n10254), .B2(n5057), .A(n9379), .ZN(n5289) );
  OAI211_X1 U6796 ( .C1(n15972), .C2(n15971), .A(n3630), .B(n1845), .ZN(n3629)
         );
  NAND2_X1 U6797 ( .A1(n15971), .A2(n1846), .ZN(n1845) );
  INV_X1 U6798 ( .A(n15638), .ZN(n1846) );
  NAND2_X1 U6799 ( .A1(n1847), .A2(n1275), .ZN(n4255) );
  NAND2_X1 U6800 ( .A1(n10110), .A2(n10107), .ZN(n1847) );
  INV_X1 U6801 ( .A(n9121), .ZN(n7895) );
  NAND2_X1 U6802 ( .A1(n7888), .A2(n7887), .ZN(n9121) );
  NAND2_X1 U6803 ( .A1(n4676), .A2(n4675), .ZN(n3555) );
  NAND2_X1 U6804 ( .A1(n1850), .A2(n1849), .ZN(n4676) );
  NAND2_X1 U6805 ( .A1(n2479), .A2(n25030), .ZN(n1849) );
  NAND2_X1 U6806 ( .A1(n2480), .A2(n24586), .ZN(n1850) );
  NAND2_X1 U6807 ( .A1(n6455), .A2(n25428), .ZN(n6507) );
  NAND3_X1 U6808 ( .A1(n17024), .A2(n2230), .A3(n1852), .ZN(n17026) );
  NAND2_X1 U6811 ( .A1(n17015), .A2(n17208), .ZN(n16557) );
  NAND2_X1 U6812 ( .A1(n19888), .A2(n20316), .ZN(n3541) );
  NAND2_X1 U6813 ( .A1(n2251), .A2(n15263), .ZN(n15264) );
  INV_X1 U6814 ( .A(n15319), .ZN(n15126) );
  INV_X1 U6815 ( .A(n13583), .ZN(n14105) );
  NAND2_X1 U6816 ( .A1(n9993), .A2(n24534), .ZN(n1857) );
  NAND2_X1 U6817 ( .A1(n9994), .A2(n422), .ZN(n1858) );
  NAND2_X1 U6820 ( .A1(n12637), .A2(n398), .ZN(n1859) );
  NAND2_X1 U6821 ( .A1(n12638), .A2(n1861), .ZN(n1860) );
  INV_X1 U6822 ( .A(n398), .ZN(n1861) );
  XNOR2_X1 U6824 ( .A(n24472), .B(n1381), .ZN(n20839) );
  NAND2_X1 U6827 ( .A1(n3324), .A2(n10757), .ZN(n9364) );
  NAND2_X1 U6828 ( .A1(n14008), .A2(n14252), .ZN(n13701) );
  NAND2_X1 U6829 ( .A1(n15925), .A2(n3778), .ZN(n1872) );
  NAND2_X1 U6830 ( .A1(n3380), .A2(n15904), .ZN(n14138) );
  OAI21_X1 U6831 ( .B1(n5246), .B2(n14042), .A(n298), .ZN(n2155) );
  NAND2_X1 U6832 ( .A1(n6755), .A2(n6673), .ZN(n6579) );
  OR3_X1 U6833 ( .A1(n7350), .A2(n7349), .A3(n7346), .ZN(n7352) );
  NAND3_X1 U6834 ( .A1(n19530), .A2(n19270), .A3(n24329), .ZN(n5654) );
  OAI22_X1 U6835 ( .A1(n13773), .A2(n14179), .B1(n13774), .B2(n24949), .ZN(
        n1866) );
  NOR2_X1 U6836 ( .A1(n14088), .A2(n14092), .ZN(n1868) );
  NAND2_X1 U6838 ( .A1(n12845), .A2(n1456), .ZN(n12846) );
  NAND2_X1 U6839 ( .A1(n12947), .A2(n12945), .ZN(n12845) );
  OAI211_X1 U6840 ( .C1(n16724), .C2(n2666), .A(n2665), .B(n2664), .ZN(n17676)
         );
  NAND3_X1 U6841 ( .A1(n312), .A2(n7636), .A3(n435), .ZN(n6495) );
  XNOR2_X1 U6842 ( .A(n15150), .B(n14414), .ZN(n3308) );
  XNOR2_X1 U6843 ( .A(n15159), .B(n15161), .ZN(n3670) );
  OAI21_X1 U6844 ( .B1(n15314), .B2(n17240), .A(n17346), .ZN(n15473) );
  NAND2_X1 U6845 ( .A1(n7580), .A2(n7573), .ZN(n3548) );
  INV_X1 U6847 ( .A(n16029), .ZN(n16273) );
  NOR2_X1 U6848 ( .A1(n6818), .A2(n6895), .ZN(n3414) );
  NAND2_X1 U6849 ( .A1(n2290), .A2(n12794), .ZN(n2048) );
  NAND2_X1 U6850 ( .A1(n12991), .A2(n4587), .ZN(n12794) );
  NAND2_X1 U6851 ( .A1(n1872), .A2(n16459), .ZN(n15704) );
  OR3_X1 U6853 ( .A1(n14130), .A2(n14127), .A3(n14126), .ZN(n13407) );
  NAND2_X1 U6854 ( .A1(n22771), .A2(n22774), .ZN(n22773) );
  NAND2_X1 U6855 ( .A1(n5498), .A2(n14256), .ZN(n14259) );
  XNOR2_X1 U6856 ( .A(n4590), .B(n12196), .ZN(n12095) );
  OR2_X1 U6857 ( .A1(n1971), .A2(n4861), .ZN(n4860) );
  NAND2_X1 U6858 ( .A1(n3616), .A2(n7747), .ZN(n1873) );
  INV_X1 U6859 ( .A(n11806), .ZN(n13963) );
  OAI21_X1 U6861 ( .B1(n271), .B2(n6752), .A(n2494), .ZN(n2496) );
  AOI21_X1 U6862 ( .B1(n16851), .B2(n16850), .A(n2105), .ZN(n16853) );
  INV_X1 U6863 ( .A(n5255), .ZN(n8671) );
  INV_X1 U6864 ( .A(n12636), .ZN(n13348) );
  INV_X1 U6865 ( .A(n10613), .ZN(n10412) );
  INV_X1 U6866 ( .A(n13305), .ZN(n12917) );
  INV_X1 U6867 ( .A(n10596), .ZN(n10936) );
  INV_X1 U6868 ( .A(n11070), .ZN(n11068) );
  INV_X1 U6869 ( .A(n13906), .ZN(n15410) );
  INV_X1 U6870 ( .A(n13868), .ZN(n14458) );
  OAI21_X1 U6871 ( .B1(n7313), .B2(n7582), .A(n7314), .ZN(n7470) );
  INV_X1 U6872 ( .A(n8667), .ZN(n8039) );
  INV_X1 U6873 ( .A(n12003), .ZN(n2917) );
  INV_X1 U6874 ( .A(n8203), .ZN(n9052) );
  INV_X1 U6875 ( .A(n223), .ZN(n15726) );
  INV_X1 U6876 ( .A(n24012), .ZN(n4477) );
  XNOR2_X1 U6877 ( .A(n14486), .B(n14485), .ZN(n15612) );
  OAI211_X1 U6878 ( .C1(n15573), .C2(n15572), .A(n2651), .B(n16274), .ZN(n2648) );
  XNOR2_X1 U6879 ( .A(n15153), .B(n1920), .ZN(n14841) );
  NAND2_X1 U6880 ( .A1(n7015), .A2(n1876), .ZN(n6828) );
  NAND2_X1 U6885 ( .A1(n7564), .A2(n6413), .ZN(n1880) );
  NAND2_X1 U6886 ( .A1(n6925), .A2(n6480), .ZN(n6923) );
  NAND2_X1 U6887 ( .A1(n20559), .A2(n20092), .ZN(n1881) );
  NAND2_X1 U6888 ( .A1(n405), .A2(n13235), .ZN(n5359) );
  NAND2_X1 U6889 ( .A1(n4617), .A2(n16461), .ZN(n14887) );
  AND3_X2 U6890 ( .A1(n12572), .A2(n12571), .A3(n12570), .ZN(n14075) );
  NAND2_X1 U6891 ( .A1(n1883), .A2(n1882), .ZN(n16669) );
  OR3_X1 U6892 ( .A1(n17347), .A2(n17241), .A3(n17342), .ZN(n1882) );
  XNOR2_X1 U6894 ( .A(n14403), .B(n14891), .ZN(n1884) );
  NAND2_X1 U6896 ( .A1(n1885), .A2(n5361), .ZN(n5360) );
  NAND2_X1 U6897 ( .A1(n407), .A2(n13264), .ZN(n1885) );
  AOI21_X1 U6898 ( .B1(n9329), .B2(n9503), .A(n1886), .ZN(n9333) );
  NAND2_X1 U6899 ( .A1(n2011), .A2(n9736), .ZN(n9430) );
  OAI21_X1 U6902 ( .B1(n10536), .B2(n4998), .A(n10535), .ZN(n1887) );
  AOI22_X1 U6905 ( .A1(n9845), .A2(n10151), .B1(n10152), .B2(n9843), .ZN(
        n10154) );
  OAI21_X1 U6906 ( .B1(n10669), .B2(n24340), .A(n1910), .ZN(n11218) );
  MUX2_X1 U6908 ( .A(n6878), .B(n6877), .S(n6876), .Z(n1888) );
  NAND3_X1 U6910 ( .A1(n385), .A2(n16448), .A3(n223), .ZN(n15728) );
  OAI21_X1 U6911 ( .B1(n7943), .B2(n4259), .A(n1892), .ZN(n7229) );
  NAND2_X1 U6912 ( .A1(n7943), .A2(n7942), .ZN(n1892) );
  NAND2_X1 U6913 ( .A1(n13460), .A2(n14307), .ZN(n13902) );
  INV_X1 U6917 ( .A(n15861), .ZN(n16116) );
  OR2_X1 U6918 ( .A1(n10303), .A2(n10302), .ZN(n5678) );
  NAND2_X1 U6919 ( .A1(n16535), .A2(n4774), .ZN(n16536) );
  XNOR2_X2 U6920 ( .A(n21628), .B(n21629), .ZN(n22832) );
  NAND2_X1 U6921 ( .A1(n13171), .A2(n11597), .ZN(n1893) );
  NAND2_X1 U6922 ( .A1(n11596), .A2(n13165), .ZN(n1894) );
  NAND3_X1 U6923 ( .A1(n7617), .A2(n7384), .A3(n1895), .ZN(n7202) );
  XNOR2_X1 U6924 ( .A(n8190), .B(n8189), .ZN(n9842) );
  NOR2_X1 U6926 ( .A1(n3817), .A2(n16974), .ZN(n3815) );
  OAI21_X1 U6927 ( .B1(n3578), .B2(n15790), .A(n1897), .ZN(n3576) );
  NAND2_X1 U6932 ( .A1(n1902), .A2(n1901), .ZN(n7603) );
  NAND2_X1 U6933 ( .A1(n7600), .A2(n7595), .ZN(n1901) );
  INV_X1 U6934 ( .A(n12541), .ZN(n4651) );
  XNOR2_X1 U6935 ( .A(n8558), .B(n3048), .ZN(n1903) );
  NAND2_X1 U6936 ( .A1(n22831), .A2(n337), .ZN(n1905) );
  XNOR2_X2 U6937 ( .A(n5937), .B(Key[1]), .ZN(n6456) );
  NAND2_X1 U6938 ( .A1(n9306), .A2(n9788), .ZN(n8455) );
  INV_X1 U6939 ( .A(n16048), .ZN(n15606) );
  NAND2_X1 U6940 ( .A1(n294), .A2(n16048), .ZN(n4624) );
  AND2_X1 U6941 ( .A1(n7749), .A2(n8012), .ZN(n7535) );
  NAND2_X1 U6944 ( .A1(n24570), .A2(n372), .ZN(n1909) );
  NAND2_X1 U6945 ( .A1(n24340), .A2(n11216), .ZN(n1910) );
  NAND2_X1 U6946 ( .A1(n16389), .A2(n1912), .ZN(n1911) );
  NOR2_X1 U6947 ( .A1(n15977), .A2(n16394), .ZN(n1912) );
  NAND2_X1 U6948 ( .A1(n14546), .A2(n15977), .ZN(n1913) );
  OAI21_X1 U6949 ( .B1(n17069), .B2(n369), .A(n1914), .ZN(n15610) );
  NAND2_X1 U6950 ( .A1(n17065), .A2(n16731), .ZN(n1914) );
  NAND2_X1 U6952 ( .A1(n1916), .A2(n1915), .ZN(n12733) );
  NAND2_X1 U6953 ( .A1(n11109), .A2(n13144), .ZN(n1916) );
  OR2_X1 U6954 ( .A1(n11210), .A2(n11209), .ZN(n1918) );
  NOR2_X1 U6956 ( .A1(n19791), .A2(n174), .ZN(n5338) );
  NOR2_X1 U6957 ( .A1(n9760), .A2(n9764), .ZN(n10076) );
  AOI22_X2 U6958 ( .A1(n10609), .A2(n10966), .B1(n10608), .B2(n1919), .ZN(
        n12031) );
  AOI21_X1 U6959 ( .B1(n10607), .B2(n10970), .A(n10606), .ZN(n1919) );
  OR2_X1 U6961 ( .A1(n10444), .A2(n10751), .ZN(n10447) );
  NAND2_X1 U6962 ( .A1(n260), .A2(n10044), .ZN(n10047) );
  OR2_X1 U6963 ( .A1(n2576), .A2(n6658), .ZN(n3110) );
  NAND2_X1 U6964 ( .A1(n24998), .A2(n23689), .ZN(n23688) );
  INV_X1 U6965 ( .A(n16962), .ZN(n17441) );
  NOR2_X1 U6966 ( .A1(n23464), .A2(n23014), .ZN(n22863) );
  OAI21_X1 U6967 ( .B1(n3422), .B2(n13051), .A(n3420), .ZN(n13386) );
  INV_X1 U6968 ( .A(n8928), .ZN(n8557) );
  INV_X1 U6969 ( .A(n17321), .ZN(n15673) );
  XNOR2_X1 U6970 ( .A(n15175), .B(n15003), .ZN(n5210) );
  NAND2_X1 U6971 ( .A1(n12526), .A2(n12796), .ZN(n3066) );
  OR2_X1 U6972 ( .A1(n10907), .A2(n10901), .ZN(n4342) );
  INV_X1 U6973 ( .A(n17386), .ZN(n17179) );
  OR2_X1 U6974 ( .A1(n11067), .A2(n11062), .ZN(n10059) );
  INV_X1 U6975 ( .A(n10128), .ZN(n10254) );
  INV_X1 U6976 ( .A(n4422), .ZN(n5559) );
  INV_X1 U6977 ( .A(n13279), .ZN(n13283) );
  INV_X1 U6978 ( .A(n8157), .ZN(n9567) );
  INV_X1 U6979 ( .A(n8119), .ZN(n9190) );
  INV_X1 U6980 ( .A(n17410), .ZN(n4487) );
  INV_X1 U6981 ( .A(n23326), .ZN(n3564) );
  NOR2_X1 U6982 ( .A1(n3544), .A2(n16202), .ZN(n3543) );
  INV_X1 U6983 ( .A(n2674), .ZN(n22420) );
  INV_X1 U6984 ( .A(n9140), .ZN(n5346) );
  AOI21_X1 U6985 ( .B1(n22948), .B2(n22947), .A(n2673), .ZN(n22949) );
  NOR2_X1 U6986 ( .A1(n17616), .A2(n17609), .ZN(n17610) );
  XNOR2_X1 U6987 ( .A(n13710), .B(n13709), .ZN(n3779) );
  XNOR2_X1 U6988 ( .A(n8615), .B(n8616), .ZN(n9090) );
  XNOR2_X1 U6989 ( .A(Plaintext[185]), .B(Key[185]), .ZN(n4866) );
  OAI22_X1 U6990 ( .A1(n24492), .A2(n23350), .B1(n23354), .B2(n23359), .ZN(
        n23363) );
  XNOR2_X1 U6991 ( .A(n12219), .B(n11542), .ZN(n11787) );
  OAI21_X2 U6992 ( .B1(n2008), .B2(n5900), .A(n5899), .ZN(n7897) );
  NAND2_X1 U6993 ( .A1(n2459), .A2(n7911), .ZN(n2458) );
  OAI22_X1 U6994 ( .A1(n25432), .A2(n16349), .B1(n16595), .B2(n24467), .ZN(
        n15671) );
  NAND2_X1 U6995 ( .A1(n16225), .A2(n15774), .ZN(n16024) );
  NAND3_X1 U6996 ( .A1(n2306), .A2(n24420), .A3(n10369), .ZN(n1921) );
  NAND2_X1 U6997 ( .A1(n2461), .A2(n7628), .ZN(n2460) );
  NAND2_X1 U6998 ( .A1(n6617), .A2(n1922), .ZN(n7787) );
  INV_X1 U6999 ( .A(n17463), .ZN(n5052) );
  NAND3_X1 U7000 ( .A1(n2721), .A2(n12635), .A3(n1923), .ZN(n14200) );
  NAND3_X1 U7001 ( .A1(n12633), .A2(n4529), .A3(n12632), .ZN(n1923) );
  NAND3_X1 U7003 ( .A1(n1459), .A2(n25445), .A3(n13417), .ZN(n13553) );
  OAI21_X2 U7004 ( .B1(n7639), .B2(n7638), .A(n1928), .ZN(n8760) );
  NAND2_X1 U7005 ( .A1(n7637), .A2(n7915), .ZN(n1928) );
  XNOR2_X1 U7006 ( .A(n1929), .B(n11991), .ZN(n10672) );
  XNOR2_X1 U7007 ( .A(n10647), .B(n10646), .ZN(n1929) );
  NAND2_X1 U7008 ( .A1(n24082), .A2(n11338), .ZN(n2675) );
  XNOR2_X1 U7010 ( .A(n1931), .B(n23401), .ZN(Ciphertext[84]) );
  NAND3_X1 U7011 ( .A1(n2630), .A2(n23400), .A3(n23399), .ZN(n1931) );
  AOI22_X1 U7013 ( .A1(n1933), .A2(n1932), .B1(n13584), .B2(n1932), .ZN(n5708)
         );
  INV_X1 U7014 ( .A(n4868), .ZN(n1932) );
  OR2_X1 U7015 ( .A1(n7358), .A2(n7412), .ZN(n7360) );
  INV_X1 U7016 ( .A(n25201), .ZN(n17211) );
  NAND2_X1 U7017 ( .A1(n4491), .A2(n4492), .ZN(n14126) );
  OAI21_X1 U7018 ( .B1(n21362), .B2(n21363), .A(n1934), .ZN(n21364) );
  INV_X1 U7019 ( .A(n16691), .ZN(n16496) );
  NOR2_X1 U7020 ( .A1(n19659), .A2(n3241), .ZN(n1936) );
  XNOR2_X1 U7021 ( .A(n17829), .B(n17830), .ZN(n19459) );
  OAI21_X1 U7023 ( .B1(n16965), .B2(n17127), .A(n17445), .ZN(n17661) );
  NAND2_X1 U7025 ( .A1(n1938), .A2(n24599), .ZN(n2398) );
  NAND2_X1 U7026 ( .A1(n25064), .A2(n10168), .ZN(n1938) );
  NAND2_X1 U7027 ( .A1(n9710), .A2(n1939), .ZN(n8886) );
  INV_X1 U7028 ( .A(n18432), .ZN(n17862) );
  OAI21_X2 U7029 ( .B1(n2653), .B2(n16744), .A(n2652), .ZN(n18432) );
  OAI211_X1 U7030 ( .C1(n10384), .C2(n11524), .A(n1940), .B(n11529), .ZN(n2124) );
  NAND2_X1 U7031 ( .A1(n11089), .A2(n11298), .ZN(n1941) );
  XNOR2_X1 U7032 ( .A(n15251), .B(n3787), .ZN(n4399) );
  INV_X1 U7033 ( .A(n13264), .ZN(n12932) );
  NAND3_X1 U7034 ( .A1(n2506), .A2(n2504), .A3(n5151), .ZN(n2503) );
  NAND3_X1 U7036 ( .A1(n14171), .A2(n14165), .A3(n14164), .ZN(n13734) );
  NAND2_X1 U7039 ( .A1(n3266), .A2(n7841), .ZN(n3265) );
  NAND3_X1 U7040 ( .A1(n3058), .A2(n1945), .A3(n1944), .ZN(n12276) );
  NAND2_X1 U7041 ( .A1(n10572), .A2(n11038), .ZN(n1944) );
  NAND2_X1 U7042 ( .A1(n10513), .A2(n10571), .ZN(n1945) );
  OR2_X1 U7044 ( .A1(n13048), .A2(n12490), .ZN(n2792) );
  NAND2_X1 U7045 ( .A1(n15687), .A2(n257), .ZN(n1946) );
  NAND2_X1 U7046 ( .A1(n1948), .A2(n16235), .ZN(n1947) );
  OAI21_X1 U7047 ( .B1(n15726), .B2(n16447), .A(n16239), .ZN(n1948) );
  INV_X1 U7048 ( .A(n14389), .ZN(n15504) );
  NAND2_X1 U7049 ( .A1(n1950), .A2(n1949), .ZN(n19801) );
  NAND2_X1 U7050 ( .A1(n19799), .A2(n20517), .ZN(n1949) );
  NAND2_X1 U7051 ( .A1(n19797), .A2(n3522), .ZN(n1950) );
  OAI211_X1 U7053 ( .C1(n22628), .C2(n21895), .A(n21897), .B(n21896), .ZN(
        n21899) );
  XOR2_X1 U7054 ( .A(n8867), .B(n8446), .Z(n3507) );
  AOI22_X2 U7055 ( .A1(n9026), .A2(n9564), .B1(n9025), .B2(n9565), .ZN(n10942)
         );
  INV_X1 U7056 ( .A(n22462), .ZN(n3938) );
  NAND2_X1 U7057 ( .A1(n1955), .A2(n1953), .ZN(n20139) );
  NAND2_X1 U7058 ( .A1(n1954), .A2(n20134), .ZN(n1953) );
  NAND2_X1 U7059 ( .A1(n4728), .A2(n20136), .ZN(n1955) );
  NOR2_X2 U7060 ( .A1(n10344), .A2(n10345), .ZN(n11951) );
  NAND3_X1 U7061 ( .A1(n1957), .A2(n1472), .A3(n1956), .ZN(n16971) );
  NAND2_X1 U7062 ( .A1(n15932), .A2(n16494), .ZN(n1956) );
  NAND2_X1 U7063 ( .A1(n15566), .A2(n16231), .ZN(n1957) );
  NAND2_X1 U7064 ( .A1(n6595), .A2(n6594), .ZN(n7782) );
  NAND3_X1 U7065 ( .A1(n21889), .A2(n5665), .A3(n22966), .ZN(n5664) );
  XNOR2_X1 U7066 ( .A(n5200), .B(n15033), .ZN(n4723) );
  NAND2_X1 U7068 ( .A1(n1959), .A2(n5893), .ZN(n1958) );
  NAND2_X1 U7069 ( .A1(n2007), .A2(n2006), .ZN(n1960) );
  NAND3_X1 U7070 ( .A1(n7350), .A2(n8508), .A3(n7347), .ZN(n6219) );
  NAND2_X1 U7071 ( .A1(n6695), .A2(n6699), .ZN(n1962) );
  OAI22_X1 U7072 ( .A1(n5616), .A2(n9897), .B1(n227), .B2(n9945), .ZN(n1963)
         );
  NAND3_X1 U7073 ( .A1(n3186), .A2(n3187), .A3(n16005), .ZN(n1965) );
  NAND2_X1 U7074 ( .A1(n17463), .A2(n16846), .ZN(n4198) );
  OR2_X1 U7075 ( .A1(n16007), .A2(n16266), .ZN(n1964) );
  NAND2_X1 U7077 ( .A1(n14231), .A2(n14230), .ZN(n13994) );
  NAND2_X1 U7078 ( .A1(n13680), .A2(n24402), .ZN(n1968) );
  NAND3_X1 U7079 ( .A1(n14231), .A2(n24402), .A3(n13682), .ZN(n1967) );
  NOR2_X2 U7080 ( .A1(n13683), .A2(n13681), .ZN(n14231) );
  NAND2_X1 U7081 ( .A1(n14232), .A2(n25434), .ZN(n1969) );
  NOR2_X1 U7083 ( .A1(n7531), .A2(n1975), .ZN(n3616) );
  NAND2_X1 U7084 ( .A1(n7277), .A2(n1975), .ZN(n8351) );
  AOI21_X1 U7085 ( .B1(n3611), .B2(n1975), .A(n2196), .ZN(n3613) );
  NAND2_X1 U7086 ( .A1(n7747), .A2(n5738), .ZN(n1973) );
  NAND2_X1 U7087 ( .A1(n3588), .A2(n1975), .ZN(n1974) );
  OAI21_X1 U7088 ( .B1(n6672), .B2(n4754), .A(n1976), .ZN(n6670) );
  NAND2_X1 U7089 ( .A1(n6669), .A2(n4754), .ZN(n1976) );
  OAI21_X1 U7092 ( .B1(n18901), .B2(n18442), .A(n1979), .ZN(n1978) );
  NAND2_X1 U7093 ( .A1(n18428), .A2(n25489), .ZN(n18901) );
  NAND2_X1 U7094 ( .A1(n1981), .A2(n19179), .ZN(n1980) );
  NAND2_X1 U7095 ( .A1(n1982), .A2(n19003), .ZN(n1981) );
  NAND2_X1 U7096 ( .A1(n18777), .A2(n19428), .ZN(n19003) );
  NAND2_X1 U7097 ( .A1(n16465), .A2(n16221), .ZN(n3778) );
  INV_X1 U7098 ( .A(n15922), .ZN(n1983) );
  NAND2_X1 U7099 ( .A1(n1985), .A2(n7682), .ZN(n7685) );
  NAND2_X1 U7100 ( .A1(n1345), .A2(n7683), .ZN(n7966) );
  NAND2_X1 U7101 ( .A1(n270), .A2(n1985), .ZN(n5684) );
  OAI21_X1 U7102 ( .B1(n270), .B2(n1985), .A(n7234), .ZN(n7036) );
  NAND2_X1 U7104 ( .A1(n1988), .A2(n19171), .ZN(n1987) );
  NAND2_X1 U7105 ( .A1(n25469), .A2(n19412), .ZN(n1990) );
  NAND2_X1 U7107 ( .A1(n19627), .A2(n20479), .ZN(n1991) );
  NAND2_X1 U7108 ( .A1(n19628), .A2(n2168), .ZN(n1993) );
  NAND2_X1 U7111 ( .A1(n25347), .A2(n20507), .ZN(n1996) );
  OAI21_X1 U7112 ( .B1(n23320), .B2(n23311), .A(n23313), .ZN(n2920) );
  NAND2_X1 U7113 ( .A1(n6274), .A2(n1509), .ZN(n6028) );
  NAND2_X1 U7116 ( .A1(n13724), .A2(n13965), .ZN(n13725) );
  NAND2_X1 U7117 ( .A1(n7771), .A2(n6126), .ZN(n2004) );
  OAI21_X1 U7118 ( .B1(n16109), .B2(n2090), .A(n2089), .ZN(n15592) );
  NAND3_X1 U7119 ( .A1(n19427), .A2(n19760), .A3(n19176), .ZN(n2663) );
  OR2_X1 U7120 ( .A1(n22734), .A2(n23014), .ZN(n2709) );
  INV_X1 U7122 ( .A(n14697), .ZN(n14809) );
  INV_X1 U7123 ( .A(n6952), .ZN(n6949) );
  OR2_X1 U7124 ( .A1(n12447), .A2(n13165), .ZN(n3442) );
  AND2_X1 U7125 ( .A1(n7953), .A2(n7952), .ZN(n7956) );
  AOI21_X1 U7126 ( .B1(n14169), .B2(n14165), .A(n14164), .ZN(n4763) );
  OAI211_X1 U7127 ( .C1(n2529), .C2(n1477), .A(n2528), .B(n2527), .ZN(n23911)
         );
  INV_X1 U7128 ( .A(n19163), .ZN(n3727) );
  XNOR2_X1 U7130 ( .A(n21343), .B(n21344), .ZN(n2415) );
  INV_X1 U7131 ( .A(n17195), .ZN(n4039) );
  OR2_X1 U7132 ( .A1(n6699), .A2(n6697), .ZN(n6415) );
  NAND2_X1 U7133 ( .A1(n6699), .A2(n6556), .ZN(n2006) );
  AOI21_X1 U7135 ( .B1(n13482), .B2(n13769), .A(n4331), .ZN(n4330) );
  NAND2_X1 U7136 ( .A1(n293), .A2(n16095), .ZN(n16146) );
  NAND2_X1 U7138 ( .A1(n2009), .A2(n22487), .ZN(n22489) );
  NAND3_X1 U7139 ( .A1(n22895), .A2(n2326), .A3(n2327), .ZN(n2009) );
  NAND3_X1 U7140 ( .A1(n23314), .A2(n2919), .A3(n23319), .ZN(n23316) );
  OAI211_X2 U7141 ( .C1(n20000), .C2(n20539), .A(n19999), .B(n2012), .ZN(n3819) );
  OAI21_X1 U7142 ( .B1(n19998), .B2(n20150), .A(n20145), .ZN(n2012) );
  NAND2_X1 U7143 ( .A1(n2015), .A2(n2013), .ZN(n11551) );
  NAND2_X1 U7144 ( .A1(n12470), .A2(n11541), .ZN(n2013) );
  NAND2_X1 U7145 ( .A1(n11549), .A2(n13066), .ZN(n2015) );
  NOR2_X1 U7146 ( .A1(n13072), .A2(n12774), .ZN(n11549) );
  NAND2_X1 U7148 ( .A1(n19572), .A2(n20369), .ZN(n2017) );
  OAI211_X1 U7150 ( .C1(n2090), .C2(n16106), .A(n24928), .B(n2020), .ZN(n15629) );
  OAI21_X1 U7153 ( .B1(n7993), .B2(n7499), .A(n7501), .ZN(n7505) );
  NOR2_X1 U7154 ( .A1(n5573), .A2(n19275), .ZN(n19542) );
  NAND2_X1 U7157 ( .A1(n7457), .A2(n2022), .ZN(n8498) );
  OR2_X1 U7158 ( .A1(n7458), .A2(n7573), .ZN(n2022) );
  XNOR2_X1 U7159 ( .A(n25481), .B(n364), .ZN(n17590) );
  NAND2_X1 U7160 ( .A1(n10595), .A2(n1430), .ZN(n10597) );
  NAND3_X1 U7161 ( .A1(n2023), .A2(n2284), .A3(n5411), .ZN(n13997) );
  OR2_X1 U7162 ( .A1(n19908), .A2(n2024), .ZN(n2568) );
  AOI21_X1 U7163 ( .B1(n20412), .B2(n25420), .A(n19741), .ZN(n19908) );
  OR2_X1 U7164 ( .A1(n413), .A2(n10518), .ZN(n9291) );
  INV_X1 U7165 ( .A(n19530), .ZN(n5480) );
  NAND2_X1 U7168 ( .A1(n3407), .A2(n6324), .ZN(n2025) );
  OR2_X2 U7169 ( .A1(n6330), .A2(n6331), .ZN(n9066) );
  OAI21_X1 U7172 ( .B1(n7568), .B2(n7641), .A(n7567), .ZN(n2026) );
  NAND2_X1 U7173 ( .A1(n6936), .A2(n6560), .ZN(n2027) );
  NAND2_X1 U7174 ( .A1(n6697), .A2(n6699), .ZN(n6936) );
  NAND2_X1 U7175 ( .A1(n6935), .A2(n6934), .ZN(n2028) );
  XNOR2_X2 U7178 ( .A(n9163), .B(n9162), .ZN(n10138) );
  OR2_X1 U7179 ( .A1(n10176), .A2(n9829), .ZN(n9584) );
  INV_X1 U7180 ( .A(n20039), .ZN(n20185) );
  XNOR2_X1 U7181 ( .A(n9199), .B(n9200), .ZN(n9398) );
  NAND2_X1 U7182 ( .A1(n2030), .A2(n9703), .ZN(n9708) );
  NAND2_X1 U7183 ( .A1(n9702), .A2(n9705), .ZN(n2030) );
  NAND2_X1 U7184 ( .A1(n3677), .A2(n4259), .ZN(n3676) );
  NAND3_X1 U7186 ( .A1(n11885), .A2(n11149), .A3(n24480), .ZN(n5000) );
  AND2_X1 U7187 ( .A1(n17048), .A2(n17050), .ZN(n15956) );
  OR3_X1 U7188 ( .A1(n25081), .A2(n22932), .A3(n24342), .ZN(n21427) );
  NAND3_X1 U7189 ( .A1(n6439), .A2(n6296), .A3(n6438), .ZN(n5947) );
  NAND3_X1 U7190 ( .A1(n3763), .A2(n6147), .A3(n6940), .ZN(n5889) );
  INV_X1 U7193 ( .A(n16604), .ZN(n3817) );
  NAND2_X1 U7196 ( .A1(n2184), .A2(n10890), .ZN(n2766) );
  NAND2_X1 U7197 ( .A1(n4308), .A2(n278), .ZN(n4307) );
  OAI21_X1 U7198 ( .B1(n4442), .B2(n4441), .A(n22274), .ZN(n2038) );
  AOI22_X1 U7199 ( .A1(n9498), .A2(n10090), .B1(n1348), .B2(n9497), .ZN(n3088)
         );
  NOR2_X1 U7200 ( .A1(n5102), .A2(n14153), .ZN(n2775) );
  OAI21_X1 U7202 ( .B1(n6088), .B2(n6372), .A(n6900), .ZN(n6087) );
  NAND2_X1 U7203 ( .A1(n6088), .A2(n6473), .ZN(n6900) );
  NAND3_X1 U7204 ( .A1(n6196), .A2(n6019), .A3(n6347), .ZN(n6020) );
  XNOR2_X1 U7205 ( .A(n18580), .B(n18581), .ZN(n2041) );
  NOR2_X1 U7207 ( .A1(n20089), .A2(n20557), .ZN(n3482) );
  OAI211_X1 U7208 ( .C1(n7292), .C2(n5202), .A(n2522), .B(n2043), .ZN(n3681)
         );
  NAND2_X1 U7209 ( .A1(n5202), .A2(n432), .ZN(n2043) );
  NAND2_X1 U7210 ( .A1(n6478), .A2(n6873), .ZN(n2045) );
  MUX2_X1 U7211 ( .A(n12820), .B(n12821), .S(n14054), .Z(n12823) );
  NAND2_X1 U7212 ( .A1(n8525), .A2(n2046), .ZN(n11168) );
  XNOR2_X1 U7213 ( .A(n21582), .B(n20777), .ZN(n3038) );
  AOI22_X2 U7214 ( .A1(n19690), .A2(n19689), .B1(n2322), .B2(n20534), .ZN(
        n21582) );
  NAND2_X1 U7215 ( .A1(n19503), .A2(n358), .ZN(n19504) );
  OR2_X1 U7216 ( .A1(n1355), .A2(n14049), .ZN(n12821) );
  OAI21_X1 U7217 ( .B1(n9500), .B2(n10000), .A(n9499), .ZN(n10775) );
  NAND2_X1 U7218 ( .A1(n9671), .A2(n9798), .ZN(n10000) );
  AND2_X2 U7219 ( .A1(n15969), .A2(n15968), .ZN(n17572) );
  NOR2_X1 U7220 ( .A1(n13159), .A2(n12440), .ZN(n13062) );
  INV_X1 U7221 ( .A(n13837), .ZN(n14271) );
  OR2_X1 U7222 ( .A1(n24974), .A2(n13907), .ZN(n13949) );
  NAND2_X1 U7223 ( .A1(n3214), .A2(n19787), .ZN(n3962) );
  INV_X1 U7224 ( .A(n9787), .ZN(n4256) );
  OR2_X1 U7225 ( .A1(n7414), .A2(n3549), .ZN(n5329) );
  XNOR2_X1 U7226 ( .A(n11658), .B(n2047), .ZN(n10949) );
  XNOR2_X1 U7227 ( .A(n10923), .B(n11942), .ZN(n2047) );
  OR2_X1 U7228 ( .A1(n13323), .A2(n2295), .ZN(n12684) );
  NAND2_X1 U7229 ( .A1(n2051), .A2(n16397), .ZN(n3628) );
  INV_X1 U7231 ( .A(n25198), .ZN(n13244) );
  XNOR2_X1 U7232 ( .A(n2052), .B(n18176), .ZN(n18180) );
  INV_X1 U7233 ( .A(n18588), .ZN(n2052) );
  OAI21_X1 U7234 ( .B1(n5704), .B2(n7329), .A(n7897), .ZN(n5703) );
  INV_X1 U7235 ( .A(n4291), .ZN(n18934) );
  XNOR2_X1 U7236 ( .A(n15219), .B(n14724), .ZN(n15319) );
  XNOR2_X1 U7237 ( .A(n24976), .B(n2242), .ZN(n14715) );
  INV_X1 U7238 ( .A(n7477), .ZN(n4144) );
  INV_X1 U7239 ( .A(n20401), .ZN(n5590) );
  INV_X1 U7240 ( .A(n21751), .ZN(n21231) );
  OAI22_X1 U7241 ( .A1(n3503), .A2(n3410), .B1(n5459), .B2(n16105), .ZN(n15798) );
  NOR2_X1 U7242 ( .A1(n13325), .A2(n13323), .ZN(n12955) );
  INV_X1 U7243 ( .A(n14667), .ZN(n3232) );
  INV_X1 U7244 ( .A(n17312), .ZN(n17599) );
  XNOR2_X1 U7245 ( .A(n8119), .B(n5328), .ZN(n8439) );
  XNOR2_X1 U7246 ( .A(n21591), .B(n4263), .ZN(n20212) );
  XNOR2_X1 U7247 ( .A(n2053), .B(n3901), .ZN(Ciphertext[12]) );
  OAI21_X1 U7248 ( .B1(n22480), .B2(n23112), .A(n22479), .ZN(n2053) );
  NAND2_X1 U7249 ( .A1(n17180), .A2(n16368), .ZN(n16205) );
  OAI21_X1 U7251 ( .B1(n17416), .B2(n17415), .A(n17419), .ZN(n2055) );
  OAI21_X1 U7253 ( .B1(n7261), .B2(n7923), .A(n2056), .ZN(n7446) );
  NAND2_X1 U7254 ( .A1(n7923), .A2(n7932), .ZN(n2056) );
  NAND2_X1 U7256 ( .A1(n16704), .A2(n16708), .ZN(n2057) );
  NAND3_X1 U7257 ( .A1(n11884), .A2(n11145), .A3(n2059), .ZN(n10535) );
  NOR2_X1 U7258 ( .A1(n11152), .A2(n2060), .ZN(n2059) );
  NAND2_X1 U7264 ( .A1(n6522), .A2(n25398), .ZN(n2061) );
  NAND2_X1 U7266 ( .A1(n16844), .A2(n16991), .ZN(n2062) );
  INV_X1 U7267 ( .A(n13260), .ZN(n3791) );
  OR2_X1 U7269 ( .A1(n25046), .A2(n10170), .ZN(n9816) );
  NAND2_X1 U7270 ( .A1(n21840), .A2(n24362), .ZN(n2066) );
  NAND2_X2 U7271 ( .A1(n19585), .A2(n2067), .ZN(n20451) );
  NAND2_X1 U7272 ( .A1(n2069), .A2(n2068), .ZN(n2067) );
  INV_X1 U7274 ( .A(n14075), .ZN(n14079) );
  NOR2_X1 U7275 ( .A1(n24586), .A2(n16109), .ZN(n5464) );
  NOR2_X1 U7277 ( .A1(n15783), .A2(n379), .ZN(n15590) );
  XNOR2_X1 U7278 ( .A(n2070), .B(n14452), .ZN(n14453) );
  XNOR2_X1 U7279 ( .A(n14451), .B(n15188), .ZN(n2070) );
  NAND3_X2 U7281 ( .A1(n10002), .A2(n9800), .A3(n9801), .ZN(n11499) );
  NAND3_X1 U7282 ( .A1(n20299), .A2(n2074), .A3(n2073), .ZN(n4932) );
  NAND2_X1 U7283 ( .A1(n19979), .A2(n20298), .ZN(n2073) );
  INV_X1 U7284 ( .A(n12717), .ZN(n10532) );
  NAND2_X1 U7285 ( .A1(n13169), .A2(n4766), .ZN(n12717) );
  NAND2_X1 U7286 ( .A1(n16683), .A2(n16681), .ZN(n17272) );
  NAND2_X1 U7287 ( .A1(n2076), .A2(n2075), .ZN(n16683) );
  NAND2_X1 U7288 ( .A1(n16082), .A2(n16102), .ZN(n2075) );
  NAND2_X1 U7289 ( .A1(n6122), .A2(n6245), .ZN(n6989) );
  XNOR2_X1 U7290 ( .A(n25234), .B(n25371), .ZN(n12372) );
  NAND3_X1 U7291 ( .A1(n10140), .A2(n10142), .A3(n10141), .ZN(n10143) );
  INV_X1 U7292 ( .A(n11905), .ZN(n2077) );
  NOR2_X1 U7294 ( .A1(n10048), .A2(n10046), .ZN(n2079) );
  NAND2_X1 U7296 ( .A1(n7982), .A2(n7985), .ZN(n2081) );
  NAND2_X1 U7297 ( .A1(n4071), .A2(n23256), .ZN(n2083) );
  NAND2_X1 U7298 ( .A1(n23218), .A2(n23217), .ZN(n2084) );
  NAND2_X1 U7299 ( .A1(n21368), .A2(n20649), .ZN(n4352) );
  OAI21_X1 U7300 ( .B1(n341), .B2(n20316), .A(n2913), .ZN(n20323) );
  NOR2_X2 U7304 ( .A1(n12589), .A2(n12588), .ZN(n14063) );
  XNOR2_X1 U7305 ( .A(n2085), .B(n8050), .ZN(n8053) );
  XNOR2_X1 U7306 ( .A(n8049), .B(n25407), .ZN(n2085) );
  OR2_X1 U7308 ( .A1(n7279), .A2(n7250), .ZN(n2749) );
  INV_X1 U7309 ( .A(n11369), .ZN(n14298) );
  INV_X1 U7310 ( .A(n23772), .ZN(n23782) );
  XNOR2_X1 U7311 ( .A(n14689), .B(n14815), .ZN(n2969) );
  MUX2_X2 U7312 ( .A(n6701), .B(n6700), .S(n6934), .Z(n7992) );
  XNOR2_X1 U7313 ( .A(n2088), .B(n22986), .ZN(Ciphertext[165]) );
  NOR2_X1 U7314 ( .A1(n22984), .A2(n22985), .ZN(n2088) );
  OR2_X1 U7315 ( .A1(n6146), .A2(n5887), .ZN(n6682) );
  XNOR2_X1 U7316 ( .A(n12212), .B(n12213), .ZN(n12215) );
  NAND2_X1 U7317 ( .A1(n6601), .A2(n6827), .ZN(n6230) );
  NAND2_X1 U7318 ( .A1(n16106), .A2(n16109), .ZN(n2089) );
  OAI21_X1 U7319 ( .B1(n22634), .B2(n24389), .A(n21943), .ZN(n21951) );
  OAI211_X1 U7321 ( .C1(n25064), .C2(n1577), .A(n24599), .B(n2091), .ZN(n2999)
         );
  NAND2_X1 U7322 ( .A1(n4933), .A2(n4932), .ZN(n19978) );
  XNOR2_X1 U7323 ( .A(n8557), .B(n8826), .ZN(n8441) );
  OR2_X1 U7324 ( .A1(n5051), .A2(n7889), .ZN(n2092) );
  NAND2_X1 U7327 ( .A1(n20143), .A2(n5445), .ZN(n5444) );
  NAND3_X1 U7329 ( .A1(n3189), .A2(n4488), .A3(n17256), .ZN(n17259) );
  NOR2_X1 U7330 ( .A1(n19446), .A2(n19449), .ZN(n5233) );
  INV_X1 U7332 ( .A(n6533), .ZN(n4199) );
  OR2_X1 U7333 ( .A1(n25046), .A2(n10166), .ZN(n9588) );
  NAND3_X1 U7334 ( .A1(n16813), .A2(n16814), .A3(n24410), .ZN(n16816) );
  NAND2_X1 U7335 ( .A1(n6755), .A2(n6757), .ZN(n6756) );
  NOR2_X1 U7336 ( .A1(n16186), .A2(n16397), .ZN(n15828) );
  NAND3_X1 U7337 ( .A1(n25061), .A2(n1353), .A3(n12454), .ZN(n3969) );
  NAND2_X1 U7338 ( .A1(n2625), .A2(n5570), .ZN(n19743) );
  NAND2_X1 U7339 ( .A1(n2095), .A2(n2094), .ZN(n13523) );
  NAND2_X1 U7340 ( .A1(n13520), .A2(n25247), .ZN(n2094) );
  NAND2_X1 U7341 ( .A1(n13519), .A2(n14054), .ZN(n2095) );
  NAND3_X1 U7343 ( .A1(n6753), .A2(n6754), .A3(n3276), .ZN(n3274) );
  NAND2_X1 U7345 ( .A1(n10648), .A2(n10649), .ZN(n10650) );
  NAND3_X1 U7346 ( .A1(n6408), .A2(n6412), .A3(n6409), .ZN(n6411) );
  NAND2_X1 U7347 ( .A1(n2096), .A2(n16036), .ZN(n5308) );
  INV_X1 U7349 ( .A(n8436), .ZN(n9001) );
  AND2_X1 U7350 ( .A1(n13940), .A2(n16397), .ZN(n16400) );
  NOR2_X1 U7351 ( .A1(n10790), .A2(n11199), .ZN(n4625) );
  OAI21_X1 U7352 ( .B1(n24092), .B2(n10053), .A(n4097), .ZN(n9870) );
  NAND3_X1 U7354 ( .A1(n15542), .A2(n15543), .A3(n15544), .ZN(n15873) );
  INV_X1 U7355 ( .A(n13418), .ZN(n4895) );
  NAND3_X1 U7356 ( .A1(n2099), .A2(n13105), .A3(n12743), .ZN(n12746) );
  NAND2_X1 U7357 ( .A1(n12741), .A2(n13183), .ZN(n2099) );
  NAND2_X1 U7358 ( .A1(n3701), .A2(n13569), .ZN(n3700) );
  OAI21_X1 U7359 ( .B1(n13713), .B2(n3699), .A(n3697), .ZN(n13396) );
  NAND3_X1 U7360 ( .A1(n5025), .A2(n5026), .A3(n425), .ZN(n4561) );
  XNOR2_X1 U7361 ( .A(n8542), .B(n9044), .ZN(n8543) );
  NAND2_X1 U7362 ( .A1(n6952), .A2(n5903), .ZN(n5905) );
  XNOR2_X2 U7363 ( .A(n5791), .B(Key[89]), .ZN(n6114) );
  INV_X1 U7364 ( .A(n2546), .ZN(n10497) );
  INV_X1 U7365 ( .A(n23342), .ZN(n22961) );
  OR2_X1 U7366 ( .A1(n15594), .A2(n24826), .ZN(n15598) );
  INV_X1 U7367 ( .A(n16901), .ZN(n2566) );
  INV_X1 U7369 ( .A(n10772), .ZN(n4281) );
  NAND2_X1 U7370 ( .A1(n2102), .A2(n2101), .ZN(n6582) );
  NAND2_X1 U7371 ( .A1(n6758), .A2(n6675), .ZN(n2101) );
  NAND2_X1 U7372 ( .A1(n5804), .A2(n6751), .ZN(n2102) );
  XNOR2_X2 U7374 ( .A(n19738), .B(n19737), .ZN(n21848) );
  INV_X1 U7377 ( .A(n19854), .ZN(n2104) );
  AND3_X2 U7379 ( .A1(n2515), .A2(n2516), .A3(n2517), .ZN(n14945) );
  NOR2_X1 U7381 ( .A1(n16848), .A2(n17140), .ZN(n2105) );
  NAND3_X1 U7382 ( .A1(n1377), .A2(n3691), .A3(n13013), .ZN(n3690) );
  NAND2_X1 U7383 ( .A1(n4177), .A2(n6616), .ZN(n6617) );
  NAND2_X1 U7385 ( .A1(n7364), .A2(n7628), .ZN(n7627) );
  OR2_X1 U7387 ( .A1(n13124), .A2(n13350), .ZN(n12873) );
  NAND3_X1 U7388 ( .A1(n10943), .A2(n3760), .A3(n10944), .ZN(n10945) );
  XNOR2_X2 U7389 ( .A(n18036), .B(n18035), .ZN(n19598) );
  XNOR2_X1 U7390 ( .A(n2106), .B(n23657), .ZN(Ciphertext[124]) );
  NAND3_X1 U7391 ( .A1(n23656), .A2(n23654), .A3(n23655), .ZN(n2106) );
  NAND3_X1 U7392 ( .A1(n11876), .A2(n11874), .A3(n11875), .ZN(n13597) );
  NAND2_X1 U7393 ( .A1(n16135), .A2(n2107), .ZN(n18277) );
  NAND2_X1 U7394 ( .A1(n17527), .A2(n17170), .ZN(n2107) );
  NAND2_X1 U7395 ( .A1(n4678), .A2(n24532), .ZN(n4677) );
  OAI21_X1 U7396 ( .B1(n8522), .B2(n9999), .A(n2108), .ZN(n3261) );
  NAND3_X1 U7397 ( .A1(n9310), .A2(n4137), .A3(n8521), .ZN(n2108) );
  NAND2_X1 U7398 ( .A1(n14002), .A2(n14003), .ZN(n14006) );
  AOI21_X1 U7400 ( .B1(n2109), .B2(n6030), .A(n6512), .ZN(n5941) );
  NAND2_X1 U7401 ( .A1(n6454), .A2(n6456), .ZN(n2109) );
  NAND3_X1 U7402 ( .A1(n3100), .A2(n10801), .A3(n10648), .ZN(n10246) );
  NAND3_X1 U7403 ( .A1(n4342), .A2(n10899), .A3(n4341), .ZN(n4343) );
  OAI21_X1 U7404 ( .B1(n2112), .B2(n285), .A(n2111), .ZN(n2110) );
  INV_X1 U7405 ( .A(n4039), .ZN(n2111) );
  INV_X1 U7406 ( .A(n4869), .ZN(n4574) );
  XNOR2_X1 U7407 ( .A(n15398), .B(n15495), .ZN(n2113) );
  NAND2_X1 U7408 ( .A1(n24532), .A2(n25030), .ZN(n2478) );
  NAND2_X1 U7410 ( .A1(n11407), .A2(n11408), .ZN(n2116) );
  NAND2_X1 U7411 ( .A1(n6734), .A2(n6730), .ZN(n2118) );
  INV_X1 U7412 ( .A(n16526), .ZN(n16832) );
  OR2_X1 U7413 ( .A1(n523), .A2(n17450), .ZN(n2121) );
  NAND2_X1 U7414 ( .A1(n16979), .A2(n17450), .ZN(n16526) );
  NAND3_X1 U7415 ( .A1(n3575), .A2(n4358), .A3(n10902), .ZN(n4357) );
  NOR2_X1 U7417 ( .A1(n5315), .A2(n2246), .ZN(n16904) );
  NAND3_X1 U7420 ( .A1(n25323), .A2(n16197), .A3(n24482), .ZN(n5165) );
  MUX2_X2 U7421 ( .A(n19718), .B(n19717), .S(n20117), .Z(n21297) );
  XNOR2_X2 U7422 ( .A(n8229), .B(n8228), .ZN(n9832) );
  AOI22_X1 U7423 ( .A1(n17323), .A2(n4426), .B1(n15673), .B2(n17320), .ZN(
        n17269) );
  NOR2_X1 U7424 ( .A1(n7013), .A2(n25045), .ZN(n6600) );
  AND2_X1 U7425 ( .A1(n3358), .A2(n7948), .ZN(n4812) );
  NOR2_X2 U7426 ( .A1(n19527), .A2(n19528), .ZN(n20370) );
  XNOR2_X1 U7427 ( .A(n24508), .B(n14805), .ZN(n3940) );
  INV_X1 U7428 ( .A(n22575), .ZN(n23202) );
  OR2_X1 U7429 ( .A1(n14205), .A2(n13549), .ZN(n2214) );
  XNOR2_X1 U7430 ( .A(n14972), .B(n14971), .ZN(n4115) );
  OAI211_X1 U7431 ( .C1(n24310), .C2(n19606), .A(n4141), .B(n19608), .ZN(n2764) );
  INV_X1 U7433 ( .A(n13978), .ZN(n13391) );
  NAND2_X1 U7435 ( .A1(n2128), .A2(n2127), .ZN(n7226) );
  NAND2_X1 U7436 ( .A1(n7225), .A2(n25251), .ZN(n2127) );
  NAND2_X1 U7437 ( .A1(n3275), .A2(n7677), .ZN(n2128) );
  INV_X1 U7438 ( .A(n13583), .ZN(n4868) );
  MUX2_X2 U7439 ( .A(n6251), .B(n6250), .S(n7734), .Z(n8806) );
  NAND2_X1 U7440 ( .A1(n2130), .A2(n2129), .ZN(n10546) );
  NAND2_X1 U7441 ( .A1(n10540), .A2(n10302), .ZN(n2129) );
  NAND2_X1 U7442 ( .A1(n10539), .A2(n2389), .ZN(n2130) );
  NAND3_X1 U7443 ( .A1(n3791), .A2(n3792), .A3(n2131), .ZN(n13450) );
  NAND2_X1 U7444 ( .A1(n13257), .A2(n13974), .ZN(n2131) );
  NAND4_X2 U7449 ( .A1(n7202), .A2(n7201), .A3(n7203), .A4(n7620), .ZN(n4378)
         );
  NOR2_X1 U7450 ( .A1(n4812), .A2(n4093), .ZN(n3359) );
  NAND2_X1 U7451 ( .A1(n19391), .A2(n19389), .ZN(n2132) );
  NAND2_X1 U7452 ( .A1(n5710), .A2(n20474), .ZN(n5711) );
  NAND2_X1 U7453 ( .A1(n5556), .A2(n5557), .ZN(n5555) );
  OR2_X1 U7454 ( .A1(n7384), .A2(n7619), .ZN(n7621) );
  NAND2_X1 U7455 ( .A1(n17063), .A2(n24385), .ZN(n2133) );
  NAND2_X1 U7456 ( .A1(n17064), .A2(n17054), .ZN(n2134) );
  NAND2_X1 U7457 ( .A1(n4692), .A2(n19681), .ZN(n2136) );
  NOR2_X1 U7460 ( .A1(n20278), .A2(n20345), .ZN(n2138) );
  NAND2_X1 U7461 ( .A1(n6810), .A2(n2139), .ZN(n8353) );
  OR2_X1 U7462 ( .A1(n436), .A2(n8530), .ZN(n2139) );
  NAND2_X1 U7463 ( .A1(n6547), .A2(n6546), .ZN(n6805) );
  NOR2_X1 U7464 ( .A1(n9796), .A2(n9798), .ZN(n2140) );
  XNOR2_X1 U7465 ( .A(n14443), .B(n3695), .ZN(n3694) );
  NAND2_X1 U7466 ( .A1(n7101), .A2(n6133), .ZN(n6134) );
  NAND2_X1 U7467 ( .A1(n2388), .A2(n10302), .ZN(n4327) );
  NAND3_X1 U7468 ( .A1(n10541), .A2(n24345), .A3(n10301), .ZN(n10213) );
  NAND2_X1 U7469 ( .A1(n2142), .A2(n2141), .ZN(n22386) );
  NAND2_X1 U7470 ( .A1(n22384), .A2(n23318), .ZN(n2141) );
  NAND2_X1 U7471 ( .A1(n2143), .A2(n23317), .ZN(n2142) );
  NAND3_X1 U7473 ( .A1(n9474), .A2(n9857), .A3(n239), .ZN(n9476) );
  NAND3_X1 U7474 ( .A1(n5402), .A2(n3339), .A3(n12631), .ZN(n3338) );
  OAI21_X1 U7475 ( .B1(n3404), .B2(n3401), .A(n14320), .ZN(n13602) );
  AOI22_X1 U7476 ( .A1(n16354), .A2(n16980), .B1(n17453), .B2(n16979), .ZN(
        n16370) );
  NAND2_X1 U7477 ( .A1(n7450), .A2(n7155), .ZN(n7630) );
  NAND2_X1 U7478 ( .A1(n4439), .A2(n19597), .ZN(n4438) );
  INV_X1 U7480 ( .A(n5649), .ZN(n5648) );
  NAND3_X1 U7481 ( .A1(n6636), .A2(n7021), .A3(n7027), .ZN(n2146) );
  NAND2_X1 U7482 ( .A1(n6638), .A2(n6637), .ZN(n2147) );
  AND2_X1 U7483 ( .A1(n7008), .A2(n7004), .ZN(n6095) );
  NAND3_X1 U7484 ( .A1(n15814), .A2(n16206), .A3(n3380), .ZN(n15643) );
  NAND2_X1 U7485 ( .A1(n11163), .A2(n10552), .ZN(n2148) );
  NAND3_X1 U7486 ( .A1(n9721), .A2(n9725), .A3(n10005), .ZN(n9654) );
  MUX2_X1 U7487 ( .A(n15673), .B(n17319), .S(n17320), .Z(n17325) );
  NAND2_X2 U7488 ( .A1(n2288), .A2(n2163), .ZN(n17320) );
  OR2_X1 U7489 ( .A1(n6325), .A2(n25398), .ZN(n2149) );
  INV_X1 U7490 ( .A(n15893), .ZN(n13374) );
  NAND2_X1 U7491 ( .A1(n24080), .A2(n16595), .ZN(n15893) );
  NAND2_X1 U7493 ( .A1(n12467), .A2(n13521), .ZN(n2150) );
  NAND2_X1 U7494 ( .A1(n13611), .A2(n14058), .ZN(n2151) );
  INV_X1 U7495 ( .A(n17686), .ZN(n17689) );
  NAND2_X1 U7496 ( .A1(n17484), .A2(n17730), .ZN(n17686) );
  INV_X1 U7497 ( .A(n17414), .ZN(n17224) );
  INV_X1 U7498 ( .A(n10064), .ZN(n9704) );
  XNOR2_X1 U7499 ( .A(n12020), .B(n12183), .ZN(n11699) );
  XNOR2_X1 U7500 ( .A(n18004), .B(n2964), .ZN(n18005) );
  NAND3_X1 U7502 ( .A1(n16235), .A2(n16449), .A3(n15725), .ZN(n15729) );
  NAND3_X1 U7503 ( .A1(n4198), .A2(n17461), .A3(n16021), .ZN(n16993) );
  OAI21_X1 U7506 ( .B1(n13026), .B2(n13029), .A(n13025), .ZN(n2153) );
  XNOR2_X1 U7507 ( .A(n18680), .B(n2154), .ZN(n18681) );
  XNOR2_X1 U7508 ( .A(n3703), .B(n18679), .ZN(n2154) );
  AND2_X1 U7509 ( .A1(n12541), .A2(n12540), .ZN(n12810) );
  NAND2_X1 U7510 ( .A1(n2157), .A2(n2156), .ZN(n10580) );
  NAND2_X1 U7511 ( .A1(n11525), .A2(n11529), .ZN(n2156) );
  NAND2_X1 U7512 ( .A1(n1332), .A2(n11026), .ZN(n2157) );
  NAND2_X1 U7514 ( .A1(n23820), .A2(n23810), .ZN(n23821) );
  NAND2_X1 U7516 ( .A1(n6697), .A2(n6560), .ZN(n5907) );
  NAND2_X1 U7517 ( .A1(n24958), .A2(n24572), .ZN(n13619) );
  NOR2_X2 U7519 ( .A1(n8752), .A2(n2159), .ZN(n11520) );
  OAI21_X1 U7520 ( .B1(n9766), .B2(n9763), .A(n8751), .ZN(n2159) );
  XNOR2_X1 U7521 ( .A(n9073), .B(n5614), .ZN(n8125) );
  XNOR2_X1 U7522 ( .A(n4025), .B(n8981), .ZN(n4024) );
  OR2_X1 U7523 ( .A1(n10886), .A2(n10887), .ZN(n3221) );
  XNOR2_X1 U7527 ( .A(n17660), .B(n18626), .ZN(n2335) );
  AND3_X2 U7528 ( .A1(n4522), .A2(n4521), .A3(n4523), .ZN(n11059) );
  OAI211_X1 U7529 ( .C1(n9507), .C2(n9786), .A(n2486), .B(n24575), .ZN(n4522)
         );
  AOI21_X2 U7530 ( .B1(n16987), .B2(n16986), .A(n2161), .ZN(n18513) );
  NOR2_X1 U7531 ( .A1(n4392), .A2(n4391), .ZN(n4390) );
  XNOR2_X1 U7532 ( .A(n2162), .B(n21448), .ZN(n19161) );
  XNOR2_X1 U7533 ( .A(n19124), .B(n21541), .ZN(n2162) );
  OR2_X1 U7534 ( .A1(n14522), .A2(n16116), .ZN(n2935) );
  INV_X1 U7535 ( .A(n16246), .ZN(n2605) );
  OR2_X1 U7536 ( .A1(n15672), .A2(n15887), .ZN(n2163) );
  OAI22_X1 U7537 ( .A1(n7126), .A2(n7581), .B1(n7879), .B2(n7582), .ZN(n7124)
         );
  NAND2_X1 U7538 ( .A1(n10054), .A2(n10053), .ZN(n10055) );
  NAND2_X1 U7539 ( .A1(n2165), .A2(n2164), .ZN(n7934) );
  OR2_X1 U7540 ( .A1(n11023), .A2(n8934), .ZN(n10920) );
  NAND2_X1 U7541 ( .A1(n6020), .A2(n6021), .ZN(n2166) );
  NAND2_X1 U7542 ( .A1(n2167), .A2(n414), .ZN(n5516) );
  NAND2_X1 U7543 ( .A1(n2675), .A2(n11206), .ZN(n2167) );
  OR2_X2 U7544 ( .A1(n3166), .A2(n10022), .ZN(n11044) );
  OAI21_X1 U7545 ( .B1(n12534), .B2(n13048), .A(n25494), .ZN(n2639) );
  NAND2_X1 U7547 ( .A1(n20194), .A2(n19744), .ZN(n2169) );
  NAND2_X1 U7548 ( .A1(n2171), .A2(n14090), .ZN(n2170) );
  NAND2_X1 U7549 ( .A1(n14088), .A2(n14089), .ZN(n2171) );
  NAND2_X1 U7550 ( .A1(n14091), .A2(n2321), .ZN(n2172) );
  XNOR2_X1 U7551 ( .A(n2174), .B(n22697), .ZN(Ciphertext[185]) );
  OAI21_X1 U7552 ( .B1(n22696), .B2(n25076), .A(n22695), .ZN(n2174) );
  INV_X1 U7554 ( .A(n13228), .ZN(n4587) );
  NAND3_X1 U7555 ( .A1(n7540), .A2(n2522), .A3(n8006), .ZN(n5203) );
  NAND2_X1 U7556 ( .A1(n17252), .A2(n17272), .ZN(n17282) );
  NOR2_X2 U7557 ( .A1(n6127), .A2(n2175), .ZN(n8824) );
  OR2_X2 U7559 ( .A1(n5141), .A2(n12072), .ZN(n14306) );
  INV_X1 U7561 ( .A(n13490), .ZN(n3071) );
  INV_X1 U7562 ( .A(n7972), .ZN(n7514) );
  INV_X1 U7563 ( .A(n18080), .ZN(n3990) );
  AND3_X2 U7564 ( .A1(n4352), .A2(n3476), .A3(n4349), .ZN(n23218) );
  NAND2_X1 U7565 ( .A1(n2177), .A2(n2176), .ZN(n4801) );
  NAND2_X1 U7566 ( .A1(n4400), .A2(n7972), .ZN(n2176) );
  NAND2_X1 U7568 ( .A1(n25360), .A2(n2178), .ZN(n12702) );
  NAND2_X1 U7569 ( .A1(n2180), .A2(n2179), .ZN(n20321) );
  OAI21_X1 U7571 ( .B1(n16869), .B2(n16870), .A(n17196), .ZN(n2183) );
  NOR2_X1 U7572 ( .A1(n2185), .A2(n11084), .ZN(n2184) );
  NAND3_X1 U7573 ( .A1(n3984), .A2(n1425), .A3(n3987), .ZN(n20533) );
  XNOR2_X1 U7574 ( .A(n2186), .B(n21696), .ZN(n18861) );
  XNOR2_X1 U7575 ( .A(n18746), .B(n21247), .ZN(n2186) );
  NAND2_X1 U7576 ( .A1(n2188), .A2(n2187), .ZN(n22458) );
  NAND2_X1 U7577 ( .A1(n22456), .A2(n22455), .ZN(n2187) );
  NAND2_X1 U7580 ( .A1(n14945), .A2(n14944), .ZN(n13801) );
  MUX2_X1 U7581 ( .A(n17346), .B(n17345), .S(n17344), .Z(n17350) );
  NAND2_X1 U7582 ( .A1(n17240), .A2(n15314), .ZN(n17344) );
  NAND2_X1 U7583 ( .A1(n20039), .A2(n25478), .ZN(n18729) );
  OR2_X1 U7584 ( .A1(n16145), .A2(n16095), .ZN(n2541) );
  INV_X1 U7586 ( .A(n12850), .ZN(n14025) );
  NAND2_X1 U7587 ( .A1(n6623), .A2(n316), .ZN(n6621) );
  NAND4_X1 U7588 ( .A1(n3708), .A2(n4707), .A3(n8351), .A4(n4706), .ZN(n4709)
         );
  XNOR2_X1 U7589 ( .A(n2194), .B(n21613), .ZN(n22027) );
  XNOR2_X1 U7590 ( .A(n21612), .B(n21611), .ZN(n2194) );
  NAND3_X1 U7591 ( .A1(n6684), .A2(n6944), .A3(n6683), .ZN(n6685) );
  NAND2_X1 U7592 ( .A1(n7582), .A2(n7313), .ZN(n7583) );
  NAND2_X1 U7593 ( .A1(n5138), .A2(n5139), .ZN(n5137) );
  NAND2_X1 U7594 ( .A1(n2195), .A2(n7598), .ZN(n7259) );
  NAND2_X1 U7595 ( .A1(n7258), .A2(n7595), .ZN(n2195) );
  NAND2_X1 U7596 ( .A1(n16122), .A2(n16123), .ZN(n15846) );
  NAND3_X1 U7600 ( .A1(n22742), .A2(n22743), .A3(n2199), .ZN(n22746) );
  XNOR2_X2 U7604 ( .A(n2203), .B(n3107), .ZN(n10128) );
  XNOR2_X1 U7605 ( .A(n7471), .B(n8703), .ZN(n2203) );
  INV_X1 U7606 ( .A(n12951), .ZN(n3256) );
  OAI21_X1 U7607 ( .B1(n19084), .B2(n24584), .A(n2204), .ZN(n19000) );
  NAND2_X1 U7608 ( .A1(n19084), .A2(n19418), .ZN(n2204) );
  NAND3_X1 U7609 ( .A1(n4159), .A2(n4163), .A3(n4162), .ZN(n4158) );
  INV_X1 U7610 ( .A(n13167), .ZN(n3688) );
  XNOR2_X1 U7611 ( .A(n2206), .B(n20628), .ZN(n20083) );
  XNOR2_X1 U7612 ( .A(n25202), .B(n20047), .ZN(n2206) );
  XNOR2_X2 U7613 ( .A(n15243), .B(n15242), .ZN(n16324) );
  NAND2_X1 U7614 ( .A1(n6588), .A2(n7029), .ZN(n6225) );
  NAND2_X1 U7615 ( .A1(n6615), .A2(n6063), .ZN(n2400) );
  INV_X1 U7616 ( .A(n14104), .ZN(n14816) );
  OAI21_X1 U7617 ( .B1(n22812), .B2(n22606), .A(n22810), .ZN(n2529) );
  OR2_X1 U7619 ( .A1(n6296), .A2(n6297), .ZN(n4865) );
  NAND3_X1 U7620 ( .A1(n2493), .A2(n13216), .A3(n4651), .ZN(n4546) );
  NAND2_X1 U7621 ( .A1(n6722), .A2(n6243), .ZN(n6721) );
  NAND2_X1 U7622 ( .A1(n16382), .A2(n15837), .ZN(n15990) );
  NAND2_X1 U7623 ( .A1(n7107), .A2(n7250), .ZN(n5928) );
  NAND2_X1 U7624 ( .A1(n24576), .A2(n7862), .ZN(n7708) );
  NAND3_X1 U7625 ( .A1(n22330), .A2(n22329), .A3(n22464), .ZN(n22331) );
  NAND2_X1 U7626 ( .A1(n6969), .A2(n6570), .ZN(n6057) );
  MUX2_X2 U7627 ( .A(n14114), .B(n14113), .S(n14112), .Z(n15082) );
  XNOR2_X2 U7628 ( .A(n8976), .B(n4070), .ZN(n9681) );
  OAI21_X1 U7629 ( .B1(n5368), .B2(n2209), .A(n2639), .ZN(n12536) );
  NAND2_X1 U7630 ( .A1(n4094), .A2(n13049), .ZN(n2209) );
  INV_X1 U7631 ( .A(n14265), .ZN(n5694) );
  INV_X1 U7632 ( .A(n8296), .ZN(n2273) );
  OAI22_X1 U7634 ( .A1(n12584), .A2(n12625), .B1(n12981), .B2(n13363), .ZN(
        n12585) );
  XNOR2_X1 U7636 ( .A(n2210), .B(n20794), .ZN(n20796) );
  XNOR2_X1 U7637 ( .A(n20793), .B(n21115), .ZN(n2210) );
  INV_X1 U7638 ( .A(n7348), .ZN(n5468) );
  OAI21_X1 U7639 ( .B1(n20823), .B2(n23217), .A(n20824), .ZN(n3086) );
  OAI21_X1 U7640 ( .B1(n4017), .B2(n20093), .A(n20023), .ZN(n20025) );
  INV_X1 U7641 ( .A(n14943), .ZN(n2684) );
  NAND2_X1 U7643 ( .A1(n3588), .A2(n7533), .ZN(n4296) );
  OAI22_X1 U7644 ( .A1(n21834), .A2(n3231), .B1(n21835), .B2(n21836), .ZN(
        n3227) );
  OAI211_X1 U7645 ( .C1(n16021), .C2(n17461), .A(n3114), .B(n5052), .ZN(n3112)
         );
  NAND3_X1 U7647 ( .A1(n15611), .A2(n15612), .A3(n16120), .ZN(n2212) );
  XNOR2_X1 U7648 ( .A(n2213), .B(n12025), .ZN(n12026) );
  XNOR2_X1 U7649 ( .A(n12184), .B(n12024), .ZN(n2213) );
  NAND2_X1 U7650 ( .A1(n2309), .A2(n10933), .ZN(n2308) );
  OR2_X1 U7651 ( .A1(n12911), .A2(n13288), .ZN(n12694) );
  NAND2_X1 U7652 ( .A1(n7961), .A2(n7683), .ZN(n7684) );
  OR2_X1 U7654 ( .A1(n16129), .A2(n16076), .ZN(n14662) );
  NAND3_X2 U7655 ( .A1(n10591), .A2(n10593), .A3(n10592), .ZN(n12127) );
  XOR2_X1 U7657 ( .A(n18149), .B(n3118), .Z(n5327) );
  NOR2_X1 U7658 ( .A1(n1353), .A2(n13162), .ZN(n5011) );
  NAND2_X1 U7659 ( .A1(n19098), .A2(n19367), .ZN(n17801) );
  NAND2_X1 U7660 ( .A1(n2219), .A2(n2218), .ZN(n2217) );
  NAND2_X1 U7661 ( .A1(n6350), .A2(n6271), .ZN(n2219) );
  NAND2_X1 U7663 ( .A1(n2221), .A2(n6346), .ZN(n6348) );
  NAND2_X1 U7664 ( .A1(n6345), .A2(n6445), .ZN(n2221) );
  NAND2_X1 U7666 ( .A1(n7124), .A2(n7123), .ZN(n2224) );
  INV_X1 U7667 ( .A(n18796), .ZN(n19281) );
  XNOR2_X1 U7669 ( .A(n14724), .B(n2145), .ZN(n13867) );
  NAND2_X1 U7670 ( .A1(n2227), .A2(n2226), .ZN(n12128) );
  OAI211_X1 U7671 ( .C1(n10282), .C2(n10856), .A(n10281), .B(n10280), .ZN(
        n2227) );
  NAND3_X2 U7672 ( .A1(n20007), .A2(n5193), .A3(n20006), .ZN(n22006) );
  OAI22_X1 U7673 ( .A1(n4968), .A2(n3218), .B1(n17501), .B2(n24441), .ZN(n2229) );
  NAND2_X1 U7674 ( .A1(n10274), .A2(n10273), .ZN(n11492) );
  NAND2_X1 U7675 ( .A1(n17186), .A2(n17389), .ZN(n2230) );
  NAND3_X1 U7676 ( .A1(n2231), .A2(n18911), .A3(n1493), .ZN(n20127) );
  OAI21_X1 U7677 ( .B1(n19140), .B2(n19560), .A(n25448), .ZN(n2231) );
  XNOR2_X1 U7678 ( .A(n2232), .B(n23489), .ZN(Ciphertext[99]) );
  NAND2_X1 U7679 ( .A1(n23487), .A2(n23488), .ZN(n2232) );
  NAND2_X1 U7680 ( .A1(n12826), .A2(n12824), .ZN(n12828) );
  NAND2_X1 U7681 ( .A1(n2566), .A2(n16539), .ZN(n16540) );
  NOR2_X1 U7683 ( .A1(n5409), .A2(n16945), .ZN(n2233) );
  NAND2_X1 U7684 ( .A1(n6828), .A2(n6829), .ZN(n6830) );
  NAND2_X1 U7685 ( .A1(n18784), .A2(n18785), .ZN(n18786) );
  NAND2_X1 U7686 ( .A1(n2235), .A2(n6265), .ZN(n6270) );
  NAND2_X1 U7687 ( .A1(n6542), .A2(n7101), .ZN(n2235) );
  NAND2_X1 U7690 ( .A1(n2238), .A2(n23321), .ZN(n23323) );
  NAND2_X1 U7693 ( .A1(n6601), .A2(n5992), .ZN(n6099) );
  INV_X1 U7699 ( .A(n18749), .ZN(n3284) );
  NAND2_X1 U7700 ( .A1(n6949), .A2(n25437), .ZN(n5881) );
  OAI21_X1 U7701 ( .B1(n12834), .B2(n4389), .A(n13278), .ZN(n4388) );
  NAND3_X1 U7702 ( .A1(n4840), .A2(n17351), .A3(n17014), .ZN(n4888) );
  OAI21_X1 U7703 ( .B1(n10553), .B2(n1447), .A(n2592), .ZN(n2762) );
  XNOR2_X1 U7704 ( .A(n2242), .B(n15347), .ZN(n15349) );
  XNOR2_X1 U7705 ( .A(n25417), .B(n2242), .ZN(n14769) );
  XNOR2_X1 U7706 ( .A(n2242), .B(n15514), .ZN(n15517) );
  NOR2_X1 U7707 ( .A1(n2243), .A2(n10831), .ZN(n10832) );
  NAND2_X1 U7708 ( .A1(n10275), .A2(n2243), .ZN(n10515) );
  NAND2_X1 U7709 ( .A1(n4779), .A2(n2243), .ZN(n10276) );
  NAND2_X1 U7710 ( .A1(n10834), .A2(n2243), .ZN(n9647) );
  NOR2_X1 U7711 ( .A1(n10850), .A2(n10720), .ZN(n10722) );
  INV_X1 U7712 ( .A(n11123), .ZN(n2244) );
  OAI211_X1 U7713 ( .C1(n17134), .C2(n25245), .A(n25226), .B(n2245), .ZN(
        n16656) );
  NAND2_X1 U7714 ( .A1(n16655), .A2(n25245), .ZN(n2245) );
  NAND2_X1 U7716 ( .A1(n21035), .A2(n20101), .ZN(n2249) );
  OAI21_X1 U7720 ( .B1(n15588), .B2(n2253), .A(n15587), .ZN(n15589) );
  NAND3_X1 U7721 ( .A1(n2255), .A2(n2256), .A3(n2254), .ZN(n10623) );
  NAND3_X1 U7722 ( .A1(n10156), .A2(n2257), .A3(n9843), .ZN(n2255) );
  NAND2_X1 U7724 ( .A1(n19370), .A2(n24968), .ZN(n5461) );
  NAND2_X1 U7725 ( .A1(n16359), .A2(n24456), .ZN(n2259) );
  NAND2_X1 U7726 ( .A1(n2262), .A2(n7676), .ZN(n2261) );
  NAND3_X1 U7727 ( .A1(n2933), .A2(n17284), .A3(n2266), .ZN(n2265) );
  NAND2_X1 U7728 ( .A1(n16950), .A2(n17293), .ZN(n2266) );
  OR2_X1 U7729 ( .A1(n2266), .A2(n17289), .ZN(n2264) );
  INV_X1 U7730 ( .A(n9236), .ZN(n2267) );
  NAND2_X1 U7732 ( .A1(n9418), .A2(n9752), .ZN(n2269) );
  OAI21_X1 U7733 ( .B1(n454), .B2(n6588), .A(n7031), .ZN(n2270) );
  INV_X1 U7734 ( .A(n6588), .ZN(n7030) );
  XNOR2_X1 U7735 ( .A(n12240), .B(n2271), .ZN(n12245) );
  XNOR2_X1 U7736 ( .A(n11917), .B(n2271), .ZN(n11919) );
  XNOR2_X1 U7737 ( .A(n8721), .B(n729), .ZN(n3797) );
  XNOR2_X1 U7738 ( .A(n8721), .B(n2273), .ZN(n8036) );
  INV_X1 U7739 ( .A(n8721), .ZN(n2274) );
  NAND2_X1 U7740 ( .A1(n13466), .A2(n13744), .ZN(n3381) );
  XNOR2_X1 U7741 ( .A(n11433), .B(n12048), .ZN(n2277) );
  XNOR2_X1 U7742 ( .A(n2277), .B(n12342), .ZN(n12348) );
  INV_X1 U7743 ( .A(n2277), .ZN(n12341) );
  NAND3_X1 U7744 ( .A1(n6926), .A2(n1175), .A3(n6291), .ZN(n2279) );
  NAND2_X1 U7746 ( .A1(n16029), .A2(n16028), .ZN(n2280) );
  NAND2_X1 U7747 ( .A1(n14927), .A2(n2281), .ZN(n5336) );
  INV_X1 U7748 ( .A(n16274), .ZN(n2281) );
  NAND2_X1 U7749 ( .A1(n17467), .A2(n2064), .ZN(n2282) );
  INV_X1 U7750 ( .A(n18633), .ZN(n2283) );
  OR2_X1 U7751 ( .A1(n13349), .A2(n25366), .ZN(n2284) );
  AND2_X1 U7752 ( .A1(n14231), .A2(n14235), .ZN(n2977) );
  NAND3_X1 U7753 ( .A1(n17284), .A2(n2285), .A3(n17283), .ZN(n17285) );
  AOI21_X2 U7754 ( .B1(n16755), .B2(n2285), .A(n16544), .ZN(n17993) );
  INV_X1 U7755 ( .A(n2285), .ZN(n17287) );
  NAND2_X1 U7756 ( .A1(n17293), .A2(n2285), .ZN(n17231) );
  AND2_X1 U7757 ( .A1(n2285), .A2(n16950), .ZN(n4986) );
  NAND3_X1 U7758 ( .A1(n2287), .A2(n16927), .A3(n17321), .ZN(n3992) );
  NAND2_X1 U7759 ( .A1(n15671), .A2(n24890), .ZN(n2288) );
  NAND2_X1 U7760 ( .A1(n2289), .A2(n12791), .ZN(n2292) );
  INV_X1 U7761 ( .A(n12993), .ZN(n2289) );
  NAND2_X1 U7762 ( .A1(n2292), .A2(n2291), .ZN(n2290) );
  OR2_X1 U7763 ( .A1(n2294), .A2(n9872), .ZN(n2444) );
  NAND3_X1 U7764 ( .A1(n9872), .A2(n24549), .A3(n2294), .ZN(n9547) );
  NAND2_X1 U7765 ( .A1(n307), .A2(n2293), .ZN(n9253) );
  NAND2_X1 U7766 ( .A1(n13330), .A2(n2295), .ZN(n5313) );
  AOI21_X1 U7767 ( .B1(n13330), .B2(n25425), .A(n2295), .ZN(n12606) );
  NAND2_X1 U7768 ( .A1(n21077), .A2(n22180), .ZN(n2297) );
  NAND2_X1 U7769 ( .A1(n2298), .A2(n25012), .ZN(n4308) );
  NOR2_X1 U7770 ( .A1(n19241), .A2(n2298), .ZN(n18836) );
  OAI21_X1 U7771 ( .B1(n2328), .B2(n2298), .A(n278), .ZN(n3055) );
  OAI21_X1 U7772 ( .B1(n3919), .B2(n1806), .A(n2298), .ZN(n18884) );
  INV_X1 U7773 ( .A(n13450), .ZN(n14911) );
  XNOR2_X1 U7774 ( .A(n15093), .B(n2299), .ZN(n14392) );
  XNOR2_X1 U7775 ( .A(n13450), .B(n2300), .ZN(n2299) );
  INV_X1 U7776 ( .A(n14737), .ZN(n2300) );
  NAND2_X1 U7777 ( .A1(n13722), .A2(n13951), .ZN(n2302) );
  INV_X1 U7778 ( .A(n20184), .ZN(n20188) );
  NAND2_X1 U7779 ( .A1(n19862), .A2(n25211), .ZN(n20184) );
  INV_X1 U7780 ( .A(n2305), .ZN(n23665) );
  NOR2_X1 U7781 ( .A1(n24998), .A2(n23666), .ZN(n5506) );
  NOR2_X1 U7782 ( .A1(n23689), .A2(n24998), .ZN(n22186) );
  NOR2_X1 U7783 ( .A1(n23690), .A2(n24998), .ZN(n23691) );
  OAI21_X1 U7784 ( .B1(n23677), .B2(n24998), .A(n23676), .ZN(n23681) );
  NAND2_X1 U7785 ( .A1(n22747), .A2(n2305), .ZN(n23676) );
  NAND3_X1 U7786 ( .A1(n25405), .A2(n23678), .A3(n24998), .ZN(n22193) );
  NAND2_X1 U7788 ( .A1(n2306), .A2(n11005), .ZN(n10363) );
  NAND2_X1 U7789 ( .A1(n10365), .A2(n2306), .ZN(n10368) );
  INV_X1 U7790 ( .A(n10930), .ZN(n2309) );
  NAND2_X1 U7791 ( .A1(n5198), .A2(n10935), .ZN(n5296) );
  AND2_X1 U7792 ( .A1(n25018), .A2(n2312), .ZN(n21765) );
  NAND2_X1 U7793 ( .A1(n2315), .A2(n25018), .ZN(n2314) );
  NAND2_X1 U7795 ( .A1(n12893), .A2(n12894), .ZN(n2316) );
  NAND2_X1 U7796 ( .A1(n12895), .A2(n12896), .ZN(n2317) );
  NAND2_X1 U7797 ( .A1(n14685), .A2(n14686), .ZN(n2320) );
  XNOR2_X1 U7798 ( .A(n14493), .B(n2320), .ZN(n11682) );
  XNOR2_X1 U7799 ( .A(n24966), .B(n2318), .ZN(n3695) );
  INV_X1 U7800 ( .A(n3696), .ZN(n2318) );
  XNOR2_X1 U7801 ( .A(n24966), .B(n2319), .ZN(n14528) );
  AND2_X1 U7802 ( .A1(n13533), .A2(n2321), .ZN(n14017) );
  NAND4_X2 U7805 ( .A1(n7190), .A2(n7189), .A3(n7188), .A4(n2323), .ZN(n9059)
         );
  NAND2_X1 U7806 ( .A1(n17224), .A2(n25433), .ZN(n2325) );
  NAND2_X1 U7807 ( .A1(n22893), .A2(n22717), .ZN(n2327) );
  INV_X1 U7808 ( .A(n22836), .ZN(n22717) );
  NAND2_X1 U7809 ( .A1(n2330), .A2(n20571), .ZN(n20619) );
  NAND2_X1 U7810 ( .A1(n3795), .A2(n2330), .ZN(n3794) );
  XNOR2_X1 U7811 ( .A(n2331), .B(n2335), .ZN(n2333) );
  XNOR2_X1 U7812 ( .A(n17528), .B(n2334), .ZN(n2331) );
  XNOR2_X1 U7813 ( .A(n17963), .B(n17672), .ZN(n2332) );
  NAND2_X1 U7814 ( .A1(n2333), .A2(n19488), .ZN(n18727) );
  NAND2_X1 U7815 ( .A1(n16211), .A2(n24080), .ZN(n2336) );
  NAND2_X1 U7818 ( .A1(n5375), .A2(n2587), .ZN(n2338) );
  NAND2_X1 U7821 ( .A1(n2341), .A2(n23443), .ZN(n4309) );
  NAND2_X1 U7822 ( .A1(n2342), .A2(n22527), .ZN(n2341) );
  NAND2_X1 U7823 ( .A1(n24989), .A2(n1370), .ZN(n2342) );
  INV_X1 U7824 ( .A(n23441), .ZN(n22506) );
  INV_X1 U7826 ( .A(n19590), .ZN(n2346) );
  NAND2_X1 U7827 ( .A1(n18806), .A2(n2347), .ZN(n18091) );
  NAND2_X1 U7828 ( .A1(n5134), .A2(n24483), .ZN(n2347) );
  INV_X1 U7829 ( .A(n5964), .ZN(n2348) );
  NAND2_X1 U7830 ( .A1(n2353), .A2(n2354), .ZN(n2352) );
  NAND2_X1 U7831 ( .A1(n2355), .A2(n1175), .ZN(n2350) );
  NAND2_X1 U7832 ( .A1(n6480), .A2(n6775), .ZN(n2354) );
  NAND2_X1 U7833 ( .A1(n2357), .A2(n20099), .ZN(n2356) );
  NAND2_X1 U7834 ( .A1(n20104), .A2(n24378), .ZN(n2357) );
  NAND3_X1 U7835 ( .A1(n15941), .A2(n25389), .A3(n2359), .ZN(n15765) );
  AOI21_X1 U7836 ( .B1(n16254), .B2(n2359), .A(n16253), .ZN(n16255) );
  NAND3_X1 U7837 ( .A1(n277), .A2(n20374), .A3(n24558), .ZN(n20305) );
  NOR2_X1 U7839 ( .A1(n20591), .A2(n5093), .ZN(n2361) );
  NAND2_X1 U7840 ( .A1(n20589), .A2(n2361), .ZN(n2360) );
  NAND2_X1 U7841 ( .A1(n20591), .A2(n1424), .ZN(n2363) );
  NAND2_X1 U7843 ( .A1(n4719), .A2(n2364), .ZN(n4718) );
  NAND2_X1 U7844 ( .A1(n22497), .A2(n2364), .ZN(n4720) );
  OAI21_X1 U7847 ( .B1(n2368), .B2(n20092), .A(n2367), .ZN(n2365) );
  NAND2_X1 U7848 ( .A1(n2369), .A2(n2370), .ZN(n2366) );
  NAND2_X1 U7849 ( .A1(n1455), .A2(n20092), .ZN(n2367) );
  NAND2_X1 U7850 ( .A1(n20090), .A2(n20555), .ZN(n2371) );
  NAND3_X2 U7852 ( .A1(n15776), .A2(n4956), .A3(n15775), .ZN(n17078) );
  NAND2_X1 U7856 ( .A1(n18998), .A2(n24584), .ZN(n18586) );
  OAI21_X1 U7857 ( .B1(n16509), .B2(n25376), .A(n16508), .ZN(n4896) );
  OAI211_X1 U7858 ( .C1(n16509), .C2(n25376), .A(n16508), .B(n4899), .ZN(
        n16510) );
  NAND2_X1 U7859 ( .A1(n294), .A2(n25376), .ZN(n4899) );
  OAI21_X1 U7860 ( .B1(n25259), .B2(n15604), .A(n25376), .ZN(n15608) );
  NAND2_X1 U7861 ( .A1(n4300), .A2(n10094), .ZN(n8381) );
  NAND2_X1 U7862 ( .A1(n9327), .A2(n4300), .ZN(n5334) );
  NAND3_X1 U7863 ( .A1(n421), .A2(n10095), .A3(n4300), .ZN(n9516) );
  NOR2_X1 U7865 ( .A1(n24043), .A2(n25471), .ZN(n22591) );
  NAND2_X1 U7866 ( .A1(n22448), .A2(n24043), .ZN(n2395) );
  NAND3_X1 U7867 ( .A1(n22448), .A2(n274), .A3(n24043), .ZN(n2677) );
  NAND3_X1 U7869 ( .A1(n2378), .A2(n2380), .A3(n2377), .ZN(n2381) );
  NAND2_X1 U7870 ( .A1(n2379), .A2(n13549), .ZN(n2377) );
  NAND2_X1 U7871 ( .A1(n14204), .A2(n3341), .ZN(n2380) );
  OAI211_X1 U7872 ( .C1(n4145), .C2(n4144), .A(n2383), .B(n3352), .ZN(n8406)
         );
  NAND2_X1 U7873 ( .A1(n7477), .A2(n2384), .ZN(n2383) );
  INV_X1 U7874 ( .A(n7953), .ZN(n2384) );
  MUX2_X1 U7876 ( .A(n10754), .B(n10755), .S(n10759), .Z(n10761) );
  INV_X1 U7877 ( .A(n10885), .ZN(n2386) );
  NOR2_X1 U7878 ( .A1(n2388), .A2(n10302), .ZN(n2387) );
  NAND2_X1 U7879 ( .A1(n9477), .A2(n2389), .ZN(n9478) );
  INV_X1 U7880 ( .A(n10302), .ZN(n2389) );
  NAND2_X1 U7881 ( .A1(n9448), .A2(n24083), .ZN(n2390) );
  NAND2_X1 U7883 ( .A1(n9447), .A2(n24054), .ZN(n2392) );
  INV_X1 U7885 ( .A(n2397), .ZN(n21371) );
  AOI21_X1 U7886 ( .B1(n2397), .B2(n22792), .A(n22791), .ZN(n22794) );
  AND2_X1 U7887 ( .A1(n22617), .A2(n2397), .ZN(n22789) );
  NOR2_X1 U7888 ( .A1(n2397), .A2(n22617), .ZN(n22618) );
  MUX2_X1 U7890 ( .A(n22617), .B(n2397), .S(n22792), .Z(n22474) );
  NOR2_X1 U7892 ( .A1(n21371), .A2(n22790), .ZN(n2396) );
  NAND2_X1 U7893 ( .A1(n22612), .A2(n2397), .ZN(n4081) );
  NAND2_X1 U7894 ( .A1(n2398), .A2(n10169), .ZN(n2399) );
  NAND2_X1 U7895 ( .A1(n2207), .A2(n10166), .ZN(n2908) );
  MUX2_X1 U7896 ( .A(n9816), .B(n9815), .S(n2207), .Z(n9819) );
  NAND2_X1 U7898 ( .A1(n7747), .A2(n2402), .ZN(n3174) );
  AND2_X1 U7900 ( .A1(n2402), .A2(n7532), .ZN(n7277) );
  NAND3_X1 U7901 ( .A1(n3615), .A2(n2402), .A3(n8021), .ZN(n4706) );
  NAND2_X1 U7902 ( .A1(n433), .A2(n2404), .ZN(n4365) );
  OAI211_X1 U7903 ( .C1(n7697), .C2(n2404), .A(n7696), .B(n2403), .ZN(n7702)
         );
  NAND3_X1 U7904 ( .A1(n7695), .A2(n1490), .A3(n2404), .ZN(n2403) );
  MUX2_X1 U7905 ( .A(n2404), .B(n7699), .S(n7148), .Z(n7152) );
  NAND3_X1 U7906 ( .A1(n2404), .A2(n7148), .A3(n7217), .ZN(n8319) );
  XNOR2_X1 U7908 ( .A(n2405), .B(n11781), .ZN(n11786) );
  XNOR2_X1 U7909 ( .A(n11242), .B(n2406), .ZN(n2405) );
  INV_X1 U7910 ( .A(n12214), .ZN(n2406) );
  XNOR2_X1 U7911 ( .A(n15296), .B(n14961), .ZN(n2408) );
  NAND2_X1 U7912 ( .A1(n4433), .A2(n2409), .ZN(n4431) );
  INV_X1 U7913 ( .A(n19522), .ZN(n2409) );
  NAND2_X1 U7914 ( .A1(n2410), .A2(n19371), .ZN(n5441) );
  OAI21_X1 U7915 ( .B1(n19223), .B2(n2410), .A(n19222), .ZN(n19224) );
  OAI22_X1 U7917 ( .A1(n23787), .A2(n2590), .B1(n2591), .B2(n2411), .ZN(n2589)
         );
  AND2_X1 U7918 ( .A1(n23786), .A2(n3201), .ZN(n2411) );
  NAND2_X1 U7919 ( .A1(n2412), .A2(n15198), .ZN(n15767) );
  NAND2_X1 U7920 ( .A1(n16010), .A2(n2173), .ZN(n15751) );
  INV_X1 U7921 ( .A(n15556), .ZN(n2412) );
  NAND2_X1 U7922 ( .A1(n2413), .A2(n24085), .ZN(n3029) );
  NAND2_X1 U7923 ( .A1(n24802), .A2(n19480), .ZN(n17894) );
  XNOR2_X1 U7925 ( .A(n21342), .B(n21345), .ZN(n2416) );
  NAND2_X1 U7926 ( .A1(n2419), .A2(n2418), .ZN(n17437) );
  NAND3_X1 U7927 ( .A1(n2420), .A2(n25502), .A3(n15973), .ZN(n2418) );
  NOR3_X1 U7928 ( .A1(n21863), .A2(n23892), .A3(n23893), .ZN(n23894) );
  OR2_X2 U7929 ( .A1(n23891), .A2(n2421), .ZN(n21863) );
  OAI22_X1 U7930 ( .A1(n22772), .A2(n22370), .B1(n22682), .B2(n22679), .ZN(
        n2421) );
  OAI211_X1 U7931 ( .C1(n25415), .C2(n398), .A(n2422), .B(n5412), .ZN(n2424)
         );
  NAND2_X1 U7932 ( .A1(n12861), .A2(n12636), .ZN(n4729) );
  NAND2_X1 U7933 ( .A1(n20460), .A2(n24460), .ZN(n20165) );
  NAND2_X1 U7935 ( .A1(n20385), .A2(n20395), .ZN(n2427) );
  NAND2_X1 U7937 ( .A1(n11302), .A2(n11297), .ZN(n10434) );
  NAND2_X1 U7938 ( .A1(n17479), .A2(n17478), .ZN(n2429) );
  INV_X1 U7939 ( .A(n17078), .ZN(n17479) );
  NAND2_X1 U7940 ( .A1(n2430), .A2(n17160), .ZN(n5225) );
  NAND2_X1 U7941 ( .A1(n10538), .A2(n10885), .ZN(n2435) );
  NAND2_X1 U7942 ( .A1(n10541), .A2(n2388), .ZN(n10544) );
  NAND2_X1 U7943 ( .A1(n10888), .A2(n2388), .ZN(n3417) );
  INV_X1 U7944 ( .A(n11722), .ZN(n12915) );
  NAND3_X1 U7945 ( .A1(n2437), .A2(n13304), .A3(n13307), .ZN(n2436) );
  NAND2_X1 U7946 ( .A1(n12904), .A2(n12915), .ZN(n2438) );
  INV_X1 U7947 ( .A(n9872), .ZN(n9251) );
  XNOR2_X2 U7948 ( .A(n8083), .B(n8082), .ZN(n9872) );
  NAND3_X1 U7949 ( .A1(n2445), .A2(n2444), .A3(n2440), .ZN(n10924) );
  NAND3_X1 U7950 ( .A1(n2442), .A2(n2441), .A3(n307), .ZN(n2440) );
  NAND2_X1 U7951 ( .A1(n2443), .A2(n9694), .ZN(n2441) );
  NAND2_X1 U7952 ( .A1(n9872), .A2(n9692), .ZN(n2442) );
  NAND3_X1 U7953 ( .A1(n9027), .A2(n9872), .A3(n2443), .ZN(n2445) );
  INV_X1 U7954 ( .A(n9692), .ZN(n2443) );
  XNOR2_X1 U7955 ( .A(n8862), .B(n8086), .ZN(n2446) );
  NAND3_X1 U7956 ( .A1(n6143), .A2(n2447), .A3(n7615), .ZN(n6151) );
  AND2_X1 U7957 ( .A1(n2448), .A2(n6142), .ZN(n2447) );
  OAI21_X1 U7958 ( .B1(n10658), .B2(n10398), .A(n2450), .ZN(n2449) );
  NAND2_X1 U7959 ( .A1(n25250), .A2(n10660), .ZN(n10658) );
  AND2_X1 U7961 ( .A1(n355), .A2(n19613), .ZN(n18837) );
  XNOR2_X1 U7962 ( .A(n18666), .B(n18491), .ZN(n18538) );
  NOR2_X2 U7963 ( .A1(n2451), .A2(n17367), .ZN(n18491) );
  NAND2_X1 U7964 ( .A1(n2452), .A2(n2453), .ZN(n2451) );
  NAND2_X1 U7966 ( .A1(n17365), .A2(n24569), .ZN(n2453) );
  NAND3_X2 U7970 ( .A1(n1390), .A2(n2887), .A3(n2456), .ZN(n23592) );
  AND2_X1 U7971 ( .A1(n24974), .A2(n14289), .ZN(n2457) );
  NAND3_X1 U7972 ( .A1(n24974), .A2(n14289), .A3(n13909), .ZN(n3069) );
  OAI21_X1 U7973 ( .B1(n13948), .B2(n2457), .A(n391), .ZN(n13910) );
  OAI21_X2 U7974 ( .B1(n5622), .B2(n7911), .A(n2458), .ZN(n9034) );
  OAI21_X1 U7975 ( .B1(n7628), .B2(n7909), .A(n2460), .ZN(n2459) );
  INV_X1 U7976 ( .A(n7155), .ZN(n2461) );
  NAND2_X1 U7978 ( .A1(n19107), .A2(n2464), .ZN(n19584) );
  NAND2_X1 U7979 ( .A1(n18445), .A2(n19875), .ZN(n2466) );
  NAND2_X1 U7980 ( .A1(n18444), .A2(n20023), .ZN(n2467) );
  NAND2_X1 U7982 ( .A1(n5051), .A2(n2471), .ZN(n3083) );
  NOR2_X1 U7983 ( .A1(n311), .A2(n7604), .ZN(n2471) );
  INV_X1 U7984 ( .A(n12955), .ZN(n2472) );
  NOR2_X1 U7985 ( .A1(n23805), .A2(n2477), .ZN(n2476) );
  NAND3_X1 U7986 ( .A1(n4533), .A2(n21837), .A3(n2474), .ZN(n2473) );
  AND2_X1 U7987 ( .A1(n24983), .A2(n21903), .ZN(n2474) );
  NAND2_X1 U7989 ( .A1(n21837), .A2(n23002), .ZN(n23787) );
  NOR2_X1 U7990 ( .A1(n25030), .A2(n16106), .ZN(n4675) );
  NAND2_X1 U7991 ( .A1(n24928), .A2(n16107), .ZN(n2479) );
  NAND2_X1 U7992 ( .A1(n16109), .A2(n16108), .ZN(n2480) );
  NAND2_X1 U7993 ( .A1(n2484), .A2(n2482), .ZN(n2481) );
  NAND2_X1 U7994 ( .A1(n25430), .A2(n2483), .ZN(n2482) );
  NOR2_X1 U7995 ( .A1(n12349), .A2(n13350), .ZN(n2483) );
  INV_X1 U7996 ( .A(n13123), .ZN(n5624) );
  INV_X1 U7997 ( .A(n25430), .ZN(n2485) );
  NAND2_X1 U7998 ( .A1(n4256), .A2(n9507), .ZN(n2486) );
  NAND2_X1 U7999 ( .A1(n21954), .A2(n24911), .ZN(n2488) );
  OAI22_X1 U8000 ( .A1(n4171), .A2(n23370), .B1(n22430), .B2(n24404), .ZN(
        n2487) );
  AOI21_X1 U8001 ( .B1(n4606), .B2(n2488), .A(n2487), .ZN(n2489) );
  XNOR2_X1 U8002 ( .A(n2489), .B(n21711), .ZN(Ciphertext[77]) );
  XNOR2_X1 U8003 ( .A(n2491), .B(n24413), .ZN(n8445) );
  NAND2_X1 U8004 ( .A1(n7223), .A2(n7952), .ZN(n2490) );
  NAND3_X1 U8005 ( .A1(n7953), .A2(n7952), .A3(n4144), .ZN(n2880) );
  OAI21_X1 U8006 ( .B1(n12767), .B2(n13216), .A(n2492), .ZN(n12811) );
  NAND2_X1 U8007 ( .A1(n24513), .A2(n13216), .ZN(n2492) );
  NAND3_X1 U8008 ( .A1(n12987), .A2(n12986), .A3(n2493), .ZN(n12988) );
  NAND2_X1 U8009 ( .A1(n6752), .A2(n6675), .ZN(n2494) );
  NAND2_X1 U8010 ( .A1(n2497), .A2(n2501), .ZN(n5101) );
  NAND2_X1 U8011 ( .A1(n2498), .A2(n2499), .ZN(n2497) );
  NAND2_X1 U8012 ( .A1(n2500), .A2(n2499), .ZN(n10838) );
  NAND2_X1 U8013 ( .A1(n9298), .A2(n9676), .ZN(n2499) );
  NAND2_X1 U8014 ( .A1(n2501), .A2(n5448), .ZN(n2500) );
  NAND3_X1 U8015 ( .A1(n298), .A2(n14327), .A3(n5230), .ZN(n2502) );
  NAND2_X1 U8016 ( .A1(n14325), .A2(n2505), .ZN(n2504) );
  INV_X1 U8017 ( .A(n13590), .ZN(n2506) );
  NAND2_X1 U8018 ( .A1(n2587), .A2(n4760), .ZN(n2509) );
  NAND2_X1 U8019 ( .A1(n2511), .A2(n17274), .ZN(n2510) );
  OR2_X1 U8021 ( .A1(n3888), .A2(n14944), .ZN(n2514) );
  NAND2_X1 U8023 ( .A1(n12621), .A2(n12622), .ZN(n2517) );
  NOR2_X2 U8024 ( .A1(n12628), .A2(n12627), .ZN(n14944) );
  NAND2_X1 U8025 ( .A1(n15857), .A2(n2518), .ZN(n15805) );
  NAND2_X1 U8026 ( .A1(n16116), .A2(n15857), .ZN(n5176) );
  NAND2_X1 U8028 ( .A1(n2520), .A2(n7757), .ZN(n2521) );
  NAND2_X1 U8029 ( .A1(n23285), .A2(n23292), .ZN(n22508) );
  NAND3_X1 U8030 ( .A1(n10698), .A2(n10952), .A3(n25232), .ZN(n2523) );
  NAND3_X1 U8031 ( .A1(n10951), .A2(n25232), .A3(n10548), .ZN(n2524) );
  NAND2_X1 U8032 ( .A1(n25038), .A2(n17330), .ZN(n17331) );
  NAND2_X1 U8033 ( .A1(n12916), .A2(n2526), .ZN(n3493) );
  NAND2_X1 U8034 ( .A1(n13311), .A2(n11722), .ZN(n2526) );
  OR2_X1 U8035 ( .A1(n13305), .A2(n12613), .ZN(n13311) );
  NAND3_X1 U8037 ( .A1(n2531), .A2(n6266), .A3(n7101), .ZN(n2533) );
  INV_X1 U8038 ( .A(n7098), .ZN(n2531) );
  NAND2_X1 U8039 ( .A1(n5916), .A2(n7103), .ZN(n2532) );
  NAND2_X1 U8040 ( .A1(n6267), .A2(n6165), .ZN(n6265) );
  NAND2_X1 U8041 ( .A1(n2536), .A2(n3181), .ZN(n2535) );
  NAND2_X1 U8042 ( .A1(n2537), .A2(n23478), .ZN(n2536) );
  NOR2_X1 U8043 ( .A1(n23479), .A2(n23499), .ZN(n2537) );
  INV_X1 U8045 ( .A(n2540), .ZN(n19211) );
  NAND2_X1 U8046 ( .A1(n24447), .A2(n19359), .ZN(n4315) );
  NAND2_X1 U8047 ( .A1(n19210), .A2(n24447), .ZN(n19215) );
  AOI22_X1 U8048 ( .A1(n3943), .A2(n4135), .B1(n18021), .B2(n24447), .ZN(
        n19878) );
  OAI21_X1 U8049 ( .B1(n6329), .B2(n6425), .A(n2542), .ZN(n6330) );
  NAND2_X1 U8051 ( .A1(n14036), .A2(n14035), .ZN(n3893) );
  NAND2_X1 U8052 ( .A1(n10971), .A2(n2546), .ZN(n10816) );
  AND2_X2 U8053 ( .A1(n3597), .A2(n3596), .ZN(n2546) );
  NAND2_X1 U8054 ( .A1(n2546), .A2(n10969), .ZN(n10495) );
  NAND2_X1 U8055 ( .A1(n10815), .A2(n2546), .ZN(n3595) );
  XNOR2_X1 U8056 ( .A(n25483), .B(n21478), .ZN(n21479) );
  INV_X1 U8059 ( .A(n17438), .ZN(n2549) );
  OAI21_X1 U8060 ( .B1(n17442), .B2(n17441), .A(n2550), .ZN(n16829) );
  NAND2_X1 U8062 ( .A1(n18808), .A2(n19590), .ZN(n19252) );
  NAND2_X1 U8064 ( .A1(n4286), .A2(n369), .ZN(n15609) );
  NOR2_X1 U8065 ( .A1(n7609), .A2(n7604), .ZN(n7608) );
  NAND2_X1 U8066 ( .A1(n7890), .A2(n7323), .ZN(n6010) );
  NAND2_X1 U8067 ( .A1(n7890), .A2(n2552), .ZN(n2551) );
  NAND2_X1 U8068 ( .A1(n7608), .A2(n7893), .ZN(n2553) );
  NAND2_X1 U8070 ( .A1(n7322), .A2(n7605), .ZN(n2555) );
  NAND3_X1 U8071 ( .A1(n4293), .A2(n13963), .A3(n13968), .ZN(n2557) );
  INV_X1 U8072 ( .A(n14732), .ZN(n15285) );
  NAND3_X1 U8073 ( .A1(n2558), .A2(n2556), .A3(n2557), .ZN(n14732) );
  NAND3_X1 U8074 ( .A1(n2559), .A2(n1771), .A3(n4305), .ZN(n2558) );
  OR2_X1 U8075 ( .A1(n13883), .A2(n11806), .ZN(n2559) );
  NAND3_X1 U8076 ( .A1(n13968), .A2(n13724), .A3(n13969), .ZN(n2556) );
  NAND2_X1 U8077 ( .A1(n11805), .A2(n13724), .ZN(n13964) );
  NAND2_X1 U8078 ( .A1(n2558), .A2(n2557), .ZN(n14397) );
  XNOR2_X1 U8079 ( .A(n8450), .B(n2560), .ZN(n8252) );
  XNOR2_X1 U8080 ( .A(n2560), .B(n8517), .ZN(n8292) );
  INV_X2 U8081 ( .A(n2562), .ZN(n17633) );
  INV_X1 U8082 ( .A(n24959), .ZN(n9372) );
  AOI21_X1 U8083 ( .B1(n10252), .B2(n9378), .A(n9211), .ZN(n2564) );
  INV_X1 U8084 ( .A(n3472), .ZN(n2565) );
  NAND3_X1 U8085 ( .A1(n17633), .A2(n16902), .A3(n2566), .ZN(n16903) );
  OR2_X1 U8086 ( .A1(n46), .A2(n2566), .ZN(n17632) );
  NAND2_X1 U8087 ( .A1(n19742), .A2(n20255), .ZN(n2567) );
  XNOR2_X1 U8088 ( .A(n2569), .B(n21084), .ZN(n20223) );
  XNOR2_X1 U8089 ( .A(n2569), .B(n21985), .ZN(n21987) );
  XNOR2_X1 U8090 ( .A(n2569), .B(n21622), .ZN(n19748) );
  XNOR2_X1 U8091 ( .A(n20815), .B(n2569), .ZN(n20817) );
  INV_X1 U8093 ( .A(n3888), .ZN(n14199) );
  INV_X1 U8094 ( .A(n14949), .ZN(n14950) );
  NAND2_X1 U8095 ( .A1(n2684), .A2(n14202), .ZN(n14949) );
  INV_X1 U8096 ( .A(n14945), .ZN(n2570) );
  NAND2_X1 U8098 ( .A1(n12660), .A2(n12272), .ZN(n2571) );
  INV_X1 U8099 ( .A(n2572), .ZN(n4921) );
  NAND2_X1 U8100 ( .A1(n13460), .A2(n13900), .ZN(n2572) );
  OAI21_X1 U8101 ( .B1(n13733), .B2(n13460), .A(n2572), .ZN(n12428) );
  NAND2_X1 U8102 ( .A1(n12499), .A2(n25033), .ZN(n2574) );
  NAND2_X1 U8103 ( .A1(n12500), .A2(n10711), .ZN(n2575) );
  AND2_X1 U8104 ( .A1(n439), .A2(n6996), .ZN(n6811) );
  NAND2_X1 U8105 ( .A1(n2576), .A2(n6658), .ZN(n4149) );
  NAND3_X1 U8106 ( .A1(n2576), .A2(n6367), .A3(n6999), .ZN(n7000) );
  NAND3_X1 U8107 ( .A1(n2576), .A2(n6658), .A3(n6367), .ZN(n6074) );
  NAND2_X1 U8108 ( .A1(n6997), .A2(n2576), .ZN(n5818) );
  INV_X1 U8109 ( .A(n6996), .ZN(n2576) );
  AOI21_X1 U8110 ( .B1(n22364), .B2(n22365), .A(n22675), .ZN(n22368) );
  XNOR2_X1 U8111 ( .A(n4978), .B(n21134), .ZN(n2577) );
  INV_X1 U8112 ( .A(n18582), .ZN(n17643) );
  INV_X1 U8116 ( .A(n17115), .ZN(n2581) );
  OAI22_X1 U8117 ( .A1(n10509), .A2(n2311), .B1(n10936), .B2(n2584), .ZN(
        n10510) );
  NAND2_X1 U8118 ( .A1(n10931), .A2(n10935), .ZN(n2584) );
  NAND2_X1 U8119 ( .A1(n10128), .A2(n2585), .ZN(n10127) );
  NAND2_X1 U8120 ( .A1(n5057), .A2(n24959), .ZN(n9212) );
  NAND2_X1 U8121 ( .A1(n10132), .A2(n24959), .ZN(n9377) );
  NAND2_X1 U8122 ( .A1(n7438), .A2(n24959), .ZN(n7439) );
  MUX2_X1 U8123 ( .A(n10251), .B(n10252), .S(n9372), .Z(n10253) );
  AND2_X1 U8125 ( .A1(n16796), .A2(n2587), .ZN(n5762) );
  NAND2_X1 U8126 ( .A1(n2586), .A2(n5375), .ZN(n16797) );
  AND2_X1 U8127 ( .A1(n2587), .A2(n16795), .ZN(n2586) );
  MUX2_X1 U8128 ( .A(n16795), .B(n2587), .S(n16796), .Z(n15737) );
  NAND2_X1 U8129 ( .A1(n5376), .A2(n2587), .ZN(n2728) );
  NAND2_X1 U8130 ( .A1(n16794), .A2(n2587), .ZN(n5242) );
  INV_X1 U8131 ( .A(n22043), .ZN(n23790) );
  XNOR2_X1 U8132 ( .A(n2589), .B(n2588), .ZN(Ciphertext[151]) );
  INV_X1 U8133 ( .A(n10985), .ZN(n2592) );
  AND2_X1 U8134 ( .A1(n6713), .A2(n2593), .ZN(n6717) );
  NAND2_X1 U8135 ( .A1(n24050), .A2(n6235), .ZN(n2593) );
  INV_X1 U8136 ( .A(n3480), .ZN(n2594) );
  AOI21_X1 U8137 ( .B1(n20555), .B2(n2594), .A(n20330), .ZN(n3478) );
  NAND2_X1 U8138 ( .A1(n20331), .A2(n2594), .ZN(n20332) );
  NAND2_X1 U8139 ( .A1(n2596), .A2(n330), .ZN(n2595) );
  NAND2_X1 U8140 ( .A1(n22677), .A2(n23997), .ZN(n2597) );
  NAND2_X1 U8141 ( .A1(n6971), .A2(n6690), .ZN(n2600) );
  NAND2_X1 U8144 ( .A1(n6974), .A2(n2600), .ZN(n4544) );
  XNOR2_X2 U8145 ( .A(n20855), .B(n20854), .ZN(n2601) );
  NAND2_X1 U8146 ( .A1(n22175), .A2(n2601), .ZN(n22198) );
  NOR2_X1 U8147 ( .A1(n23571), .A2(n2601), .ZN(n23572) );
  MUX2_X1 U8148 ( .A(n2601), .B(n23576), .S(n22175), .Z(n22080) );
  NAND2_X1 U8149 ( .A1(n22174), .A2(n2601), .ZN(n22178) );
  OAI22_X1 U8150 ( .A1(n4360), .A2(n2601), .B1(n24369), .B2(n1323), .ZN(n23577) );
  OAI22_X1 U8151 ( .A1(n21760), .A2(n2601), .B1(n23574), .B2(n22201), .ZN(
        n21761) );
  XNOR2_X1 U8152 ( .A(n2602), .B(n2222), .ZN(n11813) );
  XNOR2_X1 U8153 ( .A(n12096), .B(n2602), .ZN(n12098) );
  XNOR2_X1 U8154 ( .A(n12381), .B(n2602), .ZN(n11999) );
  XNOR2_X1 U8155 ( .A(n12241), .B(n2602), .ZN(n11432) );
  INV_X1 U8156 ( .A(n2603), .ZN(n13587) );
  NAND2_X1 U8157 ( .A1(n2629), .A2(n2603), .ZN(n13570) );
  NAND2_X1 U8160 ( .A1(n2607), .A2(n15564), .ZN(n15565) );
  NOR2_X1 U8161 ( .A1(n15933), .A2(n24387), .ZN(n15932) );
  NAND2_X1 U8162 ( .A1(n387), .A2(n24387), .ZN(n3712) );
  NAND2_X1 U8163 ( .A1(n5097), .A2(n24387), .ZN(n5096) );
  AOI21_X1 U8164 ( .B1(n387), .B2(n16232), .A(n24387), .ZN(n5024) );
  OAI21_X1 U8165 ( .B1(n387), .B2(n2607), .A(n16491), .ZN(n16493) );
  OAI211_X1 U8166 ( .C1(n24750), .C2(n25049), .A(n4587), .B(n2608), .ZN(n12999) );
  NAND2_X1 U8167 ( .A1(n25049), .A2(n12993), .ZN(n2608) );
  OAI21_X1 U8168 ( .B1(n15742), .B2(n16193), .A(n2610), .ZN(n15259) );
  NOR2_X1 U8169 ( .A1(n16324), .A2(n25447), .ZN(n15675) );
  NAND3_X1 U8170 ( .A1(n16328), .A2(n16323), .A3(n2610), .ZN(n15900) );
  MUX2_X1 U8172 ( .A(n25447), .B(n16323), .S(n16324), .Z(n16330) );
  INV_X1 U8173 ( .A(n8874), .ZN(n2612) );
  XNOR2_X1 U8174 ( .A(n2611), .B(n8874), .ZN(n8301) );
  INV_X1 U8175 ( .A(n8457), .ZN(n2611) );
  XNOR2_X1 U8176 ( .A(n2612), .B(n8897), .ZN(n8622) );
  NAND2_X1 U8177 ( .A1(n372), .A2(n17053), .ZN(n2615) );
  NAND3_X1 U8178 ( .A1(n372), .A2(n17053), .A3(n2613), .ZN(n2614) );
  NAND2_X1 U8179 ( .A1(n2615), .A2(n17051), .ZN(n3435) );
  NAND2_X1 U8180 ( .A1(n330), .A2(n23998), .ZN(n22376) );
  OR2_X1 U8181 ( .A1(n2616), .A2(n24439), .ZN(n24002) );
  NAND2_X1 U8182 ( .A1(n330), .A2(n25439), .ZN(n2617) );
  INV_X1 U8184 ( .A(n2621), .ZN(n7791) );
  OR2_X1 U8185 ( .A1(n2620), .A2(n7781), .ZN(n2621) );
  INV_X1 U8186 ( .A(n7788), .ZN(n2620) );
  NAND2_X1 U8187 ( .A1(n7441), .A2(n2621), .ZN(n7443) );
  NAND2_X1 U8188 ( .A1(n21762), .A2(n22929), .ZN(n5687) );
  NOR2_X1 U8189 ( .A1(n22188), .A2(n22715), .ZN(n21762) );
  NAND2_X1 U8190 ( .A1(n8011), .A2(n8015), .ZN(n2622) );
  INV_X1 U8191 ( .A(n8011), .ZN(n2623) );
  NAND2_X1 U8192 ( .A1(n8012), .A2(n2624), .ZN(n6207) );
  NOR2_X1 U8193 ( .A1(n2624), .A2(n7537), .ZN(n7293) );
  NAND3_X1 U8194 ( .A1(n2640), .A2(n2624), .A3(n7537), .ZN(n7538) );
  NAND2_X1 U8195 ( .A1(n8013), .A2(n2624), .ZN(n3236) );
  MUX2_X1 U8196 ( .A(n8016), .B(n8013), .S(n2624), .Z(n3238) );
  NOR2_X1 U8197 ( .A1(n20258), .A2(n5569), .ZN(n2625) );
  NAND2_X1 U8198 ( .A1(n2627), .A2(n25054), .ZN(n5570) );
  OAI21_X1 U8199 ( .B1(n5572), .B2(n19125), .A(n5571), .ZN(n2627) );
  AND2_X1 U8200 ( .A1(n15706), .A2(n16048), .ZN(n15539) );
  NAND2_X1 U8201 ( .A1(n11205), .A2(n11338), .ZN(n2628) );
  NAND2_X1 U8202 ( .A1(n2629), .A2(n14361), .ZN(n13572) );
  NOR2_X1 U8203 ( .A1(n2629), .A2(n14361), .ZN(n14363) );
  NAND2_X1 U8204 ( .A1(n13397), .A2(n1486), .ZN(n15019) );
  NAND2_X1 U8205 ( .A1(n24426), .A2(n23406), .ZN(n2630) );
  NOR2_X1 U8206 ( .A1(n24074), .A2(n23420), .ZN(n23406) );
  NOR2_X1 U8209 ( .A1(n24877), .A2(n23461), .ZN(n22491) );
  XNOR2_X1 U8210 ( .A(n21725), .B(n21722), .ZN(n2634) );
  NAND2_X1 U8211 ( .A1(n16441), .A2(n24293), .ZN(n2635) );
  INV_X1 U8212 ( .A(n16440), .ZN(n2636) );
  NAND2_X1 U8214 ( .A1(n12536), .A2(n13757), .ZN(n13837) );
  NAND3_X1 U8215 ( .A1(n25451), .A2(n8014), .A3(n2640), .ZN(n7299) );
  NAND2_X1 U8216 ( .A1(n7293), .A2(n2640), .ZN(n6214) );
  NAND3_X1 U8217 ( .A1(n8016), .A2(n8015), .A3(n2640), .ZN(n8017) );
  NAND2_X1 U8218 ( .A1(n8011), .A2(n2640), .ZN(n8020) );
  AOI21_X1 U8219 ( .B1(n7296), .B2(n7297), .A(n2640), .ZN(n7301) );
  NAND2_X1 U8221 ( .A1(n17411), .A2(n17612), .ZN(n2641) );
  NAND2_X1 U8222 ( .A1(n2645), .A2(n19233), .ZN(n2642) );
  INV_X1 U8224 ( .A(n19607), .ZN(n2644) );
  INV_X1 U8225 ( .A(n19608), .ZN(n2645) );
  NAND2_X1 U8227 ( .A1(n6838), .A2(n6991), .ZN(n2646) );
  NAND2_X1 U8228 ( .A1(n6841), .A2(n6640), .ZN(n6639) );
  NAND2_X1 U8231 ( .A1(n15574), .A2(n16273), .ZN(n2649) );
  NAND3_X1 U8232 ( .A1(n2281), .A2(n16030), .A3(n16029), .ZN(n2650) );
  NAND2_X2 U8233 ( .A1(n14786), .A2(n3067), .ZN(n17410) );
  MUX2_X1 U8234 ( .A(n17613), .B(n16743), .S(n17407), .Z(n2652) );
  INV_X1 U8235 ( .A(n17607), .ZN(n17613) );
  NAND2_X1 U8236 ( .A1(n17609), .A2(n17608), .ZN(n2653) );
  NAND3_X1 U8243 ( .A1(n24876), .A2(n24507), .A3(n24589), .ZN(n2657) );
  NAND3_X1 U8245 ( .A1(n5509), .A2(n5511), .A3(n2659), .ZN(n17515) );
  NAND2_X1 U8246 ( .A1(n16878), .A2(n17015), .ZN(n2659) );
  INV_X1 U8247 ( .A(n22901), .ZN(n5463) );
  AOI21_X1 U8249 ( .B1(n2711), .B2(n1431), .A(n2661), .ZN(n2660) );
  INV_X1 U8250 ( .A(n22848), .ZN(n2661) );
  NAND2_X1 U8251 ( .A1(n22904), .A2(n22842), .ZN(n22848) );
  INV_X1 U8253 ( .A(n19762), .ZN(n19427) );
  NOR2_X2 U8254 ( .A1(n19761), .A2(n2662), .ZN(n19953) );
  INV_X1 U8256 ( .A(n18385), .ZN(n19183) );
  NAND2_X1 U8258 ( .A1(n16724), .A2(n5484), .ZN(n2664) );
  NAND2_X1 U8259 ( .A1(n16723), .A2(n5484), .ZN(n2665) );
  OR2_X1 U8260 ( .A1(n16723), .A2(n5484), .ZN(n2666) );
  XNOR2_X1 U8261 ( .A(n18456), .B(n2667), .ZN(n18457) );
  XNOR2_X1 U8262 ( .A(n2667), .B(n18637), .ZN(n18226) );
  XNOR2_X1 U8263 ( .A(n2667), .B(n17663), .ZN(n17533) );
  XNOR2_X1 U8264 ( .A(n2667), .B(n18291), .ZN(n17804) );
  NAND2_X1 U8266 ( .A1(n2670), .A2(n23318), .ZN(n2669) );
  NAND2_X1 U8267 ( .A1(n3564), .A2(n24316), .ZN(n2670) );
  XNOR2_X2 U8270 ( .A(n21529), .B(n21528), .ZN(n2674) );
  NAND2_X1 U8271 ( .A1(n22421), .A2(n2674), .ZN(n21547) );
  NAND2_X1 U8272 ( .A1(n22422), .A2(n2674), .ZN(n21548) );
  NOR2_X1 U8274 ( .A1(n21530), .A2(n2674), .ZN(n21531) );
  INV_X1 U8277 ( .A(n10416), .ZN(n2680) );
  NAND2_X1 U8278 ( .A1(n11012), .A2(n4531), .ZN(n11010) );
  NAND2_X1 U8279 ( .A1(n4530), .A2(n2681), .ZN(n10353) );
  NAND3_X1 U8280 ( .A1(n11045), .A2(n2680), .A3(n2681), .ZN(n11049) );
  NAND2_X1 U8282 ( .A1(n2683), .A2(n14945), .ZN(n2682) );
  INV_X1 U8286 ( .A(n17192), .ZN(n17028) );
  NAND2_X1 U8287 ( .A1(n2689), .A2(n17399), .ZN(n17401) );
  NAND2_X1 U8288 ( .A1(n17398), .A2(n285), .ZN(n2689) );
  AOI22_X1 U8289 ( .A1(n3176), .A2(n23460), .B1(n2691), .B2(n23461), .ZN(n2690) );
  NAND2_X1 U8290 ( .A1(n21797), .A2(n21796), .ZN(n4000) );
  OAI211_X2 U8291 ( .C1(n24570), .C2(n4299), .A(n16776), .B(n4297), .ZN(n18660) );
  NAND4_X2 U8292 ( .A1(n19247), .A2(n2694), .A3(n2693), .A4(n19246), .ZN(
        n20599) );
  NAND2_X1 U8293 ( .A1(n2695), .A2(n19245), .ZN(n2694) );
  NAND2_X1 U8294 ( .A1(n20027), .A2(n20343), .ZN(n2696) );
  NAND2_X1 U8295 ( .A1(n19645), .A2(n20279), .ZN(n2697) );
  NAND2_X1 U8296 ( .A1(n2699), .A2(n20277), .ZN(n2698) );
  AND2_X1 U8297 ( .A1(n20346), .A2(n19809), .ZN(n20027) );
  INV_X1 U8299 ( .A(n19809), .ZN(n20280) );
  NAND2_X1 U8300 ( .A1(n2702), .A2(n2703), .ZN(n2701) );
  NAND2_X1 U8301 ( .A1(n16283), .A2(n1654), .ZN(n2703) );
  XNOR2_X1 U8302 ( .A(n17592), .B(n16574), .ZN(n2704) );
  INV_X1 U8303 ( .A(n17592), .ZN(n18374) );
  XNOR2_X1 U8304 ( .A(n18284), .B(n2704), .ZN(n16582) );
  OAI21_X1 U8307 ( .B1(n16185), .B2(n16337), .A(n16184), .ZN(n16871) );
  MUX2_X1 U8308 ( .A(n17179), .B(n3602), .S(n17389), .Z(n17190) );
  NAND3_X1 U8311 ( .A1(n25382), .A2(n22900), .A3(n25569), .ZN(n2708) );
  OAI21_X2 U8312 ( .B1(n2709), .B2(n23020), .A(n22735), .ZN(n23480) );
  NAND2_X1 U8315 ( .A1(n22896), .A2(n22835), .ZN(n2713) );
  NOR2_X1 U8316 ( .A1(n4737), .A2(n11163), .ZN(n2714) );
  NAND3_X1 U8317 ( .A1(n10053), .A2(n9244), .A3(n4096), .ZN(n3049) );
  AOI22_X2 U8319 ( .A1(n10437), .A2(n11092), .B1(n10436), .B2(n11300), .ZN(
        n11646) );
  INV_X1 U8320 ( .A(n3698), .ZN(n5526) );
  NOR2_X1 U8321 ( .A1(n17031), .A2(n4039), .ZN(n4038) );
  OR2_X1 U8323 ( .A1(n6560), .A2(n6694), .ZN(n6933) );
  INV_X1 U8324 ( .A(n19452), .ZN(n19352) );
  INV_X1 U8325 ( .A(n23505), .ZN(n23525) );
  INV_X1 U8326 ( .A(n20134), .ZN(n19755) );
  INV_X1 U8327 ( .A(n3362), .ZN(n7475) );
  XNOR2_X1 U8328 ( .A(n8591), .B(n8590), .ZN(n10006) );
  XNOR2_X1 U8329 ( .A(n8427), .B(n8238), .ZN(n8731) );
  OAI21_X2 U8330 ( .B1(n16653), .B2(n16647), .A(n15552), .ZN(n18351) );
  OAI21_X1 U8332 ( .B1(n9024), .B2(n9886), .A(n2720), .ZN(n8179) );
  OAI21_X1 U8333 ( .B1(n1376), .B2(n12768), .A(n4945), .ZN(n4943) );
  AOI21_X2 U8334 ( .B1(n19405), .B2(n19404), .A(n2722), .ZN(n20593) );
  NAND2_X1 U8335 ( .A1(n25064), .A2(n9814), .ZN(n9512) );
  NAND3_X1 U8337 ( .A1(n3734), .A2(n20176), .A3(n20588), .ZN(n2725) );
  OAI22_X1 U8338 ( .A1(n4270), .A2(n16268), .B1(n16004), .B2(n15758), .ZN(
        n3709) );
  NAND2_X1 U8340 ( .A1(n3452), .A2(n3455), .ZN(n12748) );
  NAND2_X1 U8341 ( .A1(n16146), .A2(n16145), .ZN(n16152) );
  NAND2_X1 U8342 ( .A1(n5375), .A2(n16622), .ZN(n2727) );
  NAND2_X1 U8344 ( .A1(n2732), .A2(n2731), .ZN(n2730) );
  NAND2_X1 U8345 ( .A1(n10122), .A2(n9843), .ZN(n2731) );
  NAND2_X1 U8346 ( .A1(n2868), .A2(n23236), .ZN(n3124) );
  NAND2_X1 U8347 ( .A1(n2816), .A2(n2819), .ZN(n2734) );
  NAND2_X1 U8349 ( .A1(n5087), .A2(n7022), .ZN(n2736) );
  NAND2_X1 U8352 ( .A1(n5015), .A2(n8005), .ZN(n7540) );
  OAI211_X1 U8353 ( .C1(n12582), .C2(n12844), .A(n12581), .B(n12845), .ZN(
        n13427) );
  NAND2_X1 U8354 ( .A1(n24085), .A2(n2740), .ZN(n3742) );
  AND2_X1 U8355 ( .A1(n9529), .A2(n9806), .ZN(n10114) );
  NAND3_X1 U8358 ( .A1(n7307), .A2(n7114), .A3(n6190), .ZN(n6193) );
  XOR2_X1 U8359 ( .A(n12121), .B(n12378), .Z(n3881) );
  XNOR2_X1 U8360 ( .A(n9012), .B(n8940), .ZN(n2785) );
  INV_X1 U8361 ( .A(n19952), .ZN(n3933) );
  NAND2_X1 U8362 ( .A1(n2748), .A2(n3550), .ZN(n7362) );
  NAND2_X1 U8363 ( .A1(n15688), .A2(n15471), .ZN(n3872) );
  NAND2_X1 U8364 ( .A1(n6218), .A2(n7250), .ZN(n2750) );
  XNOR2_X1 U8365 ( .A(n18675), .B(n4711), .ZN(n17716) );
  NAND3_X1 U8367 ( .A1(n12629), .A2(n3889), .A3(n14945), .ZN(n3884) );
  OAI21_X1 U8368 ( .B1(n10369), .B2(n10365), .A(n2751), .ZN(n9770) );
  INV_X1 U8370 ( .A(n7043), .ZN(n3729) );
  NAND2_X1 U8371 ( .A1(n2752), .A2(n3532), .ZN(n4577) );
  NAND2_X1 U8373 ( .A1(n15790), .A2(n16042), .ZN(n15266) );
  NAND3_X1 U8374 ( .A1(n4256), .A2(n10080), .A3(n10088), .ZN(n4521) );
  XNOR2_X1 U8377 ( .A(n17932), .B(n17756), .ZN(n17761) );
  XNOR2_X1 U8378 ( .A(n18195), .B(n18276), .ZN(n17756) );
  NAND2_X1 U8379 ( .A1(n9531), .A2(n9806), .ZN(n9335) );
  NAND3_X1 U8381 ( .A1(n3192), .A2(n24861), .A3(n7899), .ZN(n2759) );
  XNOR2_X1 U8382 ( .A(n17973), .B(n17972), .ZN(n19094) );
  INV_X1 U8383 ( .A(n13427), .ZN(n13627) );
  OR2_X1 U8384 ( .A1(n11522), .A2(n10922), .ZN(n10525) );
  OAI21_X1 U8385 ( .B1(n23138), .B2(n23143), .A(n23145), .ZN(n4631) );
  NAND2_X1 U8386 ( .A1(n23138), .A2(n23154), .ZN(n23145) );
  NAND2_X1 U8388 ( .A1(n2807), .A2(n7284), .ZN(n2806) );
  XNOR2_X1 U8389 ( .A(n2760), .B(n20625), .ZN(Ciphertext[167]) );
  OR2_X1 U8390 ( .A1(n6426), .A2(n4621), .ZN(n5449) );
  NOR2_X1 U8392 ( .A1(n16220), .A2(n16219), .ZN(n16466) );
  INV_X1 U8393 ( .A(n13317), .ZN(n12844) );
  OR2_X1 U8394 ( .A1(n5434), .A2(n17069), .ZN(n5462) );
  OR2_X1 U8396 ( .A1(n13703), .A2(n14250), .ZN(n13704) );
  OR2_X1 U8397 ( .A1(n25200), .A2(n17212), .ZN(n16556) );
  INV_X1 U8398 ( .A(n10846), .ZN(n11124) );
  XNOR2_X1 U8399 ( .A(n18448), .B(n18254), .ZN(n17990) );
  AND2_X1 U8400 ( .A1(n7268), .A2(n7843), .ZN(n3266) );
  NOR2_X1 U8401 ( .A1(n3717), .A2(n14150), .ZN(n13513) );
  INV_X1 U8402 ( .A(n17012), .ZN(n17353) );
  NOR2_X1 U8403 ( .A1(n3027), .A2(n23357), .ZN(n23358) );
  XNOR2_X1 U8404 ( .A(n18090), .B(n18089), .ZN(n19591) );
  INV_X1 U8405 ( .A(n7278), .ZN(n8023) );
  INV_X1 U8406 ( .A(n16431), .ZN(n17522) );
  INV_X1 U8407 ( .A(n12648), .ZN(n13096) );
  NOR2_X1 U8408 ( .A1(n23860), .A2(n24675), .ZN(n4904) );
  XNOR2_X1 U8409 ( .A(n21168), .B(n4455), .ZN(n22449) );
  XNOR2_X1 U8410 ( .A(n8410), .B(n8409), .ZN(n9348) );
  NAND2_X1 U8412 ( .A1(n10309), .A2(n11160), .ZN(n2763) );
  INV_X1 U8413 ( .A(n7347), .ZN(n8512) );
  NAND2_X1 U8414 ( .A1(n13063), .A2(n24601), .ZN(n13065) );
  AOI22_X2 U8415 ( .A1(n6790), .A2(n6789), .B1(n6787), .B2(n6788), .ZN(n7975)
         );
  NAND2_X1 U8416 ( .A1(n11521), .A2(n3771), .ZN(n3770) );
  XNOR2_X1 U8417 ( .A(n13906), .B(n2765), .ZN(n15167) );
  NOR2_X1 U8421 ( .A1(n367), .A2(n17356), .ZN(n2767) );
  OAI22_X1 U8422 ( .A1(n12716), .A2(n13165), .B1(n12717), .B2(n13167), .ZN(
        n12723) );
  NAND2_X1 U8423 ( .A1(n12718), .A2(n4766), .ZN(n12716) );
  NAND2_X1 U8424 ( .A1(n338), .A2(n22967), .ZN(n22129) );
  NAND2_X1 U8425 ( .A1(n7319), .A2(n3300), .ZN(n2768) );
  NAND2_X1 U8426 ( .A1(n14031), .A2(n14151), .ZN(n4963) );
  NAND2_X1 U8428 ( .A1(n284), .A2(n16628), .ZN(n16630) );
  NOR2_X1 U8429 ( .A1(n24487), .A2(n5175), .ZN(n5174) );
  NAND2_X1 U8430 ( .A1(n14146), .A2(n14198), .ZN(n14147) );
  NAND2_X1 U8431 ( .A1(n15940), .A2(n16253), .ZN(n2771) );
  NAND2_X1 U8432 ( .A1(n7950), .A2(n7949), .ZN(n2773) );
  NAND3_X1 U8433 ( .A1(n10075), .A2(n10068), .A3(n10070), .ZN(n2778) );
  OAI21_X1 U8434 ( .B1(n17712), .B2(n19352), .A(n2779), .ZN(n17713) );
  NAND3_X1 U8435 ( .A1(n17711), .A2(n19444), .A3(n25002), .ZN(n2779) );
  NAND2_X1 U8436 ( .A1(n16161), .A2(n16391), .ZN(n15621) );
  NAND2_X1 U8437 ( .A1(n15977), .A2(n16389), .ZN(n16161) );
  XNOR2_X1 U8438 ( .A(n17816), .B(n17900), .ZN(n18348) );
  NAND2_X1 U8439 ( .A1(n15792), .A2(n15791), .ZN(n16575) );
  OR2_X1 U8441 ( .A1(n12763), .A2(n11580), .ZN(n11595) );
  OR2_X1 U8442 ( .A1(n16961), .A2(n16828), .ZN(n4817) );
  AND2_X1 U8443 ( .A1(n10851), .A2(n305), .ZN(n2959) );
  OR2_X1 U8444 ( .A1(n9885), .A2(n8157), .ZN(n9024) );
  AND2_X1 U8445 ( .A1(n7023), .A2(n7021), .ZN(n5087) );
  XNOR2_X1 U8448 ( .A(n17882), .B(n18463), .ZN(n5159) );
  XNOR2_X1 U8449 ( .A(n4024), .B(n8982), .ZN(n8984) );
  NAND2_X1 U8450 ( .A1(n10524), .A2(n11529), .ZN(n10526) );
  OAI21_X1 U8451 ( .B1(n21188), .B2(n21189), .A(n24043), .ZN(n2781) );
  NAND2_X1 U8452 ( .A1(n6722), .A2(n316), .ZN(n6115) );
  BUF_X1 U8453 ( .A(n6208), .Z(n6296) );
  OAI22_X1 U8456 ( .A1(n9949), .A2(n9955), .B1(n9388), .B2(n9269), .ZN(n9360)
         );
  NAND3_X1 U8457 ( .A1(n6838), .A2(n6987), .A3(n6244), .ZN(n6839) );
  NAND2_X1 U8458 ( .A1(n4976), .A2(n7856), .ZN(n4975) );
  AOI22_X1 U8461 ( .A1(n23771), .A2(n23772), .B1(n23777), .B2(n2783), .ZN(
        n23773) );
  INV_X1 U8464 ( .A(n17312), .ZN(n2968) );
  NAND2_X1 U8466 ( .A1(n3255), .A2(n12847), .ZN(n13503) );
  NAND2_X1 U8467 ( .A1(n5910), .A2(n6146), .ZN(n6145) );
  NAND2_X1 U8468 ( .A1(n4901), .A2(n7732), .ZN(n2787) );
  OR2_X1 U8470 ( .A1(n6970), .A2(n6969), .ZN(n2788) );
  NAND2_X1 U8471 ( .A1(n11529), .A2(n11524), .ZN(n3182) );
  NAND2_X1 U8473 ( .A1(n16240), .A2(n17216), .ZN(n2789) );
  NAND2_X1 U8474 ( .A1(n3117), .A2(n9251), .ZN(n3116) );
  OAI21_X2 U8475 ( .B1(n13749), .B2(n13748), .A(n13747), .ZN(n15219) );
  XNOR2_X1 U8476 ( .A(n8674), .B(n8673), .ZN(n8677) );
  NAND2_X1 U8478 ( .A1(n2792), .A2(n2791), .ZN(n12444) );
  NAND2_X1 U8479 ( .A1(n13049), .A2(n12490), .ZN(n2791) );
  NAND2_X1 U8480 ( .A1(n13024), .A2(n12786), .ZN(n12787) );
  NAND2_X1 U8481 ( .A1(n2794), .A2(n2793), .ZN(n12790) );
  NAND2_X1 U8482 ( .A1(n12785), .A2(n302), .ZN(n2793) );
  NOR2_X1 U8485 ( .A1(n19558), .A2(n19555), .ZN(n19140) );
  NAND2_X1 U8486 ( .A1(n21476), .A2(n22965), .ZN(n21959) );
  XNOR2_X1 U8489 ( .A(n8911), .B(n8912), .ZN(n9989) );
  OR2_X1 U8490 ( .A1(n11045), .A2(n11051), .ZN(n11013) );
  AND2_X1 U8491 ( .A1(n4351), .A2(n4348), .ZN(n3476) );
  INV_X1 U8492 ( .A(n19598), .ZN(n19601) );
  XNOR2_X1 U8494 ( .A(n2797), .B(n8570), .ZN(n8571) );
  XNOR2_X1 U8495 ( .A(n8566), .B(n8567), .ZN(n2797) );
  NAND2_X1 U8496 ( .A1(n10812), .A2(n5085), .ZN(n3870) );
  NAND2_X1 U8497 ( .A1(n2799), .A2(n2798), .ZN(n23223) );
  NAND2_X1 U8498 ( .A1(n23221), .A2(n24967), .ZN(n2798) );
  NAND2_X1 U8499 ( .A1(n23222), .A2(n23218), .ZN(n2799) );
  OAI21_X1 U8500 ( .B1(n6811), .B2(n6371), .A(n7002), .ZN(n2801) );
  INV_X1 U8501 ( .A(n2803), .ZN(n2802) );
  OAI22_X1 U8502 ( .A1(n18918), .A2(n18919), .B1(n18917), .B2(n18916), .ZN(
        n2803) );
  AOI22_X1 U8503 ( .A1(n9761), .A2(n427), .B1(n9760), .B2(n1330), .ZN(n10674)
         );
  OAI211_X2 U8504 ( .C1(n1551), .C2(n1423), .A(n2804), .B(n4841), .ZN(n20289)
         );
  OR2_X1 U8506 ( .A1(n22945), .A2(n21531), .ZN(n4170) );
  INV_X1 U8507 ( .A(n20688), .ZN(n3087) );
  NOR2_X1 U8508 ( .A1(n3615), .A2(n8021), .ZN(n3614) );
  NAND2_X1 U8511 ( .A1(n2636), .A2(n2809), .ZN(n16444) );
  NAND3_X1 U8513 ( .A1(n24103), .A2(n7896), .A3(n7897), .ZN(n5901) );
  NAND2_X1 U8514 ( .A1(n9136), .A2(n2810), .ZN(n10371) );
  NAND2_X1 U8517 ( .A1(n16500), .A2(n25572), .ZN(n2811) );
  NAND3_X1 U8518 ( .A1(n11045), .A2(n4531), .A3(n11046), .ZN(n10643) );
  XNOR2_X1 U8520 ( .A(n13524), .B(n15281), .ZN(n2812) );
  OAI211_X1 U8521 ( .C1(n2814), .C2(n17085), .A(n17086), .B(n2813), .ZN(n15552) );
  INV_X1 U8523 ( .A(n17087), .ZN(n2815) );
  NAND2_X1 U8524 ( .A1(n2818), .A2(n2817), .ZN(n2816) );
  INV_X1 U8525 ( .A(n22221), .ZN(n2817) );
  NAND2_X1 U8526 ( .A1(n22214), .A2(n25461), .ZN(n2818) );
  NAND2_X1 U8527 ( .A1(n21789), .A2(n22221), .ZN(n2819) );
  NAND2_X1 U8530 ( .A1(n10907), .A2(n10901), .ZN(n10444) );
  INV_X1 U8531 ( .A(n13158), .ZN(n12666) );
  NAND2_X1 U8532 ( .A1(n13338), .A2(n13335), .ZN(n12838) );
  NOR2_X2 U8533 ( .A1(n16719), .A2(n2823), .ZN(n18637) );
  NAND2_X1 U8535 ( .A1(n13949), .A2(n13463), .ZN(n13464) );
  NAND3_X1 U8536 ( .A1(n2827), .A2(n22555), .A3(n22554), .ZN(n22557) );
  NAND3_X1 U8537 ( .A1(n22552), .A2(n22553), .A3(n22551), .ZN(n2827) );
  AOI22_X1 U8538 ( .A1(n15472), .A2(n17341), .B1(n17235), .B2(n16780), .ZN(
        n2829) );
  OR2_X1 U8539 ( .A1(n19233), .A2(n19112), .ZN(n4141) );
  NAND2_X1 U8541 ( .A1(n3985), .A2(n3986), .ZN(n3984) );
  OAI21_X1 U8544 ( .B1(n22263), .B2(n22264), .A(n22262), .ZN(n2833) );
  NAND3_X1 U8545 ( .A1(n3295), .A2(n3293), .A3(n3405), .ZN(n10482) );
  OAI22_X1 U8546 ( .A1(n23660), .A2(n23686), .B1(n23662), .B2(n23661), .ZN(
        n23664) );
  AOI21_X1 U8547 ( .B1(n10462), .B2(n10463), .A(n5077), .ZN(n4501) );
  OR2_X1 U8549 ( .A1(n10087), .A2(n10088), .ZN(n2835) );
  NAND2_X1 U8550 ( .A1(n11195), .A2(n11199), .ZN(n10479) );
  INV_X1 U8551 ( .A(n7155), .ZN(n7365) );
  OR2_X1 U8552 ( .A1(n9723), .A2(n9484), .ZN(n9655) );
  XNOR2_X1 U8553 ( .A(n14741), .B(n14740), .ZN(n5192) );
  INV_X1 U8554 ( .A(n4114), .ZN(n19367) );
  INV_X1 U8555 ( .A(n14944), .ZN(n12629) );
  XNOR2_X2 U8556 ( .A(n2839), .B(n2838), .ZN(n16106) );
  XNOR2_X1 U8557 ( .A(n15195), .B(n15447), .ZN(n2838) );
  XNOR2_X1 U8558 ( .A(n15156), .B(n14668), .ZN(n2839) );
  NAND3_X1 U8560 ( .A1(n3515), .A2(n3516), .A3(n17013), .ZN(n3514) );
  XNOR2_X1 U8561 ( .A(n3605), .B(n18541), .ZN(n18039) );
  INV_X1 U8562 ( .A(n15899), .ZN(n15676) );
  XNOR2_X1 U8564 ( .A(n8960), .B(n8244), .ZN(n8436) );
  AOI21_X1 U8565 ( .B1(n4729), .B2(n12407), .A(n13347), .ZN(n12421) );
  NAND2_X1 U8566 ( .A1(n13957), .A2(n14311), .ZN(n13904) );
  NAND3_X1 U8569 ( .A1(n12935), .A2(n13235), .A3(n2842), .ZN(n13238) );
  NOR2_X1 U8571 ( .A1(n16302), .A2(n16022), .ZN(n16299) );
  AOI21_X1 U8572 ( .B1(n15917), .B2(n25092), .A(n15916), .ZN(n15918) );
  INV_X1 U8573 ( .A(n13903), .ZN(n4525) );
  NAND3_X1 U8574 ( .A1(n6147), .A2(n6678), .A3(n2843), .ZN(n6148) );
  NAND2_X1 U8575 ( .A1(n6679), .A2(n6281), .ZN(n6147) );
  OAI21_X1 U8579 ( .B1(n18897), .B2(n18896), .A(n18895), .ZN(n2844) );
  NAND2_X1 U8581 ( .A1(n2846), .A2(n2845), .ZN(n7233) );
  NAND2_X1 U8582 ( .A1(n3469), .A2(n248), .ZN(n2845) );
  OR2_X1 U8584 ( .A1(n9753), .A2(n9613), .ZN(n9750) );
  OR2_X1 U8585 ( .A1(n4980), .A2(n14165), .ZN(n4979) );
  OR2_X1 U8586 ( .A1(n16311), .A2(n25410), .ZN(n3743) );
  OAI21_X1 U8588 ( .B1(n7648), .B2(n7651), .A(n7305), .ZN(n2848) );
  NAND4_X2 U8589 ( .A1(n7830), .A2(n7831), .A3(n7832), .A4(n7833), .ZN(n8667)
         );
  NAND2_X1 U8590 ( .A1(n16450), .A2(n223), .ZN(n15929) );
  NAND3_X1 U8591 ( .A1(n9706), .A2(n10062), .A3(n10064), .ZN(n9707) );
  NAND4_X2 U8592 ( .A1(n8017), .A2(n8020), .A3(n8018), .A4(n8019), .ZN(n9169)
         );
  NAND2_X1 U8593 ( .A1(n2850), .A2(n7005), .ZN(n5145) );
  OAI21_X1 U8594 ( .B1(n7011), .B2(n6650), .A(n6649), .ZN(n2850) );
  INV_X1 U8595 ( .A(n12017), .ZN(n4448) );
  XNOR2_X1 U8596 ( .A(n11753), .B(n12395), .ZN(n13224) );
  MUX2_X2 U8597 ( .A(n22720), .B(n22719), .S(n22893), .Z(n23499) );
  INV_X1 U8599 ( .A(n15657), .ZN(n4046) );
  AOI21_X1 U8601 ( .B1(n2851), .B2(n13313), .A(n13923), .ZN(n13314) );
  NAND2_X1 U8602 ( .A1(n14253), .A2(n13924), .ZN(n2851) );
  NAND2_X1 U8603 ( .A1(n14118), .A2(n14221), .ZN(n13403) );
  NAND2_X1 U8604 ( .A1(n13399), .A2(n14219), .ZN(n14118) );
  NAND3_X1 U8605 ( .A1(n21712), .A2(n22072), .A3(n22916), .ZN(n2853) );
  NOR2_X1 U8606 ( .A1(n19973), .A2(n19974), .ZN(n21534) );
  XOR2_X1 U8608 ( .A(n18666), .B(n18239), .Z(n4855) );
  OR2_X1 U8610 ( .A1(n25486), .A2(n9845), .ZN(n9523) );
  OR2_X1 U8611 ( .A1(n9527), .A2(n9772), .ZN(n2855) );
  OR2_X1 U8612 ( .A1(n11806), .A2(n13968), .ZN(n3425) );
  NAND2_X1 U8613 ( .A1(n12630), .A2(n13117), .ZN(n12631) );
  NAND2_X1 U8614 ( .A1(n3607), .A2(n10325), .ZN(n10330) );
  INV_X1 U8615 ( .A(n22394), .ZN(n2857) );
  NAND2_X1 U8616 ( .A1(n6121), .A2(n6642), .ZN(n6124) );
  MUX2_X1 U8620 ( .A(n20353), .B(n20476), .S(n20480), .Z(n2864) );
  NAND2_X1 U8621 ( .A1(n10759), .A2(n10757), .ZN(n2865) );
  NAND2_X1 U8622 ( .A1(n10758), .A2(n2867), .ZN(n2866) );
  XNOR2_X1 U8623 ( .A(n11868), .B(n3648), .ZN(n3647) );
  NOR2_X1 U8624 ( .A1(n23256), .A2(n2869), .ZN(n2868) );
  AND2_X1 U8626 ( .A1(n9281), .A2(n9468), .ZN(n9471) );
  OAI22_X1 U8628 ( .A1(n10512), .A2(n10570), .B1(n2870), .B2(n11038), .ZN(
        n3058) );
  OR2_X1 U8629 ( .A1(n9459), .A2(n9460), .ZN(n9465) );
  NOR2_X1 U8630 ( .A1(n20014), .A2(n20019), .ZN(n5405) );
  NOR2_X1 U8631 ( .A1(n9683), .A2(n9684), .ZN(n8978) );
  XNOR2_X1 U8633 ( .A(n12325), .B(n12144), .ZN(n11388) );
  OAI21_X2 U8634 ( .B1(n5671), .B2(n2680), .A(n10645), .ZN(n12144) );
  NAND3_X1 U8635 ( .A1(n3615), .A2(n8023), .A3(n7747), .ZN(n7745) );
  NAND2_X1 U8637 ( .A1(n12670), .A2(n12671), .ZN(n12677) );
  NAND2_X1 U8638 ( .A1(n2871), .A2(n5341), .ZN(n5340) );
  NAND2_X1 U8639 ( .A1(n9391), .A2(n9953), .ZN(n2871) );
  AOI22_X2 U8640 ( .A1(n19274), .A2(n362), .B1(n2872), .B2(n19570), .ZN(n20414) );
  NAND2_X1 U8641 ( .A1(n5632), .A2(n19569), .ZN(n2872) );
  NAND2_X1 U8642 ( .A1(n7918), .A2(n7917), .ZN(n8076) );
  NAND2_X1 U8644 ( .A1(n9325), .A2(n9788), .ZN(n5353) );
  INV_X1 U8645 ( .A(n14104), .ZN(n4875) );
  XOR2_X1 U8649 ( .A(n21324), .B(n23045), .Z(n4456) );
  XNOR2_X1 U8650 ( .A(n21455), .B(n21039), .ZN(n21041) );
  NAND2_X1 U8653 ( .A1(n11089), .A2(n419), .ZN(n2878) );
  NAND2_X1 U8654 ( .A1(n7957), .A2(n2880), .ZN(n8770) );
  AND3_X2 U8655 ( .A1(n5679), .A2(n11027), .A3(n11028), .ZN(n12234) );
  OR2_X1 U8656 ( .A1(n5673), .A2(n12928), .ZN(n4457) );
  INV_X1 U8657 ( .A(n4899), .ZN(n4898) );
  INV_X1 U8658 ( .A(n16616), .ZN(n16705) );
  INV_X1 U8659 ( .A(n13224), .ZN(n13009) );
  NAND2_X1 U8660 ( .A1(n2884), .A2(n18807), .ZN(n4550) );
  NAND2_X1 U8661 ( .A1(n4551), .A2(n19250), .ZN(n2884) );
  INV_X1 U8662 ( .A(n23748), .ZN(n22308) );
  MUX2_X2 U8664 ( .A(n14121), .B(n14120), .S(n14119), .Z(n15284) );
  NAND2_X1 U8665 ( .A1(n10411), .A2(n10612), .ZN(n10616) );
  NAND2_X1 U8666 ( .A1(n16285), .A2(n16342), .ZN(n15679) );
  NAND2_X1 U8667 ( .A1(n21762), .A2(n22926), .ZN(n2887) );
  NAND2_X1 U8668 ( .A1(n7769), .A2(n7771), .ZN(n7770) );
  NAND2_X1 U8669 ( .A1(n7767), .A2(n7527), .ZN(n7769) );
  OAI21_X1 U8670 ( .B1(n16923), .B2(n17320), .A(n16924), .ZN(n2890) );
  OAI21_X1 U8672 ( .B1(n19335), .B2(n19496), .A(n19334), .ZN(n19338) );
  NAND2_X1 U8673 ( .A1(n19335), .A2(n25459), .ZN(n19334) );
  NAND2_X1 U8674 ( .A1(n4520), .A2(n4929), .ZN(n4928) );
  OR2_X1 U8675 ( .A1(n12483), .A2(n12707), .ZN(n13076) );
  INV_X1 U8676 ( .A(n2891), .ZN(n3424) );
  OAI22_X1 U8677 ( .A1(n4922), .A2(n6871), .B1(n6876), .B2(n6874), .ZN(n5856)
         );
  NAND2_X1 U8679 ( .A1(n23941), .A2(n23937), .ZN(n23913) );
  OAI21_X1 U8680 ( .B1(n8419), .B2(n8420), .A(n8418), .ZN(n2892) );
  NAND3_X1 U8681 ( .A1(n4281), .A2(n10911), .A3(n415), .ZN(n9509) );
  INV_X1 U8682 ( .A(n6703), .ZN(n3923) );
  NAND2_X1 U8683 ( .A1(n2894), .A2(n7651), .ZN(n2893) );
  INV_X1 U8684 ( .A(n7649), .ZN(n2894) );
  NAND2_X1 U8685 ( .A1(n2895), .A2(n10370), .ZN(n10217) );
  NAND2_X1 U8686 ( .A1(n10317), .A2(n10582), .ZN(n2895) );
  NAND3_X1 U8688 ( .A1(n4825), .A2(n7908), .A3(n7365), .ZN(n2896) );
  INV_X1 U8689 ( .A(n2898), .ZN(n2897) );
  OAI21_X1 U8690 ( .B1(n7626), .B2(n7364), .A(n7627), .ZN(n2898) );
  NAND2_X1 U8691 ( .A1(n6393), .A2(n2900), .ZN(n2899) );
  OAI211_X2 U8692 ( .C1(n12444), .C2(n401), .A(n12442), .B(n12443), .ZN(n14168) );
  INV_X1 U8693 ( .A(n9844), .ZN(n3988) );
  XNOR2_X1 U8696 ( .A(n5304), .B(n16037), .ZN(n18002) );
  NAND2_X1 U8697 ( .A1(n2902), .A2(n9064), .ZN(n9689) );
  XNOR2_X2 U8698 ( .A(n9039), .B(n9038), .ZN(n9064) );
  INV_X1 U8699 ( .A(n10053), .ZN(n2902) );
  OAI21_X1 U8700 ( .B1(n5115), .B2(n19121), .A(n5467), .ZN(n5466) );
  NOR2_X1 U8701 ( .A1(n12811), .A2(n4945), .ZN(n12812) );
  AND2_X1 U8702 ( .A1(n13839), .A2(n14267), .ZN(n14276) );
  NAND2_X1 U8704 ( .A1(n12521), .A2(n13040), .ZN(n2905) );
  NAND2_X1 U8705 ( .A1(n12522), .A2(n12478), .ZN(n2906) );
  NOR2_X1 U8706 ( .A1(n19130), .A2(n3568), .ZN(n16505) );
  NAND2_X1 U8707 ( .A1(n2908), .A2(n25), .ZN(n2907) );
  NAND2_X1 U8708 ( .A1(n9512), .A2(n10168), .ZN(n2909) );
  NAND2_X1 U8709 ( .A1(n14240), .A2(n4116), .ZN(n2910) );
  NAND2_X1 U8710 ( .A1(n13932), .A2(n13933), .ZN(n2911) );
  NAND2_X1 U8711 ( .A1(n2912), .A2(n3341), .ZN(n14125) );
  NAND2_X1 U8712 ( .A1(n14124), .A2(n14205), .ZN(n2912) );
  OAI22_X1 U8713 ( .A1(n12860), .A2(n13345), .B1(n13348), .B2(n12861), .ZN(
        n5436) );
  XNOR2_X1 U8714 ( .A(n12410), .B(n12409), .ZN(n12411) );
  INV_X1 U8715 ( .A(n6072), .ZN(n7002) );
  NAND2_X1 U8716 ( .A1(n20316), .A2(n20319), .ZN(n2913) );
  OR2_X1 U8718 ( .A1(n5445), .A2(n20301), .ZN(n5443) );
  INV_X1 U8719 ( .A(n4066), .ZN(n19976) );
  XNOR2_X1 U8720 ( .A(n15040), .B(n3462), .ZN(n15332) );
  INV_X1 U8721 ( .A(n13289), .ZN(n12692) );
  NAND2_X1 U8722 ( .A1(n2914), .A2(n6893), .ZN(n6897) );
  XNOR2_X2 U8723 ( .A(Key[111]), .B(Plaintext[111]), .ZN(n6987) );
  AOI21_X1 U8724 ( .B1(n2915), .B2(n25466), .A(n12910), .ZN(n11803) );
  OR2_X1 U8725 ( .A1(n13966), .A2(n13968), .ZN(n3426) );
  AOI22_X1 U8727 ( .A1(n5497), .A2(n14009), .B1(n14251), .B2(n13923), .ZN(
        n13927) );
  NAND2_X1 U8728 ( .A1(n17179), .A2(n17185), .ZN(n16873) );
  OAI21_X1 U8730 ( .B1(n6746), .B2(n6630), .A(n6750), .ZN(n6633) );
  NAND2_X1 U8733 ( .A1(n23312), .A2(n2920), .ZN(n2919) );
  OR2_X1 U8734 ( .A1(n16706), .A2(n16708), .ZN(n5556) );
  XNOR2_X1 U8735 ( .A(n17899), .B(n4155), .ZN(n17771) );
  AOI22_X1 U8736 ( .A1(n2923), .A2(n2922), .B1(n10012), .B2(n9724), .ZN(n11172) );
  INV_X1 U8737 ( .A(n9652), .ZN(n2922) );
  NAND2_X1 U8738 ( .A1(n8609), .A2(n9725), .ZN(n2923) );
  NAND3_X1 U8739 ( .A1(n3513), .A2(n10548), .A3(n10504), .ZN(n3510) );
  NOR2_X1 U8740 ( .A1(n19499), .A2(n19498), .ZN(n18721) );
  OAI21_X1 U8741 ( .B1(n5144), .B2(n25325), .A(n6503), .ZN(n5142) );
  NAND3_X1 U8742 ( .A1(n16942), .A2(n17408), .A3(n17407), .ZN(n15025) );
  NAND2_X1 U8743 ( .A1(n3690), .A2(n2924), .ZN(n13907) );
  AOI22_X1 U8744 ( .A1(n13248), .A2(n13245), .B1(n11288), .B2(n12808), .ZN(
        n2924) );
  OAI21_X2 U8745 ( .B1(n3041), .B2(n2925), .A(n20020), .ZN(n3823) );
  NAND2_X1 U8746 ( .A1(n20015), .A2(n20016), .ZN(n2925) );
  NAND2_X1 U8747 ( .A1(n5190), .A2(n21384), .ZN(n2926) );
  OAI211_X1 U8748 ( .C1(n9928), .C2(n9600), .A(n9599), .B(n2928), .ZN(n4731)
         );
  XNOR2_X2 U8750 ( .A(n17586), .B(n17585), .ZN(n19477) );
  NAND2_X1 U8751 ( .A1(n6944), .A2(n5909), .ZN(n2930) );
  NAND2_X1 U8752 ( .A1(n2932), .A2(n6940), .ZN(n2931) );
  NAND2_X1 U8753 ( .A1(n6679), .A2(n6146), .ZN(n2932) );
  NAND2_X1 U8754 ( .A1(n16951), .A2(n17287), .ZN(n2933) );
  NAND2_X1 U8755 ( .A1(n14521), .A2(n15804), .ZN(n2934) );
  NAND2_X1 U8756 ( .A1(n2936), .A2(n12763), .ZN(n4638) );
  NAND2_X1 U8757 ( .A1(n4640), .A2(n4639), .ZN(n2936) );
  OAI21_X1 U8758 ( .B1(n13048), .B2(n13051), .A(n2940), .ZN(n2939) );
  NAND2_X1 U8759 ( .A1(n13049), .A2(n13048), .ZN(n2940) );
  NAND2_X1 U8760 ( .A1(n5368), .A2(n25408), .ZN(n2941) );
  NAND2_X1 U8761 ( .A1(n16621), .A2(n16795), .ZN(n2942) );
  NAND2_X1 U8762 ( .A1(n20225), .A2(n20269), .ZN(n20229) );
  NAND2_X1 U8763 ( .A1(n7766), .A2(n7648), .ZN(n2943) );
  XNOR2_X1 U8764 ( .A(n2944), .B(n8218), .ZN(n9845) );
  XNOR2_X1 U8765 ( .A(n8793), .B(n8217), .ZN(n2944) );
  XNOR2_X1 U8766 ( .A(n5339), .B(n21141), .ZN(n20197) );
  XNOR2_X1 U8767 ( .A(n2945), .B(n18057), .ZN(n18059) );
  XNOR2_X1 U8768 ( .A(n18056), .B(n25194), .ZN(n2945) );
  NAND3_X1 U8769 ( .A1(n19952), .A2(n19951), .A3(n20593), .ZN(n19783) );
  AOI21_X1 U8770 ( .B1(n19437), .B2(n19438), .A(n19436), .ZN(n19439) );
  NAND3_X1 U8773 ( .A1(n6499), .A2(n6500), .A3(n6498), .ZN(n6502) );
  NAND2_X1 U8775 ( .A1(n2947), .A2(n9939), .ZN(n3597) );
  NOR2_X1 U8777 ( .A1(n12770), .A2(n12769), .ZN(n12772) );
  OAI21_X2 U8778 ( .B1(n19005), .B2(n19180), .A(n19004), .ZN(n20537) );
  OAI21_X1 U8779 ( .B1(n18956), .B2(n18945), .A(n3583), .ZN(n3581) );
  INV_X1 U8781 ( .A(n7771), .ZN(n7284) );
  OAI21_X2 U8782 ( .B1(n10975), .B2(n10976), .A(n10974), .ZN(n12325) );
  NAND2_X1 U8783 ( .A1(n9946), .A2(n9945), .ZN(n9895) );
  NAND2_X1 U8784 ( .A1(n2949), .A2(n2948), .ZN(n7530) );
  NAND2_X1 U8785 ( .A1(n7524), .A2(n23), .ZN(n2948) );
  NAND2_X1 U8786 ( .A1(n16962), .A2(n24444), .ZN(n16826) );
  NAND2_X1 U8788 ( .A1(n2952), .A2(n2951), .ZN(n10209) );
  NAND2_X1 U8789 ( .A1(n9470), .A2(n262), .ZN(n2951) );
  NAND2_X1 U8790 ( .A1(n9471), .A2(n2953), .ZN(n2952) );
  INV_X1 U8791 ( .A(n9962), .ZN(n2953) );
  NAND2_X1 U8792 ( .A1(n3754), .A2(n13844), .ZN(n2955) );
  NAND2_X1 U8793 ( .A1(n24340), .A2(n10623), .ZN(n10811) );
  NAND2_X1 U8794 ( .A1(n20558), .A2(n20557), .ZN(n2956) );
  OAI21_X1 U8796 ( .B1(n13568), .B2(n13394), .A(n3698), .ZN(n13089) );
  XNOR2_X1 U8797 ( .A(n2957), .B(n14763), .ZN(n13606) );
  XNOR2_X1 U8798 ( .A(n13585), .B(n14500), .ZN(n2957) );
  AND2_X1 U8800 ( .A1(n17442), .A2(n16826), .ZN(n4819) );
  NAND3_X1 U8802 ( .A1(n6216), .A2(n8511), .A3(n7351), .ZN(n7251) );
  NAND2_X1 U8804 ( .A1(n9781), .A2(n9295), .ZN(n5082) );
  NAND2_X1 U8805 ( .A1(n9222), .A2(n9223), .ZN(n9224) );
  NAND2_X1 U8806 ( .A1(n22866), .A2(n23411), .ZN(n2960) );
  NAND2_X1 U8807 ( .A1(n8370), .A2(n3979), .ZN(n7266) );
  AND3_X1 U8808 ( .A1(n6298), .A2(n4865), .A3(n6174), .ZN(n6299) );
  OAI22_X1 U8810 ( .A1(n9430), .A2(n9737), .B1(n9978), .B2(n9429), .ZN(n2962)
         );
  NOR2_X1 U8811 ( .A1(n9431), .A2(n9982), .ZN(n2963) );
  NAND2_X1 U8812 ( .A1(n13035), .A2(n13036), .ZN(n14675) );
  XNOR2_X2 U8813 ( .A(n14899), .B(n5331), .ZN(n16029) );
  NAND2_X1 U8814 ( .A1(n24310), .A2(n4884), .ZN(n4140) );
  NAND2_X1 U8815 ( .A1(n9563), .A2(n9564), .ZN(n9570) );
  INV_X1 U8817 ( .A(n17339), .ZN(n5104) );
  OR2_X1 U8818 ( .A1(n5910), .A2(n6146), .ZN(n6945) );
  XNOR2_X2 U8819 ( .A(Key[189]), .B(Plaintext[189]), .ZN(n6445) );
  NAND2_X1 U8820 ( .A1(n16404), .A2(n16403), .ZN(n3765) );
  NAND2_X2 U8822 ( .A1(n6865), .A2(n2965), .ZN(n8987) );
  MUX2_X1 U8823 ( .A(n4951), .B(n10729), .S(n10728), .Z(n11189) );
  NAND2_X1 U8825 ( .A1(n2966), .A2(n13284), .ZN(n13286) );
  NAND2_X1 U8826 ( .A1(n13283), .A2(n13282), .ZN(n2966) );
  NAND3_X1 U8828 ( .A1(n19942), .A2(n20450), .A3(n20377), .ZN(n19943) );
  OAI21_X1 U8829 ( .B1(n2613), .B2(n17048), .A(n17049), .ZN(n16774) );
  AOI21_X2 U8830 ( .B1(n15954), .B2(n15955), .A(n16482), .ZN(n17049) );
  NAND2_X1 U8832 ( .A1(n24506), .A2(n16226), .ZN(n16298) );
  INV_X1 U8833 ( .A(n10839), .ZN(n4464) );
  NAND2_X1 U8835 ( .A1(n3499), .A2(n7580), .ZN(n3498) );
  NAND2_X1 U8836 ( .A1(n4631), .A2(n4630), .ZN(n4628) );
  INV_X1 U8838 ( .A(n7992), .ZN(n3549) );
  NOR2_X1 U8839 ( .A1(n5594), .A2(n7733), .ZN(n5593) );
  NAND2_X1 U8840 ( .A1(n15533), .A2(n15534), .ZN(n16742) );
  INV_X1 U8841 ( .A(n10518), .ZN(n4013) );
  NAND2_X1 U8842 ( .A1(n9938), .A2(n9905), .ZN(n2971) );
  NAND3_X1 U8843 ( .A1(n1485), .A2(n6618), .A3(n7419), .ZN(n2972) );
  INV_X1 U8844 ( .A(n5349), .ZN(n23449) );
  XNOR2_X2 U8845 ( .A(n20287), .B(n20288), .ZN(n22656) );
  OAI21_X2 U8847 ( .B1(n12837), .B2(n12966), .A(n12836), .ZN(n14333) );
  NAND2_X1 U8848 ( .A1(n6612), .A2(n24501), .ZN(n2973) );
  NAND3_X1 U8849 ( .A1(n6611), .A2(n6718), .A3(n6610), .ZN(n2974) );
  OR2_X1 U8850 ( .A1(n11867), .A2(n11873), .ZN(n11876) );
  NAND3_X2 U8852 ( .A1(n17097), .A2(n17095), .A3(n17096), .ZN(n18356) );
  OR2_X1 U8853 ( .A1(n13210), .A2(n5418), .ZN(n3039) );
  INV_X1 U8854 ( .A(n18902), .ZN(n19539) );
  XOR2_X1 U8855 ( .A(n18671), .B(n18083), .Z(n5135) );
  INV_X1 U8857 ( .A(n3720), .ZN(n23245) );
  NOR2_X1 U8858 ( .A1(n22279), .A2(n22280), .ZN(n22944) );
  INV_X1 U8859 ( .A(n20094), .ZN(n4017) );
  INV_X1 U8860 ( .A(n11101), .ZN(n4143) );
  INV_X1 U8861 ( .A(n20519), .ZN(n19925) );
  XNOR2_X1 U8862 ( .A(n5343), .B(n7161), .ZN(n8997) );
  NAND2_X1 U8863 ( .A1(n19372), .A2(n19376), .ZN(n19373) );
  AOI22_X1 U8864 ( .A1(n14232), .A2(n14234), .B1(n2977), .B2(n13680), .ZN(
        n14238) );
  MUX2_X1 U8865 ( .A(n4418), .B(n24249), .S(n15625), .Z(n14745) );
  XNOR2_X2 U8866 ( .A(n14572), .B(n14573), .ZN(n15625) );
  NAND2_X1 U8868 ( .A1(n18889), .A2(n25057), .ZN(n19403) );
  NAND2_X1 U8869 ( .A1(n22661), .A2(n25160), .ZN(n2978) );
  INV_X1 U8871 ( .A(n13929), .ZN(n4837) );
  NAND2_X1 U8872 ( .A1(n3926), .A2(n6956), .ZN(n4323) );
  NAND2_X1 U8873 ( .A1(n25078), .A2(n25375), .ZN(n22095) );
  NAND2_X1 U8874 ( .A1(n4322), .A2(n6960), .ZN(n4321) );
  XNOR2_X1 U8875 ( .A(n2979), .B(n14978), .ZN(n14985) );
  XNOR2_X1 U8876 ( .A(n14981), .B(n15342), .ZN(n2979) );
  NAND2_X1 U8877 ( .A1(n13118), .A2(n13117), .ZN(n2980) );
  OR2_X1 U8879 ( .A1(n1355), .A2(n14048), .ZN(n13612) );
  AOI21_X2 U8880 ( .B1(n16479), .B2(n16478), .A(n16477), .ZN(n16851) );
  NAND2_X1 U8881 ( .A1(n23554), .A2(n24057), .ZN(n23544) );
  INV_X1 U8883 ( .A(n18196), .ZN(n4666) );
  INV_X1 U8884 ( .A(n12868), .ZN(n3328) );
  NOR2_X1 U8888 ( .A1(n23766), .A2(n2982), .ZN(n23774) );
  NAND2_X1 U8889 ( .A1(n4917), .A2(n19269), .ZN(n2983) );
  INV_X1 U8890 ( .A(n4737), .ZN(n2984) );
  NOR2_X1 U8891 ( .A1(n25031), .A2(n17054), .ZN(n16721) );
  NAND2_X1 U8894 ( .A1(n2988), .A2(n2985), .ZN(n19626) );
  NAND2_X1 U8895 ( .A1(n2987), .A2(n2986), .ZN(n2985) );
  NOR2_X1 U8896 ( .A1(n22252), .A2(n21841), .ZN(n2986) );
  NAND2_X1 U8897 ( .A1(n19343), .A2(n22252), .ZN(n2988) );
  INV_X1 U8901 ( .A(n13568), .ZN(n3701) );
  NAND2_X1 U8902 ( .A1(n19764), .A2(n20591), .ZN(n19766) );
  OAI22_X1 U8903 ( .A1(n11023), .A2(n11520), .B1(n11024), .B2(n11529), .ZN(
        n11025) );
  NAND2_X1 U8904 ( .A1(n11024), .A2(n11519), .ZN(n11023) );
  INV_X1 U8905 ( .A(n7077), .ZN(n4375) );
  XNOR2_X2 U8906 ( .A(n11774), .B(n11775), .ZN(n13291) );
  NAND2_X1 U8907 ( .A1(n2993), .A2(n13790), .ZN(n13791) );
  NAND2_X1 U8908 ( .A1(n14140), .A2(n14141), .ZN(n2993) );
  OAI22_X1 U8909 ( .A1(n9229), .A2(n9709), .B1(n9711), .B2(n10039), .ZN(n2994)
         );
  INV_X1 U8910 ( .A(n5249), .ZN(n6788) );
  OAI21_X1 U8911 ( .B1(n2996), .B2(n24459), .A(n2995), .ZN(n15844) );
  NAND2_X1 U8912 ( .A1(n24459), .A2(n16125), .ZN(n2995) );
  NAND3_X1 U8913 ( .A1(n127), .A2(n6165), .A3(n6543), .ZN(n6042) );
  NOR2_X1 U8914 ( .A1(n10502), .A2(n13167), .ZN(n10531) );
  INV_X1 U8916 ( .A(n8012), .ZN(n8016) );
  NAND2_X1 U8917 ( .A1(n7002), .A2(n6815), .ZN(n5819) );
  NAND2_X1 U8919 ( .A1(n2999), .A2(n2998), .ZN(n10174) );
  NAND2_X1 U8920 ( .A1(n10171), .A2(n25046), .ZN(n2998) );
  NAND2_X1 U8923 ( .A1(n10702), .A2(n25074), .ZN(n10704) );
  OR2_X1 U8924 ( .A1(n24446), .A2(n9244), .ZN(n9688) );
  NAND2_X1 U8927 ( .A1(n16781), .A2(n17347), .ZN(n3002) );
  NAND2_X1 U8928 ( .A1(n17000), .A2(n16999), .ZN(n3005) );
  NAND3_X1 U8929 ( .A1(n4863), .A2(n22149), .A3(n4864), .ZN(n4862) );
  NAND2_X1 U8931 ( .A1(n7599), .A2(n7598), .ZN(n3006) );
  NAND2_X1 U8934 ( .A1(n15981), .A2(n16167), .ZN(n3009) );
  NAND3_X1 U8935 ( .A1(n24576), .A2(n7861), .A3(n3570), .ZN(n7872) );
  XNOR2_X1 U8936 ( .A(n18687), .B(n5304), .ZN(n5303) );
  NAND2_X1 U8937 ( .A1(n17179), .A2(n16871), .ZN(n16872) );
  NAND2_X1 U8938 ( .A1(n1324), .A2(n12725), .ZN(n12460) );
  NAND2_X1 U8939 ( .A1(n3543), .A2(n3545), .ZN(n3542) );
  NAND2_X1 U8940 ( .A1(n24386), .A2(n4435), .ZN(n16885) );
  OAI21_X2 U8941 ( .B1(n22944), .B2(n4632), .A(n3718), .ZN(n3720) );
  AND2_X1 U8942 ( .A1(n21863), .A2(n23902), .ZN(n22547) );
  NAND2_X1 U8943 ( .A1(n5290), .A2(n18765), .ZN(n19308) );
  AOI22_X2 U8944 ( .A1(n3010), .A2(n12842), .B1(n12841), .B2(n12958), .ZN(
        n14339) );
  OAI21_X1 U8945 ( .B1(n3013), .B2(n7773), .A(n3012), .ZN(n6127) );
  NAND2_X1 U8946 ( .A1(n6113), .A2(n3013), .ZN(n3012) );
  NAND2_X1 U8947 ( .A1(n25252), .A2(n7526), .ZN(n7773) );
  NAND3_X1 U8948 ( .A1(n11214), .A2(n11212), .A3(n10812), .ZN(n5627) );
  MUX2_X1 U8949 ( .A(n10555), .B(n4736), .S(n417), .Z(n4740) );
  NAND2_X1 U8951 ( .A1(n15656), .A2(n16381), .ZN(n4835) );
  AOI21_X1 U8952 ( .B1(n22290), .B2(n22291), .A(n3018), .ZN(n22292) );
  AND2_X1 U8953 ( .A1(n22289), .A2(n22387), .ZN(n3018) );
  NAND3_X1 U8954 ( .A1(n3124), .A2(n23238), .A3(n23237), .ZN(n3123) );
  XNOR2_X1 U8955 ( .A(n17756), .B(n24536), .ZN(n18049) );
  INV_X1 U8956 ( .A(n14373), .ZN(n4834) );
  NAND3_X1 U8957 ( .A1(n23743), .A2(n23748), .A3(n23740), .ZN(n3097) );
  NAND3_X1 U8958 ( .A1(n19951), .A2(n20587), .A3(n20590), .ZN(n3466) );
  NAND2_X1 U8962 ( .A1(n7514), .A2(n7977), .ZN(n7405) );
  NOR2_X1 U8963 ( .A1(n13995), .A2(n25435), .ZN(n4560) );
  INV_X1 U8964 ( .A(n10799), .ZN(n4527) );
  XNOR2_X1 U8965 ( .A(n3022), .B(n12045), .ZN(n11708) );
  XNOR2_X1 U8966 ( .A(n11705), .B(n12121), .ZN(n3022) );
  NAND2_X1 U8970 ( .A1(n22391), .A2(n22974), .ZN(n3024) );
  NAND2_X1 U8971 ( .A1(n22868), .A2(n23411), .ZN(n3025) );
  NOR2_X1 U8973 ( .A1(n23356), .A2(n23355), .ZN(n3027) );
  NOR2_X1 U8974 ( .A1(n13712), .A2(n14361), .ZN(n3030) );
  INV_X1 U8975 ( .A(n13711), .ZN(n3031) );
  NOR2_X1 U8976 ( .A1(n22415), .A2(n23300), .ZN(n23309) );
  OAI211_X1 U8977 ( .C1(n7582), .C2(n7581), .A(n7583), .B(n7882), .ZN(n5489)
         );
  NAND3_X1 U8978 ( .A1(n3796), .A2(n20569), .A3(n20570), .ZN(n3032) );
  OAI21_X1 U8979 ( .B1(n3034), .B2(n24583), .A(n3033), .ZN(n18936) );
  NAND2_X1 U8980 ( .A1(n24583), .A2(n19326), .ZN(n3033) );
  INV_X1 U8981 ( .A(n18935), .ZN(n3034) );
  OAI21_X1 U8982 ( .B1(n21915), .B2(n22404), .A(n22397), .ZN(n3035) );
  XNOR2_X1 U8983 ( .A(n3036), .B(n23191), .ZN(Ciphertext[30]) );
  XNOR2_X1 U8985 ( .A(n3038), .B(n24100), .ZN(n20779) );
  NAND2_X1 U8986 ( .A1(n3040), .A2(n23418), .ZN(n23400) );
  OAI21_X1 U8987 ( .B1(n24978), .B2(n24426), .A(n23416), .ZN(n3040) );
  NAND3_X2 U8990 ( .A1(n17303), .A2(n17302), .A3(n3376), .ZN(n18465) );
  NAND2_X1 U8991 ( .A1(n20210), .A2(n20597), .ZN(n3044) );
  NAND2_X1 U8993 ( .A1(n20209), .A2(n20208), .ZN(n3046) );
  NAND2_X1 U8994 ( .A1(n17029), .A2(n17030), .ZN(n17032) );
  NAND2_X1 U8995 ( .A1(n18968), .A2(n18967), .ZN(n3844) );
  OAI22_X1 U8997 ( .A1(n19251), .A2(n18862), .B1(n19252), .B2(n19592), .ZN(
        n3047) );
  OR2_X1 U8999 ( .A1(n6456), .A2(n6184), .ZN(n6337) );
  NAND2_X1 U9000 ( .A1(n12669), .A2(n24462), .ZN(n3562) );
  XNOR2_X1 U9001 ( .A(n8556), .B(n8557), .ZN(n3048) );
  NAND2_X1 U9002 ( .A1(n23364), .A2(n23365), .ZN(n23367) );
  OAI21_X1 U9004 ( .B1(n9867), .B2(n10053), .A(n3049), .ZN(n9245) );
  NAND2_X1 U9005 ( .A1(n3052), .A2(n5512), .ZN(n5511) );
  NOR2_X1 U9006 ( .A1(n17211), .A2(n17016), .ZN(n3052) );
  NAND2_X1 U9007 ( .A1(n3589), .A2(n12713), .ZN(n12430) );
  NAND2_X1 U9008 ( .A1(n6940), .A2(n6683), .ZN(n6144) );
  OAI21_X2 U9009 ( .B1(n7322), .B2(n7326), .A(n7325), .ZN(n8771) );
  OR2_X2 U9010 ( .A1(n6157), .A2(n6158), .ZN(n7382) );
  OAI21_X1 U9011 ( .B1(n6953), .B2(n6949), .A(n6141), .ZN(n6157) );
  OR2_X1 U9013 ( .A1(n16655), .A2(n17134), .ZN(n3053) );
  NAND2_X1 U9014 ( .A1(n17129), .A2(n16655), .ZN(n3054) );
  NAND2_X1 U9015 ( .A1(n5714), .A2(n7800), .ZN(n3056) );
  XNOR2_X1 U9016 ( .A(n3057), .B(n15303), .ZN(n14491) );
  XNOR2_X1 U9017 ( .A(n14490), .B(n15446), .ZN(n3057) );
  OAI211_X1 U9020 ( .C1(n4341), .C2(n10445), .A(n10751), .B(n9553), .ZN(n4040)
         );
  XNOR2_X1 U9021 ( .A(n18253), .B(n5327), .ZN(n5326) );
  OAI21_X1 U9022 ( .B1(n24490), .B2(n12885), .A(n3286), .ZN(n12884) );
  XOR2_X1 U9023 ( .A(n12067), .B(n3190), .Z(n3361) );
  NAND2_X1 U9024 ( .A1(n7675), .A2(n7672), .ZN(n7227) );
  OAI21_X1 U9026 ( .B1(n9403), .B2(n10734), .A(n10731), .ZN(n9404) );
  MUX2_X2 U9029 ( .A(n14134), .B(n14133), .S(n14132), .Z(n15415) );
  NAND2_X1 U9031 ( .A1(n16415), .A2(n24231), .ZN(n3060) );
  OAI21_X1 U9033 ( .B1(n13793), .B2(n13579), .A(n13769), .ZN(n4592) );
  XNOR2_X1 U9034 ( .A(n17917), .B(n17916), .ZN(n18719) );
  NAND2_X1 U9035 ( .A1(n3922), .A2(n6959), .ZN(n6958) );
  INV_X1 U9039 ( .A(n12796), .ZN(n3065) );
  NAND2_X1 U9040 ( .A1(n25370), .A2(n24569), .ZN(n3068) );
  MUX2_X2 U9042 ( .A(n17565), .B(n17564), .S(n5371), .Z(n20317) );
  NAND2_X1 U9043 ( .A1(n20054), .A2(n25089), .ZN(n20469) );
  NOR2_X1 U9044 ( .A1(n13449), .A2(n13761), .ZN(n3786) );
  INV_X1 U9045 ( .A(n7501), .ZN(n7498) );
  NAND2_X1 U9046 ( .A1(n9563), .A2(n8157), .ZN(n9248) );
  AND2_X1 U9047 ( .A1(n4117), .A2(n4118), .ZN(n12495) );
  OAI21_X1 U9048 ( .B1(n307), .B2(n4993), .A(n9872), .ZN(n3072) );
  OR2_X1 U9049 ( .A1(n13052), .A2(n13053), .ZN(n4517) );
  INV_X1 U9050 ( .A(n3717), .ZN(n14031) );
  XNOR2_X1 U9051 ( .A(n18100), .B(n18099), .ZN(n4139) );
  INV_X1 U9052 ( .A(n14245), .ZN(n13200) );
  INV_X1 U9053 ( .A(n19275), .ZN(n5572) );
  INV_X1 U9056 ( .A(n17165), .ZN(n4774) );
  INV_X1 U9057 ( .A(n15191), .ZN(n3234) );
  OAI22_X1 U9058 ( .A1(n4885), .A2(n19609), .B1(n19610), .B2(n24310), .ZN(
        n19611) );
  XNOR2_X1 U9059 ( .A(n14377), .B(n15165), .ZN(n14898) );
  NAND3_X1 U9060 ( .A1(n10989), .A2(n10406), .A3(n3606), .ZN(n3607) );
  NAND3_X1 U9061 ( .A1(n3074), .A2(n6769), .A3(n6909), .ZN(n6485) );
  NAND2_X1 U9062 ( .A1(n6910), .A2(n6918), .ZN(n3074) );
  NAND2_X1 U9063 ( .A1(n23902), .A2(n25239), .ZN(n3077) );
  NAND3_X1 U9064 ( .A1(n23903), .A2(n23902), .A3(n23904), .ZN(n3078) );
  NAND2_X1 U9065 ( .A1(n10803), .A2(n10801), .ZN(n3079) );
  NAND2_X1 U9066 ( .A1(n21377), .A2(n3080), .ZN(n23154) );
  OAI21_X1 U9067 ( .B1(n21376), .B2(n22328), .A(n22462), .ZN(n3080) );
  NAND2_X1 U9068 ( .A1(n3081), .A2(n14126), .ZN(n13899) );
  OAI22_X1 U9069 ( .A1(n13893), .A2(n14130), .B1(n13895), .B2(n4133), .ZN(
        n3081) );
  NOR2_X1 U9070 ( .A1(n16929), .A2(n24585), .ZN(n16720) );
  OAI21_X1 U9071 ( .B1(n13017), .B2(n13014), .A(n12756), .ZN(n13242) );
  XNOR2_X1 U9072 ( .A(n3086), .B(n21398), .ZN(Ciphertext[36]) );
  NAND2_X1 U9073 ( .A1(n14182), .A2(n13795), .ZN(n13773) );
  NAND3_X1 U9074 ( .A1(n6530), .A2(n6532), .A3(n6533), .ZN(n5920) );
  NAND2_X1 U9077 ( .A1(n3091), .A2(n3090), .ZN(n22260) );
  NAND2_X1 U9078 ( .A1(n25460), .A2(n22258), .ZN(n3090) );
  NAND2_X1 U9079 ( .A1(n22259), .A2(n997), .ZN(n3091) );
  XNOR2_X2 U9081 ( .A(n5940), .B(Key[5]), .ZN(n6510) );
  AOI21_X1 U9082 ( .B1(n2953), .B2(n3292), .A(n3289), .ZN(n10208) );
  AND3_X1 U9083 ( .A1(n5995), .A2(n5994), .A3(n6596), .ZN(n3167) );
  NAND2_X1 U9084 ( .A1(n20192), .A2(n3198), .ZN(n20434) );
  OAI21_X2 U9085 ( .B1(n20327), .B2(n20571), .A(n20326), .ZN(n21606) );
  NAND2_X1 U9086 ( .A1(n7602), .A2(n7257), .ZN(n7258) );
  XNOR2_X1 U9088 ( .A(n14493), .B(n21711), .ZN(n14185) );
  XNOR2_X1 U9089 ( .A(n11915), .B(n3812), .ZN(n10239) );
  NAND3_X1 U9090 ( .A1(n24286), .A2(n1357), .A3(n11151), .ZN(n4999) );
  OR2_X1 U9091 ( .A1(n6473), .A2(n6373), .ZN(n6091) );
  NAND2_X1 U9092 ( .A1(n12891), .A2(n13207), .ZN(n13210) );
  XNOR2_X2 U9093 ( .A(n11358), .B(n11359), .ZN(n13207) );
  NAND2_X1 U9095 ( .A1(n3094), .A2(n4262), .ZN(n4260) );
  INV_X1 U9096 ( .A(n7108), .ZN(n7747) );
  NAND2_X1 U9100 ( .A1(n25460), .A2(n3096), .ZN(n3095) );
  NOR2_X1 U9101 ( .A1(n23748), .A2(n23730), .ZN(n3096) );
  NAND3_X1 U9103 ( .A1(n10799), .A2(n10649), .A3(n411), .ZN(n3098) );
  INV_X1 U9104 ( .A(n10649), .ZN(n3100) );
  NAND3_X2 U9105 ( .A1(n3145), .A2(n11049), .A3(n3144), .ZN(n12197) );
  NAND2_X1 U9106 ( .A1(n3101), .A2(n22141), .ZN(n3961) );
  NAND2_X1 U9107 ( .A1(n21910), .A2(n22333), .ZN(n3101) );
  OAI21_X2 U9109 ( .B1(n3656), .B2(n20464), .A(n3102), .ZN(n21693) );
  NAND2_X1 U9110 ( .A1(n20462), .A2(n20463), .ZN(n3102) );
  OAI21_X1 U9111 ( .B1(n6323), .B2(n6523), .A(n6276), .ZN(n3407) );
  NAND2_X1 U9112 ( .A1(n19304), .A2(n19132), .ZN(n18765) );
  NAND2_X1 U9114 ( .A1(n3104), .A2(n3103), .ZN(n16650) );
  NAND2_X1 U9115 ( .A1(n16648), .A2(n17088), .ZN(n3104) );
  XNOR2_X1 U9116 ( .A(n3105), .B(n9021), .ZN(n9237) );
  XNOR2_X1 U9117 ( .A(n9019), .B(n9020), .ZN(n3105) );
  NAND2_X1 U9118 ( .A1(n2008), .A2(n6697), .ZN(n5897) );
  NAND2_X1 U9119 ( .A1(n19207), .A2(n25474), .ZN(n3106) );
  MUX2_X2 U9120 ( .A(n10289), .B(n10288), .S(n11111), .Z(n12186) );
  OR2_X1 U9121 ( .A1(n10698), .A2(n25074), .ZN(n10700) );
  INV_X1 U9123 ( .A(n18613), .ZN(n18612) );
  XNOR2_X1 U9124 ( .A(n9015), .B(n1864), .ZN(n9018) );
  XNOR2_X1 U9125 ( .A(n7276), .B(n8112), .ZN(n3107) );
  NAND2_X1 U9126 ( .A1(n7002), .A2(n6658), .ZN(n3111) );
  OR2_X1 U9127 ( .A1(n19105), .A2(n19107), .ZN(n19202) );
  OR2_X1 U9128 ( .A1(n10276), .A2(n10192), .ZN(n4777) );
  INV_X1 U9129 ( .A(n15198), .ZN(n3378) );
  INV_X1 U9130 ( .A(n13521), .ZN(n14052) );
  NAND2_X1 U9131 ( .A1(n16507), .A2(n3112), .ZN(n17041) );
  NAND2_X1 U9132 ( .A1(n16021), .A2(n16991), .ZN(n3114) );
  NAND2_X1 U9134 ( .A1(n10460), .A2(n10846), .ZN(n10464) );
  INV_X1 U9136 ( .A(n16867), .ZN(n18171) );
  NAND2_X1 U9137 ( .A1(n9978), .A2(n9980), .ZN(n9431) );
  NAND2_X1 U9138 ( .A1(n3120), .A2(n12713), .ZN(n12714) );
  OAI21_X1 U9139 ( .B1(n12712), .B2(n12711), .A(n12710), .ZN(n3120) );
  NOR2_X2 U9140 ( .A1(n4200), .A2(n13740), .ZN(n15318) );
  XNOR2_X1 U9141 ( .A(n3123), .B(n23239), .ZN(Ciphertext[42]) );
  INV_X1 U9142 ( .A(n11013), .ZN(n11011) );
  NAND3_X1 U9143 ( .A1(n6568), .A2(n6690), .A3(n6688), .ZN(n6067) );
  INV_X1 U9144 ( .A(n19084), .ZN(n19167) );
  OAI22_X1 U9145 ( .A1(n13339), .A2(n231), .B1(n13337), .B2(n13338), .ZN(n3126) );
  OAI21_X1 U9146 ( .B1(n4672), .B2(n7947), .A(n7656), .ZN(n4784) );
  NOR2_X1 U9147 ( .A1(n22458), .A2(n5584), .ZN(n5583) );
  NOR2_X1 U9149 ( .A1(n275), .A2(n20094), .ZN(n3127) );
  NOR2_X1 U9150 ( .A1(n23683), .A2(n3128), .ZN(Ciphertext[128]) );
  AND2_X1 U9151 ( .A1(n23684), .A2(n23685), .ZN(n3128) );
  NAND2_X1 U9154 ( .A1(n6906), .A2(n6372), .ZN(n5250) );
  NAND3_X1 U9155 ( .A1(n3130), .A2(n7583), .A3(n7312), .ZN(n5859) );
  OR2_X1 U9156 ( .A1(n10161), .A2(n10162), .ZN(n10163) );
  MUX2_X2 U9157 ( .A(n16330), .B(n16329), .S(n16328), .Z(n16979) );
  NAND4_X2 U9158 ( .A1(n15644), .A2(n15643), .A3(n15645), .A4(n15642), .ZN(
        n16921) );
  NOR2_X1 U9159 ( .A1(n404), .A2(n13274), .ZN(n4389) );
  XOR2_X1 U9160 ( .A(n18283), .B(n3073), .Z(n5374) );
  INV_X1 U9161 ( .A(n14459), .ZN(n13601) );
  OAI21_X1 U9162 ( .B1(n18721), .B2(n19501), .A(n4585), .ZN(n18846) );
  XNOR2_X1 U9163 ( .A(n5373), .B(n18286), .ZN(n18288) );
  INV_X1 U9165 ( .A(n4590), .ZN(n10771) );
  NAND2_X1 U9166 ( .A1(n7307), .A2(n7647), .ZN(n7765) );
  NAND2_X1 U9167 ( .A1(n19962), .A2(n20370), .ZN(n19963) );
  OAI21_X1 U9168 ( .B1(n7576), .B2(n7318), .A(n3548), .ZN(n3300) );
  AND2_X1 U9170 ( .A1(n9212), .A2(n9211), .ZN(n3134) );
  INV_X1 U9171 ( .A(n14360), .ZN(n13568) );
  OAI21_X1 U9172 ( .B1(n13587), .B2(n14359), .A(n13586), .ZN(n5527) );
  INV_X1 U9173 ( .A(n3461), .ZN(n5323) );
  OAI22_X1 U9174 ( .A1(n13627), .A2(n13843), .B1(n14063), .B2(n13847), .ZN(
        n14265) );
  NOR2_X1 U9175 ( .A1(n3324), .A2(n10756), .ZN(n10755) );
  NAND2_X1 U9176 ( .A1(n9301), .A2(n25043), .ZN(n8609) );
  NAND2_X1 U9177 ( .A1(n4140), .A2(n18120), .ZN(n18135) );
  NAND2_X1 U9178 ( .A1(n22583), .A2(n24559), .ZN(n3135) );
  NAND2_X1 U9179 ( .A1(n21238), .A2(n22803), .ZN(n3136) );
  NAND2_X1 U9180 ( .A1(n21237), .A2(n22799), .ZN(n3137) );
  NAND3_X1 U9181 ( .A1(n23507), .A2(n3139), .A3(n3138), .ZN(n23509) );
  NAND2_X1 U9182 ( .A1(n23504), .A2(n23531), .ZN(n3138) );
  NAND2_X1 U9183 ( .A1(n23513), .A2(n23503), .ZN(n3139) );
  NAND2_X1 U9184 ( .A1(n4950), .A2(n22919), .ZN(n4949) );
  NAND2_X1 U9185 ( .A1(n19657), .A2(n19850), .ZN(n3140) );
  XOR2_X1 U9186 ( .A(n15409), .B(n23620), .Z(n4636) );
  NAND3_X1 U9188 ( .A1(n5232), .A2(n9961), .A3(n3292), .ZN(n3216) );
  OR2_X1 U9189 ( .A1(n11174), .A2(n1338), .ZN(n11176) );
  MUX2_X1 U9190 ( .A(n7405), .B(n7406), .S(n4400), .Z(n7407) );
  NAND3_X1 U9191 ( .A1(n10262), .A2(n10729), .A3(n10481), .ZN(n10266) );
  XNOR2_X1 U9192 ( .A(n21029), .B(n21030), .ZN(n3141) );
  NAND2_X1 U9193 ( .A1(n11047), .A2(n11048), .ZN(n3145) );
  XNOR2_X2 U9194 ( .A(n8043), .B(n8042), .ZN(n9857) );
  AOI21_X1 U9197 ( .B1(n3147), .B2(n3146), .A(n23887), .ZN(Ciphertext[170]) );
  INV_X1 U9198 ( .A(n23877), .ZN(n3146) );
  NAND2_X1 U9199 ( .A1(n23878), .A2(n23879), .ZN(n3147) );
  OAI21_X1 U9200 ( .B1(n10095), .B2(n421), .A(n3148), .ZN(n9794) );
  NAND2_X1 U9201 ( .A1(n9790), .A2(n10095), .ZN(n3148) );
  INV_X1 U9202 ( .A(n5009), .ZN(n15351) );
  XNOR2_X1 U9205 ( .A(n3149), .B(n23973), .ZN(Ciphertext[183]) );
  NAND2_X1 U9206 ( .A1(n23971), .A2(n3150), .ZN(n3149) );
  XNOR2_X1 U9207 ( .A(n14634), .B(n15316), .ZN(n14556) );
  NAND2_X1 U9209 ( .A1(n7699), .A2(n7217), .ZN(n7215) );
  NAND2_X1 U9210 ( .A1(n6437), .A2(n5144), .ZN(n3153) );
  NAND2_X1 U9212 ( .A1(n24577), .A2(n7713), .ZN(n7719) );
  NAND2_X1 U9213 ( .A1(n5623), .A2(n7630), .ZN(n5622) );
  NAND2_X1 U9214 ( .A1(n23571), .A2(n23576), .ZN(n22201) );
  INV_X1 U9215 ( .A(n7698), .ZN(n7700) );
  OAI211_X1 U9216 ( .C1(n23418), .C2(n142), .A(n23402), .B(n3157), .ZN(n3156)
         );
  MUX2_X2 U9218 ( .A(n14177), .B(n14176), .S(n16204), .Z(n17227) );
  XNOR2_X1 U9220 ( .A(n3159), .B(n21661), .ZN(n21667) );
  XNOR2_X1 U9221 ( .A(n21663), .B(n21660), .ZN(n3159) );
  OAI21_X1 U9222 ( .B1(n25299), .B2(n22243), .A(n3160), .ZN(n22183) );
  NAND2_X1 U9223 ( .A1(n1336), .A2(n22243), .ZN(n3160) );
  XNOR2_X1 U9224 ( .A(n3162), .B(n21469), .ZN(n4657) );
  XNOR2_X1 U9225 ( .A(n21306), .B(n23798), .ZN(n3162) );
  INV_X1 U9226 ( .A(n3811), .ZN(n3810) );
  NAND2_X1 U9227 ( .A1(n19592), .A2(n19587), .ZN(n19251) );
  OR2_X2 U9228 ( .A1(n11723), .A2(n5174), .ZN(n11806) );
  NAND2_X1 U9229 ( .A1(n9523), .A2(n25207), .ZN(n4586) );
  OR3_X1 U9230 ( .A1(n17464), .A2(n17463), .A3(n16499), .ZN(n4970) );
  OR2_X1 U9232 ( .A1(n7247), .A2(n7855), .ZN(n7248) );
  OAI21_X1 U9233 ( .B1(n16943), .B2(n17613), .A(n16941), .ZN(n16944) );
  NAND3_X1 U9234 ( .A1(n16304), .A2(n16023), .A3(n15773), .ZN(n15022) );
  XNOR2_X1 U9235 ( .A(n8268), .B(n8269), .ZN(n3307) );
  NAND2_X1 U9237 ( .A1(n400), .A2(n13336), .ZN(n5505) );
  NAND2_X1 U9239 ( .A1(n6650), .A2(n7007), .ZN(n6834) );
  NAND3_X1 U9240 ( .A1(n11057), .A2(n11054), .A3(n11499), .ZN(n3163) );
  OAI211_X2 U9241 ( .C1(n13993), .C2(n14233), .A(n13377), .B(n13376), .ZN(
        n15431) );
  OAI22_X1 U9243 ( .A1(n10016), .A2(n25007), .B1(n10015), .B2(n25475), .ZN(
        n3166) );
  NAND2_X1 U9244 ( .A1(n7224), .A2(n7676), .ZN(n4376) );
  NAND2_X1 U9245 ( .A1(n10116), .A2(n10113), .ZN(n9808) );
  XNOR2_X2 U9246 ( .A(n12204), .B(n12205), .ZN(n12856) );
  NAND2_X1 U9247 ( .A1(n1149), .A2(n6975), .ZN(n6979) );
  AND2_X2 U9248 ( .A1(n20162), .A2(n20161), .ZN(n21577) );
  NAND2_X1 U9249 ( .A1(n3168), .A2(n13593), .ZN(n13594) );
  OAI21_X1 U9250 ( .B1(n14335), .B2(n25197), .A(n13877), .ZN(n3168) );
  NAND2_X1 U9251 ( .A1(n3854), .A2(n17254), .ZN(n3169) );
  XNOR2_X1 U9252 ( .A(n3170), .B(n10917), .ZN(n12510) );
  XNOR2_X1 U9253 ( .A(n12354), .B(n11639), .ZN(n3170) );
  NAND2_X1 U9254 ( .A1(n24935), .A2(n16349), .ZN(n15888) );
  INV_X1 U9255 ( .A(n7292), .ZN(n5015) );
  OR2_X1 U9258 ( .A1(n24512), .A2(n12540), .ZN(n4946) );
  NAND2_X1 U9260 ( .A1(n3172), .A2(n13103), .ZN(n13106) );
  OAI22_X1 U9261 ( .A1(n13185), .A2(n13102), .B1(n13101), .B2(n3958), .ZN(
        n3172) );
  OAI211_X1 U9265 ( .C1(n6528), .C2(n6255), .A(n6947), .B(n4757), .ZN(n4756)
         );
  OAI22_X2 U9266 ( .A1(n12332), .A2(n12331), .B1(n5625), .B2(n12350), .ZN(
        n13901) );
  XNOR2_X1 U9267 ( .A(n11564), .B(n12297), .ZN(n12028) );
  XNOR2_X1 U9269 ( .A(n14885), .B(n14886), .ZN(n15922) );
  XNOR2_X1 U9270 ( .A(n14880), .B(n14879), .ZN(n14881) );
  OR2_X1 U9271 ( .A1(n6645), .A2(n6076), .ZN(n3173) );
  INV_X1 U9272 ( .A(n9500), .ZN(n4137) );
  NAND2_X1 U9273 ( .A1(n16894), .A2(n16895), .ZN(n4612) );
  INV_X1 U9274 ( .A(n18540), .ZN(n17595) );
  XOR2_X1 U9275 ( .A(n8519), .B(n8518), .Z(n4138) );
  NAND3_X1 U9276 ( .A1(n3174), .A2(n8022), .A3(n8021), .ZN(n7746) );
  NAND2_X1 U9277 ( .A1(n17085), .A2(n17086), .ZN(n17089) );
  NAND2_X1 U9278 ( .A1(n5280), .A2(n25473), .ZN(n19024) );
  NAND2_X1 U9279 ( .A1(n313), .A2(n6651), .ZN(n6653) );
  NAND2_X1 U9280 ( .A1(n3175), .A2(n23464), .ZN(n22865) );
  OAI21_X1 U9281 ( .B1(n24364), .B2(n23016), .A(n23015), .ZN(n3175) );
  INV_X1 U9282 ( .A(n22864), .ZN(n3176) );
  OAI21_X1 U9283 ( .B1(n3177), .B2(n15539), .A(n16051), .ZN(n15309) );
  NOR2_X1 U9284 ( .A1(n4541), .A2(n16048), .ZN(n3177) );
  NOR2_X1 U9285 ( .A1(n14245), .A2(n13935), .ZN(n14243) );
  XNOR2_X1 U9286 ( .A(n11915), .B(n2145), .ZN(n11799) );
  NAND3_X1 U9288 ( .A1(n6985), .A2(n1130), .A3(n7898), .ZN(n7900) );
  XNOR2_X1 U9289 ( .A(n3179), .B(n21641), .ZN(n21643) );
  XNOR2_X1 U9290 ( .A(n21675), .B(n21638), .ZN(n3179) );
  AOI21_X1 U9291 ( .B1(n3180), .B2(n22724), .A(n22938), .ZN(n22726) );
  NAND2_X1 U9292 ( .A1(n22723), .A2(n22722), .ZN(n3180) );
  NAND3_X1 U9293 ( .A1(n23011), .A2(n23479), .A3(n23480), .ZN(n3181) );
  NOR2_X1 U9294 ( .A1(n20598), .A2(n20427), .ZN(n20425) );
  OAI211_X2 U9295 ( .C1(n7716), .C2(n7561), .A(n7560), .B(n7559), .ZN(n8880)
         );
  NAND2_X1 U9297 ( .A1(n9651), .A2(n9652), .ZN(n9656) );
  NAND4_X2 U9299 ( .A1(n9656), .A2(n9655), .A3(n3185), .A4(n9654), .ZN(n11199)
         );
  NAND2_X1 U9300 ( .A1(n9653), .A2(n10008), .ZN(n3185) );
  MUX2_X1 U9302 ( .A(n12853), .B(n12587), .S(n12854), .Z(n12589) );
  XNOR2_X2 U9303 ( .A(n12188), .B(n12187), .ZN(n12854) );
  INV_X1 U9304 ( .A(n16269), .ZN(n3186) );
  NAND2_X1 U9305 ( .A1(n16004), .A2(n16268), .ZN(n3187) );
  AOI21_X1 U9306 ( .B1(n23386), .B2(n22032), .A(n22031), .ZN(n22041) );
  OAI22_X1 U9307 ( .A1(n23033), .A2(n24972), .B1(n23034), .B2(n23830), .ZN(
        n23035) );
  NAND2_X1 U9308 ( .A1(n12758), .A2(n12784), .ZN(n12761) );
  NAND2_X1 U9309 ( .A1(n5832), .A2(n6885), .ZN(n3188) );
  XNOR2_X1 U9311 ( .A(n17984), .B(n17985), .ZN(n19381) );
  NAND2_X1 U9312 ( .A1(n10059), .A2(n10665), .ZN(n3191) );
  OR2_X1 U9313 ( .A1(n12928), .A2(n12897), .ZN(n13281) );
  XNOR2_X1 U9314 ( .A(n8950), .B(n8949), .ZN(n9550) );
  NAND2_X1 U9315 ( .A1(n6259), .A2(n24592), .ZN(n5867) );
  XNOR2_X1 U9316 ( .A(n3193), .B(n8249), .ZN(n6048) );
  XNOR2_X1 U9317 ( .A(n9175), .B(n5930), .ZN(n3193) );
  NAND3_X2 U9318 ( .A1(n16728), .A2(n3816), .A3(n16729), .ZN(n4250) );
  XNOR2_X1 U9319 ( .A(n3194), .B(n15183), .ZN(n15186) );
  XNOR2_X1 U9320 ( .A(n15184), .B(n21169), .ZN(n3194) );
  INV_X1 U9321 ( .A(n11031), .ZN(n11100) );
  NAND2_X1 U9322 ( .A1(n3196), .A2(n4739), .ZN(n4738) );
  XNOR2_X1 U9324 ( .A(n18451), .B(n3197), .ZN(n17701) );
  XNOR2_X2 U9325 ( .A(Key[123]), .B(Plaintext[123]), .ZN(n7008) );
  OAI21_X1 U9326 ( .B1(n7891), .B2(n7890), .A(n7889), .ZN(n5054) );
  NAND2_X1 U9328 ( .A1(n9804), .A2(n9805), .ZN(n10115) );
  NAND2_X1 U9329 ( .A1(n3199), .A2(n10113), .ZN(n5197) );
  NAND2_X1 U9330 ( .A1(n10115), .A2(n9533), .ZN(n3199) );
  NAND3_X1 U9331 ( .A1(n3200), .A2(n13176), .A3(n10360), .ZN(n12726) );
  NAND3_X1 U9332 ( .A1(n13177), .A2(n13178), .A3(n3200), .ZN(n13179) );
  INV_X1 U9333 ( .A(n12652), .ZN(n3200) );
  NOR2_X1 U9334 ( .A1(n22043), .A2(n3201), .ZN(n22044) );
  NAND3_X1 U9335 ( .A1(n21837), .A2(n24983), .A3(n4533), .ZN(n21900) );
  OR2_X1 U9337 ( .A1(n19389), .A2(n19386), .ZN(n3202) );
  NAND2_X1 U9339 ( .A1(n19388), .A2(n19389), .ZN(n3203) );
  XNOR2_X2 U9340 ( .A(n17719), .B(n17718), .ZN(n19389) );
  XNOR2_X1 U9342 ( .A(n12133), .B(n3207), .ZN(n3205) );
  OAI21_X1 U9346 ( .B1(n24881), .B2(n22973), .A(n22387), .ZN(n3211) );
  NOR2_X1 U9347 ( .A1(n3213), .A2(n22977), .ZN(n3212) );
  OR2_X1 U9349 ( .A1(n18952), .A2(n24441), .ZN(n3215) );
  NAND2_X1 U9350 ( .A1(n3217), .A2(n3216), .ZN(n11004) );
  NAND2_X1 U9351 ( .A1(n7572), .A2(n8140), .ZN(n3217) );
  MUX2_X1 U9352 ( .A(n17472), .B(n17633), .S(n16901), .Z(n16793) );
  INV_X1 U9353 ( .A(n19135), .ZN(n18949) );
  NAND2_X1 U9354 ( .A1(n3218), .A2(n19304), .ZN(n19135) );
  INV_X1 U9355 ( .A(n19133), .ZN(n3218) );
  NAND2_X1 U9358 ( .A1(n4327), .A2(n3221), .ZN(n3220) );
  NAND2_X1 U9359 ( .A1(n399), .A2(n12956), .ZN(n13339) );
  OAI21_X1 U9361 ( .B1(n16400), .B2(n3223), .A(n15972), .ZN(n3222) );
  NOR2_X1 U9362 ( .A1(n17453), .A2(n5072), .ZN(n17454) );
  AOI22_X2 U9363 ( .A1(n3225), .A2(n16368), .B1(n3224), .B2(n17180), .ZN(
        n17450) );
  NAND2_X1 U9364 ( .A1(n3299), .A2(n16367), .ZN(n3224) );
  NAND2_X1 U9365 ( .A1(n16365), .A2(n16366), .ZN(n3225) );
  NAND2_X1 U9366 ( .A1(n3229), .A2(n3231), .ZN(n3228) );
  OAI21_X1 U9367 ( .B1(n22233), .B2(n22234), .A(n3230), .ZN(n3229) );
  XNOR2_X1 U9368 ( .A(n3232), .B(n15191), .ZN(n13928) );
  XNOR2_X1 U9369 ( .A(n15374), .B(n3234), .ZN(n15377) );
  OAI211_X2 U9370 ( .C1(n3238), .C2(n8014), .A(n3237), .B(n3235), .ZN(n9035)
         );
  NAND3_X1 U9371 ( .A1(n7749), .A2(n8014), .A3(n25451), .ZN(n3237) );
  INV_X1 U9372 ( .A(n19851), .ZN(n3240) );
  OR2_X1 U9373 ( .A1(n18847), .A2(n19334), .ZN(n3239) );
  NAND2_X1 U9374 ( .A1(n13486), .A2(n14000), .ZN(n12678) );
  AOI21_X1 U9375 ( .B1(n299), .B2(n13485), .A(n14000), .ZN(n13490) );
  NAND2_X1 U9376 ( .A1(n13262), .A2(n14000), .ZN(n4226) );
  XNOR2_X1 U9377 ( .A(n11644), .B(n11643), .ZN(n12440) );
  INV_X1 U9378 ( .A(n12440), .ZN(n13162) );
  NAND3_X1 U9381 ( .A1(n5347), .A2(n5350), .A3(n1480), .ZN(n5349) );
  NAND2_X1 U9383 ( .A1(n5106), .A2(n5621), .ZN(n3243) );
  AND3_X2 U9386 ( .A1(n3247), .A2(n3246), .A3(n4120), .ZN(n10558) );
  NAND2_X1 U9387 ( .A1(n9592), .A2(n10160), .ZN(n3246) );
  NAND2_X1 U9388 ( .A1(n10164), .A2(n10163), .ZN(n3247) );
  NAND2_X1 U9389 ( .A1(n3249), .A2(n9066), .ZN(n3248) );
  INV_X1 U9390 ( .A(n12028), .ZN(n12029) );
  OR2_X1 U9391 ( .A1(n10939), .A2(n24591), .ZN(n3250) );
  NAND2_X1 U9392 ( .A1(n3253), .A2(n3386), .ZN(n3251) );
  NAND2_X1 U9393 ( .A1(n10313), .A2(n11168), .ZN(n3253) );
  NAND2_X1 U9394 ( .A1(n12955), .A2(n13330), .ZN(n3255) );
  XNOR2_X2 U9395 ( .A(n12035), .B(n12034), .ZN(n13323) );
  XNOR2_X2 U9396 ( .A(n18107), .B(n18108), .ZN(n19112) );
  XNOR2_X1 U9397 ( .A(n4679), .B(n18133), .ZN(n19608) );
  AOI21_X1 U9399 ( .B1(n3263), .B2(n8497), .A(n9310), .ZN(n3262) );
  NAND2_X1 U9400 ( .A1(n9998), .A2(n25453), .ZN(n3263) );
  AOI21_X2 U9401 ( .B1(n3264), .B2(n22958), .A(n22861), .ZN(n23416) );
  NAND3_X1 U9403 ( .A1(n9658), .A2(n9747), .A3(n24535), .ZN(n9663) );
  NAND2_X1 U9404 ( .A1(n24577), .A2(n8370), .ZN(n7841) );
  MUX2_X1 U9405 ( .A(n24878), .B(n7713), .S(n8368), .Z(n3267) );
  XNOR2_X1 U9407 ( .A(n12275), .B(n3269), .ZN(n11167) );
  NAND2_X1 U9408 ( .A1(n3271), .A2(n3270), .ZN(n16222) );
  NAND3_X1 U9409 ( .A1(n389), .A2(n16220), .A3(n16460), .ZN(n3270) );
  XNOR2_X1 U9412 ( .A(n8731), .B(n8421), .ZN(n8425) );
  OAI21_X1 U9414 ( .B1(n7479), .B2(n7954), .A(n7478), .ZN(n3272) );
  NAND3_X1 U9415 ( .A1(n6756), .A2(n3276), .A3(n5805), .ZN(n3273) );
  NAND3_X1 U9416 ( .A1(n19352), .A2(n19445), .A3(n25002), .ZN(n3277) );
  NAND2_X1 U9419 ( .A1(n3281), .A2(n23714), .ZN(n22084) );
  NOR2_X1 U9420 ( .A1(n23727), .A2(n22082), .ZN(n3281) );
  NAND3_X1 U9421 ( .A1(n23705), .A2(n23715), .A3(n3283), .ZN(n23706) );
  AOI21_X1 U9422 ( .B1(n23698), .B2(n3283), .A(n3282), .ZN(n23709) );
  NAND3_X1 U9423 ( .A1(n22147), .A2(n22148), .A3(n3283), .ZN(n4863) );
  NAND2_X1 U9425 ( .A1(n12885), .A2(n13224), .ZN(n3286) );
  NAND2_X1 U9426 ( .A1(n13292), .A2(n13291), .ZN(n3287) );
  MUX2_X1 U9427 ( .A(n12827), .B(n13291), .S(n12824), .Z(n12825) );
  NAND3_X1 U9428 ( .A1(n24482), .A2(n16191), .A3(n16328), .ZN(n3288) );
  NAND2_X1 U9429 ( .A1(n3291), .A2(n3290), .ZN(n3289) );
  OAI211_X1 U9430 ( .C1(n9349), .C2(n9850), .A(n3294), .B(n3305), .ZN(n3293)
         );
  NAND2_X1 U9431 ( .A1(n9349), .A2(n9384), .ZN(n3294) );
  NAND2_X1 U9432 ( .A1(n9383), .A2(n9592), .ZN(n3295) );
  NAND2_X1 U9433 ( .A1(n18987), .A2(n3296), .ZN(n3297) );
  XNOR2_X2 U9434 ( .A(n17904), .B(n17903), .ZN(n19500) );
  NAND2_X1 U9435 ( .A1(n13728), .A2(n24588), .ZN(n3298) );
  NAND2_X1 U9436 ( .A1(n15640), .A2(n16206), .ZN(n3299) );
  NAND2_X1 U9438 ( .A1(n3300), .A2(n7575), .ZN(n7457) );
  NAND2_X1 U9439 ( .A1(n3303), .A2(n3301), .ZN(n14826) );
  NAND2_X1 U9441 ( .A1(n3304), .A2(n13952), .ZN(n14157) );
  NAND2_X1 U9442 ( .A1(n5080), .A2(n13775), .ZN(n3304) );
  AND2_X1 U9443 ( .A1(n10728), .A2(n10482), .ZN(n11184) );
  NAND2_X1 U9444 ( .A1(n9385), .A2(n9520), .ZN(n10257) );
  NAND2_X1 U9445 ( .A1(n9386), .A2(n9832), .ZN(n10259) );
  NAND3_X1 U9446 ( .A1(n9522), .A2(n9521), .A3(n2257), .ZN(n5492) );
  NAND2_X1 U9447 ( .A1(n22390), .A2(n24881), .ZN(n3309) );
  MUX2_X1 U9448 ( .A(n20960), .B(n20961), .S(n20451), .Z(n20963) );
  OAI21_X1 U9449 ( .B1(n20451), .B2(n20159), .A(n3310), .ZN(n19945) );
  NAND2_X1 U9450 ( .A1(n20159), .A2(n20377), .ZN(n3310) );
  NAND2_X1 U9451 ( .A1(n3313), .A2(n10595), .ZN(n3312) );
  NAND2_X1 U9452 ( .A1(n10425), .A2(n2311), .ZN(n3313) );
  INV_X1 U9453 ( .A(n12530), .ZN(n3314) );
  NAND3_X1 U9455 ( .A1(n12773), .A2(n12471), .A3(n12470), .ZN(n3315) );
  NAND2_X1 U9457 ( .A1(n16327), .A2(n16197), .ZN(n3318) );
  NAND2_X1 U9458 ( .A1(n16196), .A2(n16195), .ZN(n3319) );
  NAND2_X1 U9459 ( .A1(n3321), .A2(n6652), .ZN(n3320) );
  MUX2_X1 U9460 ( .A(n6895), .B(n6651), .S(n6358), .Z(n3321) );
  NAND2_X1 U9461 ( .A1(n6895), .A2(n6086), .ZN(n6357) );
  XNOR2_X2 U9462 ( .A(n18593), .B(n18592), .ZN(n19418) );
  NAND2_X1 U9463 ( .A1(n9374), .A2(n3324), .ZN(n9375) );
  NAND2_X1 U9464 ( .A1(n3325), .A2(n4909), .ZN(n21481) );
  NAND2_X1 U9465 ( .A1(n25388), .A2(n20109), .ZN(n19885) );
  NAND2_X1 U9466 ( .A1(n3327), .A2(n12865), .ZN(n4181) );
  INV_X1 U9467 ( .A(n12272), .ZN(n3327) );
  NAND2_X1 U9468 ( .A1(n3330), .A2(n14166), .ZN(n3329) );
  MUX2_X1 U9469 ( .A(n13744), .B(n14165), .S(n13742), .Z(n3330) );
  NOR2_X2 U9470 ( .A1(n12449), .A2(n12448), .ZN(n13742) );
  XNOR2_X1 U9472 ( .A(n12113), .B(n12114), .ZN(n12115) );
  XNOR2_X1 U9474 ( .A(n19832), .B(n19833), .ZN(n21847) );
  INV_X1 U9475 ( .A(n21847), .ZN(n3336) );
  OAI21_X1 U9476 ( .B1(n21848), .B2(n22686), .A(n3335), .ZN(n21850) );
  NAND2_X1 U9477 ( .A1(n3336), .A2(n21848), .ZN(n3335) );
  INV_X1 U9478 ( .A(n3339), .ZN(n3337) );
  AND2_X1 U9479 ( .A1(n14205), .A2(n3341), .ZN(n3340) );
  OR2_X2 U9480 ( .A1(n12962), .A2(n12961), .ZN(n3341) );
  NAND2_X1 U9481 ( .A1(n25209), .A2(n13931), .ZN(n14247) );
  NAND2_X1 U9482 ( .A1(n4059), .A2(n4057), .ZN(n3342) );
  NAND2_X1 U9483 ( .A1(n4057), .A2(n24573), .ZN(n3343) );
  NAND2_X1 U9484 ( .A1(n414), .A2(n11207), .ZN(n10633) );
  INV_X1 U9485 ( .A(n7449), .ZN(n3348) );
  INV_X1 U9486 ( .A(n25253), .ZN(n3347) );
  NAND3_X1 U9487 ( .A1(n3346), .A2(n7635), .A3(n6486), .ZN(n3345) );
  NAND2_X1 U9488 ( .A1(n13983), .A2(n13982), .ZN(n3349) );
  NAND2_X1 U9489 ( .A1(n13984), .A2(n13922), .ZN(n3350) );
  MUX2_X1 U9491 ( .A(n13225), .B(n13226), .S(n24490), .Z(n3351) );
  NAND2_X1 U9492 ( .A1(n14221), .A2(n14222), .ZN(n3353) );
  NAND2_X1 U9493 ( .A1(n3357), .A2(n11754), .ZN(n3356) );
  NAND2_X1 U9494 ( .A1(n13009), .A2(n24965), .ZN(n3357) );
  NAND3_X1 U9495 ( .A1(n19446), .A2(n19452), .A3(n19445), .ZN(n19356) );
  INV_X1 U9497 ( .A(n4672), .ZN(n3358) );
  OAI211_X2 U9498 ( .C1(n3359), .C2(n6931), .A(n6929), .B(n6930), .ZN(n8897)
         );
  XNOR2_X1 U9499 ( .A(n11420), .B(n3361), .ZN(n3360) );
  NAND2_X1 U9500 ( .A1(n3362), .A2(n7474), .ZN(n7066) );
  NOR2_X1 U9501 ( .A1(n3362), .A2(n7421), .ZN(n7954) );
  NAND2_X1 U9502 ( .A1(n7423), .A2(n3362), .ZN(n7220) );
  NAND2_X1 U9503 ( .A1(n7477), .A2(n7475), .ZN(n3363) );
  NAND2_X1 U9504 ( .A1(n1380), .A2(n7573), .ZN(n3365) );
  NAND2_X1 U9505 ( .A1(n3366), .A2(n7580), .ZN(n7319) );
  NAND3_X1 U9506 ( .A1(n3366), .A2(n7580), .A3(n7575), .ZN(n4347) );
  NAND2_X1 U9507 ( .A1(n5809), .A2(n3366), .ZN(n5815) );
  NAND2_X1 U9508 ( .A1(n10005), .A2(n10007), .ZN(n9723) );
  INV_X1 U9510 ( .A(n9481), .ZN(n10005) );
  NAND3_X1 U9511 ( .A1(n14317), .A2(n14458), .A3(n14319), .ZN(n3367) );
  NAND2_X1 U9512 ( .A1(n13868), .A2(n13500), .ZN(n3368) );
  XNOR2_X1 U9514 ( .A(n15177), .B(n14815), .ZN(n14402) );
  NAND2_X1 U9515 ( .A1(n5522), .A2(n3371), .ZN(n15998) );
  NOR2_X1 U9516 ( .A1(n17043), .A2(n3374), .ZN(n17576) );
  AOI22_X1 U9517 ( .A1(n17372), .A2(n3371), .B1(n17373), .B2(n3374), .ZN(
        n17374) );
  AOI22_X1 U9518 ( .A1(n16678), .A2(n3374), .B1(n17572), .B2(n16677), .ZN(
        n16679) );
  OAI211_X1 U9519 ( .C1(n16767), .C2(n3374), .A(n3373), .B(n3372), .ZN(n18233)
         );
  NAND2_X1 U9520 ( .A1(n16766), .A2(n3374), .ZN(n3373) );
  OR2_X2 U9521 ( .A1(n15964), .A2(n15963), .ZN(n5522) );
  NAND3_X1 U9522 ( .A1(n1055), .A2(n11092), .A3(n11302), .ZN(n3375) );
  OAI211_X1 U9523 ( .C1(n11302), .C2(n9536), .A(n3375), .B(n1056), .ZN(n9537)
         );
  INV_X1 U9524 ( .A(n16708), .ZN(n3377) );
  NAND2_X1 U9525 ( .A1(n1473), .A2(n16708), .ZN(n3376) );
  NAND3_X1 U9527 ( .A1(n16615), .A2(n17296), .A3(n3377), .ZN(n15731) );
  NAND2_X1 U9528 ( .A1(n3378), .A2(n25410), .ZN(n16009) );
  OAI21_X1 U9529 ( .B1(n16315), .B2(n3378), .A(n16311), .ZN(n15768) );
  OAI21_X1 U9530 ( .B1(n16309), .B2(n3378), .A(n3554), .ZN(n16314) );
  AOI21_X1 U9531 ( .B1(n15752), .B2(n3378), .A(n16312), .ZN(n15753) );
  NAND3_X1 U9532 ( .A1(n19390), .A2(n19630), .A3(n24909), .ZN(n3379) );
  OAI21_X1 U9533 ( .B1(n16206), .B2(n3380), .A(n17182), .ZN(n14177) );
  OR2_X1 U9534 ( .A1(n16367), .A2(n15640), .ZN(n17182) );
  NAND3_X1 U9535 ( .A1(n16367), .A2(n17180), .A3(n3380), .ZN(n15910) );
  NAND3_X1 U9537 ( .A1(n13529), .A2(n3382), .A3(n3381), .ZN(n14892) );
  OAI21_X1 U9538 ( .B1(n12445), .B2(n3383), .A(n13526), .ZN(n3382) );
  XNOR2_X1 U9539 ( .A(n11957), .B(n11959), .ZN(n12320) );
  NAND2_X1 U9540 ( .A1(n11169), .A2(n11168), .ZN(n11174) );
  NAND3_X1 U9541 ( .A1(n3386), .A2(n11175), .A3(n24591), .ZN(n3385) );
  NAND3_X1 U9542 ( .A1(n3387), .A2(n10586), .A3(n10587), .ZN(n10593) );
  NAND2_X1 U9543 ( .A1(n10582), .A2(n10583), .ZN(n3387) );
  NAND3_X1 U9544 ( .A1(n18037), .A2(n19602), .A3(n19596), .ZN(n3389) );
  NAND2_X1 U9545 ( .A1(n16577), .A2(n17131), .ZN(n3392) );
  NAND2_X1 U9546 ( .A1(n5337), .A2(n3393), .ZN(n19248) );
  NAND2_X1 U9547 ( .A1(n3394), .A2(n19575), .ZN(n3393) );
  INV_X1 U9548 ( .A(n19578), .ZN(n3394) );
  NAND2_X1 U9549 ( .A1(n25072), .A2(n19248), .ZN(n4425) );
  XNOR2_X1 U9550 ( .A(n17592), .B(n18283), .ZN(n3397) );
  NAND3_X1 U9551 ( .A1(n4774), .A2(n16375), .A3(n16262), .ZN(n3395) );
  NAND2_X1 U9552 ( .A1(n16089), .A2(n17165), .ZN(n3396) );
  XNOR2_X1 U9553 ( .A(n3397), .B(n18375), .ZN(n18044) );
  XNOR2_X1 U9554 ( .A(n3398), .B(n1466), .ZN(n9365) );
  XNOR2_X1 U9555 ( .A(n9137), .B(n9138), .ZN(n3398) );
  INV_X1 U9557 ( .A(n14320), .ZN(n3402) );
  INV_X1 U9558 ( .A(n14321), .ZN(n3404) );
  NAND2_X1 U9560 ( .A1(n3402), .A2(n3401), .ZN(n3400) );
  NAND2_X1 U9561 ( .A1(n3404), .A2(n14320), .ZN(n3403) );
  NAND2_X1 U9562 ( .A1(n9382), .A2(n10162), .ZN(n3405) );
  NAND2_X1 U9563 ( .A1(n15933), .A2(n16231), .ZN(n3406) );
  NAND3_X1 U9564 ( .A1(n17662), .A2(n3131), .A3(n17661), .ZN(n16969) );
  NAND3_X1 U9565 ( .A1(n16105), .A2(n25409), .A3(n3410), .ZN(n3408) );
  INV_X1 U9566 ( .A(n16102), .ZN(n3410) );
  NAND2_X1 U9568 ( .A1(n22800), .A2(n22798), .ZN(n3411) );
  XNOR2_X2 U9569 ( .A(n21197), .B(n21196), .ZN(n22803) );
  INV_X1 U9571 ( .A(n3414), .ZN(n6892) );
  OR2_X1 U9572 ( .A1(n6651), .A2(n6893), .ZN(n3413) );
  NAND3_X1 U9573 ( .A1(n24345), .A2(n10302), .A3(n2386), .ZN(n3415) );
  NAND3_X1 U9574 ( .A1(n3419), .A2(n19254), .A3(n25001), .ZN(n5027) );
  NAND2_X1 U9575 ( .A1(n25244), .A2(n19596), .ZN(n3419) );
  NOR2_X1 U9576 ( .A1(n3419), .A2(n18870), .ZN(n18873) );
  OAI21_X1 U9577 ( .B1(n5561), .B2(n3421), .A(n13051), .ZN(n3420) );
  NOR2_X1 U9578 ( .A1(n25408), .A2(n13049), .ZN(n3421) );
  AND2_X1 U9579 ( .A1(n4850), .A2(n13050), .ZN(n5561) );
  NOR2_X1 U9580 ( .A1(n13049), .A2(n12490), .ZN(n3423) );
  NAND2_X1 U9581 ( .A1(n13968), .A2(n13969), .ZN(n3427) );
  NAND2_X1 U9582 ( .A1(n3767), .A2(n3428), .ZN(n5764) );
  INV_X1 U9583 ( .A(n3767), .ZN(n3429) );
  MUX2_X1 U9585 ( .A(n17050), .B(n17049), .S(n17048), .Z(n3432) );
  NAND2_X1 U9586 ( .A1(n3435), .A2(n3434), .ZN(n3433) );
  NAND2_X1 U9587 ( .A1(n17053), .A2(n17048), .ZN(n17052) );
  NAND2_X1 U9588 ( .A1(n24162), .A2(n16016), .ZN(n15941) );
  NAND2_X1 U9589 ( .A1(n24162), .A2(n3436), .ZN(n3437) );
  AND2_X1 U9590 ( .A1(n16246), .A2(n16016), .ZN(n3436) );
  NAND3_X1 U9592 ( .A1(n392), .A2(n13080), .A3(n13081), .ZN(n13559) );
  AOI21_X1 U9593 ( .B1(n24984), .B2(n9384), .A(n3438), .ZN(n9854) );
  AND2_X1 U9594 ( .A1(n9348), .A2(n10158), .ZN(n3438) );
  NAND2_X1 U9597 ( .A1(n12719), .A2(n13167), .ZN(n12447) );
  NAND2_X1 U9598 ( .A1(n3445), .A2(n24051), .ZN(n3444) );
  NAND2_X1 U9599 ( .A1(n24051), .A2(n24500), .ZN(n6719) );
  NAND2_X1 U9600 ( .A1(n9410), .A2(n10452), .ZN(n3446) );
  NAND2_X1 U9601 ( .A1(n9411), .A2(n10290), .ZN(n3447) );
  XNOR2_X1 U9602 ( .A(n3448), .B(n4670), .ZN(n11504) );
  XNOR2_X1 U9603 ( .A(n11504), .B(n11505), .ZN(n11508) );
  OAI22_X1 U9604 ( .A1(n4496), .A2(n24841), .B1(n16359), .B2(n3450), .ZN(n3449) );
  NAND2_X1 U9605 ( .A1(n3451), .A2(n16355), .ZN(n3450) );
  INV_X1 U9606 ( .A(n16356), .ZN(n3451) );
  INV_X1 U9607 ( .A(n1355), .ZN(n3453) );
  OAI21_X1 U9608 ( .B1(n13518), .B2(n13521), .A(n3453), .ZN(n3452) );
  NAND2_X1 U9609 ( .A1(n14050), .A2(n1355), .ZN(n3455) );
  INV_X1 U9610 ( .A(n3456), .ZN(n22055) );
  NAND2_X1 U9611 ( .A1(n336), .A2(n21829), .ZN(n3456) );
  NOR2_X1 U9613 ( .A1(n25244), .A2(n19071), .ZN(n18831) );
  NOR2_X1 U9614 ( .A1(n3461), .A2(n13094), .ZN(n13095) );
  NOR2_X1 U9615 ( .A1(n3461), .A2(n3492), .ZN(n12505) );
  NOR2_X1 U9616 ( .A1(n4405), .A2(n3461), .ZN(n10199) );
  OAI21_X1 U9617 ( .B1(n13093), .B2(n3461), .A(n3460), .ZN(n4906) );
  NAND2_X1 U9618 ( .A1(n3461), .A2(n12648), .ZN(n3460) );
  XNOR2_X1 U9619 ( .A(n25394), .B(n14816), .ZN(n14115) );
  XNOR2_X1 U9620 ( .A(n25394), .B(n15002), .ZN(n15004) );
  XNOR2_X1 U9621 ( .A(n14889), .B(n25394), .ZN(n15084) );
  NAND2_X1 U9622 ( .A1(n3464), .A2(n13788), .ZN(n3463) );
  NAND2_X1 U9623 ( .A1(n14188), .A2(n14142), .ZN(n3464) );
  INV_X1 U9625 ( .A(n19953), .ZN(n20587) );
  NAND2_X1 U9626 ( .A1(n4143), .A2(n10772), .ZN(n10910) );
  NAND2_X1 U9628 ( .A1(n7897), .A2(n3469), .ZN(n7140) );
  NAND3_X1 U9629 ( .A1(n7898), .A2(n7232), .A3(n3469), .ZN(n5236) );
  INV_X1 U9630 ( .A(n3471), .ZN(n14599) );
  NAND2_X1 U9631 ( .A1(n9211), .A2(n3472), .ZN(n9380) );
  NAND2_X1 U9632 ( .A1(n10125), .A2(n3472), .ZN(n10126) );
  NAND2_X1 U9633 ( .A1(n5057), .A2(n3472), .ZN(n9597) );
  AOI21_X1 U9634 ( .B1(n10130), .B2(n9211), .A(n3472), .ZN(n10131) );
  OAI21_X1 U9635 ( .B1(n5057), .B2(n3472), .A(n7437), .ZN(n7438) );
  INV_X1 U9636 ( .A(n13274), .ZN(n12963) );
  MUX2_X1 U9637 ( .A(n12695), .B(n404), .S(n13274), .Z(n12697) );
  NOR2_X1 U9638 ( .A1(n24967), .A2(n23220), .ZN(n3475) );
  NOR2_X1 U9639 ( .A1(n23212), .A2(n3475), .ZN(n23232) );
  NAND2_X1 U9640 ( .A1(n7991), .A2(n7993), .ZN(n7414) );
  OAI21_X2 U9641 ( .B1(n6677), .B2(n271), .A(n6676), .ZN(n7993) );
  XNOR2_X1 U9642 ( .A(n21559), .B(n2120), .ZN(n21127) );
  NAND2_X1 U9646 ( .A1(n20330), .A2(n3482), .ZN(n3481) );
  NAND2_X1 U9647 ( .A1(n18136), .A2(n20089), .ZN(n3483) );
  XNOR2_X1 U9648 ( .A(n3484), .B(n24009), .ZN(Ciphertext[189]) );
  OAI211_X1 U9649 ( .C1(n24018), .C2(n24008), .A(n3487), .B(n3485), .ZN(n3484)
         );
  NAND2_X1 U9650 ( .A1(n24008), .A2(n5773), .ZN(n3487) );
  NAND2_X1 U9651 ( .A1(n806), .A2(n3488), .ZN(n7073) );
  NAND2_X1 U9652 ( .A1(n9247), .A2(n3489), .ZN(n4594) );
  NAND2_X1 U9653 ( .A1(n9326), .A2(n9787), .ZN(n10087) );
  NAND2_X1 U9654 ( .A1(n9507), .A2(n9787), .ZN(n4208) );
  MUX2_X1 U9655 ( .A(n10080), .B(n9507), .S(n9787), .Z(n8466) );
  NAND2_X1 U9656 ( .A1(n9789), .A2(n9787), .ZN(n9307) );
  NAND3_X1 U9657 ( .A1(n3491), .A2(n19412), .A3(n19173), .ZN(n19174) );
  MUX2_X1 U9658 ( .A(n5324), .B(n5323), .S(n4405), .Z(n13098) );
  NAND2_X1 U9659 ( .A1(n15795), .A2(n15794), .ZN(n3494) );
  NAND2_X1 U9661 ( .A1(n3495), .A2(n4533), .ZN(n4953) );
  NAND2_X1 U9662 ( .A1(n4533), .A2(n22043), .ZN(n23792) );
  NAND2_X1 U9663 ( .A1(n3497), .A2(n7789), .ZN(n3496) );
  NAND2_X1 U9664 ( .A1(n7441), .A2(n7788), .ZN(n3497) );
  NAND2_X1 U9665 ( .A1(n7781), .A2(n7787), .ZN(n7441) );
  MUX2_X1 U9666 ( .A(n7579), .B(n7578), .S(n7577), .Z(n3499) );
  OAI21_X1 U9667 ( .B1(n14038), .B2(n3501), .A(n14319), .ZN(n5058) );
  AOI21_X1 U9668 ( .B1(n14461), .B2(n14460), .A(n1474), .ZN(n14463) );
  XNOR2_X1 U9669 ( .A(n11660), .B(n12391), .ZN(n10196) );
  NAND3_X1 U9671 ( .A1(n10283), .A2(n10859), .A3(n10855), .ZN(n3502) );
  NOR2_X2 U9672 ( .A1(n15798), .A2(n15787), .ZN(n17134) );
  XNOR2_X1 U9674 ( .A(n8112), .B(n8115), .ZN(n3504) );
  XNOR2_X1 U9675 ( .A(n8114), .B(n8113), .ZN(n3505) );
  NAND2_X1 U9677 ( .A1(n19206), .A2(n19381), .ZN(n3508) );
  NAND2_X1 U9679 ( .A1(n20131), .A2(n55), .ZN(n19671) );
  NAND2_X1 U9680 ( .A1(n3509), .A2(n4671), .ZN(n3511) );
  INV_X1 U9681 ( .A(n10699), .ZN(n3509) );
  NAND2_X1 U9683 ( .A1(n2754), .A2(n25233), .ZN(n3513) );
  NAND2_X1 U9684 ( .A1(n266), .A2(n17012), .ZN(n3515) );
  INV_X1 U9685 ( .A(n19094), .ZN(n18877) );
  NOR2_X2 U9686 ( .A1(n3518), .A2(n17986), .ZN(n20554) );
  OAI21_X1 U9687 ( .B1(n20518), .B2(n3519), .A(n20517), .ZN(n3520) );
  INV_X1 U9688 ( .A(n20516), .ZN(n3519) );
  NAND2_X1 U9690 ( .A1(n20273), .A2(n3522), .ZN(n3521) );
  NAND2_X1 U9691 ( .A1(n17078), .A2(n17075), .ZN(n16892) );
  XNOR2_X1 U9692 ( .A(n15170), .B(n14973), .ZN(n3525) );
  XNOR2_X2 U9693 ( .A(n3525), .B(n4115), .ZN(n16449) );
  NAND2_X1 U9694 ( .A1(n24911), .A2(n23375), .ZN(n3527) );
  XNOR2_X1 U9695 ( .A(n3526), .B(n22440), .ZN(Ciphertext[76]) );
  NAND3_X1 U9696 ( .A1(n3528), .A2(n22439), .A3(n3527), .ZN(n3526) );
  NAND3_X1 U9697 ( .A1(n18944), .A2(n19472), .A3(n19322), .ZN(n3529) );
  NAND3_X1 U9698 ( .A1(n19471), .A2(n19322), .A3(n18956), .ZN(n3530) );
  OAI22_X1 U9699 ( .A1(n11116), .A2(n3532), .B1(n11111), .B2(n10725), .ZN(
        n5335) );
  AOI21_X1 U9700 ( .B1(n6235), .B2(n5784), .A(n6232), .ZN(n5785) );
  MUX2_X1 U9701 ( .A(n6717), .B(n6716), .S(n6232), .Z(n7074) );
  NAND2_X1 U9702 ( .A1(n3533), .A2(n14064), .ZN(n13430) );
  OAI21_X1 U9703 ( .B1(n5694), .B2(n3533), .A(n5693), .ZN(n5692) );
  INV_X1 U9704 ( .A(n18073), .ZN(n17899) );
  XNOR2_X1 U9705 ( .A(n18073), .B(n3535), .ZN(n3534) );
  INV_X1 U9706 ( .A(n18523), .ZN(n3535) );
  NAND2_X1 U9709 ( .A1(n13806), .A2(n13805), .ZN(n3539) );
  NAND2_X1 U9710 ( .A1(n341), .A2(n20320), .ZN(n3540) );
  INV_X1 U9711 ( .A(n24062), .ZN(n3545) );
  NAND2_X1 U9713 ( .A1(n16171), .A2(n244), .ZN(n3547) );
  OAI21_X1 U9714 ( .B1(n3366), .B2(n7579), .A(n3548), .ZN(n4345) );
  NAND2_X1 U9715 ( .A1(n7359), .A2(n7993), .ZN(n3550) );
  OR2_X2 U9718 ( .A1(n3552), .A2(n3551), .ZN(n10411) );
  AOI21_X1 U9719 ( .B1(n9591), .B2(n9590), .A(n10168), .ZN(n3552) );
  NAND2_X1 U9721 ( .A1(n4677), .A2(n4676), .ZN(n3556) );
  XNOR2_X1 U9722 ( .A(n14907), .B(n23523), .ZN(n14413) );
  AND2_X1 U9723 ( .A1(n14240), .A2(n25209), .ZN(n3557) );
  NAND2_X1 U9724 ( .A1(n12805), .A2(n13017), .ZN(n3559) );
  OR2_X1 U9727 ( .A1(n12669), .A2(n3561), .ZN(n12671) );
  NOR2_X1 U9728 ( .A1(n12668), .A2(n13488), .ZN(n3561) );
  AND2_X1 U9729 ( .A1(n299), .A2(n12669), .ZN(n13667) );
  OR2_X1 U9730 ( .A1(n12669), .A2(n299), .ZN(n5221) );
  NAND2_X1 U9732 ( .A1(n14001), .A2(n3562), .ZN(n14007) );
  OAI21_X1 U9733 ( .B1(n23320), .B2(n23317), .A(n3564), .ZN(n21895) );
  MUX2_X1 U9734 ( .A(n23311), .B(n24316), .S(n23326), .Z(n22384) );
  OR2_X2 U9735 ( .A1(n21877), .A2(n21876), .ZN(n23326) );
  XNOR2_X1 U9736 ( .A(n11628), .B(n445), .ZN(n3565) );
  INV_X1 U9737 ( .A(n7516), .ZN(n7404) );
  NAND2_X1 U9741 ( .A1(n3571), .A2(n3570), .ZN(n3569) );
  NAND2_X1 U9742 ( .A1(n7554), .A2(n7863), .ZN(n3572) );
  INV_X1 U9743 ( .A(n6922), .ZN(n4042) );
  XNOR2_X2 U9744 ( .A(Key[167]), .B(Plaintext[167]), .ZN(n6198) );
  NAND2_X1 U9745 ( .A1(n11000), .A2(n3573), .ZN(n11001) );
  INV_X1 U9746 ( .A(n10907), .ZN(n10747) );
  NAND2_X1 U9747 ( .A1(n10902), .A2(n10907), .ZN(n3574) );
  INV_X1 U9748 ( .A(n10751), .ZN(n10902) );
  NAND2_X1 U9749 ( .A1(n10747), .A2(n10746), .ZN(n3575) );
  NAND3_X1 U9750 ( .A1(n25409), .A2(n16101), .A3(n5100), .ZN(n3592) );
  INV_X1 U9753 ( .A(n14625), .ZN(n16038) );
  AND3_X2 U9754 ( .A1(n3580), .A2(n3584), .A3(n3579), .ZN(n20071) );
  NAND2_X1 U9755 ( .A1(n3581), .A2(n19470), .ZN(n3580) );
  NAND2_X1 U9757 ( .A1(n22564), .A2(n21934), .ZN(n22132) );
  AOI22_X1 U9759 ( .A1(n22297), .A2(n25373), .B1(n3586), .B2(n3585), .ZN(
        Ciphertext[44]) );
  NAND2_X1 U9760 ( .A1(n22294), .A2(n189), .ZN(n3585) );
  NAND2_X1 U9761 ( .A1(n3588), .A2(n7531), .ZN(n3708) );
  NAND2_X1 U9762 ( .A1(n3590), .A2(n12707), .ZN(n12429) );
  NAND2_X1 U9763 ( .A1(n13078), .A2(n24573), .ZN(n3589) );
  NAND3_X1 U9764 ( .A1(n12712), .A2(n12431), .A3(n3590), .ZN(n12432) );
  NAND2_X1 U9765 ( .A1(n11589), .A2(n3590), .ZN(n11594) );
  NAND2_X1 U9766 ( .A1(n24585), .A2(n17054), .ZN(n17057) );
  OAI21_X1 U9767 ( .B1(n16722), .B2(n24398), .A(n3593), .ZN(n16723) );
  NAND2_X1 U9768 ( .A1(n10814), .A2(n10967), .ZN(n3594) );
  NAND2_X1 U9769 ( .A1(n9909), .A2(n9935), .ZN(n3596) );
  NAND2_X1 U9770 ( .A1(n17023), .A2(n3598), .ZN(n3600) );
  NAND2_X1 U9771 ( .A1(n16627), .A2(n17389), .ZN(n3599) );
  XNOR2_X1 U9772 ( .A(n18261), .B(n2717), .ZN(n3605) );
  INV_X1 U9773 ( .A(n10326), .ZN(n3606) );
  NAND3_X1 U9775 ( .A1(n9814), .A2(n10169), .A3(n25046), .ZN(n9589) );
  MUX2_X1 U9776 ( .A(n9814), .B(n9817), .S(n25046), .Z(n8332) );
  NAND3_X1 U9777 ( .A1(n16324), .A2(n24482), .A3(n16197), .ZN(n16198) );
  NAND2_X1 U9778 ( .A1(n15258), .A2(n24482), .ZN(n5408) );
  INV_X1 U9779 ( .A(n8022), .ZN(n3615) );
  NOR2_X1 U9780 ( .A1(n7532), .A2(n8024), .ZN(n3611) );
  NAND2_X1 U9781 ( .A1(n3614), .A2(n7532), .ZN(n3612) );
  XNOR2_X1 U9782 ( .A(n18467), .B(n21335), .ZN(n17430) );
  XNOR2_X1 U9783 ( .A(n18467), .B(n729), .ZN(n17797) );
  XNOR2_X1 U9784 ( .A(n18467), .B(n2049), .ZN(n18153) );
  INV_X1 U9785 ( .A(n19366), .ZN(n19219) );
  OAI21_X1 U9786 ( .B1(n24424), .B2(n24361), .A(n3617), .ZN(n5682) );
  NAND2_X1 U9787 ( .A1(n24424), .A2(n19371), .ZN(n3617) );
  OR2_X1 U9788 ( .A1(n6878), .A2(n6768), .ZN(n3618) );
  NAND3_X1 U9789 ( .A1(n12917), .A2(n12612), .A3(n25248), .ZN(n11714) );
  NOR2_X1 U9791 ( .A1(n12612), .A2(n25248), .ZN(n4789) );
  NAND2_X1 U9792 ( .A1(n19060), .A2(n19059), .ZN(n3620) );
  OR2_X1 U9794 ( .A1(n22510), .A2(n23303), .ZN(n3622) );
  NAND2_X1 U9795 ( .A1(n22763), .A2(n22509), .ZN(n3624) );
  INV_X1 U9796 ( .A(n23306), .ZN(n3625) );
  NOR2_X1 U9798 ( .A1(n12508), .A2(n12652), .ZN(n3631) );
  OR2_X1 U9800 ( .A1(n13614), .A2(n13610), .ZN(n3634) );
  NAND2_X1 U9802 ( .A1(n3635), .A2(n3634), .ZN(n13616) );
  NAND2_X1 U9803 ( .A1(n13611), .A2(n13614), .ZN(n3635) );
  OAI211_X1 U9804 ( .C1(n16130), .C2(n1365), .A(n24826), .B(n3636), .ZN(n3639)
         );
  NAND2_X1 U9807 ( .A1(n3638), .A2(n15800), .ZN(n3637) );
  NOR2_X1 U9808 ( .A1(n1365), .A2(n14664), .ZN(n3638) );
  NAND2_X1 U9809 ( .A1(n7663), .A2(n7662), .ZN(n7670) );
  NAND2_X1 U9810 ( .A1(n23999), .A2(n25079), .ZN(n3641) );
  NOR2_X1 U9811 ( .A1(n23994), .A2(n25079), .ZN(n22676) );
  INV_X1 U9814 ( .A(n16670), .ZN(n3645) );
  NAND3_X1 U9817 ( .A1(n9899), .A2(n9286), .A3(n9287), .ZN(n8139) );
  NAND2_X1 U9819 ( .A1(n25021), .A2(n9898), .ZN(n9286) );
  XNOR2_X1 U9820 ( .A(n21106), .B(n23983), .ZN(n21107) );
  NAND3_X1 U9821 ( .A1(n19818), .A2(n20243), .A3(n20244), .ZN(n3650) );
  NAND2_X1 U9822 ( .A1(n3652), .A2(n3651), .ZN(n19510) );
  NAND2_X1 U9823 ( .A1(n19298), .A2(n19297), .ZN(n3651) );
  NAND2_X1 U9824 ( .A1(n19299), .A2(n3653), .ZN(n3652) );
  NAND2_X1 U9825 ( .A1(n1344), .A2(n19939), .ZN(n19818) );
  NAND2_X1 U9826 ( .A1(n9380), .A2(n9379), .ZN(n10255) );
  OR2_X1 U9827 ( .A1(n20462), .A2(n3656), .ZN(n20396) );
  NAND2_X1 U9828 ( .A1(n20393), .A2(n20394), .ZN(n3657) );
  INV_X1 U9829 ( .A(n16004), .ZN(n3658) );
  NAND2_X1 U9830 ( .A1(n3658), .A2(n15758), .ZN(n16270) );
  NOR2_X1 U9834 ( .A1(n19275), .A2(n3773), .ZN(n3661) );
  INV_X1 U9835 ( .A(n5573), .ZN(n3662) );
  OAI21_X1 U9837 ( .B1(n22358), .B2(n3664), .A(n4203), .ZN(n22045) );
  NAND2_X1 U9838 ( .A1(n21348), .A2(n21782), .ZN(n3664) );
  INV_X1 U9839 ( .A(n17300), .ZN(n16704) );
  NAND2_X1 U9840 ( .A1(n20422), .A2(n20399), .ZN(n4265) );
  AOI21_X1 U9841 ( .B1(n3667), .B2(n3666), .A(n23860), .ZN(n23855) );
  NAND3_X1 U9842 ( .A1(n23851), .A2(n3183), .A3(n24428), .ZN(n3666) );
  OR2_X1 U9843 ( .A1(n23851), .A2(n3183), .ZN(n3667) );
  NAND2_X1 U9844 ( .A1(n23839), .A2(n23862), .ZN(n23851) );
  OAI211_X1 U9845 ( .C1(n5371), .C2(n4874), .A(n3673), .B(n3672), .ZN(n3671)
         );
  NAND2_X1 U9846 ( .A1(n18747), .A2(n18923), .ZN(n3672) );
  NAND2_X1 U9847 ( .A1(n18748), .A2(n19315), .ZN(n3673) );
  OAI21_X1 U9848 ( .B1(n3674), .B2(n10064), .A(n10060), .ZN(n5609) );
  INV_X1 U9850 ( .A(n10063), .ZN(n3674) );
  NAND2_X1 U9851 ( .A1(n3676), .A2(n3675), .ZN(n7493) );
  NAND2_X1 U9852 ( .A1(n7489), .A2(n24475), .ZN(n3675) );
  NAND2_X1 U9853 ( .A1(n7947), .A2(n7942), .ZN(n7489) );
  NAND2_X1 U9855 ( .A1(n3681), .A2(n3679), .ZN(n8132) );
  NAND3_X1 U9856 ( .A1(n5015), .A2(n7754), .A3(n5202), .ZN(n3680) );
  INV_X1 U9857 ( .A(n22270), .ZN(n22324) );
  NAND4_X1 U9860 ( .A1(n15920), .A2(n3685), .A3(n17366), .A4(n3684), .ZN(n3683) );
  OR2_X1 U9861 ( .A1(n17039), .A2(n25058), .ZN(n3684) );
  NAND2_X1 U9862 ( .A1(n25058), .A2(n16770), .ZN(n17366) );
  AND2_X1 U9863 ( .A1(n13164), .A2(n1353), .ZN(n3686) );
  NAND2_X1 U9864 ( .A1(n24601), .A2(n13061), .ZN(n13164) );
  XNOR2_X2 U9866 ( .A(n20959), .B(n20958), .ZN(n22072) );
  NOR2_X1 U9867 ( .A1(n22917), .A2(n22072), .ZN(n4948) );
  INV_X1 U9868 ( .A(n12719), .ZN(n3689) );
  NAND2_X1 U9870 ( .A1(n13011), .A2(n13014), .ZN(n3691) );
  NAND2_X1 U9871 ( .A1(n19438), .A2(n361), .ZN(n19246) );
  NAND2_X1 U9872 ( .A1(n6076), .A2(n6795), .ZN(n6362) );
  NAND2_X1 U9875 ( .A1(n17370), .A2(n17369), .ZN(n3693) );
  NAND2_X1 U9876 ( .A1(n13395), .A2(n3698), .ZN(n3697) );
  NAND2_X1 U9877 ( .A1(n3700), .A2(n24995), .ZN(n3699) );
  XNOR2_X1 U9878 ( .A(n12225), .B(n20609), .ZN(n11543) );
  XNOR2_X1 U9879 ( .A(n18301), .B(n3703), .ZN(n18567) );
  XNOR2_X1 U9880 ( .A(n3703), .B(n18294), .ZN(n16946) );
  NAND2_X1 U9881 ( .A1(n13081), .A2(n13080), .ZN(n13647) );
  NOR2_X1 U9882 ( .A1(n13078), .A2(n24573), .ZN(n3704) );
  XNOR2_X1 U9884 ( .A(n3706), .B(n18233), .ZN(n18613) );
  XNOR2_X1 U9885 ( .A(n14916), .B(n14915), .ZN(n3707) );
  INV_X1 U9886 ( .A(n16030), .ZN(n4092) );
  MUX2_X1 U9887 ( .A(n16274), .B(n24403), .S(n16030), .Z(n4091) );
  NAND2_X1 U9888 ( .A1(n21841), .A2(n22252), .ZN(n22254) );
  NOR2_X1 U9891 ( .A1(n17320), .A2(n4426), .ZN(n16710) );
  NAND2_X1 U9892 ( .A1(n17079), .A2(n17075), .ZN(n17482) );
  NAND3_X1 U9894 ( .A1(n22282), .A2(n3714), .A3(n2673), .ZN(n3713) );
  NAND2_X1 U9895 ( .A1(n22947), .A2(n22946), .ZN(n3714) );
  XNOR2_X1 U9896 ( .A(n3715), .B(n2847), .ZN(n7494) );
  XNOR2_X1 U9897 ( .A(n3715), .B(n889), .ZN(n8996) );
  XNOR2_X1 U9898 ( .A(n3715), .B(n22886), .ZN(n8422) );
  XNOR2_X1 U9899 ( .A(n3715), .B(n21533), .ZN(n8629) );
  NAND3_X1 U9900 ( .A1(n3717), .A2(n1028), .A3(n14150), .ZN(n3892) );
  NAND2_X1 U9901 ( .A1(n5102), .A2(n3716), .ZN(n14032) );
  NAND2_X1 U9902 ( .A1(n13805), .A2(n3717), .ZN(n4962) );
  NAND2_X1 U9903 ( .A1(n3720), .A2(n23250), .ZN(n4072) );
  NOR2_X1 U9904 ( .A1(n23236), .A2(n25373), .ZN(n22648) );
  NAND3_X1 U9905 ( .A1(n23241), .A2(n24914), .A3(n3719), .ZN(n23244) );
  INV_X1 U9906 ( .A(n9220), .ZN(n3722) );
  NAND2_X1 U9907 ( .A1(n4806), .A2(n24586), .ZN(n3723) );
  XNOR2_X1 U9908 ( .A(n3725), .B(n921), .ZN(n4873) );
  XNOR2_X1 U9909 ( .A(n18239), .B(n3725), .ZN(n17982) );
  XNOR2_X1 U9910 ( .A(n3725), .B(n17840), .ZN(n18537) );
  XNOR2_X1 U9911 ( .A(n3725), .B(n18621), .ZN(n17261) );
  INV_X1 U9912 ( .A(n24407), .ZN(n3726) );
  AOI21_X1 U9913 ( .B1(n3727), .B2(n3726), .A(n19393), .ZN(n19399) );
  NAND2_X1 U9914 ( .A1(n25198), .A2(n13246), .ZN(n12807) );
  NAND2_X1 U9915 ( .A1(n13015), .A2(n25199), .ZN(n12561) );
  NOR2_X1 U9916 ( .A1(n10685), .A2(n4481), .ZN(n11007) );
  NAND2_X1 U9917 ( .A1(n11007), .A2(n11004), .ZN(n3728) );
  NAND2_X1 U9920 ( .A1(n3734), .A2(n3733), .ZN(n3732) );
  NOR2_X1 U9921 ( .A1(n19953), .A2(n20588), .ZN(n3733) );
  INV_X1 U9922 ( .A(n20590), .ZN(n3734) );
  INV_X1 U9923 ( .A(n16686), .ZN(n3735) );
  NAND2_X1 U9924 ( .A1(n16686), .A2(n25030), .ZN(n3736) );
  NAND3_X1 U9925 ( .A1(n17279), .A2(n17275), .A3(n17252), .ZN(n17253) );
  OAI21_X1 U9926 ( .B1(n16106), .B2(n16109), .A(n2090), .ZN(n15855) );
  XNOR2_X1 U9929 ( .A(n3738), .B(n23841), .ZN(Ciphertext[163]) );
  NAND3_X1 U9930 ( .A1(n3739), .A2(n4816), .A3(n23840), .ZN(n3738) );
  XNOR2_X1 U9931 ( .A(n17913), .B(n23602), .ZN(n16947) );
  NAND2_X1 U9932 ( .A1(n3740), .A2(n20444), .ZN(n23843) );
  OAI21_X1 U9933 ( .B1(n9340), .B2(n10148), .A(n3742), .ZN(n8225) );
  NOR2_X2 U9934 ( .A1(n12578), .A2(n12579), .ZN(n13843) );
  NAND3_X1 U9935 ( .A1(n5099), .A2(n3749), .A3(n3747), .ZN(n19697) );
  NAND2_X1 U9936 ( .A1(n19325), .A2(n19472), .ZN(n3747) );
  NOR2_X1 U9937 ( .A1(n10202), .A2(n3750), .ZN(n9411) );
  MUX2_X1 U9938 ( .A(n4733), .B(n10752), .S(n3750), .Z(n4732) );
  NAND2_X1 U9939 ( .A1(n19125), .A2(n19539), .ZN(n3752) );
  INV_X1 U9940 ( .A(n14063), .ZN(n3756) );
  AND2_X1 U9941 ( .A1(n13627), .A2(n14063), .ZN(n3754) );
  AOI21_X1 U9942 ( .B1(n3760), .B2(n3761), .A(n3758), .ZN(n3757) );
  NOR2_X1 U9944 ( .A1(n10941), .A2(n11038), .ZN(n3762) );
  NAND2_X1 U9945 ( .A1(n6939), .A2(n5908), .ZN(n3763) );
  NAND2_X1 U9946 ( .A1(n3544), .A2(n24062), .ZN(n3764) );
  NAND2_X1 U9947 ( .A1(n11026), .A2(n3769), .ZN(n3768) );
  NOR2_X1 U9948 ( .A1(n11520), .A2(n10922), .ZN(n3769) );
  NAND2_X1 U9949 ( .A1(n3773), .A2(n19276), .ZN(n3772) );
  AND2_X1 U9950 ( .A1(n19278), .A2(n19126), .ZN(n19276) );
  NAND2_X1 U9952 ( .A1(n16371), .A2(n16616), .ZN(n3774) );
  AOI21_X1 U9953 ( .B1(n24556), .B2(n14510), .A(n14439), .ZN(n3776) );
  NAND2_X1 U9954 ( .A1(n24062), .A2(n3779), .ZN(n15647) );
  MUX2_X1 U9955 ( .A(n16404), .B(n16202), .S(n3544), .Z(n15813) );
  NAND2_X1 U9956 ( .A1(n1130), .A2(n7230), .ZN(n6982) );
  NOR2_X1 U9957 ( .A1(n3780), .A2(n7327), .ZN(n7329) );
  INV_X1 U9958 ( .A(n7232), .ZN(n3780) );
  MUX2_X1 U9959 ( .A(n24543), .B(n3783), .S(n17312), .Z(n17318) );
  NAND2_X1 U9960 ( .A1(n16716), .A2(n3783), .ZN(n16717) );
  NAND2_X1 U9961 ( .A1(n3785), .A2(n17410), .ZN(n3784) );
  NAND2_X1 U9962 ( .A1(n3822), .A2(n17409), .ZN(n3785) );
  NOR2_X1 U9963 ( .A1(n14165), .A2(n14167), .ZN(n13466) );
  NAND2_X1 U9964 ( .A1(n14268), .A2(n13840), .ZN(n3789) );
  NAND2_X1 U9966 ( .A1(n12739), .A2(n14436), .ZN(n3792) );
  AND2_X1 U9967 ( .A1(n20617), .A2(n20615), .ZN(n3795) );
  OR2_X1 U9968 ( .A1(n20614), .A2(n20571), .ZN(n3796) );
  XNOR2_X1 U9969 ( .A(n3797), .B(n8722), .ZN(n8723) );
  INV_X1 U9970 ( .A(n729), .ZN(n3798) );
  OAI21_X1 U9971 ( .B1(n9978), .B2(n9986), .A(n9665), .ZN(n3800) );
  NAND2_X1 U9972 ( .A1(n3799), .A2(n9664), .ZN(n9986) );
  INV_X1 U9973 ( .A(n9429), .ZN(n3799) );
  INV_X1 U9974 ( .A(n9429), .ZN(n9740) );
  NAND2_X1 U9977 ( .A1(n21290), .A2(n21848), .ZN(n3804) );
  NAND2_X1 U9978 ( .A1(n21289), .A2(n25395), .ZN(n3805) );
  NAND2_X2 U9980 ( .A1(n11595), .A2(n11590), .ZN(n13394) );
  NAND2_X1 U9981 ( .A1(n20193), .A2(n20432), .ZN(n5205) );
  NAND2_X1 U9983 ( .A1(n19214), .A2(n19215), .ZN(n3809) );
  NAND3_X1 U9985 ( .A1(n404), .A2(n12695), .A3(n12834), .ZN(n12696) );
  NAND3_X1 U9986 ( .A1(n12964), .A2(n12963), .A3(n404), .ZN(n12969) );
  NAND2_X1 U9987 ( .A1(n7960), .A2(n437), .ZN(n7964) );
  INV_X1 U9988 ( .A(n3818), .ZN(n16976) );
  XNOR2_X1 U9990 ( .A(n3819), .B(n21738), .ZN(n20741) );
  XNOR2_X1 U9991 ( .A(n3819), .B(n451), .ZN(n20811) );
  XNOR2_X1 U9992 ( .A(n3819), .B(n2215), .ZN(n21431) );
  XNOR2_X1 U9993 ( .A(n3819), .B(n21273), .ZN(n20984) );
  XNOR2_X1 U9994 ( .A(n3819), .B(n21633), .ZN(n20679) );
  NAND3_X1 U9995 ( .A1(n19171), .A2(n19169), .A3(n19170), .ZN(n3821) );
  XNOR2_X1 U9996 ( .A(n3823), .B(n20021), .ZN(n20033) );
  XNOR2_X1 U9997 ( .A(n3823), .B(n21160), .ZN(n20551) );
  XNOR2_X1 U9998 ( .A(n3823), .B(n23663), .ZN(n21344) );
  XNOR2_X1 U9999 ( .A(n3823), .B(n22525), .ZN(n21424) );
  NAND2_X1 U10001 ( .A1(n3828), .A2(n12854), .ZN(n3826) );
  INV_X1 U10002 ( .A(n12854), .ZN(n3827) );
  INV_X1 U10003 ( .A(n12853), .ZN(n3828) );
  NAND2_X1 U10006 ( .A1(n3832), .A2(n20131), .ZN(n3831) );
  MUX2_X1 U10007 ( .A(n21008), .B(n20522), .S(n20289), .Z(n3832) );
  NOR2_X1 U10009 ( .A1(n1449), .A2(n3835), .ZN(n3834) );
  OAI21_X1 U10010 ( .B1(n20126), .B2(n20125), .A(n20130), .ZN(n3835) );
  NAND3_X1 U10011 ( .A1(n3837), .A2(n22727), .A3(n3836), .ZN(n22730) );
  AND2_X1 U10013 ( .A1(n6967), .A2(n6576), .ZN(n3839) );
  OAI21_X1 U10014 ( .B1(n23969), .B2(n3841), .A(n3842), .ZN(n3840) );
  NAND2_X1 U10015 ( .A1(n23967), .A2(n23966), .ZN(n3841) );
  NAND2_X1 U10016 ( .A1(n22827), .A2(n23969), .ZN(n3842) );
  XNOR2_X1 U10017 ( .A(n3843), .B(n2126), .ZN(Ciphertext[184]) );
  NAND2_X1 U10018 ( .A1(n16023), .A2(n4957), .ZN(n16025) );
  OAI21_X1 U10019 ( .B1(n18969), .B2(n18970), .A(n3844), .ZN(n18982) );
  OAI22_X1 U10020 ( .A1(n19300), .A2(n19297), .B1(n18927), .B2(n19295), .ZN(
        n18968) );
  INV_X1 U10021 ( .A(n1363), .ZN(n3845) );
  NAND2_X1 U10022 ( .A1(n13513), .A2(n14153), .ZN(n13514) );
  NAND2_X1 U10024 ( .A1(n13304), .A2(n12914), .ZN(n3848) );
  INV_X1 U10026 ( .A(n14122), .ZN(n3851) );
  XNOR2_X1 U10028 ( .A(n18704), .B(n18701), .ZN(n3852) );
  XNOR2_X1 U10029 ( .A(n18703), .B(n18702), .ZN(n3853) );
  NAND2_X1 U10030 ( .A1(n3855), .A2(n17248), .ZN(n3854) );
  INV_X1 U10031 ( .A(n17272), .ZN(n3855) );
  OAI22_X1 U10032 ( .A1(n335), .A2(n3856), .B1(n21826), .B2(n22252), .ZN(n3890) );
  NOR2_X1 U10033 ( .A1(n23744), .A2(n1462), .ZN(n23731) );
  NAND2_X1 U10034 ( .A1(n23735), .A2(n3857), .ZN(n23737) );
  INV_X1 U10035 ( .A(n23744), .ZN(n3857) );
  NAND3_X1 U10036 ( .A1(n13311), .A2(n24487), .A3(n3859), .ZN(n3858) );
  NOR2_X1 U10037 ( .A1(n3866), .A2(n10111), .ZN(n3863) );
  NAND2_X1 U10038 ( .A1(n3865), .A2(n8644), .ZN(n3864) );
  AOI21_X1 U10039 ( .B1(n10107), .B2(n10106), .A(n8644), .ZN(n3866) );
  NAND3_X1 U10041 ( .A1(n3868), .A2(n11214), .A3(n233), .ZN(n3867) );
  NAND3_X1 U10042 ( .A1(n24340), .A2(n10810), .A3(n11212), .ZN(n3869) );
  NAND3_X1 U10043 ( .A1(n25082), .A2(n245), .A3(n22356), .ZN(n4203) );
  INV_X1 U10044 ( .A(n17341), .ZN(n17347) );
  NAND3_X1 U10045 ( .A1(n24307), .A2(n24895), .A3(n22043), .ZN(n3878) );
  OAI21_X1 U10046 ( .B1(n3876), .B2(n12673), .A(n13661), .ZN(n3873) );
  NAND2_X1 U10048 ( .A1(n13111), .A2(n4923), .ZN(n3874) );
  NAND2_X1 U10049 ( .A1(n3876), .A2(n13107), .ZN(n3875) );
  INV_X1 U10050 ( .A(n13110), .ZN(n3876) );
  XNOR2_X1 U10051 ( .A(n3877), .B(n22049), .ZN(Ciphertext[150]) );
  NAND3_X1 U10052 ( .A1(n3879), .A2(n22048), .A3(n3878), .ZN(n3877) );
  OAI21_X1 U10053 ( .B1(n22047), .B2(n24307), .A(n3880), .ZN(n3879) );
  NAND2_X1 U10054 ( .A1(n24307), .A2(n24983), .ZN(n3880) );
  XNOR2_X1 U10055 ( .A(n11798), .B(n3881), .ZN(n12126) );
  INV_X1 U10058 ( .A(n14200), .ZN(n3887) );
  NAND2_X1 U10060 ( .A1(n3886), .A2(n3888), .ZN(n3885) );
  NOR2_X1 U10061 ( .A1(n14945), .A2(n3887), .ZN(n3886) );
  INV_X1 U10062 ( .A(n14200), .ZN(n3889) );
  NAND2_X1 U10064 ( .A1(n3893), .A2(n3892), .ZN(n3891) );
  INV_X1 U10065 ( .A(n3894), .ZN(n5832) );
  NAND2_X1 U10066 ( .A1(n3894), .A2(n6791), .ZN(n6798) );
  NAND2_X1 U10067 ( .A1(n24362), .A2(n332), .ZN(n3895) );
  NAND2_X1 U10068 ( .A1(n21840), .A2(n22257), .ZN(n3896) );
  NAND2_X1 U10071 ( .A1(n7881), .A2(n7884), .ZN(n3898) );
  NAND2_X1 U10073 ( .A1(n3904), .A2(n341), .ZN(n3903) );
  MUX2_X1 U10074 ( .A(n18994), .B(n20319), .S(n19889), .Z(n3904) );
  INV_X1 U10076 ( .A(n22465), .ZN(n21929) );
  XNOR2_X2 U10077 ( .A(n20814), .B(n20813), .ZN(n22465) );
  NAND2_X1 U10078 ( .A1(n3907), .A2(n3906), .ZN(n21377) );
  NAND2_X1 U10080 ( .A1(n22463), .A2(n1363), .ZN(n22329) );
  NAND2_X1 U10083 ( .A1(n23042), .A2(n23048), .ZN(n3910) );
  INV_X1 U10084 ( .A(n23048), .ZN(n23059) );
  NOR2_X1 U10087 ( .A1(n20602), .A2(n3916), .ZN(n19848) );
  AND2_X1 U10088 ( .A1(n25476), .A2(n20597), .ZN(n3916) );
  INV_X1 U10089 ( .A(n19615), .ZN(n3919) );
  INV_X1 U10090 ( .A(n7380), .ZN(n7386) );
  NAND2_X1 U10091 ( .A1(n5656), .A2(n3923), .ZN(n3920) );
  XNOR2_X1 U10092 ( .A(n18605), .B(n896), .ZN(n17504) );
  AND2_X2 U10093 ( .A1(n3928), .A2(n3927), .ZN(n18605) );
  NAND2_X1 U10094 ( .A1(n16519), .A2(n17139), .ZN(n3927) );
  XNOR2_X1 U10095 ( .A(n15482), .B(n15481), .ZN(n3931) );
  NAND2_X1 U10096 ( .A1(n3933), .A2(n20591), .ZN(n3932) );
  NOR2_X1 U10099 ( .A1(n22465), .A2(n3938), .ZN(n3937) );
  INV_X1 U10100 ( .A(n22464), .ZN(n22461) );
  NAND3_X1 U10101 ( .A1(n22459), .A2(n3845), .A3(n22464), .ZN(n3939) );
  XNOR2_X1 U10102 ( .A(n15431), .B(n14805), .ZN(n15268) );
  XNOR2_X1 U10103 ( .A(n3941), .B(n3940), .ZN(n3942) );
  XNOR2_X1 U10104 ( .A(n15410), .B(n15431), .ZN(n3941) );
  XNOR2_X2 U10105 ( .A(n3942), .B(n13393), .ZN(n15667) );
  OAI21_X1 U10106 ( .B1(n12853), .B2(n3945), .A(n3944), .ZN(n13663) );
  NAND2_X1 U10107 ( .A1(n12673), .A2(n12856), .ZN(n3944) );
  OR2_X1 U10108 ( .A1(n12672), .A2(n12856), .ZN(n3945) );
  NAND2_X1 U10109 ( .A1(n25455), .A2(n15667), .ZN(n15670) );
  OAI21_X1 U10111 ( .B1(n267), .B2(n3947), .A(n3946), .ZN(n15669) );
  NAND2_X1 U10112 ( .A1(n267), .A2(n25455), .ZN(n3946) );
  INV_X1 U10113 ( .A(n15667), .ZN(n3947) );
  INV_X1 U10114 ( .A(n17039), .ZN(n3950) );
  NAND2_X1 U10115 ( .A1(n3955), .A2(n25215), .ZN(n3948) );
  NAND2_X1 U10116 ( .A1(n3950), .A2(n25058), .ZN(n3949) );
  NAND2_X1 U10117 ( .A1(n17037), .A2(n3951), .ZN(n3956) );
  NAND2_X1 U10118 ( .A1(n3953), .A2(n3952), .ZN(n18023) );
  NAND2_X1 U10119 ( .A1(n3956), .A2(n370), .ZN(n3952) );
  XNOR2_X2 U10120 ( .A(n10988), .B(n10987), .ZN(n3958) );
  NAND2_X1 U10121 ( .A1(n3958), .A2(n13102), .ZN(n12511) );
  NAND2_X1 U10122 ( .A1(n12742), .A2(n3958), .ZN(n13104) );
  NAND2_X1 U10123 ( .A1(n12744), .A2(n3958), .ZN(n12741) );
  MUX2_X1 U10124 ( .A(n13187), .B(n3958), .S(n13102), .Z(n11020) );
  OR2_X1 U10125 ( .A1(n13191), .A2(n3958), .ZN(n3957) );
  OAI22_X1 U10126 ( .A1(n2321), .A2(n13609), .B1(n14090), .B2(n3959), .ZN(
        n13542) );
  OAI21_X2 U10127 ( .B1(n22143), .B2(n22142), .A(n3960), .ZN(n23275) );
  NAND2_X1 U10128 ( .A1(n3961), .A2(n22274), .ZN(n3960) );
  INV_X1 U10129 ( .A(n19784), .ZN(n21068) );
  OAI21_X1 U10130 ( .B1(n24588), .B2(n3966), .A(n3965), .ZN(n3964) );
  NAND2_X1 U10131 ( .A1(n24588), .A2(n13888), .ZN(n3965) );
  NAND3_X1 U10132 ( .A1(n9919), .A2(n9914), .A3(n9920), .ZN(n9274) );
  NAND2_X1 U10134 ( .A1(n13062), .A2(n12439), .ZN(n3970) );
  MUX2_X1 U10135 ( .A(n12454), .B(n1353), .S(n13061), .Z(n3971) );
  NAND2_X1 U10136 ( .A1(n3973), .A2(n12459), .ZN(n3972) );
  NAND2_X1 U10137 ( .A1(n12460), .A2(n12652), .ZN(n3973) );
  NAND2_X1 U10138 ( .A1(n16741), .A2(n16742), .ZN(n3976) );
  NAND2_X1 U10139 ( .A1(n17090), .A2(n16740), .ZN(n3977) );
  INV_X1 U10140 ( .A(n16649), .ZN(n17085) );
  NAND2_X1 U10142 ( .A1(n4947), .A2(n4949), .ZN(n3978) );
  NAND3_X1 U10143 ( .A1(n3978), .A2(n22920), .A3(n23018), .ZN(n5465) );
  NAND2_X1 U10144 ( .A1(n3979), .A2(n24878), .ZN(n7268) );
  MUX2_X1 U10145 ( .A(n3979), .B(n24878), .S(n8370), .Z(n7840) );
  NAND2_X1 U10148 ( .A1(n3982), .A2(n5072), .ZN(n3981) );
  INV_X1 U10149 ( .A(n19245), .ZN(n3986) );
  XNOR2_X1 U10151 ( .A(n3990), .B(n18435), .ZN(n18620) );
  NAND2_X1 U10152 ( .A1(n10954), .A2(n10548), .ZN(n10958) );
  OAI21_X1 U10153 ( .B1(n3996), .B2(n3995), .A(n3994), .ZN(n19730) );
  NAND2_X1 U10154 ( .A1(n363), .A2(n18340), .ZN(n3994) );
  NAND2_X1 U10155 ( .A1(n3997), .A2(n24446), .ZN(n9086) );
  INV_X1 U10156 ( .A(n4096), .ZN(n3997) );
  OAI21_X1 U10157 ( .B1(n4096), .B2(n10058), .A(n3998), .ZN(n9691) );
  NOR3_X1 U10158 ( .A1(n24921), .A2(n23752), .A3(n4000), .ZN(n22524) );
  INV_X1 U10159 ( .A(n7481), .ZN(n7575) );
  MUX2_X1 U10160 ( .A(n7577), .B(n7573), .S(n7481), .Z(n4002) );
  NAND3_X1 U10162 ( .A1(n17012), .A2(n17356), .A3(n4004), .ZN(n4003) );
  NAND4_X2 U10163 ( .A1(n4007), .A2(n19378), .A3(n4006), .A4(n4008), .ZN(
        n20459) );
  NAND3_X1 U10164 ( .A1(n19377), .A2(n25067), .A3(n18876), .ZN(n4006) );
  NAND2_X1 U10165 ( .A1(n4010), .A2(n20022), .ZN(n4009) );
  NAND2_X1 U10166 ( .A1(n19727), .A2(n19728), .ZN(n4010) );
  NAND2_X1 U10167 ( .A1(n4012), .A2(n4011), .ZN(n10837) );
  NAND2_X1 U10168 ( .A1(n10829), .A2(n4013), .ZN(n4011) );
  NAND2_X1 U10169 ( .A1(n10830), .A2(n10518), .ZN(n4012) );
  NAND3_X1 U10170 ( .A1(n10829), .A2(n10275), .A3(n4013), .ZN(n10193) );
  NAND3_X1 U10171 ( .A1(n13728), .A2(n24588), .A3(n13945), .ZN(n4014) );
  NAND2_X1 U10172 ( .A1(n13909), .A2(n13951), .ZN(n4016) );
  NAND2_X1 U10175 ( .A1(n14218), .A2(n4019), .ZN(n13400) );
  MUX2_X1 U10176 ( .A(n14218), .B(n4019), .S(n14219), .Z(n14121) );
  NAND2_X1 U10177 ( .A1(n4020), .A2(n21046), .ZN(n4022) );
  NAND2_X1 U10178 ( .A1(n4022), .A2(n4021), .ZN(n4025) );
  NAND3_X1 U10179 ( .A1(n5162), .A2(n7237), .A3(n4023), .ZN(n4021) );
  NAND3_X1 U10180 ( .A1(n16175), .A2(n4027), .A3(n4026), .ZN(n16180) );
  NAND2_X1 U10181 ( .A1(n15655), .A2(n15656), .ZN(n4027) );
  OR2_X1 U10182 ( .A1(n15993), .A2(n4027), .ZN(n4645) );
  OR2_X1 U10183 ( .A1(n22529), .A2(n4034), .ZN(n4031) );
  OAI211_X1 U10184 ( .C1(n4031), .C2(n4030), .A(n4029), .B(n4028), .ZN(
        Ciphertext[93]) );
  NAND2_X1 U10185 ( .A1(n22529), .A2(n4034), .ZN(n4028) );
  INV_X1 U10186 ( .A(n4032), .ZN(n4030) );
  NAND3_X1 U10187 ( .A1(n4033), .A2(n3242), .A3(n23437), .ZN(n4032) );
  NAND2_X1 U10188 ( .A1(n285), .A2(n25003), .ZN(n4037) );
  INV_X1 U10189 ( .A(n17840), .ZN(n17726) );
  NAND2_X1 U10190 ( .A1(n4038), .A2(n285), .ZN(n4035) );
  NAND3_X1 U10191 ( .A1(n4037), .A2(n16661), .A3(n17399), .ZN(n4036) );
  NAND2_X1 U10192 ( .A1(n20437), .A2(n20194), .ZN(n5209) );
  INV_X1 U10193 ( .A(n10445), .ZN(n10905) );
  NAND2_X1 U10194 ( .A1(n13266), .A2(n24443), .ZN(n13268) );
  OAI21_X1 U10195 ( .B1(n12932), .B2(n25015), .A(n24443), .ZN(n12933) );
  AOI22_X1 U10198 ( .A1(n6480), .A2(n4042), .B1(n6479), .B2(n6924), .ZN(n6482)
         );
  NAND2_X1 U10199 ( .A1(n4043), .A2(n14130), .ZN(n13410) );
  INV_X1 U10200 ( .A(n15656), .ZN(n4045) );
  NAND2_X1 U10201 ( .A1(n15839), .A2(n15655), .ZN(n4044) );
  OAI21_X1 U10202 ( .B1(n10630), .B2(n11201), .A(n4047), .ZN(n4050) );
  NAND2_X1 U10204 ( .A1(n4050), .A2(n11195), .ZN(n4048) );
  XNOR2_X1 U10205 ( .A(n8520), .B(n4138), .ZN(n9500) );
  NAND2_X1 U10206 ( .A1(n10003), .A2(n9668), .ZN(n9670) );
  OR2_X1 U10207 ( .A1(n9500), .A2(n1796), .ZN(n10003) );
  OAI22_X1 U10208 ( .A1(n19252), .A2(n4052), .B1(n5134), .B2(n19250), .ZN(
        n4549) );
  INV_X1 U10209 ( .A(n19587), .ZN(n4052) );
  NAND2_X1 U10210 ( .A1(n25480), .A2(n6198), .ZN(n4053) );
  NAND3_X1 U10212 ( .A1(n25446), .A2(n15694), .A3(n16063), .ZN(n4054) );
  INV_X1 U10213 ( .A(n12482), .ZN(n4061) );
  NAND2_X1 U10214 ( .A1(n4055), .A2(n4057), .ZN(n13636) );
  NAND2_X1 U10215 ( .A1(n4058), .A2(n4056), .ZN(n4055) );
  NAND2_X1 U10216 ( .A1(n12482), .A2(n24573), .ZN(n4056) );
  NAND2_X1 U10217 ( .A1(n12483), .A2(n12710), .ZN(n4060) );
  NAND2_X1 U10218 ( .A1(n11024), .A2(n11518), .ZN(n11522) );
  NAND2_X1 U10219 ( .A1(n24902), .A2(n22166), .ZN(n4062) );
  NOR2_X1 U10221 ( .A1(n4064), .A2(n22166), .ZN(n4063) );
  NAND3_X1 U10222 ( .A1(n22117), .A2(n22170), .A3(n4064), .ZN(n22118) );
  INV_X1 U10223 ( .A(n20480), .ZN(n4065) );
  NOR2_X1 U10226 ( .A1(n20296), .A2(n4066), .ZN(n19047) );
  OAI21_X1 U10227 ( .B1(n20298), .B2(n4066), .A(n20140), .ZN(n19035) );
  AOI21_X1 U10228 ( .B1(n20296), .B2(n4066), .A(n20142), .ZN(n20143) );
  NAND3_X1 U10229 ( .A1(n10048), .A2(n10046), .A3(n4069), .ZN(n4068) );
  INV_X1 U10230 ( .A(n8977), .ZN(n4070) );
  NAND2_X1 U10231 ( .A1(n22298), .A2(n4072), .ZN(n4071) );
  NAND2_X1 U10232 ( .A1(n24914), .A2(n23251), .ZN(n22298) );
  NAND2_X1 U10234 ( .A1(n4075), .A2(n19296), .ZN(n4077) );
  INV_X1 U10236 ( .A(n19295), .ZN(n4075) );
  NAND2_X1 U10237 ( .A1(n4077), .A2(n18970), .ZN(n4076) );
  NAND2_X1 U10238 ( .A1(n6924), .A2(n4078), .ZN(n6779) );
  NAND3_X1 U10240 ( .A1(n24953), .A2(n4081), .A3(n4080), .ZN(n4079) );
  NAND2_X1 U10241 ( .A1(n17465), .A2(n25572), .ZN(n4082) );
  NOR2_X1 U10242 ( .A1(n16021), .A2(n287), .ZN(n4083) );
  XNOR2_X1 U10243 ( .A(n18197), .B(n17959), .ZN(n18692) );
  AND2_X2 U10244 ( .A1(n4084), .A2(n1492), .ZN(n18197) );
  OAI21_X1 U10245 ( .B1(n16988), .B2(n4085), .A(n5763), .ZN(n4084) );
  INV_X1 U10246 ( .A(n17363), .ZN(n4085) );
  XNOR2_X1 U10248 ( .A(n18044), .B(n4087), .ZN(n4086) );
  XNOR2_X1 U10249 ( .A(n18285), .B(n18562), .ZN(n4087) );
  INV_X1 U10250 ( .A(n11003), .ZN(n4088) );
  NAND2_X1 U10251 ( .A1(n10681), .A2(n10682), .ZN(n11003) );
  NAND2_X1 U10254 ( .A1(n10558), .A2(n10660), .ZN(n10397) );
  NAND2_X1 U10255 ( .A1(n13235), .A2(n12902), .ZN(n4490) );
  NAND3_X1 U10256 ( .A1(n24403), .A2(n15572), .A3(n4092), .ZN(n4090) );
  INV_X1 U10257 ( .A(n7657), .ZN(n4093) );
  INV_X1 U10258 ( .A(n12490), .ZN(n4094) );
  XNOR2_X1 U10259 ( .A(n4095), .B(n15016), .ZN(n14387) );
  NAND2_X1 U10260 ( .A1(n12649), .A2(n4405), .ZN(n12179) );
  OAI21_X1 U10261 ( .B1(n5323), .B2(n4405), .A(n13094), .ZN(n12870) );
  AND2_X1 U10262 ( .A1(n10053), .A2(n4096), .ZN(n10051) );
  NAND2_X1 U10263 ( .A1(n2902), .A2(n9866), .ZN(n9247) );
  XNOR2_X1 U10265 ( .A(n20677), .B(n20679), .ZN(n4101) );
  NAND2_X1 U10266 ( .A1(n20684), .A2(n4109), .ZN(n4102) );
  INV_X1 U10268 ( .A(n22389), .ZN(n4098) );
  NAND2_X1 U10269 ( .A1(n4372), .A2(n22387), .ZN(n4099) );
  OAI211_X2 U10271 ( .C1(n19426), .C2(n19177), .A(n18598), .B(n4103), .ZN(
        n20615) );
  NAND2_X1 U10272 ( .A1(n4104), .A2(n19427), .ZN(n4103) );
  OAI21_X1 U10273 ( .B1(n19177), .B2(n18597), .A(n1361), .ZN(n4104) );
  NAND2_X1 U10274 ( .A1(n5495), .A2(n5493), .ZN(n16549) );
  NAND2_X1 U10275 ( .A1(n6924), .A2(n6775), .ZN(n4106) );
  INV_X1 U10276 ( .A(n6292), .ZN(n6924) );
  XNOR2_X1 U10277 ( .A(n24027), .B(n8761), .ZN(n11447) );
  XNOR2_X1 U10278 ( .A(n24027), .B(n4107), .ZN(n11321) );
  NAND2_X1 U10279 ( .A1(n13935), .A2(n14245), .ZN(n13932) );
  AND2_X1 U10281 ( .A1(n23320), .A2(n4108), .ZN(n22628) );
  NAND2_X1 U10282 ( .A1(n19948), .A2(n20460), .ZN(n4110) );
  INV_X1 U10283 ( .A(n20394), .ZN(n19948) );
  NAND4_X1 U10284 ( .A1(n4113), .A2(n23193), .A3(n23202), .A4(n2903), .ZN(
        n4112) );
  NAND2_X1 U10285 ( .A1(n19376), .A2(n25010), .ZN(n17803) );
  NAND2_X1 U10287 ( .A1(n25128), .A2(n14241), .ZN(n4118) );
  NAND2_X1 U10290 ( .A1(n10159), .A2(n10162), .ZN(n4120) );
  NOR2_X1 U10291 ( .A1(n7734), .A2(n7642), .ZN(n5594) );
  NAND2_X1 U10293 ( .A1(n6600), .A2(n6824), .ZN(n4121) );
  OR2_X1 U10294 ( .A1(n2793), .A2(n13030), .ZN(n4124) );
  OR2_X2 U10295 ( .A1(n5786), .A2(n5785), .ZN(n7580) );
  NOR2_X1 U10297 ( .A1(n23359), .A2(n22961), .ZN(n23355) );
  NAND2_X1 U10299 ( .A1(n22956), .A2(n4128), .ZN(n4126) );
  NAND2_X1 U10300 ( .A1(n22955), .A2(n22954), .ZN(n4127) );
  INV_X1 U10301 ( .A(n22954), .ZN(n4128) );
  NAND2_X1 U10302 ( .A1(n4844), .A2(n4130), .ZN(n4129) );
  NAND2_X1 U10303 ( .A1(n14130), .A2(n13895), .ZN(n4130) );
  NAND2_X1 U10304 ( .A1(n13826), .A2(n4132), .ZN(n4131) );
  NAND2_X1 U10305 ( .A1(n4133), .A2(n1331), .ZN(n4132) );
  INV_X1 U10306 ( .A(n14127), .ZN(n4133) );
  NAND2_X1 U10307 ( .A1(n12885), .A2(n13223), .ZN(n12918) );
  XNOR2_X1 U10308 ( .A(n12400), .B(n11757), .ZN(n4134) );
  XNOR2_X1 U10309 ( .A(n11740), .B(n11739), .ZN(n11755) );
  INV_X1 U10310 ( .A(n19210), .ZN(n4135) );
  NAND3_X1 U10311 ( .A1(n9797), .A2(n9796), .A3(n4137), .ZN(n9801) );
  NAND2_X1 U10312 ( .A1(n9795), .A2(n4137), .ZN(n10002) );
  NAND2_X1 U10313 ( .A1(n9314), .A2(n4137), .ZN(n9312) );
  NAND2_X1 U10314 ( .A1(n19607), .A2(n4139), .ZN(n18864) );
  NAND2_X1 U10315 ( .A1(n4143), .A2(n11099), .ZN(n4142) );
  XNOR2_X2 U10316 ( .A(n14813), .B(n14812), .ZN(n16232) );
  NAND2_X1 U10317 ( .A1(n7476), .A2(n7423), .ZN(n4145) );
  XNOR2_X1 U10318 ( .A(n4146), .B(n8084), .ZN(n8416) );
  INV_X1 U10319 ( .A(n8411), .ZN(n4146) );
  XNOR2_X1 U10320 ( .A(n4147), .B(n8084), .ZN(n8750) );
  INV_X1 U10321 ( .A(n8745), .ZN(n4147) );
  NAND2_X1 U10322 ( .A1(n4148), .A2(n6659), .ZN(n7155) );
  NAND3_X1 U10323 ( .A1(n4150), .A2(n4151), .A3(n4149), .ZN(n4148) );
  NAND2_X1 U10324 ( .A1(n6657), .A2(n6072), .ZN(n4151) );
  NOR2_X1 U10325 ( .A1(n11338), .A2(n25025), .ZN(n4152) );
  XNOR2_X1 U10328 ( .A(n16799), .B(n4153), .ZN(n17328) );
  XNOR2_X1 U10329 ( .A(n4154), .B(n16799), .ZN(n18076) );
  INV_X1 U10330 ( .A(n18096), .ZN(n4154) );
  XNOR2_X1 U10331 ( .A(n18700), .B(n4155), .ZN(n18702) );
  INV_X1 U10332 ( .A(n16799), .ZN(n4155) );
  OAI211_X1 U10335 ( .C1(n11214), .C2(n233), .A(n10810), .B(n11215), .ZN(n4156) );
  INV_X1 U10336 ( .A(n11216), .ZN(n10810) );
  XNOR2_X1 U10337 ( .A(n4157), .B(n21537), .ZN(n21539) );
  XNOR2_X1 U10338 ( .A(n21535), .B(n4158), .ZN(n4157) );
  NAND2_X1 U10339 ( .A1(n4161), .A2(n4160), .ZN(n4159) );
  INV_X1 U10340 ( .A(n19973), .ZN(n4160) );
  NOR2_X1 U10341 ( .A1(n19974), .A2(n4164), .ZN(n4161) );
  NAND2_X1 U10342 ( .A1(n19973), .A2(n4164), .ZN(n4162) );
  NAND2_X1 U10343 ( .A1(n19974), .A2(n4164), .ZN(n4163) );
  XNOR2_X1 U10344 ( .A(n18334), .B(n4761), .ZN(n18615) );
  NAND2_X1 U10345 ( .A1(n17089), .A2(n17088), .ZN(n4165) );
  NAND3_X1 U10346 ( .A1(n262), .A2(n9468), .A3(n9281), .ZN(n4166) );
  NAND2_X1 U10349 ( .A1(n19235), .A2(n19237), .ZN(n4167) );
  NAND2_X1 U10350 ( .A1(n19235), .A2(n19112), .ZN(n18869) );
  NAND2_X1 U10351 ( .A1(n1428), .A2(n4168), .ZN(n4282) );
  NAND2_X1 U10352 ( .A1(n23372), .A2(n24412), .ZN(n4171) );
  NAND2_X1 U10353 ( .A1(n4170), .A2(n4632), .ZN(n4633) );
  NAND2_X1 U10354 ( .A1(n4171), .A2(n24404), .ZN(n22993) );
  NAND2_X1 U10355 ( .A1(n22610), .A2(n22611), .ZN(n23048) );
  INV_X1 U10356 ( .A(n18761), .ZN(n4172) );
  NAND2_X1 U10357 ( .A1(n4172), .A2(n24329), .ZN(n17554) );
  XNOR2_X1 U10358 ( .A(n21729), .B(n1854), .ZN(n20733) );
  NAND4_X2 U10359 ( .A1(n4174), .A2(n19692), .A3(n19693), .A4(n4173), .ZN(
        n21729) );
  NAND3_X1 U10360 ( .A1(n20322), .A2(n24917), .A3(n19889), .ZN(n4173) );
  NAND2_X1 U10362 ( .A1(n1327), .A2(n24460), .ZN(n4175) );
  NAND3_X1 U10363 ( .A1(n19948), .A2(n20460), .A3(n20395), .ZN(n4176) );
  NAND2_X1 U10364 ( .A1(n4177), .A2(n6395), .ZN(n6399) );
  OAI21_X1 U10366 ( .B1(n13172), .B2(n13171), .A(n13170), .ZN(n4179) );
  XNOR2_X1 U10367 ( .A(n8988), .B(n9041), .ZN(n8621) );
  XNOR2_X1 U10368 ( .A(n4180), .B(n9041), .ZN(n8287) );
  INV_X1 U10369 ( .A(n8498), .ZN(n4180) );
  XNOR2_X1 U10370 ( .A(n12269), .B(n12270), .ZN(n4182) );
  NAND2_X1 U10371 ( .A1(n20413), .A2(n20264), .ZN(n4184) );
  INV_X1 U10372 ( .A(n4190), .ZN(n4193) );
  OR2_X1 U10373 ( .A1(n23867), .A2(n4189), .ZN(n4187) );
  NAND4_X1 U10374 ( .A1(n4191), .A2(n23867), .A3(n4190), .A4(n4189), .ZN(n4188) );
  INV_X1 U10375 ( .A(n4192), .ZN(n4191) );
  NAND2_X1 U10376 ( .A1(n20476), .A2(n20353), .ZN(n20354) );
  OR2_X1 U10377 ( .A1(n19420), .A2(n19418), .ZN(n4195) );
  NAND2_X1 U10378 ( .A1(n4196), .A2(n13110), .ZN(n12632) );
  NAND2_X1 U10379 ( .A1(n4196), .A2(n13108), .ZN(n4924) );
  NAND2_X1 U10380 ( .A1(n5211), .A2(n16404), .ZN(n4197) );
  MUX2_X1 U10381 ( .A(n16956), .B(n17414), .S(n17413), .Z(n14353) );
  NAND2_X1 U10382 ( .A1(n4198), .A2(n25572), .ZN(n16506) );
  INV_X1 U10383 ( .A(n13281), .ZN(n12698) );
  NAND2_X1 U10384 ( .A1(n4202), .A2(n4201), .ZN(n4200) );
  NAND3_X1 U10385 ( .A1(n14191), .A2(n14189), .A3(n14142), .ZN(n4201) );
  NOR2_X1 U10386 ( .A1(n8023), .A2(n8022), .ZN(n4206) );
  NAND3_X1 U10387 ( .A1(n4209), .A2(n9506), .A3(n4208), .ZN(n4207) );
  NAND2_X1 U10388 ( .A1(n10088), .A2(n9507), .ZN(n4209) );
  NAND2_X1 U10389 ( .A1(n24575), .A2(n9786), .ZN(n4210) );
  NAND2_X1 U10390 ( .A1(n10508), .A2(n10931), .ZN(n10425) );
  NAND4_X1 U10391 ( .A1(n4216), .A2(n4217), .A3(n4218), .A4(n21357), .ZN(n4215) );
  NAND2_X1 U10392 ( .A1(n21351), .A2(n21352), .ZN(n4217) );
  AND2_X1 U10393 ( .A1(n21350), .A2(n21349), .ZN(n4218) );
  NAND2_X1 U10394 ( .A1(n4221), .A2(n21844), .ZN(n4219) );
  OAI211_X2 U10396 ( .C1(n14060), .C2(n14415), .A(n4224), .B(n4222), .ZN(
        n15133) );
  NAND3_X1 U10398 ( .A1(n4225), .A2(n14849), .A3(n14415), .ZN(n4224) );
  OAI211_X2 U10399 ( .C1(n13263), .C2(n13484), .A(n4226), .B(n1407), .ZN(
        n15062) );
  XNOR2_X1 U10400 ( .A(n4227), .B(n20982), .ZN(n21430) );
  XNOR2_X1 U10401 ( .A(n4227), .B(n889), .ZN(n20847) );
  XNOR2_X1 U10402 ( .A(n4227), .B(n21630), .ZN(n21631) );
  XNOR2_X1 U10403 ( .A(n4227), .B(n4294), .ZN(n20700) );
  NAND2_X1 U10406 ( .A1(n4234), .A2(n4236), .ZN(n4231) );
  NOR2_X1 U10407 ( .A1(n20520), .A2(n20515), .ZN(n19797) );
  NAND4_X2 U10408 ( .A1(n4239), .A2(n19111), .A3(n4238), .A4(n4977), .ZN(
        n20272) );
  NAND2_X1 U10409 ( .A1(n19110), .A2(n24908), .ZN(n4238) );
  NAND2_X1 U10410 ( .A1(n19108), .A2(n19384), .ZN(n4239) );
  NAND2_X1 U10411 ( .A1(n12688), .A2(n13318), .ZN(n4240) );
  OAI21_X1 U10412 ( .B1(n12946), .B2(n13318), .A(n4240), .ZN(n12582) );
  NOR2_X1 U10413 ( .A1(n4241), .A2(n13318), .ZN(n12944) );
  NAND2_X1 U10414 ( .A1(n13317), .A2(n4241), .ZN(n12687) );
  XNOR2_X1 U10415 ( .A(n15504), .B(n15503), .ZN(n15511) );
  XNOR2_X1 U10416 ( .A(n4242), .B(n23257), .ZN(Ciphertext[47]) );
  OAI211_X1 U10417 ( .C1(n23256), .C2(n23255), .A(n4244), .B(n4243), .ZN(n4242) );
  NAND2_X1 U10418 ( .A1(n23256), .A2(n23254), .ZN(n4244) );
  NOR2_X2 U10419 ( .A1(n22287), .A2(n22286), .ZN(n23256) );
  OAI21_X1 U10421 ( .B1(n16269), .B2(n24366), .A(n4249), .ZN(n15162) );
  XNOR2_X1 U10422 ( .A(n4250), .B(n18289), .ZN(n18086) );
  XNOR2_X1 U10423 ( .A(n4250), .B(n18190), .ZN(n17788) );
  XNOR2_X1 U10424 ( .A(n4250), .B(n20609), .ZN(n18228) );
  XNOR2_X1 U10425 ( .A(n4250), .B(n3158), .ZN(n18638) );
  XNOR2_X1 U10426 ( .A(n4250), .B(n21711), .ZN(n18414) );
  XNOR2_X1 U10427 ( .A(n4250), .B(n17851), .ZN(n17852) );
  NAND2_X1 U10428 ( .A1(n11058), .A2(n11057), .ZN(n4251) );
  NAND2_X1 U10429 ( .A1(n9808), .A2(n9809), .ZN(n4252) );
  NAND2_X1 U10430 ( .A1(n9776), .A2(n4254), .ZN(n4253) );
  AOI21_X1 U10431 ( .B1(n9836), .B2(n428), .A(n4257), .ZN(n9840) );
  AND2_X1 U10432 ( .A1(n8359), .A2(n10094), .ZN(n4257) );
  NAND2_X1 U10434 ( .A1(n9515), .A2(n9837), .ZN(n4258) );
  OAI21_X1 U10435 ( .B1(n9514), .B2(n428), .A(n10097), .ZN(n9518) );
  INV_X1 U10436 ( .A(n7948), .ZN(n4259) );
  OAI211_X2 U10437 ( .C1(n19289), .C2(n25448), .A(n4261), .B(n4260), .ZN(
        n20419) );
  INV_X1 U10438 ( .A(n19559), .ZN(n4262) );
  XNOR2_X1 U10439 ( .A(n21227), .B(n4263), .ZN(n22004) );
  XNOR2_X1 U10440 ( .A(n21231), .B(n4263), .ZN(n21233) );
  XNOR2_X1 U10441 ( .A(n24485), .B(n4263), .ZN(n21270) );
  XNOR2_X1 U10442 ( .A(n4263), .B(n1935), .ZN(n21544) );
  NAND2_X1 U10443 ( .A1(n17054), .A2(n25031), .ZN(n4266) );
  NAND2_X1 U10444 ( .A1(n16609), .A2(n16722), .ZN(n4267) );
  NOR2_X1 U10445 ( .A1(n16001), .A2(n16266), .ZN(n4270) );
  NAND2_X1 U10446 ( .A1(n5447), .A2(n16266), .ZN(n16272) );
  NAND2_X1 U10447 ( .A1(n24385), .A2(n17059), .ZN(n16722) );
  NOR2_X1 U10450 ( .A1(n22657), .A2(n4273), .ZN(n22363) );
  NAND2_X1 U10452 ( .A1(n20442), .A2(n4273), .ZN(n20443) );
  AND2_X1 U10453 ( .A1(n22657), .A2(n4273), .ZN(n4272) );
  OAI21_X1 U10454 ( .B1(n1457), .B2(n22609), .A(n4273), .ZN(n4283) );
  NAND2_X1 U10456 ( .A1(n4276), .A2(n20669), .ZN(n20340) );
  OAI21_X1 U10457 ( .B1(n20338), .B2(n20666), .A(n20671), .ZN(n4276) );
  INV_X1 U10459 ( .A(n7989), .ZN(n7826) );
  NAND3_X1 U10460 ( .A1(n7827), .A2(n7982), .A3(n7826), .ZN(n4277) );
  NAND3_X1 U10461 ( .A1(n7828), .A2(n7989), .A3(n7825), .ZN(n4278) );
  OAI21_X2 U10465 ( .B1(n22815), .B2(n22816), .A(n22814), .ZN(n24011) );
  NAND3_X1 U10466 ( .A1(n4281), .A2(n24753), .A3(n11101), .ZN(n11103) );
  NAND2_X1 U10467 ( .A1(n4286), .A2(n17069), .ZN(n17070) );
  NAND2_X1 U10468 ( .A1(n17944), .A2(n4290), .ZN(n4289) );
  OR2_X1 U10469 ( .A1(n19327), .A2(n4291), .ZN(n4290) );
  OAI21_X1 U10470 ( .B1(n20666), .B2(n20670), .A(n4292), .ZN(n20351) );
  NAND2_X1 U10471 ( .A1(n20336), .A2(n20668), .ZN(n4292) );
  OAI21_X2 U10472 ( .B1(n17310), .B2(n18933), .A(n17309), .ZN(n20668) );
  AOI22_X2 U10473 ( .A1(n20351), .A2(n20341), .B1(n20670), .B2(n18745), .ZN(
        n21247) );
  XNOR2_X1 U10474 ( .A(n4294), .B(n22697), .ZN(n20047) );
  XNOR2_X1 U10475 ( .A(n4294), .B(n2036), .ZN(n20983) );
  XNOR2_X1 U10476 ( .A(n4294), .B(n21699), .ZN(n21221) );
  XNOR2_X1 U10477 ( .A(n21054), .B(n4294), .ZN(n21564) );
  NAND2_X1 U10479 ( .A1(n4295), .A2(n20302), .ZN(n4692) );
  INV_X1 U10480 ( .A(n20009), .ZN(n4295) );
  NAND2_X1 U10481 ( .A1(n4298), .A2(n24570), .ZN(n4297) );
  INV_X1 U10482 ( .A(n16774), .ZN(n4299) );
  AND2_X1 U10484 ( .A1(n4303), .A2(n17114), .ZN(n5429) );
  NOR2_X1 U10485 ( .A1(n17100), .A2(n17114), .ZN(n5760) );
  INV_X1 U10486 ( .A(n17118), .ZN(n4303) );
  OAI21_X1 U10487 ( .B1(n16573), .B2(n25357), .A(n4304), .ZN(n4714) );
  MUX2_X1 U10489 ( .A(n13965), .B(n11806), .S(n13966), .Z(n13885) );
  NAND2_X1 U10490 ( .A1(n13965), .A2(n11806), .ZN(n4305) );
  MUX2_X1 U10491 ( .A(n13725), .B(n13883), .S(n11806), .Z(n13726) );
  NOR2_X1 U10492 ( .A1(n20478), .A2(n20003), .ZN(n19627) );
  NOR2_X2 U10493 ( .A1(n18838), .A2(n4306), .ZN(n20478) );
  AOI21_X1 U10494 ( .B1(n19239), .B2(n19064), .A(n4307), .ZN(n4306) );
  NAND2_X1 U10496 ( .A1(n19213), .A2(n4315), .ZN(n4314) );
  XNOR2_X1 U10497 ( .A(n11615), .B(n11614), .ZN(n4316) );
  OAI21_X1 U10498 ( .B1(n19363), .B2(n24424), .A(n24968), .ZN(n4317) );
  NAND3_X1 U10499 ( .A1(n13065), .A2(n4319), .A3(n4318), .ZN(n13385) );
  NAND3_X1 U10500 ( .A1(n13064), .A2(n13063), .A3(n12737), .ZN(n4318) );
  INV_X1 U10501 ( .A(n13159), .ZN(n12737) );
  OAI21_X1 U10502 ( .B1(n13062), .B2(n4320), .A(n13163), .ZN(n4319) );
  INV_X1 U10503 ( .A(n6956), .ZN(n6702) );
  OAI21_X1 U10504 ( .B1(n3926), .B2(n6703), .A(n4323), .ZN(n4322) );
  INV_X1 U10505 ( .A(n11009), .ZN(n4326) );
  NOR2_X1 U10506 ( .A1(n1218), .A2(n11009), .ZN(n11055) );
  INV_X1 U10507 ( .A(n13796), .ZN(n13774) );
  XNOR2_X1 U10508 ( .A(n4334), .B(n8914), .ZN(n8131) );
  XNOR2_X1 U10509 ( .A(n8914), .B(n4335), .ZN(n8197) );
  NAND2_X1 U10510 ( .A1(n4336), .A2(n13072), .ZN(n12775) );
  NAND3_X1 U10511 ( .A1(n23179), .A2(n23167), .A3(n25488), .ZN(n22555) );
  NAND3_X1 U10512 ( .A1(n4344), .A2(n4347), .A3(n7130), .ZN(n8826) );
  NAND2_X1 U10513 ( .A1(n4345), .A2(n7320), .ZN(n4344) );
  NAND2_X1 U10514 ( .A1(n20650), .A2(n24415), .ZN(n4348) );
  NAND2_X1 U10516 ( .A1(n20648), .A2(n22141), .ZN(n4351) );
  OR2_X1 U10518 ( .A1(n15802), .A2(n1365), .ZN(n15594) );
  INV_X1 U10519 ( .A(n24826), .ZN(n4353) );
  NAND2_X1 U10520 ( .A1(n4355), .A2(n14160), .ZN(n4354) );
  XNOR2_X1 U10521 ( .A(n12048), .B(n1792), .ZN(n11916) );
  NAND2_X1 U10522 ( .A1(n10899), .A2(n4341), .ZN(n4358) );
  NAND2_X1 U10523 ( .A1(n23722), .A2(n23727), .ZN(n23726) );
  NAND2_X1 U10525 ( .A1(n22081), .A2(n4360), .ZN(n4359) );
  INV_X1 U10526 ( .A(n22079), .ZN(n4360) );
  NAND2_X1 U10527 ( .A1(n22080), .A2(n22079), .ZN(n4361) );
  NAND2_X1 U10528 ( .A1(n4364), .A2(n3726), .ZN(n4363) );
  MUX2_X1 U10529 ( .A(n19163), .B(n19393), .S(n19162), .Z(n4364) );
  NAND2_X1 U10531 ( .A1(n8316), .A2(n8315), .ZN(n4366) );
  NAND3_X1 U10534 ( .A1(n24532), .A2(n24586), .A3(n16107), .ZN(n15628) );
  NAND2_X1 U10535 ( .A1(n6942), .A2(n6941), .ZN(n4369) );
  NAND2_X1 U10536 ( .A1(n5560), .A2(n6947), .ZN(n4370) );
  NOR3_X1 U10537 ( .A1(n22974), .A2(n22975), .A3(n22387), .ZN(n4371) );
  NOR2_X1 U10538 ( .A1(n4373), .A2(n21822), .ZN(n19343) );
  NOR2_X1 U10539 ( .A1(n332), .A2(n21822), .ZN(n4374) );
  XNOR2_X1 U10540 ( .A(n8039), .B(n8452), .ZN(n9114) );
  XNOR2_X1 U10541 ( .A(n9114), .B(n9115), .ZN(n9119) );
  OAI21_X1 U10542 ( .B1(n7535), .B2(n7536), .A(n8013), .ZN(n4377) );
  XNOR2_X1 U10543 ( .A(n4378), .B(n2034), .ZN(n7204) );
  XNOR2_X1 U10544 ( .A(n4378), .B(n2193), .ZN(n8264) );
  XNOR2_X1 U10545 ( .A(n8485), .B(n4378), .ZN(n8246) );
  XNOR2_X1 U10546 ( .A(n8698), .B(n4378), .ZN(n7778) );
  NAND2_X1 U10547 ( .A1(n12107), .A2(n400), .ZN(n4379) );
  NAND2_X1 U10548 ( .A1(n4381), .A2(n13335), .ZN(n4380) );
  INV_X1 U10549 ( .A(n13337), .ZN(n4381) );
  NAND2_X1 U10550 ( .A1(n14005), .A2(n24462), .ZN(n4383) );
  XNOR2_X1 U10551 ( .A(n17648), .B(n4384), .ZN(n4385) );
  INV_X1 U10552 ( .A(n17918), .ZN(n4384) );
  XNOR2_X1 U10553 ( .A(n8697), .B(n8696), .ZN(n4386) );
  INV_X1 U10554 ( .A(n12834), .ZN(n13273) );
  NAND3_X1 U10555 ( .A1(n4394), .A2(n4393), .A3(n4390), .ZN(n11736) );
  NAND3_X1 U10556 ( .A1(n4326), .A2(n11057), .A3(n10694), .ZN(n4393) );
  NOR2_X2 U10557 ( .A1(n9794), .A2(n9793), .ZN(n11052) );
  NAND2_X1 U10558 ( .A1(n11055), .A2(n11054), .ZN(n4394) );
  XNOR2_X1 U10559 ( .A(n21092), .B(n24453), .ZN(n21095) );
  XNOR2_X1 U10560 ( .A(n21542), .B(n24453), .ZN(n21546) );
  XNOR2_X1 U10561 ( .A(n21611), .B(n4396), .ZN(n20035) );
  NOR2_X1 U10564 ( .A1(n4525), .A2(n13901), .ZN(n14309) );
  OAI21_X1 U10565 ( .B1(n7972), .B2(n7977), .A(n4400), .ZN(n7817) );
  MUX2_X1 U10566 ( .A(n7972), .B(n7973), .S(n4400), .Z(n7979) );
  AOI21_X1 U10567 ( .B1(n7049), .B2(n7819), .A(n4400), .ZN(n7050) );
  XNOR2_X1 U10568 ( .A(n8881), .B(n4401), .ZN(n8883) );
  OAI21_X1 U10569 ( .B1(n20069), .B2(n20068), .A(n20067), .ZN(n20070) );
  NAND2_X1 U10570 ( .A1(n20068), .A2(n19849), .ZN(n20067) );
  NAND2_X1 U10571 ( .A1(n18849), .A2(n18848), .ZN(n4404) );
  NAND2_X1 U10575 ( .A1(n23397), .A2(n23396), .ZN(n4406) );
  NOR2_X1 U10579 ( .A1(n23396), .A2(n23394), .ZN(n4411) );
  AND2_X1 U10580 ( .A1(n17172), .A2(n17175), .ZN(n4414) );
  XNOR2_X1 U10583 ( .A(n15191), .B(n15112), .ZN(n14937) );
  XNOR2_X1 U10584 ( .A(n15246), .B(n14937), .ZN(n14583) );
  NAND2_X1 U10585 ( .A1(n4419), .A2(n4417), .ZN(n4416) );
  NAND2_X1 U10586 ( .A1(n16148), .A2(n4418), .ZN(n4417) );
  AOI21_X1 U10587 ( .B1(n16097), .B2(n16096), .A(n213), .ZN(n4419) );
  AND2_X1 U10588 ( .A1(n4422), .A2(n412), .ZN(n10439) );
  NAND2_X1 U10589 ( .A1(n10438), .A2(n4422), .ZN(n10442) );
  NAND2_X1 U10591 ( .A1(n14154), .A2(n14153), .ZN(n4424) );
  NAND2_X1 U10592 ( .A1(n4426), .A2(n17320), .ZN(n17324) );
  INV_X1 U10593 ( .A(n16607), .ZN(n4426) );
  NAND2_X2 U10594 ( .A1(n4428), .A2(n6378), .ZN(n7843) );
  NAND2_X1 U10595 ( .A1(n6790), .A2(n6089), .ZN(n4428) );
  OR2_X1 U10597 ( .A1(n19283), .A2(n19127), .ZN(n4429) );
  NAND3_X1 U10598 ( .A1(n4432), .A2(n19518), .A3(n4431), .ZN(n4430) );
  NAND2_X1 U10599 ( .A1(n4433), .A2(n19526), .ZN(n4432) );
  OAI211_X1 U10601 ( .C1(n21814), .C2(n22063), .A(n21813), .B(n21812), .ZN(
        n4434) );
  XNOR2_X2 U10603 ( .A(n16785), .B(n16786), .ZN(n4436) );
  AND2_X1 U10604 ( .A1(n19266), .A2(n4436), .ZN(n5239) );
  NAND2_X1 U10605 ( .A1(n1299), .A2(n4436), .ZN(n16822) );
  NAND2_X1 U10607 ( .A1(n18916), .A2(n4436), .ZN(n19149) );
  NAND3_X1 U10608 ( .A1(n1336), .A2(n22244), .A3(n4437), .ZN(n22246) );
  INV_X1 U10609 ( .A(n22059), .ZN(n4437) );
  AOI21_X1 U10610 ( .B1(n19601), .B2(n18037), .A(n4438), .ZN(n19603) );
  NAND2_X1 U10611 ( .A1(n19255), .A2(n19598), .ZN(n4439) );
  NAND3_X1 U10613 ( .A1(n16075), .A2(n1365), .A3(n16077), .ZN(n4440) );
  NOR2_X1 U10614 ( .A1(n22334), .A2(n22333), .ZN(n4441) );
  NAND2_X1 U10616 ( .A1(n4449), .A2(n13266), .ZN(n4443) );
  NAND2_X1 U10617 ( .A1(n14301), .A2(n13888), .ZN(n13944) );
  INV_X1 U10620 ( .A(n12835), .ZN(n4445) );
  NAND2_X1 U10621 ( .A1(n4930), .A2(n12680), .ZN(n4449) );
  NAND2_X1 U10622 ( .A1(n4450), .A2(n24391), .ZN(n5295) );
  NAND2_X1 U10624 ( .A1(n12819), .A2(n4451), .ZN(n4721) );
  NAND2_X1 U10625 ( .A1(n14168), .A2(n13742), .ZN(n4452) );
  OAI211_X2 U10627 ( .C1(n10185), .C2(n10186), .A(n10184), .B(n10183), .ZN(
        n10660) );
  INV_X1 U10628 ( .A(n20434), .ZN(n19225) );
  MUX2_X2 U10629 ( .A(n9583), .B(n9582), .S(n25463), .Z(n10617) );
  INV_X1 U10630 ( .A(n4882), .ZN(n18028) );
  MUX2_X2 U10633 ( .A(n10067), .B(n10066), .S(n10065), .Z(n11070) );
  OAI21_X1 U10635 ( .B1(n239), .B2(n9864), .A(n4453), .ZN(n8064) );
  NAND2_X1 U10636 ( .A1(n9864), .A2(n9857), .ZN(n4453) );
  INV_X1 U10637 ( .A(n9859), .ZN(n4454) );
  MUX2_X1 U10638 ( .A(n9860), .B(n9559), .S(n239), .Z(n9262) );
  XNOR2_X1 U10640 ( .A(n4456), .B(n21167), .ZN(n4455) );
  NAND2_X1 U10641 ( .A1(n19276), .A2(n1334), .ZN(n4458) );
  NAND2_X1 U10643 ( .A1(n19125), .A2(n5573), .ZN(n4459) );
  INV_X1 U10644 ( .A(n10713), .ZN(n4463) );
  OAI21_X1 U10645 ( .B1(n5744), .B2(n11131), .A(n11129), .ZN(n4465) );
  NOR2_X1 U10646 ( .A1(n4463), .A2(n10838), .ZN(n4462) );
  OAI21_X1 U10647 ( .B1(n22656), .B2(n331), .A(n4466), .ZN(n4473) );
  NAND2_X1 U10648 ( .A1(n22813), .A2(n22656), .ZN(n4466) );
  OAI21_X1 U10649 ( .B1(n22656), .B2(n22657), .A(n25241), .ZN(n4467) );
  INV_X1 U10650 ( .A(n22658), .ZN(n4470) );
  XNOR2_X2 U10651 ( .A(n20408), .B(n20407), .ZN(n22813) );
  NAND2_X1 U10652 ( .A1(n24015), .A2(n4478), .ZN(n4474) );
  NAND2_X1 U10653 ( .A1(n4478), .A2(n23993), .ZN(n23987) );
  NAND2_X1 U10654 ( .A1(n23982), .A2(n4478), .ZN(n23981) );
  AOI21_X1 U10655 ( .B1(n24954), .B2(n4477), .A(n23983), .ZN(n4476) );
  NAND4_X2 U10656 ( .A1(n12436), .A2(n12437), .A3(n12438), .A4(n12435), .ZN(
        n14167) );
  NOR2_X2 U10657 ( .A1(n19593), .A2(n4479), .ZN(n20377) );
  MUX2_X1 U10658 ( .A(n24483), .B(n19591), .S(n19077), .Z(n4480) );
  NOR2_X1 U10659 ( .A1(n10365), .A2(n4481), .ZN(n10321) );
  OAI21_X1 U10660 ( .B1(n10684), .B2(n11004), .A(n4481), .ZN(n11008) );
  NAND2_X1 U10661 ( .A1(n17012), .A2(n25491), .ZN(n4482) );
  OAI21_X1 U10662 ( .B1(n7956), .B2(n4483), .A(n7955), .ZN(n7957) );
  NAND2_X1 U10663 ( .A1(n4486), .A2(n4484), .ZN(n12887) );
  NAND3_X1 U10665 ( .A1(n17613), .A2(n17409), .A3(n17608), .ZN(n4488) );
  NAND3_X1 U10666 ( .A1(n19948), .A2(n4489), .A3(n20461), .ZN(n19949) );
  MUX2_X1 U10667 ( .A(n20383), .B(n20384), .S(n20459), .Z(n20398) );
  NAND2_X1 U10669 ( .A1(n12937), .A2(n4490), .ZN(n4492) );
  NAND2_X1 U10671 ( .A1(n11006), .A2(n24420), .ZN(n4495) );
  NAND2_X1 U10672 ( .A1(n11836), .A2(n12902), .ZN(n4497) );
  NAND2_X1 U10674 ( .A1(n17416), .A2(n16565), .ZN(n4502) );
  AOI21_X1 U10675 ( .B1(n4503), .B2(n6678), .A(n6281), .ZN(n6282) );
  XNOR2_X1 U10676 ( .A(n14843), .B(n14842), .ZN(n4504) );
  INV_X1 U10677 ( .A(n10753), .ZN(n4505) );
  NAND2_X1 U10678 ( .A1(n9364), .A2(n4506), .ZN(n10204) );
  INV_X1 U10679 ( .A(n17297), .ZN(n4508) );
  INV_X1 U10680 ( .A(n4510), .ZN(n14021) );
  NAND2_X1 U10681 ( .A1(n4510), .A2(n14022), .ZN(n12513) );
  NAND2_X1 U10682 ( .A1(n14086), .A2(n4510), .ZN(n14087) );
  NAND2_X1 U10683 ( .A1(n2008), .A2(n6933), .ZN(n4512) );
  NAND2_X1 U10684 ( .A1(n11113), .A2(n11116), .ZN(n5351) );
  NAND2_X1 U10685 ( .A1(n9789), .A2(n24575), .ZN(n5354) );
  NAND2_X1 U10686 ( .A1(n22151), .A2(n4513), .ZN(n22152) );
  OR2_X1 U10687 ( .A1(n23647), .A2(n23612), .ZN(n4514) );
  OR2_X1 U10688 ( .A1(n24366), .A2(n4516), .ZN(n4515) );
  INV_X1 U10689 ( .A(n16001), .ZN(n4516) );
  OAI21_X1 U10690 ( .B1(n13055), .B2(n13054), .A(n4517), .ZN(n12484) );
  OR2_X1 U10691 ( .A1(n13053), .A2(n13055), .ZN(n12753) );
  NAND2_X1 U10693 ( .A1(n4523), .A2(n4522), .ZN(n9811) );
  NAND2_X1 U10694 ( .A1(n9789), .A2(n9788), .ZN(n4523) );
  NAND2_X1 U10695 ( .A1(n13901), .A2(n4525), .ZN(n4524) );
  NOR2_X1 U10698 ( .A1(n10244), .A2(n10799), .ZN(n10804) );
  NAND3_X1 U10699 ( .A1(n10651), .A2(n10800), .A3(n4527), .ZN(n10248) );
  NAND3_X1 U10700 ( .A1(n10244), .A2(n10651), .A3(n4527), .ZN(n9966) );
  AOI21_X1 U10701 ( .B1(n411), .B2(n4527), .A(n10805), .ZN(n10428) );
  NAND2_X1 U10702 ( .A1(n5427), .A2(n20269), .ZN(n20230) );
  NOR2_X1 U10703 ( .A1(n16845), .A2(n16846), .ZN(n4528) );
  INV_X1 U10704 ( .A(n13353), .ZN(n5626) );
  AND2_X1 U10705 ( .A1(n5626), .A2(n5624), .ZN(n5625) );
  NOR2_X1 U10706 ( .A1(n4531), .A2(n11044), .ZN(n4530) );
  INV_X1 U10707 ( .A(n11051), .ZN(n4531) );
  OAI21_X1 U10708 ( .B1(n11046), .B2(n2680), .A(n4532), .ZN(n11047) );
  MUX2_X1 U10709 ( .A(n11046), .B(n11045), .S(n11044), .Z(n10418) );
  NAND2_X1 U10711 ( .A1(n7867), .A2(n7862), .ZN(n4534) );
  NAND2_X1 U10713 ( .A1(n22832), .A2(n22936), .ZN(n4609) );
  XNOR2_X1 U10714 ( .A(n12200), .B(n12201), .ZN(n12202) );
  INV_X1 U10716 ( .A(n19386), .ZN(n4543) );
  NAND2_X2 U10717 ( .A1(n4544), .A2(n6569), .ZN(n7923) );
  OAI21_X1 U10718 ( .B1(n13219), .B2(n13220), .A(n4546), .ZN(n4548) );
  NOR2_X1 U10719 ( .A1(n4052), .A2(n18808), .ZN(n4551) );
  INV_X1 U10720 ( .A(n18808), .ZN(n5134) );
  INV_X1 U10722 ( .A(n16795), .ZN(n4554) );
  NOR2_X1 U10724 ( .A1(n4553), .A2(n16551), .ZN(n4552) );
  XNOR2_X1 U10725 ( .A(n4556), .B(n14430), .ZN(n15308) );
  INV_X1 U10726 ( .A(n15303), .ZN(n4556) );
  XNOR2_X1 U10727 ( .A(n4557), .B(n14430), .ZN(n13499) );
  XNOR2_X1 U10728 ( .A(n3990), .B(n18579), .ZN(n18581) );
  NAND2_X1 U10729 ( .A1(n17596), .A2(n17597), .ZN(n4563) );
  AND2_X1 U10730 ( .A1(n17600), .A2(n2968), .ZN(n4566) );
  NOR2_X1 U10731 ( .A1(n4567), .A2(n13335), .ZN(n4822) );
  XNOR2_X2 U10732 ( .A(n4820), .B(n4568), .ZN(n13335) );
  INV_X1 U10733 ( .A(n13341), .ZN(n4567) );
  NAND3_X2 U10734 ( .A1(n4570), .A2(n18913), .A3(n4569), .ZN(n21678) );
  INV_X1 U10736 ( .A(n20125), .ZN(n20545) );
  NAND2_X1 U10738 ( .A1(n17226), .A2(n17227), .ZN(n4573) );
  AOI21_X2 U10739 ( .B1(n4576), .B2(n10459), .A(n10458), .ZN(n11653) );
  MUX2_X1 U10740 ( .A(n10730), .B(n10734), .S(n11190), .Z(n4576) );
  NAND2_X1 U10741 ( .A1(n19420), .A2(n19418), .ZN(n19168) );
  XNOR2_X1 U10742 ( .A(n14654), .B(n14799), .ZN(n4582) );
  XNOR2_X1 U10743 ( .A(n14599), .B(n14909), .ZN(n4583) );
  AOI21_X1 U10744 ( .B1(n24499), .B2(n403), .A(n1324), .ZN(n13175) );
  NAND3_X1 U10745 ( .A1(n12727), .A2(n12726), .A3(n4584), .ZN(n13975) );
  NAND2_X1 U10746 ( .A1(n13178), .A2(n12506), .ZN(n4584) );
  MUX2_X1 U10747 ( .A(n12652), .B(n12651), .S(n12506), .Z(n13668) );
  NAND2_X1 U10748 ( .A1(n19501), .A2(n19500), .ZN(n4585) );
  NAND2_X1 U10749 ( .A1(n4586), .A2(n10148), .ZN(n5355) );
  AOI21_X1 U10750 ( .B1(n3317), .B2(n17390), .A(n3604), .ZN(n16875) );
  NAND2_X1 U10751 ( .A1(n25465), .A2(n17185), .ZN(n17390) );
  NAND2_X1 U10752 ( .A1(n15880), .A2(n24385), .ZN(n15635) );
  OR2_X1 U10753 ( .A1(n7155), .A2(n4588), .ZN(n7912) );
  NAND2_X1 U10754 ( .A1(n5636), .A2(n5635), .ZN(n4588) );
  XNOR2_X1 U10756 ( .A(n10771), .B(n11913), .ZN(n10564) );
  XNOR2_X1 U10757 ( .A(n10771), .B(n4589), .ZN(n9217) );
  XNOR2_X1 U10758 ( .A(n4590), .B(n11582), .ZN(n11512) );
  NAND2_X1 U10759 ( .A1(n3653), .A2(n19300), .ZN(n18932) );
  INV_X1 U10760 ( .A(n22406), .ZN(n4591) );
  XNOR2_X1 U10761 ( .A(n15054), .B(n14500), .ZN(n15267) );
  NAND2_X1 U10762 ( .A1(n13364), .A2(n13363), .ZN(n4595) );
  NAND2_X1 U10763 ( .A1(n12977), .A2(n13365), .ZN(n4596) );
  INV_X1 U10764 ( .A(n24503), .ZN(n4597) );
  NAND2_X1 U10765 ( .A1(n4602), .A2(n19014), .ZN(n4601) );
  NAND2_X1 U10767 ( .A1(n25489), .A2(n24407), .ZN(n4602) );
  NAND2_X1 U10770 ( .A1(n23370), .A2(n24404), .ZN(n22991) );
  NAND3_X1 U10771 ( .A1(n23370), .A2(n24404), .A3(n4606), .ZN(n4607) );
  INV_X1 U10772 ( .A(n23379), .ZN(n4606) );
  NAND2_X1 U10773 ( .A1(n4609), .A2(n4608), .ZN(n21657) );
  XNOR2_X1 U10774 ( .A(n11435), .B(n11665), .ZN(n4610) );
  INV_X1 U10775 ( .A(n11665), .ZN(n11764) );
  XNOR2_X1 U10776 ( .A(n9217), .B(n11061), .ZN(n4611) );
  XNOR2_X1 U10777 ( .A(n18540), .B(n18080), .ZN(n18183) );
  NAND2_X1 U10779 ( .A1(n16893), .A2(n17481), .ZN(n4613) );
  NAND2_X1 U10780 ( .A1(n16739), .A2(n16578), .ZN(n16740) );
  INV_X1 U10781 ( .A(n15873), .ZN(n16739) );
  INV_X1 U10782 ( .A(n20140), .ZN(n4616) );
  NOR2_X1 U10783 ( .A1(n5269), .A2(n16217), .ZN(n4617) );
  AND2_X1 U10784 ( .A1(n16219), .A2(n15921), .ZN(n16217) );
  NOR2_X1 U10785 ( .A1(n10149), .A2(n25486), .ZN(n5357) );
  NAND3_X1 U10786 ( .A1(n6314), .A2(n4620), .A3(n6470), .ZN(n4619) );
  NAND2_X1 U10788 ( .A1(n9857), .A2(n239), .ZN(n4622) );
  NAND2_X1 U10790 ( .A1(n4625), .A2(n44), .ZN(n10796) );
  AOI22_X1 U10791 ( .A1(n24526), .A2(n11199), .B1(n4625), .B2(n11201), .ZN(
        n11202) );
  NAND2_X1 U10792 ( .A1(n23160), .A2(n24325), .ZN(n4626) );
  INV_X1 U10795 ( .A(n22424), .ZN(n4632) );
  XNOR2_X1 U10796 ( .A(n15269), .B(n4636), .ZN(n4635) );
  XNOR2_X1 U10797 ( .A(n14721), .B(n15055), .ZN(n15269) );
  XNOR2_X1 U10798 ( .A(n15268), .B(n15267), .ZN(n4637) );
  INV_X1 U10799 ( .A(n12797), .ZN(n4640) );
  NAND2_X1 U10800 ( .A1(n13792), .A2(n13795), .ZN(n14181) );
  NAND2_X1 U10801 ( .A1(n4644), .A2(n7022), .ZN(n4642) );
  INV_X1 U10802 ( .A(n7266), .ZN(n7193) );
  NOR2_X1 U10803 ( .A1(n442), .A2(n4643), .ZN(n4644) );
  NAND2_X1 U10804 ( .A1(n4645), .A2(n4646), .ZN(n17368) );
  NAND2_X1 U10805 ( .A1(n19201), .A2(n4647), .ZN(n19843) );
  XNOR2_X2 U10810 ( .A(n21682), .B(n21683), .ZN(n22901) );
  NAND2_X1 U10811 ( .A1(n4651), .A2(n24513), .ZN(n12987) );
  NAND2_X1 U10813 ( .A1(n13220), .A2(n24513), .ZN(n4652) );
  NAND2_X1 U10814 ( .A1(n17896), .A2(n19479), .ZN(n4653) );
  NAND2_X1 U10815 ( .A1(n20117), .A2(n20109), .ZN(n20113) );
  OAI22_X1 U10816 ( .A1(n11081), .A2(n10766), .B1(n3119), .B2(n4654), .ZN(
        n10770) );
  NAND2_X1 U10817 ( .A1(n4656), .A2(n309), .ZN(n4655) );
  XNOR2_X1 U10818 ( .A(n4657), .B(n21023), .ZN(n21026) );
  OAI21_X1 U10819 ( .B1(n17124), .B2(n17123), .A(n4664), .ZN(n4658) );
  OAI21_X1 U10820 ( .B1(n17124), .B2(n4663), .A(n4658), .ZN(n17587) );
  NAND2_X1 U10821 ( .A1(n4661), .A2(n4659), .ZN(n18430) );
  NAND3_X1 U10822 ( .A1(n17117), .A2(n17824), .A3(n4660), .ZN(n4659) );
  INV_X1 U10823 ( .A(n17123), .ZN(n4660) );
  XNOR2_X1 U10824 ( .A(n4665), .B(n18049), .ZN(n4667) );
  XNOR2_X1 U10825 ( .A(n4666), .B(n17588), .ZN(n4665) );
  XNOR2_X1 U10827 ( .A(n4670), .B(n4669), .ZN(n12192) );
  INV_X1 U10828 ( .A(n2746), .ZN(n4669) );
  NAND2_X1 U10829 ( .A1(n7942), .A2(n4672), .ZN(n7944) );
  NAND2_X1 U10830 ( .A1(n6889), .A2(n6888), .ZN(n4673) );
  NAND2_X1 U10831 ( .A1(n6887), .A2(n6886), .ZN(n4674) );
  NAND2_X1 U10832 ( .A1(n16106), .A2(n16109), .ZN(n4678) );
  XNOR2_X1 U10833 ( .A(n18560), .B(n18464), .ZN(n4679) );
  INV_X1 U10834 ( .A(n18560), .ZN(n18130) );
  NAND2_X1 U10835 ( .A1(n4680), .A2(n12993), .ZN(n12890) );
  NAND2_X1 U10836 ( .A1(n6526), .A2(n6952), .ZN(n4682) );
  OAI211_X1 U10837 ( .C1(n4684), .C2(n17130), .A(n17134), .B(n25226), .ZN(
        n4683) );
  INV_X1 U10839 ( .A(n17134), .ZN(n4686) );
  NAND2_X1 U10841 ( .A1(n24407), .A2(n18788), .ZN(n18443) );
  NAND2_X1 U10843 ( .A1(n5149), .A2(n19395), .ZN(n5501) );
  INV_X1 U10844 ( .A(n10992), .ZN(n4691) );
  NAND2_X1 U10846 ( .A1(n6053), .A2(n5775), .ZN(n4694) );
  INV_X1 U10847 ( .A(n5774), .ZN(n6409) );
  INV_X1 U10848 ( .A(n6744), .ZN(n4696) );
  NAND2_X1 U10849 ( .A1(n5777), .A2(n6628), .ZN(n4697) );
  NAND4_X1 U10850 ( .A1(n4699), .A2(n4698), .A3(n4704), .A4(n2744), .ZN(n4702)
         );
  INV_X1 U10851 ( .A(n22999), .ZN(n4698) );
  INV_X1 U10852 ( .A(n23000), .ZN(n4699) );
  OAI21_X1 U10853 ( .B1(n4701), .B2(n22999), .A(n444), .ZN(n4700) );
  INV_X1 U10854 ( .A(n4704), .ZN(n4701) );
  NAND2_X1 U10855 ( .A1(n23000), .A2(n444), .ZN(n4703) );
  NAND3_X1 U10856 ( .A1(n22749), .A2(n22998), .A3(n1442), .ZN(n4704) );
  OAI21_X1 U10857 ( .B1(n10095), .B2(n10098), .A(n8359), .ZN(n8384) );
  INV_X1 U10858 ( .A(n8351), .ZN(n4705) );
  OAI211_X1 U10860 ( .C1(n8352), .C2(n4711), .A(n4710), .B(n4709), .ZN(n8354)
         );
  NAND2_X1 U10861 ( .A1(n16418), .A2(n16408), .ZN(n15866) );
  XNOR2_X1 U10862 ( .A(n14729), .B(n14444), .ZN(n4712) );
  NAND2_X1 U10864 ( .A1(n5774), .A2(n6050), .ZN(n6052) );
  NAND2_X1 U10865 ( .A1(n5774), .A2(n6744), .ZN(n6629) );
  NAND2_X1 U10866 ( .A1(n5774), .A2(n6630), .ZN(n5775) );
  NAND2_X1 U10867 ( .A1(n6628), .A2(n5774), .ZN(n6748) );
  NAND3_X1 U10868 ( .A1(n6051), .A2(n5774), .A3(n4696), .ZN(n6410) );
  AOI21_X1 U10869 ( .B1(n6566), .B2(n6746), .A(n5774), .ZN(n7927) );
  NAND2_X1 U10870 ( .A1(n20301), .A2(n20009), .ZN(n19049) );
  MUX2_X1 U10871 ( .A(n14458), .B(n3404), .S(n3401), .Z(n14318) );
  NAND2_X1 U10872 ( .A1(n24079), .A2(n4715), .ZN(n4716) );
  NAND2_X1 U10873 ( .A1(n5439), .A2(n24079), .ZN(n4717) );
  XNOR2_X1 U10874 ( .A(n18041), .B(n18040), .ZN(n19071) );
  NAND2_X1 U10875 ( .A1(n4720), .A2(n4718), .ZN(n23425) );
  OAI22_X1 U10876 ( .A1(n22528), .A2(n23425), .B1(n1370), .B2(n23442), .ZN(
        n23453) );
  XNOR2_X1 U10877 ( .A(n4723), .B(n14579), .ZN(n14840) );
  NOR2_X2 U10878 ( .A1(n4722), .A2(n4721), .ZN(n14579) );
  AOI21_X1 U10879 ( .B1(n12818), .B2(n14172), .A(n13526), .ZN(n4722) );
  NAND3_X1 U10880 ( .A1(n16461), .A2(n16462), .A3(n16460), .ZN(n4725) );
  OAI211_X2 U10881 ( .C1(n9453), .C2(n9935), .A(n9451), .B(n9452), .ZN(n10885)
         );
  NAND2_X1 U10883 ( .A1(n6429), .A2(n6785), .ZN(n4727) );
  NAND3_X1 U10884 ( .A1(n25242), .A2(n20136), .A3(n4728), .ZN(n19756) );
  NAND2_X1 U10885 ( .A1(n5566), .A2(n4728), .ZN(n5565) );
  AOI21_X1 U10886 ( .B1(n20135), .B2(n4728), .A(n19755), .ZN(n19758) );
  NAND2_X1 U10887 ( .A1(n5436), .A2(n4729), .ZN(n12862) );
  OAI21_X1 U10888 ( .B1(n10759), .B2(n10757), .A(n10756), .ZN(n4733) );
  XNOR2_X2 U10889 ( .A(n5981), .B(Key[125]), .ZN(n7007) );
  NAND3_X1 U10890 ( .A1(n15130), .A2(n4735), .A3(n4734), .ZN(n17381) );
  NAND2_X1 U10891 ( .A1(n15118), .A2(n24919), .ZN(n4734) );
  OAI21_X1 U10892 ( .B1(n1434), .B2(n15117), .A(n24841), .ZN(n4735) );
  NOR2_X1 U10893 ( .A1(n10985), .A2(n10552), .ZN(n4736) );
  NAND2_X1 U10894 ( .A1(n10554), .A2(n4737), .ZN(n4739) );
  NOR2_X1 U10896 ( .A1(n11160), .A2(n11163), .ZN(n10553) );
  NOR2_X2 U10897 ( .A1(n4740), .A2(n4738), .ZN(n11761) );
  MUX2_X1 U10898 ( .A(n24490), .B(n13222), .S(n24965), .Z(n4741) );
  NAND2_X1 U10899 ( .A1(n17426), .A2(n17379), .ZN(n4742) );
  NAND2_X1 U10900 ( .A1(n4745), .A2(n25014), .ZN(n4744) );
  NAND2_X1 U10901 ( .A1(n4746), .A2(n4747), .ZN(n4745) );
  NAND2_X1 U10902 ( .A1(n6530), .A2(n24067), .ZN(n4747) );
  XNOR2_X2 U10903 ( .A(Key[27]), .B(Plaintext[27]), .ZN(n6530) );
  NOR2_X1 U10904 ( .A1(n19500), .A2(n4748), .ZN(n18720) );
  NOR2_X1 U10905 ( .A1(n19502), .A2(n3296), .ZN(n18983) );
  NAND2_X1 U10906 ( .A1(n19497), .A2(n3296), .ZN(n19495) );
  OAI21_X1 U10907 ( .B1(n19335), .B2(n19500), .A(n3296), .ZN(n17924) );
  AOI21_X1 U10908 ( .B1(n18987), .B2(n17938), .A(n4748), .ZN(n17939) );
  NAND3_X1 U10910 ( .A1(n20236), .A2(n20170), .A3(n20239), .ZN(n4750) );
  NAND2_X1 U10912 ( .A1(n5802), .A2(n5801), .ZN(n4753) );
  NAND2_X1 U10913 ( .A1(n14157), .A2(n14156), .ZN(n14163) );
  XNOR2_X1 U10915 ( .A(n4759), .B(n11838), .ZN(n12239) );
  OAI211_X2 U10916 ( .C1(n10550), .C2(n3509), .A(n10551), .B(n4758), .ZN(
        n11838) );
  NOR2_X1 U10918 ( .A1(n5376), .A2(n16796), .ZN(n4760) );
  OAI21_X1 U10919 ( .B1(n19597), .B2(n19598), .A(n19255), .ZN(n19075) );
  MUX2_X1 U10920 ( .A(n19255), .B(n19596), .S(n19597), .Z(n18054) );
  NAND2_X1 U10921 ( .A1(n4764), .A2(n24919), .ZN(n15897) );
  NAND2_X1 U10922 ( .A1(n15748), .A2(n16293), .ZN(n4764) );
  NAND2_X1 U10923 ( .A1(n16357), .A2(n16356), .ZN(n15748) );
  NOR2_X1 U10924 ( .A1(n4766), .A2(n13170), .ZN(n12720) );
  NOR2_X1 U10925 ( .A1(n4766), .A2(n13165), .ZN(n13166) );
  XNOR2_X2 U10926 ( .A(n18180), .B(n18179), .ZN(n19522) );
  OR2_X1 U10927 ( .A1(n14278), .A2(n24572), .ZN(n4771) );
  NAND3_X1 U10928 ( .A1(n4225), .A2(n14850), .A3(n4767), .ZN(n4769) );
  XNOR2_X1 U10929 ( .A(n14980), .B(n14789), .ZN(n15338) );
  NAND2_X1 U10932 ( .A1(n14416), .A2(n13617), .ZN(n4770) );
  NAND2_X1 U10933 ( .A1(n16484), .A2(n16481), .ZN(n4772) );
  INV_X1 U10934 ( .A(n25218), .ZN(n4775) );
  NAND2_X1 U10937 ( .A1(n24927), .A2(n262), .ZN(n7572) );
  INV_X1 U10938 ( .A(n10518), .ZN(n4779) );
  OAI211_X1 U10939 ( .C1(n10520), .C2(n10829), .A(n4778), .B(n4777), .ZN(
        n10279) );
  NAND2_X1 U10940 ( .A1(n10830), .A2(n10275), .ZN(n10520) );
  NAND2_X1 U10941 ( .A1(n19838), .A2(n20194), .ZN(n4780) );
  NAND2_X1 U10942 ( .A1(n25078), .A2(n22093), .ZN(n4781) );
  INV_X1 U10943 ( .A(n4781), .ZN(n21772) );
  OAI211_X1 U10944 ( .C1(n22642), .C2(n22641), .A(n22640), .B(n4782), .ZN(
        Ciphertext[118]) );
  MUX2_X1 U10946 ( .A(n7660), .B(n7659), .S(n7947), .Z(n4785) );
  AOI22_X1 U10947 ( .A1(n9695), .A2(n10026), .B1(n9699), .B2(n9639), .ZN(n4787) );
  OAI21_X2 U10948 ( .B1(n4787), .B2(n9240), .A(n9239), .ZN(n11123) );
  NAND3_X1 U10950 ( .A1(n4794), .A2(n14317), .A3(n13868), .ZN(n4793) );
  NAND2_X1 U10951 ( .A1(n14322), .A2(n14458), .ZN(n4795) );
  NAND2_X2 U10952 ( .A1(n5172), .A2(n5170), .ZN(n14317) );
  NAND2_X1 U10953 ( .A1(n12870), .A2(n13097), .ZN(n4796) );
  NAND2_X1 U10954 ( .A1(n12867), .A2(n13117), .ZN(n4797) );
  NAND2_X1 U10955 ( .A1(n4800), .A2(n7739), .ZN(n4799) );
  INV_X1 U10957 ( .A(n8913), .ZN(n4802) );
  OAI211_X2 U10958 ( .C1(n4801), .C2(n7820), .A(n6799), .B(n7821), .ZN(n8913)
         );
  NAND2_X1 U10959 ( .A1(n8219), .A2(n7809), .ZN(n4804) );
  NAND2_X1 U10961 ( .A1(n14702), .A2(n24586), .ZN(n4806) );
  OAI22_X1 U10964 ( .A1(n19016), .A2(n19162), .B1(n19164), .B2(n4809), .ZN(
        n18791) );
  XNOR2_X1 U10965 ( .A(n18434), .B(n18478), .ZN(n4810) );
  XNOR2_X1 U10967 ( .A(n18441), .B(n18440), .ZN(n19163) );
  NAND2_X1 U10968 ( .A1(n7229), .A2(n7946), .ZN(n4813) );
  INV_X1 U10970 ( .A(n10553), .ZN(n4815) );
  NAND2_X1 U10971 ( .A1(n16830), .A2(n17445), .ZN(n4818) );
  NAND2_X1 U10972 ( .A1(n12957), .A2(n13336), .ZN(n4823) );
  XNOR2_X1 U10973 ( .A(n4821), .B(n12105), .ZN(n4820) );
  INV_X1 U10974 ( .A(n12106), .ZN(n4821) );
  NAND2_X1 U10975 ( .A1(n11022), .A2(n13775), .ZN(n4824) );
  INV_X1 U10976 ( .A(n7358), .ZN(n7415) );
  NAND2_X1 U10977 ( .A1(n4827), .A2(n7358), .ZN(n7994) );
  OR2_X1 U10978 ( .A1(n6690), .A2(n6686), .ZN(n4830) );
  INV_X1 U10979 ( .A(n9423), .ZN(n9746) );
  NAND2_X1 U10982 ( .A1(n4833), .A2(n9747), .ZN(n4832) );
  AND2_X1 U10983 ( .A1(n9991), .A2(n9990), .ZN(n4833) );
  OAI21_X1 U10985 ( .B1(n16383), .B2(n15656), .A(n4835), .ZN(n16387) );
  OAI22_X2 U10987 ( .A1(n4837), .A2(n14236), .B1(n13994), .B2(n13930), .ZN(
        n15112) );
  NAND2_X1 U10988 ( .A1(n7022), .A2(n6846), .ZN(n4839) );
  NAND3_X1 U10989 ( .A1(n6001), .A2(n250), .A3(n4839), .ZN(n4838) );
  AOI21_X1 U10990 ( .B1(n16316), .B2(n17013), .A(n4840), .ZN(n16317) );
  INV_X1 U10991 ( .A(n17356), .ZN(n4840) );
  OAI21_X1 U10992 ( .B1(n19077), .B2(n24483), .A(n4843), .ZN(n4842) );
  NAND2_X1 U10993 ( .A1(n24483), .A2(n19078), .ZN(n4843) );
  INV_X1 U10994 ( .A(n21812), .ZN(n4845) );
  NAND2_X1 U10995 ( .A1(n22059), .A2(n22245), .ZN(n21812) );
  NOR2_X1 U10996 ( .A1(n21786), .A2(n4845), .ZN(n21788) );
  NOR2_X1 U10998 ( .A1(n7382), .A2(n7619), .ZN(n4848) );
  OAI211_X2 U10999 ( .C1(n4848), .C2(n7304), .A(n7303), .B(n7302), .ZN(n8916)
         );
  INV_X1 U11000 ( .A(n12534), .ZN(n4850) );
  NAND3_X1 U11001 ( .A1(n401), .A2(n13051), .A3(n12534), .ZN(n12443) );
  NAND2_X1 U11002 ( .A1(n19211), .A2(n4853), .ZN(n4852) );
  INV_X1 U11004 ( .A(n4854), .ZN(n23762) );
  NAND2_X1 U11005 ( .A1(n23767), .A2(n23769), .ZN(n4854) );
  OAI22_X1 U11006 ( .A1(n23783), .A2(n22523), .B1(n22524), .B2(n4854), .ZN(
        n22526) );
  INV_X1 U11007 ( .A(n23769), .ZN(n23778) );
  XNOR2_X1 U11008 ( .A(n18381), .B(n4855), .ZN(n16664) );
  XNOR2_X1 U11009 ( .A(n18381), .B(n4856), .ZN(n18013) );
  INV_X1 U11010 ( .A(n18183), .ZN(n4856) );
  NAND2_X1 U11011 ( .A1(n19210), .A2(n18816), .ZN(n4857) );
  XNOR2_X1 U11012 ( .A(n15282), .B(n15174), .ZN(n4859) );
  NAND3_X1 U11014 ( .A1(n23723), .A2(n23714), .A3(n23727), .ZN(n4864) );
  NAND2_X1 U11015 ( .A1(n23721), .A2(n23720), .ZN(n22148) );
  XNOR2_X1 U11016 ( .A(n4862), .B(n22150), .ZN(Ciphertext[135]) );
  NAND2_X1 U11017 ( .A1(n438), .A2(n6295), .ZN(n6211) );
  MUX2_X1 U11018 ( .A(n5946), .B(n6173), .S(n6174), .Z(n5948) );
  NAND2_X1 U11019 ( .A1(n16202), .A2(n16200), .ZN(n4870) );
  MUX2_X1 U11020 ( .A(n11205), .B(n11338), .S(n11209), .Z(n9645) );
  NAND2_X1 U11023 ( .A1(n264), .A2(n18841), .ZN(n4874) );
  NAND2_X1 U11024 ( .A1(n6174), .A2(n6335), .ZN(n6176) );
  NAND2_X1 U11026 ( .A1(n9880), .A2(n4993), .ZN(n9252) );
  NAND2_X1 U11028 ( .A1(n4878), .A2(n4881), .ZN(n4880) );
  OAI21_X1 U11029 ( .B1(n7647), .B2(n7761), .A(n4879), .ZN(n7766) );
  NAND2_X1 U11030 ( .A1(n7646), .A2(n4880), .ZN(n4879) );
  XNOR2_X1 U11031 ( .A(n18704), .B(n4882), .ZN(n17035) );
  XNOR2_X1 U11032 ( .A(n17900), .B(n17817), .ZN(n4882) );
  INV_X1 U11033 ( .A(n19237), .ZN(n18863) );
  INV_X1 U11034 ( .A(n19112), .ZN(n4884) );
  INV_X1 U11035 ( .A(n24310), .ZN(n4885) );
  NAND2_X1 U11036 ( .A1(n5446), .A2(n16269), .ZN(n4886) );
  NAND2_X1 U11037 ( .A1(n16270), .A2(n16271), .ZN(n4887) );
  XNOR2_X1 U11038 ( .A(n18123), .B(n18124), .ZN(n18492) );
  XNOR2_X1 U11039 ( .A(n18184), .B(n18492), .ZN(n18127) );
  OAI21_X1 U11040 ( .B1(n7228), .B2(n7080), .A(n7943), .ZN(n4889) );
  XNOR2_X1 U11041 ( .A(n18383), .B(n1410), .ZN(n4890) );
  OAI21_X1 U11042 ( .B1(n25445), .B2(n4892), .A(n4891), .ZN(n4893) );
  NAND2_X1 U11044 ( .A1(n14211), .A2(n24376), .ZN(n4892) );
  AOI21_X2 U11045 ( .B1(n4895), .B2(n1391), .A(n4893), .ZN(n14834) );
  INV_X1 U11046 ( .A(n24375), .ZN(n4894) );
  NAND3_X1 U11047 ( .A1(n16050), .A2(n294), .A3(n15606), .ZN(n4900) );
  AOI21_X1 U11048 ( .B1(n24574), .B2(n11111), .A(n10868), .ZN(n10877) );
  NAND2_X1 U11049 ( .A1(n19704), .A2(n20615), .ZN(n4991) );
  NAND2_X1 U11050 ( .A1(n20616), .A2(n20617), .ZN(n19704) );
  NAND2_X1 U11051 ( .A1(n4902), .A2(n7376), .ZN(n4901) );
  NAND2_X1 U11052 ( .A1(n5432), .A2(n7735), .ZN(n4902) );
  AOI22_X1 U11053 ( .A1(n4904), .A2(n25240), .B1(n23866), .B2(n23857), .ZN(
        n4903) );
  NAND3_X1 U11054 ( .A1(n13093), .A2(n13096), .A3(n12871), .ZN(n4907) );
  NAND2_X1 U11055 ( .A1(n4910), .A2(n4912), .ZN(n4909) );
  NAND2_X1 U11056 ( .A1(n20117), .A2(n25034), .ZN(n4910) );
  INV_X1 U11057 ( .A(n17951), .ZN(n20848) );
  AOI21_X1 U11058 ( .B1(n25262), .B2(n19883), .A(n20109), .ZN(n4912) );
  XNOR2_X1 U11059 ( .A(n9124), .B(n4913), .ZN(n9125) );
  XNOR2_X1 U11060 ( .A(n8236), .B(n4913), .ZN(n5504) );
  XNOR2_X1 U11061 ( .A(n8843), .B(n4913), .ZN(n8833) );
  NAND2_X1 U11062 ( .A1(n15815), .A2(n4914), .ZN(n15818) );
  NAND2_X1 U11063 ( .A1(n4919), .A2(n19532), .ZN(n4915) );
  INV_X1 U11064 ( .A(n19270), .ZN(n19529) );
  NOR2_X1 U11065 ( .A1(n24393), .A2(n4918), .ZN(n4917) );
  INV_X1 U11066 ( .A(n19537), .ZN(n4918) );
  OAI21_X1 U11067 ( .B1(n19530), .B2(n19270), .A(n19269), .ZN(n4919) );
  INV_X1 U11069 ( .A(n6874), .ZN(n4922) );
  NAND2_X1 U11070 ( .A1(n314), .A2(n6767), .ZN(n6878) );
  NAND2_X1 U11071 ( .A1(n6876), .A2(n314), .ZN(n6764) );
  NAND3_X1 U11072 ( .A1(n6309), .A2(n6768), .A3(n314), .ZN(n6312) );
  MUX2_X1 U11073 ( .A(n5855), .B(n5854), .S(n314), .Z(n5858) );
  NOR2_X1 U11075 ( .A1(n10942), .A2(n5392), .ZN(n10513) );
  NOR2_X1 U11076 ( .A1(n10571), .A2(n5392), .ZN(n10572) );
  NAND2_X1 U11077 ( .A1(n13109), .A2(n12856), .ZN(n4925) );
  NAND2_X1 U11078 ( .A1(n13265), .A2(n13267), .ZN(n4930) );
  NOR2_X2 U11079 ( .A1(n19046), .A2(n19045), .ZN(n19979) );
  NAND2_X1 U11080 ( .A1(n19977), .A2(n20140), .ZN(n4933) );
  INV_X1 U11081 ( .A(n17485), .ZN(n17733) );
  NOR2_X1 U11082 ( .A1(n17485), .A2(n4934), .ZN(n17484) );
  NAND2_X1 U11083 ( .A1(n3978), .A2(n23531), .ZN(n23009) );
  NAND3_X1 U11084 ( .A1(n23013), .A2(n23533), .A3(n3978), .ZN(n23024) );
  OR2_X2 U11085 ( .A1(n9402), .A2(n9401), .ZN(n11190) );
  NAND2_X1 U11086 ( .A1(n10457), .A2(n10728), .ZN(n4936) );
  NAND2_X1 U11087 ( .A1(n4951), .A2(n10728), .ZN(n4937) );
  NAND2_X1 U11089 ( .A1(n4353), .A2(n14663), .ZN(n4939) );
  INV_X1 U11090 ( .A(n14267), .ZN(n14274) );
  NAND2_X1 U11092 ( .A1(n12984), .A2(n12541), .ZN(n4944) );
  INV_X1 U11093 ( .A(n13220), .ZN(n4945) );
  INV_X1 U11094 ( .A(n23515), .ZN(n4947) );
  MUX2_X1 U11095 ( .A(n22916), .B(n4948), .S(n22918), .Z(n23515) );
  OAI22_X1 U11096 ( .A1(n21712), .A2(n22918), .B1(n22916), .B2(n22917), .ZN(
        n4950) );
  AND2_X1 U11097 ( .A1(n4951), .A2(n11190), .ZN(n9403) );
  INV_X1 U11098 ( .A(n10730), .ZN(n4951) );
  INV_X1 U11099 ( .A(n4957), .ZN(n16304) );
  OAI22_X1 U11101 ( .A1(n16300), .A2(n16299), .B1(n16303), .B2(n4957), .ZN(
        n16308) );
  NAND2_X1 U11102 ( .A1(n7666), .A2(n436), .ZN(n6551) );
  NAND3_X1 U11103 ( .A1(n7666), .A2(n436), .A3(n269), .ZN(n8533) );
  NAND2_X1 U11104 ( .A1(n12925), .A2(n4958), .ZN(n12609) );
  INV_X1 U11105 ( .A(n12899), .ZN(n4958) );
  OAI21_X1 U11107 ( .B1(n20317), .B2(n4961), .A(n4960), .ZN(n19716) );
  INV_X1 U11108 ( .A(n20316), .ZN(n4961) );
  NAND2_X1 U11109 ( .A1(n12898), .A2(n12897), .ZN(n4964) );
  XNOR2_X1 U11110 ( .A(n14429), .B(n14430), .ZN(n4967) );
  OR2_X1 U11111 ( .A1(n19128), .A2(n19304), .ZN(n4968) );
  XNOR2_X1 U11113 ( .A(n4971), .B(n25481), .ZN(n18173) );
  NAND3_X1 U11114 ( .A1(n16027), .A2(n2062), .A3(n4970), .ZN(n4969) );
  OAI21_X1 U11117 ( .B1(n24089), .B2(n6965), .A(n4973), .ZN(n7184) );
  NAND2_X1 U11118 ( .A1(n19109), .A2(n25052), .ZN(n4977) );
  XNOR2_X1 U11119 ( .A(n21463), .B(n25040), .ZN(n4978) );
  NOR2_X1 U11120 ( .A1(n14168), .A2(n13742), .ZN(n4980) );
  NAND2_X1 U11122 ( .A1(n4982), .A2(n4981), .ZN(n16950) );
  NAND2_X1 U11123 ( .A1(n4984), .A2(n4983), .ZN(n4982) );
  NAND2_X1 U11124 ( .A1(n1382), .A2(n16417), .ZN(n4983) );
  NAND2_X1 U11125 ( .A1(n17289), .A2(n4986), .ZN(n17541) );
  NAND3_X1 U11126 ( .A1(n23079), .A2(n23064), .A3(n25024), .ZN(n4989) );
  NAND2_X1 U11129 ( .A1(n4991), .A2(n24338), .ZN(n19873) );
  NAND2_X1 U11130 ( .A1(n13171), .A2(n3688), .ZN(n4992) );
  INV_X1 U11131 ( .A(n10534), .ZN(n11884) );
  NAND4_X1 U11132 ( .A1(n6808), .A2(n6807), .A3(n6809), .A4(n4994), .ZN(n6810)
         );
  XNOR2_X1 U11133 ( .A(n12106), .B(n11849), .ZN(n4996) );
  NAND2_X1 U11134 ( .A1(n1357), .A2(n10534), .ZN(n10308) );
  NAND2_X1 U11135 ( .A1(n1357), .A2(n4997), .ZN(n10965) );
  AND2_X1 U11136 ( .A1(n10534), .A2(n24479), .ZN(n4997) );
  OR2_X1 U11138 ( .A1(n6392), .A2(n6238), .ZN(n5002) );
  XNOR2_X2 U11139 ( .A(n18210), .B(n18211), .ZN(n19526) );
  NAND2_X1 U11140 ( .A1(n19523), .A2(n19284), .ZN(n5496) );
  NAND2_X1 U11141 ( .A1(n19526), .A2(n19522), .ZN(n5003) );
  INV_X1 U11142 ( .A(n9064), .ZN(n10058) );
  INV_X1 U11143 ( .A(n10052), .ZN(n5004) );
  NAND2_X1 U11144 ( .A1(n19433), .A2(n25423), .ZN(n5006) );
  NAND2_X1 U11145 ( .A1(n19438), .A2(n18834), .ZN(n19433) );
  NAND2_X1 U11147 ( .A1(n21958), .A2(n21959), .ZN(n21961) );
  XNOR2_X1 U11149 ( .A(n295), .B(n15244), .ZN(n5009) );
  NAND2_X1 U11150 ( .A1(n13064), .A2(n5011), .ZN(n5010) );
  XNOR2_X1 U11151 ( .A(n8595), .B(n8594), .ZN(n9481) );
  XNOR2_X1 U11152 ( .A(n5014), .B(n2241), .ZN(n8777) );
  XNOR2_X1 U11153 ( .A(n8446), .B(n5014), .ZN(n8447) );
  XNOR2_X1 U11154 ( .A(n8172), .B(n5014), .ZN(n8174) );
  INV_X1 U11158 ( .A(n14188), .ZN(n5020) );
  OR2_X1 U11160 ( .A1(n12694), .A2(n13292), .ZN(n5021) );
  NAND2_X1 U11161 ( .A1(n19691), .A2(n20316), .ZN(n19692) );
  NAND2_X1 U11163 ( .A1(n12650), .A2(n12505), .ZN(n5022) );
  INV_X1 U11164 ( .A(n17607), .ZN(n16942) );
  NAND2_X1 U11165 ( .A1(n5066), .A2(n5065), .ZN(n5064) );
  NAND2_X1 U11166 ( .A1(n10090), .A2(n24505), .ZN(n5026) );
  MUX2_X1 U11168 ( .A(n13294), .B(n13295), .S(n12827), .Z(n13296) );
  NAND2_X1 U11172 ( .A1(n5033), .A2(n5030), .ZN(n5029) );
  NOR2_X1 U11173 ( .A1(n23089), .A2(n5131), .ZN(n5030) );
  NAND4_X1 U11174 ( .A1(n5035), .A2(n24941), .A3(n20975), .A4(n5037), .ZN(
        n5031) );
  OR2_X1 U11175 ( .A1(n23112), .A2(n24993), .ZN(n5037) );
  NAND3_X1 U11176 ( .A1(n23089), .A2(n24498), .A3(n5131), .ZN(n5032) );
  NAND2_X1 U11177 ( .A1(n5040), .A2(n5038), .ZN(n16486) );
  NAND2_X1 U11178 ( .A1(n16482), .A2(n15951), .ZN(n5040) );
  AND2_X1 U11179 ( .A1(n13231), .A2(n5041), .ZN(n13232) );
  NAND2_X1 U11180 ( .A1(n9443), .A2(n10584), .ZN(n5042) );
  NAND2_X1 U11181 ( .A1(n5042), .A2(n10317), .ZN(n10319) );
  OAI22_X1 U11182 ( .A1(n5042), .A2(n25507), .B1(n10370), .B2(n10372), .ZN(
        n9215) );
  OAI211_X1 U11183 ( .C1(n20426), .C2(n276), .A(n24883), .B(n5044), .ZN(n5043)
         );
  OR2_X1 U11186 ( .A1(n22592), .A2(n22317), .ZN(n5046) );
  NAND2_X1 U11187 ( .A1(n21378), .A2(n274), .ZN(n5047) );
  NAND3_X1 U11189 ( .A1(n23143), .A2(n1349), .A3(n22442), .ZN(n5049) );
  NAND2_X1 U11190 ( .A1(n7129), .A2(n7606), .ZN(n5050) );
  INV_X1 U11191 ( .A(n7893), .ZN(n5051) );
  NOR2_X1 U11192 ( .A1(n16844), .A2(n5052), .ZN(n17467) );
  NAND2_X1 U11193 ( .A1(n5054), .A2(n5051), .ZN(n5053) );
  NAND2_X1 U11194 ( .A1(n7609), .A2(n7604), .ZN(n7889) );
  NAND2_X1 U11195 ( .A1(n7894), .A2(n7893), .ZN(n5055) );
  NOR2_X1 U11196 ( .A1(n5056), .A2(n17130), .ZN(n17129) );
  INV_X1 U11197 ( .A(n25225), .ZN(n5056) );
  NOR2_X1 U11199 ( .A1(n10487), .A2(n10486), .ZN(n5060) );
  NAND2_X1 U11200 ( .A1(n10488), .A2(n5060), .ZN(n5059) );
  NAND2_X1 U11201 ( .A1(n5730), .A2(n10614), .ZN(n5061) );
  NAND2_X1 U11202 ( .A1(n10531), .A2(n304), .ZN(n5063) );
  NAND3_X1 U11203 ( .A1(n10465), .A2(n10855), .A3(n10858), .ZN(n10466) );
  NAND2_X1 U11204 ( .A1(n9456), .A2(n9565), .ZN(n5065) );
  NOR2_X1 U11206 ( .A1(n16832), .A2(n17152), .ZN(n16834) );
  NAND2_X1 U11210 ( .A1(n18734), .A2(n19477), .ZN(n5070) );
  OAI21_X1 U11211 ( .B1(n20173), .B2(n19803), .A(n5071), .ZN(n19508) );
  NAND2_X1 U11212 ( .A1(n19507), .A2(n20173), .ZN(n5071) );
  NAND2_X1 U11213 ( .A1(n5072), .A2(n16980), .ZN(n5073) );
  INV_X1 U11214 ( .A(n17450), .ZN(n5072) );
  INV_X1 U11216 ( .A(n23765), .ZN(n23766) );
  NAND2_X1 U11217 ( .A1(n23779), .A2(n23757), .ZN(n23765) );
  NAND2_X1 U11219 ( .A1(n21793), .A2(n22231), .ZN(n5076) );
  NAND2_X1 U11220 ( .A1(n5077), .A2(n1481), .ZN(n5078) );
  NAND2_X1 U11221 ( .A1(n5078), .A2(n11127), .ZN(n12219) );
  NAND2_X1 U11222 ( .A1(n13953), .A2(n13954), .ZN(n5079) );
  INV_X1 U11223 ( .A(n13954), .ZN(n5080) );
  NAND2_X1 U11224 ( .A1(n395), .A2(n13953), .ZN(n13718) );
  NAND2_X1 U11225 ( .A1(n14156), .A2(n395), .ZN(n13719) );
  NAND2_X1 U11226 ( .A1(n5081), .A2(n23256), .ZN(n22649) );
  NAND2_X1 U11227 ( .A1(n425), .A2(n25454), .ZN(n9298) );
  OR2_X1 U11228 ( .A1(n5082), .A2(n1348), .ZN(n8574) );
  NAND2_X1 U11229 ( .A1(n5083), .A2(n10089), .ZN(n10091) );
  NAND2_X1 U11230 ( .A1(n9779), .A2(n8571), .ZN(n5083) );
  OAI21_X1 U11231 ( .B1(n9780), .B2(n25454), .A(n425), .ZN(n9674) );
  INV_X1 U11232 ( .A(n5084), .ZN(n21885) );
  NAND2_X1 U11233 ( .A1(n5084), .A2(n22396), .ZN(n22267) );
  NOR2_X1 U11234 ( .A1(n22261), .A2(n5084), .ZN(n22264) );
  AOI21_X1 U11235 ( .B1(n22398), .B2(n5084), .A(n22265), .ZN(n21914) );
  MUX2_X1 U11236 ( .A(n22400), .B(n5084), .S(n25381), .Z(n22136) );
  AND2_X1 U11237 ( .A1(n7023), .A2(n7025), .ZN(n5088) );
  NAND2_X1 U11238 ( .A1(n5089), .A2(n7027), .ZN(n5086) );
  XNOR2_X1 U11241 ( .A(n18290), .B(n24886), .ZN(n17792) );
  XNOR2_X1 U11242 ( .A(n24886), .B(n2319), .ZN(n18460) );
  NAND2_X1 U11243 ( .A1(n10772), .A2(n11101), .ZN(n10218) );
  NAND2_X1 U11244 ( .A1(n11031), .A2(n10772), .ZN(n11034) );
  OAI22_X1 U11245 ( .A1(n1552), .A2(n10772), .B1(n24753), .B2(n415), .ZN(
        n11035) );
  NAND2_X1 U11246 ( .A1(n23194), .A2(n24889), .ZN(n5090) );
  INV_X1 U11247 ( .A(n11684), .ZN(n12891) );
  NAND2_X1 U11248 ( .A1(n19442), .A2(n20588), .ZN(n5091) );
  NAND2_X1 U11249 ( .A1(n5094), .A2(n5093), .ZN(n5092) );
  AND3_X2 U11251 ( .A1(n5670), .A2(n19416), .A3(n5669), .ZN(n20586) );
  NAND3_X1 U11252 ( .A1(n5218), .A2(n23974), .A3(n5095), .ZN(n5217) );
  NAND2_X1 U11253 ( .A1(n1488), .A2(n24440), .ZN(n5095) );
  NAND2_X1 U11254 ( .A1(n5098), .A2(n5096), .ZN(n16234) );
  NOR2_X1 U11255 ( .A1(n16491), .A2(n16232), .ZN(n5097) );
  NAND2_X1 U11256 ( .A1(n16233), .A2(n16232), .ZN(n5098) );
  NAND2_X1 U11258 ( .A1(n5100), .A2(n16100), .ZN(n16104) );
  NAND2_X1 U11261 ( .A1(n15576), .A2(n5104), .ZN(n5103) );
  OAI211_X1 U11262 ( .C1(n10699), .C2(n2754), .A(n5109), .B(n10955), .ZN(n5108) );
  NAND2_X1 U11263 ( .A1(n10699), .A2(n10548), .ZN(n5109) );
  NAND2_X1 U11264 ( .A1(n5111), .A2(n5110), .ZN(n14172) );
  NAND2_X1 U11265 ( .A1(n5113), .A2(n5112), .ZN(n5110) );
  NAND2_X1 U11266 ( .A1(n12441), .A2(n12737), .ZN(n5111) );
  NAND2_X1 U11268 ( .A1(n5115), .A2(n20060), .ZN(n5114) );
  NOR2_X1 U11270 ( .A1(n7221), .A2(n5117), .ZN(n5116) );
  INV_X1 U11271 ( .A(n7222), .ZN(n5117) );
  NAND2_X1 U11273 ( .A1(n11062), .A2(n11070), .ZN(n5119) );
  XNOR2_X1 U11274 ( .A(n5120), .B(n2743), .ZN(n18570) );
  XNOR2_X1 U11275 ( .A(n5120), .B(n18295), .ZN(n18087) );
  XNOR2_X1 U11276 ( .A(n5120), .B(n18188), .ZN(n15810) );
  NAND2_X1 U11277 ( .A1(n13227), .A2(n13224), .ZN(n13225) );
  INV_X1 U11278 ( .A(n25367), .ZN(n20822) );
  NOR2_X1 U11279 ( .A1(n20803), .A2(n21928), .ZN(n5121) );
  XNOR2_X1 U11280 ( .A(n21647), .B(n21106), .ZN(n21184) );
  XNOR2_X1 U11282 ( .A(n21184), .B(n5124), .ZN(n20978) );
  XNOR2_X1 U11283 ( .A(n21332), .B(n5125), .ZN(n5124) );
  NAND2_X1 U11284 ( .A1(n5127), .A2(n5129), .ZN(n5125) );
  OAI21_X1 U11285 ( .B1(n19260), .B2(n5131), .A(n5126), .ZN(n5128) );
  NAND3_X1 U11286 ( .A1(n276), .A2(n24463), .A3(n20975), .ZN(n5126) );
  INV_X1 U11287 ( .A(n5128), .ZN(n5127) );
  NAND2_X1 U11288 ( .A1(n5130), .A2(n19260), .ZN(n5129) );
  NAND2_X1 U11289 ( .A1(n19260), .A2(n5132), .ZN(n21583) );
  OAI21_X1 U11291 ( .B1(n19589), .B2(n5134), .A(n19588), .ZN(n19593) );
  NOR2_X1 U11292 ( .A1(n24422), .A2(n13323), .ZN(n13326) );
  OAI21_X1 U11293 ( .B1(n12062), .B2(n5140), .A(n5137), .ZN(n5141) );
  NOR2_X1 U11294 ( .A1(n3256), .A2(n13323), .ZN(n5138) );
  INV_X1 U11295 ( .A(n24422), .ZN(n5139) );
  NAND3_X1 U11296 ( .A1(n416), .A2(n10941), .A3(n3760), .ZN(n10379) );
  INV_X1 U11297 ( .A(n441), .ZN(n5144) );
  XNOR2_X1 U11298 ( .A(n21455), .B(n1891), .ZN(n21260) );
  OAI21_X2 U11300 ( .B1(n5148), .B2(n5146), .A(n5145), .ZN(n7628) );
  NAND2_X1 U11301 ( .A1(n5147), .A2(n7007), .ZN(n5146) );
  NAND2_X1 U11302 ( .A1(n6647), .A2(n7008), .ZN(n5147) );
  INV_X1 U11303 ( .A(n18428), .ZN(n5149) );
  NAND2_X1 U11304 ( .A1(n19164), .A2(n18788), .ZN(n18428) );
  XNOR2_X1 U11305 ( .A(n18388), .B(n17663), .ZN(n18413) );
  INV_X1 U11306 ( .A(n14327), .ZN(n5151) );
  NAND3_X1 U11307 ( .A1(n5151), .A2(n13864), .A3(n14044), .ZN(n5150) );
  AOI21_X1 U11308 ( .B1(n25072), .B2(n1443), .A(n5153), .ZN(n5152) );
  NOR2_X1 U11309 ( .A1(n280), .A2(n19578), .ZN(n5153) );
  NAND2_X1 U11310 ( .A1(n12931), .A2(n12897), .ZN(n5156) );
  XNOR2_X1 U11311 ( .A(n8297), .B(n8034), .ZN(n5157) );
  OAI21_X1 U11313 ( .B1(n19476), .B2(n18734), .A(n19478), .ZN(n17640) );
  XNOR2_X1 U11315 ( .A(n18372), .B(n17710), .ZN(n5160) );
  NAND2_X1 U11316 ( .A1(n311), .A2(n7604), .ZN(n7324) );
  NOR2_X2 U11318 ( .A1(n15678), .A2(n5164), .ZN(n17326) );
  NAND2_X1 U11319 ( .A1(n5166), .A2(n5165), .ZN(n5164) );
  NAND2_X1 U11320 ( .A1(n15675), .A2(n16328), .ZN(n5166) );
  INV_X1 U11321 ( .A(n16232), .ZN(n15933) );
  OAI21_X1 U11322 ( .B1(n5169), .B2(n15932), .A(n5168), .ZN(n5167) );
  AOI21_X1 U11323 ( .B1(n5405), .B2(n20134), .A(n5566), .ZN(n5404) );
  NAND3_X1 U11324 ( .A1(n12873), .A2(n12872), .A3(n13123), .ZN(n5170) );
  NAND2_X1 U11325 ( .A1(n12875), .A2(n5624), .ZN(n5172) );
  OAI21_X1 U11326 ( .B1(n13305), .B2(n12555), .A(n5173), .ZN(n5175) );
  NAND2_X1 U11327 ( .A1(n12555), .A2(n12611), .ZN(n5173) );
  NAND2_X1 U11328 ( .A1(n16115), .A2(n16120), .ZN(n5177) );
  XNOR2_X1 U11329 ( .A(n5179), .B(n8755), .ZN(n5255) );
  XNOR2_X1 U11330 ( .A(n5179), .B(n9052), .ZN(n9054) );
  XNOR2_X1 U11331 ( .A(n5179), .B(n8754), .ZN(n8559) );
  XNOR2_X1 U11332 ( .A(n5179), .B(n9190), .ZN(n8121) );
  MUX2_X1 U11334 ( .A(n20118), .B(n25514), .S(n19883), .Z(n19718) );
  INV_X1 U11335 ( .A(n11433), .ZN(n12376) );
  XNOR2_X1 U11336 ( .A(n5180), .B(n10689), .ZN(n11343) );
  XNOR2_X1 U11337 ( .A(n5181), .B(n10689), .ZN(n11658) );
  XNOR2_X1 U11338 ( .A(n10689), .B(n5182), .ZN(n12011) );
  XNOR2_X1 U11339 ( .A(n5183), .B(n8734), .ZN(n7310) );
  INV_X1 U11340 ( .A(n8329), .ZN(n5183) );
  XNOR2_X1 U11341 ( .A(n8734), .B(n5184), .ZN(n8357) );
  NAND2_X1 U11343 ( .A1(n20410), .A2(n20411), .ZN(n5187) );
  NAND2_X1 U11344 ( .A1(n20409), .A2(n20264), .ZN(n5188) );
  INV_X1 U11345 ( .A(n22452), .ZN(n5190) );
  NAND2_X1 U11346 ( .A1(n5191), .A2(n12626), .ZN(n12627) );
  MUX2_X1 U11347 ( .A(n16100), .B(n16101), .S(n15583), .Z(n16103) );
  NAND2_X1 U11348 ( .A1(n8005), .A2(n7292), .ZN(n7541) );
  XNOR2_X1 U11349 ( .A(n22006), .B(n2805), .ZN(n21752) );
  NAND2_X1 U11350 ( .A1(n20362), .A2(n24078), .ZN(n5193) );
  INV_X1 U11354 ( .A(n24909), .ZN(n5196) );
  OAI21_X1 U11355 ( .B1(n17764), .B2(n5196), .A(n17763), .ZN(n17765) );
  INV_X1 U11356 ( .A(n10505), .ZN(n5198) );
  NAND2_X1 U11357 ( .A1(n9809), .A2(n9338), .ZN(n5199) );
  INV_X1 U11358 ( .A(n5200), .ZN(n15374) );
  XNOR2_X1 U11359 ( .A(n5200), .B(n14454), .ZN(n14456) );
  OAI21_X1 U11360 ( .B1(n12816), .B2(n12815), .A(n12814), .ZN(n5200) );
  XNOR2_X1 U11361 ( .A(n15374), .B(n3232), .ZN(n14547) );
  NAND3_X1 U11362 ( .A1(n24908), .A2(n19389), .A3(n25052), .ZN(n19111) );
  OAI21_X1 U11363 ( .B1(n5202), .B2(n432), .A(n5201), .ZN(n5204) );
  NAND2_X1 U11364 ( .A1(n432), .A2(n7292), .ZN(n5201) );
  XNOR2_X1 U11365 ( .A(n21043), .B(n641), .ZN(n5339) );
  XNOR2_X1 U11366 ( .A(n5210), .B(n15477), .ZN(n5513) );
  XNOR2_X1 U11367 ( .A(n5210), .B(n14374), .ZN(n14375) );
  XNOR2_X1 U11368 ( .A(n5210), .B(n13691), .ZN(n13710) );
  NOR2_X1 U11369 ( .A1(n15646), .A2(n24061), .ZN(n5211) );
  OAI21_X1 U11370 ( .B1(n19326), .B2(n24516), .A(n19329), .ZN(n17945) );
  OAI211_X1 U11371 ( .C1(n19328), .C2(n18933), .A(n19326), .B(n24516), .ZN(
        n17498) );
  AOI21_X1 U11373 ( .B1(n19330), .B2(n24516), .A(n5213), .ZN(n19332) );
  NAND2_X1 U11374 ( .A1(n18938), .A2(n24583), .ZN(n18853) );
  INV_X1 U11377 ( .A(n13532), .ZN(n5216) );
  XNOR2_X1 U11378 ( .A(n5217), .B(n450), .ZN(Ciphertext[186]) );
  NAND2_X1 U11379 ( .A1(n5220), .A2(n5219), .ZN(n5218) );
  NAND2_X1 U11380 ( .A1(n23984), .A2(n24014), .ZN(n5219) );
  OAI21_X1 U11381 ( .B1(n24448), .B2(n23978), .A(n23993), .ZN(n5220) );
  NAND2_X1 U11382 ( .A1(n22322), .A2(n24496), .ZN(n5222) );
  NAND2_X1 U11383 ( .A1(n23228), .A2(n23227), .ZN(n23221) );
  INV_X1 U11384 ( .A(n21766), .ZN(n22064) );
  NAND2_X1 U11386 ( .A1(n15958), .A2(n5229), .ZN(n17434) );
  AND2_X1 U11387 ( .A1(n16170), .A2(n16426), .ZN(n5229) );
  NAND2_X1 U11388 ( .A1(n15958), .A2(n16170), .ZN(n16172) );
  NAND2_X1 U11389 ( .A1(n21917), .A2(n1352), .ZN(n5231) );
  NOR2_X1 U11390 ( .A1(n329), .A2(n22455), .ZN(n21917) );
  NAND2_X1 U11391 ( .A1(n9468), .A2(n9963), .ZN(n5232) );
  NAND2_X1 U11392 ( .A1(n19036), .A2(n19451), .ZN(n5234) );
  OAI211_X2 U11393 ( .C1(n17561), .C2(n5238), .A(n5237), .B(n17560), .ZN(
        n20316) );
  NAND3_X1 U11394 ( .A1(n4554), .A2(n5243), .A3(n5242), .ZN(n5241) );
  AOI21_X1 U11395 ( .B1(n16100), .B2(n16101), .A(n15583), .ZN(n15632) );
  NAND2_X1 U11396 ( .A1(n15780), .A2(n15583), .ZN(n16681) );
  NAND2_X1 U11397 ( .A1(n5458), .A2(n5245), .ZN(n5459) );
  INV_X1 U11398 ( .A(n10623), .ZN(n10669) );
  NAND2_X1 U11399 ( .A1(n5824), .A2(n6473), .ZN(n5249) );
  NAND2_X1 U11401 ( .A1(n13392), .A2(n13975), .ZN(n5252) );
  AOI21_X1 U11402 ( .B1(n13391), .B2(n13974), .A(n13390), .ZN(n5253) );
  OAI21_X2 U11403 ( .B1(n5254), .B2(n9316), .A(n9317), .ZN(n11128) );
  OAI21_X1 U11404 ( .B1(n422), .B2(n9989), .A(n25444), .ZN(n5254) );
  XNOR2_X1 U11405 ( .A(n5255), .B(n8672), .ZN(n8679) );
  NAND2_X1 U11406 ( .A1(n14320), .A2(n13868), .ZN(n5256) );
  NAND2_X1 U11408 ( .A1(n22591), .A2(n21921), .ZN(n5258) );
  OAI211_X2 U11409 ( .C1(n20311), .C2(n25101), .A(n5262), .B(n5261), .ZN(
        n21324) );
  NAND3_X1 U11410 ( .A1(n20309), .A2(n25101), .A3(n20549), .ZN(n5261) );
  NAND2_X1 U11412 ( .A1(n20309), .A2(n20549), .ZN(n20544) );
  INV_X1 U11413 ( .A(n7175), .ZN(n5264) );
  NAND2_X1 U11414 ( .A1(n7418), .A2(n7789), .ZN(n7175) );
  NAND2_X1 U11415 ( .A1(n5264), .A2(n7782), .ZN(n5263) );
  NAND3_X1 U11416 ( .A1(n5267), .A2(n5266), .A3(n7783), .ZN(n5265) );
  NAND2_X1 U11417 ( .A1(n7784), .A2(n7787), .ZN(n5267) );
  NAND2_X1 U11418 ( .A1(n7420), .A2(n7419), .ZN(n5268) );
  AOI21_X1 U11419 ( .B1(n6468), .B2(n6469), .A(n6467), .ZN(n5270) );
  NAND3_X1 U11420 ( .A1(n7638), .A2(n312), .A3(n7915), .ZN(n7396) );
  NAND2_X1 U11421 ( .A1(n9670), .A2(n9669), .ZN(n5273) );
  NOR2_X1 U11422 ( .A1(n9730), .A2(n9729), .ZN(n5275) );
  NAND2_X1 U11423 ( .A1(n10020), .A2(n5275), .ZN(n5274) );
  NAND2_X1 U11424 ( .A1(n9650), .A2(n9730), .ZN(n5276) );
  NAND2_X1 U11425 ( .A1(n9730), .A2(n25475), .ZN(n5278) );
  NOR2_X1 U11426 ( .A1(n5280), .A2(n20388), .ZN(n20387) );
  NOR2_X1 U11427 ( .A1(n5280), .A2(n19490), .ZN(n19349) );
  NAND3_X1 U11428 ( .A1(n25473), .A2(n19490), .A3(n5280), .ZN(n19492) );
  OAI21_X1 U11429 ( .B1(n23728), .B2(n24381), .A(n5286), .ZN(n5283) );
  NAND3_X1 U11430 ( .A1(n22091), .A2(n5282), .A3(n5281), .ZN(n5285) );
  NAND3_X1 U11431 ( .A1(n5284), .A2(n24374), .A3(n23714), .ZN(n5281) );
  INV_X1 U11432 ( .A(n5283), .ZN(n5282) );
  OR2_X1 U11434 ( .A1(n22091), .A2(Key[60]), .ZN(n5287) );
  NAND2_X1 U11435 ( .A1(n5289), .A2(n9372), .ZN(n5288) );
  NAND2_X1 U11436 ( .A1(n19302), .A2(n19128), .ZN(n5290) );
  NAND2_X1 U11438 ( .A1(n7053), .A2(n7803), .ZN(n5291) );
  OAI211_X2 U11439 ( .C1(n7434), .C2(n7054), .A(n5294), .B(n5292), .ZN(n8896)
         );
  OR2_X1 U11440 ( .A1(n5293), .A2(n7795), .ZN(n5292) );
  NAND2_X1 U11441 ( .A1(n7798), .A2(n7166), .ZN(n5293) );
  NAND2_X1 U11442 ( .A1(n7166), .A2(n6280), .ZN(n7053) );
  NAND2_X1 U11443 ( .A1(n17173), .A2(n16434), .ZN(n16432) );
  NAND2_X1 U11444 ( .A1(n13478), .A2(n5299), .ZN(n5298) );
  XNOR2_X1 U11445 ( .A(n5300), .B(n16037), .ZN(n5302) );
  XNOR2_X1 U11446 ( .A(n18374), .B(n18513), .ZN(n5304) );
  NAND2_X1 U11447 ( .A1(n16970), .A2(n16969), .ZN(n5305) );
  NOR2_X1 U11448 ( .A1(n22506), .A2(n22528), .ZN(n5306) );
  NAND2_X1 U11449 ( .A1(n3240), .A2(n19849), .ZN(n19855) );
  INV_X1 U11450 ( .A(n12683), .ZN(n5311) );
  NOR2_X1 U11452 ( .A1(n2561), .A2(n5316), .ZN(n5315) );
  NAND2_X1 U11453 ( .A1(n5318), .A2(n7761), .ZN(n5689) );
  INV_X1 U11454 ( .A(n13094), .ZN(n12649) );
  XNOR2_X2 U11455 ( .A(n9680), .B(n9679), .ZN(n13094) );
  NAND2_X1 U11456 ( .A1(n5319), .A2(n5325), .ZN(n13675) );
  NAND2_X1 U11457 ( .A1(n5320), .A2(n5323), .ZN(n5319) );
  NAND2_X1 U11458 ( .A1(n5322), .A2(n5321), .ZN(n5320) );
  NAND2_X1 U11459 ( .A1(n12649), .A2(n12648), .ZN(n5322) );
  INV_X1 U11460 ( .A(n12648), .ZN(n5324) );
  NOR2_X2 U11461 ( .A1(n13791), .A2(n5330), .ZN(n15484) );
  XNOR2_X1 U11463 ( .A(n14898), .B(n1411), .ZN(n5331) );
  NAND2_X1 U11464 ( .A1(n5333), .A2(n5709), .ZN(n5332) );
  AND2_X1 U11465 ( .A1(n13565), .A2(n14108), .ZN(n5709) );
  NAND2_X1 U11466 ( .A1(n19061), .A2(n24982), .ZN(n5337) );
  NAND2_X1 U11467 ( .A1(n9390), .A2(n9389), .ZN(n5341) );
  NAND2_X1 U11468 ( .A1(n25203), .A2(n11069), .ZN(n5342) );
  XNOR2_X1 U11469 ( .A(n5344), .B(n7161), .ZN(n8430) );
  XNOR2_X1 U11470 ( .A(n5346), .B(n7161), .ZN(n8149) );
  INV_X1 U11471 ( .A(n22493), .ZN(n5347) );
  NAND3_X1 U11472 ( .A1(n5349), .A2(n22528), .A3(n23443), .ZN(n5348) );
  NAND2_X1 U11473 ( .A1(n22491), .A2(n22733), .ZN(n5350) );
  NAND2_X1 U11474 ( .A1(n23442), .A2(n25042), .ZN(n22527) );
  INV_X1 U11475 ( .A(n10871), .ZN(n5352) );
  OAI21_X1 U11476 ( .B1(n11115), .B2(n11117), .A(n5351), .ZN(n10878) );
  NAND2_X1 U11477 ( .A1(n5357), .A2(n10120), .ZN(n5356) );
  NAND2_X1 U11478 ( .A1(n24096), .A2(n5359), .ZN(n11837) );
  NAND3_X1 U11479 ( .A1(n23810), .A2(n25391), .A3(n23811), .ZN(n22540) );
  NAND2_X1 U11480 ( .A1(n10114), .A2(n9338), .ZN(n5362) );
  NOR2_X1 U11482 ( .A1(n20600), .A2(n5364), .ZN(n5363) );
  NOR2_X1 U11483 ( .A1(n276), .A2(n5365), .ZN(n5364) );
  NAND2_X1 U11484 ( .A1(n266), .A2(n17356), .ZN(n5367) );
  INV_X1 U11485 ( .A(n12533), .ZN(n5368) );
  XNOR2_X1 U11486 ( .A(n24337), .B(n18499), .ZN(n18225) );
  XNOR2_X1 U11487 ( .A(n17850), .B(n18289), .ZN(n5369) );
  OAI211_X1 U11488 ( .C1(n19322), .C2(n19472), .A(n19467), .B(n18959), .ZN(
        n19323) );
  NAND2_X1 U11489 ( .A1(n18959), .A2(n17872), .ZN(n18962) );
  OAI21_X1 U11490 ( .B1(n19467), .B2(n18959), .A(n19466), .ZN(n19468) );
  AND2_X1 U11492 ( .A1(n19314), .A2(n5370), .ZN(n19320) );
  NAND3_X1 U11493 ( .A1(n19309), .A2(n24912), .A3(n5371), .ZN(n5370) );
  NAND2_X1 U11494 ( .A1(n5372), .A2(n9493), .ZN(n10776) );
  NAND2_X1 U11496 ( .A1(n5372), .A2(n9732), .ZN(n9733) );
  INV_X1 U11497 ( .A(n18397), .ZN(n18284) );
  XNOR2_X1 U11498 ( .A(n18397), .B(n5374), .ZN(n5373) );
  INV_X1 U11499 ( .A(n16551), .ZN(n5375) );
  AOI22_X1 U11500 ( .A1(n16554), .A2(n16553), .B1(n16552), .B2(n5376), .ZN(
        n17680) );
  INV_X1 U11501 ( .A(n5378), .ZN(n22370) );
  NAND2_X1 U11502 ( .A1(n5378), .A2(n22769), .ZN(n21292) );
  NAND2_X1 U11503 ( .A1(n22680), .A2(n5378), .ZN(n20605) );
  AOI21_X1 U11504 ( .B1(n5378), .B2(n22770), .A(n22769), .ZN(n22775) );
  AOI21_X1 U11505 ( .B1(n22773), .B2(n22772), .A(n5378), .ZN(n5611) );
  NAND3_X1 U11507 ( .A1(n1552), .A2(n415), .A3(n11101), .ZN(n5379) );
  OAI21_X1 U11508 ( .B1(n11101), .B2(n5380), .A(n10912), .ZN(n5381) );
  NAND2_X1 U11509 ( .A1(n1552), .A2(n10772), .ZN(n5380) );
  NAND3_X1 U11511 ( .A1(n15773), .A2(n16024), .A3(n5383), .ZN(n15776) );
  NAND2_X1 U11512 ( .A1(n5385), .A2(n16923), .ZN(n5384) );
  NOR2_X1 U11513 ( .A1(n17320), .A2(n16927), .ZN(n5385) );
  AND2_X1 U11514 ( .A1(n16809), .A2(n17077), .ZN(n5386) );
  AND2_X1 U11515 ( .A1(n7364), .A2(n7909), .ZN(n5387) );
  NAND2_X1 U11517 ( .A1(n7365), .A2(n7908), .ZN(n5389) );
  NAND2_X1 U11519 ( .A1(n10574), .A2(n11039), .ZN(n5393) );
  AOI21_X1 U11520 ( .B1(n25071), .B2(n24893), .A(n323), .ZN(n5396) );
  AOI22_X1 U11521 ( .A1(n22710), .A2(n323), .B1(n5397), .B2(n5396), .ZN(n5398)
         );
  XNOR2_X1 U11522 ( .A(n5398), .B(n3798), .ZN(Ciphertext[110]) );
  XNOR2_X1 U11523 ( .A(n5399), .B(n21079), .ZN(Ciphertext[125]) );
  OAI211_X1 U11524 ( .C1(n21078), .C2(n23650), .A(n5401), .B(n5400), .ZN(n5399) );
  NAND3_X1 U11525 ( .A1(n23637), .A2(n23640), .A3(n23629), .ZN(n5400) );
  NAND2_X1 U11526 ( .A1(n23651), .A2(n23649), .ZN(n5401) );
  NAND2_X1 U11530 ( .A1(n15259), .A2(n25323), .ZN(n5407) );
  NAND2_X1 U11531 ( .A1(n16191), .A2(n16197), .ZN(n15901) );
  INV_X1 U11532 ( .A(n17424), .ZN(n5409) );
  OAI21_X1 U11533 ( .B1(n12861), .B2(n12636), .A(n5410), .ZN(n12638) );
  NAND2_X1 U11534 ( .A1(n12636), .A2(n13345), .ZN(n5410) );
  NAND2_X1 U11535 ( .A1(n5731), .A2(n5412), .ZN(n5411) );
  OR2_X1 U11536 ( .A1(n7583), .A2(n7584), .ZN(n5490) );
  NAND3_X1 U11537 ( .A1(n7475), .A2(n7952), .A3(n5413), .ZN(n7424) );
  OAI21_X1 U11538 ( .B1(n23206), .B2(n22820), .A(n5769), .ZN(n5415) );
  NOR2_X1 U11539 ( .A1(n13988), .A2(n13987), .ZN(n13917) );
  NAND2_X1 U11540 ( .A1(n13242), .A2(n5417), .ZN(n5416) );
  INV_X1 U11541 ( .A(n13248), .ZN(n5417) );
  INV_X1 U11542 ( .A(n13211), .ZN(n5418) );
  OAI211_X1 U11543 ( .C1(n25004), .C2(n24341), .A(n5420), .B(n25081), .ZN(
        n5419) );
  NAND2_X1 U11544 ( .A1(n5421), .A2(n24342), .ZN(n5420) );
  INV_X1 U11545 ( .A(n22932), .ZN(n5421) );
  NAND2_X1 U11546 ( .A1(n22931), .A2(n22499), .ZN(n5422) );
  NAND2_X1 U11547 ( .A1(n343), .A2(n20499), .ZN(n5423) );
  NAND2_X1 U11548 ( .A1(n16572), .A2(n5429), .ZN(n5428) );
  NAND2_X1 U11550 ( .A1(n16303), .A2(n24506), .ZN(n16305) );
  XNOR2_X1 U11552 ( .A(n24568), .B(n5433), .ZN(n16784) );
  INV_X1 U11553 ( .A(n17065), .ZN(n5434) );
  NAND2_X1 U11554 ( .A1(n5436), .A2(n13347), .ZN(n12973) );
  NAND2_X1 U11555 ( .A1(n1328), .A2(n5437), .ZN(n23586) );
  NAND3_X1 U11556 ( .A1(n1328), .A2(n23592), .A3(n22633), .ZN(n21777) );
  AND2_X1 U11558 ( .A1(n19255), .A2(n19596), .ZN(n5439) );
  INV_X1 U11559 ( .A(n14317), .ZN(n5440) );
  NOR2_X1 U11560 ( .A1(n13601), .A2(n13600), .ZN(n13604) );
  NAND2_X1 U11561 ( .A1(n18724), .A2(n19367), .ZN(n19222) );
  NOR2_X1 U11562 ( .A1(n24366), .A2(n5447), .ZN(n5446) );
  INV_X1 U11563 ( .A(n16268), .ZN(n5447) );
  INV_X1 U11564 ( .A(n9296), .ZN(n5448) );
  XNOR2_X1 U11566 ( .A(n12073), .B(n12005), .ZN(n10421) );
  NAND3_X1 U11570 ( .A1(n5454), .A2(n25474), .A3(n240), .ZN(n5456) );
  XNOR2_X1 U11572 ( .A(n5457), .B(n21139), .ZN(n21140) );
  XNOR2_X1 U11573 ( .A(n1461), .B(n21664), .ZN(n5457) );
  XNOR2_X1 U11574 ( .A(n24305), .B(n21138), .ZN(n21664) );
  NAND3_X1 U11576 ( .A1(n5460), .A2(n7924), .A3(n7923), .ZN(n7373) );
  NAND2_X1 U11577 ( .A1(n5461), .A2(n24424), .ZN(n19100) );
  AND2_X1 U11578 ( .A1(n25382), .A2(n22901), .ZN(n22482) );
  NOR2_X1 U11579 ( .A1(n5463), .A2(n22907), .ZN(n22908) );
  NAND2_X1 U11580 ( .A1(n22921), .A2(n5465), .ZN(n23008) );
  AOI21_X1 U11582 ( .B1(n19121), .B2(n20054), .A(n25089), .ZN(n5467) );
  OAI22_X1 U11583 ( .A1(n5469), .A2(n13628), .B1(n14079), .B2(n14083), .ZN(
        n12705) );
  MUX2_X1 U11584 ( .A(n14077), .B(n13852), .S(n14075), .Z(n5469) );
  NAND2_X1 U11585 ( .A1(n5476), .A2(n5474), .ZN(n20259) );
  NAND2_X1 U11586 ( .A1(n5477), .A2(n19531), .ZN(n5476) );
  NAND2_X1 U11588 ( .A1(n19530), .A2(n19145), .ZN(n5478) );
  OR2_X1 U11590 ( .A1(n19531), .A2(n19534), .ZN(n5481) );
  NAND2_X1 U11591 ( .A1(n5487), .A2(n5484), .ZN(n5482) );
  NAND2_X1 U11592 ( .A1(n14397), .A2(n5484), .ZN(n5483) );
  NAND2_X1 U11594 ( .A1(n5486), .A2(n2215), .ZN(n5485) );
  INV_X1 U11595 ( .A(n14397), .ZN(n5486) );
  OAI22_X1 U11596 ( .A1(n10178), .A2(n9832), .B1(n10175), .B2(n10177), .ZN(
        n9385) );
  NAND2_X1 U11597 ( .A1(n6600), .A2(n7019), .ZN(n5488) );
  XNOR2_X1 U11598 ( .A(n21208), .B(n21209), .ZN(n21210) );
  OAI21_X1 U11602 ( .B1(n19521), .B2(n19523), .A(n5496), .ZN(n18894) );
  XNOR2_X2 U11603 ( .A(n18194), .B(n18193), .ZN(n19523) );
  INV_X1 U11605 ( .A(n13924), .ZN(n5497) );
  NOR2_X1 U11606 ( .A1(n14250), .A2(n13924), .ZN(n5498) );
  MUX2_X1 U11607 ( .A(n14008), .B(n14254), .S(n13924), .Z(n14012) );
  NAND3_X1 U11608 ( .A1(n15655), .A2(n16381), .A3(n15656), .ZN(n5502) );
  NOR2_X1 U11609 ( .A1(n20054), .A2(n20055), .ZN(n20471) );
  OAI21_X1 U11610 ( .B1(n13336), .B2(n12958), .A(n5505), .ZN(n13342) );
  AND2_X1 U11611 ( .A1(n23670), .A2(n5506), .ZN(n23668) );
  OR3_X1 U11612 ( .A1(n23667), .A2(n5508), .A3(n23679), .ZN(n5507) );
  NOR2_X1 U11613 ( .A1(n22157), .A2(n25018), .ZN(n5508) );
  INV_X1 U11614 ( .A(n7798), .ZN(n7167) );
  NAND3_X1 U11615 ( .A1(n7432), .A2(n7167), .A3(n7166), .ZN(n7168) );
  OAI211_X1 U11616 ( .C1(n17214), .C2(n17216), .A(n17212), .B(n5510), .ZN(
        n5509) );
  AOI21_X1 U11618 ( .B1(n12694), .B2(n13289), .A(n12824), .ZN(n11804) );
  NAND2_X1 U11619 ( .A1(n5533), .A2(n10060), .ZN(n5519) );
  INV_X1 U11620 ( .A(n10060), .ZN(n5518) );
  OAI21_X2 U11621 ( .B1(n13727), .B2(n5520), .A(n13726), .ZN(n15074) );
  NAND2_X1 U11622 ( .A1(n16766), .A2(n5522), .ZN(n5521) );
  NAND3_X1 U11623 ( .A1(n9897), .A2(n24083), .A3(n5524), .ZN(n8138) );
  OR2_X1 U11624 ( .A1(n9944), .A2(n9899), .ZN(n5523) );
  NAND2_X1 U11625 ( .A1(n9896), .A2(n5524), .ZN(n9902) );
  INV_X1 U11626 ( .A(n9899), .ZN(n5524) );
  NAND2_X1 U11627 ( .A1(n24995), .A2(n13569), .ZN(n5525) );
  NAND2_X1 U11628 ( .A1(n6255), .A2(n5903), .ZN(n6953) );
  NOR2_X1 U11629 ( .A1(n25550), .A2(n23275), .ZN(n5531) );
  NAND2_X1 U11630 ( .A1(n5531), .A2(n24907), .ZN(n5530) );
  NAND2_X1 U11632 ( .A1(n309), .A2(n9218), .ZN(n5533) );
  OAI21_X1 U11633 ( .B1(n10062), .B2(n5533), .A(n9220), .ZN(n9128) );
  MUX2_X1 U11634 ( .A(n5533), .B(n9414), .S(n10060), .Z(n9415) );
  NAND2_X1 U11635 ( .A1(n9519), .A2(n5536), .ZN(n5535) );
  NAND2_X1 U11636 ( .A1(n5537), .A2(n10176), .ZN(n5536) );
  NAND2_X1 U11637 ( .A1(n10186), .A2(n10179), .ZN(n5537) );
  AOI21_X1 U11638 ( .B1(n13210), .B2(n13212), .A(n13213), .ZN(n5538) );
  NAND2_X1 U11639 ( .A1(n23165), .A2(n23181), .ZN(n22552) );
  NAND2_X1 U11640 ( .A1(n22336), .A2(n24415), .ZN(n5539) );
  NAND2_X1 U11642 ( .A1(n20156), .A2(n24558), .ZN(n5541) );
  OAI21_X1 U11643 ( .B1(n12433), .B2(n13140), .A(n5542), .ZN(n5545) );
  NAND2_X1 U11644 ( .A1(n11109), .A2(n12455), .ZN(n5542) );
  INV_X1 U11645 ( .A(n12455), .ZN(n12729) );
  INV_X1 U11646 ( .A(n11109), .ZN(n13139) );
  NAND2_X1 U11647 ( .A1(n5545), .A2(n13143), .ZN(n5544) );
  NAND2_X1 U11648 ( .A1(n15720), .A2(n5546), .ZN(n15721) );
  XNOR2_X1 U11649 ( .A(n8506), .B(n9011), .ZN(n8250) );
  NAND2_X1 U11650 ( .A1(n5550), .A2(n7591), .ZN(n5547) );
  NOR2_X1 U11651 ( .A1(n5549), .A2(n5972), .ZN(n5548) );
  NAND2_X1 U11652 ( .A1(n5552), .A2(n5551), .ZN(n5550) );
  NAND2_X1 U11653 ( .A1(n5971), .A2(n7592), .ZN(n5551) );
  XNOR2_X1 U11654 ( .A(n5553), .B(n8739), .ZN(n8489) );
  XNOR2_X1 U11655 ( .A(n5554), .B(n8739), .ZN(n9062) );
  INV_X1 U11656 ( .A(n9146), .ZN(n5554) );
  XNOR2_X1 U11657 ( .A(n18326), .B(n18214), .ZN(n18576) );
  NAND2_X1 U11659 ( .A1(n16513), .A2(n16708), .ZN(n5557) );
  XNOR2_X1 U11660 ( .A(n12214), .B(n12324), .ZN(n11088) );
  NAND2_X1 U11661 ( .A1(n11083), .A2(n5559), .ZN(n5558) );
  OAI21_X1 U11662 ( .B1(n6949), .B2(n25437), .A(n24994), .ZN(n5560) );
  NAND2_X1 U11663 ( .A1(n5561), .A2(n12535), .ZN(n13757) );
  NAND2_X1 U11664 ( .A1(n20507), .A2(n25224), .ZN(n20511) );
  OAI211_X1 U11666 ( .C1(n3554), .C2(n15557), .A(n16312), .B(n15556), .ZN(
        n16641) );
  NAND2_X1 U11667 ( .A1(n20017), .A2(n25242), .ZN(n5564) );
  NAND2_X1 U11668 ( .A1(n5570), .A2(n5568), .ZN(n20256) );
  INV_X1 U11669 ( .A(n6721), .ZN(n5576) );
  NAND2_X1 U11670 ( .A1(n6727), .A2(n6723), .ZN(n5575) );
  NAND2_X1 U11671 ( .A1(n5575), .A2(n5576), .ZN(n5574) );
  INV_X1 U11673 ( .A(n12233), .ZN(n5577) );
  INV_X1 U11674 ( .A(n12089), .ZN(n5578) );
  XNOR2_X1 U11675 ( .A(n11907), .B(n5577), .ZN(n12236) );
  XNOR2_X1 U11676 ( .A(n5578), .B(n11907), .ZN(n12091) );
  XNOR2_X1 U11677 ( .A(n11907), .B(n24514), .ZN(n11911) );
  OAI211_X1 U11679 ( .C1(n15958), .C2(n707), .A(n5579), .B(n15825), .ZN(n5581)
         );
  NAND2_X1 U11680 ( .A1(n16424), .A2(n707), .ZN(n5579) );
  NAND2_X1 U11681 ( .A1(n15958), .A2(n1329), .ZN(n15962) );
  NAND2_X1 U11683 ( .A1(n5585), .A2(n22456), .ZN(n5582) );
  INV_X1 U11684 ( .A(n22451), .ZN(n5585) );
  NAND2_X1 U11686 ( .A1(n18908), .A2(n19565), .ZN(n5586) );
  NAND2_X1 U11687 ( .A1(n5589), .A2(n13350), .ZN(n5588) );
  NAND2_X1 U11688 ( .A1(n12349), .A2(n13124), .ZN(n5589) );
  NOR2_X1 U11689 ( .A1(n5591), .A2(n20401), .ZN(n20402) );
  NAND2_X1 U11690 ( .A1(n20419), .A2(n5591), .ZN(n19291) );
  AOI21_X1 U11691 ( .B1(n20419), .B2(n20415), .A(n25108), .ZN(n19860) );
  NAND2_X1 U11694 ( .A1(n4463), .A2(n10838), .ZN(n11135) );
  XNOR2_X1 U11695 ( .A(n17817), .B(n8347), .ZN(n18575) );
  XNOR2_X1 U11696 ( .A(n17817), .B(n5598), .ZN(n18701) );
  XNOR2_X1 U11697 ( .A(n8428), .B(n8690), .ZN(n9124) );
  NAND3_X1 U11698 ( .A1(n7736), .A2(n7734), .A3(n7735), .ZN(n5600) );
  NAND3_X1 U11699 ( .A1(n25151), .A2(n7736), .A3(n7731), .ZN(n5601) );
  NAND2_X1 U11700 ( .A1(n7730), .A2(n7733), .ZN(n5602) );
  NAND2_X1 U11701 ( .A1(n7165), .A2(n5603), .ZN(n8428) );
  INV_X1 U11702 ( .A(n7642), .ZN(n7736) );
  NOR2_X1 U11703 ( .A1(n7924), .A2(n7923), .ZN(n5605) );
  INV_X1 U11704 ( .A(n7932), .ZN(n7372) );
  NAND2_X1 U11705 ( .A1(n5613), .A2(n5612), .ZN(n20374) );
  NAND2_X1 U11706 ( .A1(n19545), .A2(n279), .ZN(n5612) );
  NAND2_X1 U11707 ( .A1(n19544), .A2(n19543), .ZN(n5613) );
  XNOR2_X1 U11708 ( .A(n5614), .B(n21662), .ZN(n8599) );
  XNOR2_X1 U11709 ( .A(n8313), .B(n5614), .ZN(n7379) );
  XNOR2_X1 U11710 ( .A(n8517), .B(n5614), .ZN(n8519) );
  XNOR2_X1 U11711 ( .A(n8223), .B(n5614), .ZN(n8793) );
  XNOR2_X1 U11712 ( .A(n9008), .B(n5614), .ZN(n9009) );
  NAND3_X1 U11713 ( .A1(n14315), .A2(n13460), .A3(n14311), .ZN(n14312) );
  NAND2_X1 U11714 ( .A1(n13901), .A2(n13460), .ZN(n13458) );
  NAND2_X1 U11715 ( .A1(n13904), .A2(n5615), .ZN(n15103) );
  OR2_X1 U11716 ( .A1(n13905), .A2(n13460), .ZN(n5615) );
  NAND2_X1 U11717 ( .A1(n25021), .A2(n9945), .ZN(n5616) );
  INV_X1 U11718 ( .A(n9893), .ZN(n9946) );
  NAND3_X1 U11720 ( .A1(n1429), .A2(n5618), .A3(n19169), .ZN(n5617) );
  INV_X1 U11721 ( .A(n19408), .ZN(n19171) );
  NAND2_X1 U11722 ( .A1(n19412), .A2(n19408), .ZN(n5618) );
  XNOR2_X1 U11723 ( .A(n9092), .B(n1414), .ZN(n5619) );
  OR2_X1 U11724 ( .A1(n10063), .A2(n10064), .ZN(n9702) );
  MUX2_X1 U11725 ( .A(n14059), .B(n14278), .S(n14850), .Z(n5620) );
  XNOR2_X1 U11726 ( .A(n18659), .B(n18334), .ZN(n17092) );
  NAND2_X1 U11727 ( .A1(n7365), .A2(n7629), .ZN(n5623) );
  OAI22_X1 U11728 ( .A1(n406), .A2(n13125), .B1(n13126), .B2(n5626), .ZN(
        n13127) );
  OAI21_X1 U11729 ( .B1(n10623), .B2(n10810), .A(n3868), .ZN(n5630) );
  INV_X1 U11731 ( .A(n19273), .ZN(n5633) );
  NAND2_X1 U11732 ( .A1(n19570), .A2(n5634), .ZN(n19567) );
  OAI21_X1 U11733 ( .B1(n1053), .B2(n19191), .A(n5631), .ZN(n18909) );
  NAND2_X1 U11734 ( .A1(n5633), .A2(n19192), .ZN(n5631) );
  NAND3_X1 U11736 ( .A1(n20545), .A2(n20546), .A3(n20124), .ZN(n5637) );
  XNOR2_X1 U11738 ( .A(n14858), .B(n15056), .ZN(n15427) );
  NAND2_X1 U11739 ( .A1(n14140), .A2(n5641), .ZN(n5640) );
  NAND3_X1 U11740 ( .A1(n14142), .A2(n14141), .A3(n5641), .ZN(n5642) );
  NAND2_X1 U11741 ( .A1(n12933), .A2(n12934), .ZN(n5643) );
  NOR2_X1 U11742 ( .A1(n20480), .A2(n20476), .ZN(n19628) );
  OAI211_X1 U11743 ( .C1(n19413), .C2(n19173), .A(n5647), .B(n19170), .ZN(
        n5646) );
  NAND2_X1 U11744 ( .A1(n19173), .A2(n19171), .ZN(n5647) );
  OAI211_X1 U11745 ( .C1(n6909), .C2(n6918), .A(n6774), .B(n24037), .ZN(n5649)
         );
  OR2_X1 U11746 ( .A1(n6773), .A2(n6770), .ZN(n5651) );
  NAND2_X1 U11747 ( .A1(n5650), .A2(n5649), .ZN(n7974) );
  NOR2_X1 U11748 ( .A1(n24393), .A2(n19531), .ZN(n5655) );
  NAND4_X2 U11749 ( .A1(n19271), .A2(n5652), .A3(n5654), .A4(n5653), .ZN(
        n20400) );
  NAND2_X1 U11750 ( .A1(n5655), .A2(n19269), .ZN(n5653) );
  AND2_X1 U11751 ( .A1(n5924), .A2(n6956), .ZN(n5656) );
  NAND2_X1 U11752 ( .A1(n5658), .A2(n23326), .ZN(n23328) );
  NAND2_X1 U11753 ( .A1(n5660), .A2(n5659), .ZN(n5658) );
  NAND2_X1 U11755 ( .A1(n21956), .A2(n5663), .ZN(n5662) );
  INV_X1 U11756 ( .A(n22128), .ZN(n5663) );
  NAND2_X1 U11758 ( .A1(n338), .A2(n21467), .ZN(n5665) );
  NAND3_X1 U11759 ( .A1(n407), .A2(n25015), .A3(n12680), .ZN(n12608) );
  MUX2_X1 U11760 ( .A(n13266), .B(n13264), .S(n12680), .Z(n13271) );
  NAND2_X1 U11761 ( .A1(n19414), .A2(n19413), .ZN(n5669) );
  NAND3_X1 U11762 ( .A1(n5673), .A2(n13283), .A3(n12899), .ZN(n12700) );
  NAND2_X1 U11763 ( .A1(n25191), .A2(n12897), .ZN(n5673) );
  NAND3_X2 U11764 ( .A1(n16735), .A2(n5675), .A3(n5674), .ZN(n18190) );
  NAND2_X1 U11765 ( .A1(n5676), .A2(n16730), .ZN(n5675) );
  NOR2_X1 U11766 ( .A1(n16731), .A2(n369), .ZN(n5676) );
  MUX2_X1 U11767 ( .A(n23278), .B(n23281), .S(n24349), .Z(n22537) );
  INV_X1 U11768 ( .A(n11025), .ZN(n5679) );
  XNOR2_X1 U11769 ( .A(n11310), .B(n12234), .ZN(n11851) );
  NAND2_X1 U11770 ( .A1(n19225), .A2(n5680), .ZN(n19226) );
  NAND2_X1 U11771 ( .A1(n20193), .A2(n20576), .ZN(n5680) );
  NAND2_X1 U11772 ( .A1(n5682), .A2(n25243), .ZN(n5681) );
  NAND2_X1 U11773 ( .A1(n5683), .A2(n7962), .ZN(n7963) );
  NAND2_X1 U11774 ( .A1(n5684), .A2(n7961), .ZN(n5683) );
  NAND2_X1 U11775 ( .A1(n18848), .A2(n19477), .ZN(n5686) );
  NAND3_X1 U11776 ( .A1(n18848), .A2(n19482), .A3(n19477), .ZN(n18973) );
  INV_X1 U11777 ( .A(n9231), .ZN(n9763) );
  OAI21_X1 U11778 ( .B1(n10070), .B2(n9231), .A(n5688), .ZN(n9622) );
  NAND2_X1 U11780 ( .A1(n9622), .A2(n1330), .ZN(n9413) );
  XNOR2_X1 U11781 ( .A(n8616), .B(n5690), .ZN(n8102) );
  NAND2_X1 U11782 ( .A1(n15937), .A2(n387), .ZN(n15934) );
  OAI21_X1 U11785 ( .B1(n5697), .B2(n6323), .A(n5696), .ZN(n5695) );
  NOR2_X1 U11787 ( .A1(n25398), .A2(n943), .ZN(n5697) );
  AOI21_X1 U11788 ( .B1(n5700), .B2(n5699), .A(n23528), .ZN(n23534) );
  NAND3_X1 U11789 ( .A1(n23533), .A2(n23531), .A3(n23532), .ZN(n5699) );
  NAND2_X1 U11790 ( .A1(n5701), .A2(n5702), .ZN(n5700) );
  NAND2_X1 U11791 ( .A1(n23505), .A2(n24351), .ZN(n5702) );
  INV_X1 U11794 ( .A(n11761), .ZN(n11913) );
  NOR2_X1 U11796 ( .A1(n13373), .A2(n15888), .ZN(n5706) );
  NAND2_X1 U11797 ( .A1(n17413), .A2(n17225), .ZN(n5707) );
  INV_X1 U11798 ( .A(n14108), .ZN(n13582) );
  INV_X1 U11799 ( .A(n20471), .ZN(n5710) );
  NAND2_X1 U11800 ( .A1(n25088), .A2(n20060), .ZN(n20468) );
  INV_X1 U11801 ( .A(n22770), .ZN(n5712) );
  MUX2_X1 U11802 ( .A(n22370), .B(n22774), .S(n21856), .Z(n22371) );
  OR2_X1 U11803 ( .A1(n7434), .A2(n7800), .ZN(n5713) );
  OAI21_X1 U11804 ( .B1(n7799), .B2(n7794), .A(n5715), .ZN(n5714) );
  NAND2_X1 U11805 ( .A1(n7794), .A2(n7802), .ZN(n5715) );
  INV_X1 U11806 ( .A(n16100), .ZN(n16085) );
  INV_X1 U11807 ( .A(n15584), .ZN(n5716) );
  NAND2_X1 U11808 ( .A1(n5716), .A2(n16101), .ZN(n15582) );
  NAND2_X1 U11809 ( .A1(n16957), .A2(n17414), .ZN(n16954) );
  NAND2_X1 U11812 ( .A1(n6638), .A2(n6848), .ZN(n5719) );
  NAND2_X1 U11813 ( .A1(n6109), .A2(n250), .ZN(n5720) );
  XNOR2_X1 U11816 ( .A(n5722), .B(n18509), .ZN(n18165) );
  INV_X1 U11817 ( .A(n18218), .ZN(n5722) );
  AOI21_X1 U11818 ( .B1(n18782), .B2(n18783), .A(n19411), .ZN(n18787) );
  NAND3_X1 U11819 ( .A1(n12759), .A2(n13030), .A3(n13024), .ZN(n5723) );
  NAND2_X1 U11820 ( .A1(n12760), .A2(n13028), .ZN(n5724) );
  NAND2_X1 U11823 ( .A1(n10190), .A2(n25230), .ZN(n10857) );
  NAND2_X1 U11824 ( .A1(n10190), .A2(n5727), .ZN(n10865) );
  AND3_X1 U11825 ( .A1(n22587), .A2(n22804), .A3(n22586), .ZN(n22588) );
  OR2_X1 U11827 ( .A1(n19313), .A2(n19312), .ZN(n18842) );
  OR2_X1 U11829 ( .A1(n20450), .A2(n20377), .ZN(n19772) );
  OR2_X1 U11830 ( .A1(n20401), .A2(n20414), .ZN(n20203) );
  AND2_X1 U11831 ( .A1(n20414), .A2(n20401), .ZN(n19857) );
  XNOR2_X1 U11832 ( .A(n16960), .B(n18089), .ZN(n17562) );
  XNOR2_X1 U11834 ( .A(n20639), .B(n20638), .ZN(n22139) );
  OAI21_X1 U11835 ( .B1(n21413), .B2(n22932), .A(n24309), .ZN(n21428) );
  INV_X1 U11836 ( .A(n19560), .ZN(n19141) );
  INV_X1 U11837 ( .A(n23305), .ZN(n22762) );
  NOR2_X1 U11839 ( .A1(n19238), .A2(n25086), .ZN(n18546) );
  AND2_X1 U11840 ( .A1(n22027), .A2(n24932), .ZN(n22934) );
  AND2_X1 U11843 ( .A1(n14327), .A2(n14325), .ZN(n13525) );
  OR2_X1 U11844 ( .A1(n21806), .A2(n23779), .ZN(n21807) );
  OR2_X1 U11845 ( .A1(n21467), .A2(n22968), .ZN(n21486) );
  AND2_X1 U11849 ( .A1(n23958), .A2(n22826), .ZN(n22827) );
  AND2_X1 U11850 ( .A1(n22940), .A2(n22938), .ZN(n22831) );
  OAI211_X1 U11852 ( .C1(n22675), .C2(n22674), .A(n22673), .B(n22672), .ZN(
        n23958) );
  AND2_X1 U11854 ( .A1(n25479), .A2(n25070), .ZN(n22190) );
  OR2_X1 U11855 ( .A1(n7541), .A2(n7757), .ZN(n7546) );
  AND2_X1 U11856 ( .A1(n22983), .A2(n23860), .ZN(n22984) );
  MUX2_X2 U11857 ( .A(n18760), .B(n18759), .S(n19265), .Z(n20343) );
  INV_X1 U11858 ( .A(n11955), .ZN(n11400) );
  NOR2_X1 U11859 ( .A1(n13828), .A2(n14116), .ZN(n13833) );
  INV_X1 U11860 ( .A(n23612), .ZN(n23648) );
  OAI21_X1 U11861 ( .B1(n12874), .B2(n13352), .A(n12330), .ZN(n13354) );
  XNOR2_X1 U11862 ( .A(n18471), .B(n18470), .ZN(n19578) );
  INV_X1 U11863 ( .A(n23361), .ZN(n23362) );
  OAI211_X1 U11864 ( .C1(n24941), .C2(n24059), .A(n23123), .B(n23091), .ZN(
        n23096) );
  INV_X1 U11865 ( .A(n17572), .ZN(n17371) );
  XNOR2_X1 U11866 ( .A(n7063), .B(n7062), .ZN(n7183) );
  AND2_X1 U11867 ( .A1(n18009), .A2(n19210), .ZN(n19042) );
  AND2_X1 U11869 ( .A1(n20556), .A2(n3480), .ZN(n19700) );
  NOR2_X1 U11870 ( .A1(n14318), .A2(n14317), .ZN(n14323) );
  AOI21_X1 U11873 ( .B1(n406), .B2(n13351), .A(n25430), .ZN(n12621) );
  XNOR2_X2 U11875 ( .A(n21991), .B(n21990), .ZN(n22893) );
  OR2_X1 U11876 ( .A1(n9531), .A2(n9805), .ZN(n10117) );
  OAI21_X1 U11877 ( .B1(n19616), .B2(n18546), .A(n19613), .ZN(n18547) );
  XNOR2_X1 U11878 ( .A(n11786), .B(n11785), .ZN(n12911) );
  AOI22_X1 U11879 ( .A1(n9360), .A2(n9950), .B1(n2876), .B2(n9270), .ZN(n10192) );
  AND2_X1 U11880 ( .A1(n19279), .A2(n19526), .ZN(n19282) );
  AND2_X1 U11881 ( .A1(n18795), .A2(n19526), .ZN(n18897) );
  OR2_X1 U11882 ( .A1(n10280), .A2(n10190), .ZN(n9268) );
  OR2_X1 U11883 ( .A1(n23157), .A2(n23129), .ZN(n23133) );
  INV_X1 U11884 ( .A(n19986), .ZN(n19684) );
  XNOR2_X1 U11885 ( .A(n20735), .B(n21110), .ZN(n22453) );
  OR2_X1 U11886 ( .A1(n25375), .A2(n22728), .ZN(n20892) );
  OR2_X1 U11887 ( .A1(n9462), .A2(n9461), .ZN(n9464) );
  OR2_X1 U11890 ( .A1(n13358), .A2(n12976), .ZN(n12584) );
  XNOR2_X2 U11891 ( .A(n18339), .B(n18338), .ZN(n19192) );
  NOR2_X2 U11892 ( .A1(n14197), .A2(n14196), .ZN(n15282) );
  MUX2_X2 U11893 ( .A(n10581), .B(n10580), .S(n10922), .Z(n12129) );
  NOR2_X1 U11894 ( .A1(n13272), .A2(n13275), .ZN(n12835) );
  OAI21_X2 U11895 ( .B1(n22716), .B2(n22715), .A(n22714), .ZN(n23479) );
  MUX2_X2 U11896 ( .A(n13362), .B(n13361), .S(n13364), .Z(n13683) );
  OR2_X1 U11898 ( .A1(n22842), .A2(n22847), .ZN(n21692) );
  OR2_X1 U11899 ( .A1(n24475), .A2(n7657), .ZN(n7660) );
  OR2_X1 U11900 ( .A1(n23720), .A2(n23714), .ZN(n22147) );
  OR2_X1 U11901 ( .A1(n20289), .A2(n20131), .ZN(n5728) );
  AND2_X1 U11902 ( .A1(n6621), .A2(n6619), .ZN(n5729) );
  AND2_X1 U11903 ( .A1(n10489), .A2(n10613), .ZN(n5730) );
  AND2_X1 U11904 ( .A1(n13347), .A2(n13348), .ZN(n5731) );
  OR3_X1 U11905 ( .A1(n23805), .A2(n21837), .A3(n24895), .ZN(n5732) );
  OR2_X1 U11906 ( .A1(n20062), .A2(n20055), .ZN(n5734) );
  AND2_X1 U11907 ( .A1(n11057), .A2(n11009), .ZN(n5735) );
  AND2_X1 U11908 ( .A1(n18933), .A2(n19327), .ZN(n5736) );
  OR2_X1 U11909 ( .A1(n7464), .A2(n7590), .ZN(n5737) );
  AND2_X1 U11910 ( .A1(n7278), .A2(n8021), .ZN(n5738) );
  INV_X1 U11911 ( .A(n9991), .ZN(n9657) );
  OR2_X1 U11912 ( .A1(n10127), .A2(n10132), .ZN(n5740) );
  OR3_X1 U11913 ( .A1(n9837), .A2(n10094), .A3(n10098), .ZN(n5741) );
  AND2_X1 U11914 ( .A1(n9820), .A2(n25463), .ZN(n5742) );
  XOR2_X1 U11915 ( .A(n9061), .B(n9060), .Z(n5743) );
  INV_X1 U11916 ( .A(n11069), .ZN(n10347) );
  XOR2_X1 U11917 ( .A(n11838), .B(n1835), .Z(n5745) );
  AND2_X1 U11918 ( .A1(n10364), .A2(n10682), .ZN(n5746) );
  OR2_X1 U11919 ( .A1(n13228), .A2(n12995), .ZN(n5747) );
  OR2_X1 U11920 ( .A1(n12794), .A2(n12792), .ZN(n5748) );
  INV_X1 U11921 ( .A(n12800), .ZN(n11580) );
  OR2_X1 U11922 ( .A1(n14326), .A2(n5230), .ZN(n5750) );
  NOR2_X1 U11923 ( .A1(n14127), .A2(n1331), .ZN(n5751) );
  AND2_X1 U11924 ( .A1(n14439), .A2(n13974), .ZN(n5752) );
  INV_X1 U11925 ( .A(n14439), .ZN(n14440) );
  AND4_X1 U11926 ( .A1(n13666), .A2(n13665), .A3(n14000), .A4(n13664), .ZN(
        n5753) );
  AND2_X1 U11927 ( .A1(n25033), .A2(n13132), .ZN(n5754) );
  OR2_X1 U11928 ( .A1(n13796), .A2(n13795), .ZN(n5755) );
  OR2_X1 U11929 ( .A1(n16067), .A2(n16060), .ZN(n5756) );
  XOR2_X1 U11930 ( .A(n15499), .B(n13405), .Z(n5757) );
  AND2_X1 U11931 ( .A1(n15977), .A2(n16394), .ZN(n5758) );
  OR2_X1 U11932 ( .A1(n17368), .A2(n17572), .ZN(n5759) );
  AND2_X1 U11933 ( .A1(n17069), .A2(n17067), .ZN(n5761) );
  XNOR2_X1 U11934 ( .A(n17999), .B(n17998), .ZN(n19041) );
  OR2_X1 U11935 ( .A1(n21370), .A2(n22615), .ZN(n5765) );
  AND2_X1 U11936 ( .A1(n22837), .A2(n22836), .ZN(n5766) );
  AND2_X1 U11937 ( .A1(n22333), .A2(n22137), .ZN(n5767) );
  AND2_X1 U11939 ( .A1(n21816), .A2(n22688), .ZN(n5770) );
  OR3_X1 U11940 ( .A1(n22939), .A2(n22832), .A3(n22027), .ZN(n5771) );
  OR2_X1 U11941 ( .A1(n23394), .A2(n24449), .ZN(n5772) );
  AND2_X1 U11942 ( .A1(n24954), .A2(n24011), .ZN(n5773) );
  OR2_X1 U11943 ( .A1(n24067), .A2(n4199), .ZN(n6261) );
  OR2_X1 U11944 ( .A1(n6919), .A2(n6915), .ZN(n5846) );
  INV_X1 U11945 ( .A(n6812), .ZN(n6371) );
  BUF_X1 U11946 ( .A(n6392), .Z(n6730) );
  OR2_X1 U11947 ( .A1(n6334), .A2(n6209), .ZN(n5949) );
  OAI22_X1 U11948 ( .A1(n6946), .A2(n6253), .B1(n5903), .B2(n5904), .ZN(n6526)
         );
  OR2_X1 U11949 ( .A1(n5863), .A2(n6531), .ZN(n6012) );
  OR2_X1 U11950 ( .A1(n6817), .A2(n6893), .ZN(n5830) );
  NOR2_X1 U11951 ( .A1(n6445), .A2(n6195), .ZN(n6344) );
  BUF_X1 U11952 ( .A(n6184), .Z(n6457) );
  OR2_X1 U11953 ( .A1(n7031), .A2(n7035), .ZN(n6227) );
  OR2_X1 U11954 ( .A1(n8514), .A2(n17960), .ZN(n8212) );
  BUF_X1 U11955 ( .A(n6497), .Z(n6503) );
  BUF_X1 U11956 ( .A(n6280), .Z(n7802) );
  AND2_X1 U11960 ( .A1(n6852), .A2(n6853), .ZN(n6854) );
  OR2_X1 U11961 ( .A1(n7821), .A2(n7820), .ZN(n7822) );
  INV_X1 U11962 ( .A(n8596), .ZN(n8597) );
  OR2_X1 U11963 ( .A1(n7345), .A2(n7256), .ZN(n7260) );
  INV_X1 U11964 ( .A(n8786), .ZN(n8552) );
  INV_X1 U11966 ( .A(n9711), .ZN(n9713) );
  OR2_X1 U11967 ( .A1(n24222), .A2(n10104), .ZN(n10106) );
  OR2_X1 U11968 ( .A1(n8534), .A2(n7667), .ZN(n7668) );
  XNOR2_X1 U11969 ( .A(n7706), .B(n7705), .ZN(n9345) );
  XNOR2_X1 U11970 ( .A(n8300), .B(n8299), .ZN(n8327) );
  AND2_X1 U11971 ( .A1(n9285), .A2(n9898), .ZN(n9288) );
  XNOR2_X1 U11972 ( .A(n8992), .B(n8993), .ZN(n9696) );
  AND2_X1 U11974 ( .A1(n9945), .A2(n9899), .ZN(n9445) );
  OR2_X1 U11976 ( .A1(n9934), .A2(n9599), .ZN(n9205) );
  INV_X1 U11978 ( .A(n9972), .ZN(n9975) );
  XNOR2_X1 U11980 ( .A(n8267), .B(n8266), .ZN(n8523) );
  OR2_X1 U11981 ( .A1(n9458), .A2(n9916), .ZN(n9275) );
  OR2_X1 U11982 ( .A1(n2953), .A2(n8142), .ZN(n8143) );
  OR2_X1 U11983 ( .A1(n10176), .A2(n10177), .ZN(n9830) );
  AND2_X1 U11984 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  BUF_X1 U11985 ( .A(n9462), .Z(n9920) );
  INV_X1 U11986 ( .A(n10836), .ZN(n9279) );
  OR2_X1 U11987 ( .A1(n10163), .A2(n24984), .ZN(n9593) );
  OR2_X1 U11988 ( .A1(n9864), .A2(n9860), .ZN(n9556) );
  INV_X1 U11989 ( .A(n9762), .ZN(n10072) );
  INV_X1 U11990 ( .A(n11143), .ZN(n11885) );
  INV_X1 U11991 ( .A(n9955), .ZN(n9959) );
  AND2_X1 U11992 ( .A1(n2244), .A2(n11122), .ZN(n11126) );
  INV_X1 U11993 ( .A(n10444), .ZN(n10749) );
  AND2_X1 U11994 ( .A1(n10969), .A2(n10967), .ZN(n9903) );
  INV_X1 U11995 ( .A(n10590), .ZN(n10372) );
  INV_X1 U11996 ( .A(n10405), .ZN(n10927) );
  OR2_X1 U11997 ( .A1(n11092), .A2(n11297), .ZN(n10895) );
  AND2_X1 U11998 ( .A1(n11059), .A2(n5735), .ZN(n10978) );
  NAND4_X1 U11999 ( .A1(n10965), .A2(n10964), .A3(n10963), .A4(n10962), .ZN(
        n12101) );
  OR2_X1 U12000 ( .A1(n10243), .A2(n10800), .ZN(n10249) );
  OAI21_X1 U12002 ( .B1(n11306), .B2(n11305), .A(n11304), .ZN(n11308) );
  INV_X1 U12003 ( .A(n13207), .ZN(n11360) );
  XNOR2_X1 U12004 ( .A(n11839), .B(n5745), .ZN(n11844) );
  XNOR2_X1 U12006 ( .A(n10640), .B(n10639), .ZN(n12663) );
  INV_X1 U12008 ( .A(n11965), .ZN(n13272) );
  AND2_X1 U12009 ( .A1(n12462), .A2(n13077), .ZN(n12709) );
  INV_X1 U12010 ( .A(n12892), .ZN(n12895) );
  OR2_X1 U12011 ( .A1(n4587), .A2(n12991), .ZN(n12998) );
  XNOR2_X1 U12012 ( .A(n11780), .B(n11779), .ZN(n12594) );
  INV_X1 U12013 ( .A(n14362), .ZN(n13088) );
  OR2_X1 U12014 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  INV_X1 U12015 ( .A(n14000), .ZN(n13487) );
  INV_X1 U12017 ( .A(n13236), .ZN(n13237) );
  OR2_X1 U12018 ( .A1(n13990), .A2(n13989), .ZN(n13991) );
  INV_X1 U12019 ( .A(n14153), .ZN(n13805) );
  OR2_X1 U12020 ( .A1(n13829), .A2(n13830), .ZN(n13401) );
  AND2_X1 U12022 ( .A1(n13997), .A2(n13995), .ZN(n14232) );
  INV_X1 U12023 ( .A(n2847), .ZN(n14879) );
  INV_X1 U12026 ( .A(n14880), .ZN(n15417) );
  OR2_X1 U12027 ( .A1(n13573), .A2(n13089), .ZN(n13091) );
  INV_X1 U12029 ( .A(n15454), .ZN(n15069) );
  XNOR2_X1 U12030 ( .A(n14985), .B(n14984), .ZN(n15774) );
  XNOR2_X1 U12031 ( .A(n15529), .B(n15530), .ZN(n15707) );
  OR2_X1 U12032 ( .A1(n16131), .A2(n15801), .ZN(n15595) );
  XNOR2_X1 U12034 ( .A(n15223), .B(n15002), .ZN(n15331) );
  OR2_X1 U12035 ( .A1(n16393), .A2(n16391), .ZN(n15980) );
  OR2_X1 U12036 ( .A1(n16030), .A2(n16029), .ZN(n16276) );
  OR2_X1 U12037 ( .A1(n16449), .A2(n16451), .ZN(n16239) );
  OR2_X1 U12038 ( .A1(n24366), .A2(n16266), .ZN(n16005) );
  INV_X1 U12039 ( .A(n17208), .ZN(n17207) );
  AND2_X1 U12040 ( .A1(n16422), .A2(n707), .ZN(n16174) );
  AOI21_X1 U12041 ( .B1(n15541), .B2(n294), .A(n15540), .ZN(n15542) );
  NOR2_X1 U12042 ( .A1(n16897), .A2(n17081), .ZN(n16898) );
  OR2_X1 U12043 ( .A1(n2636), .A2(n16241), .ZN(n15711) );
  OR2_X1 U12044 ( .A1(n17051), .A2(n17053), .ZN(n17002) );
  AOI22_X1 U12045 ( .A1(n15989), .A2(n15988), .B1(n15987), .B2(n16414), .ZN(
        n16765) );
  NOR2_X1 U12046 ( .A1(n16899), .A2(n16898), .ZN(n16900) );
  OAI21_X1 U12047 ( .B1(n17242), .B2(n17241), .A(n15314), .ZN(n16781) );
  OR2_X1 U12048 ( .A1(n17141), .A2(n17138), .ZN(n16694) );
  XNOR2_X1 U12049 ( .A(n18146), .B(n17772), .ZN(n17577) );
  AND2_X1 U12052 ( .A1(n20386), .A2(n19485), .ZN(n19344) );
  XNOR2_X1 U12053 ( .A(n17577), .B(n17578), .ZN(n17579) );
  INV_X1 U12054 ( .A(n19061), .ZN(n19056) );
  XNOR2_X1 U12055 ( .A(n18362), .B(n18361), .ZN(n18596) );
  XNOR2_X1 U12056 ( .A(n18664), .B(n18663), .ZN(n18690) );
  XNOR2_X1 U12057 ( .A(n18209), .B(n18208), .ZN(n18210) );
  XNOR2_X1 U12058 ( .A(n18059), .B(n18058), .ZN(n19587) );
  XNOR2_X1 U12059 ( .A(n18504), .B(n18503), .ZN(n19065) );
  AND2_X1 U12062 ( .A1(n19560), .A2(n19290), .ZN(n18752) );
  XNOR2_X1 U12063 ( .A(n18464), .B(n18463), .ZN(n18471) );
  OR2_X1 U12064 ( .A1(n20359), .A2(n20484), .ZN(n20487) );
  NOR2_X1 U12065 ( .A1(n24940), .A2(n20192), .ZN(n19744) );
  AND2_X1 U12066 ( .A1(n20560), .A2(n19731), .ZN(n19732) );
  NOR2_X1 U12067 ( .A1(n25012), .A2(n19065), .ZN(n19612) );
  OR2_X1 U12068 ( .A1(n19680), .A2(n19035), .ZN(n19050) );
  XNOR2_X1 U12070 ( .A(n17685), .B(n17684), .ZN(n19353) );
  NOR2_X1 U12071 ( .A1(n20409), .A2(n20411), .ZN(n19910) );
  OR2_X1 U12072 ( .A1(n19288), .A2(n19857), .ZN(n19292) );
  OAI21_X1 U12073 ( .B1(n19671), .B2(n24581), .A(n5728), .ZN(n19672) );
  OAI21_X1 U12074 ( .B1(n20337), .B2(n19708), .A(n19707), .ZN(n19712) );
  OAI211_X1 U12075 ( .C1(n18855), .C2(n18934), .A(n18854), .B(n18853), .ZN(
        n19195) );
  INV_X1 U12076 ( .A(n20173), .ZN(n20170) );
  INV_X1 U12077 ( .A(n20354), .ZN(n20355) );
  OR2_X1 U12078 ( .A1(n20141), .A2(n19975), .ZN(n20144) );
  XNOR2_X1 U12079 ( .A(n24434), .B(n21431), .ZN(n21432) );
  INV_X1 U12081 ( .A(n20222), .ZN(n19927) );
  INV_X1 U12082 ( .A(n22798), .ZN(n22584) );
  OR2_X1 U12085 ( .A1(n21920), .A2(n22752), .ZN(n22561) );
  BUF_X1 U12086 ( .A(n21908), .Z(n21910) );
  NOR2_X1 U12087 ( .A1(n22947), .A2(n22282), .ZN(n22945) );
  AND2_X1 U12089 ( .A1(n22209), .A2(n24333), .ZN(n20932) );
  AOI211_X1 U12090 ( .C1(n22800), .C2(n24559), .A(n22803), .B(n22798), .ZN(
        n22476) );
  BUF_X1 U12091 ( .A(n20776), .Z(n22400) );
  AND2_X1 U12092 ( .A1(n22952), .A2(n22954), .ZN(n22857) );
  NOR2_X1 U12093 ( .A1(n22726), .A2(n22725), .ZN(n23470) );
  AND3_X1 U12094 ( .A1(n22187), .A2(n22929), .A3(n22111), .ZN(n22112) );
  OR2_X1 U12095 ( .A1(n20940), .A2(n22066), .ZN(n20941) );
  OR2_X1 U12097 ( .A1(n22794), .A2(n24953), .ZN(n22795) );
  AND2_X1 U12098 ( .A1(n23052), .A2(n23040), .ZN(n22643) );
  INV_X1 U12102 ( .A(n23499), .ZN(n23484) );
  AND2_X1 U12103 ( .A1(n23647), .A2(n20896), .ZN(n20981) );
  OAI21_X1 U12104 ( .B1(n22598), .B2(n21855), .A(n21854), .ZN(n23869) );
  OAI21_X1 U12106 ( .B1(n22304), .B2(n5772), .A(n22303), .ZN(n22305) );
  OR2_X1 U12107 ( .A1(n23386), .A2(n24879), .ZN(n22884) );
  INV_X1 U12109 ( .A(n187), .ZN(n22049) );
  XNOR2_X1 U12110 ( .A(Key[76]), .B(Plaintext[76]), .ZN(n6744) );
  XNOR2_X1 U12111 ( .A(Key[73]), .B(Plaintext[73]), .ZN(n6050) );
  XNOR2_X1 U12112 ( .A(Key[72]), .B(Plaintext[72]), .ZN(n6407) );
  NAND2_X1 U12113 ( .A1(n6630), .A2(n6407), .ZN(n5776) );
  OAI21_X1 U12114 ( .B1(n453), .B2(n6630), .A(n5776), .ZN(n5777) );
  INV_X1 U12116 ( .A(n6051), .ZN(n6628) );
  INV_X1 U12117 ( .A(Plaintext[90]), .ZN(n5778) );
  XNOR2_X1 U12118 ( .A(n5778), .B(Key[90]), .ZN(n6235) );
  INV_X1 U12119 ( .A(Plaintext[91]), .ZN(n5779) );
  NAND2_X1 U12120 ( .A1(n6235), .A2(n6712), .ZN(n6112) );
  INV_X1 U12121 ( .A(Plaintext[95]), .ZN(n5780) );
  INV_X1 U12123 ( .A(Plaintext[92]), .ZN(n5781) );
  XNOR2_X1 U12124 ( .A(n5781), .B(Key[92]), .ZN(n6234) );
  INV_X1 U12125 ( .A(n6234), .ZN(n6232) );
  INV_X1 U12126 ( .A(Plaintext[94]), .ZN(n5782) );
  INV_X1 U12128 ( .A(n6233), .ZN(n6714) );
  INV_X1 U12130 ( .A(Plaintext[93]), .ZN(n5783) );
  NAND2_X1 U12131 ( .A1(n24051), .A2(n6712), .ZN(n5784) );
  INV_X1 U12132 ( .A(Plaintext[84]), .ZN(n5787) );
  XNOR2_X1 U12133 ( .A(n5787), .B(Key[84]), .ZN(n5795) );
  INV_X1 U12134 ( .A(Plaintext[87]), .ZN(n5788) );
  XNOR2_X1 U12135 ( .A(n5788), .B(Key[87]), .ZN(n5794) );
  NAND2_X1 U12136 ( .A1(n6619), .A2(n6623), .ZN(n5793) );
  INV_X1 U12137 ( .A(Plaintext[88]), .ZN(n5789) );
  INV_X1 U12138 ( .A(Plaintext[86]), .ZN(n5790) );
  NAND2_X1 U12139 ( .A1(n6622), .A2(n6049), .ZN(n5792) );
  INV_X1 U12140 ( .A(Plaintext[89]), .ZN(n5791) );
  INV_X1 U12141 ( .A(n6114), .ZN(n6723) );
  MUX2_X1 U12142 ( .A(n5793), .B(n5792), .S(n6723), .Z(n5799) );
  INV_X1 U12143 ( .A(n5795), .ZN(n6724) );
  MUX2_X1 U12144 ( .A(n6722), .B(n6243), .S(n6724), .Z(n5797) );
  NAND2_X1 U12145 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  OAI21_X1 U12149 ( .B1(n443), .B2(n6963), .A(n5800), .ZN(n5802) );
  NAND2_X1 U12151 ( .A1(n6965), .A2(n6964), .ZN(n5801) );
  XNOR2_X1 U12152 ( .A(Key[69]), .B(Plaintext[69]), .ZN(n6577) );
  INV_X1 U12153 ( .A(Plaintext[67]), .ZN(n5803) );
  NAND2_X1 U12154 ( .A1(n6752), .A2(n271), .ZN(n6754) );
  XNOR2_X1 U12155 ( .A(Key[70]), .B(Plaintext[70]), .ZN(n6757) );
  AND2_X1 U12156 ( .A1(n6757), .A2(n6578), .ZN(n5808) );
  XNOR2_X1 U12157 ( .A(Key[66]), .B(Plaintext[66]), .ZN(n6751) );
  NAND3_X1 U12159 ( .A1(n6675), .A2(n5804), .A3(n6578), .ZN(n5807) );
  XNOR2_X1 U12160 ( .A(Key[68]), .B(Plaintext[68]), .ZN(n6400) );
  NAND2_X1 U12161 ( .A1(n5805), .A2(n6755), .ZN(n5806) );
  NAND2_X1 U12162 ( .A1(n7576), .A2(n7579), .ZN(n5809) );
  XNOR2_X1 U12163 ( .A(Key[83]), .B(Plaintext[83]), .ZN(n6060) );
  INV_X1 U12164 ( .A(n6060), .ZN(n6393) );
  INV_X1 U12165 ( .A(Plaintext[81]), .ZN(n5810) );
  XNOR2_X1 U12166 ( .A(n5810), .B(Key[81]), .ZN(n6062) );
  INV_X1 U12167 ( .A(n6062), .ZN(n6729) );
  NAND2_X1 U12169 ( .A1(n6729), .A2(n6396), .ZN(n6736) );
  XNOR2_X1 U12171 ( .A(Key[80]), .B(Plaintext[80]), .ZN(n6392) );
  NAND2_X1 U12172 ( .A1(n6732), .A2(n6392), .ZN(n5812) );
  NAND2_X1 U12173 ( .A1(n5812), .A2(n6393), .ZN(n5811) );
  OAI21_X1 U12174 ( .B1(n6393), .B2(n6736), .A(n5811), .ZN(n5814) );
  INV_X1 U12175 ( .A(n6392), .ZN(n6615) );
  XNOR2_X1 U12176 ( .A(Key[82]), .B(Plaintext[82]), .ZN(n6238) );
  NAND3_X1 U12177 ( .A1(n6393), .A2(n6615), .A3(n6238), .ZN(n6242) );
  NOR2_X1 U12178 ( .A1(n5812), .A2(n2119), .ZN(n5813) );
  OR2_X1 U12179 ( .A1(n7577), .A2(n7576), .ZN(n7483) );
  MUX2_X1 U12180 ( .A(n4136), .B(n5815), .S(n7483), .Z(n5816) );
  XNOR2_X1 U12181 ( .A(Key[131]), .B(Plaintext[131]), .ZN(n6071) );
  INV_X1 U12182 ( .A(n6071), .ZN(n6815) );
  XNOR2_X1 U12183 ( .A(Key[130]), .B(Plaintext[130]), .ZN(n6369) );
  INV_X1 U12184 ( .A(n6369), .ZN(n6999) );
  INV_X1 U12185 ( .A(Plaintext[126]), .ZN(n5817) );
  XNOR2_X1 U12186 ( .A(Key[129]), .B(Plaintext[129]), .ZN(n6368) );
  AOI21_X1 U12187 ( .B1(n7003), .B2(n439), .A(n6997), .ZN(n5821) );
  XNOR2_X1 U12189 ( .A(Key[127]), .B(Plaintext[127]), .ZN(n6996) );
  AOI21_X1 U12190 ( .B1(n5819), .B2(n5818), .A(n6999), .ZN(n5820) );
  INV_X1 U12191 ( .A(Plaintext[146]), .ZN(n5822) );
  INV_X1 U12192 ( .A(Plaintext[149]), .ZN(n5823) );
  XNOR2_X1 U12193 ( .A(n5823), .B(Key[149]), .ZN(n6375) );
  NAND2_X1 U12194 ( .A1(n6377), .A2(n6375), .ZN(n6789) );
  XNOR2_X1 U12195 ( .A(Key[147]), .B(Plaintext[147]), .ZN(n6473) );
  INV_X1 U12196 ( .A(n6377), .ZN(n6374) );
  NAND3_X1 U12197 ( .A1(n6473), .A2(n6373), .A3(n6906), .ZN(n5825) );
  INV_X1 U12198 ( .A(n7887), .ZN(n5861) );
  XNOR2_X1 U12199 ( .A(Key[132]), .B(Plaintext[132]), .ZN(n6890) );
  INV_X1 U12200 ( .A(n6890), .ZN(n6819) );
  XNOR2_X1 U12201 ( .A(Key[133]), .B(Plaintext[133]), .ZN(n6086) );
  INV_X1 U12202 ( .A(n6086), .ZN(n6818) );
  NAND2_X1 U12203 ( .A1(n6819), .A2(n6818), .ZN(n6817) );
  INV_X1 U12204 ( .A(Plaintext[137]), .ZN(n5826) );
  INV_X1 U12205 ( .A(Plaintext[136]), .ZN(n5827) );
  XNOR2_X1 U12206 ( .A(n5827), .B(Key[136]), .ZN(n6651) );
  INV_X1 U12207 ( .A(Plaintext[135]), .ZN(n5828) );
  XNOR2_X2 U12208 ( .A(n5828), .B(Key[135]), .ZN(n6895) );
  INV_X1 U12209 ( .A(Plaintext[134]), .ZN(n5829) );
  INV_X1 U12211 ( .A(n6076), .ZN(n6882) );
  INV_X1 U12212 ( .A(Plaintext[142]), .ZN(n5831) );
  INV_X1 U12213 ( .A(n6795), .ZN(n6884) );
  XNOR2_X1 U12214 ( .A(Key[143]), .B(Plaintext[143]), .ZN(n5833) );
  BUF_X2 U12215 ( .A(n5833), .Z(n6885) );
  INV_X1 U12216 ( .A(n5833), .ZN(n6881) );
  INV_X1 U12217 ( .A(Plaintext[141]), .ZN(n5834) );
  XNOR2_X1 U12218 ( .A(n5834), .B(Key[141]), .ZN(n5835) );
  NAND3_X1 U12219 ( .A1(n6881), .A2(n6793), .A3(n6794), .ZN(n5838) );
  INV_X1 U12220 ( .A(n5835), .ZN(n6075) );
  INV_X1 U12221 ( .A(Key[140]), .ZN(n23151) );
  INV_X1 U12222 ( .A(Plaintext[140]), .ZN(n5836) );
  NAND4_X1 U12223 ( .A1(n6075), .A2(n6885), .A3(n23151), .A4(n5836), .ZN(n5837) );
  AND2_X1 U12224 ( .A1(n5837), .A2(n5838), .ZN(n5843) );
  INV_X1 U12225 ( .A(Plaintext[138]), .ZN(n5839) );
  NAND3_X1 U12226 ( .A1(n5833), .A2(Key[140]), .A3(Plaintext[140]), .ZN(n5840)
         );
  OAI21_X1 U12227 ( .B1(n6078), .B2(n6885), .A(n5840), .ZN(n5841) );
  NAND2_X1 U12228 ( .A1(n5841), .A2(n6075), .ZN(n5842) );
  OAI21_X1 U12229 ( .B1(n7879), .B2(n7585), .A(n7313), .ZN(n5860) );
  INV_X1 U12230 ( .A(Plaintext[160]), .ZN(n5844) );
  XNOR2_X1 U12231 ( .A(Key[156]), .B(Plaintext[156]), .ZN(n6917) );
  INV_X1 U12232 ( .A(n6917), .ZN(n6916) );
  AOI21_X1 U12233 ( .B1(n5846), .B2(n5845), .A(n6918), .ZN(n5850) );
  INV_X1 U12234 ( .A(Plaintext[161]), .ZN(n5847) );
  NAND3_X1 U12235 ( .A1(n6912), .A2(n6770), .A3(n6919), .ZN(n5848) );
  OAI21_X1 U12236 ( .B1(n6916), .B2(n24037), .A(n5848), .ZN(n5849) );
  INV_X1 U12237 ( .A(Plaintext[154]), .ZN(n5851) );
  XNOR2_X1 U12238 ( .A(Key[155]), .B(Plaintext[155]), .ZN(n6081) );
  NAND2_X1 U12239 ( .A1(n6767), .A2(n6876), .ZN(n5855) );
  INV_X1 U12240 ( .A(Plaintext[150]), .ZN(n5852) );
  XNOR2_X1 U12241 ( .A(n5852), .B(Key[150]), .ZN(n6083) );
  INV_X1 U12242 ( .A(n6083), .ZN(n6875) );
  INV_X1 U12243 ( .A(Plaintext[151]), .ZN(n5853) );
  XNOR2_X1 U12244 ( .A(n5853), .B(Key[151]), .ZN(n6310) );
  INV_X1 U12245 ( .A(n6310), .ZN(n6870) );
  NAND2_X1 U12246 ( .A1(n6875), .A2(n6870), .ZN(n5854) );
  XNOR2_X1 U12247 ( .A(Key[152]), .B(Plaintext[152]), .ZN(n6871) );
  NAND2_X1 U12249 ( .A1(n5856), .A2(n6083), .ZN(n5857) );
  AND2_X1 U12250 ( .A1(n5858), .A2(n5857), .ZN(n7584) );
  XNOR2_X1 U12252 ( .A(n8596), .B(n8666), .ZN(n8249) );
  INV_X1 U12253 ( .A(Plaintext[28]), .ZN(n5862) );
  INV_X1 U12254 ( .A(n6532), .ZN(n5863) );
  INV_X1 U12255 ( .A(Plaintext[24]), .ZN(n5864) );
  XNOR2_X1 U12256 ( .A(n5864), .B(Key[24]), .ZN(n6013) );
  INV_X1 U12257 ( .A(n6013), .ZN(n6538) );
  AOI21_X1 U12258 ( .B1(n6012), .B2(n6538), .A(n6530), .ZN(n5869) );
  INV_X1 U12259 ( .A(Plaintext[26]), .ZN(n5865) );
  INV_X1 U12260 ( .A(n6531), .ZN(n6259) );
  NAND2_X1 U12262 ( .A1(n4199), .A2(n6530), .ZN(n5866) );
  AOI21_X1 U12263 ( .B1(n5867), .B2(n5866), .A(n6532), .ZN(n5868) );
  INV_X1 U12264 ( .A(Plaintext[46]), .ZN(n5870) );
  XNOR2_X1 U12266 ( .A(Key[43]), .B(Plaintext[43]), .ZN(n6703) );
  XNOR2_X1 U12267 ( .A(Key[47]), .B(Plaintext[47]), .ZN(n6705) );
  INV_X1 U12268 ( .A(n6705), .ZN(n6960) );
  INV_X1 U12269 ( .A(Plaintext[42]), .ZN(n5871) );
  INV_X1 U12270 ( .A(n5924), .ZN(n6957) );
  XNOR2_X2 U12271 ( .A(Key[45]), .B(Plaintext[45]), .ZN(n6959) );
  XNOR2_X1 U12273 ( .A(Key[57]), .B(Plaintext[57]), .ZN(n6066) );
  INV_X1 U12274 ( .A(n6066), .ZN(n6971) );
  INV_X1 U12275 ( .A(Plaintext[55]), .ZN(n5872) );
  INV_X1 U12278 ( .A(Plaintext[56]), .ZN(n5873) );
  INV_X1 U12279 ( .A(Plaintext[58]), .ZN(n5874) );
  NAND2_X1 U12282 ( .A1(n6692), .A2(n6977), .ZN(n5875) );
  INV_X1 U12283 ( .A(Plaintext[30]), .ZN(n5877) );
  INV_X1 U12284 ( .A(n6529), .ZN(n6946) );
  INV_X1 U12285 ( .A(Plaintext[31]), .ZN(n5878) );
  XNOR2_X1 U12286 ( .A(n5878), .B(Key[31]), .ZN(n5902) );
  INV_X1 U12287 ( .A(n5902), .ZN(n6253) );
  INV_X1 U12288 ( .A(Plaintext[32]), .ZN(n5879) );
  INV_X1 U12289 ( .A(n5904), .ZN(n6255) );
  XNOR2_X1 U12290 ( .A(Key[33]), .B(Plaintext[33]), .ZN(n6948) );
  NAND2_X1 U12291 ( .A1(n6253), .A2(n6948), .ZN(n6139) );
  INV_X1 U12292 ( .A(n6139), .ZN(n5882) );
  INV_X1 U12293 ( .A(Plaintext[34]), .ZN(n5880) );
  AOI22_X1 U12295 ( .A1(n6526), .A2(n6953), .B1(n5882), .B2(n5881), .ZN(n7327)
         );
  XNOR2_X1 U12296 ( .A(Key[39]), .B(Plaintext[39]), .ZN(n5887) );
  INV_X1 U12297 ( .A(n5887), .ZN(n6684) );
  XNOR2_X1 U12298 ( .A(Key[37]), .B(Plaintext[37]), .ZN(n5910) );
  INV_X1 U12299 ( .A(n5910), .ZN(n6680) );
  XNOR2_X1 U12300 ( .A(Key[36]), .B(Plaintext[36]), .ZN(n6146) );
  NOR2_X1 U12301 ( .A1(n6684), .A2(n6146), .ZN(n5883) );
  XNOR2_X1 U12302 ( .A(Key[41]), .B(Plaintext[41]), .ZN(n5888) );
  INV_X1 U12303 ( .A(n5888), .ZN(n6944) );
  OAI21_X1 U12304 ( .B1(n5884), .B2(n5883), .A(n6944), .ZN(n5890) );
  INV_X1 U12305 ( .A(Plaintext[38]), .ZN(n5885) );
  XNOR2_X1 U12306 ( .A(n5885), .B(Key[38]), .ZN(n5908) );
  INV_X1 U12307 ( .A(Plaintext[40]), .ZN(n5886) );
  INV_X1 U12309 ( .A(n5908), .ZN(n6281) );
  INV_X1 U12310 ( .A(Plaintext[51]), .ZN(n5891) );
  XNOR2_X1 U12311 ( .A(n5891), .B(Key[51]), .ZN(n6414) );
  XNOR2_X1 U12313 ( .A(Key[49]), .B(Plaintext[49]), .ZN(n6694) );
  INV_X1 U12314 ( .A(n6694), .ZN(n5893) );
  INV_X1 U12315 ( .A(Plaintext[48]), .ZN(n5892) );
  INV_X1 U12316 ( .A(n6556), .ZN(n6693) );
  MUX2_X1 U12317 ( .A(n6695), .B(n5893), .S(n6693), .Z(n5900) );
  INV_X1 U12318 ( .A(Plaintext[50]), .ZN(n5894) );
  NAND2_X1 U12319 ( .A1(n6695), .A2(n6556), .ZN(n5898) );
  INV_X1 U12320 ( .A(Plaintext[52]), .ZN(n5895) );
  INV_X1 U12321 ( .A(Plaintext[53]), .ZN(n5896) );
  MUX2_X1 U12322 ( .A(n5898), .B(n5897), .S(n6934), .Z(n5899) );
  XNOR2_X1 U12323 ( .A(n8412), .B(n860), .ZN(n5930) );
  INV_X1 U12324 ( .A(n5903), .ZN(n6528) );
  INV_X1 U12325 ( .A(n6948), .ZN(n6947) );
  NAND2_X1 U12326 ( .A1(n5908), .A2(n6683), .ZN(n5909) );
  MUX2_X1 U12327 ( .A(n7250), .B(n8508), .S(n8512), .Z(n8209) );
  INV_X1 U12328 ( .A(Plaintext[18]), .ZN(n5913) );
  XNOR2_X1 U12329 ( .A(Key[21]), .B(Plaintext[21]), .ZN(n6267) );
  INV_X1 U12330 ( .A(Plaintext[19]), .ZN(n5914) );
  XNOR2_X1 U12331 ( .A(n5914), .B(Key[19]), .ZN(n5915) );
  INV_X1 U12332 ( .A(n5915), .ZN(n6539) );
  XNOR2_X1 U12333 ( .A(Key[23]), .B(Plaintext[23]), .ZN(n6133) );
  INV_X1 U12334 ( .A(n6267), .ZN(n7103) );
  XNOR2_X1 U12335 ( .A(Key[22]), .B(Plaintext[22]), .ZN(n7101) );
  INV_X1 U12336 ( .A(n5916), .ZN(n6266) );
  NAND2_X1 U12338 ( .A1(n127), .A2(n6164), .ZN(n5917) );
  NAND2_X1 U12339 ( .A1(n6530), .A2(n6533), .ZN(n5918) );
  AOI21_X1 U12340 ( .B1(n5918), .B2(n24067), .A(n6531), .ZN(n5923) );
  NAND3_X1 U12341 ( .A1(n4199), .A2(n25014), .A3(n6531), .ZN(n5921) );
  NAND2_X1 U12342 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  AND2_X1 U12343 ( .A1(n7350), .A2(n7346), .ZN(n5929) );
  NAND2_X1 U12344 ( .A1(n6956), .A2(n24405), .ZN(n6137) );
  INV_X1 U12345 ( .A(n6959), .ZN(n6553) );
  NAND2_X1 U12346 ( .A1(n6553), .A2(n6705), .ZN(n5925) );
  NAND2_X1 U12347 ( .A1(n24405), .A2(n6959), .ZN(n6954) );
  NAND3_X1 U12348 ( .A1(n5925), .A2(n6954), .A3(n5924), .ZN(n5927) );
  NAND3_X1 U12349 ( .A1(n3926), .A2(n6703), .A3(n3922), .ZN(n5926) );
  OAI211_X1 U12350 ( .C1(n6137), .C2(n6960), .A(n5927), .B(n5926), .ZN(n7348)
         );
  OAI21_X1 U12351 ( .B1(n7250), .B2(n5929), .A(n5928), .ZN(n8514) );
  OAI21_X1 U12352 ( .B1(n8209), .B2(n7350), .A(n8514), .ZN(n9175) );
  INV_X1 U12353 ( .A(n6445), .ZN(n6019) );
  XNOR2_X1 U12354 ( .A(Key[186]), .B(Plaintext[186]), .ZN(n6444) );
  INV_X1 U12355 ( .A(n6444), .ZN(n6345) );
  INV_X1 U12356 ( .A(n6021), .ZN(n5935) );
  INV_X1 U12358 ( .A(n6452), .ZN(n6341) );
  OAI21_X1 U12359 ( .B1(n6345), .B2(n6195), .A(n6341), .ZN(n5934) );
  XNOR2_X1 U12360 ( .A(Key[190]), .B(Plaintext[190]), .ZN(n6447) );
  INV_X1 U12361 ( .A(n6447), .ZN(n6196) );
  NAND2_X1 U12362 ( .A1(n6196), .A2(n6452), .ZN(n5932) );
  INV_X1 U12363 ( .A(Plaintext[191]), .ZN(n5931) );
  INV_X1 U12365 ( .A(n6187), .ZN(n6449) );
  MUX2_X1 U12366 ( .A(n6021), .B(n5932), .S(n6449), .Z(n5933) );
  INV_X1 U12367 ( .A(n7464), .ZN(n7587) );
  INV_X1 U12368 ( .A(Plaintext[3]), .ZN(n5936) );
  INV_X1 U12370 ( .A(Plaintext[1]), .ZN(n5937) );
  AND2_X1 U12371 ( .A1(n6513), .A2(n6456), .ZN(n6183) );
  INV_X1 U12372 ( .A(n6183), .ZN(n5939) );
  INV_X1 U12373 ( .A(n6455), .ZN(n6454) );
  INV_X1 U12374 ( .A(Plaintext[2]), .ZN(n5938) );
  XNOR2_X1 U12375 ( .A(n5938), .B(Key[2]), .ZN(n6184) );
  INV_X1 U12376 ( .A(n6184), .ZN(n6509) );
  AOI21_X1 U12377 ( .B1(n5939), .B2(n6454), .A(n6509), .ZN(n5942) );
  INV_X1 U12378 ( .A(Plaintext[5]), .ZN(n5940) );
  NAND2_X1 U12379 ( .A1(n6509), .A2(n6510), .ZN(n6030) );
  XNOR2_X1 U12380 ( .A(Key[4]), .B(Plaintext[4]), .ZN(n6512) );
  NOR2_X1 U12381 ( .A1(n7587), .A2(n7590), .ZN(n5970) );
  INV_X1 U12382 ( .A(Plaintext[182]), .ZN(n5943) );
  INV_X1 U12383 ( .A(Plaintext[181]), .ZN(n5944) );
  INV_X1 U12385 ( .A(n6297), .ZN(n6209) );
  INV_X1 U12386 ( .A(Plaintext[184]), .ZN(n5945) );
  XNOR2_X1 U12387 ( .A(n5945), .B(Key[184]), .ZN(n6332) );
  NAND2_X1 U12388 ( .A1(n6335), .A2(n6332), .ZN(n6173) );
  XNOR2_X1 U12389 ( .A(Key[180]), .B(Plaintext[180]), .ZN(n6208) );
  INV_X1 U12390 ( .A(n6335), .ZN(n6439) );
  XNOR2_X2 U12391 ( .A(Key[173]), .B(Plaintext[173]), .ZN(n6493) );
  INV_X1 U12392 ( .A(Plaintext[170]), .ZN(n5950) );
  INV_X1 U12394 ( .A(Plaintext[171]), .ZN(n5951) );
  INV_X1 U12395 ( .A(n6427), .ZN(n6301) );
  INV_X1 U12396 ( .A(Plaintext[169]), .ZN(n5952) );
  INV_X1 U12397 ( .A(n6488), .ZN(n6304) );
  NAND2_X1 U12398 ( .A1(n6781), .A2(n5953), .ZN(n5956) );
  INV_X1 U12399 ( .A(Plaintext[172]), .ZN(n5954) );
  INV_X1 U12401 ( .A(n6490), .ZN(n6780) );
  NAND2_X1 U12402 ( .A1(n6493), .A2(n6780), .ZN(n5955) );
  NAND2_X1 U12403 ( .A1(n5956), .A2(n5955), .ZN(n5960) );
  INV_X1 U12404 ( .A(Plaintext[168]), .ZN(n5957) );
  XNOR2_X1 U12405 ( .A(n5957), .B(Key[168]), .ZN(n6784) );
  NAND2_X1 U12406 ( .A1(n6784), .A2(n6488), .ZN(n6782) );
  INV_X1 U12407 ( .A(n6782), .ZN(n5958) );
  NAND2_X1 U12408 ( .A1(n5958), .A2(n6493), .ZN(n5959) );
  NAND2_X1 U12409 ( .A1(n5960), .A2(n5959), .ZN(n7335) );
  XNOR2_X1 U12410 ( .A(Key[162]), .B(Plaintext[162]), .ZN(n6777) );
  INV_X1 U12411 ( .A(Plaintext[163]), .ZN(n5961) );
  INV_X1 U12412 ( .A(Plaintext[164]), .ZN(n5962) );
  INV_X1 U12413 ( .A(Plaintext[166]), .ZN(n5963) );
  XNOR2_X1 U12414 ( .A(n5963), .B(Key[166]), .ZN(n6776) );
  INV_X1 U12415 ( .A(Plaintext[177]), .ZN(n5965) );
  INV_X1 U12416 ( .A(n5966), .ZN(n6315) );
  INV_X1 U12418 ( .A(Plaintext[174]), .ZN(n5967) );
  XNOR2_X1 U12419 ( .A(n5967), .B(Key[174]), .ZN(n6470) );
  INV_X1 U12420 ( .A(n6470), .ZN(n6329) );
  INV_X1 U12421 ( .A(Plaintext[175]), .ZN(n5968) );
  NAND2_X1 U12422 ( .A1(n4621), .A2(n6426), .ZN(n6471) );
  INV_X1 U12423 ( .A(Plaintext[179]), .ZN(n5969) );
  NOR2_X1 U12424 ( .A1(n7593), .A2(n5971), .ZN(n5972) );
  XNOR2_X1 U12425 ( .A(Key[110]), .B(Plaintext[110]), .ZN(n6245) );
  AND2_X1 U12426 ( .A1(n6245), .A2(n6244), .ZN(n5975) );
  XNOR2_X1 U12427 ( .A(Key[113]), .B(Plaintext[113]), .ZN(n6122) );
  XNOR2_X1 U12428 ( .A(Key[108]), .B(Plaintext[108]), .ZN(n6119) );
  NAND2_X1 U12429 ( .A1(n6122), .A2(n6119), .ZN(n5973) );
  NAND2_X1 U12430 ( .A1(n5973), .A2(n6987), .ZN(n5974) );
  INV_X1 U12431 ( .A(n6245), .ZN(n6841) );
  XNOR2_X1 U12432 ( .A(Key[112]), .B(Plaintext[112]), .ZN(n6640) );
  INV_X1 U12433 ( .A(n5975), .ZN(n5976) );
  INV_X1 U12434 ( .A(n6122), .ZN(n6986) );
  NAND3_X1 U12435 ( .A1(n6639), .A2(n5976), .A3(n6986), .ZN(n5977) );
  INV_X1 U12436 ( .A(Plaintext[121]), .ZN(n5979) );
  INV_X1 U12437 ( .A(Plaintext[120]), .ZN(n5980) );
  XNOR2_X1 U12438 ( .A(n5980), .B(Key[120]), .ZN(n6647) );
  AND2_X1 U12439 ( .A1(n6647), .A2(n7004), .ZN(n6384) );
  XNOR2_X1 U12440 ( .A(Key[124]), .B(Plaintext[124]), .ZN(n6094) );
  INV_X1 U12441 ( .A(n6094), .ZN(n6650) );
  NAND2_X1 U12442 ( .A1(n6384), .A2(n6650), .ZN(n5985) );
  NAND3_X1 U12443 ( .A1(n7006), .A2(n7004), .A3(n448), .ZN(n5984) );
  INV_X1 U12444 ( .A(Plaintext[125]), .ZN(n5981) );
  AND2_X1 U12445 ( .A1(n7007), .A2(n6648), .ZN(n6836) );
  NAND2_X1 U12446 ( .A1(n6836), .A2(n6650), .ZN(n5983) );
  INV_X1 U12447 ( .A(n6647), .ZN(n7009) );
  NAND3_X1 U12449 ( .A1(n24051), .A2(n6233), .A3(n24500), .ZN(n5988) );
  NAND3_X1 U12450 ( .A1(n6234), .A2(n24501), .A3(n6714), .ZN(n5987) );
  INV_X1 U12451 ( .A(n24050), .ZN(n6611) );
  NAND3_X1 U12452 ( .A1(n6712), .A2(n6611), .A3(n6714), .ZN(n5986) );
  INV_X1 U12453 ( .A(n5992), .ZN(n7019) );
  INV_X1 U12454 ( .A(Plaintext[102]), .ZN(n5989) );
  XNOR2_X1 U12455 ( .A(n5989), .B(Key[102]), .ZN(n6598) );
  INV_X1 U12456 ( .A(Plaintext[105]), .ZN(n5990) );
  INV_X1 U12457 ( .A(n6823), .ZN(n7015) );
  NAND3_X1 U12458 ( .A1(n7019), .A2(n6598), .A3(n7015), .ZN(n5996) );
  INV_X1 U12459 ( .A(Plaintext[104]), .ZN(n5991) );
  NAND2_X1 U12460 ( .A1(n25044), .A2(n5992), .ZN(n5995) );
  NAND2_X1 U12461 ( .A1(n6823), .A2(n5992), .ZN(n5994) );
  INV_X1 U12462 ( .A(Plaintext[103]), .ZN(n5993) );
  XNOR2_X1 U12463 ( .A(Key[106]), .B(Plaintext[106]), .ZN(n7013) );
  NAND2_X1 U12464 ( .A1(n6100), .A2(n6824), .ZN(n5997) );
  INV_X1 U12466 ( .A(n7026), .ZN(n6846) );
  XNOR2_X1 U12467 ( .A(Key[117]), .B(Plaintext[117]), .ZN(n6845) );
  INV_X1 U12468 ( .A(n6845), .ZN(n7022) );
  INV_X1 U12469 ( .A(Plaintext[119]), .ZN(n5999) );
  XNOR2_X1 U12470 ( .A(n5999), .B(Key[119]), .ZN(n6381) );
  INV_X1 U12471 ( .A(Plaintext[116]), .ZN(n6000) );
  INV_X1 U12473 ( .A(n7021), .ZN(n7024) );
  NAND2_X1 U12474 ( .A1(n7024), .A2(n7026), .ZN(n6001) );
  INV_X1 U12475 ( .A(Plaintext[118]), .ZN(n6002) );
  INV_X1 U12476 ( .A(n6849), .ZN(n7023) );
  NAND3_X1 U12477 ( .A1(n6848), .A2(n7023), .A3(n442), .ZN(n6003) );
  XNOR2_X1 U12479 ( .A(Key[98]), .B(Plaintext[98]), .ZN(n6104) );
  INV_X1 U12480 ( .A(Plaintext[101]), .ZN(n6004) );
  OAI21_X1 U12481 ( .B1(n7032), .B2(n6588), .A(n6005), .ZN(n6740) );
  NAND2_X1 U12483 ( .A1(n6740), .A2(n7031), .ZN(n6006) );
  NAND2_X1 U12484 ( .A1(n6006), .A2(n6225), .ZN(n6009) );
  INV_X1 U12485 ( .A(n6740), .ZN(n6007) );
  NAND3_X1 U12486 ( .A1(n6007), .A2(n7033), .A3(n7035), .ZN(n6008) );
  NAND2_X1 U12487 ( .A1(n24067), .A2(n6538), .ZN(n6011) );
  OAI21_X1 U12488 ( .B1(n6012), .B2(n24592), .A(n6011), .ZN(n6017) );
  NAND2_X1 U12489 ( .A1(n6532), .A2(n25014), .ZN(n6014) );
  AOI21_X1 U12490 ( .B1(n6015), .B2(n6014), .A(n24254), .ZN(n6016) );
  OR2_X2 U12491 ( .A1(n6017), .A2(n6016), .ZN(n7600) );
  INV_X1 U12493 ( .A(n6195), .ZN(n6450) );
  NAND2_X1 U12494 ( .A1(n6450), .A2(n6445), .ZN(n6018) );
  AOI21_X1 U12495 ( .B1(n6448), .B2(n6018), .A(n6196), .ZN(n6022) );
  INV_X1 U12496 ( .A(Plaintext[17]), .ZN(n6023) );
  INV_X1 U12498 ( .A(Plaintext[16]), .ZN(n6024) );
  XNOR2_X1 U12499 ( .A(n6024), .B(Key[16]), .ZN(n6324) );
  INV_X1 U12500 ( .A(Plaintext[15]), .ZN(n6025) );
  INV_X1 U12501 ( .A(n6519), .ZN(n6156) );
  INV_X1 U12502 ( .A(Plaintext[12]), .ZN(n6026) );
  XNOR2_X1 U12503 ( .A(n6026), .B(Key[12]), .ZN(n6179) );
  INV_X1 U12504 ( .A(n6179), .ZN(n6323) );
  INV_X1 U12505 ( .A(n6518), .ZN(n6027) );
  INV_X1 U12506 ( .A(n6275), .ZN(n6274) );
  NAND2_X1 U12507 ( .A1(n6027), .A2(n6274), .ZN(n6029) );
  XNOR2_X1 U12508 ( .A(Key[13]), .B(Plaintext[13]), .ZN(n6523) );
  NAND2_X1 U12509 ( .A1(n7595), .A2(n7602), .ZN(n6802) );
  NOR2_X1 U12510 ( .A1(n7135), .A2(n7602), .ZN(n6039) );
  INV_X1 U12511 ( .A(n6510), .ZN(n6459) );
  INV_X1 U12513 ( .A(n6512), .ZN(n6460) );
  NOR2_X1 U12514 ( .A1(n6513), .A2(n6456), .ZN(n6506) );
  OAI21_X1 U12515 ( .B1(n6510), .B2(n6460), .A(n6506), .ZN(n6031) );
  NOR2_X1 U12516 ( .A1(n7595), .A2(n7257), .ZN(n6038) );
  INV_X1 U12517 ( .A(Plaintext[10]), .ZN(n6033) );
  XNOR2_X1 U12518 ( .A(n6033), .B(Key[10]), .ZN(n6496) );
  NAND2_X1 U12519 ( .A1(n6271), .A2(n6034), .ZN(n6169) );
  INV_X1 U12520 ( .A(Plaintext[7]), .ZN(n6035) );
  OAI21_X1 U12521 ( .B1(n6351), .B2(n6498), .A(n6168), .ZN(n6037) );
  INV_X1 U12522 ( .A(Plaintext[11]), .ZN(n6036) );
  XNOR2_X1 U12523 ( .A(n6036), .B(Key[11]), .ZN(n6497) );
  OAI21_X1 U12524 ( .B1(n6039), .B2(n6038), .A(n7598), .ZN(n6045) );
  INV_X1 U12525 ( .A(n6133), .ZN(n6136) );
  OAI211_X1 U12526 ( .C1(n6136), .C2(n6164), .A(n6265), .B(n7097), .ZN(n6043)
         );
  NAND2_X1 U12527 ( .A1(n6266), .A2(n6539), .ZN(n6040) );
  NAND3_X1 U12528 ( .A1(n7255), .A2(n24772), .A3(n7597), .ZN(n6044) );
  XNOR2_X1 U12529 ( .A(n310), .B(n9181), .ZN(n6046) );
  XNOR2_X1 U12530 ( .A(n9011), .B(n6046), .ZN(n6047) );
  XNOR2_X1 U12531 ( .A(n6048), .B(n6047), .ZN(n9460) );
  OAI211_X1 U12532 ( .C1(n6750), .C2(n6409), .A(n6054), .B(n6053), .ZN(n6056)
         );
  NAND3_X1 U12533 ( .A1(n6630), .A2(n6407), .A3(n6051), .ZN(n6055) );
  OAI21_X1 U12534 ( .B1(n6964), .B2(n6963), .A(n6057), .ZN(n6967) );
  NAND2_X1 U12536 ( .A1(n6570), .A2(n24089), .ZN(n6576) );
  NAND2_X1 U12537 ( .A1(n5800), .A2(n6963), .ZN(n6572) );
  NAND2_X1 U12538 ( .A1(n4754), .A2(n6575), .ZN(n6059) );
  MUX2_X1 U12539 ( .A(n7747), .B(n8021), .S(n8022), .Z(n6070) );
  NAND2_X1 U12540 ( .A1(n6393), .A2(n6396), .ZN(n6061) );
  MUX2_X1 U12543 ( .A(n6729), .B(n6732), .S(n6396), .Z(n6063) );
  NAND2_X1 U12544 ( .A1(n6692), .A2(n6975), .ZN(n6069) );
  INV_X1 U12545 ( .A(n6976), .ZN(n6568) );
  AND2_X1 U12547 ( .A1(n6368), .A2(n6996), .ZN(n6657) );
  NAND2_X1 U12548 ( .A1(n6815), .A2(n6072), .ZN(n6073) );
  NAND2_X1 U12549 ( .A1(n6075), .A2(n6794), .ZN(n6883) );
  INV_X1 U12550 ( .A(n6794), .ZN(n6644) );
  NAND2_X1 U12551 ( .A1(n6644), .A2(n6885), .ZN(n6077) );
  NAND3_X1 U12552 ( .A1(n6882), .A2(n6881), .A3(n6795), .ZN(n6080) );
  INV_X1 U12553 ( .A(n6078), .ZN(n6792) );
  NAND3_X1 U12554 ( .A1(n6075), .A2(n6885), .A3(n6792), .ZN(n6079) );
  NOR2_X1 U12555 ( .A1(n7754), .A2(n7292), .ZN(n7755) );
  INV_X1 U12556 ( .A(n6081), .ZN(n6768) );
  NAND2_X1 U12557 ( .A1(n6768), .A2(n6871), .ZN(n6873) );
  AND2_X1 U12558 ( .A1(n6083), .A2(n6310), .ZN(n6477) );
  INV_X1 U12559 ( .A(n6477), .ZN(n6082) );
  NAND2_X1 U12560 ( .A1(n6873), .A2(n6082), .ZN(n6085) );
  OAI21_X1 U12561 ( .B1(n6874), .B2(n6870), .A(n6083), .ZN(n6084) );
  OAI21_X1 U12562 ( .B1(n2522), .B2(n7542), .A(n432), .ZN(n6098) );
  INV_X1 U12563 ( .A(n6373), .ZN(n6088) );
  NAND2_X1 U12564 ( .A1(n6087), .A2(n6377), .ZN(n6093) );
  INV_X1 U12565 ( .A(n6473), .ZN(n6902) );
  MUX2_X1 U12567 ( .A(n6091), .B(n6090), .S(n6906), .Z(n6092) );
  NAND2_X1 U12568 ( .A1(n7006), .A2(n7007), .ZN(n6383) );
  INV_X1 U12569 ( .A(n6383), .ZN(n6096) );
  INV_X1 U12570 ( .A(n7004), .ZN(n6832) );
  OAI21_X1 U12571 ( .B1(n6096), .B2(n6095), .A(n6094), .ZN(n6097) );
  XNOR2_X1 U12572 ( .A(n8674), .B(n8604), .ZN(n8256) );
  INV_X1 U12573 ( .A(n6602), .ZN(n7012) );
  INV_X1 U12574 ( .A(n6827), .ZN(n7014) );
  NAND2_X1 U12575 ( .A1(n7012), .A2(n7014), .ZN(n6101) );
  INV_X1 U12576 ( .A(n6598), .ZN(n6601) );
  MUX2_X1 U12577 ( .A(n6101), .B(n6099), .S(n7015), .Z(n6103) );
  NAND3_X1 U12578 ( .A1(n6826), .A2(n6101), .A3(n7019), .ZN(n6102) );
  NAND2_X1 U12579 ( .A1(n6104), .A2(n7029), .ZN(n6593) );
  NAND2_X1 U12580 ( .A1(n6593), .A2(n6105), .ZN(n6108) );
  NAND2_X1 U12581 ( .A1(n7029), .A2(n7032), .ZN(n6106) );
  OAI21_X1 U12582 ( .B1(n7030), .B2(n7029), .A(n6106), .ZN(n6107) );
  AND2_X1 U12583 ( .A1(n7768), .A2(n7526), .ZN(n6113) );
  OAI21_X1 U12584 ( .B1(n6845), .B2(n7021), .A(n6846), .ZN(n6109) );
  INV_X1 U12585 ( .A(n6715), .ZN(n6610) );
  INV_X1 U12586 ( .A(n6712), .ZN(n6606) );
  NAND2_X1 U12587 ( .A1(n5796), .A2(n6114), .ZN(n6728) );
  AOI21_X1 U12588 ( .B1(n6728), .B2(n6115), .A(n6622), .ZN(n6118) );
  NAND2_X1 U12589 ( .A1(n6622), .A2(n6114), .ZN(n6116) );
  AOI21_X1 U12590 ( .B1(n6116), .B2(n6724), .A(n6722), .ZN(n6117) );
  NOR2_X1 U12591 ( .A1(n7768), .A2(n7527), .ZN(n6126) );
  INV_X1 U12592 ( .A(n6987), .ZN(n6991) );
  INV_X1 U12593 ( .A(n6119), .ZN(n6988) );
  INV_X1 U12594 ( .A(n6642), .ZN(n6120) );
  NAND2_X1 U12595 ( .A1(n6120), .A2(n6990), .ZN(n6125) );
  OAI21_X1 U12596 ( .B1(n6988), .B2(n6244), .A(n6841), .ZN(n6121) );
  INV_X1 U12597 ( .A(n6640), .ZN(n6838) );
  INV_X1 U12598 ( .A(n6989), .ZN(n6123) );
  INV_X1 U12600 ( .A(n24592), .ZN(n6128) );
  AOI21_X1 U12602 ( .B1(n6264), .B2(n6130), .A(n6531), .ZN(n6131) );
  AOI21_X1 U12603 ( .B1(n5916), .B2(n6543), .A(n6539), .ZN(n6135) );
  NAND2_X1 U12604 ( .A1(n6136), .A2(n6165), .ZN(n6540) );
  INV_X1 U12605 ( .A(n7384), .ZN(n7618) );
  OAI21_X1 U12606 ( .B1(n7385), .B2(n7618), .A(n7386), .ZN(n6152) );
  NAND2_X1 U12607 ( .A1(n6950), .A2(n25437), .ZN(n6138) );
  AND3_X1 U12608 ( .A1(n6139), .A2(n6528), .A3(n6138), .ZN(n6158) );
  INV_X1 U12609 ( .A(n6158), .ZN(n6140) );
  AND2_X1 U12610 ( .A1(n6540), .A2(n6140), .ZN(n6143) );
  NAND3_X1 U12611 ( .A1(n25437), .A2(n6948), .A3(n24994), .ZN(n6141) );
  INV_X1 U12612 ( .A(n6157), .ZN(n6142) );
  MUX2_X1 U12613 ( .A(n6145), .B(n6144), .S(n6281), .Z(n6149) );
  INV_X1 U12614 ( .A(n6146), .ZN(n6678) );
  NAND2_X1 U12615 ( .A1(n7385), .A2(n7619), .ZN(n6150) );
  NAND3_X1 U12616 ( .A1(n6152), .A2(n6151), .A3(n6150), .ZN(n6160) );
  NAND2_X1 U12617 ( .A1(n1509), .A2(n6156), .ZN(n6153) );
  NAND3_X1 U12618 ( .A1(n7622), .A2(n1895), .A3(n7386), .ZN(n6159) );
  XNOR2_X1 U12619 ( .A(n9194), .B(n8824), .ZN(n6161) );
  XNOR2_X1 U12620 ( .A(n8256), .B(n6161), .ZN(n6222) );
  OAI21_X1 U12621 ( .B1(n6164), .B2(n6539), .A(n5916), .ZN(n6166) );
  INV_X1 U12622 ( .A(n6165), .ZN(n6542) );
  INV_X1 U12623 ( .A(n7761), .ZN(n7307) );
  OAI22_X1 U12624 ( .A1(n6351), .A2(n6169), .B1(n6168), .B2(n6503), .ZN(n6172)
         );
  NAND2_X1 U12625 ( .A1(n6351), .A2(n6034), .ZN(n6170) );
  INV_X1 U12626 ( .A(n6497), .ZN(n6350) );
  INV_X1 U12627 ( .A(n7760), .ZN(n7305) );
  AOI21_X1 U12628 ( .B1(n6173), .B2(n6296), .A(n6438), .ZN(n6178) );
  NAND2_X1 U12629 ( .A1(n6297), .A2(n6438), .ZN(n6175) );
  AOI21_X1 U12630 ( .B1(n6176), .B2(n6175), .A(n6332), .ZN(n6177) );
  NAND2_X1 U12631 ( .A1(n6524), .A2(n944), .ZN(n6181) );
  NOR2_X1 U12632 ( .A1(n25427), .A2(n6455), .ZN(n6182) );
  OAI21_X1 U12633 ( .B1(n6183), .B2(n6182), .A(n6510), .ZN(n6186) );
  NAND2_X1 U12634 ( .A1(n6457), .A2(n6512), .ZN(n6338) );
  OAI211_X1 U12635 ( .C1(n25427), .C2(n6457), .A(n6338), .B(n6459), .ZN(n6185)
         );
  INV_X1 U12637 ( .A(n7647), .ZN(n6191) );
  NAND2_X1 U12638 ( .A1(n6187), .A2(n6452), .ZN(n6188) );
  NAND2_X1 U12639 ( .A1(n6449), .A2(n6447), .ZN(n6189) );
  NAND2_X1 U12640 ( .A1(n6191), .A2(n7651), .ZN(n6190) );
  NAND3_X1 U12641 ( .A1(n6191), .A2(n7651), .A3(n7760), .ZN(n6192) );
  OAI211_X1 U12642 ( .C1(n7307), .C2(n6194), .A(n6193), .B(n6192), .ZN(n9196)
         );
  OAI21_X1 U12643 ( .B1(n6344), .B2(n6444), .A(n6341), .ZN(n6197) );
  NAND2_X1 U12644 ( .A1(n25401), .A2(n6488), .ZN(n6785) );
  INV_X1 U12645 ( .A(n6493), .ZN(n6429) );
  NAND2_X1 U12646 ( .A1(n6489), .A2(n6490), .ZN(n6303) );
  INV_X1 U12647 ( .A(n6777), .ZN(n6925) );
  INV_X1 U12648 ( .A(n7294), .ZN(n7749) );
  NAND2_X1 U12649 ( .A1(n6915), .A2(n6918), .ZN(n6774) );
  INV_X1 U12650 ( .A(n6915), .ZN(n6910) );
  NAND2_X1 U12651 ( .A1(n6910), .A2(n24509), .ZN(n6201) );
  INV_X1 U12652 ( .A(n6912), .ZN(n6771) );
  NAND2_X1 U12653 ( .A1(n24037), .A2(n6771), .ZN(n6200) );
  NOR2_X1 U12654 ( .A1(n6910), .A2(n6771), .ZN(n6202) );
  NAND2_X1 U12655 ( .A1(n7749), .A2(n7537), .ZN(n6206) );
  INV_X1 U12657 ( .A(n6467), .ZN(n6326) );
  NAND2_X1 U12658 ( .A1(n6326), .A2(n6315), .ZN(n6204) );
  MUX2_X1 U12659 ( .A(n6204), .B(n6203), .S(n5451), .Z(n6205) );
  MUX2_X1 U12660 ( .A(n6207), .B(n6206), .S(n8014), .Z(n6215) );
  INV_X1 U12661 ( .A(n6208), .ZN(n6294) );
  NAND2_X1 U12662 ( .A1(n6294), .A2(n6438), .ZN(n6298) );
  NAND2_X1 U12663 ( .A1(n6298), .A2(n6335), .ZN(n6443) );
  INV_X1 U12665 ( .A(n6332), .ZN(n6295) );
  NAND3_X1 U12666 ( .A1(n6212), .A2(n6334), .A3(n6211), .ZN(n6213) );
  XNOR2_X1 U12667 ( .A(n8935), .B(n9196), .ZN(n8034) );
  INV_X1 U12668 ( .A(n7347), .ZN(n6216) );
  NAND2_X1 U12669 ( .A1(n6216), .A2(n7346), .ZN(n6217) );
  OAI21_X1 U12670 ( .B1(n8508), .B2(n7346), .A(n6217), .ZN(n6218) );
  XNOR2_X1 U12671 ( .A(n8341), .B(n1863), .ZN(n6220) );
  XNOR2_X1 U12672 ( .A(n8034), .B(n6220), .ZN(n6221) );
  INV_X1 U12673 ( .A(n7619), .ZN(n7617) );
  MUX2_X1 U12674 ( .A(n7617), .B(n7382), .S(n7615), .Z(n6224) );
  MUX2_X2 U12676 ( .A(n6224), .B(n6223), .S(n7380), .Z(n8333) );
  NAND3_X1 U12677 ( .A1(n6226), .A2(n6225), .A3(n6104), .ZN(n6229) );
  NAND3_X1 U12678 ( .A1(n7032), .A2(n7029), .A3(n7033), .ZN(n6228) );
  NAND2_X1 U12679 ( .A1(n6823), .A2(n6598), .ZN(n6829) );
  INV_X1 U12680 ( .A(n7013), .ZN(n6822) );
  NAND3_X1 U12681 ( .A1(n6829), .A2(n25044), .A3(n6230), .ZN(n6231) );
  NAND2_X1 U12682 ( .A1(n6234), .A2(n6233), .ZN(n6609) );
  INV_X1 U12683 ( .A(n6235), .ZN(n6718) );
  INV_X1 U12685 ( .A(n6238), .ZN(n6395) );
  INV_X1 U12686 ( .A(n6732), .ZN(n6397) );
  NAND3_X1 U12687 ( .A1(n6397), .A2(n6729), .A3(n6238), .ZN(n6241) );
  INV_X1 U12688 ( .A(n6396), .ZN(n6239) );
  NAND2_X1 U12689 ( .A1(n6733), .A2(n6239), .ZN(n6240) );
  INV_X1 U12690 ( .A(n6622), .ZN(n6727) );
  MUX2_X1 U12691 ( .A(n7732), .B(n7731), .S(n7733), .Z(n6250) );
  NAND2_X1 U12692 ( .A1(n6986), .A2(n6245), .ZN(n6246) );
  AOI21_X1 U12693 ( .B1(n6840), .B2(n6246), .A(n6640), .ZN(n6249) );
  AOI21_X1 U12694 ( .B1(n6247), .B2(n6988), .A(n6245), .ZN(n6248) );
  INV_X1 U12695 ( .A(n8806), .ZN(n6252) );
  XNOR2_X1 U12696 ( .A(n8333), .B(n6252), .ZN(n8398) );
  INV_X1 U12697 ( .A(n8398), .ZN(n6322) );
  NAND2_X1 U12698 ( .A1(n6253), .A2(n24994), .ZN(n6254) );
  NAND3_X1 U12699 ( .A1(n6255), .A2(n6947), .A3(n6529), .ZN(n6257) );
  NAND3_X1 U12700 ( .A1(n6952), .A2(n25437), .A3(n6528), .ZN(n6256) );
  NAND3_X1 U12702 ( .A1(n6530), .A2(n6531), .A3(n6538), .ZN(n6262) );
  OAI211_X1 U12703 ( .C1(n6264), .C2(n24067), .A(n6263), .B(n6262), .ZN(n6280)
         );
  NAND2_X1 U12704 ( .A1(n6164), .A2(n6266), .ZN(n6544) );
  NAND2_X1 U12705 ( .A1(n7103), .A2(n6539), .ZN(n6268) );
  NAND2_X1 U12706 ( .A1(n6544), .A2(n6268), .ZN(n6269) );
  MUX2_X1 U12708 ( .A(n7798), .B(n7802), .S(n7800), .Z(n6285) );
  INV_X1 U12709 ( .A(n6280), .ZN(n7432) );
  NAND2_X1 U12710 ( .A1(n6351), .A2(n441), .ZN(n6272) );
  MUX2_X1 U12711 ( .A(n6434), .B(n6272), .S(n6498), .Z(n6273) );
  NAND2_X1 U12712 ( .A1(n7432), .A2(n7803), .ZN(n7797) );
  AND2_X1 U12713 ( .A1(n440), .A2(n6274), .ZN(n6279) );
  NAND2_X1 U12714 ( .A1(n6275), .A2(n6521), .ZN(n6276) );
  NAND2_X1 U12715 ( .A1(n7797), .A2(n7053), .ZN(n6284) );
  AOI21_X1 U12717 ( .B1(n6945), .B2(n6943), .A(n6939), .ZN(n6283) );
  INV_X1 U12718 ( .A(n6770), .ZN(n6911) );
  AND2_X1 U12719 ( .A1(n6771), .A2(n6911), .ZN(n6289) );
  INV_X1 U12720 ( .A(n6918), .ZN(n6286) );
  NAND2_X1 U12722 ( .A1(n6909), .A2(n24037), .ZN(n6287) );
  OAI211_X2 U12723 ( .C1(n6289), .C2(n6774), .A(n6288), .B(n6287), .ZN(n7707)
         );
  INV_X1 U12724 ( .A(n7707), .ZN(n7867) );
  NAND2_X1 U12726 ( .A1(n6925), .A2(n6775), .ZN(n6291) );
  NAND2_X1 U12727 ( .A1(n6294), .A2(n6297), .ZN(n6336) );
  AOI21_X1 U12728 ( .B1(n6334), .B2(n6336), .A(n6295), .ZN(n6300) );
  INV_X1 U12729 ( .A(n6784), .ZN(n6487) );
  MUX2_X1 U12730 ( .A(n6303), .B(n6302), .S(n6493), .Z(n6307) );
  INV_X1 U12731 ( .A(n7863), .ZN(n7860) );
  INV_X1 U12732 ( .A(n6767), .ZN(n6309) );
  OAI21_X1 U12733 ( .B1(n6876), .B2(n6309), .A(n6875), .ZN(n6308) );
  NAND2_X1 U12734 ( .A1(n6308), .A2(n4922), .ZN(n6313) );
  NAND3_X1 U12735 ( .A1(n6310), .A2(n6874), .A3(n6309), .ZN(n6311) );
  NAND2_X1 U12736 ( .A1(n3570), .A2(n7861), .ZN(n6319) );
  NAND3_X1 U12737 ( .A1(n6315), .A2(n6329), .A3(n25404), .ZN(n6317) );
  NAND3_X1 U12738 ( .A1(n6326), .A2(n5451), .A3(n5966), .ZN(n6316) );
  XNOR2_X1 U12740 ( .A(n9155), .B(n25235), .ZN(n6321) );
  XNOR2_X1 U12741 ( .A(n6322), .B(n6321), .ZN(n6423) );
  AOI21_X1 U12742 ( .B1(n6519), .B2(n1509), .A(n6323), .ZN(n6325) );
  OAI21_X1 U12743 ( .B1(n6328), .B2(n5451), .A(n6327), .ZN(n6331) );
  NAND3_X1 U12744 ( .A1(n6440), .A2(n6209), .A3(n6438), .ZN(n6333) );
  OAI211_X1 U12745 ( .C1(n6336), .C2(n6335), .A(n6334), .B(n6333), .ZN(n7057)
         );
  INV_X1 U12746 ( .A(n6456), .ZN(n6339) );
  NAND3_X1 U12747 ( .A1(n25428), .A2(n6339), .A3(n6509), .ZN(n6340) );
  MUX2_X1 U12748 ( .A(n9066), .B(n7057), .S(n9067), .Z(n6355) );
  NAND2_X1 U12749 ( .A1(n6341), .A2(n6447), .ZN(n6343) );
  NAND2_X1 U12750 ( .A1(n6452), .A2(n6445), .ZN(n6342) );
  AND2_X1 U12751 ( .A1(n6343), .A2(n6342), .ZN(n6349) );
  INV_X1 U12752 ( .A(n6344), .ZN(n6346) );
  NOR2_X1 U12753 ( .A1(n7809), .A2(n8219), .ZN(n7814) );
  NAND2_X1 U12754 ( .A1(n6496), .A2(n6350), .ZN(n6353) );
  INV_X1 U12755 ( .A(n6351), .ZN(n6499) );
  NOR2_X1 U12757 ( .A1(n7813), .A2(n8219), .ZN(n7196) );
  INV_X1 U12758 ( .A(n9067), .ZN(n7738) );
  OAI22_X1 U12759 ( .A1(n7814), .A2(n7196), .B1(n7738), .B2(n7809), .ZN(n6354)
         );
  OAI21_X2 U12760 ( .B1(n6355), .B2(n7812), .A(n6354), .ZN(n8278) );
  NAND2_X1 U12761 ( .A1(n6818), .A2(n6893), .ZN(n6356) );
  AOI21_X1 U12762 ( .B1(n6357), .B2(n6356), .A(n6358), .ZN(n6361) );
  NAND3_X1 U12763 ( .A1(n6651), .A2(n6358), .A3(n6893), .ZN(n6360) );
  OR3_X1 U12764 ( .A1(n6819), .A2(n6895), .A3(n6893), .ZN(n6359) );
  NAND2_X1 U12765 ( .A1(n6793), .A2(n6078), .ZN(n6363) );
  INV_X1 U12766 ( .A(n6363), .ZN(n6366) );
  OAI21_X1 U12767 ( .B1(n6078), .B2(n6794), .A(n6882), .ZN(n6365) );
  MUX2_X1 U12768 ( .A(n6363), .B(n6362), .S(n6885), .Z(n6364) );
  OAI21_X1 U12771 ( .B1(n6072), .B2(n6369), .A(n6071), .ZN(n6370) );
  OAI21_X1 U12772 ( .B1(n6899), .B2(n6373), .A(n6377), .ZN(n6378) );
  OAI21_X1 U12774 ( .B1(n6848), .B2(n7021), .A(n6845), .ZN(n6380) );
  NAND2_X1 U12775 ( .A1(n7022), .A2(n7026), .ZN(n6379) );
  NAND3_X1 U12776 ( .A1(n7025), .A2(n250), .A3(n4643), .ZN(n6382) );
  AND2_X1 U12777 ( .A1(n6094), .A2(n7005), .ZN(n6387) );
  NAND2_X1 U12778 ( .A1(n6832), .A2(n7008), .ZN(n6386) );
  OAI21_X1 U12779 ( .B1(n6384), .B2(n7007), .A(n6383), .ZN(n6385) );
  XNOR2_X1 U12780 ( .A(n8278), .B(n8615), .ZN(n6421) );
  OAI21_X1 U12781 ( .B1(n6975), .B2(n1149), .A(n24395), .ZN(n6391) );
  AND2_X1 U12782 ( .A1(n1149), .A2(n6688), .ZN(n6389) );
  NAND2_X1 U12783 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  AOI21_X1 U12784 ( .B1(n6397), .B2(n6733), .A(n6396), .ZN(n6398) );
  NAND2_X1 U12785 ( .A1(n271), .A2(n6400), .ZN(n6403) );
  INV_X1 U12786 ( .A(n6400), .ZN(n6674) );
  NAND2_X1 U12787 ( .A1(n6674), .A2(n6757), .ZN(n6401) );
  NAND2_X1 U12788 ( .A1(n7563), .A2(n7721), .ZN(n7858) );
  NAND2_X1 U12789 ( .A1(n6965), .A2(n6963), .ZN(n6405) );
  NAND2_X1 U12790 ( .A1(n6964), .A2(n5800), .ZN(n6404) );
  OAI21_X1 U12791 ( .B1(n7184), .B2(n4752), .A(n6406), .ZN(n6413) );
  INV_X1 U12792 ( .A(n6630), .ZN(n6565) );
  INV_X1 U12793 ( .A(n6407), .ZN(n6746) );
  NAND2_X1 U12794 ( .A1(n453), .A2(n6407), .ZN(n6408) );
  INV_X1 U12795 ( .A(n7853), .ZN(n7564) );
  INV_X1 U12796 ( .A(n7563), .ZN(n7854) );
  INV_X1 U12797 ( .A(n6414), .ZN(n6698) );
  NAND2_X1 U12798 ( .A1(n6698), .A2(n6694), .ZN(n6558) );
  INV_X1 U12799 ( .A(n6697), .ZN(n6559) );
  NOR2_X1 U12800 ( .A1(n6695), .A2(n6559), .ZN(n6416) );
  NOR2_X1 U12801 ( .A1(n7857), .A2(n7721), .ZN(n7849) );
  NAND2_X1 U12802 ( .A1(n7849), .A2(n7563), .ZN(n6418) );
  OAI211_X1 U12803 ( .C1(n24072), .C2(n7858), .A(n6419), .B(n6418), .ZN(n8588)
         );
  XNOR2_X1 U12804 ( .A(n8588), .B(n1739), .ZN(n6420) );
  XNOR2_X1 U12805 ( .A(n6421), .B(n6420), .ZN(n6422) );
  XNOR2_X1 U12806 ( .A(n6423), .B(n6422), .ZN(n9462) );
  NAND2_X1 U12809 ( .A1(n6470), .A2(n6426), .ZN(n6469) );
  NAND2_X1 U12810 ( .A1(n25401), .A2(n6784), .ZN(n6494) );
  NAND2_X1 U12811 ( .A1(n6429), .A2(n6490), .ZN(n6428) );
  AOI21_X1 U12812 ( .B1(n6494), .B2(n6428), .A(n6301), .ZN(n6433) );
  NAND2_X1 U12813 ( .A1(n6429), .A2(n6489), .ZN(n6431) );
  AOI21_X1 U12814 ( .B1(n6431), .B2(n6430), .A(n6490), .ZN(n6432) );
  NAND2_X1 U12816 ( .A1(n6497), .A2(n6034), .ZN(n6501) );
  OAI21_X1 U12817 ( .B1(n6499), .B2(n6498), .A(n24466), .ZN(n6436) );
  NOR2_X1 U12818 ( .A1(n6438), .A2(n6209), .ZN(n6442) );
  NAND2_X1 U12819 ( .A1(n7085), .A2(n433), .ZN(n6466) );
  NAND3_X1 U12820 ( .A1(n6445), .A2(n6449), .A3(n6444), .ZN(n6446) );
  OAI21_X1 U12821 ( .B1(n6448), .B2(n6447), .A(n6446), .ZN(n7689) );
  NOR2_X1 U12823 ( .A1(n7689), .A2(n7691), .ZN(n7147) );
  INV_X1 U12824 ( .A(n7147), .ZN(n8317) );
  NOR2_X1 U12825 ( .A1(n8317), .A2(n8315), .ZN(n6465) );
  INV_X1 U12826 ( .A(n25428), .ZN(n6464) );
  NAND2_X1 U12827 ( .A1(n6454), .A2(n6510), .ZN(n6463) );
  NAND2_X1 U12828 ( .A1(n6456), .A2(n6455), .ZN(n6458) );
  OAI211_X1 U12829 ( .C1(n6455), .C2(n6464), .A(n6458), .B(n6457), .ZN(n6462)
         );
  NAND3_X1 U12830 ( .A1(n6460), .A2(n6459), .A3(n6509), .ZN(n6461) );
  INV_X1 U12833 ( .A(n9147), .ZN(n8152) );
  AOI21_X1 U12834 ( .B1(n6471), .B2(n6470), .A(n5966), .ZN(n6472) );
  NAND2_X1 U12835 ( .A1(n6372), .A2(n6473), .ZN(n6474) );
  NAND2_X1 U12836 ( .A1(n6477), .A2(n6876), .ZN(n6478) );
  AND2_X1 U12837 ( .A1(n6874), .A2(n6870), .ZN(n6879) );
  NOR2_X1 U12838 ( .A1(n6480), .A2(n6775), .ZN(n6479) );
  NAND2_X1 U12839 ( .A1(n6915), .A2(n24509), .ZN(n6769) );
  NAND2_X1 U12840 ( .A1(n24037), .A2(n6915), .ZN(n6483) );
  OAI211_X1 U12841 ( .C1(n6912), .C2(n24037), .A(n6483), .B(n6911), .ZN(n6484)
         );
  NAND2_X1 U12842 ( .A1(n7638), .A2(n7917), .ZN(n7635) );
  INV_X1 U12843 ( .A(n6489), .ZN(n6783) );
  NAND3_X1 U12844 ( .A1(n6490), .A2(n6783), .A3(n6493), .ZN(n6491) );
  XNOR2_X1 U12845 ( .A(n8152), .B(n8908), .ZN(n8050) );
  OR2_X1 U12846 ( .A1(n6497), .A2(n6496), .ZN(n6500) );
  INV_X1 U12848 ( .A(n6506), .ZN(n6508) );
  NAND2_X1 U12849 ( .A1(n6508), .A2(n6507), .ZN(n6516) );
  NAND2_X1 U12850 ( .A1(n6509), .A2(n6512), .ZN(n6511) );
  NAND2_X1 U12851 ( .A1(n6511), .A2(n6510), .ZN(n6515) );
  NOR2_X1 U12852 ( .A1(n25427), .A2(n6512), .ZN(n6514) );
  INV_X1 U12853 ( .A(n6806), .ZN(n8531) );
  NAND2_X1 U12854 ( .A1(n6519), .A2(n25398), .ZN(n6520) );
  NAND2_X1 U12855 ( .A1(n6524), .A2(n6523), .ZN(n6525) );
  NAND3_X1 U12856 ( .A1(n6947), .A2(n5903), .A3(n6950), .ZN(n6527) );
  OAI21_X1 U12857 ( .B1(n7087), .B2(n8531), .A(n6548), .ZN(n6860) );
  NAND2_X1 U12858 ( .A1(n6532), .A2(n6531), .ZN(n6536) );
  NAND2_X1 U12859 ( .A1(n24254), .A2(n6538), .ZN(n6535) );
  MUX2_X1 U12860 ( .A(n6536), .B(n6535), .S(n24067), .Z(n6537) );
  MUX2_X1 U12861 ( .A(n6540), .B(n7098), .S(n6539), .Z(n6547) );
  MUX2_X1 U12862 ( .A(n6545), .B(n6544), .S(n6543), .Z(n6546) );
  OAI211_X1 U12863 ( .C1(n8531), .C2(n7663), .A(n6549), .B(n6548), .ZN(n6550)
         );
  NAND2_X1 U12867 ( .A1(n6553), .A2(n5924), .ZN(n6555) );
  NAND3_X1 U12868 ( .A1(n3923), .A2(n6702), .A3(n6959), .ZN(n6554) );
  INV_X1 U12870 ( .A(n6933), .ZN(n6557) );
  NAND2_X1 U12871 ( .A1(n6557), .A2(n6556), .ZN(n6563) );
  INV_X1 U12872 ( .A(n6558), .ZN(n6937) );
  NAND2_X1 U12873 ( .A1(n6560), .A2(n2008), .ZN(n6561) );
  NAND2_X1 U12874 ( .A1(n7445), .A2(n7444), .ZN(n7262) );
  NAND2_X1 U12875 ( .A1(n6746), .A2(n453), .ZN(n6564) );
  AOI21_X1 U12876 ( .B1(n6748), .B2(n6564), .A(n6744), .ZN(n7928) );
  NAND2_X1 U12877 ( .A1(n6565), .A2(n453), .ZN(n6566) );
  OR2_X1 U12878 ( .A1(n7262), .A2(n5607), .ZN(n6586) );
  AOI21_X1 U12879 ( .B1(n24579), .B2(n6688), .A(n6687), .ZN(n6974) );
  OAI211_X1 U12880 ( .C1(n6977), .C2(n6568), .A(n6567), .B(n24395), .ZN(n6569)
         );
  NAND3_X1 U12881 ( .A1(n6572), .A2(n6969), .A3(n6571), .ZN(n6574) );
  NAND3_X1 U12882 ( .A1(n4754), .A2(n6964), .A3(n5800), .ZN(n6573) );
  OAI211_X2 U12883 ( .C1(n6576), .C2(n6575), .A(n6574), .B(n6573), .ZN(n7932)
         );
  NOR2_X1 U12884 ( .A1(n7444), .A2(n7932), .ZN(n6583) );
  NAND2_X1 U12885 ( .A1(n6583), .A2(n5607), .ZN(n6585) );
  INV_X1 U12886 ( .A(n6577), .ZN(n6758) );
  NAND2_X1 U12887 ( .A1(n6675), .A2(n6758), .ZN(n6580) );
  INV_X1 U12888 ( .A(n6757), .ZN(n6673) );
  MUX2_X1 U12889 ( .A(n6580), .B(n6579), .S(n6578), .Z(n6581) );
  NAND2_X1 U12890 ( .A1(n6583), .A2(n7924), .ZN(n6584) );
  XNOR2_X1 U12891 ( .A(n8484), .B(n8634), .ZN(n6587) );
  XNOR2_X1 U12892 ( .A(n8050), .B(n6587), .ZN(n6666) );
  INV_X1 U12893 ( .A(n7035), .ZN(n6739) );
  NAND2_X1 U12894 ( .A1(n6588), .A2(n7032), .ZN(n6590) );
  MUX2_X1 U12895 ( .A(n6591), .B(n6590), .S(n25424), .Z(n6595) );
  INV_X1 U12896 ( .A(n7032), .ZN(n6592) );
  NAND2_X1 U12898 ( .A1(n6597), .A2(n25045), .ZN(n6605) );
  NAND2_X1 U12901 ( .A1(n24090), .A2(n6822), .ZN(n6604) );
  NAND2_X1 U12902 ( .A1(n25044), .A2(n6601), .ZN(n6603) );
  INV_X1 U12903 ( .A(n6609), .ZN(n6612) );
  NAND2_X1 U12904 ( .A1(n6393), .A2(n6615), .ZN(n6616) );
  INV_X1 U12905 ( .A(n7787), .ZN(n6618) );
  NAND2_X1 U12906 ( .A1(n6619), .A2(n6722), .ZN(n6620) );
  AOI21_X1 U12907 ( .B1(n6621), .B2(n6620), .A(n6723), .ZN(n6627) );
  NAND2_X1 U12908 ( .A1(n6622), .A2(n5796), .ZN(n6625) );
  AOI21_X1 U12909 ( .B1(n6625), .B2(n6624), .A(n6114), .ZN(n6626) );
  INV_X1 U12910 ( .A(n7789), .ZN(n7783) );
  NAND2_X1 U12911 ( .A1(n6629), .A2(n6628), .ZN(n6632) );
  AND2_X1 U12912 ( .A1(n6630), .A2(n4696), .ZN(n6631) );
  AOI22_X1 U12913 ( .A1(n7783), .A2(n7418), .B1(n7787), .B2(n7788), .ZN(n7045)
         );
  NAND2_X1 U12916 ( .A1(n7025), .A2(n250), .ZN(n6637) );
  NAND2_X1 U12917 ( .A1(n442), .A2(n4643), .ZN(n6636) );
  INV_X1 U12918 ( .A(n7908), .ZN(n7450) );
  NAND2_X1 U12919 ( .A1(n7450), .A2(n7629), .ZN(n7626) );
  OAI21_X1 U12920 ( .B1(n6794), .B2(n6792), .A(n6643), .ZN(n6889) );
  NAND2_X1 U12921 ( .A1(n6889), .A2(n6795), .ZN(n6646) );
  AOI21_X1 U12922 ( .B1(n6793), .B2(n6644), .A(n6792), .ZN(n6645) );
  NAND2_X1 U12923 ( .A1(n6648), .A2(n7008), .ZN(n6649) );
  MUX2_X1 U12924 ( .A(n6895), .B(n6818), .S(n6890), .Z(n6656) );
  NAND2_X1 U12925 ( .A1(n6819), .A2(n6895), .ZN(n6654) );
  INV_X1 U12926 ( .A(n6893), .ZN(n6652) );
  MUX2_X1 U12927 ( .A(n6654), .B(n6653), .S(n6652), .Z(n6655) );
  OAI21_X1 U12928 ( .B1(n6656), .B2(n313), .A(n6655), .ZN(n7909) );
  NAND3_X1 U12929 ( .A1(n6658), .A2(n6997), .A3(n439), .ZN(n6659) );
  XNOR2_X1 U12930 ( .A(n8635), .B(n8699), .ZN(n6664) );
  INV_X1 U12931 ( .A(n7801), .ZN(n7799) );
  NAND3_X1 U12932 ( .A1(n7799), .A2(n7803), .A3(n7166), .ZN(n6662) );
  INV_X1 U12933 ( .A(n7166), .ZN(n7794) );
  OAI211_X1 U12934 ( .C1(n7801), .C2(n7798), .A(n7432), .B(n7794), .ZN(n6661)
         );
  NAND2_X1 U12935 ( .A1(n7800), .A2(n7801), .ZN(n6660) );
  NAND3_X1 U12936 ( .A1(n6662), .A2(n6661), .A3(n6660), .ZN(n8361) );
  XNOR2_X1 U12937 ( .A(n8361), .B(n447), .ZN(n6663) );
  XNOR2_X1 U12938 ( .A(n6664), .B(n6663), .ZN(n6665) );
  XNOR2_X1 U12939 ( .A(n6666), .B(n6665), .ZN(n9463) );
  NAND2_X1 U12940 ( .A1(n24944), .A2(n9463), .ZN(n9921) );
  INV_X1 U12941 ( .A(n6964), .ZN(n6668) );
  OAI21_X1 U12942 ( .B1(n6668), .B2(n6963), .A(n24089), .ZN(n6671) );
  NAND2_X1 U12943 ( .A1(n443), .A2(n6969), .ZN(n6669) );
  AOI22_X1 U12944 ( .A1(n6673), .A2(n6675), .B1(n6758), .B2(n6674), .ZN(n6677)
         );
  NAND3_X1 U12945 ( .A1(n6680), .A2(n6679), .A3(n6939), .ZN(n6681) );
  AND2_X1 U12946 ( .A1(n7414), .A2(n7415), .ZN(n6711) );
  NAND3_X1 U12947 ( .A1(n6688), .A2(n6975), .A3(n6687), .ZN(n6689) );
  INV_X1 U12948 ( .A(n7413), .ZN(n7998) );
  NAND2_X1 U12949 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  AND2_X1 U12950 ( .A1(n6696), .A2(n6935), .ZN(n6701) );
  OAI21_X1 U12951 ( .B1(n6699), .B2(n6698), .A(n6936), .ZN(n6700) );
  NAND2_X1 U12954 ( .A1(n6960), .A2(n24405), .ZN(n6707) );
  NAND3_X1 U12955 ( .A1(n3923), .A2(n5924), .A3(n6705), .ZN(n6706) );
  NAND3_X1 U12956 ( .A1(n6708), .A2(n6707), .A3(n6706), .ZN(n7412) );
  INV_X1 U12957 ( .A(n7412), .ZN(n7990) );
  NOR2_X1 U12958 ( .A1(n7413), .A2(n7990), .ZN(n6709) );
  OAI21_X1 U12959 ( .B1(n7498), .B2(n6709), .A(n7357), .ZN(n6710) );
  INV_X1 U12960 ( .A(n8846), .ZN(n8576) );
  NOR2_X1 U12961 ( .A1(n24501), .A2(n6714), .ZN(n6716) );
  NAND3_X1 U12962 ( .A1(n6724), .A2(n6723), .A3(n6722), .ZN(n6725) );
  NAND2_X1 U12963 ( .A1(n6869), .A2(n25251), .ZN(n6743) );
  INV_X1 U12964 ( .A(n6868), .ZN(n6738) );
  NAND2_X1 U12965 ( .A1(n6733), .A2(n6732), .ZN(n6735) );
  INV_X1 U12966 ( .A(n6867), .ZN(n6737) );
  NAND4_X1 U12967 ( .A1(n7506), .A2(n6738), .A3(n1379), .A4(n6737), .ZN(n7672)
         );
  AOI21_X1 U12968 ( .B1(n7030), .B2(n454), .A(n7032), .ZN(n6742) );
  AOI21_X1 U12969 ( .B1(n6743), .B2(n7672), .A(n7676), .ZN(n6761) );
  INV_X1 U12970 ( .A(n25251), .ZN(n7677) );
  AND2_X1 U12971 ( .A1(n6744), .A2(n6051), .ZN(n6749) );
  NAND2_X1 U12972 ( .A1(n7677), .A2(n7674), .ZN(n6759) );
  OAI22_X1 U12973 ( .A1(n6869), .A2(n6759), .B1(n7677), .B2(n3275), .ZN(n6760)
         );
  NAND2_X1 U12975 ( .A1(n7591), .A2(n7590), .ZN(n7337) );
  OAI21_X1 U12976 ( .B1(n7464), .B2(n7592), .A(n7462), .ZN(n6762) );
  OAI21_X1 U12977 ( .B1(n6876), .B2(n6875), .A(n6874), .ZN(n6766) );
  NAND3_X1 U12978 ( .A1(n6768), .A2(n4922), .A3(n6870), .ZN(n6765) );
  INV_X1 U12979 ( .A(n6769), .ZN(n6773) );
  NAND3_X1 U12980 ( .A1(n6292), .A2(n6290), .A3(n6777), .ZN(n6778) );
  AOI21_X1 U12981 ( .B1(n6785), .B2(n6784), .A(n6783), .ZN(n6786) );
  INV_X1 U12982 ( .A(n7977), .ZN(n7820) );
  INV_X1 U12984 ( .A(n7975), .ZN(n7816) );
  NAND3_X1 U12985 ( .A1(n7973), .A2(n7972), .A3(n7816), .ZN(n6799) );
  NAND2_X1 U12986 ( .A1(n6793), .A2(n6795), .ZN(n6791) );
  NAND2_X1 U12987 ( .A1(n6793), .A2(n6792), .ZN(n6797) );
  OAI21_X1 U12988 ( .B1(n6795), .B2(n6794), .A(n6075), .ZN(n6796) );
  AOI22_X1 U12989 ( .A1(n6798), .A2(n6881), .B1(n6797), .B2(n6796), .ZN(n7976)
         );
  INV_X1 U12990 ( .A(n7976), .ZN(n7819) );
  NAND2_X1 U12991 ( .A1(n7819), .A2(n7974), .ZN(n7821) );
  XNOR2_X1 U12992 ( .A(n8913), .B(n9140), .ZN(n6800) );
  XNOR2_X1 U12993 ( .A(n8628), .B(n6800), .ZN(n6859) );
  AOI22_X1 U12995 ( .A1(n7598), .A2(n7600), .B1(n25037), .B2(n7257), .ZN(n6804) );
  NAND3_X1 U12996 ( .A1(n7597), .A2(n7600), .A3(n7602), .ZN(n6801) );
  AND2_X1 U12997 ( .A1(n6802), .A2(n6801), .ZN(n6803) );
  OAI21_X2 U12998 ( .B1(n6804), .B2(n7597), .A(n6803), .ZN(n9141) );
  XNOR2_X1 U12999 ( .A(n9141), .B(n2318), .ZN(n6857) );
  NAND2_X1 U13000 ( .A1(n7665), .A2(n8527), .ZN(n6809) );
  NAND2_X1 U13001 ( .A1(n6805), .A2(n7667), .ZN(n6808) );
  NAND2_X1 U13002 ( .A1(n7664), .A2(n8528), .ZN(n6807) );
  NAND2_X1 U13003 ( .A1(n6999), .A2(n6072), .ZN(n6814) );
  NAND2_X1 U13006 ( .A1(n6818), .A2(n6895), .ZN(n6820) );
  AOI21_X1 U13007 ( .B1(n6820), .B2(n6819), .A(n313), .ZN(n6821) );
  INV_X1 U13008 ( .A(n7985), .ZN(n7828) );
  NAND2_X1 U13009 ( .A1(n6823), .A2(n6822), .ZN(n6825) );
  AOI21_X1 U13010 ( .B1(n6826), .B2(n6825), .A(n6824), .ZN(n6831) );
  INV_X1 U13011 ( .A(n7984), .ZN(n7825) );
  MUX2_X1 U13012 ( .A(n6834), .B(n6833), .S(n7011), .Z(n6837) );
  AND2_X1 U13013 ( .A1(n7009), .A2(n7008), .ZN(n6835) );
  OAI21_X1 U13014 ( .B1(n6840), .B2(n6986), .A(n6839), .ZN(n6844) );
  NAND2_X1 U13015 ( .A1(n6244), .A2(n6987), .ZN(n6842) );
  AOI21_X1 U13016 ( .B1(n6842), .B2(n6841), .A(n6990), .ZN(n6843) );
  NOR2_X1 U13017 ( .A1(n6844), .A2(n6843), .ZN(n7409) );
  INV_X1 U13018 ( .A(n7409), .ZN(n7046) );
  NAND3_X1 U13019 ( .A1(n7989), .A2(n7048), .A3(n7046), .ZN(n6853) );
  NAND2_X1 U13020 ( .A1(n6846), .A2(n6845), .ZN(n6847) );
  OAI211_X1 U13021 ( .C1(n7027), .C2(n7021), .A(n6847), .B(n7025), .ZN(n6851)
         );
  OAI211_X1 U13022 ( .C1(n250), .C2(n7027), .A(n7028), .B(n442), .ZN(n6850) );
  XNOR2_X1 U13023 ( .A(n8353), .B(n8687), .ZN(n6856) );
  XNOR2_X1 U13024 ( .A(n6857), .B(n6856), .ZN(n6858) );
  XNOR2_X1 U13025 ( .A(n6859), .B(n6858), .ZN(n9459) );
  NAND2_X1 U13026 ( .A1(n9461), .A2(n9459), .ZN(n9913) );
  NAND2_X1 U13027 ( .A1(n9921), .A2(n9913), .ZN(n7043) );
  NAND2_X1 U13028 ( .A1(n6860), .A2(n7664), .ZN(n6863) );
  NOR2_X1 U13029 ( .A1(n7087), .A2(n7662), .ZN(n6861) );
  AOI22_X1 U13030 ( .A1(n6861), .A2(n8530), .B1(n269), .B2(n8531), .ZN(n6862)
         );
  AOI21_X1 U13031 ( .B1(n8317), .B2(n8315), .A(n8314), .ZN(n6866) );
  XNOR2_X1 U13032 ( .A(n8987), .B(n9167), .ZN(n8058) );
  NAND2_X1 U13033 ( .A1(n6871), .A2(n6870), .ZN(n6872) );
  AND2_X1 U13034 ( .A1(n6873), .A2(n6872), .ZN(n6880) );
  NAND2_X1 U13035 ( .A1(n6875), .A2(n6874), .ZN(n6877) );
  NAND2_X1 U13036 ( .A1(n6882), .A2(n6881), .ZN(n6888) );
  INV_X1 U13037 ( .A(n6883), .ZN(n6887) );
  NAND2_X1 U13038 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  NAND2_X1 U13039 ( .A1(n6895), .A2(n6890), .ZN(n6891) );
  NAND2_X1 U13040 ( .A1(n6892), .A2(n6891), .ZN(n6898) );
  NOR2_X1 U13041 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  AOI21_X2 U13042 ( .B1(n6897), .B2(n6898), .A(n6896), .ZN(n7657) );
  INV_X1 U13043 ( .A(n6899), .ZN(n6901) );
  NAND2_X1 U13044 ( .A1(n6901), .A2(n6900), .ZN(n6908) );
  OAI21_X1 U13045 ( .B1(n6905), .B2(n6904), .A(n6903), .ZN(n6907) );
  MUX2_X2 U13046 ( .A(n6908), .B(n6907), .S(n6906), .Z(n7943) );
  NAND3_X1 U13047 ( .A1(n6910), .A2(n6909), .A3(n6916), .ZN(n6914) );
  NAND3_X1 U13048 ( .A1(n6912), .A2(n24037), .A3(n6911), .ZN(n6913) );
  NAND2_X1 U13049 ( .A1(n6916), .A2(n6915), .ZN(n6921) );
  NAND2_X1 U13050 ( .A1(n6918), .A2(n24509), .ZN(n6920) );
  NAND3_X1 U13051 ( .A1(n7945), .A2(n7657), .A3(n7942), .ZN(n6930) );
  AOI21_X1 U13052 ( .B1(n6926), .B2(n6925), .A(n6924), .ZN(n6927) );
  INV_X1 U13055 ( .A(n6938), .ZN(n6942) );
  NAND2_X1 U13056 ( .A1(n6940), .A2(n6939), .ZN(n6941) );
  NAND3_X1 U13057 ( .A1(n6950), .A2(n6949), .A3(n6948), .ZN(n6951) );
  OAI21_X1 U13058 ( .B1(n6956), .B2(n24257), .A(n6954), .ZN(n6962) );
  OAI21_X1 U13059 ( .B1(n3923), .B2(n6959), .A(n6958), .ZN(n6961) );
  INV_X1 U13060 ( .A(n6963), .ZN(n6966) );
  AOI21_X1 U13061 ( .B1(n6966), .B2(n6965), .A(n6964), .ZN(n6970) );
  NAND2_X1 U13062 ( .A1(n6967), .A2(n443), .ZN(n6968) );
  NOR2_X1 U13064 ( .A1(n6971), .A2(n6977), .ZN(n6973) );
  OAI21_X1 U13065 ( .B1(n6973), .B2(n6974), .A(n24579), .ZN(n6981) );
  NAND2_X1 U13066 ( .A1(n6976), .A2(n24395), .ZN(n6978) );
  MUX2_X1 U13067 ( .A(n6979), .B(n6978), .S(n6977), .Z(n6980) );
  INV_X1 U13068 ( .A(n7897), .ZN(n6985) );
  NAND2_X1 U13069 ( .A1(n6982), .A2(n7232), .ZN(n6983) );
  NAND2_X1 U13070 ( .A1(n6983), .A2(n24861), .ZN(n6984) );
  XNOR2_X1 U13071 ( .A(n8499), .B(n8088), .ZN(n7040) );
  OAI21_X1 U13072 ( .B1(n6838), .B2(n6986), .A(n6989), .ZN(n6995) );
  AOI21_X1 U13073 ( .B1(n6988), .B2(n6987), .A(n6990), .ZN(n6994) );
  OAI21_X1 U13074 ( .B1(n6244), .B2(n6990), .A(n6989), .ZN(n6992) );
  NAND2_X1 U13075 ( .A1(n6992), .A2(n6991), .ZN(n6993) );
  INV_X1 U13076 ( .A(n7961), .ZN(n7070) );
  OAI21_X1 U13077 ( .B1(n6368), .B2(n6996), .A(n6367), .ZN(n6998) );
  NAND2_X1 U13078 ( .A1(n6998), .A2(n7002), .ZN(n7001) );
  NAND2_X1 U13079 ( .A1(n7070), .A2(n7962), .ZN(n7069) );
  OAI21_X1 U13080 ( .B1(n7009), .B2(n7008), .A(n7007), .ZN(n7010) );
  NAND2_X1 U13081 ( .A1(n5992), .A2(n7013), .ZN(n7016) );
  OAI21_X1 U13082 ( .B1(n7033), .B2(n7035), .A(n7032), .ZN(n7034) );
  NAND2_X1 U13083 ( .A1(n7036), .A2(n7961), .ZN(n7038) );
  AND2_X1 U13084 ( .A1(n7234), .A2(n7965), .ZN(n7960) );
  NAND2_X1 U13085 ( .A1(n7960), .A2(n7683), .ZN(n7037) );
  OAI211_X2 U13086 ( .C1(n7069), .C2(n7235), .A(n7038), .B(n7037), .ZN(n8813)
         );
  XNOR2_X1 U13087 ( .A(n8813), .B(n2772), .ZN(n7039) );
  XNOR2_X1 U13088 ( .A(n7040), .B(n7039), .ZN(n7041) );
  AOI21_X1 U13089 ( .B1(n7046), .B2(n7826), .A(n7825), .ZN(n7047) );
  XNOR2_X1 U13090 ( .A(n8812), .B(n24056), .ZN(n8459) );
  AOI21_X1 U13091 ( .B1(n7517), .B2(n7516), .A(n7972), .ZN(n7051) );
  NAND2_X1 U13092 ( .A1(n7816), .A2(n7974), .ZN(n7049) );
  XNOR2_X1 U13093 ( .A(n8764), .B(n8406), .ZN(n7052) );
  XNOR2_X1 U13094 ( .A(n8459), .B(n7052), .ZN(n7063) );
  INV_X1 U13095 ( .A(n7800), .ZN(n7054) );
  NAND2_X1 U13096 ( .A1(n7801), .A2(n7798), .ZN(n7434) );
  INV_X1 U13097 ( .A(n3118), .ZN(n23448) );
  XNOR2_X1 U13098 ( .A(n8896), .B(n23448), .ZN(n7061) );
  AND2_X1 U13099 ( .A1(n7412), .A2(n7358), .ZN(n7499) );
  AOI22_X1 U13100 ( .A1(n7499), .A2(n7991), .B1(n7992), .B2(n7415), .ZN(n7056)
         );
  NAND3_X1 U13101 ( .A1(n7992), .A2(n7413), .A3(n7412), .ZN(n7055) );
  OAI211_X1 U13102 ( .C1(n7414), .C2(n7992), .A(n7056), .B(n7055), .ZN(n8285)
         );
  NAND2_X1 U13103 ( .A1(n7813), .A2(n8219), .ZN(n7059) );
  NAND3_X1 U13104 ( .A1(n7813), .A2(n9068), .A3(n9066), .ZN(n7058) );
  XNOR2_X1 U13105 ( .A(n8285), .B(n9044), .ZN(n7060) );
  XNOR2_X1 U13106 ( .A(n7061), .B(n7060), .ZN(n7062) );
  INV_X1 U13107 ( .A(n7183), .ZN(n9951) );
  NOR2_X1 U13108 ( .A1(n7421), .A2(n7474), .ZN(n7064) );
  NAND2_X1 U13109 ( .A1(n7423), .A2(n7477), .ZN(n7067) );
  MUX2_X1 U13110 ( .A(n7067), .B(n7066), .S(n7476), .Z(n7068) );
  OAI211_X1 U13111 ( .C1(n7071), .C2(n7070), .A(n7485), .B(n7069), .ZN(n7072)
         );
  OR2_X1 U13112 ( .A1(n7078), .A2(n7674), .ZN(n7076) );
  OAI21_X1 U13113 ( .B1(n7076), .B2(n7224), .A(n7075), .ZN(n7077) );
  NAND3_X1 U13114 ( .A1(n434), .A2(n7677), .A3(n7078), .ZN(n7079) );
  INV_X1 U13115 ( .A(n8452), .ZN(n8820) );
  INV_X1 U13116 ( .A(n7947), .ZN(n7946) );
  NAND2_X1 U13117 ( .A1(n7946), .A2(n7942), .ZN(n7081) );
  NOR2_X1 U13118 ( .A1(n7945), .A2(n7657), .ZN(n7080) );
  XNOR2_X1 U13119 ( .A(n8820), .B(n8787), .ZN(n7082) );
  XNOR2_X1 U13120 ( .A(n7083), .B(n7082), .ZN(n7095) );
  NAND2_X1 U13121 ( .A1(n8317), .A2(n8316), .ZN(n7149) );
  NAND2_X1 U13122 ( .A1(n8315), .A2(n8314), .ZN(n7084) );
  NAND3_X1 U13123 ( .A1(n7149), .A2(n7085), .A3(n7084), .ZN(n7086) );
  OAI211_X1 U13124 ( .C1(n7149), .C2(n7217), .A(n7086), .B(n8319), .ZN(n9073)
         );
  NAND3_X1 U13125 ( .A1(n8530), .A2(n7667), .A3(n8528), .ZN(n7091) );
  NAND3_X1 U13126 ( .A1(n7665), .A2(n7667), .A3(n269), .ZN(n7090) );
  NAND3_X1 U13128 ( .A1(n7664), .A2(n7666), .A3(n7662), .ZN(n7088) );
  NAND4_X2 U13129 ( .A1(n7088), .A2(n7091), .A3(n7090), .A4(n7089), .ZN(n8651)
         );
  XNOR2_X1 U13130 ( .A(n9073), .B(n8651), .ZN(n7093) );
  INV_X1 U13131 ( .A(n21204), .ZN(n22150) );
  XNOR2_X1 U13132 ( .A(n8412), .B(n22150), .ZN(n7092) );
  XNOR2_X1 U13133 ( .A(n7093), .B(n7092), .ZN(n7094) );
  XNOR2_X1 U13134 ( .A(n7095), .B(n7094), .ZN(n9950) );
  NAND2_X1 U13135 ( .A1(n9951), .A2(n9950), .ZN(n9387) );
  NOR2_X1 U13137 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  NAND4_X1 U13138 ( .A1(n7105), .A2(n7347), .A3(n7349), .A4(n7104), .ZN(n7106)
         );
  XNOR2_X1 U13139 ( .A(n8333), .B(n8280), .ZN(n7113) );
  NAND2_X1 U13140 ( .A1(n7526), .A2(n7771), .ZN(n7110) );
  NAND2_X1 U13141 ( .A1(n7284), .A2(n7527), .ZN(n7109) );
  INV_X1 U13142 ( .A(n7768), .ZN(n7288) );
  MUX2_X1 U13143 ( .A(n7110), .B(n7109), .S(n7288), .Z(n7112) );
  AOI22_X1 U13145 ( .A1(n7522), .A2(n23), .B1(n7525), .B2(n7767), .ZN(n7111)
         );
  XNOR2_X1 U13147 ( .A(n8891), .B(n8807), .ZN(n8444) );
  XNOR2_X1 U13148 ( .A(n8444), .B(n7113), .ZN(n7120) );
  NAND2_X1 U13149 ( .A1(n7754), .A2(n7292), .ZN(n8006) );
  NAND2_X1 U13150 ( .A1(n7760), .A2(n7651), .ZN(n7115) );
  NOR2_X1 U13151 ( .A1(n7761), .A2(n7646), .ZN(n7116) );
  OAI21_X1 U13152 ( .B1(n7391), .B2(n7116), .A(n7305), .ZN(n7117) );
  XNOR2_X1 U13153 ( .A(n8400), .B(n923), .ZN(n7118) );
  XNOR2_X1 U13154 ( .A(n25020), .B(n7118), .ZN(n7119) );
  OAI21_X1 U13155 ( .B1(n7592), .B2(n7590), .A(n268), .ZN(n7122) );
  NAND3_X1 U13156 ( .A1(n7462), .A2(n2035), .A3(n5971), .ZN(n7121) );
  INV_X1 U13157 ( .A(n7882), .ZN(n7126) );
  INV_X1 U13159 ( .A(n7313), .ZN(n7123) );
  INV_X1 U13160 ( .A(n7585), .ZN(n7125) );
  NAND3_X1 U13161 ( .A1(n7126), .A2(n7125), .A3(n7582), .ZN(n7127) );
  INV_X1 U13162 ( .A(n7604), .ZN(n7128) );
  NOR2_X1 U13163 ( .A1(n7604), .A2(n7323), .ZN(n7129) );
  INV_X1 U13164 ( .A(n7579), .ZN(n7318) );
  NAND2_X1 U13165 ( .A1(n7577), .A2(n7318), .ZN(n7320) );
  NAND3_X1 U13166 ( .A1(n7577), .A2(n4136), .A3(n7576), .ZN(n7130) );
  NAND2_X1 U13169 ( .A1(n7600), .A2(n7597), .ZN(n7132) );
  NAND2_X1 U13171 ( .A1(n7596), .A2(n7255), .ZN(n7133) );
  NAND3_X1 U13172 ( .A1(n25037), .A2(n24772), .A3(n7135), .ZN(n7138) );
  NAND3_X1 U13173 ( .A1(n7255), .A2(n7600), .A3(n7257), .ZN(n7137) );
  XNOR2_X1 U13174 ( .A(n8647), .B(n8341), .ZN(n8387) );
  NAND2_X1 U13175 ( .A1(n248), .A2(n7230), .ZN(n7139) );
  NAND2_X1 U13176 ( .A1(n7140), .A2(n24861), .ZN(n7142) );
  NOR2_X1 U13177 ( .A1(n7230), .A2(n7232), .ZN(n7141) );
  INV_X1 U13178 ( .A(n8168), .ZN(n8270) );
  XNOR2_X1 U13179 ( .A(n8270), .B(n3089), .ZN(n7144) );
  XNOR2_X1 U13180 ( .A(n8387), .B(n7144), .ZN(n7145) );
  XNOR2_X1 U13181 ( .A(n7146), .B(n7145), .ZN(n9134) );
  INV_X1 U13182 ( .A(n9134), .ZN(n9389) );
  NAND3_X1 U13183 ( .A1(n7699), .A2(n7688), .A3(n8315), .ZN(n7150) );
  XNOR2_X1 U13186 ( .A(n24547), .B(n8353), .ZN(n8421) );
  INV_X1 U13187 ( .A(n7909), .ZN(n7625) );
  NAND2_X1 U13188 ( .A1(n7625), .A2(n7628), .ZN(n7154) );
  NAND2_X1 U13189 ( .A1(n7365), .A2(n7909), .ZN(n7153) );
  NAND3_X1 U13190 ( .A1(n7154), .A2(n7153), .A3(n7364), .ZN(n7158) );
  XNOR2_X1 U13194 ( .A(n7161), .B(n9082), .ZN(n8689) );
  INV_X1 U13195 ( .A(n8689), .ZN(n7162) );
  XNOR2_X1 U13196 ( .A(n7162), .B(n8421), .ZN(n7182) );
  NOR2_X1 U13197 ( .A1(n7163), .A2(n7932), .ZN(n7164) );
  INV_X1 U13198 ( .A(n7924), .ZN(n7261) );
  AOI22_X1 U13199 ( .A1(n7164), .A2(n7261), .B1(n7445), .B2(n7932), .ZN(n7165)
         );
  NAND2_X1 U13200 ( .A1(n7167), .A2(n7801), .ZN(n7169) );
  OAI21_X1 U13201 ( .B1(n7169), .B2(n7800), .A(n7168), .ZN(n7171) );
  AOI21_X1 U13202 ( .B1(n7434), .B2(n7795), .A(n7432), .ZN(n7170) );
  OR2_X1 U13203 ( .A1(n7171), .A2(n7170), .ZN(n8237) );
  XNOR2_X1 U13204 ( .A(n8428), .B(n8237), .ZN(n7180) );
  NAND2_X1 U13205 ( .A1(n7782), .A2(n7418), .ZN(n7172) );
  NAND2_X1 U13206 ( .A1(n7172), .A2(n2620), .ZN(n7173) );
  NAND2_X1 U13207 ( .A1(n7173), .A2(n7781), .ZN(n7178) );
  NAND3_X1 U13208 ( .A1(n7419), .A2(n7174), .A3(n7787), .ZN(n7177) );
  XNOR2_X1 U13209 ( .A(n8917), .B(n2120), .ZN(n7179) );
  XNOR2_X1 U13210 ( .A(n7180), .B(n7179), .ZN(n7181) );
  XNOR2_X1 U13211 ( .A(n7182), .B(n7181), .ZN(n9269) );
  OR2_X1 U13212 ( .A1(n9133), .A2(n9951), .ZN(n7210) );
  NAND2_X1 U13213 ( .A1(n7184), .A2(n4754), .ZN(n7185) );
  OAI21_X1 U13214 ( .B1(n24072), .B2(n7857), .A(n7562), .ZN(n7245) );
  INV_X1 U13215 ( .A(n7246), .ZN(n7565) );
  NAND2_X1 U13216 ( .A1(n7565), .A2(n7563), .ZN(n7186) );
  NAND2_X1 U13219 ( .A1(n24578), .A2(n7732), .ZN(n7187) );
  XNOR2_X1 U13220 ( .A(n9107), .B(n8909), .ZN(n7195) );
  NAND3_X1 U13221 ( .A1(n3570), .A2(n7867), .A3(n7865), .ZN(n7190) );
  NAND3_X1 U13222 ( .A1(n7860), .A2(n7867), .A3(n7862), .ZN(n7189) );
  NAND2_X1 U13223 ( .A1(n7271), .A2(n4536), .ZN(n7188) );
  NAND2_X1 U13224 ( .A1(n7843), .A2(n24577), .ZN(n7191) );
  NAND2_X1 U13225 ( .A1(n7719), .A2(n7191), .ZN(n7192) );
  NAND2_X1 U13226 ( .A1(n7843), .A2(n8368), .ZN(n7716) );
  OAI21_X1 U13227 ( .B1(n7193), .B2(n7843), .A(n7716), .ZN(n7194) );
  XNOR2_X1 U13228 ( .A(n8772), .B(n9059), .ZN(n8696) );
  XNOR2_X1 U13229 ( .A(n8696), .B(n7195), .ZN(n7207) );
  OR2_X1 U13230 ( .A1(n9067), .A2(n7057), .ZN(n7430) );
  OAI21_X1 U13231 ( .B1(n7812), .B2(n7809), .A(n7430), .ZN(n7198) );
  INV_X1 U13232 ( .A(n7057), .ZN(n7810) );
  NAND2_X1 U13233 ( .A1(n7196), .A2(n7810), .ZN(n7197) );
  INV_X1 U13235 ( .A(n8361), .ZN(n7200) );
  XNOR2_X1 U13236 ( .A(n8633), .B(n7200), .ZN(n8395) );
  INV_X1 U13237 ( .A(n8395), .ZN(n7205) );
  NAND2_X1 U13238 ( .A1(n7615), .A2(n7380), .ZN(n7620) );
  XNOR2_X1 U13239 ( .A(n7205), .B(n7204), .ZN(n7206) );
  NAND2_X1 U13240 ( .A1(n9134), .A2(n9388), .ZN(n9132) );
  OAI21_X1 U13241 ( .B1(n9949), .B2(n9388), .A(n9132), .ZN(n7208) );
  NAND2_X1 U13242 ( .A1(n7208), .A2(n9959), .ZN(n7209) );
  NOR2_X1 U13243 ( .A1(n7666), .A2(n8527), .ZN(n7212) );
  INV_X1 U13244 ( .A(n8533), .ZN(n7213) );
  OAI21_X1 U13246 ( .B1(n8315), .B2(n7217), .A(n8317), .ZN(n7218) );
  OAI21_X1 U13247 ( .B1(n7698), .B2(n8317), .A(n7218), .ZN(n7219) );
  XNOR2_X1 U13248 ( .A(n24946), .B(n8172), .ZN(n7448) );
  OAI21_X1 U13249 ( .B1(n7423), .B2(n4144), .A(n7220), .ZN(n7223) );
  INV_X1 U13250 ( .A(n7674), .ZN(n7225) );
  XNOR2_X1 U13251 ( .A(n8491), .B(n9159), .ZN(n8947) );
  XNOR2_X1 U13252 ( .A(n8947), .B(n7448), .ZN(n7241) );
  INV_X1 U13253 ( .A(n7230), .ZN(n7898) );
  XNOR2_X1 U13254 ( .A(n8867), .B(n8612), .ZN(n7239) );
  XNOR2_X1 U13255 ( .A(n8980), .B(n1767), .ZN(n7238) );
  XNOR2_X1 U13256 ( .A(n7239), .B(n7238), .ZN(n7240) );
  AOI21_X1 U13257 ( .B1(n7773), .B2(n7769), .A(n7776), .ZN(n7244) );
  NAND2_X1 U13258 ( .A1(n7768), .A2(n7767), .ZN(n7242) );
  AOI21_X1 U13259 ( .B1(n7242), .B2(n7527), .A(n7526), .ZN(n7243) );
  NAND2_X1 U13260 ( .A1(n7245), .A2(n7853), .ZN(n7249) );
  INV_X1 U13261 ( .A(n7850), .ZN(n7725) );
  AOI21_X1 U13262 ( .B1(n7725), .B2(n7721), .A(n7857), .ZN(n7247) );
  XNOR2_X1 U13263 ( .A(n8460), .B(n8501), .ZN(n8703) );
  NAND2_X1 U13264 ( .A1(n8511), .A2(n7350), .ZN(n7252) );
  NAND2_X1 U13265 ( .A1(n7255), .A2(n7600), .ZN(n7344) );
  NAND2_X1 U13266 ( .A1(n7595), .A2(n7257), .ZN(n7345) );
  INV_X1 U13267 ( .A(n7597), .ZN(n7256) );
  XNOR2_X1 U13269 ( .A(n8542), .B(n8345), .ZN(n7471) );
  NAND2_X1 U13270 ( .A1(n7444), .A2(n7932), .ZN(n7263) );
  AOI21_X1 U13271 ( .B1(n7445), .B2(n7263), .A(n7923), .ZN(n7264) );
  XNOR2_X1 U13272 ( .A(n8899), .B(n20995), .ZN(n7276) );
  INV_X1 U13273 ( .A(n8368), .ZN(n7714) );
  NAND2_X1 U13274 ( .A1(n7714), .A2(n7843), .ZN(n7267) );
  INV_X1 U13275 ( .A(n7713), .ZN(n7561) );
  AOI21_X1 U13276 ( .B1(n7267), .B2(n7266), .A(n7561), .ZN(n7270) );
  AOI21_X1 U13277 ( .B1(n7268), .B2(n8370), .A(n7714), .ZN(n7269) );
  NAND2_X1 U13278 ( .A1(n7553), .A2(n7865), .ZN(n7275) );
  NAND2_X1 U13279 ( .A1(n7868), .A2(n24576), .ZN(n7274) );
  NAND3_X1 U13280 ( .A1(n7863), .A2(n24576), .A3(n7707), .ZN(n7273) );
  NAND2_X1 U13281 ( .A1(n7271), .A2(n7865), .ZN(n7272) );
  XNOR2_X1 U13282 ( .A(n8989), .B(n8875), .ZN(n8112) );
  NAND2_X1 U13283 ( .A1(n7279), .A2(n7350), .ZN(n7280) );
  NAND3_X1 U13284 ( .A1(n7347), .A2(n5468), .A3(n7351), .ZN(n7282) );
  NAND3_X1 U13285 ( .A1(n8511), .A2(n5468), .A3(n7349), .ZN(n7281) );
  XNOR2_X1 U13286 ( .A(n9139), .B(n8952), .ZN(n7291) );
  INV_X1 U13287 ( .A(n7776), .ZN(n7283) );
  AOI21_X1 U13288 ( .B1(n7283), .B2(n25252), .A(n7527), .ZN(n7289) );
  NAND3_X1 U13289 ( .A1(n23), .A2(n7776), .A3(n7284), .ZN(n7286) );
  XNOR2_X1 U13290 ( .A(n8798), .B(n2743), .ZN(n7290) );
  XNOR2_X1 U13291 ( .A(n7291), .B(n7290), .ZN(n7311) );
  INV_X1 U13292 ( .A(n7293), .ZN(n7297) );
  INV_X1 U13293 ( .A(n8014), .ZN(n7295) );
  NAND2_X1 U13294 ( .A1(n7295), .A2(n8015), .ZN(n7296) );
  NAND2_X1 U13295 ( .A1(n8014), .A2(n8016), .ZN(n7298) );
  NAND2_X1 U13296 ( .A1(n7299), .A2(n7298), .ZN(n7300) );
  XNOR2_X1 U13298 ( .A(n8147), .B(n8132), .ZN(n8734) );
  OAI21_X1 U13299 ( .B1(n7385), .B2(n7617), .A(n7380), .ZN(n7304) );
  NAND3_X1 U13300 ( .A1(n1895), .A2(n7619), .A3(n7618), .ZN(n7302) );
  NAND2_X1 U13301 ( .A1(n7390), .A2(n7760), .ZN(n7306) );
  NAND3_X1 U13302 ( .A1(n7760), .A2(n7307), .A3(n7648), .ZN(n7308) );
  XNOR2_X1 U13304 ( .A(n8799), .B(n8916), .ZN(n8329) );
  NOR2_X1 U13307 ( .A1(n7575), .A2(n7580), .ZN(n7321) );
  XNOR2_X1 U13308 ( .A(n8853), .B(n8959), .ZN(n8363) );
  INV_X1 U13309 ( .A(n8363), .ZN(n7334) );
  INV_X1 U13310 ( .A(n7323), .ZN(n7605) );
  AND2_X1 U13311 ( .A1(n7898), .A2(n248), .ZN(n7328) );
  NAND2_X1 U13312 ( .A1(n7328), .A2(n3469), .ZN(n7333) );
  NAND2_X1 U13313 ( .A1(n7329), .A2(n24103), .ZN(n7331) );
  NAND4_X2 U13314 ( .A1(n7332), .A2(n7333), .A3(n7331), .A4(n7330), .ZN(n8962)
         );
  XNOR2_X1 U13315 ( .A(n8771), .B(n8962), .ZN(n8192) );
  XNOR2_X1 U13316 ( .A(n7334), .B(n8192), .ZN(n7356) );
  NAND2_X1 U13317 ( .A1(n7335), .A2(n7461), .ZN(n7463) );
  NAND2_X1 U13318 ( .A1(n7463), .A2(n2035), .ZN(n7336) );
  NAND2_X1 U13319 ( .A1(n7337), .A2(n7336), .ZN(n7340) );
  NAND2_X1 U13320 ( .A1(n5737), .A2(n7338), .ZN(n7339) );
  NAND2_X1 U13321 ( .A1(n7340), .A2(n7339), .ZN(n8360) );
  OAI211_X1 U13322 ( .C1(n7600), .C2(n7597), .A(n25037), .B(n7341), .ZN(n7343)
         );
  XNOR2_X1 U13323 ( .A(n8964), .B(n8360), .ZN(n7518) );
  OAI211_X1 U13324 ( .C1(n7349), .C2(n7348), .A(n7347), .B(n7346), .ZN(n7353)
         );
  INV_X1 U13325 ( .A(n7350), .ZN(n8509) );
  OAI211_X1 U13326 ( .C1(n8508), .C2(n8511), .A(n7353), .B(n7352), .ZN(n8638)
         );
  XNOR2_X1 U13327 ( .A(n8638), .B(n187), .ZN(n7354) );
  XNOR2_X1 U13328 ( .A(n7518), .B(n7354), .ZN(n7355) );
  AND2_X1 U13329 ( .A1(n7358), .A2(n7413), .ZN(n7359) );
  AOI21_X1 U13330 ( .B1(n7994), .B2(n7360), .A(n3549), .ZN(n7361) );
  NOR2_X2 U13331 ( .A1(n7362), .A2(n7361), .ZN(n8313) );
  NAND2_X1 U13332 ( .A1(n7363), .A2(n7364), .ZN(n7369) );
  NAND3_X1 U13333 ( .A1(n7909), .A2(n7911), .A3(n7628), .ZN(n7368) );
  NAND3_X1 U13334 ( .A1(n7913), .A2(n7910), .A3(n7908), .ZN(n7367) );
  NAND3_X1 U13335 ( .A1(n7913), .A2(n7365), .A3(n7629), .ZN(n7366) );
  INV_X1 U13336 ( .A(n7923), .ZN(n7370) );
  NAND2_X1 U13337 ( .A1(n7370), .A2(n7163), .ZN(n7375) );
  NAND2_X1 U13338 ( .A1(n7372), .A2(n7923), .ZN(n7371) );
  OAI211_X1 U13339 ( .C1(n7372), .C2(n5607), .A(n7371), .B(n7445), .ZN(n7374)
         );
  NAND2_X1 U13341 ( .A1(n5595), .A2(n7640), .ZN(n7378) );
  NAND2_X1 U13342 ( .A1(n7734), .A2(n7733), .ZN(n7376) );
  NAND3_X1 U13343 ( .A1(n7641), .A2(n24578), .A3(n7642), .ZN(n7377) );
  XNOR2_X1 U13344 ( .A(n9182), .B(n8517), .ZN(n8940) );
  XNOR2_X1 U13345 ( .A(n8940), .B(n7379), .ZN(n7402) );
  NAND3_X1 U13348 ( .A1(n7622), .A2(n7385), .A3(n7384), .ZN(n7388) );
  NAND3_X1 U13349 ( .A1(n7617), .A2(n7386), .A3(n7615), .ZN(n7387) );
  NAND3_X2 U13350 ( .A1(n7389), .A2(n7388), .A3(n7387), .ZN(n8786) );
  NAND2_X1 U13351 ( .A1(n7391), .A2(n7648), .ZN(n7394) );
  OAI211_X1 U13352 ( .C1(n7647), .C2(n7760), .A(n7392), .B(n7646), .ZN(n7393)
         );
  XNOR2_X1 U13353 ( .A(n8375), .B(n8786), .ZN(n7400) );
  NAND3_X1 U13354 ( .A1(n7634), .A2(n3347), .A3(n7917), .ZN(n7397) );
  NAND3_X1 U13355 ( .A1(n7449), .A2(n25253), .A3(n7918), .ZN(n7395) );
  XNOR2_X1 U13356 ( .A(n8860), .B(n21169), .ZN(n7399) );
  XNOR2_X1 U13357 ( .A(n7400), .B(n7399), .ZN(n7401) );
  XNOR2_X1 U13358 ( .A(n7402), .B(n7401), .ZN(n10129) );
  NOR2_X1 U13359 ( .A1(n7819), .A2(n7974), .ZN(n7403) );
  AOI22_X1 U13360 ( .A1(n7404), .A2(n7816), .B1(n7403), .B2(n7820), .ZN(n7408)
         );
  NAND2_X1 U13361 ( .A1(n7975), .A2(n7974), .ZN(n7406) );
  NAND2_X1 U13362 ( .A1(n7829), .A2(n7983), .ZN(n7987) );
  OAI21_X1 U13363 ( .B1(n7983), .B2(n7982), .A(n7987), .ZN(n7410) );
  NAND2_X1 U13364 ( .A1(n7410), .A2(n7985), .ZN(n7411) );
  XNOR2_X1 U13365 ( .A(n9015), .B(n8476), .ZN(n8117) );
  OR2_X1 U13366 ( .A1(n7413), .A2(n7412), .ZN(n7502) );
  OAI211_X1 U13367 ( .C1(n7990), .C2(n7993), .A(n7502), .B(n3549), .ZN(n7417)
         );
  INV_X1 U13368 ( .A(n7993), .ZN(n7500) );
  NAND3_X1 U13369 ( .A1(n7500), .A2(n7415), .A3(n7998), .ZN(n7416) );
  INV_X1 U13370 ( .A(n7418), .ZN(n7784) );
  NOR2_X1 U13371 ( .A1(n7788), .A2(n7418), .ZN(n7420) );
  XNOR2_X1 U13372 ( .A(n8119), .B(n8477), .ZN(n8937) );
  INV_X1 U13373 ( .A(n8937), .ZN(n8672) );
  XNOR2_X1 U13374 ( .A(n8672), .B(n8117), .ZN(n7436) );
  INV_X1 U13375 ( .A(n7421), .ZN(n7422) );
  OAI21_X1 U13376 ( .B1(n7422), .B2(n7476), .A(n7423), .ZN(n7426) );
  OAI211_X1 U13377 ( .C1(n7954), .C2(n7426), .A(n7425), .B(n7424), .ZN(n8296)
         );
  INV_X1 U13378 ( .A(n3131), .ZN(n23347) );
  XNOR2_X1 U13379 ( .A(n8296), .B(n23347), .ZN(n7435) );
  NAND2_X1 U13380 ( .A1(n7809), .A2(n7813), .ZN(n7429) );
  MUX2_X1 U13381 ( .A(n7429), .B(n7428), .S(n7812), .Z(n7431) );
  INV_X1 U13382 ( .A(n7809), .ZN(n9071) );
  NAND3_X1 U13383 ( .A1(n7795), .A2(n7432), .A3(n7799), .ZN(n7433) );
  XNOR2_X1 U13384 ( .A(n8754), .B(n8339), .ZN(n7552) );
  MUX2_X1 U13385 ( .A(n7781), .B(n7782), .S(n7789), .Z(n7442) );
  MUX2_X1 U13386 ( .A(n7443), .B(n7442), .S(n7784), .Z(n8780) );
  MUX2_X1 U13387 ( .A(n7445), .B(n7444), .S(n7932), .Z(n7447) );
  XNOR2_X1 U13388 ( .A(n8780), .B(n8492), .ZN(n8279) );
  XNOR2_X1 U13389 ( .A(n7448), .B(n8279), .ZN(n7454) );
  INV_X1 U13390 ( .A(n9034), .ZN(n7451) );
  XNOR2_X1 U13391 ( .A(n7451), .B(n8613), .ZN(n8399) );
  XNOR2_X1 U13392 ( .A(n9155), .B(n3125), .ZN(n7452) );
  XNOR2_X1 U13393 ( .A(n8399), .B(n7452), .ZN(n7453) );
  AOI21_X1 U13394 ( .B1(n7322), .B2(n7890), .A(n7605), .ZN(n7456) );
  INV_X1 U13395 ( .A(n7577), .ZN(n7574) );
  AOI21_X1 U13396 ( .B1(n7574), .B2(n7579), .A(n7576), .ZN(n7458) );
  XNOR2_X1 U13397 ( .A(n8499), .B(n1789), .ZN(n7459) );
  XNOR2_X1 U13398 ( .A(n8287), .B(n7459), .ZN(n7473) );
  OAI211_X1 U13399 ( .C1(n7462), .C2(n7592), .A(n7591), .B(n7461), .ZN(n7466)
         );
  INV_X1 U13400 ( .A(n7463), .ZN(n7465) );
  AOI22_X1 U13401 ( .A1(n7467), .A2(n7466), .B1(n7465), .B2(n7464), .ZN(n8620)
         );
  INV_X1 U13402 ( .A(n8620), .ZN(n8988) );
  INV_X1 U13403 ( .A(n7584), .ZN(n7884) );
  NAND2_X1 U13404 ( .A1(n7581), .A2(n7882), .ZN(n7468) );
  NAND2_X1 U13405 ( .A1(n7468), .A2(n7585), .ZN(n7469) );
  XNOR2_X1 U13407 ( .A(n8988), .B(n25228), .ZN(n8405) );
  XNOR2_X1 U13408 ( .A(n8405), .B(n7471), .ZN(n7472) );
  NOR2_X1 U13409 ( .A1(n7475), .A2(n7474), .ZN(n7479) );
  NAND2_X1 U13410 ( .A1(n7477), .A2(n7476), .ZN(n7478) );
  INV_X1 U13411 ( .A(n9141), .ZN(n7480) );
  XNOR2_X1 U13412 ( .A(n7480), .B(n8238), .ZN(n8467) );
  NAND3_X1 U13413 ( .A1(n7481), .A2(n7577), .A3(n7579), .ZN(n7482) );
  AND2_X1 U13414 ( .A1(n7483), .A2(n7482), .ZN(n7484) );
  XNOR2_X1 U13415 ( .A(n8795), .B(n8147), .ZN(n8580) );
  XNOR2_X1 U13416 ( .A(n8467), .B(n8580), .ZN(n7497) );
  NAND2_X1 U13417 ( .A1(n7485), .A2(n7962), .ZN(n7488) );
  INV_X1 U13418 ( .A(n7966), .ZN(n7486) );
  XNOR2_X1 U13419 ( .A(n9081), .B(n8799), .ZN(n7495) );
  INV_X1 U13420 ( .A(n7942), .ZN(n7490) );
  NAND3_X1 U13421 ( .A1(n7943), .A2(n7490), .A3(n7947), .ZN(n7492) );
  NAND2_X1 U13422 ( .A1(n24475), .A2(n7657), .ZN(n7491) );
  XNOR2_X1 U13423 ( .A(n7495), .B(n7494), .ZN(n7496) );
  XNOR2_X1 U13424 ( .A(n8484), .B(n21623), .ZN(n7511) );
  INV_X1 U13425 ( .A(n7502), .ZN(n7503) );
  OAI21_X1 U13426 ( .B1(n7991), .B2(n7993), .A(n7503), .ZN(n7504) );
  NAND2_X1 U13427 ( .A1(n7505), .A2(n7504), .ZN(n8093) );
  INV_X1 U13428 ( .A(n8093), .ZN(n8485) );
  NOR2_X1 U13429 ( .A1(n25251), .A2(n7674), .ZN(n7508) );
  XNOR2_X1 U13430 ( .A(n8485), .B(n8769), .ZN(n8265) );
  XNOR2_X1 U13431 ( .A(n7511), .B(n8265), .ZN(n7520) );
  OAI211_X1 U13432 ( .C1(n7985), .C2(n7829), .A(n7989), .B(n7982), .ZN(n7512)
         );
  OAI211_X1 U13433 ( .C1(n7977), .C2(n7514), .A(n7975), .B(n7973), .ZN(n7515)
         );
  OAI211_X1 U13434 ( .C1(n7517), .C2(n7977), .A(n7516), .B(n7515), .ZN(n8639)
         );
  XNOR2_X1 U13435 ( .A(n9058), .B(n8639), .ZN(n8391) );
  XNOR2_X1 U13436 ( .A(n7518), .B(n8391), .ZN(n7519) );
  XNOR2_X1 U13437 ( .A(n7520), .B(n7519), .ZN(n8141) );
  OAI22_X1 U13438 ( .A1(n9962), .A2(n9468), .B1(n9964), .B2(n9961), .ZN(n8140)
         );
  INV_X1 U13439 ( .A(n7527), .ZN(n7521) );
  NAND2_X1 U13440 ( .A1(n3013), .A2(n7521), .ZN(n7524) );
  XNOR2_X1 U13442 ( .A(n8790), .B(n8506), .ZN(n8291) );
  XNOR2_X1 U13443 ( .A(n9175), .B(n8786), .ZN(n7534) );
  XNOR2_X1 U13444 ( .A(n7534), .B(n8291), .ZN(n7550) );
  NOR2_X1 U13445 ( .A1(n8014), .A2(n8012), .ZN(n7536) );
  NAND3_X1 U13446 ( .A1(n8014), .A2(n8016), .A3(n25451), .ZN(n7539) );
  NAND3_X1 U13447 ( .A1(n7543), .A2(n7542), .A3(n7758), .ZN(n7545) );
  XNOR2_X1 U13449 ( .A(n9007), .B(n9075), .ZN(n8411) );
  XNOR2_X1 U13450 ( .A(n8375), .B(n763), .ZN(n7548) );
  XNOR2_X1 U13451 ( .A(n8411), .B(n7548), .ZN(n7549) );
  XNOR2_X1 U13452 ( .A(n9194), .B(n16574), .ZN(n7551) );
  XNOR2_X1 U13453 ( .A(n7552), .B(n7551), .ZN(n7571) );
  AOI22_X1 U13454 ( .A1(n7710), .A2(n24576), .B1(n7553), .B2(n7707), .ZN(n7556) );
  NAND2_X1 U13455 ( .A1(n7867), .A2(n7864), .ZN(n7554) );
  INV_X1 U13457 ( .A(n7843), .ZN(n7718) );
  INV_X1 U13458 ( .A(n8370), .ZN(n7715) );
  OAI211_X1 U13459 ( .C1(n8371), .C2(n7843), .A(n7558), .B(n7714), .ZN(n7559)
         );
  XNOR2_X1 U13460 ( .A(n9016), .B(n8880), .ZN(n8385) );
  INV_X1 U13461 ( .A(n7857), .ZN(n7722) );
  NAND3_X1 U13462 ( .A1(n7565), .A2(n7564), .A3(n7563), .ZN(n7724) );
  INV_X1 U13463 ( .A(n7730), .ZN(n7568) );
  XNOR2_X1 U13464 ( .A(n8478), .B(n9191), .ZN(n8269) );
  XNOR2_X1 U13465 ( .A(n8269), .B(n8385), .ZN(n7570) );
  NAND3_X1 U13466 ( .A1(n7887), .A2(n7585), .A3(n7883), .ZN(n7586) );
  XNOR2_X1 U13467 ( .A(n7594), .B(n8889), .ZN(n7614) );
  NOR2_X1 U13469 ( .A1(n7600), .A2(n7597), .ZN(n7599) );
  XNOR2_X1 U13470 ( .A(n8280), .B(n8446), .ZN(n7612) );
  NAND2_X1 U13471 ( .A1(n7890), .A2(n7604), .ZN(n7892) );
  AND2_X1 U13472 ( .A1(n7605), .A2(n7604), .ZN(n7607) );
  XNOR2_X1 U13474 ( .A(n8682), .B(n1810), .ZN(n7611) );
  XNOR2_X1 U13475 ( .A(n7612), .B(n7611), .ZN(n7613) );
  OAI22_X1 U13476 ( .A1(n7622), .A2(n7621), .B1(n7620), .B2(n7619), .ZN(n7623)
         );
  XNOR2_X1 U13477 ( .A(n8285), .B(n8458), .ZN(n8230) );
  AOI21_X1 U13478 ( .B1(n7627), .B2(n7626), .A(n7625), .ZN(n7632) );
  AOI21_X1 U13479 ( .B1(n7630), .B2(n7629), .A(n7628), .ZN(n7631) );
  XNOR2_X1 U13481 ( .A(n8899), .B(n8706), .ZN(n7633) );
  XNOR2_X1 U13482 ( .A(n8230), .B(n7633), .ZN(n7655) );
  AOI21_X1 U13483 ( .B1(n7634), .B2(n3348), .A(n25253), .ZN(n7639) );
  NAND2_X1 U13484 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  NAND3_X1 U13485 ( .A1(n7731), .A2(n7642), .A3(n7732), .ZN(n7643) );
  XNOR2_X1 U13486 ( .A(n8760), .B(n8898), .ZN(n7653) );
  NAND2_X1 U13487 ( .A1(n7760), .A2(n7647), .ZN(n7650) );
  INV_X1 U13488 ( .A(n1754), .ZN(n23225) );
  XNOR2_X1 U13489 ( .A(n9043), .B(n23225), .ZN(n7652) );
  XNOR2_X1 U13490 ( .A(n7653), .B(n7652), .ZN(n7654) );
  NOR2_X1 U13491 ( .A1(n24474), .A2(n7945), .ZN(n7661) );
  INV_X1 U13492 ( .A(n7943), .ZN(n7656) );
  NAND2_X1 U13493 ( .A1(n7943), .A2(n7942), .ZN(n7659) );
  XNOR2_X1 U13494 ( .A(n8721), .B(n8673), .ZN(n7681) );
  OAI211_X1 U13495 ( .C1(n7675), .C2(n7674), .A(n7673), .B(n7672), .ZN(n7679)
         );
  NAND3_X1 U13496 ( .A1(n7677), .A2(n7676), .A3(n3275), .ZN(n7678) );
  XNOR2_X1 U13497 ( .A(n8116), .B(n8296), .ZN(n9020) );
  INV_X1 U13498 ( .A(n9020), .ZN(n7680) );
  XNOR2_X1 U13499 ( .A(n7680), .B(n7681), .ZN(n7706) );
  MUX2_X1 U13500 ( .A(n7685), .B(n7684), .S(n7962), .Z(n7686) );
  OAI21_X2 U13501 ( .B1(n7687), .B2(n7961), .A(n7686), .ZN(n8675) );
  XNOR2_X1 U13502 ( .A(n8270), .B(n8675), .ZN(n7704) );
  NOR2_X1 U13503 ( .A1(n7217), .A2(n7688), .ZN(n7697) );
  NOR2_X1 U13504 ( .A1(n7690), .A2(n7689), .ZN(n7695) );
  INV_X1 U13505 ( .A(n7691), .ZN(n7694) );
  INV_X1 U13506 ( .A(n7692), .ZN(n7693) );
  NAND2_X1 U13507 ( .A1(n8315), .A2(n7217), .ZN(n7696) );
  NAND3_X1 U13508 ( .A1(n7700), .A2(n7699), .A3(n8314), .ZN(n7701) );
  XNOR2_X1 U13509 ( .A(n8203), .B(n23620), .ZN(n7703) );
  XNOR2_X1 U13510 ( .A(n7704), .B(n7703), .ZN(n7705) );
  MUX2_X1 U13511 ( .A(n25217), .B(n9599), .S(n9927), .Z(n7839) );
  NAND2_X1 U13512 ( .A1(n7860), .A2(n7707), .ZN(n7709) );
  AOI21_X1 U13513 ( .B1(n7709), .B2(n7708), .A(n7865), .ZN(n7712) );
  NAND2_X1 U13514 ( .A1(n7714), .A2(n7713), .ZN(n7844) );
  OAI211_X1 U13515 ( .C1(n7718), .C2(n7844), .A(n7717), .B(n7716), .ZN(n7720)
         );
  NAND2_X1 U13516 ( .A1(n7722), .A2(n7721), .ZN(n7723) );
  AND2_X1 U13517 ( .A1(n7724), .A2(n7723), .ZN(n7729) );
  MUX2_X1 U13519 ( .A(n7727), .B(n7858), .S(n7853), .Z(n7728) );
  XNOR2_X1 U13520 ( .A(n8914), .B(n8916), .ZN(n8995) );
  XNOR2_X1 U13521 ( .A(n8797), .B(n8995), .ZN(n7744) );
  NAND2_X1 U13522 ( .A1(n7733), .A2(n7732), .ZN(n7737) );
  XNOR2_X1 U13523 ( .A(n8237), .B(n8690), .ZN(n7742) );
  INV_X1 U13524 ( .A(n7813), .ZN(n7739) );
  NAND3_X1 U13525 ( .A1(n7813), .A2(n8219), .A3(n9067), .ZN(n7740) );
  INV_X1 U13526 ( .A(n2881), .ZN(n23283) );
  XNOR2_X1 U13527 ( .A(n8691), .B(n23283), .ZN(n7741) );
  XNOR2_X1 U13528 ( .A(n7742), .B(n7741), .ZN(n7743) );
  INV_X1 U13530 ( .A(n9925), .ZN(n9346) );
  NOR2_X1 U13531 ( .A1(n25217), .A2(n9925), .ZN(n9929) );
  XNOR2_X1 U13532 ( .A(n9002), .B(n8638), .ZN(n8907) );
  OR2_X1 U13533 ( .A1(n7748), .A2(n8015), .ZN(n7752) );
  OAI21_X1 U13534 ( .B1(n25451), .B2(n8012), .A(n8015), .ZN(n7751) );
  NAND2_X1 U13536 ( .A1(n5202), .A2(n7757), .ZN(n7756) );
  OR2_X1 U13537 ( .A1(n7758), .A2(n7757), .ZN(n8004) );
  XNOR2_X1 U13538 ( .A(n9057), .B(n8965), .ZN(n8191) );
  INV_X1 U13539 ( .A(n8191), .ZN(n7759) );
  XNOR2_X1 U13540 ( .A(n7759), .B(n8907), .ZN(n7780) );
  NOR2_X1 U13541 ( .A1(n7760), .A2(n4880), .ZN(n7764) );
  NAND2_X1 U13542 ( .A1(n7762), .A2(n7761), .ZN(n7763) );
  AOI22_X1 U13543 ( .A1(n7766), .A2(n7765), .B1(n7764), .B2(n7763), .ZN(n8244)
         );
  NOR2_X1 U13544 ( .A1(n7768), .A2(n7767), .ZN(n7772) );
  INV_X1 U13545 ( .A(n7772), .ZN(n7775) );
  OAI21_X1 U13546 ( .B1(n7772), .B2(n7771), .A(n7770), .ZN(n7774) );
  XNOR2_X1 U13548 ( .A(n9106), .B(n3155), .ZN(n7777) );
  XNOR2_X1 U13549 ( .A(n7778), .B(n7777), .ZN(n7779) );
  NAND2_X1 U13550 ( .A1(n7781), .A2(n7788), .ZN(n7786) );
  NAND2_X1 U13551 ( .A1(n7783), .A2(n7782), .ZN(n7785) );
  MUX2_X1 U13552 ( .A(n7786), .B(n7785), .S(n7784), .Z(n7793) );
  NOR2_X1 U13553 ( .A1(n7788), .A2(n7787), .ZN(n7790) );
  OAI21_X1 U13554 ( .B1(n7791), .B2(n7790), .A(n7789), .ZN(n7792) );
  XNOR2_X1 U13555 ( .A(n8313), .B(n8366), .ZN(n9010) );
  INV_X1 U13556 ( .A(n9010), .ZN(n7808) );
  NAND2_X1 U13557 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  AOI21_X1 U13558 ( .B1(n7797), .B2(n7796), .A(n7800), .ZN(n7807) );
  NAND3_X1 U13559 ( .A1(n7800), .A2(n7799), .A3(n7798), .ZN(n7805) );
  NAND3_X1 U13560 ( .A1(n7803), .A2(n7802), .A3(n7801), .ZN(n7804) );
  NAND2_X1 U13561 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  XNOR2_X1 U13562 ( .A(n7808), .B(n8252), .ZN(n7837) );
  OAI21_X1 U13563 ( .B1(n7810), .B2(n9066), .A(n7809), .ZN(n8220) );
  NAND2_X1 U13564 ( .A1(n7814), .A2(n7813), .ZN(n9070) );
  OAI21_X1 U13565 ( .B1(n7819), .B2(n7816), .A(n7971), .ZN(n7818) );
  NAND2_X1 U13566 ( .A1(n7818), .A2(n7817), .ZN(n7824) );
  NAND3_X1 U13567 ( .A1(n7819), .A2(n7973), .A3(n7971), .ZN(n7823) );
  NAND3_X2 U13568 ( .A1(n7824), .A2(n7823), .A3(n7822), .ZN(n8746) );
  XNOR2_X1 U13569 ( .A(n8746), .B(n8507), .ZN(n7835) );
  NAND3_X1 U13570 ( .A1(n7989), .A2(n7983), .A3(n7984), .ZN(n7833) );
  NAND3_X1 U13571 ( .A1(n7983), .A2(n7982), .A3(n7825), .ZN(n7832) );
  XNOR2_X1 U13573 ( .A(n8667), .B(n1891), .ZN(n7834) );
  XNOR2_X1 U13574 ( .A(n7835), .B(n7834), .ZN(n7836) );
  INV_X1 U13575 ( .A(n9599), .ZN(n9604) );
  NOR2_X1 U13576 ( .A1(n9603), .A2(n9604), .ZN(n7838) );
  NOR2_X1 U13577 ( .A1(n7840), .A2(n7714), .ZN(n7845) );
  OAI21_X1 U13578 ( .B1(n7844), .B2(n7843), .A(n7842), .ZN(n8374) );
  INV_X1 U13579 ( .A(n9176), .ZN(n7846) );
  XNOR2_X1 U13580 ( .A(n7846), .B(n8507), .ZN(n7848) );
  XNOR2_X1 U13581 ( .A(n8786), .B(n8517), .ZN(n7847) );
  XNOR2_X1 U13582 ( .A(n7848), .B(n7847), .ZN(n7876) );
  INV_X1 U13583 ( .A(n8450), .ZN(n8126) );
  INV_X1 U13584 ( .A(n7849), .ZN(n7852) );
  NAND2_X1 U13585 ( .A1(n7857), .A2(n24072), .ZN(n7851) );
  AOI21_X1 U13586 ( .B1(n7852), .B2(n7851), .A(n7855), .ZN(n7859) );
  NAND3_X1 U13587 ( .A1(n7855), .A2(n7854), .A3(n7853), .ZN(n7856) );
  XNOR2_X1 U13588 ( .A(n8126), .B(n8789), .ZN(n7874) );
  NAND3_X1 U13589 ( .A1(n4537), .A2(n7862), .A3(n7861), .ZN(n7871) );
  NAND3_X1 U13590 ( .A1(n7865), .A2(n4536), .A3(n7864), .ZN(n7870) );
  NAND3_X1 U13591 ( .A1(n7868), .A2(n7867), .A3(n24576), .ZN(n7869) );
  XNOR2_X1 U13592 ( .A(n9179), .B(n20284), .ZN(n7873) );
  XNOR2_X1 U13593 ( .A(n7874), .B(n7873), .ZN(n7875) );
  XNOR2_X1 U13594 ( .A(n8952), .B(n8799), .ZN(n7878) );
  XNOR2_X1 U13595 ( .A(n8691), .B(n21711), .ZN(n7877) );
  XNOR2_X1 U13596 ( .A(n7878), .B(n7877), .ZN(n7907) );
  INV_X1 U13598 ( .A(n7892), .ZN(n7894) );
  XNOR2_X1 U13599 ( .A(n7895), .B(n8951), .ZN(n9138) );
  INV_X1 U13602 ( .A(n8468), .ZN(n7904) );
  XNOR2_X1 U13603 ( .A(n8796), .B(n7904), .ZN(n7905) );
  XNOR2_X1 U13604 ( .A(n9138), .B(n7905), .ZN(n7906) );
  XNOR2_X1 U13605 ( .A(n8673), .B(n9188), .ZN(n7922) );
  AND2_X1 U13606 ( .A1(n7915), .A2(n7918), .ZN(n7916) );
  MUX2_X1 U13607 ( .A(n430), .B(n7916), .S(n7917), .Z(n7921) );
  NAND2_X1 U13608 ( .A1(n7917), .A2(n3348), .ZN(n7919) );
  AOI21_X1 U13609 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n8078) );
  XNOR2_X1 U13610 ( .A(n9189), .B(n2191), .ZN(n8268) );
  XNOR2_X1 U13611 ( .A(n8268), .B(n7922), .ZN(n7940) );
  INV_X1 U13612 ( .A(n7933), .ZN(n7936) );
  OAI21_X1 U13613 ( .B1(n7924), .B2(n7923), .A(n5607), .ZN(n7935) );
  NOR2_X1 U13614 ( .A1(n7927), .A2(n7926), .ZN(n7931) );
  INV_X1 U13615 ( .A(n7928), .ZN(n7929) );
  XNOR2_X1 U13616 ( .A(n8203), .B(n24445), .ZN(n7938) );
  XNOR2_X1 U13617 ( .A(n8754), .B(n1777), .ZN(n7937) );
  XNOR2_X1 U13618 ( .A(n7938), .B(n7937), .ZN(n7939) );
  XNOR2_X1 U13619 ( .A(n7940), .B(n7939), .ZN(n7941) );
  MUX2_X1 U13620 ( .A(n9939), .B(n9449), .S(n9276), .Z(n8030) );
  INV_X1 U13621 ( .A(n7941), .ZN(n9908) );
  OAI22_X1 U13622 ( .A1(n7944), .A2(n24474), .B1(n7946), .B2(n7943), .ZN(n7951) );
  XNOR2_X1 U13623 ( .A(n9149), .B(n8959), .ZN(n8263) );
  INV_X1 U13624 ( .A(n7954), .ZN(n7955) );
  INV_X1 U13625 ( .A(n9057), .ZN(n7958) );
  XNOR2_X1 U13626 ( .A(n8770), .B(n7958), .ZN(n7959) );
  XNOR2_X1 U13627 ( .A(n8263), .B(n7959), .ZN(n7970) );
  XNOR2_X1 U13629 ( .A(n8698), .B(n8961), .ZN(n7968) );
  XNOR2_X1 U13630 ( .A(n8964), .B(n20825), .ZN(n7967) );
  XNOR2_X1 U13631 ( .A(n7968), .B(n7967), .ZN(n7969) );
  XNOR2_X1 U13632 ( .A(n7969), .B(n7970), .ZN(n9907) );
  AND2_X1 U13633 ( .A1(n9907), .A2(n9908), .ZN(n9937) );
  MUX2_X1 U13634 ( .A(n7976), .B(n7975), .S(n7974), .Z(n7978) );
  XNOR2_X1 U13635 ( .A(n24946), .B(n8069), .ZN(n7981) );
  XNOR2_X1 U13636 ( .A(n7981), .B(n7980), .ZN(n8002) );
  NAND2_X1 U13637 ( .A1(n7989), .A2(n7984), .ZN(n7986) );
  MUX2_X1 U13638 ( .A(n7987), .B(n7986), .S(n7985), .Z(n7988) );
  MUX2_X1 U13639 ( .A(n7992), .B(n7990), .S(n7993), .Z(n7997) );
  NAND2_X1 U13640 ( .A1(n7992), .A2(n7991), .ZN(n7995) );
  XNOR2_X1 U13642 ( .A(n8779), .B(n9158), .ZN(n8000) );
  XNOR2_X1 U13643 ( .A(n8446), .B(n1757), .ZN(n7999) );
  XNOR2_X1 U13644 ( .A(n8000), .B(n7999), .ZN(n8001) );
  MUX2_X1 U13645 ( .A(n9905), .B(n9908), .S(n9939), .Z(n8029) );
  AOI21_X1 U13646 ( .B1(n8004), .B2(n8003), .A(n5202), .ZN(n8008) );
  AOI21_X1 U13647 ( .B1(n8006), .B2(n8005), .A(n432), .ZN(n8007) );
  XNOR2_X1 U13648 ( .A(n8458), .B(n8970), .ZN(n8010) );
  XNOR2_X1 U13649 ( .A(n9043), .B(n92), .ZN(n8009) );
  XNOR2_X1 U13650 ( .A(n8010), .B(n8009), .ZN(n8028) );
  NAND3_X1 U13652 ( .A1(n8013), .A2(n8014), .A3(n8015), .ZN(n8018) );
  XNOR2_X1 U13653 ( .A(n9169), .B(n8501), .ZN(n8288) );
  NAND3_X1 U13654 ( .A1(n3615), .A2(n8024), .A3(n8023), .ZN(n8025) );
  XNOR2_X1 U13655 ( .A(n8542), .B(n9040), .ZN(n8766) );
  XNOR2_X1 U13656 ( .A(n8288), .B(n8766), .ZN(n8027) );
  OAI21_X1 U13658 ( .B1(n10369), .B2(n10363), .A(n8031), .ZN(n8032) );
  XNOR2_X1 U13660 ( .A(n8826), .B(n8675), .ZN(n8297) );
  XNOR2_X1 U13661 ( .A(n8647), .B(n3178), .ZN(n8035) );
  XNOR2_X1 U13662 ( .A(n8036), .B(n8035), .ZN(n8037) );
  XNOR2_X1 U13663 ( .A(n8746), .B(n2033), .ZN(n8038) );
  XNOR2_X1 U13664 ( .A(n8038), .B(n8313), .ZN(n8040) );
  XNOR2_X1 U13665 ( .A(n9114), .B(n8040), .ZN(n8043) );
  XNOR2_X1 U13666 ( .A(n9181), .B(n8651), .ZN(n8041) );
  XNOR2_X1 U13667 ( .A(n9011), .B(n8041), .ZN(n8042) );
  XNOR2_X1 U13668 ( .A(n8782), .B(n25235), .ZN(n8044) );
  XNOR2_X1 U13669 ( .A(n8807), .B(n8682), .ZN(n9092) );
  XNOR2_X1 U13670 ( .A(n9092), .B(n8044), .ZN(n8048) );
  XNOR2_X1 U13671 ( .A(n8278), .B(n8612), .ZN(n8046) );
  XNOR2_X1 U13672 ( .A(n8400), .B(n2042), .ZN(n8045) );
  XNOR2_X1 U13673 ( .A(n8046), .B(n8045), .ZN(n8047) );
  XNOR2_X1 U13675 ( .A(n8965), .B(n1758), .ZN(n8049) );
  XNOR2_X1 U13676 ( .A(n9106), .B(n8638), .ZN(n8052) );
  INV_X1 U13677 ( .A(n9107), .ZN(n8051) );
  XNOR2_X1 U13678 ( .A(n8052), .B(n8051), .ZN(n8310) );
  XNOR2_X1 U13679 ( .A(n8053), .B(n8310), .ZN(n9856) );
  XNOR2_X1 U13680 ( .A(n8913), .B(n8730), .ZN(n8953) );
  XNOR2_X1 U13681 ( .A(n8953), .B(n9124), .ZN(n8057) );
  XNOR2_X1 U13682 ( .A(n24547), .B(n9140), .ZN(n8055) );
  XNOR2_X1 U13683 ( .A(n8916), .B(n20046), .ZN(n8054) );
  XNOR2_X1 U13684 ( .A(n8055), .B(n8054), .ZN(n8056) );
  XNOR2_X1 U13685 ( .A(n8057), .B(n8056), .ZN(n9560) );
  MUX2_X1 U13686 ( .A(n9856), .B(n9560), .S(n238), .Z(n8063) );
  XNOR2_X1 U13687 ( .A(n8812), .B(n8706), .ZN(n9095) );
  XNOR2_X1 U13688 ( .A(n8058), .B(n9095), .ZN(n8062) );
  XNOR2_X1 U13689 ( .A(n8899), .B(n8760), .ZN(n8060) );
  INV_X1 U13690 ( .A(n16), .ZN(n21861) );
  XNOR2_X1 U13691 ( .A(n8896), .B(n21861), .ZN(n8059) );
  XNOR2_X1 U13692 ( .A(n8060), .B(n8059), .ZN(n8061) );
  XNOR2_X1 U13693 ( .A(n8062), .B(n8061), .ZN(n9554) );
  MUX2_X1 U13695 ( .A(n9905), .B(n24511), .S(n9276), .Z(n8068) );
  NAND2_X1 U13696 ( .A1(n9449), .A2(n9907), .ZN(n8066) );
  NAND2_X1 U13697 ( .A1(n9939), .A2(n24511), .ZN(n8065) );
  MUX2_X1 U13698 ( .A(n8066), .B(n8065), .S(n9905), .Z(n8067) );
  OAI21_X1 U13699 ( .B1(n8068), .B2(n9449), .A(n8067), .ZN(n10990) );
  XNOR2_X1 U13700 ( .A(n8865), .B(n8714), .ZN(n8073) );
  XNOR2_X1 U13701 ( .A(n8071), .B(n8070), .ZN(n8072) );
  XNOR2_X1 U13702 ( .A(n8073), .B(n8072), .ZN(n9694) );
  XNOR2_X1 U13703 ( .A(n8478), .B(n8824), .ZN(n8720) );
  OAI21_X1 U13704 ( .B1(n8076), .B2(n435), .A(n8075), .ZN(n8077) );
  NOR2_X1 U13705 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  XNOR2_X1 U13706 ( .A(n8341), .B(n8079), .ZN(n8882) );
  XNOR2_X1 U13707 ( .A(n8720), .B(n8882), .ZN(n8083) );
  XNOR2_X1 U13708 ( .A(n8674), .B(n8339), .ZN(n8081) );
  XNOR2_X1 U13709 ( .A(n8203), .B(n23883), .ZN(n8080) );
  XNOR2_X1 U13710 ( .A(n8081), .B(n8080), .ZN(n8082) );
  XNOR2_X1 U13711 ( .A(n8666), .B(n8507), .ZN(n8085) );
  XNOR2_X1 U13712 ( .A(n8084), .B(n8085), .ZN(n8087) );
  XNOR2_X1 U13713 ( .A(n8375), .B(n19392), .ZN(n8086) );
  XNOR2_X1 U13714 ( .A(n9179), .B(n8412), .ZN(n8862) );
  XNOR2_X1 U13715 ( .A(n8498), .B(n8813), .ZN(n8726) );
  XNOR2_X1 U13716 ( .A(n8088), .B(n9169), .ZN(n8872) );
  XNOR2_X1 U13717 ( .A(n8726), .B(n8872), .ZN(n8092) );
  XNOR2_X1 U13718 ( .A(n8345), .B(n8897), .ZN(n8090) );
  XNOR2_X1 U13719 ( .A(n9043), .B(n853), .ZN(n8089) );
  XNOR2_X1 U13720 ( .A(n8090), .B(n8089), .ZN(n8091) );
  XNOR2_X1 U13721 ( .A(n8635), .B(n8093), .ZN(n8741) );
  XNOR2_X1 U13722 ( .A(n9149), .B(n8361), .ZN(n8855) );
  INV_X1 U13723 ( .A(n8855), .ZN(n8585) );
  XNOR2_X1 U13724 ( .A(n8585), .B(n8741), .ZN(n8097) );
  XNOR2_X1 U13725 ( .A(n8360), .B(n9057), .ZN(n8095) );
  XNOR2_X1 U13726 ( .A(n8699), .B(n912), .ZN(n8094) );
  XNOR2_X1 U13727 ( .A(n8095), .B(n8094), .ZN(n8096) );
  XNOR2_X1 U13729 ( .A(n8353), .B(n9121), .ZN(n8844) );
  INV_X1 U13730 ( .A(n8844), .ZN(n8578) );
  XNOR2_X1 U13731 ( .A(n8578), .B(n8731), .ZN(n8101) );
  XNOR2_X1 U13732 ( .A(n8468), .B(n8687), .ZN(n8099) );
  XNOR2_X1 U13733 ( .A(n8147), .B(n3158), .ZN(n8098) );
  XNOR2_X1 U13734 ( .A(n8099), .B(n8098), .ZN(n8100) );
  XNOR2_X1 U13735 ( .A(n8980), .B(n9035), .ZN(n8103) );
  XNOR2_X1 U13736 ( .A(n8103), .B(n8102), .ZN(n8104) );
  XNOR2_X1 U13737 ( .A(n8698), .B(n9002), .ZN(n8106) );
  INV_X1 U13738 ( .A(n2211), .ZN(n23432) );
  XNOR2_X1 U13739 ( .A(n8962), .B(n23432), .ZN(n8105) );
  XNOR2_X1 U13740 ( .A(n8106), .B(n8105), .ZN(n8111) );
  XNOR2_X1 U13741 ( .A(n25407), .B(n9059), .ZN(n8109) );
  INV_X1 U13742 ( .A(n8853), .ZN(n8107) );
  XNOR2_X1 U13743 ( .A(n8107), .B(n8771), .ZN(n8108) );
  XNOR2_X1 U13744 ( .A(n8108), .B(n8109), .ZN(n8110) );
  XNOR2_X1 U13745 ( .A(n8460), .B(n8458), .ZN(n8113) );
  INV_X1 U13746 ( .A(n2040), .ZN(n22635) );
  XNOR2_X1 U13747 ( .A(n8896), .B(n22635), .ZN(n8115) );
  XNOR2_X1 U13748 ( .A(n8898), .B(n9044), .ZN(n8114) );
  INV_X1 U13749 ( .A(n8116), .ZN(n8340) );
  XNOR2_X1 U13750 ( .A(n8340), .B(n8673), .ZN(n8118) );
  XNOR2_X1 U13751 ( .A(n8118), .B(n8117), .ZN(n8123) );
  XNOR2_X1 U13752 ( .A(n8647), .B(n2746), .ZN(n8120) );
  XNOR2_X1 U13753 ( .A(n8121), .B(n8120), .ZN(n8122) );
  INV_X1 U13754 ( .A(n9182), .ZN(n8124) );
  XNOR2_X1 U13755 ( .A(n8366), .B(n8124), .ZN(n8216) );
  XNOR2_X1 U13756 ( .A(n8125), .B(n8216), .ZN(n8130) );
  XNOR2_X1 U13757 ( .A(n8126), .B(n8651), .ZN(n8128) );
  XNOR2_X1 U13758 ( .A(n8860), .B(n3129), .ZN(n8127) );
  XNOR2_X1 U13759 ( .A(n8128), .B(n8127), .ZN(n8129) );
  XNOR2_X1 U13760 ( .A(n8131), .B(n8198), .ZN(n8136) );
  XNOR2_X1 U13761 ( .A(n8132), .B(n9082), .ZN(n8134) );
  XNOR2_X1 U13762 ( .A(n8691), .B(n2228), .ZN(n8133) );
  XNOR2_X1 U13763 ( .A(n8134), .B(n8133), .ZN(n8135) );
  NAND3_X1 U13764 ( .A1(n9945), .A2(n227), .A3(n24054), .ZN(n8137) );
  INV_X1 U13765 ( .A(n10993), .ZN(n10327) );
  NOR2_X1 U13766 ( .A1(n10924), .A2(n10327), .ZN(n8145) );
  NAND2_X1 U13767 ( .A1(n8140), .A2(n9281), .ZN(n8144) );
  INV_X1 U13768 ( .A(n8141), .ZN(n9469) );
  MUX2_X1 U13769 ( .A(n8146), .B(n8145), .S(n10405), .Z(n8181) );
  XNOR2_X1 U13770 ( .A(n8846), .B(n8917), .ZN(n8236) );
  XNOR2_X1 U13771 ( .A(n8147), .B(n2190), .ZN(n8148) );
  XNOR2_X1 U13772 ( .A(n8149), .B(n8148), .ZN(n8150) );
  XNOR2_X1 U13773 ( .A(n8634), .B(n8909), .ZN(n8852) );
  INV_X1 U13774 ( .A(n9111), .ZN(n8151) );
  XNOR2_X1 U13775 ( .A(n8151), .B(n8852), .ZN(n8156) );
  XNOR2_X1 U13776 ( .A(n8772), .B(n8152), .ZN(n8154) );
  INV_X1 U13777 ( .A(n3133), .ZN(n23072) );
  XNOR2_X1 U13778 ( .A(n8360), .B(n23072), .ZN(n8153) );
  XNOR2_X1 U13779 ( .A(n8154), .B(n8153), .ZN(n8155) );
  XNOR2_X1 U13780 ( .A(n8285), .B(n8620), .ZN(n9096) );
  INV_X1 U13781 ( .A(n9096), .ZN(n8158) );
  XNOR2_X1 U13782 ( .A(n8158), .B(n8301), .ZN(n8162) );
  XNOR2_X1 U13783 ( .A(n9167), .B(n8345), .ZN(n8160) );
  XNOR2_X1 U13784 ( .A(n24056), .B(n4233), .ZN(n8159) );
  XNOR2_X1 U13785 ( .A(n8160), .B(n8159), .ZN(n8161) );
  XNOR2_X2 U13786 ( .A(n8162), .B(n8161), .ZN(n9886) );
  XNOR2_X1 U13787 ( .A(n8596), .B(n8923), .ZN(n8859) );
  XNOR2_X1 U13788 ( .A(n8859), .B(n9115), .ZN(n8166) );
  XNOR2_X1 U13789 ( .A(n8787), .B(n8375), .ZN(n8164) );
  INV_X1 U13790 ( .A(n2087), .ZN(n22745) );
  XNOR2_X1 U13791 ( .A(n9181), .B(n22745), .ZN(n8163) );
  XNOR2_X1 U13792 ( .A(n8164), .B(n8163), .ZN(n8165) );
  INV_X1 U13793 ( .A(Key[44]), .ZN(n21942) );
  INV_X1 U13794 ( .A(n21942), .ZN(n21944) );
  XNOR2_X1 U13795 ( .A(n8755), .B(n21944), .ZN(n8167) );
  XNOR2_X1 U13796 ( .A(n8167), .B(n8339), .ZN(n8169) );
  XNOR2_X1 U13797 ( .A(n9016), .B(n8168), .ZN(n9101) );
  XNOR2_X1 U13798 ( .A(n8169), .B(n9101), .ZN(n8171) );
  XNOR2_X1 U13799 ( .A(n8928), .B(n9196), .ZN(n8170) );
  XNOR2_X1 U13800 ( .A(n8604), .B(n8170), .ZN(n8884) );
  XNOR2_X1 U13801 ( .A(n8171), .B(n8884), .ZN(n9454) );
  NAND2_X1 U13802 ( .A1(n9454), .A2(n25069), .ZN(n8177) );
  XNOR2_X1 U13803 ( .A(n8891), .B(n8588), .ZN(n8868) );
  XNOR2_X1 U13804 ( .A(n8868), .B(n9089), .ZN(n8176) );
  XNOR2_X1 U13805 ( .A(n8278), .B(n641), .ZN(n8173) );
  XNOR2_X1 U13806 ( .A(n8174), .B(n8173), .ZN(n8175) );
  XNOR2_X2 U13807 ( .A(n8176), .B(n8175), .ZN(n9565) );
  AOI21_X1 U13809 ( .B1(n8177), .B2(n9565), .A(n9563), .ZN(n8178) );
  INV_X1 U13810 ( .A(n10994), .ZN(n10326) );
  AND2_X1 U13811 ( .A1(n10326), .A2(n10405), .ZN(n10925) );
  NOR2_X2 U13813 ( .A1(n8181), .A2(n8180), .ZN(n12378) );
  XNOR2_X1 U13814 ( .A(n11914), .B(n12378), .ZN(n11061) );
  XNOR2_X1 U13815 ( .A(n9155), .B(n8782), .ZN(n8713) );
  XNOR2_X1 U13818 ( .A(n8807), .B(n2222), .ZN(n8184) );
  XNOR2_X1 U13819 ( .A(n8778), .B(n8184), .ZN(n8185) );
  XNOR2_X1 U13820 ( .A(n8185), .B(n8186), .ZN(n9843) );
  INV_X1 U13821 ( .A(n8460), .ZN(n8971) );
  XNOR2_X1 U13822 ( .A(n8971), .B(n8499), .ZN(n9165) );
  XNOR2_X1 U13823 ( .A(n8989), .B(n9043), .ZN(n8503) );
  XNOR2_X1 U13824 ( .A(n9165), .B(n8503), .ZN(n8190) );
  XNOR2_X1 U13825 ( .A(n8812), .B(n8898), .ZN(n8188) );
  INV_X1 U13826 ( .A(n2050), .ZN(n21309) );
  XNOR2_X1 U13827 ( .A(n8760), .B(n21309), .ZN(n8187) );
  XNOR2_X1 U13828 ( .A(n8188), .B(n8187), .ZN(n8189) );
  XNOR2_X1 U13829 ( .A(n8191), .B(n8192), .ZN(n8196) );
  XNOR2_X1 U13830 ( .A(n8484), .B(n9107), .ZN(n8194) );
  XNOR2_X1 U13831 ( .A(n9002), .B(n836), .ZN(n8193) );
  XNOR2_X1 U13832 ( .A(n8193), .B(n8194), .ZN(n8195) );
  XNOR2_X1 U13833 ( .A(n8797), .B(n8197), .ZN(n8202) );
  INV_X1 U13834 ( .A(n8198), .ZN(n8200) );
  XNOR2_X1 U13835 ( .A(n9141), .B(n22702), .ZN(n8199) );
  XNOR2_X1 U13836 ( .A(n8200), .B(n8199), .ZN(n8201) );
  XNOR2_X1 U13837 ( .A(n8721), .B(n8340), .ZN(n8204) );
  XNOR2_X1 U13838 ( .A(n8203), .B(n9015), .ZN(n8753) );
  XNOR2_X1 U13840 ( .A(n8826), .B(n9190), .ZN(n8206) );
  XNOR2_X1 U13841 ( .A(n9194), .B(n21335), .ZN(n8205) );
  INV_X1 U13843 ( .A(n8209), .ZN(n8211) );
  INV_X1 U13844 ( .A(n17960), .ZN(n23750) );
  AOI21_X1 U13845 ( .B1(n8211), .B2(n8509), .A(n23750), .ZN(n8210) );
  NAND2_X1 U13846 ( .A1(n8210), .A2(n8514), .ZN(n8214) );
  NAND3_X1 U13847 ( .A1(n8211), .A2(n8509), .A3(n23750), .ZN(n8213) );
  NAND3_X1 U13848 ( .A1(n8214), .A2(n8213), .A3(n8212), .ZN(n8215) );
  XNOR2_X1 U13849 ( .A(n8820), .B(n8215), .ZN(n8218) );
  INV_X1 U13850 ( .A(n8216), .ZN(n8217) );
  NAND2_X1 U13851 ( .A1(n8221), .A2(n8219), .ZN(n9069) );
  OAI211_X1 U13852 ( .C1(n8221), .C2(n8220), .A(n9070), .B(n9069), .ZN(n8222)
         );
  XNOR2_X1 U13853 ( .A(n8222), .B(n8746), .ZN(n8223) );
  AND2_X1 U13854 ( .A1(n25486), .A2(n9845), .ZN(n10122) );
  XNOR2_X1 U13855 ( .A(n8492), .B(n25235), .ZN(n8226) );
  XNOR2_X1 U13856 ( .A(n8868), .B(n8226), .ZN(n8229) );
  XNOR2_X1 U13857 ( .A(n8615), .B(n8446), .ZN(n8684) );
  XNOR2_X1 U13858 ( .A(n8280), .B(n688), .ZN(n8227) );
  XNOR2_X1 U13859 ( .A(n8684), .B(n8227), .ZN(n8228) );
  XNOR2_X1 U13860 ( .A(n8498), .B(n8897), .ZN(n8231) );
  XNOR2_X1 U13861 ( .A(n8231), .B(n8230), .ZN(n8235) );
  XNOR2_X1 U13862 ( .A(n8987), .B(n8874), .ZN(n8233) );
  XNOR2_X1 U13863 ( .A(n24056), .B(n859), .ZN(n8232) );
  XNOR2_X1 U13864 ( .A(n8233), .B(n8232), .ZN(n8234) );
  XNOR2_X1 U13865 ( .A(n8235), .B(n8234), .ZN(n9829) );
  NAND2_X1 U13866 ( .A1(n9832), .A2(n9829), .ZN(n10185) );
  INV_X1 U13867 ( .A(n8236), .ZN(n8239) );
  XNOR2_X1 U13868 ( .A(n8238), .B(n8237), .ZN(n8274) );
  XNOR2_X1 U13869 ( .A(n8239), .B(n8274), .ZN(n8243) );
  XNOR2_X1 U13870 ( .A(n8913), .B(n8687), .ZN(n8241) );
  XNOR2_X1 U13871 ( .A(n8691), .B(n20744), .ZN(n8240) );
  XNOR2_X1 U13872 ( .A(n8241), .B(n8240), .ZN(n8242) );
  XNOR2_X1 U13873 ( .A(n8243), .B(n8242), .ZN(n10175) );
  XNOR2_X1 U13874 ( .A(n9001), .B(n8852), .ZN(n8248) );
  XNOR2_X1 U13875 ( .A(n8699), .B(n2834), .ZN(n8245) );
  XNOR2_X1 U13876 ( .A(n8246), .B(n8245), .ZN(n8247) );
  XNOR2_X1 U13877 ( .A(n8250), .B(n8249), .ZN(n8254) );
  XNOR2_X1 U13878 ( .A(n8923), .B(n876), .ZN(n8251) );
  XNOR2_X1 U13879 ( .A(n8251), .B(n8252), .ZN(n8253) );
  NAND2_X1 U13880 ( .A1(n10186), .A2(n10178), .ZN(n8262) );
  XNOR2_X1 U13881 ( .A(n8928), .B(n8478), .ZN(n8255) );
  XNOR2_X1 U13882 ( .A(n8256), .B(n8255), .ZN(n8260) );
  XNOR2_X1 U13883 ( .A(n8935), .B(n23476), .ZN(n8258) );
  XNOR2_X1 U13884 ( .A(n8673), .B(n8270), .ZN(n8257) );
  XNOR2_X1 U13885 ( .A(n8258), .B(n8257), .ZN(n8259) );
  NAND2_X1 U13886 ( .A1(n10176), .A2(n10177), .ZN(n10181) );
  INV_X1 U13887 ( .A(n10181), .ZN(n8261) );
  XNOR2_X1 U13888 ( .A(n9147), .B(n9058), .ZN(n8851) );
  XNOR2_X1 U13889 ( .A(n8265), .B(n8264), .ZN(n8266) );
  INV_X1 U13890 ( .A(n8523), .ZN(n9804) );
  XNOR2_X1 U13891 ( .A(n9196), .B(n8880), .ZN(n8827) );
  XNOR2_X1 U13892 ( .A(n8270), .B(n2735), .ZN(n8271) );
  XNOR2_X1 U13893 ( .A(n8271), .B(n8827), .ZN(n8272) );
  XNOR2_X1 U13894 ( .A(n8952), .B(n681), .ZN(n8273) );
  XNOR2_X1 U13895 ( .A(n9140), .B(n9081), .ZN(n8843) );
  XNOR2_X1 U13896 ( .A(n8843), .B(n8273), .ZN(n8277) );
  XNOR2_X1 U13897 ( .A(n9121), .B(n8795), .ZN(n8275) );
  XNOR2_X1 U13898 ( .A(n8275), .B(n8274), .ZN(n8276) );
  XNOR2_X1 U13899 ( .A(n8277), .B(n8276), .ZN(n9531) );
  INV_X1 U13900 ( .A(n9531), .ZN(n9533) );
  XNOR2_X1 U13901 ( .A(n8278), .B(n9034), .ZN(n8866) );
  INV_X1 U13902 ( .A(n8866), .ZN(n8805) );
  XNOR2_X1 U13903 ( .A(n8805), .B(n8279), .ZN(n8284) );
  XNOR2_X1 U13904 ( .A(n8491), .B(n8069), .ZN(n8282) );
  XNOR2_X1 U13905 ( .A(n8280), .B(n1935), .ZN(n8281) );
  XNOR2_X1 U13906 ( .A(n8282), .B(n8281), .ZN(n8283) );
  XNOR2_X1 U13908 ( .A(n8285), .B(n2126), .ZN(n8286) );
  XNOR2_X1 U13909 ( .A(n8287), .B(n8286), .ZN(n8290) );
  XNOR2_X1 U13910 ( .A(n25228), .B(n9167), .ZN(n8873) );
  XNOR2_X1 U13911 ( .A(n8873), .B(n8288), .ZN(n8289) );
  OAI22_X1 U13912 ( .A1(n9531), .A2(n8523), .B1(n10113), .B2(n9806), .ZN(n9809) );
  XNOR2_X1 U13913 ( .A(n8292), .B(n8291), .ZN(n8295) );
  XNOR2_X1 U13914 ( .A(n9181), .B(n9075), .ZN(n8858) );
  INV_X1 U13915 ( .A(n1875), .ZN(n21500) );
  XNOR2_X1 U13916 ( .A(n9179), .B(n21500), .ZN(n8293) );
  XNOR2_X1 U13917 ( .A(n8858), .B(n8293), .ZN(n8294) );
  XNOR2_X1 U13918 ( .A(n8295), .B(n8294), .ZN(n9807) );
  INV_X1 U13919 ( .A(n9807), .ZN(n9338) );
  XNOR2_X1 U13920 ( .A(n8604), .B(n8296), .ZN(n8648) );
  XNOR2_X1 U13921 ( .A(n8671), .B(n8648), .ZN(n8300) );
  XNOR2_X1 U13922 ( .A(n8754), .B(n2137), .ZN(n8298) );
  XNOR2_X1 U13923 ( .A(n8297), .B(n8298), .ZN(n8299) );
  INV_X1 U13924 ( .A(n8327), .ZN(n9817) );
  INV_X1 U13925 ( .A(n8301), .ZN(n8302) );
  XNOR2_X1 U13926 ( .A(n8302), .B(n9095), .ZN(n8306) );
  XNOR2_X1 U13927 ( .A(n8899), .B(n9044), .ZN(n8304) );
  XNOR2_X1 U13928 ( .A(n8542), .B(n896), .ZN(n8303) );
  XNOR2_X1 U13929 ( .A(n8304), .B(n8303), .ZN(n8305) );
  XNOR2_X2 U13930 ( .A(n8306), .B(n8305), .ZN(n10169) );
  NAND2_X1 U13931 ( .A1(n9817), .A2(n10169), .ZN(n10172) );
  XNOR2_X1 U13932 ( .A(n8964), .B(n1855), .ZN(n8308) );
  INV_X1 U13933 ( .A(n8634), .ZN(n8307) );
  XNOR2_X1 U13934 ( .A(n8308), .B(n8307), .ZN(n8309) );
  XNOR2_X1 U13935 ( .A(n8309), .B(n8696), .ZN(n8312) );
  INV_X1 U13936 ( .A(n8310), .ZN(n8311) );
  XNOR2_X1 U13938 ( .A(n8596), .B(n8313), .ZN(n8652) );
  XNOR2_X1 U13939 ( .A(n9114), .B(n8652), .ZN(n8324) );
  MUX2_X1 U13940 ( .A(n8317), .B(n8315), .S(n8314), .Z(n8320) );
  NAND3_X1 U13941 ( .A1(n8317), .A2(n8316), .A3(n433), .ZN(n8318) );
  XNOR2_X1 U13942 ( .A(n8551), .B(n20690), .ZN(n8322) );
  XNOR2_X1 U13943 ( .A(n8787), .B(n8786), .ZN(n8321) );
  XNOR2_X1 U13944 ( .A(n8322), .B(n8321), .ZN(n8323) );
  XNOR2_X1 U13945 ( .A(n8324), .B(n8323), .ZN(n10170) );
  INV_X1 U13946 ( .A(n10170), .ZN(n9814) );
  XNOR2_X1 U13947 ( .A(n8781), .B(n8612), .ZN(n8325) );
  XNOR2_X1 U13948 ( .A(n25020), .B(n8325), .ZN(n8326) );
  XNOR2_X1 U13949 ( .A(n8846), .B(n20609), .ZN(n8328) );
  XNOR2_X1 U13950 ( .A(n8689), .B(n8328), .ZN(n8331) );
  XNOR2_X1 U13951 ( .A(n8329), .B(n9124), .ZN(n8330) );
  XNOR2_X1 U13953 ( .A(n8333), .B(n8867), .ZN(n8335) );
  XNOR2_X1 U13954 ( .A(n8491), .B(n1827), .ZN(n8334) );
  XNOR2_X1 U13955 ( .A(n8335), .B(n8334), .ZN(n8338) );
  XNOR2_X1 U13956 ( .A(n8779), .B(n8981), .ZN(n8539) );
  XNOR2_X1 U13957 ( .A(n8336), .B(n9158), .ZN(n8715) );
  XNOR2_X1 U13958 ( .A(n8715), .B(n8539), .ZN(n8337) );
  XNOR2_X1 U13959 ( .A(n8339), .B(n9188), .ZN(n8719) );
  XNOR2_X1 U13960 ( .A(n8340), .B(n9195), .ZN(n8558) );
  XNOR2_X1 U13961 ( .A(n8558), .B(n8719), .ZN(n8344) );
  XNOR2_X1 U13962 ( .A(n8341), .B(n23679), .ZN(n8342) );
  BUF_X2 U13963 ( .A(n10100), .Z(n10095) );
  XNOR2_X1 U13965 ( .A(n8501), .B(n8406), .ZN(n8346) );
  XNOR2_X1 U13966 ( .A(n8725), .B(n8346), .ZN(n8350) );
  XNOR2_X1 U13967 ( .A(n9040), .B(n8898), .ZN(n8544) );
  INV_X1 U13968 ( .A(n663), .ZN(n8347) );
  XNOR2_X1 U13969 ( .A(n8875), .B(n8347), .ZN(n8348) );
  XNOR2_X1 U13970 ( .A(n8544), .B(n8348), .ZN(n8349) );
  XNOR2_X1 U13971 ( .A(n8350), .B(n8349), .ZN(n9515) );
  XNOR2_X1 U13972 ( .A(n8354), .B(n8353), .ZN(n8356) );
  XNOR2_X1 U13973 ( .A(n8796), .B(n8914), .ZN(n8561) );
  INV_X1 U13974 ( .A(n8561), .ZN(n8355) );
  XNOR2_X1 U13975 ( .A(n8355), .B(n8356), .ZN(n8358) );
  XNOR2_X1 U13976 ( .A(n8358), .B(n8357), .ZN(n8359) );
  XNOR2_X1 U13977 ( .A(n8961), .B(n8360), .ZN(n8738) );
  XNOR2_X1 U13978 ( .A(n8361), .B(n2761), .ZN(n8362) );
  XNOR2_X1 U13979 ( .A(n8738), .B(n8362), .ZN(n8365) );
  XNOR2_X1 U13980 ( .A(n8770), .B(n9002), .ZN(n8567) );
  XNOR2_X1 U13981 ( .A(n8363), .B(n8567), .ZN(n8364) );
  XNOR2_X2 U13982 ( .A(n8365), .B(n8364), .ZN(n10099) );
  NAND2_X1 U13984 ( .A1(n24878), .A2(n8370), .ZN(n8369) );
  OAI211_X1 U13985 ( .C1(n8371), .C2(n8370), .A(n8369), .B(n8368), .ZN(n8372)
         );
  INV_X1 U13986 ( .A(n8372), .ZN(n8373) );
  OR2_X1 U13987 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  XNOR2_X1 U13988 ( .A(n8376), .B(n8375), .ZN(n8745) );
  XNOR2_X1 U13989 ( .A(n8745), .B(n8549), .ZN(n8380) );
  XNOR2_X1 U13990 ( .A(n8517), .B(n8860), .ZN(n8378) );
  XNOR2_X1 U13991 ( .A(n8412), .B(n1896), .ZN(n8377) );
  XNOR2_X1 U13992 ( .A(n8378), .B(n8377), .ZN(n8379) );
  INV_X1 U13994 ( .A(n8385), .ZN(n8386) );
  XNOR2_X1 U13995 ( .A(n8720), .B(n8386), .ZN(n8390) );
  XNOR2_X1 U13996 ( .A(n9195), .B(n2236), .ZN(n8388) );
  XNOR2_X1 U13997 ( .A(n8388), .B(n8387), .ZN(n8389) );
  XNOR2_X1 U13998 ( .A(n8770), .B(n2990), .ZN(n8393) );
  INV_X1 U13999 ( .A(n8391), .ZN(n8392) );
  XNOR2_X1 U14000 ( .A(n8393), .B(n8392), .ZN(n8397) );
  INV_X1 U14001 ( .A(n8741), .ZN(n8394) );
  XNOR2_X1 U14002 ( .A(n8394), .B(n8395), .ZN(n8396) );
  XNOR2_X1 U14003 ( .A(n8396), .B(n8397), .ZN(n9384) );
  INV_X1 U14004 ( .A(n9384), .ZN(n9849) );
  NOR2_X1 U14005 ( .A1(n10161), .A2(n9849), .ZN(n8420) );
  XNOR2_X1 U14006 ( .A(n8398), .B(n8399), .ZN(n8404) );
  XNOR2_X1 U14007 ( .A(n8779), .B(n8492), .ZN(n8402) );
  XNOR2_X1 U14008 ( .A(n8400), .B(n881), .ZN(n8401) );
  XNOR2_X1 U14009 ( .A(n8402), .B(n8401), .ZN(n8403) );
  XNOR2_X1 U14010 ( .A(n8403), .B(n8404), .ZN(n10158) );
  XNOR2_X1 U14011 ( .A(n8405), .B(n8726), .ZN(n8410) );
  XNOR2_X1 U14012 ( .A(n9040), .B(n8406), .ZN(n8408) );
  XNOR2_X1 U14013 ( .A(n8896), .B(n3115), .ZN(n8407) );
  XNOR2_X1 U14014 ( .A(n8408), .B(n8407), .ZN(n8409) );
  INV_X1 U14015 ( .A(n9348), .ZN(n9592) );
  XNOR2_X1 U14017 ( .A(n8789), .B(n8651), .ZN(n8414) );
  XNOR2_X1 U14018 ( .A(n8412), .B(n1826), .ZN(n8413) );
  XNOR2_X1 U14019 ( .A(n8414), .B(n8413), .ZN(n8415) );
  NAND2_X1 U14022 ( .A1(n8417), .A2(n9851), .ZN(n8418) );
  XNOR2_X1 U14023 ( .A(n8796), .B(n9081), .ZN(n8423) );
  XNOR2_X1 U14024 ( .A(n8423), .B(n8422), .ZN(n8424) );
  XNOR2_X1 U14025 ( .A(n8425), .B(n8424), .ZN(n9349) );
  NAND3_X1 U14026 ( .A1(n2311), .A2(n24470), .A3(n10935), .ZN(n8426) );
  INV_X1 U14027 ( .A(n11464), .ZN(n8664) );
  XNOR2_X1 U14028 ( .A(n8427), .B(n8428), .ZN(n8831) );
  XNOR2_X1 U14029 ( .A(n8994), .B(n8831), .ZN(n8432) );
  XNOR2_X1 U14030 ( .A(n8917), .B(n2031), .ZN(n8429) );
  XNOR2_X1 U14031 ( .A(n8430), .B(n8429), .ZN(n8431) );
  XNOR2_X1 U14032 ( .A(n8432), .B(n8431), .ZN(n10080) );
  XNOR2_X1 U14033 ( .A(n8635), .B(n9107), .ZN(n8835) );
  INV_X1 U14034 ( .A(n8772), .ZN(n8433) );
  XNOR2_X1 U14035 ( .A(n8433), .B(n8909), .ZN(n8434) );
  XNOR2_X1 U14036 ( .A(n8835), .B(n8434), .ZN(n8438) );
  XNOR2_X1 U14037 ( .A(n8962), .B(n673), .ZN(n8435) );
  XNOR2_X1 U14038 ( .A(n8436), .B(n8435), .ZN(n8437) );
  XNOR2_X1 U14039 ( .A(n8439), .B(n8824), .ZN(n8440) );
  XNOR2_X1 U14040 ( .A(n8440), .B(n8441), .ZN(n8443) );
  XNOR2_X1 U14041 ( .A(n8755), .B(n8935), .ZN(n8442) );
  XNOR2_X1 U14042 ( .A(n8442), .B(n8673), .ZN(n9021) );
  XNOR2_X1 U14043 ( .A(n8443), .B(n9021), .ZN(n9787) );
  XNOR2_X1 U14044 ( .A(n8445), .B(n8444), .ZN(n8448) );
  XNOR2_X1 U14045 ( .A(n8447), .B(n25235), .ZN(n8983) );
  NAND2_X1 U14047 ( .A1(n24575), .A2(n4256), .ZN(n8456) );
  XNOR2_X1 U14048 ( .A(n9182), .B(n21553), .ZN(n8449) );
  XNOR2_X1 U14049 ( .A(n8449), .B(n8923), .ZN(n8451) );
  XNOR2_X1 U14050 ( .A(n8452), .B(n8818), .ZN(n8453) );
  XNOR2_X1 U14051 ( .A(n8453), .B(n9011), .ZN(n8454) );
  INV_X1 U14052 ( .A(n10082), .ZN(n9306) );
  NAND2_X1 U14053 ( .A1(n8456), .A2(n8455), .ZN(n8465) );
  XNOR2_X1 U14054 ( .A(n8458), .B(n8457), .ZN(n8985) );
  INV_X1 U14055 ( .A(n8985), .ZN(n8704) );
  XNOR2_X1 U14056 ( .A(n8704), .B(n8459), .ZN(n8464) );
  XNOR2_X1 U14057 ( .A(n8460), .B(n8987), .ZN(n8462) );
  INV_X1 U14058 ( .A(n869), .ZN(n22440) );
  XNOR2_X1 U14059 ( .A(n8813), .B(n22440), .ZN(n8461) );
  XNOR2_X1 U14060 ( .A(n8462), .B(n8461), .ZN(n8463) );
  MUX2_X2 U14061 ( .A(n8466), .B(n8465), .S(n10088), .Z(n11178) );
  INV_X1 U14062 ( .A(n8467), .ZN(n8470) );
  XNOR2_X1 U14063 ( .A(n8468), .B(n8845), .ZN(n9080) );
  INV_X1 U14064 ( .A(n9080), .ZN(n8469) );
  XNOR2_X1 U14065 ( .A(n8470), .B(n8469), .ZN(n8474) );
  XNOR2_X1 U14066 ( .A(n8798), .B(n8952), .ZN(n8472) );
  XNOR2_X1 U14067 ( .A(n8690), .B(n2215), .ZN(n8471) );
  XNOR2_X1 U14068 ( .A(n8472), .B(n8471), .ZN(n8473) );
  XNOR2_X1 U14069 ( .A(n8474), .B(n8473), .ZN(n8483) );
  INV_X1 U14070 ( .A(n8483), .ZN(n9797) );
  XNOR2_X1 U14071 ( .A(n8475), .B(n8476), .ZN(n8722) );
  INV_X1 U14072 ( .A(n8722), .ZN(n9051) );
  XNOR2_X1 U14073 ( .A(n9051), .B(n8753), .ZN(n8482) );
  XNOR2_X1 U14074 ( .A(n8477), .B(n8478), .ZN(n8480) );
  XNOR2_X1 U14075 ( .A(n8675), .B(n2757), .ZN(n8479) );
  XNOR2_X1 U14076 ( .A(n8480), .B(n8479), .ZN(n8481) );
  NAND2_X1 U14077 ( .A1(n9797), .A2(n246), .ZN(n8497) );
  XNOR2_X1 U14078 ( .A(n8484), .B(n8853), .ZN(n8739) );
  XNOR2_X1 U14079 ( .A(n8771), .B(n9057), .ZN(n8487) );
  XNOR2_X1 U14080 ( .A(n8485), .B(n5286), .ZN(n8486) );
  XNOR2_X1 U14081 ( .A(n8487), .B(n8486), .ZN(n8488) );
  XNOR2_X1 U14082 ( .A(n8489), .B(n8488), .ZN(n9998) );
  INV_X1 U14083 ( .A(n9998), .ZN(n9796) );
  INV_X1 U14084 ( .A(n9796), .ZN(n9669) );
  INV_X1 U14085 ( .A(n9155), .ZN(n8490) );
  XNOR2_X1 U14086 ( .A(n8867), .B(n8490), .ZN(n9033) );
  XNOR2_X1 U14087 ( .A(n9033), .B(n8778), .ZN(n8496) );
  XNOR2_X1 U14088 ( .A(n8492), .B(n8491), .ZN(n8494) );
  XNOR2_X1 U14089 ( .A(n8682), .B(n494), .ZN(n8493) );
  XNOR2_X1 U14090 ( .A(n8494), .B(n8493), .ZN(n8495) );
  INV_X1 U14091 ( .A(n9798), .ZN(n9310) );
  XNOR2_X1 U14092 ( .A(n8498), .B(n8706), .ZN(n8500) );
  XNOR2_X1 U14093 ( .A(n8499), .B(n8875), .ZN(n9042) );
  XNOR2_X1 U14094 ( .A(n9042), .B(n8500), .ZN(n8505) );
  INV_X1 U14095 ( .A(n891), .ZN(n21359) );
  XNOR2_X1 U14096 ( .A(n8501), .B(n21359), .ZN(n8502) );
  XNOR2_X1 U14097 ( .A(n8503), .B(n8502), .ZN(n8504) );
  INV_X1 U14098 ( .A(n8521), .ZN(n9671) );
  NAND2_X1 U14099 ( .A1(n1796), .A2(n9671), .ZN(n8522) );
  XNOR2_X1 U14100 ( .A(n8506), .B(n8507), .ZN(n8516) );
  NAND2_X1 U14101 ( .A1(n8508), .A2(n8512), .ZN(n8510) );
  OAI211_X1 U14102 ( .C1(n8512), .C2(n8511), .A(n8510), .B(n8509), .ZN(n8513)
         );
  NAND2_X1 U14103 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  XNOR2_X1 U14104 ( .A(n8515), .B(n8860), .ZN(n8748) );
  INV_X1 U14105 ( .A(n8748), .ZN(n9065) );
  XNOR2_X1 U14106 ( .A(n8516), .B(n9065), .ZN(n8520) );
  XNOR2_X1 U14107 ( .A(n8667), .B(n3062), .ZN(n8518) );
  NOR2_X1 U14108 ( .A1(n11178), .A2(n24591), .ZN(n8611) );
  OAI21_X1 U14109 ( .B1(n9533), .B2(n9338), .A(n9805), .ZN(n8526) );
  INV_X1 U14110 ( .A(n9806), .ZN(n10116) );
  NOR2_X1 U14111 ( .A1(n9805), .A2(n9530), .ZN(n8524) );
  OAI21_X1 U14112 ( .B1(n9339), .B2(n8524), .A(n9807), .ZN(n8525) );
  NAND2_X1 U14113 ( .A1(n8530), .A2(n8527), .ZN(n8529) );
  OAI211_X1 U14114 ( .C1(n8531), .C2(n8530), .A(n8529), .B(n8528), .ZN(n8532)
         );
  OAI211_X1 U14115 ( .C1(n269), .C2(n8534), .A(n8533), .B(n8532), .ZN(n8535)
         );
  XNOR2_X1 U14116 ( .A(n9035), .B(n8535), .ZN(n8536) );
  XNOR2_X1 U14117 ( .A(n8537), .B(n8536), .ZN(n8950) );
  INV_X1 U14118 ( .A(n8950), .ZN(n8541) );
  XNOR2_X1 U14119 ( .A(n8682), .B(n21423), .ZN(n8538) );
  INV_X1 U14120 ( .A(n9495), .ZN(n9782) );
  XNOR2_X1 U14121 ( .A(n8543), .B(n8760), .ZN(n8977) );
  XNOR2_X1 U14122 ( .A(n8977), .B(n8544), .ZN(n8547) );
  XNOR2_X1 U14123 ( .A(n24056), .B(n886), .ZN(n8545) );
  XNOR2_X1 U14124 ( .A(n8706), .B(n8545), .ZN(n8546) );
  XNOR2_X1 U14126 ( .A(n8667), .B(n2039), .ZN(n8548) );
  XNOR2_X1 U14127 ( .A(n8548), .B(n8923), .ZN(n8550) );
  XNOR2_X1 U14128 ( .A(n8549), .B(n8550), .ZN(n8555) );
  XNOR2_X1 U14129 ( .A(n8746), .B(n8551), .ZN(n8553) );
  XNOR2_X1 U14130 ( .A(n8553), .B(n8552), .ZN(n8941) );
  INV_X1 U14131 ( .A(n8941), .ZN(n8554) );
  XNOR2_X1 U14132 ( .A(n8554), .B(n8555), .ZN(n9297) );
  NAND2_X1 U14133 ( .A1(n9676), .A2(n9780), .ZN(n8575) );
  XNOR2_X1 U14134 ( .A(n8675), .B(n2100), .ZN(n8556) );
  XNOR2_X1 U14135 ( .A(n8730), .B(n8690), .ZN(n8560) );
  XNOR2_X1 U14136 ( .A(n8561), .B(n8560), .ZN(n8564) );
  XNOR2_X1 U14137 ( .A(n9082), .B(n8799), .ZN(n8955) );
  XNOR2_X1 U14138 ( .A(n8917), .B(n1856), .ZN(n8562) );
  XNOR2_X1 U14139 ( .A(n8955), .B(n8562), .ZN(n8563) );
  XNOR2_X1 U14140 ( .A(n8563), .B(n8564), .ZN(n9496) );
  INV_X1 U14141 ( .A(n9496), .ZN(n9295) );
  INV_X1 U14142 ( .A(n9059), .ZN(n8565) );
  XNOR2_X1 U14143 ( .A(n8565), .B(n8909), .ZN(n8566) );
  XNOR2_X1 U14144 ( .A(n8964), .B(n9106), .ZN(n8569) );
  XNOR2_X1 U14145 ( .A(n8965), .B(n1833), .ZN(n8568) );
  XNOR2_X1 U14146 ( .A(n8569), .B(n8568), .ZN(n8570) );
  NAND3_X1 U14148 ( .A1(n9782), .A2(n25454), .A3(n1348), .ZN(n8573) );
  NOR2_X1 U14149 ( .A1(n11168), .A2(n24957), .ZN(n8610) );
  XNOR2_X1 U14150 ( .A(n8576), .B(n8951), .ZN(n8577) );
  XNOR2_X1 U14152 ( .A(n8798), .B(n14398), .ZN(n8579) );
  XNOR2_X1 U14153 ( .A(n8580), .B(n8579), .ZN(n8581) );
  XNOR2_X1 U14154 ( .A(n8582), .B(n8581), .ZN(n9485) );
  XNOR2_X1 U14155 ( .A(n8771), .B(n8634), .ZN(n8583) );
  XNOR2_X1 U14156 ( .A(n8738), .B(n8583), .ZN(n8587) );
  XNOR2_X1 U14157 ( .A(n8769), .B(n677), .ZN(n8584) );
  XNOR2_X1 U14158 ( .A(n8585), .B(n8584), .ZN(n8586) );
  XNOR2_X1 U14159 ( .A(n8586), .B(n8587), .ZN(n9484) );
  XNOR2_X1 U14160 ( .A(n8588), .B(n8780), .ZN(n8614) );
  XNOR2_X1 U14161 ( .A(n8865), .B(n8614), .ZN(n8591) );
  XNOR2_X1 U14162 ( .A(n8980), .B(n925), .ZN(n8589) );
  XNOR2_X1 U14163 ( .A(n8715), .B(n8589), .ZN(n8590) );
  XNOR2_X1 U14164 ( .A(n1337), .B(n8725), .ZN(n8595) );
  XNOR2_X1 U14165 ( .A(n8874), .B(n9041), .ZN(n8593) );
  XNOR2_X1 U14166 ( .A(n8989), .B(n2739), .ZN(n8592) );
  XNOR2_X1 U14167 ( .A(n8593), .B(n8592), .ZN(n8594) );
  OAI22_X1 U14168 ( .A1(n9485), .A2(n9484), .B1(n10006), .B2(n10008), .ZN(
        n10012) );
  XNOR2_X1 U14169 ( .A(n8790), .B(n8597), .ZN(n8598) );
  XNOR2_X1 U14170 ( .A(n8745), .B(n8598), .ZN(n8601) );
  XNOR2_X1 U14171 ( .A(n8599), .B(n8862), .ZN(n8600) );
  XNOR2_X1 U14172 ( .A(n8601), .B(n8600), .ZN(n9299) );
  INV_X1 U14173 ( .A(n9299), .ZN(n9724) );
  INV_X1 U14174 ( .A(n9485), .ZN(n9725) );
  INV_X1 U14175 ( .A(n8719), .ZN(n8602) );
  XNOR2_X1 U14176 ( .A(n8602), .B(n8882), .ZN(n8608) );
  INV_X1 U14177 ( .A(n9191), .ZN(n8603) );
  XNOR2_X1 U14178 ( .A(n8604), .B(n8603), .ZN(n8606) );
  XNOR2_X1 U14179 ( .A(n9015), .B(n23983), .ZN(n8605) );
  XNOR2_X1 U14180 ( .A(n8606), .B(n8605), .ZN(n8607) );
  INV_X1 U14181 ( .A(n9484), .ZN(n9301) );
  MUX2_X1 U14182 ( .A(n8611), .B(n8610), .S(n1338), .Z(n8663) );
  XNOR2_X1 U14183 ( .A(n8613), .B(n8612), .ZN(n8982) );
  XNOR2_X1 U14184 ( .A(n8982), .B(n8614), .ZN(n8619) );
  XNOR2_X1 U14185 ( .A(n8806), .B(n2826), .ZN(n8617) );
  XNOR2_X1 U14186 ( .A(n8617), .B(n9090), .ZN(n8618) );
  XNOR2_X1 U14187 ( .A(n8619), .B(n8618), .ZN(n9772) );
  INV_X1 U14188 ( .A(n9772), .ZN(n8644) );
  XNOR2_X1 U14189 ( .A(n8622), .B(n8621), .ZN(n8626) );
  XNOR2_X1 U14190 ( .A(n8899), .B(n8896), .ZN(n8624) );
  XNOR2_X1 U14191 ( .A(n8813), .B(n2744), .ZN(n8623) );
  XNOR2_X1 U14192 ( .A(n8624), .B(n8623), .ZN(n8625) );
  XNOR2_X1 U14193 ( .A(n24547), .B(n8687), .ZN(n9122) );
  XNOR2_X1 U14194 ( .A(n9122), .B(n8628), .ZN(n8632) );
  XNOR2_X1 U14195 ( .A(n8795), .B(n8916), .ZN(n8630) );
  INV_X1 U14196 ( .A(Key[119]), .ZN(n21533) );
  XNOR2_X1 U14197 ( .A(n8630), .B(n8629), .ZN(n8631) );
  XNOR2_X1 U14198 ( .A(n8633), .B(n8699), .ZN(n9110) );
  INV_X1 U14199 ( .A(n9110), .ZN(n8637) );
  XNOR2_X1 U14200 ( .A(n8635), .B(n8634), .ZN(n8636) );
  XNOR2_X1 U14201 ( .A(n8637), .B(n8636), .ZN(n8642) );
  XNOR2_X1 U14202 ( .A(n8639), .B(n8638), .ZN(n9003) );
  XNOR2_X1 U14203 ( .A(n8769), .B(n1745), .ZN(n8640) );
  XNOR2_X1 U14204 ( .A(n9003), .B(n8640), .ZN(n8641) );
  OAI21_X1 U14205 ( .B1(n8644), .B2(n4254), .A(n8643), .ZN(n9525) );
  NAND2_X1 U14206 ( .A1(n8644), .A2(n10109), .ZN(n8659) );
  XNOR2_X1 U14207 ( .A(n8824), .B(n9016), .ZN(n8646) );
  XNOR2_X1 U14208 ( .A(n9191), .B(n3190), .ZN(n8645) );
  XNOR2_X1 U14209 ( .A(n8646), .B(n8645), .ZN(n8650) );
  XNOR2_X1 U14210 ( .A(n8647), .B(n8674), .ZN(n9102) );
  XNOR2_X1 U14211 ( .A(n9102), .B(n8648), .ZN(n8649) );
  XNOR2_X1 U14212 ( .A(n8649), .B(n8650), .ZN(n9328) );
  INV_X1 U14213 ( .A(n9328), .ZN(n9775) );
  INV_X1 U14214 ( .A(n10104), .ZN(n9526) );
  NOR2_X1 U14215 ( .A1(n9775), .A2(n9526), .ZN(n8658) );
  XNOR2_X1 U14216 ( .A(n8666), .B(n8651), .ZN(n9117) );
  INV_X1 U14217 ( .A(n9117), .ZN(n8922) );
  XNOR2_X1 U14218 ( .A(n8652), .B(n8922), .ZN(n8656) );
  XNOR2_X1 U14219 ( .A(n8790), .B(n8818), .ZN(n8654) );
  XNOR2_X1 U14220 ( .A(n9007), .B(n1724), .ZN(n8653) );
  XNOR2_X1 U14221 ( .A(n8654), .B(n8653), .ZN(n8655) );
  NAND2_X1 U14222 ( .A1(n25393), .A2(n4254), .ZN(n8657) );
  AOI22_X1 U14223 ( .A1(n9525), .A2(n8659), .B1(n8658), .B2(n8657), .ZN(n8660)
         );
  INV_X1 U14224 ( .A(n8660), .ZN(n11170) );
  NOR2_X1 U14225 ( .A1(n11170), .A2(n24957), .ZN(n10937) );
  INV_X1 U14226 ( .A(n11172), .ZN(n11175) );
  OAI21_X1 U14227 ( .B1(n8660), .B2(n11175), .A(n11178), .ZN(n8661) );
  NOR2_X1 U14228 ( .A1(n10937), .A2(n8661), .ZN(n8662) );
  XNOR2_X1 U14230 ( .A(n8664), .B(n11840), .ZN(n11435) );
  XNOR2_X1 U14231 ( .A(n8666), .B(n9073), .ZN(n8669) );
  XNOR2_X1 U14232 ( .A(n8667), .B(n887), .ZN(n8668) );
  XNOR2_X1 U14233 ( .A(n8669), .B(n8668), .ZN(n8670) );
  INV_X1 U14234 ( .A(n9664), .ZN(n9221) );
  XNOR2_X1 U14235 ( .A(n8675), .B(n2005), .ZN(n8676) );
  XNOR2_X1 U14236 ( .A(n8677), .B(n8676), .ZN(n8678) );
  INV_X1 U14237 ( .A(n9981), .ZN(n9736) );
  XNOR2_X1 U14239 ( .A(n24598), .B(n8947), .ZN(n8686) );
  XNOR2_X1 U14240 ( .A(n8682), .B(n1768), .ZN(n8683) );
  XNOR2_X1 U14241 ( .A(n8684), .B(n8683), .ZN(n8685) );
  XNOR2_X1 U14242 ( .A(n8686), .B(n8685), .ZN(n9429) );
  MUX2_X1 U14243 ( .A(n9221), .B(n9736), .S(n3799), .Z(n8712) );
  XNOR2_X1 U14244 ( .A(n8687), .B(n8952), .ZN(n8688) );
  XNOR2_X1 U14245 ( .A(n8689), .B(n8688), .ZN(n8695) );
  XNOR2_X1 U14246 ( .A(n9139), .B(n8690), .ZN(n8693) );
  XNOR2_X1 U14247 ( .A(n8691), .B(n2747), .ZN(n8692) );
  XNOR2_X1 U14248 ( .A(n8693), .B(n8692), .ZN(n8694) );
  INV_X1 U14250 ( .A(n9980), .ZN(n9984) );
  XNOR2_X1 U14251 ( .A(n8698), .B(n8962), .ZN(n8701) );
  XNOR2_X1 U14252 ( .A(n8699), .B(n1364), .ZN(n8700) );
  XNOR2_X1 U14253 ( .A(n8701), .B(n8700), .ZN(n8702) );
  MUX2_X1 U14254 ( .A(n9984), .B(n9982), .S(n9981), .Z(n8711) );
  INV_X1 U14255 ( .A(n8703), .ZN(n8705) );
  XNOR2_X1 U14256 ( .A(n8704), .B(n8705), .ZN(n8710) );
  XNOR2_X1 U14257 ( .A(n8897), .B(n8706), .ZN(n8708) );
  XNOR2_X1 U14258 ( .A(n9044), .B(n2970), .ZN(n8707) );
  XOR2_X1 U14259 ( .A(n8708), .B(n8707), .Z(n8709) );
  XNOR2_X2 U14260 ( .A(n8710), .B(n8709), .ZN(n9985) );
  XNOR2_X1 U14262 ( .A(n8714), .B(n8713), .ZN(n8718) );
  XNOR2_X1 U14263 ( .A(n8867), .B(n1815), .ZN(n8716) );
  XNOR2_X1 U14264 ( .A(n8716), .B(n8715), .ZN(n8717) );
  XNOR2_X1 U14265 ( .A(n8720), .B(n8719), .ZN(n8724) );
  XNOR2_X1 U14266 ( .A(n8723), .B(n8724), .ZN(n10069) );
  NOR2_X1 U14267 ( .A1(n427), .A2(n25457), .ZN(n9232) );
  INV_X1 U14268 ( .A(n10069), .ZN(n10075) );
  XNOR2_X1 U14269 ( .A(n8726), .B(n8725), .ZN(n8729) );
  XNOR2_X1 U14270 ( .A(n8760), .B(n812), .ZN(n8727) );
  XNOR2_X1 U14271 ( .A(n9042), .B(n8727), .ZN(n8728) );
  XNOR2_X1 U14272 ( .A(n8729), .B(n8728), .ZN(n8744) );
  INV_X1 U14273 ( .A(n8744), .ZN(n9620) );
  XNOR2_X1 U14274 ( .A(n8730), .B(n8951), .ZN(n8732) );
  XNOR2_X1 U14275 ( .A(n8731), .B(n8732), .ZN(n8736) );
  XNOR2_X1 U14276 ( .A(n9141), .B(n2036), .ZN(n8733) );
  XNOR2_X1 U14277 ( .A(n8734), .B(n8733), .ZN(n8735) );
  XNOR2_X1 U14278 ( .A(n8736), .B(n8735), .ZN(n10068) );
  INV_X1 U14279 ( .A(n10068), .ZN(n9764) );
  OAI21_X1 U14280 ( .B1(n10075), .B2(n9620), .A(n9764), .ZN(n8737) );
  NOR2_X1 U14281 ( .A1(n9232), .A2(n8737), .ZN(n8752) );
  NAND2_X1 U14282 ( .A1(n427), .A2(n10068), .ZN(n9766) );
  XNOR2_X1 U14283 ( .A(n8739), .B(n8738), .ZN(n8743) );
  XNOR2_X1 U14284 ( .A(n8965), .B(n3084), .ZN(n8740) );
  XNOR2_X1 U14285 ( .A(n8741), .B(n8740), .ZN(n8742) );
  XNOR2_X1 U14286 ( .A(n8746), .B(n1804), .ZN(n8747) );
  XOR2_X1 U14287 ( .A(n8748), .B(n8747), .Z(n8749) );
  NAND3_X1 U14288 ( .A1(n1330), .A2(n10070), .A3(n9762), .ZN(n8751) );
  XNOR2_X1 U14289 ( .A(n9191), .B(n24445), .ZN(n9050) );
  XNOR2_X1 U14290 ( .A(n9050), .B(n8753), .ZN(n8759) );
  XNOR2_X1 U14291 ( .A(n8754), .B(n3183), .ZN(n8757) );
  XNOR2_X1 U14292 ( .A(n8756), .B(n8757), .ZN(n8758) );
  XNOR2_X1 U14293 ( .A(n8759), .B(n8758), .ZN(n9419) );
  INV_X1 U14294 ( .A(n9419), .ZN(n9617) );
  XNOR2_X1 U14295 ( .A(n9043), .B(n8760), .ZN(n8763) );
  INV_X1 U14296 ( .A(n173), .ZN(n8761) );
  XNOR2_X1 U14297 ( .A(n8989), .B(n8761), .ZN(n8762) );
  XNOR2_X1 U14298 ( .A(n8763), .B(n8762), .ZN(n8768) );
  XNOR2_X1 U14299 ( .A(n9041), .B(n8764), .ZN(n8765) );
  XNOR2_X1 U14300 ( .A(n8766), .B(n8765), .ZN(n8767) );
  XNOR2_X1 U14301 ( .A(n8770), .B(n8769), .ZN(n9146) );
  XNOR2_X1 U14302 ( .A(n8771), .B(n8772), .ZN(n9000) );
  XNOR2_X1 U14303 ( .A(n9146), .B(n9000), .ZN(n8776) );
  XNOR2_X1 U14304 ( .A(n8964), .B(n9057), .ZN(n8774) );
  XNOR2_X1 U14305 ( .A(n8965), .B(n1924), .ZN(n8773) );
  XNOR2_X1 U14306 ( .A(n8774), .B(n8773), .ZN(n8775) );
  XNOR2_X1 U14307 ( .A(n8776), .B(n8775), .ZN(n9613) );
  MUX2_X1 U14308 ( .A(n9617), .B(n25005), .S(n9613), .Z(n8804) );
  XNOR2_X1 U14309 ( .A(n8778), .B(n8777), .ZN(n8785) );
  XNOR2_X1 U14310 ( .A(n8779), .B(n8780), .ZN(n9154) );
  XNOR2_X1 U14311 ( .A(n8782), .B(n8781), .ZN(n8783) );
  XNOR2_X1 U14312 ( .A(n9154), .B(n8783), .ZN(n8784) );
  XNOR2_X1 U14313 ( .A(n8786), .B(n3164), .ZN(n8788) );
  XNOR2_X1 U14314 ( .A(n8788), .B(n8787), .ZN(n8792) );
  XNOR2_X1 U14315 ( .A(n8790), .B(n8789), .ZN(n9177) );
  INV_X1 U14316 ( .A(n9177), .ZN(n8791) );
  XNOR2_X1 U14317 ( .A(n8791), .B(n8792), .ZN(n8794) );
  XNOR2_X1 U14318 ( .A(n8794), .B(n8793), .ZN(n9977) );
  INV_X1 U14319 ( .A(n9977), .ZN(n9757) );
  XNOR2_X1 U14320 ( .A(n9137), .B(n8797), .ZN(n8802) );
  INV_X1 U14321 ( .A(n2240), .ZN(n20864) );
  XNOR2_X1 U14322 ( .A(n8799), .B(n20864), .ZN(n8800) );
  XNOR2_X1 U14323 ( .A(n8997), .B(n8800), .ZN(n8801) );
  XNOR2_X1 U14324 ( .A(n8802), .B(n8801), .ZN(n9753) );
  INV_X1 U14325 ( .A(n9753), .ZN(n9974) );
  NAND3_X1 U14326 ( .A1(n9617), .A2(n9974), .A3(n25005), .ZN(n8803) );
  XNOR2_X1 U14327 ( .A(n8805), .B(n9089), .ZN(n8811) );
  XNOR2_X1 U14328 ( .A(n9158), .B(n1874), .ZN(n8809) );
  XNOR2_X1 U14329 ( .A(n8806), .B(n8807), .ZN(n8808) );
  XNOR2_X1 U14330 ( .A(n8809), .B(n8808), .ZN(n8810) );
  INV_X1 U14332 ( .A(n8970), .ZN(n9168) );
  XNOR2_X1 U14333 ( .A(n9168), .B(n8812), .ZN(n8815) );
  XNOR2_X1 U14334 ( .A(n8813), .B(Key[172]), .ZN(n8814) );
  XNOR2_X1 U14335 ( .A(n8815), .B(n8814), .ZN(n8817) );
  XNOR2_X1 U14336 ( .A(n8873), .B(n9096), .ZN(n8816) );
  NAND2_X1 U14337 ( .A1(n10020), .A2(n24495), .ZN(n9732) );
  INV_X1 U14338 ( .A(n9732), .ZN(n8842) );
  XNOR2_X1 U14339 ( .A(n8818), .B(n4034), .ZN(n8819) );
  XNOR2_X1 U14340 ( .A(n8858), .B(n8819), .ZN(n8823) );
  XNOR2_X1 U14341 ( .A(n8820), .B(n9176), .ZN(n8821) );
  XNOR2_X1 U14342 ( .A(n8821), .B(n9115), .ZN(n8822) );
  INV_X1 U14343 ( .A(n10018), .ZN(n9730) );
  XNOR2_X1 U14344 ( .A(n8824), .B(n9188), .ZN(n8825) );
  XNOR2_X1 U14345 ( .A(n9101), .B(n8825), .ZN(n8830) );
  XNOR2_X1 U14346 ( .A(n8826), .B(n23699), .ZN(n8828) );
  XNOR2_X1 U14347 ( .A(n8828), .B(n8827), .ZN(n8829) );
  XNOR2_X1 U14348 ( .A(n8830), .B(n8829), .ZN(n8839) );
  XNOR2_X1 U14349 ( .A(n8951), .B(n21703), .ZN(n8832) );
  XNOR2_X1 U14350 ( .A(n8832), .B(n8831), .ZN(n8834) );
  XNOR2_X1 U14351 ( .A(n8833), .B(n8834), .ZN(n10019) );
  INV_X1 U14352 ( .A(n10019), .ZN(n9320) );
  OAI211_X1 U14353 ( .C1(n9729), .C2(n9730), .A(n8839), .B(n9320), .ZN(n8841)
         );
  INV_X1 U14354 ( .A(n9729), .ZN(n9493) );
  XNOR2_X1 U14355 ( .A(n8961), .B(n1952), .ZN(n8836) );
  XNOR2_X1 U14356 ( .A(n9111), .B(n8836), .ZN(n8837) );
  INV_X1 U14357 ( .A(n8839), .ZN(n9731) );
  XNOR2_X1 U14358 ( .A(n8843), .B(n8844), .ZN(n8850) );
  XNOR2_X1 U14359 ( .A(n8846), .B(n8845), .ZN(n8848) );
  XNOR2_X1 U14360 ( .A(n8917), .B(n2989), .ZN(n8847) );
  XNOR2_X1 U14361 ( .A(n8848), .B(n8847), .ZN(n8849) );
  XNOR2_X1 U14362 ( .A(n8850), .B(n8849), .ZN(n9634) );
  XNOR2_X1 U14363 ( .A(n8852), .B(n8851), .ZN(n8857) );
  XNOR2_X1 U14364 ( .A(n8853), .B(n921), .ZN(n8854) );
  XNOR2_X1 U14365 ( .A(n8855), .B(n8854), .ZN(n8856) );
  XNOR2_X1 U14366 ( .A(n8857), .B(n8856), .ZN(n9435) );
  XNOR2_X1 U14368 ( .A(n8858), .B(n8859), .ZN(n8864) );
  XNOR2_X1 U14369 ( .A(n8860), .B(n2745), .ZN(n8861) );
  XNOR2_X1 U14370 ( .A(n8862), .B(n8861), .ZN(n8863) );
  XNOR2_X1 U14371 ( .A(n8864), .B(n8863), .ZN(n9711) );
  OR2_X1 U14372 ( .A1(n10038), .A2(n9711), .ZN(n8888) );
  XNOR2_X1 U14373 ( .A(n8866), .B(n8865), .ZN(n8871) );
  XNOR2_X1 U14374 ( .A(n8867), .B(n899), .ZN(n8869) );
  XNOR2_X1 U14375 ( .A(n8868), .B(n8869), .ZN(n8870) );
  XNOR2_X1 U14376 ( .A(n8873), .B(n8872), .ZN(n8879) );
  XNOR2_X1 U14377 ( .A(n8874), .B(n24056), .ZN(n8877) );
  XNOR2_X1 U14378 ( .A(n8875), .B(n4189), .ZN(n8876) );
  XNOR2_X1 U14379 ( .A(n8877), .B(n8876), .ZN(n8878) );
  XNOR2_X1 U14380 ( .A(n8879), .B(n8878), .ZN(n10037) );
  NOR2_X1 U14381 ( .A1(n9635), .A2(n10037), .ZN(n9228) );
  NAND2_X1 U14382 ( .A1(n9228), .A2(n9713), .ZN(n8887) );
  INV_X1 U14383 ( .A(n9634), .ZN(n9718) );
  XNOR2_X1 U14384 ( .A(n8880), .B(n1854), .ZN(n8881) );
  XNOR2_X1 U14385 ( .A(n8883), .B(n8882), .ZN(n8885) );
  INV_X1 U14387 ( .A(n9433), .ZN(n9710) );
  INV_X1 U14388 ( .A(n9090), .ZN(n8890) );
  XNOR2_X1 U14389 ( .A(n8890), .B(n8889), .ZN(n8895) );
  XNOR2_X1 U14390 ( .A(n9034), .B(n25235), .ZN(n8893) );
  XNOR2_X1 U14391 ( .A(n8891), .B(n2805), .ZN(n8892) );
  XNOR2_X1 U14392 ( .A(n8893), .B(n8892), .ZN(n8894) );
  XNOR2_X1 U14393 ( .A(n8897), .B(n8896), .ZN(n9098) );
  XNOR2_X1 U14394 ( .A(n8899), .B(n8898), .ZN(n8986) );
  XNOR2_X1 U14395 ( .A(n9098), .B(n8986), .ZN(n8905) );
  XNOR2_X1 U14396 ( .A(n25228), .B(n8987), .ZN(n8903) );
  XNOR2_X1 U14398 ( .A(n24056), .B(n24280), .ZN(n8902) );
  XNOR2_X1 U14399 ( .A(n8903), .B(n8902), .ZN(n8904) );
  XNOR2_X2 U14400 ( .A(n8905), .B(n8904), .ZN(n9990) );
  INV_X1 U14401 ( .A(n9990), .ZN(n9996) );
  XNOR2_X1 U14402 ( .A(n9058), .B(n1726), .ZN(n8906) );
  XNOR2_X1 U14403 ( .A(n8907), .B(n8906), .ZN(n8912) );
  XNOR2_X1 U14404 ( .A(n8908), .B(n8909), .ZN(n8910) );
  XNOR2_X1 U14405 ( .A(n9110), .B(n8910), .ZN(n8911) );
  XNOR2_X1 U14406 ( .A(n8913), .B(n8914), .ZN(n8915) );
  XNOR2_X1 U14407 ( .A(n9122), .B(n8915), .ZN(n8921) );
  XNOR2_X1 U14408 ( .A(n9081), .B(n8916), .ZN(n8919) );
  XNOR2_X1 U14409 ( .A(n8917), .B(n21964), .ZN(n8918) );
  XNOR2_X1 U14410 ( .A(n8919), .B(n8918), .ZN(n8920) );
  XNOR2_X1 U14411 ( .A(n8921), .B(n8920), .ZN(n9658) );
  INV_X1 U14412 ( .A(n9658), .ZN(n9745) );
  AOI21_X1 U14413 ( .B1(n9745), .B2(n9989), .A(n9990), .ZN(n9316) );
  XNOR2_X1 U14414 ( .A(n8922), .B(n9011), .ZN(n8927) );
  XNOR2_X1 U14415 ( .A(n9075), .B(n21742), .ZN(n8924) );
  XNOR2_X1 U14416 ( .A(n8924), .B(n8923), .ZN(n8925) );
  XNOR2_X1 U14417 ( .A(n9010), .B(n8925), .ZN(n8926) );
  XNOR2_X1 U14418 ( .A(n8926), .B(n8927), .ZN(n9423) );
  XNOR2_X1 U14419 ( .A(n9102), .B(n9020), .ZN(n8932) );
  XNOR2_X1 U14420 ( .A(n8928), .B(n8880), .ZN(n8930) );
  XNOR2_X1 U14421 ( .A(n8935), .B(n3152), .ZN(n8929) );
  XNOR2_X1 U14422 ( .A(n8930), .B(n8929), .ZN(n8931) );
  XNOR2_X2 U14423 ( .A(n8932), .B(n8931), .ZN(n9991) );
  OAI211_X1 U14424 ( .C1(n25444), .C2(n9990), .A(n9657), .B(n9747), .ZN(n8933)
         );
  OAI21_X1 U14425 ( .B1(n9425), .B2(n9316), .A(n8933), .ZN(n11519) );
  INV_X1 U14426 ( .A(n25060), .ZN(n10384) );
  XNOR2_X1 U14427 ( .A(n8935), .B(n2049), .ZN(n8936) );
  XNOR2_X1 U14428 ( .A(n8940), .B(n8941), .ZN(n8944) );
  XNOR2_X1 U14429 ( .A(n9176), .B(n1870), .ZN(n8942) );
  XNOR2_X1 U14430 ( .A(n9011), .B(n8942), .ZN(n8943) );
  XNOR2_X1 U14431 ( .A(n9158), .B(n1951), .ZN(n8946) );
  XNOR2_X1 U14432 ( .A(n8946), .B(n25235), .ZN(n8948) );
  XNOR2_X1 U14433 ( .A(n8948), .B(n8947), .ZN(n8949) );
  INV_X1 U14434 ( .A(n9550), .ZN(n9682) );
  MUX2_X1 U14435 ( .A(n260), .B(n10046), .S(n9682), .Z(n8979) );
  XNOR2_X1 U14436 ( .A(n8952), .B(n8951), .ZN(n8954) );
  XNOR2_X1 U14437 ( .A(n8954), .B(n8953), .ZN(n8958) );
  XNOR2_X1 U14438 ( .A(n9139), .B(n3093), .ZN(n8956) );
  XNOR2_X1 U14439 ( .A(n8956), .B(n8955), .ZN(n8957) );
  XNOR2_X1 U14440 ( .A(n8960), .B(n8959), .ZN(n8963) );
  XNOR2_X1 U14441 ( .A(n8962), .B(n8961), .ZN(n9144) );
  XNOR2_X1 U14442 ( .A(n9144), .B(n8963), .ZN(n8969) );
  XNOR2_X1 U14443 ( .A(n9059), .B(n8964), .ZN(n8967) );
  XNOR2_X1 U14444 ( .A(n8965), .B(n2717), .ZN(n8966) );
  XNOR2_X1 U14445 ( .A(n8967), .B(n8966), .ZN(n8968) );
  XNOR2_X1 U14446 ( .A(n8969), .B(n8968), .ZN(n10045) );
  INV_X1 U14447 ( .A(n10045), .ZN(n9627) );
  AND2_X1 U14448 ( .A1(n261), .A2(n9627), .ZN(n9684) );
  XNOR2_X1 U14449 ( .A(n8970), .B(n765), .ZN(n8972) );
  XNOR2_X1 U14450 ( .A(n8971), .B(n8972), .ZN(n8975) );
  XNOR2_X1 U14451 ( .A(n8987), .B(n8973), .ZN(n8974) );
  XNOR2_X1 U14452 ( .A(n8975), .B(n8974), .ZN(n8976) );
  MUX2_X2 U14453 ( .A(n8979), .B(n8978), .S(n9681), .Z(n11038) );
  INV_X1 U14454 ( .A(n11038), .ZN(n10570) );
  XNOR2_X1 U14455 ( .A(n8985), .B(n8986), .ZN(n8993) );
  XNOR2_X1 U14456 ( .A(n8987), .B(n8988), .ZN(n8991) );
  XNOR2_X1 U14457 ( .A(n8989), .B(n24287), .ZN(n8990) );
  XNOR2_X1 U14458 ( .A(n8991), .B(n8990), .ZN(n8992) );
  INV_X1 U14459 ( .A(n9696), .ZN(n9699) );
  XNOR2_X1 U14460 ( .A(n8994), .B(n8995), .ZN(n8999) );
  XNOR2_X1 U14461 ( .A(n8997), .B(n8996), .ZN(n8998) );
  XNOR2_X1 U14462 ( .A(n8998), .B(n8999), .ZN(n10029) );
  INV_X1 U14463 ( .A(n10029), .ZN(n9695) );
  XNOR2_X1 U14464 ( .A(n9000), .B(n9001), .ZN(n9006) );
  XNOR2_X1 U14465 ( .A(n9002), .B(n2795), .ZN(n9004) );
  XNOR2_X1 U14466 ( .A(n9003), .B(n9004), .ZN(n9005) );
  NOR2_X1 U14467 ( .A1(n9639), .A2(n24332), .ZN(n10028) );
  XNOR2_X1 U14468 ( .A(n9007), .B(n2882), .ZN(n9008) );
  XNOR2_X1 U14469 ( .A(n9010), .B(n9009), .ZN(n9014) );
  XNOR2_X1 U14470 ( .A(n9012), .B(n9011), .ZN(n9013) );
  INV_X1 U14471 ( .A(n9016), .ZN(n9017) );
  XNOR2_X1 U14472 ( .A(n9018), .B(n9017), .ZN(n9019) );
  INV_X1 U14473 ( .A(n10026), .ZN(n9022) );
  OAI211_X1 U14474 ( .C1(n9699), .C2(n10027), .A(n10031), .B(n9022), .ZN(n9023) );
  OAI21_X1 U14475 ( .B1(n9565), .B2(n9563), .A(n9024), .ZN(n9026) );
  OAI21_X1 U14476 ( .B1(n9454), .B2(n9885), .A(n9567), .ZN(n9025) );
  AOI21_X1 U14477 ( .B1(n10570), .B2(n10944), .A(n10942), .ZN(n9131) );
  NAND3_X1 U14478 ( .A1(n4993), .A2(n9872), .A3(n9875), .ZN(n9031) );
  NAND2_X1 U14479 ( .A1(n9694), .A2(n9028), .ZN(n9030) );
  NAND3_X1 U14480 ( .A1(n9875), .A2(n307), .A3(n9251), .ZN(n9029) );
  XNOR2_X1 U14482 ( .A(n9033), .B(n9154), .ZN(n9039) );
  XNOR2_X1 U14483 ( .A(n9035), .B(n1792), .ZN(n9036) );
  XNOR2_X1 U14484 ( .A(n9037), .B(n9036), .ZN(n9038) );
  XNOR2_X1 U14485 ( .A(n9040), .B(n9041), .ZN(n9164) );
  XNOR2_X1 U14486 ( .A(n9164), .B(n9042), .ZN(n9049) );
  XNOR2_X1 U14487 ( .A(n9043), .B(n62), .ZN(n9047) );
  XNOR2_X1 U14488 ( .A(n25228), .B(n9044), .ZN(n9046) );
  XNOR2_X1 U14489 ( .A(n9047), .B(n9046), .ZN(n9048) );
  XNOR2_X1 U14490 ( .A(n9049), .B(n9048), .ZN(n9244) );
  XNOR2_X1 U14492 ( .A(n9051), .B(n9050), .ZN(n9056) );
  XNOR2_X1 U14493 ( .A(n8880), .B(n2903), .ZN(n9053) );
  XNOR2_X1 U14494 ( .A(n9054), .B(n9053), .ZN(n9055) );
  NAND2_X1 U14495 ( .A1(n10058), .A2(n24092), .ZN(n9063) );
  XNOR2_X1 U14496 ( .A(n9058), .B(n9057), .ZN(n9061) );
  XNOR2_X1 U14497 ( .A(n9059), .B(n1801), .ZN(n9060) );
  XNOR2_X2 U14498 ( .A(n9062), .B(n5743), .ZN(n10053) );
  XNOR2_X1 U14499 ( .A(n9065), .B(n9177), .ZN(n9079) );
  MUX2_X1 U14500 ( .A(n9068), .B(n9067), .S(n9066), .Z(n9072) );
  OAI211_X1 U14501 ( .C1(n9072), .C2(n9071), .A(n9070), .B(n9069), .ZN(n9074)
         );
  XNOR2_X1 U14502 ( .A(n9074), .B(n9073), .ZN(n9077) );
  XNOR2_X1 U14503 ( .A(n9075), .B(n2044), .ZN(n9076) );
  XNOR2_X1 U14504 ( .A(n9077), .B(n9076), .ZN(n9078) );
  XNOR2_X1 U14505 ( .A(n9137), .B(n9080), .ZN(n9085) );
  XNOR2_X1 U14506 ( .A(n9081), .B(n9141), .ZN(n9084) );
  XNOR2_X1 U14507 ( .A(n9082), .B(n2782), .ZN(n9083) );
  MUX2_X1 U14508 ( .A(n9539), .B(n9086), .S(n9244), .Z(n9087) );
  XNOR2_X1 U14509 ( .A(n9089), .B(n9090), .ZN(n9094) );
  XNOR2_X1 U14510 ( .A(n8069), .B(n1835), .ZN(n9091) );
  XNOR2_X1 U14511 ( .A(n9092), .B(n9091), .ZN(n9093) );
  XNOR2_X1 U14512 ( .A(n9096), .B(n9095), .ZN(n9100) );
  XNOR2_X1 U14513 ( .A(n9169), .B(n1920), .ZN(n9097) );
  XNOR2_X1 U14514 ( .A(n9098), .B(n9097), .ZN(n9099) );
  XNOR2_X1 U14515 ( .A(n9100), .B(n9099), .ZN(n9218) );
  NAND2_X1 U14516 ( .A1(n10060), .A2(n10065), .ZN(n9703) );
  XNOR2_X1 U14517 ( .A(n9102), .B(n9101), .ZN(n9105) );
  XNOR2_X1 U14518 ( .A(n9189), .B(n3073), .ZN(n9103) );
  XNOR2_X1 U14519 ( .A(n8297), .B(n9103), .ZN(n9104) );
  XNOR2_X1 U14520 ( .A(n9106), .B(n9107), .ZN(n9109) );
  XNOR2_X1 U14521 ( .A(n9149), .B(n2208), .ZN(n9108) );
  XNOR2_X1 U14522 ( .A(n9109), .B(n9108), .ZN(n9113) );
  XNOR2_X1 U14523 ( .A(n9110), .B(n9111), .ZN(n9112) );
  NAND2_X1 U14524 ( .A1(n9127), .A2(n9704), .ZN(n9120) );
  XNOR2_X1 U14525 ( .A(n9179), .B(n2477), .ZN(n9116) );
  XNOR2_X1 U14526 ( .A(n9117), .B(n9116), .ZN(n9118) );
  XNOR2_X1 U14527 ( .A(n9119), .B(n9118), .ZN(n10061) );
  AOI21_X1 U14528 ( .B1(n9703), .B2(n9120), .A(n309), .ZN(n9129) );
  XNOR2_X1 U14529 ( .A(n9121), .B(n2991), .ZN(n9123) );
  XNOR2_X1 U14530 ( .A(n9122), .B(n9123), .ZN(n9126) );
  XNOR2_X1 U14531 ( .A(n9125), .B(n9126), .ZN(n10063) );
  INV_X1 U14533 ( .A(n9460), .ZN(n9919) );
  INV_X1 U14534 ( .A(n9459), .ZN(n9271) );
  INV_X1 U14535 ( .A(n9918), .ZN(n9914) );
  INV_X1 U14536 ( .A(n9463), .ZN(n9916) );
  NOR2_X1 U14538 ( .A1(n10583), .A2(n10371), .ZN(n9210) );
  XNOR2_X1 U14539 ( .A(n9140), .B(n9139), .ZN(n9143) );
  INV_X1 U14542 ( .A(n9144), .ZN(n9145) );
  XNOR2_X1 U14543 ( .A(n9145), .B(n9146), .ZN(n9153) );
  XNOR2_X1 U14544 ( .A(n9147), .B(n8484), .ZN(n9151) );
  XNOR2_X1 U14545 ( .A(n9149), .B(n1865), .ZN(n9150) );
  XNOR2_X1 U14546 ( .A(n9151), .B(n9150), .ZN(n9152) );
  INV_X1 U14547 ( .A(n24025), .ZN(n10140) );
  NOR2_X1 U14548 ( .A1(n10146), .A2(n10140), .ZN(n9187) );
  INV_X1 U14549 ( .A(n9154), .ZN(n9157) );
  XNOR2_X1 U14550 ( .A(n9155), .B(n8069), .ZN(n9156) );
  XNOR2_X1 U14551 ( .A(n9157), .B(n9156), .ZN(n9163) );
  XNOR2_X1 U14552 ( .A(n9159), .B(n9158), .ZN(n9161) );
  XNOR2_X1 U14553 ( .A(n8278), .B(n2726), .ZN(n9160) );
  XNOR2_X1 U14554 ( .A(n9161), .B(n9160), .ZN(n9162) );
  INV_X1 U14555 ( .A(n9164), .ZN(n9166) );
  XNOR2_X1 U14556 ( .A(n9165), .B(n9166), .ZN(n9173) );
  XNOR2_X1 U14557 ( .A(n9167), .B(n9168), .ZN(n9171) );
  XNOR2_X1 U14558 ( .A(n9169), .B(n1746), .ZN(n9170) );
  XNOR2_X1 U14559 ( .A(n9171), .B(n9170), .ZN(n9172) );
  INV_X1 U14562 ( .A(n9174), .ZN(n9397) );
  XNOR2_X1 U14563 ( .A(n9175), .B(n9176), .ZN(n9178) );
  XNOR2_X1 U14564 ( .A(n9177), .B(n9178), .ZN(n9186) );
  INV_X1 U14565 ( .A(n9179), .ZN(n9180) );
  XNOR2_X1 U14566 ( .A(n9181), .B(n9180), .ZN(n9184) );
  INV_X1 U14567 ( .A(n22986), .ZN(n20805) );
  XNOR2_X1 U14568 ( .A(n9182), .B(n20805), .ZN(n9183) );
  XNOR2_X1 U14569 ( .A(n9184), .B(n9183), .ZN(n9185) );
  XNOR2_X1 U14570 ( .A(n9186), .B(n9185), .ZN(n9820) );
  XNOR2_X1 U14571 ( .A(n9189), .B(n9188), .ZN(n9193) );
  XNOR2_X1 U14572 ( .A(n9190), .B(n9191), .ZN(n9192) );
  XNOR2_X1 U14573 ( .A(n9193), .B(n9192), .ZN(n9200) );
  XNOR2_X1 U14574 ( .A(n9194), .B(n24445), .ZN(n9198) );
  XNOR2_X1 U14575 ( .A(n9196), .B(n5131), .ZN(n9197) );
  XNOR2_X1 U14576 ( .A(n9198), .B(n9197), .ZN(n9199) );
  NOR2_X1 U14578 ( .A1(n10584), .A2(n10585), .ZN(n9209) );
  INV_X1 U14579 ( .A(n25216), .ZN(n9928) );
  NAND2_X1 U14580 ( .A1(n9930), .A2(n9928), .ZN(n9208) );
  INV_X1 U14581 ( .A(n9345), .ZN(n9600) );
  NAND2_X1 U14586 ( .A1(n2565), .A2(n10254), .ZN(n10252) );
  NAND2_X1 U14587 ( .A1(n10250), .A2(n9372), .ZN(n9213) );
  INV_X1 U14589 ( .A(n9218), .ZN(n9705) );
  NAND2_X1 U14590 ( .A1(n309), .A2(n9705), .ZN(n9219) );
  NAND2_X1 U14591 ( .A1(n9221), .A2(n9985), .ZN(n9225) );
  NAND3_X1 U14592 ( .A1(n9984), .A2(n9742), .A3(n9981), .ZN(n9223) );
  OAI21_X1 U14593 ( .B1(n9664), .B2(n9982), .A(n9736), .ZN(n9222) );
  NOR2_X1 U14594 ( .A1(n9635), .A2(n9435), .ZN(n9227) );
  INV_X1 U14595 ( .A(n10037), .ZN(n9633) );
  NOR2_X1 U14596 ( .A1(n9634), .A2(n9633), .ZN(n9226) );
  MUX2_X1 U14597 ( .A(n9227), .B(n9226), .S(n9433), .Z(n9230) );
  INV_X1 U14598 ( .A(n9228), .ZN(n9229) );
  INV_X1 U14599 ( .A(n9435), .ZN(n9709) );
  MUX2_X1 U14600 ( .A(n9231), .B(n10068), .S(n10075), .Z(n9235) );
  INV_X1 U14601 ( .A(n9232), .ZN(n9234) );
  AOI21_X1 U14602 ( .B1(n427), .B2(n10072), .A(n9620), .ZN(n9233) );
  INV_X1 U14604 ( .A(n10848), .ZN(n11125) );
  INV_X1 U14605 ( .A(n10027), .ZN(n9240) );
  AOI21_X1 U14606 ( .B1(n9697), .B2(n10026), .A(n10029), .ZN(n9238) );
  OR2_X1 U14607 ( .A1(n9238), .A2(n9639), .ZN(n9239) );
  NAND2_X1 U14608 ( .A1(n11121), .A2(n11123), .ZN(n10847) );
  INV_X1 U14609 ( .A(n10847), .ZN(n9241) );
  NAND2_X1 U14610 ( .A1(n24446), .A2(n10050), .ZN(n9867) );
  INV_X1 U14611 ( .A(n9245), .ZN(n9246) );
  INV_X1 U14612 ( .A(n9564), .ZN(n9456) );
  INV_X1 U14613 ( .A(n9565), .ZN(n9883) );
  NAND2_X1 U14614 ( .A1(n9883), .A2(n9885), .ZN(n9249) );
  MUX2_X1 U14615 ( .A(n9249), .B(n9248), .S(n9887), .Z(n9250) );
  INV_X1 U14616 ( .A(n9255), .ZN(n9628) );
  AOI22_X1 U14617 ( .A1(n9682), .A2(n9681), .B1(n9628), .B2(n10045), .ZN(n9257) );
  NAND2_X1 U14618 ( .A1(n261), .A2(n9681), .ZN(n9256) );
  MUX2_X1 U14619 ( .A(n9257), .B(n9256), .S(n10046), .Z(n9258) );
  INV_X1 U14620 ( .A(n10740), .ZN(n10856) );
  NAND2_X1 U14621 ( .A1(n10856), .A2(n10861), .ZN(n10743) );
  INV_X1 U14622 ( .A(n9864), .ZN(n9559) );
  INV_X1 U14623 ( .A(n9554), .ZN(n9860) );
  INV_X1 U14624 ( .A(n9560), .ZN(n9858) );
  NAND2_X1 U14625 ( .A1(n9857), .A2(n9860), .ZN(n9260) );
  INV_X1 U14626 ( .A(n9856), .ZN(n9474) );
  NAND2_X1 U14627 ( .A1(n9474), .A2(n9858), .ZN(n9259) );
  MUX2_X1 U14628 ( .A(n9260), .B(n9259), .S(n9864), .Z(n9261) );
  NAND3_X1 U14629 ( .A1(n10740), .A2(n10737), .A3(n10858), .ZN(n9267) );
  AOI21_X1 U14630 ( .B1(n9942), .B2(n25021), .A(n227), .ZN(n9265) );
  NOR2_X1 U14631 ( .A1(n9893), .A2(n9943), .ZN(n9263) );
  OAI21_X1 U14632 ( .B1(n9289), .B2(n9263), .A(n9897), .ZN(n9264) );
  AND2_X1 U14633 ( .A1(n25229), .A2(n10737), .ZN(n10862) );
  NAND2_X1 U14634 ( .A1(n10862), .A2(n10190), .ZN(n9266) );
  NAND4_X2 U14635 ( .A1(n9268), .A2(n9266), .A3(n10743), .A4(n9267), .ZN(
        n12364) );
  XNOR2_X1 U14636 ( .A(n12364), .B(n12089), .ZN(n11734) );
  INV_X1 U14638 ( .A(n9269), .ZN(n9952) );
  INV_X1 U14639 ( .A(n9388), .ZN(n9948) );
  OAI21_X1 U14640 ( .B1(n9389), .B2(n9388), .A(n9952), .ZN(n9270) );
  INV_X1 U14641 ( .A(n10192), .ZN(n10831) );
  INV_X1 U14642 ( .A(n9462), .ZN(n9354) );
  NAND2_X1 U14643 ( .A1(n9354), .A2(n9459), .ZN(n9458) );
  NAND3_X1 U14644 ( .A1(n9354), .A2(n9271), .A3(n9461), .ZN(n9273) );
  NAND3_X1 U14645 ( .A1(n24944), .A2(n9271), .A3(n9355), .ZN(n9272) );
  NAND4_X1 U14646 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n10277) );
  AND2_X1 U14647 ( .A1(n10277), .A2(n10831), .ZN(n10834) );
  INV_X1 U14648 ( .A(n9449), .ZN(n9906) );
  INV_X1 U14649 ( .A(n9907), .ZN(n9904) );
  MUX2_X1 U14650 ( .A(n9906), .B(n9904), .S(n9276), .Z(n9278) );
  MUX2_X1 U14651 ( .A(n9939), .B(n9276), .S(n9905), .Z(n9277) );
  NAND2_X1 U14652 ( .A1(n10834), .A2(n9279), .ZN(n9293) );
  INV_X1 U14653 ( .A(n9857), .ZN(n9555) );
  NAND2_X1 U14654 ( .A1(n9555), .A2(n9558), .ZN(n9280) );
  NAND3_X1 U14655 ( .A1(n3292), .A2(n9468), .A3(n9964), .ZN(n9284) );
  NAND2_X1 U14656 ( .A1(n9469), .A2(n9468), .ZN(n9282) );
  INV_X1 U14657 ( .A(n9944), .ZN(n9285) );
  OAI22_X1 U14658 ( .A1(n9288), .A2(n9287), .B1(n9286), .B2(n227), .ZN(n9290)
         );
  NOR2_X2 U14659 ( .A1(n9290), .A2(n9289), .ZN(n10518) );
  INV_X1 U14661 ( .A(n10275), .ZN(n10833) );
  OAI22_X1 U14662 ( .A1(n10090), .A2(n24505), .B1(n9295), .B2(n25454), .ZN(
        n9296) );
  AND2_X1 U14664 ( .A1(n9781), .A2(n10093), .ZN(n9498) );
  NOR2_X1 U14665 ( .A1(n9652), .A2(n9299), .ZN(n9653) );
  NOR2_X1 U14666 ( .A1(n9725), .A2(n25043), .ZN(n9300) );
  MUX2_X1 U14667 ( .A(n9653), .B(n9300), .S(n10008), .Z(n9304) );
  INV_X1 U14668 ( .A(n10007), .ZN(n9721) );
  MUX2_X1 U14669 ( .A(n9721), .B(n10008), .S(n9301), .Z(n9302) );
  NOR2_X1 U14670 ( .A1(n9302), .A2(n2922), .ZN(n9303) );
  INV_X1 U14673 ( .A(n10080), .ZN(n9326) );
  NAND3_X1 U14674 ( .A1(n4256), .A2(n10079), .A3(n9306), .ZN(n9308) );
  NAND4_X1 U14675 ( .A1(n9309), .A2(n10087), .A3(n9308), .A4(n9307), .ZN(
        n11130) );
  OAI21_X1 U14676 ( .B1(n9796), .B2(n8521), .A(n1796), .ZN(n9313) );
  NAND2_X1 U14677 ( .A1(n9671), .A2(n246), .ZN(n9668) );
  INV_X1 U14678 ( .A(n10714), .ZN(n10839) );
  OAI21_X1 U14679 ( .B1(n9657), .B2(n9747), .A(n9745), .ZN(n9315) );
  NAND2_X1 U14680 ( .A1(n9315), .A2(n24534), .ZN(n9317) );
  NOR2_X1 U14681 ( .A1(n10019), .A2(n25475), .ZN(n9319) );
  NOR2_X1 U14682 ( .A1(n9729), .A2(n24495), .ZN(n9318) );
  MUX2_X1 U14684 ( .A(n9319), .B(n9318), .S(n25007), .Z(n9323) );
  NAND2_X1 U14685 ( .A1(n10020), .A2(n9731), .ZN(n9321) );
  AOI21_X1 U14687 ( .B1(n9321), .B2(n10015), .A(n9320), .ZN(n9322) );
  INV_X1 U14688 ( .A(n10470), .ZN(n11129) );
  XNOR2_X1 U14689 ( .A(n24328), .B(n11356), .ZN(n9409) );
  OAI21_X1 U14690 ( .B1(n4256), .B2(n9507), .A(n9326), .ZN(n9325) );
  NOR2_X1 U14693 ( .A1(n9774), .A2(n4254), .ZN(n9329) );
  INV_X1 U14694 ( .A(n9773), .ZN(n9503) );
  INV_X1 U14698 ( .A(n10113), .ZN(n9529) );
  NAND2_X1 U14699 ( .A1(n9529), .A2(n8523), .ZN(n9336) );
  INV_X1 U14700 ( .A(n9805), .ZN(n10112) );
  MUX2_X1 U14701 ( .A(n9336), .B(n9335), .S(n10112), .Z(n10873) );
  NOR2_X1 U14702 ( .A1(n9806), .A2(n9530), .ZN(n9337) );
  INV_X1 U14703 ( .A(n9845), .ZN(n10156) );
  AND2_X1 U14708 ( .A1(n9384), .A2(n10161), .ZN(n10159) );
  OAI21_X1 U14709 ( .B1(n10159), .B2(n9349), .A(n3305), .ZN(n9350) );
  NOR2_X1 U14712 ( .A1(n9950), .A2(n9951), .ZN(n9363) );
  NAND2_X1 U14713 ( .A1(n9389), .A2(n9388), .ZN(n9362) );
  NAND2_X1 U14714 ( .A1(n9955), .A2(n9951), .ZN(n9359) );
  NAND2_X1 U14715 ( .A1(n9360), .A2(n9359), .ZN(n9361) );
  INV_X1 U14716 ( .A(n9365), .ZN(n9368) );
  NAND2_X1 U14719 ( .A1(n9365), .A2(n24025), .ZN(n9366) );
  INV_X1 U14720 ( .A(n10137), .ZN(n10134) );
  NAND3_X1 U14721 ( .A1(n9368), .A2(n25463), .A3(n10136), .ZN(n9369) );
  OR2_X1 U14722 ( .A1(n9380), .A2(n10128), .ZN(n9373) );
  INV_X1 U14723 ( .A(n10129), .ZN(n10132) );
  NAND2_X1 U14724 ( .A1(n10756), .A2(n10757), .ZN(n9374) );
  INV_X1 U14725 ( .A(n12249), .ZN(n9376) );
  XNOR2_X1 U14726 ( .A(n25090), .B(n9376), .ZN(n9407) );
  NAND2_X1 U14727 ( .A1(n9378), .A2(n9377), .ZN(n9381) );
  INV_X1 U14728 ( .A(n10729), .ZN(n10731) );
  NOR2_X1 U14729 ( .A1(n3305), .A2(n10157), .ZN(n9383) );
  INV_X1 U14730 ( .A(n10175), .ZN(n9585) );
  NAND2_X1 U14731 ( .A1(n9830), .A2(n9585), .ZN(n9386) );
  NAND2_X1 U14732 ( .A1(n9387), .A2(n9947), .ZN(n9391) );
  NOR2_X1 U14733 ( .A1(n9950), .A2(n9388), .ZN(n9390) );
  INV_X1 U14734 ( .A(n10734), .ZN(n10271) );
  INV_X1 U14735 ( .A(n9603), .ZN(n9926) );
  OAI211_X1 U14736 ( .C1(n9926), .C2(n9604), .A(n9600), .B(n9934), .ZN(n9396)
         );
  NAND2_X1 U14737 ( .A1(n25217), .A2(n9604), .ZN(n9395) );
  NAND3_X1 U14738 ( .A1(n9925), .A2(n24084), .A3(n9599), .ZN(n9394) );
  NAND3_X1 U14739 ( .A1(n10271), .A2(n4951), .A3(n10482), .ZN(n9405) );
  INV_X1 U14740 ( .A(n9398), .ZN(n10142) );
  NAND3_X1 U14741 ( .A1(n10146), .A2(n10142), .A3(n10134), .ZN(n9399) );
  OAI21_X1 U14742 ( .B1(n9174), .B2(n10140), .A(n9399), .ZN(n9402) );
  NOR2_X1 U14743 ( .A1(n10142), .A2(n24026), .ZN(n9400) );
  AOI21_X1 U14744 ( .B1(n10291), .B2(n10757), .A(n10753), .ZN(n9410) );
  NAND2_X1 U14745 ( .A1(n9760), .A2(n427), .ZN(n9412) );
  AOI21_X1 U14746 ( .B1(n9704), .B2(n429), .A(n10063), .ZN(n9414) );
  NAND2_X1 U14747 ( .A1(n9417), .A2(n9416), .ZN(n9422) );
  NAND2_X1 U14748 ( .A1(n9418), .A2(n9754), .ZN(n9421) );
  NAND2_X1 U14749 ( .A1(n9617), .A2(n9753), .ZN(n9751) );
  AND2_X1 U14750 ( .A1(n9972), .A2(n9752), .ZN(n9420) );
  NAND2_X1 U14751 ( .A1(n11084), .A2(n10890), .ZN(n9428) );
  NOR2_X1 U14752 ( .A1(n9991), .A2(n9747), .ZN(n9424) );
  OAI21_X1 U14753 ( .B1(n9425), .B2(n9424), .A(n9746), .ZN(n9427) );
  AND2_X1 U14754 ( .A1(n9423), .A2(n9990), .ZN(n9993) );
  OAI21_X1 U14755 ( .B1(n9993), .B2(n9745), .A(n9991), .ZN(n9426) );
  NAND2_X1 U14756 ( .A1(n9427), .A2(n9426), .ZN(n10889) );
  AOI21_X1 U14757 ( .B1(n11082), .B2(n9428), .A(n418), .ZN(n9439) );
  INV_X1 U14758 ( .A(n9985), .ZN(n9978) );
  NAND2_X1 U14759 ( .A1(n10890), .A2(n418), .ZN(n10441) );
  INV_X1 U14760 ( .A(n9635), .ZN(n9434) );
  INV_X1 U14761 ( .A(n10439), .ZN(n9437) );
  OAI22_X1 U14762 ( .A1(n10891), .A2(n10441), .B1(n9437), .B2(n10767), .ZN(
        n9438) );
  XNOR2_X1 U14763 ( .A(n11295), .B(n12108), .ZN(n9480) );
  AND2_X1 U14765 ( .A1(n10375), .A2(n10584), .ZN(n10589) );
  NAND2_X1 U14766 ( .A1(n10589), .A2(n10585), .ZN(n9442) );
  NOR2_X1 U14767 ( .A1(n10583), .A2(n10584), .ZN(n9440) );
  NAND2_X1 U14768 ( .A1(n10590), .A2(n9440), .ZN(n9441) );
  MUX2_X1 U14769 ( .A(n25021), .B(n9946), .S(n9945), .Z(n9448) );
  NOR2_X1 U14770 ( .A1(n9899), .A2(n9944), .ZN(n9446) );
  NOR2_X1 U14771 ( .A1(n9446), .A2(n9445), .ZN(n9447) );
  MUX2_X1 U14772 ( .A(n9908), .B(n24511), .S(n9904), .Z(n9453) );
  INV_X1 U14773 ( .A(n9905), .ZN(n9935) );
  NAND3_X1 U14774 ( .A1(n9449), .A2(n24511), .A3(n9908), .ZN(n9452) );
  INV_X1 U14775 ( .A(n9450), .ZN(n9938) );
  NAND3_X1 U14776 ( .A1(n9935), .A2(n9939), .A3(n9938), .ZN(n9451) );
  INV_X1 U14777 ( .A(n9454), .ZN(n9882) );
  INV_X1 U14778 ( .A(n25069), .ZN(n9455) );
  NAND3_X1 U14779 ( .A1(n9564), .A2(n9882), .A3(n9886), .ZN(n9457) );
  OAI21_X1 U14780 ( .B1(n9460), .B2(n9912), .A(n9458), .ZN(n9467) );
  AOI21_X1 U14781 ( .B1(n9465), .B2(n9464), .A(n9463), .ZN(n9466) );
  NOR2_X1 U14782 ( .A1(n3290), .A2(n9469), .ZN(n9470) );
  NAND3_X1 U14783 ( .A1(n24168), .A2(n24345), .A3(n10302), .ZN(n9479) );
  NAND2_X1 U14784 ( .A1(n9474), .A2(n239), .ZN(n9473) );
  NAND3_X1 U14785 ( .A1(n9558), .A2(n9560), .A3(n9860), .ZN(n9475) );
  XNOR2_X1 U14786 ( .A(n9480), .B(n11167), .ZN(n9573) );
  OAI21_X1 U14787 ( .B1(n25043), .B2(n9652), .A(n9723), .ZN(n9482) );
  NAND2_X1 U14788 ( .A1(n9482), .A2(n9725), .ZN(n9490) );
  NAND2_X1 U14789 ( .A1(n9724), .A2(n10008), .ZN(n9483) );
  NAND2_X1 U14790 ( .A1(n9483), .A2(n9652), .ZN(n9488) );
  NAND2_X1 U14791 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  OAI21_X1 U14792 ( .B1(n9731), .B2(n426), .A(n10019), .ZN(n9494) );
  NOR2_X1 U14794 ( .A1(n24505), .A2(n8571), .ZN(n9497) );
  OR3_X1 U14795 ( .A1(n9798), .A2(n9998), .A3(n8521), .ZN(n9499) );
  INV_X1 U14796 ( .A(n10775), .ZN(n9502) );
  NOR2_X1 U14797 ( .A1(n9797), .A2(n9671), .ZN(n9501) );
  NOR2_X1 U14798 ( .A1(n9775), .A2(n10104), .ZN(n9504) );
  AOI22_X1 U14799 ( .A1(n9504), .A2(n25393), .B1(n9775), .B2(n9503), .ZN(n9505) );
  OAI21_X1 U14800 ( .B1(n10080), .B2(n9786), .A(n10079), .ZN(n9506) );
  NAND3_X1 U14801 ( .A1(n4256), .A2(n9507), .A3(n10082), .ZN(n9508) );
  NAND2_X1 U14802 ( .A1(n10100), .A2(n10099), .ZN(n9514) );
  OAI21_X2 U14803 ( .B1(n9517), .B2(n9518), .A(n9516), .ZN(n11298) );
  INV_X1 U14804 ( .A(n10176), .ZN(n9831) );
  OAI211_X1 U14805 ( .C1(n10186), .C2(n10178), .A(n9831), .B(n10175), .ZN(
        n9519) );
  MUX2_X1 U14806 ( .A(n11301), .B(n11298), .S(n10762), .Z(n9536) );
  NAND2_X1 U14809 ( .A1(n9841), .A2(n25207), .ZN(n9521) );
  NAND2_X1 U14810 ( .A1(n9525), .A2(n9524), .ZN(n9528) );
  AOI21_X1 U14811 ( .B1(n9526), .B2(n9775), .A(n9773), .ZN(n9527) );
  NAND2_X1 U14812 ( .A1(n9532), .A2(n10113), .ZN(n9535) );
  NAND3_X1 U14813 ( .A1(n9533), .A2(n9805), .A3(n10116), .ZN(n9534) );
  XNOR2_X1 U14814 ( .A(n11396), .B(n9537), .ZN(n11420) );
  NAND2_X1 U14815 ( .A1(n4096), .A2(n24446), .ZN(n9538) );
  MUX2_X1 U14816 ( .A(n9539), .B(n9538), .S(n9866), .Z(n9540) );
  INV_X1 U14817 ( .A(n10028), .ZN(n9543) );
  NAND2_X1 U14818 ( .A1(n10031), .A2(n10026), .ZN(n9542) );
  AOI21_X1 U14819 ( .B1(n9543), .B2(n9542), .A(n10027), .ZN(n9546) );
  NAND2_X1 U14820 ( .A1(n9697), .A2(n9695), .ZN(n9643) );
  NAND3_X1 U14821 ( .A1(n9697), .A2(n9699), .A3(n10027), .ZN(n9544) );
  NAND2_X1 U14822 ( .A1(n9643), .A2(n9544), .ZN(n9545) );
  NAND3_X1 U14823 ( .A1(n1517), .A2(n307), .A3(n9692), .ZN(n9548) );
  OAI211_X2 U14824 ( .C1(n9549), .C2(n4993), .A(n9548), .B(n9547), .ZN(n10904)
         );
  NAND2_X1 U14825 ( .A1(n10445), .A2(n10904), .ZN(n9553) );
  NAND2_X1 U14826 ( .A1(n10044), .A2(n10045), .ZN(n9625) );
  OAI211_X1 U14827 ( .C1(n10046), .C2(n9681), .A(n9628), .B(n9627), .ZN(n9552)
         );
  NAND2_X1 U14828 ( .A1(n10048), .A2(n9681), .ZN(n9551) );
  NAND2_X1 U14829 ( .A1(n9558), .A2(n9560), .ZN(n9557) );
  NAND3_X1 U14830 ( .A1(n10445), .A2(n10907), .A3(n10904), .ZN(n9572) );
  NAND3_X1 U14831 ( .A1(n9882), .A2(n9886), .A3(n9567), .ZN(n9569) );
  OAI211_X1 U14832 ( .C1(n25069), .C2(n9567), .A(n9566), .B(n9565), .ZN(n9568)
         );
  NAND3_X1 U14833 ( .A1(n10902), .A2(n10747), .A3(n10901), .ZN(n9571) );
  INV_X1 U14834 ( .A(n12402), .ZN(n12067) );
  NOR2_X1 U14835 ( .A1(n10885), .A2(n10886), .ZN(n9574) );
  AOI22_X1 U14836 ( .A1(n10884), .A2(n9574), .B1(n10301), .B2(n10885), .ZN(
        n9575) );
  OAI22_X1 U14837 ( .A1(n10902), .A2(n10747), .B1(n4341), .B2(n10904), .ZN(
        n9579) );
  INV_X1 U14838 ( .A(n10901), .ZN(n9578) );
  NAND2_X1 U14839 ( .A1(n10444), .A2(n10905), .ZN(n9577) );
  XNOR2_X1 U14840 ( .A(n11845), .B(n12150), .ZN(n11087) );
  INV_X1 U14841 ( .A(n11087), .ZN(n9612) );
  INV_X1 U14843 ( .A(n10284), .ZN(n10286) );
  INV_X1 U14844 ( .A(n11385), .ZN(n9611) );
  INV_X1 U14845 ( .A(n10617), .ZN(n10610) );
  INV_X1 U14846 ( .A(n9832), .ZN(n10182) );
  OAI211_X1 U14847 ( .C1(n9832), .C2(n9831), .A(n9585), .B(n9584), .ZN(n9587)
         );
  NAND3_X1 U14848 ( .A1(n9832), .A2(n10177), .A3(n10175), .ZN(n9586) );
  INV_X1 U14849 ( .A(n10612), .ZN(n10341) );
  NAND2_X1 U14850 ( .A1(n9814), .A2(n10166), .ZN(n9590) );
  NAND2_X1 U14851 ( .A1(n10341), .A2(n10411), .ZN(n9610) );
  INV_X1 U14852 ( .A(n10161), .ZN(n9850) );
  INV_X1 U14853 ( .A(n10157), .ZN(n9851) );
  NAND3_X1 U14854 ( .A1(n3305), .A2(n10162), .A3(n9851), .ZN(n9594) );
  INV_X1 U14855 ( .A(n10486), .ZN(n10410) );
  NOR2_X1 U14856 ( .A1(n10129), .A2(n10128), .ZN(n9598) );
  NAND2_X1 U14857 ( .A1(n9595), .A2(n10127), .ZN(n9596) );
  NAND3_X1 U14858 ( .A1(n10410), .A2(n10614), .A3(n10341), .ZN(n9609) );
  OAI21_X1 U14859 ( .B1(n9927), .B2(n9934), .A(n9603), .ZN(n9602) );
  OAI21_X1 U14860 ( .B1(n9600), .B2(n9599), .A(n9926), .ZN(n9601) );
  NAND3_X1 U14861 ( .A1(n9928), .A2(n9604), .A3(n9603), .ZN(n9606) );
  NAND2_X1 U14862 ( .A1(n9927), .A2(n9925), .ZN(n9605) );
  XNOR2_X1 U14864 ( .A(n9611), .B(n12143), .ZN(n11446) );
  XNOR2_X1 U14865 ( .A(n11446), .B(n9612), .ZN(n9680) );
  AOI21_X1 U14866 ( .B1(n9757), .B2(n9752), .A(n9753), .ZN(n9618) );
  INV_X1 U14867 ( .A(n9613), .ZN(n9749) );
  NOR2_X1 U14868 ( .A1(n9754), .A2(n9749), .ZN(n9614) );
  OAI21_X1 U14869 ( .B1(n9615), .B2(n9614), .A(n9977), .ZN(n9616) );
  NOR2_X1 U14870 ( .A1(n9762), .A2(n9620), .ZN(n9619) );
  MUX2_X1 U14871 ( .A(n10068), .B(n9619), .S(n9231), .Z(n9623) );
  NAND2_X1 U14872 ( .A1(n1330), .A2(n9620), .ZN(n9621) );
  OAI21_X2 U14873 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n11338) );
  NAND2_X1 U14874 ( .A1(n10062), .A2(n9705), .ZN(n9624) );
  INV_X1 U14875 ( .A(n9625), .ZN(n9626) );
  OAI21_X1 U14877 ( .B1(n9628), .B2(n9627), .A(n10044), .ZN(n9629) );
  NAND2_X1 U14878 ( .A1(n9629), .A2(n9682), .ZN(n9631) );
  NAND3_X1 U14879 ( .A1(n10048), .A2(n9681), .A3(n10046), .ZN(n9630) );
  MUX2_X1 U14880 ( .A(n9635), .B(n9634), .S(n9633), .Z(n9638) );
  INV_X1 U14881 ( .A(n9714), .ZN(n9636) );
  AND2_X1 U14882 ( .A1(n9711), .A2(n10037), .ZN(n10043) );
  AOI22_X1 U14883 ( .A1(n9636), .A2(n9709), .B1(n9635), .B2(n10043), .ZN(n9637) );
  OAI21_X1 U14884 ( .B1(n9638), .B2(n9710), .A(n9637), .ZN(n10632) );
  INV_X1 U14885 ( .A(n9639), .ZN(n10034) );
  NAND2_X1 U14886 ( .A1(n10029), .A2(n10026), .ZN(n9640) );
  NAND3_X1 U14887 ( .A1(n9643), .A2(n10034), .A3(n9640), .ZN(n9642) );
  NAND3_X1 U14888 ( .A1(n9639), .A2(n24332), .A3(n10027), .ZN(n9641) );
  NAND2_X1 U14890 ( .A1(n10233), .A2(n10633), .ZN(n9644) );
  NAND2_X1 U14891 ( .A1(n25025), .A2(n11207), .ZN(n11340) );
  OAI21_X2 U14892 ( .B1(n9644), .B2(n9645), .A(n11340), .ZN(n12409) );
  NAND2_X1 U14893 ( .A1(n413), .A2(n10831), .ZN(n9649) );
  AND2_X1 U14894 ( .A1(n10515), .A2(n9646), .ZN(n9648) );
  XNOR2_X1 U14895 ( .A(n24980), .B(n12409), .ZN(n9678) );
  NOR2_X1 U14896 ( .A1(n10019), .A2(n8839), .ZN(n9650) );
  NOR2_X1 U14897 ( .A1(n9721), .A2(n10005), .ZN(n9651) );
  NAND2_X1 U14898 ( .A1(n9996), .A2(n9991), .ZN(n9660) );
  NOR2_X1 U14900 ( .A1(n9746), .A2(n9990), .ZN(n9661) );
  NAND3_X1 U14902 ( .A1(n9980), .A2(n9737), .A3(n9664), .ZN(n9665) );
  NAND2_X1 U14903 ( .A1(n9737), .A2(n9981), .ZN(n9666) );
  AOI21_X1 U14904 ( .B1(n9980), .B2(n9666), .A(n9740), .ZN(n9667) );
  NOR2_X1 U14905 ( .A1(n25453), .A2(n9671), .ZN(n9672) );
  NAND2_X1 U14906 ( .A1(n9672), .A2(n9796), .ZN(n9673) );
  NOR2_X1 U14907 ( .A1(n9798), .A2(n8521), .ZN(n9795) );
  OAI211_X1 U14908 ( .C1(n9781), .C2(n10093), .A(n9295), .B(n1348), .ZN(n9675)
         );
  NOR2_X1 U14909 ( .A1(n11201), .A2(n11196), .ZN(n10788) );
  XNOR2_X1 U14910 ( .A(n12102), .B(n859), .ZN(n9677) );
  XNOR2_X1 U14911 ( .A(n9678), .B(n9677), .ZN(n9679) );
  AOI21_X1 U14912 ( .B1(n12648), .B2(n12871), .A(n13094), .ZN(n10201) );
  OAI21_X1 U14913 ( .B1(n9682), .B2(n10045), .A(n9681), .ZN(n9687) );
  NAND2_X1 U14914 ( .A1(n9684), .A2(n10048), .ZN(n9685) );
  MUX2_X1 U14915 ( .A(n9689), .B(n9688), .S(n4096), .Z(n9690) );
  NOR2_X1 U14916 ( .A1(n10026), .A2(n24332), .ZN(n9698) );
  NOR2_X1 U14917 ( .A1(n9639), .A2(n9699), .ZN(n9700) );
  NAND2_X1 U14918 ( .A1(n10061), .A2(n9705), .ZN(n9706) );
  NAND2_X1 U14919 ( .A1(n9708), .A2(n9707), .ZN(n11143) );
  NAND2_X1 U14920 ( .A1(n10304), .A2(n11151), .ZN(n9719) );
  OR2_X1 U14922 ( .A1(n9712), .A2(n9713), .ZN(n9717) );
  INV_X1 U14923 ( .A(n10039), .ZN(n9716) );
  NAND2_X1 U14924 ( .A1(n9714), .A2(n9713), .ZN(n9715) );
  OR2_X1 U14925 ( .A1(n9718), .A2(n9433), .ZN(n11146) );
  MUX2_X1 U14926 ( .A(n9723), .B(n9722), .S(n9299), .Z(n9728) );
  NOR2_X1 U14927 ( .A1(n9724), .A2(n10008), .ZN(n9726) );
  NAND2_X1 U14929 ( .A1(n9730), .A2(n9729), .ZN(n10016) );
  INV_X1 U14930 ( .A(n10016), .ZN(n9735) );
  NAND2_X1 U14931 ( .A1(n9731), .A2(n426), .ZN(n9734) );
  OAI21_X1 U14932 ( .B1(n9735), .B2(n9734), .A(n9733), .ZN(n11159) );
  NAND3_X1 U14933 ( .A1(n9740), .A2(n9737), .A3(n9985), .ZN(n9738) );
  AND2_X1 U14934 ( .A1(n9739), .A2(n9738), .ZN(n9744) );
  NAND2_X1 U14935 ( .A1(n9982), .A2(n9981), .ZN(n9741) );
  MUX2_X1 U14936 ( .A(n9742), .B(n9741), .S(n9740), .Z(n9743) );
  NAND2_X2 U14937 ( .A1(n9743), .A2(n9744), .ZN(n11157) );
  MUX2_X1 U14938 ( .A(n1358), .B(n4737), .S(n11157), .Z(n9768) );
  NAND2_X1 U14940 ( .A1(n9751), .A2(n9750), .ZN(n9756) );
  AND3_X1 U14941 ( .A1(n9753), .A2(n9754), .A3(n9752), .ZN(n9755) );
  AOI21_X1 U14942 ( .B1(n9756), .B2(n9973), .A(n9755), .ZN(n10675) );
  NAND2_X1 U14943 ( .A1(n9758), .A2(n9757), .ZN(n10673) );
  NAND2_X1 U14944 ( .A1(n10985), .A2(n11160), .ZN(n9759) );
  OAI21_X1 U14945 ( .B1(n11160), .B2(n11157), .A(n9759), .ZN(n9767) );
  NOR2_X1 U14946 ( .A1(n10075), .A2(n9231), .ZN(n9761) );
  NAND3_X1 U14947 ( .A1(n9764), .A2(n9763), .A3(n9762), .ZN(n9765) );
  XNOR2_X1 U14948 ( .A(n12002), .B(n11967), .ZN(n11642) );
  INV_X1 U14949 ( .A(n11642), .ZN(n11725) );
  OAI21_X1 U14950 ( .B1(n10681), .B2(n24622), .A(n11003), .ZN(n9771) );
  MUX2_X2 U14951 ( .A(n9771), .B(n9770), .S(n10685), .Z(n11289) );
  MUX2_X1 U14952 ( .A(n10108), .B(n9774), .S(n9772), .Z(n9776) );
  NAND2_X1 U14953 ( .A1(n9774), .A2(n9773), .ZN(n10110) );
  NAND2_X1 U14954 ( .A1(n9775), .A2(n10104), .ZN(n10107) );
  NAND2_X1 U14955 ( .A1(n1348), .A2(n10089), .ZN(n9778) );
  NAND2_X1 U14956 ( .A1(n8571), .A2(n9295), .ZN(n9777) );
  NAND3_X1 U14957 ( .A1(n10090), .A2(n9778), .A3(n9777), .ZN(n9785) );
  NAND3_X1 U14958 ( .A1(n9782), .A2(n24505), .A3(n9780), .ZN(n9783) );
  NOR2_X1 U14959 ( .A1(n11054), .A2(n11009), .ZN(n9803) );
  NOR2_X1 U14960 ( .A1(n10094), .A2(n10099), .ZN(n9790) );
  INV_X1 U14961 ( .A(n10094), .ZN(n9791) );
  NAND2_X1 U14962 ( .A1(n9791), .A2(n10098), .ZN(n9792) );
  OAI22_X1 U14963 ( .A1(n9838), .A2(n10095), .B1(n9792), .B2(n9837), .ZN(n9793) );
  NOR3_X1 U14964 ( .A1(n9811), .A2(n11052), .A3(n9810), .ZN(n9802) );
  NOR2_X1 U14965 ( .A1(n9997), .A2(n9998), .ZN(n9799) );
  OAI21_X1 U14966 ( .B1(n9799), .B2(n9999), .A(n9798), .ZN(n9800) );
  INV_X1 U14967 ( .A(n11440), .ZN(n9812) );
  XNOR2_X1 U14968 ( .A(n11289), .B(n9812), .ZN(n9813) );
  XNOR2_X1 U14969 ( .A(n11725), .B(n9813), .ZN(n9971) );
  INV_X1 U14970 ( .A(n9820), .ZN(n9821) );
  NAND2_X1 U14971 ( .A1(n25463), .A2(n9821), .ZN(n9824) );
  NAND3_X1 U14972 ( .A1(n10136), .A2(n9820), .A3(n25463), .ZN(n9823) );
  OAI211_X1 U14974 ( .C1(n10138), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9826)
         );
  INV_X1 U14975 ( .A(n9827), .ZN(n9828) );
  NAND2_X1 U14976 ( .A1(n9828), .A2(n10176), .ZN(n9835) );
  OAI211_X1 U14977 ( .C1(n9831), .C2(n10175), .A(n9830), .B(n9829), .ZN(n9834)
         );
  NAND3_X1 U14978 ( .A1(n10186), .A2(n9832), .A3(n10178), .ZN(n9833) );
  INV_X1 U14979 ( .A(n10703), .ZN(n10699) );
  OAI21_X1 U14980 ( .B1(n25206), .B2(n25486), .A(n9841), .ZN(n9848) );
  NAND2_X1 U14981 ( .A1(n9844), .A2(n10148), .ZN(n9847) );
  NAND3_X1 U14982 ( .A1(n1210), .A2(n24085), .A3(n9845), .ZN(n9846) );
  OAI211_X1 U14983 ( .C1(n9851), .C2(n10162), .A(n9850), .B(n9849), .ZN(n9852)
         );
  OAI21_X1 U14984 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n10953) );
  INV_X1 U14985 ( .A(n11637), .ZN(n9855) );
  XNOR2_X1 U14986 ( .A(n9855), .B(n2761), .ZN(n9969) );
  MUX2_X1 U14987 ( .A(n239), .B(n9860), .S(n9856), .Z(n9865) );
  NAND2_X1 U14988 ( .A1(n9857), .A2(n9864), .ZN(n9862) );
  MUX2_X1 U14989 ( .A(n9862), .B(n9861), .S(n9860), .Z(n9863) );
  INV_X1 U14991 ( .A(n10971), .ZN(n9871) );
  INV_X1 U14992 ( .A(n9867), .ZN(n9868) );
  NAND2_X1 U14993 ( .A1(n9871), .A2(n10970), .ZN(n10608) );
  NAND3_X1 U14994 ( .A1(n9875), .A2(n24549), .A3(n9027), .ZN(n9878) );
  INV_X1 U14995 ( .A(n9876), .ZN(n9877) );
  NAND2_X1 U14996 ( .A1(n25497), .A2(n10968), .ZN(n9881) );
  NAND2_X1 U14997 ( .A1(n10608), .A2(n9881), .ZN(n9911) );
  NAND2_X1 U14998 ( .A1(n8157), .A2(n9886), .ZN(n9888) );
  NAND2_X1 U14999 ( .A1(n9891), .A2(n9890), .ZN(n9892) );
  INV_X1 U15000 ( .A(n9892), .ZN(n10967) );
  NAND2_X1 U15001 ( .A1(n227), .A2(n9943), .ZN(n9894) );
  NAND2_X1 U15002 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  NAND3_X1 U15003 ( .A1(n9899), .A2(n24054), .A3(n9897), .ZN(n9901) );
  NAND3_X1 U15004 ( .A1(n9942), .A2(n9946), .A3(n24083), .ZN(n9900) );
  NOR2_X1 U15005 ( .A1(n10818), .A2(n9903), .ZN(n9910) );
  OAI21_X1 U15006 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(n9909) );
  INV_X1 U15007 ( .A(n9912), .ZN(n9917) );
  INV_X1 U15008 ( .A(n9913), .ZN(n9915) );
  AOI22_X1 U15009 ( .A1(n9917), .A2(n9916), .B1(n9915), .B2(n9914), .ZN(n9924)
         );
  NAND2_X1 U15010 ( .A1(n24844), .A2(n9918), .ZN(n9922) );
  INV_X1 U15012 ( .A(n9929), .ZN(n9933) );
  INV_X1 U15013 ( .A(n9930), .ZN(n9932) );
  OAI21_X1 U15015 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(n9940) );
  NAND2_X1 U15016 ( .A1(n10804), .A2(n411), .ZN(n9968) );
  NAND3_X1 U15017 ( .A1(n10798), .A2(n10799), .A3(n10648), .ZN(n9967) );
  MUX2_X1 U15018 ( .A(n9953), .B(n9948), .S(n9947), .Z(n9960) );
  NAND2_X1 U15019 ( .A1(n9950), .A2(n9949), .ZN(n9956) );
  OAI21_X1 U15020 ( .B1(n9956), .B2(n9955), .A(n9954), .ZN(n9957) );
  INV_X1 U15021 ( .A(n9957), .ZN(n9958) );
  OAI21_X1 U15022 ( .B1(n9960), .B2(n9959), .A(n9958), .ZN(n10426) );
  INV_X1 U15023 ( .A(n10426), .ZN(n10649) );
  NOR2_X1 U15024 ( .A1(n10649), .A2(n10648), .ZN(n10803) );
  INV_X1 U15025 ( .A(n10651), .ZN(n10801) );
  INV_X1 U15026 ( .A(n10245), .ZN(n10244) );
  XNOR2_X1 U15027 ( .A(n11194), .B(n9969), .ZN(n9970) );
  OAI21_X1 U15028 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(n9976) );
  NAND2_X1 U15029 ( .A1(n9978), .A2(n9981), .ZN(n9979) );
  MUX2_X1 U15031 ( .A(n9991), .B(n9990), .S(n9989), .Z(n9994) );
  INV_X1 U15032 ( .A(n11045), .ZN(n10642) );
  AOI21_X1 U15033 ( .B1(n2680), .B2(n11046), .A(n10642), .ZN(n10014) );
  NAND2_X1 U15034 ( .A1(n10006), .A2(n10005), .ZN(n10011) );
  NOR2_X1 U15035 ( .A1(n25043), .A2(n9301), .ZN(n10010) );
  NAND2_X1 U15036 ( .A1(n9299), .A2(n10008), .ZN(n10009) );
  AOI22_X1 U15037 ( .A1(n10012), .A2(n10011), .B1(n10010), .B2(n10009), .ZN(
        n11051) );
  MUX2_X1 U15038 ( .A(n10020), .B(n10019), .S(n10018), .Z(n10021) );
  NOR2_X1 U15039 ( .A1(n10021), .A2(n8839), .ZN(n10022) );
  NAND2_X1 U15040 ( .A1(n11044), .A2(n10416), .ZN(n11050) );
  NAND2_X1 U15041 ( .A1(n10801), .A2(n10648), .ZN(n10025) );
  OAI21_X1 U15042 ( .B1(n10426), .B2(n10245), .A(n10799), .ZN(n10023) );
  NOR2_X1 U15043 ( .A1(n10023), .A2(n411), .ZN(n10024) );
  AOI21_X2 U15044 ( .B1(n10427), .B2(n10025), .A(n10024), .ZN(n11542) );
  XNOR2_X1 U15045 ( .A(n11542), .B(n12082), .ZN(n10124) );
  MUX2_X1 U15046 ( .A(n10031), .B(n24332), .S(n10026), .Z(n10035) );
  NAND2_X1 U15047 ( .A1(n10028), .A2(n10027), .ZN(n10033) );
  NAND3_X1 U15048 ( .A1(n10031), .A2(n24332), .A3(n10029), .ZN(n10032) );
  OAI211_X2 U15049 ( .C1(n10035), .C2(n10034), .A(n10033), .B(n10032), .ZN(
        n11064) );
  NAND2_X1 U15050 ( .A1(n9433), .A2(n9709), .ZN(n10042) );
  NAND2_X1 U15051 ( .A1(n10038), .A2(n10037), .ZN(n10040) );
  NAND2_X1 U15052 ( .A1(n10040), .A2(n10039), .ZN(n10041) );
  NOR2_X1 U15053 ( .A1(n11064), .A2(n11069), .ZN(n10665) );
  MUX2_X1 U15054 ( .A(n10045), .B(n260), .S(n10044), .Z(n10049) );
  OAI21_X1 U15055 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(n10056) );
  MUX2_X1 U15056 ( .A(n10064), .B(n10063), .S(n9127), .Z(n10066) );
  OAI22_X1 U15057 ( .A1(n1330), .A2(n10070), .B1(n25457), .B2(n9231), .ZN(
        n10073) );
  NAND2_X1 U15058 ( .A1(n10073), .A2(n10072), .ZN(n10074) );
  INV_X1 U15060 ( .A(n11062), .ZN(n11071) );
  NOR2_X1 U15061 ( .A1(n11070), .A2(n11071), .ZN(n10078) );
  INV_X1 U15062 ( .A(n10665), .ZN(n10077) );
  NAND2_X1 U15063 ( .A1(n10080), .A2(n10079), .ZN(n10081) );
  NAND2_X1 U15064 ( .A1(n10087), .A2(n10081), .ZN(n10085) );
  NAND2_X1 U15065 ( .A1(n10082), .A2(n10088), .ZN(n10084) );
  MUX2_X1 U15066 ( .A(n10085), .B(n10084), .S(n24575), .Z(n10086) );
  NAND2_X1 U15067 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  NAND3_X1 U15068 ( .A1(n10100), .A2(n10094), .A3(n10099), .ZN(n10096) );
  OAI21_X1 U15069 ( .B1(n421), .B2(n10097), .A(n10096), .ZN(n10103) );
  NOR2_X1 U15072 ( .A1(n10110), .A2(n10109), .ZN(n10111) );
  OAI22_X1 U15073 ( .A1(n10114), .A2(n1406), .B1(n10113), .B2(n10112), .ZN(
        n10119) );
  NAND3_X1 U15074 ( .A1(n10117), .A2(n10116), .A3(n10115), .ZN(n10118) );
  XNOR2_X1 U15075 ( .A(n12053), .B(n11424), .ZN(n11391) );
  XNOR2_X1 U15076 ( .A(n11391), .B(n10124), .ZN(n10198) );
  NAND2_X1 U15077 ( .A1(n10127), .A2(n10126), .ZN(n10133) );
  NAND2_X1 U15078 ( .A1(n10129), .A2(n10128), .ZN(n10130) );
  INV_X1 U15080 ( .A(n10559), .ZN(n10659) );
  NOR2_X1 U15082 ( .A1(n9398), .A2(n24026), .ZN(n10139) );
  OAI21_X1 U15083 ( .B1(n10139), .B2(n10138), .A(n25463), .ZN(n10144) );
  NAND2_X1 U15084 ( .A1(n10659), .A2(n10654), .ZN(n10314) );
  NOR2_X1 U15085 ( .A1(n25206), .A2(n10148), .ZN(n10152) );
  NOR2_X1 U15086 ( .A1(n10149), .A2(n10148), .ZN(n10151) );
  NOR2_X1 U15087 ( .A1(n10158), .A2(n10157), .ZN(n10160) );
  OAI22_X1 U15088 ( .A1(n3305), .A2(n10162), .B1(n10161), .B2(n9349), .ZN(
        n10164) );
  OAI21_X1 U15089 ( .B1(n10165), .B2(n25250), .A(n10657), .ZN(n10189) );
  NOR2_X1 U15090 ( .A1(n10170), .A2(n10169), .ZN(n10171) );
  NOR2_X1 U15091 ( .A1(n10172), .A2(n1577), .ZN(n10173) );
  NAND3_X1 U15092 ( .A1(n10176), .A2(n10178), .A3(n10175), .ZN(n10184) );
  INV_X1 U15093 ( .A(n10177), .ZN(n10179) );
  NOR2_X1 U15094 ( .A1(n10654), .A2(n10660), .ZN(n10187) );
  OAI21_X1 U15095 ( .B1(n10661), .B2(n25250), .A(n10187), .ZN(n10188) );
  NAND2_X1 U15096 ( .A1(n10189), .A2(n10188), .ZN(n11660) );
  INV_X1 U15097 ( .A(n25229), .ZN(n10854) );
  INV_X1 U15099 ( .A(n10737), .ZN(n10465) );
  OAI211_X1 U15100 ( .C1(n10831), .C2(n10277), .A(n10830), .B(n10518), .ZN(
        n10194) );
  XNOR2_X1 U15101 ( .A(n12255), .B(n22702), .ZN(n10195) );
  XNOR2_X1 U15102 ( .A(n10196), .B(n10195), .ZN(n10197) );
  INV_X1 U15103 ( .A(n14158), .ZN(n10396) );
  NOR2_X1 U15104 ( .A1(n10756), .A2(n10757), .ZN(n10203) );
  NOR2_X1 U15105 ( .A1(n11298), .A2(n11301), .ZN(n10205) );
  NAND2_X1 U15106 ( .A1(n10895), .A2(n10205), .ZN(n10207) );
  NAND3_X1 U15107 ( .A1(n11091), .A2(n11301), .A3(n10762), .ZN(n10206) );
  XNOR2_X1 U15108 ( .A(n12314), .B(n11263), .ZN(n11829) );
  INV_X1 U15109 ( .A(n10208), .ZN(n10211) );
  INV_X1 U15110 ( .A(n10209), .ZN(n10210) );
  NAND3_X1 U15111 ( .A1(n10211), .A2(n10538), .A3(n10210), .ZN(n10212) );
  NAND2_X1 U15112 ( .A1(n10585), .A2(n10371), .ZN(n10317) );
  INV_X1 U15113 ( .A(n10584), .ZN(n10582) );
  AND2_X1 U15114 ( .A1(n10587), .A2(n25507), .ZN(n10215) );
  OAI21_X1 U15115 ( .B1(n10590), .B2(n10584), .A(n10215), .ZN(n10216) );
  NAND2_X1 U15116 ( .A1(n10217), .A2(n10216), .ZN(n11747) );
  XNOR2_X1 U15117 ( .A(n12218), .B(n11747), .ZN(n11481) );
  XNOR2_X1 U15118 ( .A(n11829), .B(n11481), .ZN(n10226) );
  INV_X1 U15119 ( .A(n10891), .ZN(n11081) );
  NAND2_X1 U15120 ( .A1(n10767), .A2(n412), .ZN(n10766) );
  XNOR2_X1 U15122 ( .A(n11616), .B(n12313), .ZN(n10224) );
  INV_X1 U15123 ( .A(n10904), .ZN(n10899) );
  XNOR2_X1 U15124 ( .A(n12159), .B(n2228), .ZN(n10223) );
  XNOR2_X1 U15125 ( .A(n10224), .B(n10223), .ZN(n10225) );
  XNOR2_X1 U15126 ( .A(n10226), .B(n10225), .ZN(n12724) );
  INV_X1 U15127 ( .A(n12724), .ZN(n13176) );
  NAND2_X1 U15129 ( .A1(n44), .A2(n11199), .ZN(n10228) );
  NAND2_X1 U15130 ( .A1(n11201), .A2(n11196), .ZN(n10227) );
  INV_X1 U15132 ( .A(n10789), .ZN(n11195) );
  OAI211_X1 U15133 ( .C1(n10793), .C2(n11195), .A(n10477), .B(n10229), .ZN(
        n10230) );
  AND2_X1 U15134 ( .A1(n10632), .A2(n11338), .ZN(n10232) );
  INV_X1 U15135 ( .A(n10411), .ZN(n10489) );
  AOI22_X1 U15136 ( .A1(n10617), .A2(n10616), .B1(n10489), .B2(n10614), .ZN(
        n10237) );
  NOR2_X1 U15137 ( .A1(n10614), .A2(n10486), .ZN(n10234) );
  NAND2_X1 U15138 ( .A1(n10610), .A2(n10234), .ZN(n10236) );
  NOR3_X1 U15139 ( .A1(n10486), .A2(n10411), .A3(n10613), .ZN(n10235) );
  NAND3_X1 U15140 ( .A1(n233), .A2(n11212), .A3(n11216), .ZN(n10238) );
  XNOR2_X1 U15141 ( .A(n10239), .B(n12046), .ZN(n10270) );
  INV_X1 U15142 ( .A(n10968), .ZN(n10607) );
  OAI21_X1 U15143 ( .B1(n10497), .B2(n10607), .A(n10606), .ZN(n10240) );
  NOR2_X1 U15144 ( .A1(n25497), .A2(n10968), .ZN(n10496) );
  NOR2_X1 U15145 ( .A1(n10606), .A2(n10969), .ZN(n10242) );
  NOR2_X1 U15146 ( .A1(n25497), .A2(n10970), .ZN(n10241) );
  NAND3_X1 U15147 ( .A1(n10805), .A2(n10799), .A3(n10244), .ZN(n10247) );
  NAND4_X2 U15148 ( .A1(n10246), .A2(n10248), .A3(n10249), .A4(n10247), .ZN(
        n12201) );
  XNOR2_X1 U15149 ( .A(n12122), .B(n12201), .ZN(n12242) );
  INV_X1 U15150 ( .A(n10256), .ZN(n10258) );
  AND2_X1 U15151 ( .A1(n10257), .A2(n10258), .ZN(n10260) );
  NAND4_X1 U15152 ( .A1(n10261), .A2(n10480), .A3(n10260), .A4(n10259), .ZN(
        n10265) );
  INV_X1 U15153 ( .A(n10262), .ZN(n10263) );
  NAND2_X1 U15154 ( .A1(n10263), .A2(n11190), .ZN(n10264) );
  XNOR2_X1 U15156 ( .A(n12383), .B(n3125), .ZN(n10268) );
  XNOR2_X1 U15157 ( .A(n12242), .B(n10268), .ZN(n10269) );
  INV_X1 U15158 ( .A(n12459), .ZN(n13177) );
  NAND2_X1 U15159 ( .A1(n11189), .A2(n11190), .ZN(n11371) );
  NOR2_X1 U15160 ( .A1(n11190), .A2(n10728), .ZN(n11185) );
  NAND2_X1 U15161 ( .A1(n11371), .A2(n11370), .ZN(n11809) );
  MUX2_X1 U15163 ( .A(n10464), .B(n10272), .S(n11123), .Z(n10274) );
  INV_X1 U15164 ( .A(n11123), .ZN(n10720) );
  AND2_X1 U15165 ( .A1(n10850), .A2(n2244), .ZN(n10851) );
  AOI22_X1 U15166 ( .A1(n10851), .A2(n11124), .B1(n10722), .B2(n10848), .ZN(
        n10273) );
  XNOR2_X1 U15167 ( .A(n11809), .B(n11492), .ZN(n12303) );
  NAND2_X1 U15168 ( .A1(n10829), .A2(n10277), .ZN(n10514) );
  NOR2_X1 U15169 ( .A1(n9279), .A2(n10514), .ZN(n10278) );
  NOR2_X2 U15170 ( .A1(n10279), .A2(n10278), .ZN(n12184) );
  OAI21_X1 U15171 ( .B1(n10860), .B2(n10861), .A(n10854), .ZN(n10281) );
  XNOR2_X1 U15172 ( .A(n12184), .B(n12128), .ZN(n12269) );
  MUX2_X1 U15174 ( .A(n10284), .B(n24574), .S(n11117), .Z(n10289) );
  INV_X1 U15175 ( .A(n10285), .ZN(n10287) );
  NAND2_X1 U15176 ( .A1(n10287), .A2(n10727), .ZN(n10288) );
  INV_X1 U15177 ( .A(n10451), .ZN(n10752) );
  XNOR2_X1 U15178 ( .A(n11966), .B(n12186), .ZN(n10298) );
  NAND2_X1 U15179 ( .A1(n10713), .A2(n11128), .ZN(n10296) );
  AND2_X1 U15180 ( .A1(n11128), .A2(n11130), .ZN(n10712) );
  INV_X1 U15181 ( .A(n10712), .ZN(n10292) );
  XNOR2_X1 U15183 ( .A(n11698), .B(n20825), .ZN(n10297) );
  XNOR2_X1 U15184 ( .A(n10298), .B(n10297), .ZN(n10299) );
  AOI21_X1 U15185 ( .B1(n10541), .B2(n10885), .A(n10887), .ZN(n10303) );
  INV_X1 U15186 ( .A(n10304), .ZN(n10305) );
  NAND3_X1 U15187 ( .A1(n714), .A2(n11143), .A3(n1357), .ZN(n10307) );
  XNOR2_X1 U15188 ( .A(n11310), .B(n11776), .ZN(n11536) );
  INV_X1 U15189 ( .A(n11157), .ZN(n10676) );
  OAI21_X1 U15190 ( .B1(n10676), .B2(n4737), .A(n11158), .ZN(n10309) );
  XNOR2_X1 U15191 ( .A(n11607), .B(n21204), .ZN(n10310) );
  NAND2_X1 U15192 ( .A1(n10548), .A2(n2754), .ZN(n10311) );
  OAI211_X1 U15193 ( .C1(n10548), .C2(n10950), .A(n10312), .B(n10311), .ZN(
        n12297) );
  NAND2_X1 U15194 ( .A1(n11170), .A2(n11168), .ZN(n10940) );
  OAI21_X1 U15196 ( .B1(n10587), .B2(n25507), .A(n10585), .ZN(n10318) );
  XNOR2_X1 U15197 ( .A(n12248), .B(n25371), .ZN(n11489) );
  XNOR2_X1 U15198 ( .A(n11489), .B(n12028), .ZN(n10320) );
  NOR2_X1 U15199 ( .A1(n10360), .A2(n12724), .ZN(n10361) );
  INV_X1 U15200 ( .A(n11005), .ZN(n10365) );
  MUX2_X1 U15201 ( .A(n5746), .B(n10321), .S(n10685), .Z(n10324) );
  NAND2_X1 U15202 ( .A1(n10684), .A2(n24622), .ZN(n10322) );
  AOI21_X1 U15203 ( .B1(n11003), .B2(n10322), .A(n10369), .ZN(n10323) );
  INV_X1 U15205 ( .A(n10924), .ZN(n10989) );
  NAND3_X1 U15207 ( .A1(n24118), .A2(n10405), .A3(n10990), .ZN(n10325) );
  NAND2_X1 U15208 ( .A1(n10924), .A2(n10993), .ZN(n10407) );
  OAI21_X1 U15209 ( .B1(n10407), .B2(n24118), .A(n10328), .ZN(n10329) );
  XNOR2_X1 U15210 ( .A(n12109), .B(n12189), .ZN(n12274) );
  AOI21_X1 U15211 ( .B1(n11052), .B2(n11057), .A(n11054), .ZN(n11500) );
  NAND2_X1 U15212 ( .A1(n11500), .A2(n11059), .ZN(n10335) );
  NAND2_X1 U15213 ( .A1(n11500), .A2(n11052), .ZN(n10334) );
  INV_X1 U15214 ( .A(n11052), .ZN(n10694) );
  OR2_X1 U15216 ( .A1(n11059), .A2(n10331), .ZN(n10333) );
  NOR2_X1 U15217 ( .A1(n11499), .A2(n11009), .ZN(n10332) );
  NAND2_X1 U15218 ( .A1(n11054), .A2(n10332), .ZN(n11501) );
  NAND4_X1 U15219 ( .A1(n10335), .A2(n10334), .A3(n10333), .A4(n11501), .ZN(
        n11274) );
  OAI22_X1 U15220 ( .A1(n10337), .A2(n10398), .B1(n10658), .B2(n10559), .ZN(
        n10340) );
  OR2_X1 U15221 ( .A1(n10559), .A2(n10660), .ZN(n10400) );
  INV_X1 U15222 ( .A(n10654), .ZN(n10557) );
  NAND2_X1 U15223 ( .A1(n10559), .A2(n10557), .ZN(n10338) );
  AOI21_X1 U15224 ( .B1(n10400), .B2(n10338), .A(n10558), .ZN(n10339) );
  XNOR2_X1 U15226 ( .A(n11622), .B(n11274), .ZN(n12063) );
  XNOR2_X1 U15227 ( .A(n12274), .B(n12063), .ZN(n10359) );
  AND2_X1 U15228 ( .A1(n10486), .A2(n10613), .ZN(n10342) );
  NOR2_X1 U15229 ( .A1(n10488), .A2(n10613), .ZN(n10343) );
  NOR3_X1 U15230 ( .A1(n10343), .A2(n10342), .A3(n10610), .ZN(n10344) );
  MUX2_X1 U15231 ( .A(n11068), .B(n11062), .S(n11064), .Z(n10346) );
  NAND2_X1 U15232 ( .A1(n10346), .A2(n25203), .ZN(n10350) );
  NAND3_X1 U15233 ( .A1(n11070), .A2(n11071), .A3(n11067), .ZN(n10349) );
  INV_X1 U15234 ( .A(n25203), .ZN(n10662) );
  AND3_X2 U15235 ( .A1(n10350), .A2(n10349), .A3(n10348), .ZN(n12333) );
  XNOR2_X1 U15236 ( .A(n11951), .B(n12333), .ZN(n10357) );
  NOR2_X1 U15237 ( .A1(n11045), .A2(n2680), .ZN(n10352) );
  NOR2_X1 U15238 ( .A1(n10642), .A2(n11044), .ZN(n10351) );
  OAI21_X1 U15239 ( .B1(n10352), .B2(n10351), .A(n11012), .ZN(n10355) );
  NAND3_X1 U15240 ( .A1(n11044), .A2(n2680), .A3(n10641), .ZN(n10354) );
  NAND3_X1 U15241 ( .A1(n10355), .A2(n10354), .A3(n10353), .ZN(n11686) );
  XNOR2_X1 U15242 ( .A(n11686), .B(n1863), .ZN(n10356) );
  XNOR2_X1 U15243 ( .A(n10357), .B(n10356), .ZN(n10358) );
  XNOR2_X1 U15244 ( .A(n10359), .B(n10358), .ZN(n12725) );
  INV_X1 U15245 ( .A(n12460), .ZN(n12651) );
  OAI22_X1 U15246 ( .A1(n10362), .A2(n10361), .B1(n12651), .B2(n12506), .ZN(
        n10395) );
  NAND3_X1 U15247 ( .A1(n10365), .A2(n10681), .A3(n11004), .ZN(n10366) );
  XNOR2_X1 U15249 ( .A(n11960), .B(n4233), .ZN(n10378) );
  INV_X1 U15250 ( .A(n10370), .ZN(n10374) );
  AND2_X1 U15251 ( .A1(n10587), .A2(n10371), .ZN(n10373) );
  OAI21_X1 U15252 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(n10377) );
  AOI22_X1 U15253 ( .A1(n10589), .A2(n10590), .B1(n10375), .B2(n10585), .ZN(
        n10376) );
  XNOR2_X1 U15254 ( .A(n10378), .B(n12324), .ZN(n10381) );
  INV_X1 U15255 ( .A(n10942), .ZN(n10574) );
  OAI21_X1 U15256 ( .B1(n10406), .B2(n10990), .A(n10927), .ZN(n10380) );
  XNOR2_X1 U15257 ( .A(n12151), .B(n12207), .ZN(n12288) );
  XNOR2_X1 U15258 ( .A(n12288), .B(n10381), .ZN(n10392) );
  NAND3_X1 U15259 ( .A1(n11175), .A2(n11171), .A3(n24957), .ZN(n10383) );
  AOI21_X1 U15260 ( .B1(n11529), .B2(n11520), .A(n10922), .ZN(n10386) );
  OAI21_X1 U15261 ( .B1(n10384), .B2(n11525), .A(n11522), .ZN(n10385) );
  OAI22_X1 U15262 ( .A1(n10386), .A2(n10385), .B1(n11520), .B2(n11525), .ZN(
        n10387) );
  XNOR2_X1 U15263 ( .A(n11959), .B(n10387), .ZN(n10391) );
  NOR2_X1 U15264 ( .A1(n10935), .A2(n10931), .ZN(n10389) );
  NOR2_X1 U15265 ( .A1(n10931), .A2(n10505), .ZN(n10388) );
  AOI22_X1 U15266 ( .A1(n10936), .A2(n10389), .B1(n10388), .B2(n24470), .ZN(
        n10390) );
  INV_X1 U15267 ( .A(n10594), .ZN(n10595) );
  XNOR2_X1 U15268 ( .A(n10391), .B(n12213), .ZN(n11284) );
  OAI21_X1 U15270 ( .B1(n10398), .B2(n10558), .A(n10397), .ZN(n10402) );
  NAND2_X1 U15271 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  MUX2_X1 U15272 ( .A(n11067), .B(n11064), .S(n11070), .Z(n10404) );
  MUX2_X1 U15273 ( .A(n25203), .B(n11069), .S(n11064), .Z(n10403) );
  MUX2_X1 U15274 ( .A(n10404), .B(n10403), .S(n11062), .Z(n12130) );
  MUX2_X1 U15275 ( .A(n10994), .B(n10406), .S(n10405), .Z(n10409) );
  OAI21_X1 U15276 ( .B1(n10993), .B2(n10409), .A(n10408), .ZN(n12351) );
  XNOR2_X1 U15277 ( .A(n12130), .B(n12351), .ZN(n12005) );
  NAND2_X1 U15278 ( .A1(n10410), .A2(n10489), .ZN(n10414) );
  NOR2_X1 U15279 ( .A1(n10411), .A2(n10612), .ZN(n10487) );
  NAND2_X1 U15280 ( .A1(n10617), .A2(n10487), .ZN(n10413) );
  XNOR2_X1 U15281 ( .A(n11237), .B(n11289), .ZN(n11494) );
  NOR2_X1 U15282 ( .A1(n11011), .A2(n10415), .ZN(n10417) );
  XNOR2_X1 U15283 ( .A(n11771), .B(n673), .ZN(n10419) );
  XNOR2_X1 U15284 ( .A(n11494), .B(n10419), .ZN(n10420) );
  NOR2_X1 U15285 ( .A1(n10594), .A2(n10505), .ZN(n10422) );
  OAI21_X1 U15286 ( .B1(n10422), .B2(n2311), .A(n10936), .ZN(n10424) );
  NAND3_X1 U15287 ( .A1(n10934), .A2(n5198), .A3(n10931), .ZN(n10423) );
  OAI211_X1 U15288 ( .C1(n10936), .C2(n10425), .A(n10424), .B(n10423), .ZN(
        n12233) );
  NAND2_X2 U15291 ( .A1(n10429), .A2(n10430), .ZN(n12362) );
  XNOR2_X1 U15292 ( .A(n12233), .B(n12362), .ZN(n10432) );
  XNOR2_X1 U15293 ( .A(n10432), .B(n10431), .ZN(n10450) );
  NAND2_X1 U15294 ( .A1(n11301), .A2(n10762), .ZN(n10433) );
  NAND2_X1 U15295 ( .A1(n10434), .A2(n10433), .ZN(n10437) );
  NAND2_X1 U15297 ( .A1(n10435), .A2(n10762), .ZN(n10436) );
  XNOR2_X1 U15298 ( .A(n11414), .B(n11646), .ZN(n12087) );
  NAND2_X1 U15299 ( .A1(n10439), .A2(n10767), .ZN(n10440) );
  NAND2_X1 U15302 ( .A1(n10443), .A2(n10751), .ZN(n10448) );
  NAND3_X1 U15303 ( .A1(n10445), .A2(n10746), .A3(n10901), .ZN(n10446) );
  XNOR2_X1 U15304 ( .A(n11908), .B(n11412), .ZN(n11355) );
  XNOR2_X1 U15305 ( .A(n12087), .B(n11355), .ZN(n10449) );
  NAND2_X1 U15307 ( .A1(n10752), .A2(n10757), .ZN(n10453) );
  XNOR2_X1 U15309 ( .A(n12209), .B(n11782), .ZN(n11515) );
  NAND2_X1 U15310 ( .A1(n10729), .A2(n10457), .ZN(n10456) );
  NAND2_X1 U15311 ( .A1(n10456), .A2(n10481), .ZN(n10459) );
  NOR2_X1 U15312 ( .A1(n10457), .A2(n11190), .ZN(n10458) );
  XNOR2_X1 U15313 ( .A(n11515), .B(n11848), .ZN(n10476) );
  OAI21_X1 U15314 ( .B1(n10850), .B2(n11122), .A(n10460), .ZN(n10463) );
  NAND2_X1 U15316 ( .A1(n10740), .A2(n10860), .ZN(n10469) );
  NAND2_X1 U15317 ( .A1(n10862), .A2(n10860), .ZN(n10468) );
  NAND3_X1 U15318 ( .A1(n10465), .A2(n10861), .A3(n25230), .ZN(n10467) );
  XNOR2_X1 U15319 ( .A(n12147), .B(n11741), .ZN(n11992) );
  AOI21_X1 U15320 ( .B1(n11129), .B2(n11128), .A(n11130), .ZN(n10473) );
  AND2_X1 U15321 ( .A1(n11128), .A2(n10714), .ZN(n10841) );
  NAND2_X1 U15322 ( .A1(n10841), .A2(n10470), .ZN(n10471) );
  XNOR2_X1 U15323 ( .A(n12286), .B(n663), .ZN(n10474) );
  XNOR2_X1 U15324 ( .A(n11992), .B(n10474), .ZN(n10475) );
  XNOR2_X1 U15325 ( .A(n10475), .B(n10476), .ZN(n13170) );
  INV_X1 U15326 ( .A(n13170), .ZN(n10502) );
  XNOR2_X1 U15329 ( .A(n11542), .B(n12257), .ZN(n10485) );
  NAND2_X1 U15330 ( .A1(n10729), .A2(n10481), .ZN(n10483) );
  XNOR2_X1 U15331 ( .A(n12224), .B(n4164), .ZN(n10484) );
  XNOR2_X1 U15332 ( .A(n10485), .B(n10484), .ZN(n10501) );
  XNOR2_X1 U15333 ( .A(n10490), .B(n11659), .ZN(n11861) );
  OAI21_X1 U15334 ( .B1(n11340), .B2(n11338), .A(n10493), .ZN(n10494) );
  NAND2_X1 U15335 ( .A1(n11935), .A2(n10494), .ZN(n10499) );
  NAND2_X1 U15336 ( .A1(n10970), .A2(n10968), .ZN(n10604) );
  NAND2_X1 U15337 ( .A1(n10496), .A2(n10495), .ZN(n10498) );
  NAND2_X1 U15338 ( .A1(n10497), .A2(n10606), .ZN(n10605) );
  OAI211_X1 U15339 ( .C1(n10497), .C2(n10604), .A(n10498), .B(n10605), .ZN(
        n11746) );
  XNOR2_X1 U15340 ( .A(n10499), .B(n11746), .ZN(n11429) );
  XNOR2_X1 U15341 ( .A(n11861), .B(n11429), .ZN(n10500) );
  XNOR2_X2 U15342 ( .A(n10501), .B(n10500), .ZN(n13167) );
  NAND2_X1 U15343 ( .A1(n10951), .A2(n10952), .ZN(n10504) );
  NAND3_X1 U15344 ( .A1(n5107), .A2(n10698), .A3(n10702), .ZN(n10503) );
  NAND2_X1 U15345 ( .A1(n10934), .A2(n24470), .ZN(n10507) );
  NAND2_X1 U15346 ( .A1(n2311), .A2(n10505), .ZN(n10506) );
  AOI21_X1 U15347 ( .B1(n10507), .B2(n10506), .A(n10596), .ZN(n10511) );
  XNOR2_X1 U15349 ( .A(n11672), .B(n11396), .ZN(n12110) );
  XNOR2_X1 U15350 ( .A(n11504), .B(n12110), .ZN(n10530) );
  NOR2_X1 U15351 ( .A1(n11036), .A2(n10941), .ZN(n10512) );
  OAI22_X1 U15352 ( .A1(n10515), .A2(n10829), .B1(n10836), .B2(n10514), .ZN(
        n10522) );
  NAND3_X1 U15353 ( .A1(n10518), .A2(n10517), .A3(n10516), .ZN(n10519) );
  AOI21_X1 U15354 ( .B1(n10520), .B2(n10519), .A(n9279), .ZN(n10521) );
  NOR2_X1 U15355 ( .A1(n10522), .A2(n10521), .ZN(n11756) );
  XNOR2_X1 U15356 ( .A(n12276), .B(n11756), .ZN(n11975) );
  MUX2_X1 U15357 ( .A(n11518), .B(n11519), .S(n10523), .Z(n10527) );
  NOR2_X1 U15358 ( .A1(n11520), .A2(n11524), .ZN(n10524) );
  XNOR2_X1 U15359 ( .A(n12277), .B(n2757), .ZN(n10528) );
  XNOR2_X1 U15360 ( .A(n11975), .B(n10528), .ZN(n10529) );
  INV_X1 U15361 ( .A(n13165), .ZN(n11597) );
  OAI21_X1 U15362 ( .B1(n10532), .B2(n10531), .A(n11597), .ZN(n10569) );
  NAND2_X1 U15363 ( .A1(n11151), .A2(n11143), .ZN(n10536) );
  AND2_X1 U15364 ( .A1(n10885), .A2(n10886), .ZN(n10540) );
  NOR2_X1 U15365 ( .A1(n10884), .A2(n24345), .ZN(n10539) );
  OR2_X2 U15367 ( .A1(n10546), .A2(n10545), .ZN(n11433) );
  XNOR2_X1 U15368 ( .A(n12241), .B(n11433), .ZN(n11995) );
  NAND2_X1 U15369 ( .A1(n5107), .A2(n25233), .ZN(n10705) );
  NOR2_X1 U15370 ( .A1(n10951), .A2(n25231), .ZN(n10701) );
  INV_X1 U15371 ( .A(n10701), .ZN(n10547) );
  NAND2_X1 U15372 ( .A1(n10955), .A2(n2754), .ZN(n10550) );
  NAND2_X1 U15373 ( .A1(n10548), .A2(n10698), .ZN(n10549) );
  XNOR2_X1 U15374 ( .A(n11840), .B(n11838), .ZN(n12094) );
  XNOR2_X1 U15375 ( .A(n11995), .B(n12094), .ZN(n10566) );
  AND2_X1 U15376 ( .A1(n10552), .A2(n11157), .ZN(n10554) );
  NOR2_X1 U15377 ( .A1(n11157), .A2(n11158), .ZN(n10555) );
  NOR2_X1 U15378 ( .A1(n10661), .A2(n10558), .ZN(n10562) );
  OAI21_X1 U15379 ( .B1(n10556), .B2(n10654), .A(n25250), .ZN(n10561) );
  NAND3_X1 U15380 ( .A1(n10558), .A2(n10557), .A3(n10660), .ZN(n10560) );
  INV_X1 U15381 ( .A(n10660), .ZN(n10655) );
  XNOR2_X1 U15382 ( .A(n12200), .B(n21423), .ZN(n10563) );
  XNOR2_X1 U15383 ( .A(n10564), .B(n10563), .ZN(n10565) );
  NOR3_X1 U15384 ( .A1(n24373), .A2(n12719), .A3(n13167), .ZN(n10567) );
  NOR2_X1 U15385 ( .A1(n24373), .A2(n13170), .ZN(n13168) );
  NOR2_X1 U15386 ( .A1(n10567), .A2(n13168), .ZN(n10568) );
  INV_X1 U15387 ( .A(n10572), .ZN(n10573) );
  MUX2_X2 U15388 ( .A(n10576), .B(n10575), .S(n10574), .Z(n12019) );
  XNOR2_X1 U15389 ( .A(n12019), .B(n12351), .ZN(n12302) );
  MUX2_X1 U15390 ( .A(n11171), .B(n24957), .S(n11178), .Z(n10578) );
  MUX2_X1 U15391 ( .A(n11168), .B(n11170), .S(n24957), .Z(n10577) );
  XNOR2_X1 U15392 ( .A(n11289), .B(n11638), .ZN(n10579) );
  XNOR2_X1 U15393 ( .A(n12302), .B(n10579), .ZN(n10603) );
  NAND2_X1 U15394 ( .A1(n10585), .A2(n10584), .ZN(n10586) );
  NAND2_X1 U15395 ( .A1(n10589), .A2(n25507), .ZN(n10592) );
  XNOR2_X1 U15396 ( .A(n12129), .B(n12127), .ZN(n10601) );
  NAND3_X1 U15397 ( .A1(n10934), .A2(n24470), .A3(n10508), .ZN(n10599) );
  XNOR2_X1 U15398 ( .A(n10602), .B(n10603), .ZN(n13132) );
  NAND2_X1 U15399 ( .A1(n10605), .A2(n10604), .ZN(n10609) );
  INV_X1 U15400 ( .A(n10969), .ZN(n10966) );
  XNOR2_X1 U15401 ( .A(n12031), .B(n12362), .ZN(n12293) );
  AOI21_X1 U15402 ( .B1(n10613), .B2(n10611), .A(n10610), .ZN(n10619) );
  NAND3_X1 U15403 ( .A1(n10614), .A2(n10613), .A3(n10612), .ZN(n10615) );
  OAI21_X1 U15404 ( .B1(n10617), .B2(n10616), .A(n10615), .ZN(n10618) );
  NAND3_X1 U15406 ( .A1(n24340), .A2(n3868), .A3(n11216), .ZN(n10625) );
  XNOR2_X1 U15407 ( .A(n12370), .B(n10627), .ZN(n11986) );
  XNOR2_X1 U15408 ( .A(n11986), .B(n12293), .ZN(n10640) );
  NOR2_X1 U15409 ( .A1(n10793), .A2(n11201), .ZN(n11204) );
  OAI21_X1 U15410 ( .B1(n11204), .B2(n11196), .A(n11199), .ZN(n10629) );
  INV_X1 U15412 ( .A(n10632), .ZN(n11210) );
  NAND3_X1 U15413 ( .A1(n11205), .A2(n11207), .A3(n11338), .ZN(n10635) );
  OAI21_X1 U15414 ( .B1(n11205), .B2(n10819), .A(n10635), .ZN(n10636) );
  XNOR2_X1 U15415 ( .A(n12167), .B(n3164), .ZN(n10637) );
  XNOR2_X1 U15416 ( .A(n10638), .B(n10637), .ZN(n10639) );
  XNOR2_X1 U15417 ( .A(n24980), .B(n886), .ZN(n10647) );
  NAND2_X1 U15418 ( .A1(n10642), .A2(n11012), .ZN(n10644) );
  AND2_X1 U15419 ( .A1(n10643), .A2(n10644), .ZN(n10645) );
  INV_X1 U15420 ( .A(n12144), .ZN(n10646) );
  NAND2_X1 U15421 ( .A1(n10655), .A2(n10654), .ZN(n10656) );
  XNOR2_X1 U15422 ( .A(n12146), .B(n12414), .ZN(n11991) );
  INV_X1 U15423 ( .A(n11067), .ZN(n10667) );
  AND2_X1 U15424 ( .A1(n11064), .A2(n10662), .ZN(n10664) );
  NOR2_X1 U15425 ( .A1(n11068), .A2(n11067), .ZN(n10663) );
  OAI22_X1 U15426 ( .A1(n10665), .A2(n10664), .B1(n10663), .B2(n11071), .ZN(
        n10666) );
  OAI21_X1 U15427 ( .B1(n10667), .B2(n11064), .A(n10666), .ZN(n11243) );
  INV_X1 U15428 ( .A(n11243), .ZN(n12039) );
  NAND2_X1 U15430 ( .A1(n11215), .A2(n11216), .ZN(n10670) );
  XNOR2_X1 U15431 ( .A(n12152), .B(n12322), .ZN(n10671) );
  XNOR2_X1 U15432 ( .A(n10672), .B(n10671), .ZN(n12498) );
  NAND2_X1 U15433 ( .A1(n11163), .A2(n11158), .ZN(n10680) );
  NAND3_X1 U15434 ( .A1(n10674), .A2(n1453), .A3(n10673), .ZN(n10678) );
  INV_X1 U15435 ( .A(n10675), .ZN(n10677) );
  OAI21_X1 U15436 ( .B1(n10678), .B2(n10677), .A(n10676), .ZN(n10679) );
  INV_X1 U15437 ( .A(n11007), .ZN(n10688) );
  OAI211_X1 U15438 ( .C1(n2306), .C2(n24420), .A(n24622), .B(n10681), .ZN(
        n10687) );
  INV_X1 U15439 ( .A(n10682), .ZN(n10684) );
  NAND2_X1 U15440 ( .A1(n11006), .A2(n10685), .ZN(n10686) );
  XNOR2_X1 U15441 ( .A(n11717), .B(n10689), .ZN(n12156) );
  NAND2_X1 U15442 ( .A1(n11149), .A2(n11151), .ZN(n11888) );
  NAND3_X1 U15443 ( .A1(n714), .A2(n11884), .A3(n11143), .ZN(n10692) );
  NAND3_X1 U15444 ( .A1(n10690), .A2(n11147), .A3(n11885), .ZN(n10691) );
  NAND3_X1 U15445 ( .A1(n11888), .A2(n10692), .A3(n10691), .ZN(n11247) );
  XNOR2_X1 U15446 ( .A(n11247), .B(n11746), .ZN(n12311) );
  XNOR2_X1 U15447 ( .A(n12156), .B(n12311), .ZN(n10709) );
  NAND2_X1 U15448 ( .A1(n11054), .A2(n11499), .ZN(n10696) );
  NOR2_X1 U15449 ( .A1(n11057), .A2(n11009), .ZN(n10693) );
  NAND2_X1 U15450 ( .A1(n11059), .A2(n10693), .ZN(n10695) );
  INV_X1 U15451 ( .A(n11499), .ZN(n11053) );
  INV_X1 U15452 ( .A(n10698), .ZN(n10954) );
  XNOR2_X1 U15453 ( .A(n10707), .B(n10706), .ZN(n10708) );
  NOR2_X1 U15454 ( .A1(n12498), .A2(n13130), .ZN(n10710) );
  NOR2_X1 U15455 ( .A1(n5754), .A2(n10710), .ZN(n12426) );
  INV_X1 U15456 ( .A(n12663), .ZN(n10711) );
  NAND2_X1 U15457 ( .A1(n10713), .A2(n10712), .ZN(n10718) );
  NAND3_X1 U15459 ( .A1(n10838), .A2(n420), .A3(n10714), .ZN(n10715) );
  NAND4_X2 U15460 ( .A1(n10716), .A2(n10717), .A3(n10715), .A4(n10718), .ZN(
        n11795) );
  XNOR2_X1 U15461 ( .A(n11795), .B(n2005), .ZN(n10719) );
  AND2_X1 U15463 ( .A1(n10720), .A2(n11121), .ZN(n10721) );
  NAND2_X1 U15465 ( .A1(n11110), .A2(n10875), .ZN(n10726) );
  MUX2_X1 U15466 ( .A(n10729), .B(n10728), .S(n11190), .Z(n10735) );
  NAND2_X1 U15467 ( .A1(n11184), .A2(n10729), .ZN(n10733) );
  NAND3_X1 U15468 ( .A1(n10731), .A2(n10730), .A3(n10734), .ZN(n10732) );
  XNOR2_X1 U15469 ( .A(n12404), .B(n25236), .ZN(n11981) );
  AND2_X1 U15470 ( .A1(n10860), .A2(n25230), .ZN(n10739) );
  NOR2_X1 U15471 ( .A1(n10861), .A2(n25230), .ZN(n10738) );
  AOI22_X1 U15472 ( .A1(n10739), .A2(n10740), .B1(n10738), .B2(n10737), .ZN(
        n10742) );
  NAND3_X1 U15473 ( .A1(n10740), .A2(n10855), .A3(n10861), .ZN(n10741) );
  XNOR2_X1 U15474 ( .A(n12066), .B(n11756), .ZN(n12338) );
  XNOR2_X1 U15475 ( .A(n11981), .B(n12338), .ZN(n10744) );
  INV_X1 U15476 ( .A(n13150), .ZN(n13157) );
  NOR2_X1 U15477 ( .A1(n10904), .A2(n10907), .ZN(n10748) );
  AOI22_X1 U15478 ( .A1(n10749), .A2(n10751), .B1(n10748), .B2(n10905), .ZN(
        n10750) );
  NOR2_X1 U15479 ( .A1(n10753), .A2(n10752), .ZN(n10754) );
  INV_X1 U15480 ( .A(n10756), .ZN(n10758) );
  NOR2_X2 U15481 ( .A1(n10761), .A2(n10760), .ZN(n11581) );
  INV_X1 U15482 ( .A(n11301), .ZN(n11089) );
  INV_X1 U15483 ( .A(n10762), .ZN(n11305) );
  MUX2_X1 U15484 ( .A(n10764), .B(n10763), .S(n11091), .Z(n10765) );
  XNOR2_X1 U15485 ( .A(n11581), .B(n12375), .ZN(n11996) );
  XNOR2_X1 U15486 ( .A(n12341), .B(n11996), .ZN(n10786) );
  NOR2_X1 U15487 ( .A1(n11084), .A2(n10891), .ZN(n10768) );
  NOR2_X2 U15488 ( .A1(n10770), .A2(n10769), .ZN(n12121) );
  XNOR2_X1 U15489 ( .A(n10771), .B(n12121), .ZN(n10784) );
  OAI21_X1 U15490 ( .B1(n11101), .B2(n10911), .A(n10772), .ZN(n10781) );
  INV_X1 U15491 ( .A(n10773), .ZN(n10774) );
  NOR2_X1 U15492 ( .A1(n10775), .A2(n10774), .ZN(n10777) );
  NAND4_X1 U15493 ( .A1(n10778), .A2(n415), .A3(n10777), .A4(n10776), .ZN(
        n10780) );
  OAI211_X2 U15494 ( .C1(n10781), .C2(n10782), .A(n10780), .B(n10779), .ZN(
        n11765) );
  XNOR2_X1 U15495 ( .A(n11765), .B(n2805), .ZN(n10783) );
  XNOR2_X1 U15496 ( .A(n10784), .B(n10783), .ZN(n10785) );
  XNOR2_X1 U15497 ( .A(n10786), .B(n10785), .ZN(n13151) );
  OAI211_X1 U15499 ( .C1(n13157), .C2(n13152), .A(n13148), .B(n13130), .ZN(
        n10787) );
  NAND2_X1 U15500 ( .A1(n10788), .A2(n11195), .ZN(n10797) );
  INV_X1 U15501 ( .A(n10789), .ZN(n10790) );
  INV_X1 U15502 ( .A(n11196), .ZN(n10792) );
  NAND3_X1 U15503 ( .A1(n11201), .A2(n11199), .A3(n10792), .ZN(n10795) );
  NAND3_X1 U15504 ( .A1(n10793), .A2(n11196), .A3(n11199), .ZN(n10794) );
  XNOR2_X1 U15505 ( .A(n11951), .B(n12401), .ZN(n10809) );
  MUX2_X1 U15506 ( .A(n10800), .B(n10799), .S(n10798), .Z(n10802) );
  MUX2_X1 U15507 ( .A(n10803), .B(n10802), .S(n10801), .Z(n10807) );
  NOR2_X2 U15508 ( .A1(n10807), .A2(n10806), .ZN(n12334) );
  INV_X1 U15509 ( .A(n12334), .ZN(n10808) );
  XNOR2_X1 U15510 ( .A(n10809), .B(n10808), .ZN(n10828) );
  XNOR2_X1 U15512 ( .A(n11619), .B(n25236), .ZN(n10826) );
  NOR2_X1 U15513 ( .A1(n10967), .A2(n10969), .ZN(n10815) );
  NOR2_X1 U15514 ( .A1(n10970), .A2(n10968), .ZN(n10814) );
  NAND2_X1 U15515 ( .A1(n10816), .A2(n10970), .ZN(n10817) );
  XNOR2_X1 U15516 ( .A(n12112), .B(n2903), .ZN(n10824) );
  MUX2_X1 U15517 ( .A(n11342), .B(n10819), .S(n25025), .Z(n10823) );
  INV_X1 U15518 ( .A(n11205), .ZN(n11339) );
  NAND2_X1 U15519 ( .A1(n11342), .A2(n11207), .ZN(n10820) );
  MUX2_X1 U15520 ( .A(n10821), .B(n10820), .S(n10819), .Z(n10822) );
  OAI21_X2 U15521 ( .B1(n10823), .B2(n11339), .A(n10822), .ZN(n12397) );
  XNOR2_X1 U15522 ( .A(n10824), .B(n12397), .ZN(n10825) );
  XNOR2_X1 U15523 ( .A(n10825), .B(n10826), .ZN(n10827) );
  XNOR2_X1 U15524 ( .A(n10827), .B(n10828), .ZN(n12740) );
  INV_X1 U15525 ( .A(n12740), .ZN(n13101) );
  AOI22_X1 U15526 ( .A1(n10836), .A2(n10834), .B1(n10833), .B2(n10832), .ZN(
        n10835) );
  OAI21_X1 U15527 ( .B1(n10837), .B2(n10836), .A(n10835), .ZN(n12344) );
  XNOR2_X1 U15528 ( .A(n12344), .B(n11581), .ZN(n11666) );
  NAND2_X1 U15529 ( .A1(n10841), .A2(n11129), .ZN(n10842) );
  XNOR2_X1 U15530 ( .A(n12381), .B(n1951), .ZN(n10845) );
  XNOR2_X1 U15531 ( .A(n11666), .B(n10845), .ZN(n10883) );
  OR2_X1 U15532 ( .A1(n10848), .A2(n2244), .ZN(n10849) );
  OAI211_X1 U15533 ( .C1(n11125), .C2(n10850), .A(n10849), .B(n11124), .ZN(
        n10852) );
  NAND3_X1 U15534 ( .A1(n10856), .A2(n10855), .A3(n10854), .ZN(n10866) );
  NAND2_X1 U15536 ( .A1(n10862), .A2(n10861), .ZN(n10863) );
  XNOR2_X1 U15537 ( .A(n11703), .B(n12096), .ZN(n11602) );
  NAND4_X1 U15539 ( .A1(n10873), .A2(n10870), .A3(n10867), .A4(n9340), .ZN(
        n11115) );
  INV_X1 U15540 ( .A(n10870), .ZN(n10872) );
  NOR2_X1 U15541 ( .A1(n10872), .A2(n10871), .ZN(n10874) );
  NAND4_X1 U15542 ( .A1(n10875), .A2(n1494), .A3(n10874), .A4(n10873), .ZN(
        n10876) );
  OAI21_X2 U15543 ( .B1(n10877), .B2(n10878), .A(n10876), .ZN(n11766) );
  INV_X1 U15544 ( .A(n12383), .ZN(n10879) );
  XNOR2_X1 U15545 ( .A(n10879), .B(n11766), .ZN(n10880) );
  MUX2_X1 U15547 ( .A(n10887), .B(n10886), .S(n10885), .Z(n10888) );
  XNOR2_X1 U15548 ( .A(n12306), .B(n12127), .ZN(n11639) );
  INV_X1 U15549 ( .A(n11966), .ZN(n11457) );
  INV_X1 U15550 ( .A(n11086), .ZN(n10893) );
  NOR2_X1 U15551 ( .A1(n11085), .A2(n10891), .ZN(n10892) );
  XNOR2_X1 U15552 ( .A(n11457), .B(n12020), .ZN(n12354) );
  NAND2_X1 U15553 ( .A1(n11302), .A2(n11298), .ZN(n10897) );
  OAI21_X1 U15554 ( .B1(n10902), .B2(n10901), .A(n10900), .ZN(n10909) );
  OAI21_X1 U15555 ( .B1(n10905), .B2(n10904), .A(n10903), .ZN(n10906) );
  INV_X1 U15556 ( .A(n10906), .ZN(n10908) );
  XNOR2_X1 U15558 ( .A(n11627), .B(n12183), .ZN(n10916) );
  NAND3_X1 U15559 ( .A1(n11099), .A2(n10911), .A3(n11101), .ZN(n10912) );
  INV_X1 U15560 ( .A(n2795), .ZN(n23191) );
  XNOR2_X1 U15561 ( .A(n12357), .B(n23191), .ZN(n10915) );
  XNOR2_X1 U15562 ( .A(n10916), .B(n10915), .ZN(n10917) );
  MUX2_X1 U15563 ( .A(n13101), .B(n13102), .S(n13185), .Z(n11021) );
  NAND2_X1 U15564 ( .A1(n10922), .A2(n11520), .ZN(n10919) );
  INV_X1 U15566 ( .A(n2991), .ZN(n21079) );
  XNOR2_X1 U15567 ( .A(n12388), .B(n21079), .ZN(n10923) );
  INV_X1 U15568 ( .A(n11747), .ZN(n11942) );
  NAND2_X1 U15569 ( .A1(n10925), .A2(n10924), .ZN(n10929) );
  OAI21_X1 U15570 ( .B1(n10927), .B2(n10990), .A(n10926), .ZN(n10928) );
  INV_X1 U15571 ( .A(n10931), .ZN(n10932) );
  NAND2_X1 U15572 ( .A1(n10932), .A2(n10935), .ZN(n10933) );
  OAI21_X1 U15573 ( .B1(n11171), .B2(n11175), .A(n10937), .ZN(n10938) );
  XNOR2_X1 U15574 ( .A(n11749), .B(n12389), .ZN(n10947) );
  INV_X1 U15575 ( .A(n11040), .ZN(n10946) );
  NAND2_X1 U15576 ( .A1(n416), .A2(n10942), .ZN(n10943) );
  XNOR2_X1 U15577 ( .A(n10947), .B(n24915), .ZN(n10948) );
  XNOR2_X1 U15578 ( .A(n10949), .B(n10948), .ZN(n13187) );
  NAND3_X1 U15579 ( .A1(n10955), .A2(n10954), .A3(n25232), .ZN(n10956) );
  XNOR2_X1 U15581 ( .A(n24401), .B(n812), .ZN(n10959) );
  INV_X1 U15582 ( .A(n12146), .ZN(n11555) );
  XNOR2_X1 U15583 ( .A(n10959), .B(n11555), .ZN(n10977) );
  NAND2_X1 U15584 ( .A1(n714), .A2(n24480), .ZN(n10964) );
  NOR2_X1 U15585 ( .A1(n10961), .A2(n11884), .ZN(n10960) );
  INV_X1 U15587 ( .A(n10961), .ZN(n11148) );
  NOR2_X1 U15588 ( .A1(n25497), .A2(n10969), .ZN(n10976) );
  OAI21_X1 U15589 ( .B1(n10967), .B2(n10966), .A(n10497), .ZN(n10975) );
  NAND2_X1 U15590 ( .A1(n10969), .A2(n10968), .ZN(n10973) );
  INV_X1 U15591 ( .A(n10970), .ZN(n10972) );
  MUX2_X1 U15592 ( .A(n10973), .B(n10972), .S(n25497), .Z(n10974) );
  XNOR2_X1 U15593 ( .A(n11897), .B(n12325), .ZN(n12210) );
  XNOR2_X1 U15594 ( .A(n10977), .B(n12210), .ZN(n10988) );
  NOR2_X1 U15595 ( .A1(n11059), .A2(n11052), .ZN(n11498) );
  NOR2_X1 U15596 ( .A1(n10978), .A2(n11498), .ZN(n10981) );
  AOI21_X1 U15597 ( .B1(n11054), .B2(n11009), .A(n11053), .ZN(n10979) );
  OAI21_X1 U15598 ( .B1(n11009), .B2(n410), .A(n10979), .ZN(n10980) );
  NAND2_X1 U15599 ( .A1(n417), .A2(n11157), .ZN(n11166) );
  NOR2_X1 U15600 ( .A1(n4737), .A2(n11157), .ZN(n10982) );
  AOI22_X1 U15601 ( .A1(n10982), .A2(n10985), .B1(n11158), .B2(n11157), .ZN(
        n10984) );
  NAND3_X1 U15602 ( .A1(n417), .A2(n10985), .A3(n11160), .ZN(n10983) );
  OAI211_X2 U15603 ( .C1(n11166), .C2(n10985), .A(n10984), .B(n10983), .ZN(
        n12413) );
  XNOR2_X1 U15604 ( .A(n11960), .B(n12413), .ZN(n10986) );
  XNOR2_X1 U15605 ( .A(n12410), .B(n10986), .ZN(n10987) );
  NOR2_X1 U15606 ( .A1(n10989), .A2(n10994), .ZN(n10991) );
  OAI21_X1 U15607 ( .B1(n10992), .B2(n10991), .A(n10990), .ZN(n10999) );
  NOR3_X1 U15608 ( .A1(n24118), .A2(n3606), .A3(n10993), .ZN(n10997) );
  NOR2_X1 U15609 ( .A1(n10997), .A2(n10996), .ZN(n10998) );
  NAND3_X1 U15610 ( .A1(n11068), .A2(n11069), .A3(n11064), .ZN(n11000) );
  XNOR2_X1 U15611 ( .A(n11907), .B(n25234), .ZN(n11608) );
  XNOR2_X1 U15612 ( .A(n11563), .B(n12295), .ZN(n11648) );
  XNOR2_X1 U15613 ( .A(n11608), .B(n11648), .ZN(n11019) );
  XNOR2_X1 U15614 ( .A(n11736), .B(n19392), .ZN(n11017) );
  AOI21_X1 U15615 ( .B1(n11010), .B2(n11050), .A(n11046), .ZN(n11015) );
  AOI21_X1 U15616 ( .B1(n11013), .B2(n11012), .A(n11044), .ZN(n11014) );
  NOR2_X2 U15617 ( .A1(n11015), .A2(n11014), .ZN(n12363) );
  XNOR2_X1 U15618 ( .A(n12363), .B(n25371), .ZN(n11016) );
  XNOR2_X1 U15619 ( .A(n11017), .B(n11016), .ZN(n11018) );
  NAND3_X1 U15622 ( .A1(n11026), .A2(n11525), .A3(n25060), .ZN(n11028) );
  NAND3_X1 U15623 ( .A1(n11529), .A2(n1332), .A3(n11524), .ZN(n11027) );
  XNOR2_X1 U15624 ( .A(n12234), .B(n17960), .ZN(n11030) );
  XNOR2_X1 U15625 ( .A(n12249), .B(n12297), .ZN(n11029) );
  XNOR2_X1 U15626 ( .A(n11030), .B(n11029), .ZN(n11043) );
  XNOR2_X1 U15627 ( .A(n12233), .B(n11561), .ZN(n11692) );
  XNOR2_X1 U15628 ( .A(n11983), .B(n12365), .ZN(n11041) );
  XNOR2_X1 U15629 ( .A(n11692), .B(n11041), .ZN(n11042) );
  XNOR2_X2 U15630 ( .A(n11042), .B(n11043), .ZN(n13144) );
  INV_X1 U15631 ( .A(n13144), .ZN(n13138) );
  OAI21_X1 U15632 ( .B1(n11045), .B2(n4531), .A(n11044), .ZN(n11048) );
  NAND3_X1 U15633 ( .A1(n11059), .A2(n11053), .A3(n11052), .ZN(n11056) );
  XNOR2_X1 U15634 ( .A(n12197), .B(n11706), .ZN(n11060) );
  XNOR2_X1 U15635 ( .A(n11060), .B(n11061), .ZN(n11080) );
  NAND2_X1 U15636 ( .A1(n10347), .A2(n11064), .ZN(n11066) );
  OR3_X1 U15637 ( .A1(n11064), .A2(n25203), .A3(n11062), .ZN(n11065) );
  NAND2_X1 U15639 ( .A1(n11068), .A2(n11067), .ZN(n11073) );
  NAND2_X1 U15640 ( .A1(n11070), .A2(n11069), .ZN(n11072) );
  AOI21_X1 U15641 ( .B1(n11073), .B2(n11072), .A(n11071), .ZN(n11074) );
  INV_X1 U15642 ( .A(n11076), .ZN(n12343) );
  XNOR2_X1 U15643 ( .A(n12343), .B(n12196), .ZN(n11078) );
  XNOR2_X1 U15644 ( .A(n12200), .B(n688), .ZN(n11077) );
  XNOR2_X1 U15645 ( .A(n11078), .B(n11077), .ZN(n11079) );
  XNOR2_X1 U15646 ( .A(n11079), .B(n11080), .ZN(n13140) );
  INV_X1 U15647 ( .A(n13140), .ZN(n12728) );
  NOR2_X1 U15648 ( .A1(n3119), .A2(n11081), .ZN(n11083) );
  XNOR2_X1 U15649 ( .A(n11087), .B(n11088), .ZN(n11108) );
  OAI21_X1 U15650 ( .B1(n11089), .B2(n11092), .A(n419), .ZN(n11095) );
  OAI211_X1 U15651 ( .C1(n11090), .C2(n11091), .A(n11305), .B(n11298), .ZN(
        n11094) );
  NOR2_X1 U15652 ( .A1(n11092), .A2(n11091), .ZN(n11093) );
  XNOR2_X1 U15653 ( .A(n24027), .B(n12209), .ZN(n11900) );
  NAND2_X1 U15654 ( .A1(n11096), .A2(n1552), .ZN(n11098) );
  NAND2_X1 U15655 ( .A1(n11099), .A2(n415), .ZN(n11097) );
  NAND2_X1 U15657 ( .A1(n11100), .A2(n11099), .ZN(n11104) );
  XNOR2_X1 U15658 ( .A(n12212), .B(n1754), .ZN(n11106) );
  XNOR2_X1 U15659 ( .A(n11900), .B(n11106), .ZN(n11107) );
  XNOR2_X1 U15660 ( .A(n11108), .B(n11107), .ZN(n11109) );
  NAND2_X1 U15661 ( .A1(n12728), .A2(n11109), .ZN(n12437) );
  AOI21_X1 U15662 ( .B1(n11117), .B2(n11111), .A(n11110), .ZN(n11120) );
  AOI21_X1 U15663 ( .B1(n11116), .B2(n11112), .A(n11113), .ZN(n11119) );
  OAI211_X1 U15664 ( .C1(n11117), .C2(n11116), .A(n11115), .B(n11114), .ZN(
        n11118) );
  XNOR2_X1 U15665 ( .A(n12314), .B(n11715), .ZN(n11137) );
  AOI22_X1 U15666 ( .A1(n11126), .A2(n11125), .B1(n11124), .B2(n11123), .ZN(
        n11127) );
  NOR2_X1 U15667 ( .A1(n11129), .A2(n11128), .ZN(n11134) );
  INV_X1 U15668 ( .A(n11131), .ZN(n11132) );
  OAI211_X2 U15669 ( .C1(n11135), .C2(n11134), .A(n11133), .B(n11132), .ZN(
        n12221) );
  XNOR2_X1 U15670 ( .A(n12221), .B(n12219), .ZN(n11136) );
  XNOR2_X1 U15671 ( .A(n11137), .B(n11136), .ZN(n11141) );
  XNOR2_X1 U15672 ( .A(n12391), .B(n12224), .ZN(n11139) );
  XNOR2_X1 U15673 ( .A(n12255), .B(n1869), .ZN(n11138) );
  XNOR2_X1 U15674 ( .A(n11139), .B(n11138), .ZN(n11140) );
  XNOR2_X1 U15675 ( .A(n11141), .B(n11140), .ZN(n13136) );
  INV_X1 U15676 ( .A(n13136), .ZN(n13143) );
  NAND2_X1 U15677 ( .A1(n13139), .A2(n13143), .ZN(n11142) );
  NAND3_X1 U15679 ( .A1(n11145), .A2(n11146), .A3(n11143), .ZN(n11144) );
  OAI21_X1 U15680 ( .B1(n11147), .B2(n11145), .A(n11144), .ZN(n11156) );
  OAI21_X1 U15681 ( .B1(n11147), .B2(n11146), .A(n4998), .ZN(n11155) );
  NOR2_X1 U15682 ( .A1(n11148), .A2(n11151), .ZN(n11150) );
  NAND2_X1 U15683 ( .A1(n11150), .A2(n11149), .ZN(n11154) );
  NAND3_X1 U15684 ( .A1(n714), .A2(n24479), .A3(n11151), .ZN(n11153) );
  NOR2_X1 U15685 ( .A1(n1358), .A2(n11157), .ZN(n11162) );
  NOR2_X1 U15686 ( .A1(n11159), .A2(n11158), .ZN(n11161) );
  OAI21_X1 U15687 ( .B1(n11162), .B2(n11161), .A(n11160), .ZN(n11165) );
  XNOR2_X1 U15688 ( .A(n12065), .B(n11977), .ZN(n12193) );
  XNOR2_X1 U15689 ( .A(n11167), .B(n12193), .ZN(n11183) );
  AND2_X1 U15691 ( .A1(n11171), .A2(n1338), .ZN(n11173) );
  NAND2_X1 U15692 ( .A1(n11178), .A2(n11173), .ZN(n11177) );
  OAI211_X2 U15693 ( .C1(n11179), .C2(n11178), .A(n11177), .B(n11176), .ZN(
        n11689) );
  XNOR2_X1 U15696 ( .A(n11181), .B(n11180), .ZN(n11182) );
  NAND2_X1 U15698 ( .A1(n13138), .A2(n12455), .ZN(n11222) );
  INV_X1 U15699 ( .A(n11370), .ZN(n11191) );
  INV_X1 U15700 ( .A(n11184), .ZN(n11187) );
  INV_X1 U15701 ( .A(n11185), .ZN(n11186) );
  NAND2_X1 U15702 ( .A1(n11187), .A2(n11186), .ZN(n11188) );
  OAI22_X1 U15703 ( .A1(n11191), .A2(n11190), .B1(n11189), .B2(n11188), .ZN(
        n11192) );
  XNOR2_X1 U15704 ( .A(n11192), .B(n2990), .ZN(n11193) );
  XNOR2_X1 U15705 ( .A(n11194), .B(n11193), .ZN(n11221) );
  INV_X1 U15706 ( .A(n11201), .ZN(n11197) );
  OAI21_X1 U15707 ( .B1(n11197), .B2(n11196), .A(n10790), .ZN(n11203) );
  NAND2_X1 U15709 ( .A1(n25025), .A2(n11205), .ZN(n11206) );
  NAND2_X1 U15710 ( .A1(n11210), .A2(n11207), .ZN(n11208) );
  MUX2_X1 U15711 ( .A(n11214), .B(n24340), .S(n11212), .Z(n11219) );
  XNOR2_X1 U15712 ( .A(n12181), .B(n11880), .ZN(n11220) );
  XNOR2_X1 U15713 ( .A(n11220), .B(n11221), .ZN(n12433) );
  INV_X1 U15715 ( .A(n14156), .ZN(n13780) );
  XNOR2_X1 U15717 ( .A(n12189), .B(n12397), .ZN(n12064) );
  XNOR2_X1 U15718 ( .A(n11619), .B(n11795), .ZN(n11759) );
  XNOR2_X1 U15719 ( .A(n12064), .B(n11759), .ZN(n11227) );
  XNOR2_X1 U15720 ( .A(n12066), .B(n12401), .ZN(n11816) );
  INV_X1 U15721 ( .A(n23476), .ZN(n20840) );
  XNOR2_X1 U15722 ( .A(n11816), .B(n11225), .ZN(n11226) );
  XNOR2_X1 U15723 ( .A(n11227), .B(n11226), .ZN(n12541) );
  XNOR2_X1 U15724 ( .A(n12031), .B(n12363), .ZN(n11833) );
  INV_X1 U15725 ( .A(n11833), .ZN(n11228) );
  XNOR2_X1 U15726 ( .A(n12248), .B(n25234), .ZN(n12030) );
  XNOR2_X1 U15727 ( .A(n11228), .B(n12030), .ZN(n11231) );
  XNOR2_X1 U15728 ( .A(n12233), .B(n11736), .ZN(n11535) );
  XNOR2_X1 U15729 ( .A(n11735), .B(n20690), .ZN(n11229) );
  XNOR2_X1 U15730 ( .A(n11535), .B(n11229), .ZN(n11230) );
  INV_X1 U15731 ( .A(n11703), .ZN(n12377) );
  XNOR2_X1 U15732 ( .A(n12377), .B(n11766), .ZN(n11232) );
  XNOR2_X1 U15733 ( .A(n11232), .B(n11812), .ZN(n11236) );
  XNOR2_X1 U15734 ( .A(n11765), .B(n12201), .ZN(n11234) );
  XNOR2_X1 U15735 ( .A(n12200), .B(n881), .ZN(n11233) );
  XNOR2_X1 U15736 ( .A(n11234), .B(n11233), .ZN(n11235) );
  XNOR2_X1 U15737 ( .A(n11627), .B(n11638), .ZN(n11724) );
  XNOR2_X1 U15738 ( .A(n12019), .B(n12357), .ZN(n11456) );
  XNOR2_X1 U15739 ( .A(n11456), .B(n11724), .ZN(n11241) );
  XNOR2_X1 U15740 ( .A(n12184), .B(n12020), .ZN(n11239) );
  INV_X1 U15741 ( .A(n11237), .ZN(n12180) );
  XNOR2_X1 U15742 ( .A(n12180), .B(n1865), .ZN(n11238) );
  XNOR2_X1 U15743 ( .A(n11239), .B(n11238), .ZN(n11240) );
  XNOR2_X1 U15744 ( .A(n11240), .B(n11241), .ZN(n12540) );
  XNOR2_X1 U15745 ( .A(n24401), .B(n11242), .ZN(n11745) );
  XNOR2_X1 U15746 ( .A(n12410), .B(n11243), .ZN(n11822) );
  XNOR2_X1 U15747 ( .A(n11822), .B(n11745), .ZN(n11246) );
  XNOR2_X1 U15748 ( .A(n12209), .B(n3118), .ZN(n11244) );
  XNOR2_X1 U15749 ( .A(n12413), .B(n12207), .ZN(n12038) );
  XNOR2_X1 U15750 ( .A(n12038), .B(n11244), .ZN(n11245) );
  XNOR2_X1 U15751 ( .A(n12218), .B(n12388), .ZN(n11718) );
  XNOR2_X1 U15752 ( .A(n11718), .B(n11827), .ZN(n11250) );
  XNOR2_X1 U15753 ( .A(n11749), .B(n12224), .ZN(n11545) );
  XNOR2_X1 U15754 ( .A(n11248), .B(n11545), .ZN(n11249) );
  MUX2_X1 U15755 ( .A(n13217), .B(n13216), .S(n12767), .Z(n11251) );
  NOR2_X1 U15756 ( .A1(n11251), .A2(n24512), .ZN(n11252) );
  XNOR2_X1 U15757 ( .A(n11253), .B(n11914), .ZN(n11842) );
  XNOR2_X1 U15758 ( .A(n12096), .B(n11582), .ZN(n12198) );
  XNOR2_X1 U15759 ( .A(n11842), .B(n12198), .ZN(n11257) );
  XNOR2_X1 U15760 ( .A(n11838), .B(n1831), .ZN(n11255) );
  XNOR2_X1 U15761 ( .A(n11704), .B(n12381), .ZN(n11254) );
  XNOR2_X1 U15762 ( .A(n11255), .B(n11254), .ZN(n11256) );
  XNOR2_X1 U15763 ( .A(n12249), .B(n11776), .ZN(n11905) );
  XNOR2_X1 U15764 ( .A(n11607), .B(n11907), .ZN(n11693) );
  XNOR2_X1 U15765 ( .A(n11693), .B(n11905), .ZN(n11261) );
  XNOR2_X1 U15766 ( .A(n12363), .B(n3062), .ZN(n11259) );
  XNOR2_X1 U15767 ( .A(n11646), .B(n11564), .ZN(n11258) );
  XNOR2_X1 U15768 ( .A(n11259), .B(n11258), .ZN(n11260) );
  XNOR2_X1 U15769 ( .A(n11261), .B(n11260), .ZN(n11287) );
  INV_X1 U15770 ( .A(n11616), .ZN(n11262) );
  XNOR2_X1 U15771 ( .A(n12226), .B(n11262), .ZN(n11716) );
  XNOR2_X1 U15772 ( .A(n12313), .B(n12255), .ZN(n11893) );
  XNOR2_X1 U15773 ( .A(n11716), .B(n11893), .ZN(n11267) );
  XNOR2_X1 U15774 ( .A(n11659), .B(n12389), .ZN(n11265) );
  XNOR2_X1 U15775 ( .A(n12225), .B(n681), .ZN(n11264) );
  XNOR2_X1 U15776 ( .A(n11265), .B(n11264), .ZN(n11266) );
  XNOR2_X1 U15777 ( .A(n11267), .B(n11266), .ZN(n13011) );
  XNOR2_X1 U15778 ( .A(n12186), .B(n11640), .ZN(n11269) );
  XNOR2_X1 U15779 ( .A(n11268), .B(n11492), .ZN(n11878) );
  INV_X1 U15780 ( .A(n11878), .ZN(n11858) );
  XNOR2_X1 U15781 ( .A(n11858), .B(n11269), .ZN(n11273) );
  XNOR2_X1 U15782 ( .A(n12183), .B(n12357), .ZN(n11271) );
  XNOR2_X1 U15783 ( .A(n11698), .B(n1745), .ZN(n11270) );
  XNOR2_X1 U15784 ( .A(n11271), .B(n11270), .ZN(n11272) );
  INV_X1 U15785 ( .A(n13013), .ZN(n13017) );
  XNOR2_X1 U15787 ( .A(n12333), .B(n12275), .ZN(n11924) );
  INV_X1 U15788 ( .A(n11924), .ZN(n11275) );
  XNOR2_X1 U15789 ( .A(n25027), .B(n11274), .ZN(n12190) );
  XNOR2_X1 U15790 ( .A(n11275), .B(n12190), .ZN(n11279) );
  INV_X1 U15791 ( .A(n11686), .ZN(n11618) );
  XNOR2_X1 U15792 ( .A(n11672), .B(n11618), .ZN(n11277) );
  XNOR2_X1 U15793 ( .A(n12401), .B(n2100), .ZN(n11276) );
  XNOR2_X1 U15794 ( .A(n11277), .B(n11276), .ZN(n11278) );
  XNOR2_X2 U15795 ( .A(n11279), .B(n11278), .ZN(n13245) );
  XNOR2_X1 U15796 ( .A(n12101), .B(n2050), .ZN(n11280) );
  XNOR2_X1 U15797 ( .A(n11280), .B(n12410), .ZN(n11283) );
  INV_X1 U15798 ( .A(n11653), .ZN(n11281) );
  XNOR2_X1 U15799 ( .A(n12283), .B(n11281), .ZN(n11282) );
  XNOR2_X1 U15800 ( .A(n11282), .B(n11283), .ZN(n11286) );
  INV_X1 U15801 ( .A(n11284), .ZN(n11285) );
  XNOR2_X1 U15802 ( .A(n11285), .B(n11286), .ZN(n12560) );
  INV_X1 U15803 ( .A(n12560), .ZN(n12808) );
  NOR2_X1 U15804 ( .A1(n25199), .A2(n13246), .ZN(n11288) );
  XNOR2_X1 U15805 ( .A(n12003), .B(n11289), .ZN(n12074) );
  XNOR2_X1 U15807 ( .A(n11637), .B(n11568), .ZN(n11439) );
  XNOR2_X1 U15808 ( .A(n24990), .B(n11439), .ZN(n11293) );
  XNOR2_X1 U15809 ( .A(n12023), .B(n12128), .ZN(n11856) );
  XNOR2_X1 U15810 ( .A(n11698), .B(n1364), .ZN(n11291) );
  XNOR2_X1 U15811 ( .A(n11856), .B(n11291), .ZN(n11292) );
  XNOR2_X1 U15812 ( .A(n11292), .B(n11293), .ZN(n13228) );
  XNOR2_X1 U15814 ( .A(n11689), .B(n729), .ZN(n11294) );
  XNOR2_X1 U15815 ( .A(n11294), .B(n11618), .ZN(n11296) );
  XNOR2_X1 U15816 ( .A(n11296), .B(n12114), .ZN(n11309) );
  NOR2_X1 U15817 ( .A1(n11302), .A2(n11301), .ZN(n11303) );
  NAND2_X1 U15818 ( .A1(n11303), .A2(n11305), .ZN(n11304) );
  XNOR2_X1 U15819 ( .A(n12065), .B(n12134), .ZN(n11868) );
  XNOR2_X1 U15820 ( .A(n25090), .B(n11561), .ZN(n11413) );
  XNOR2_X1 U15821 ( .A(n12088), .B(n11413), .ZN(n11313) );
  XNOR2_X1 U15822 ( .A(n11607), .B(n2745), .ZN(n11311) );
  XNOR2_X1 U15823 ( .A(n11851), .B(n11311), .ZN(n11312) );
  INV_X1 U15824 ( .A(n12197), .ZN(n11314) );
  XNOR2_X1 U15825 ( .A(n11314), .B(n12122), .ZN(n11510) );
  INV_X1 U15826 ( .A(n11510), .ZN(n11839) );
  XNOR2_X1 U15827 ( .A(n11839), .B(n12095), .ZN(n11318) );
  XNOR2_X1 U15828 ( .A(n11704), .B(n11706), .ZN(n11316) );
  XNOR2_X1 U15829 ( .A(n11316), .B(n11315), .ZN(n11317) );
  NOR2_X1 U15830 ( .A1(n12993), .A2(n24750), .ZN(n11319) );
  XNOR2_X1 U15832 ( .A(n25087), .B(n11959), .ZN(n11320) );
  XNOR2_X1 U15833 ( .A(n12151), .B(n12212), .ZN(n11516) );
  INV_X1 U15834 ( .A(n11516), .ZN(n11849) );
  INV_X1 U15835 ( .A(n11782), .ZN(n11322) );
  XNOR2_X1 U15836 ( .A(n12214), .B(n11322), .ZN(n12106) );
  INV_X1 U15837 ( .A(n12159), .ZN(n12260) );
  XNOR2_X1 U15838 ( .A(n12221), .B(n12260), .ZN(n11863) );
  XNOR2_X1 U15840 ( .A(n11616), .B(n21964), .ZN(n11324) );
  XNOR2_X1 U15841 ( .A(n25048), .B(n11324), .ZN(n11327) );
  XNOR2_X1 U15842 ( .A(n11715), .B(n11660), .ZN(n11426) );
  XNOR2_X1 U15843 ( .A(n11787), .B(n11426), .ZN(n11326) );
  NOR2_X1 U15844 ( .A1(n4587), .A2(n12791), .ZN(n11329) );
  NAND2_X1 U15845 ( .A1(n11329), .A2(n25080), .ZN(n11330) );
  INV_X1 U15846 ( .A(n11771), .ZN(n11879) );
  XNOR2_X1 U15847 ( .A(n11879), .B(n12130), .ZN(n12267) );
  XNOR2_X1 U15848 ( .A(n11628), .B(n11440), .ZN(n11332) );
  XNOR2_X1 U15849 ( .A(n12267), .B(n11332), .ZN(n11335) );
  XNOR2_X1 U15850 ( .A(n12355), .B(n12127), .ZN(n11570) );
  XNOR2_X1 U15851 ( .A(n12023), .B(n1801), .ZN(n11333) );
  XNOR2_X1 U15852 ( .A(n11570), .B(n11333), .ZN(n11334) );
  XNOR2_X2 U15853 ( .A(n11335), .B(n11334), .ZN(n13211) );
  XNOR2_X1 U15854 ( .A(n11892), .B(n12391), .ZN(n11789) );
  XNOR2_X1 U15855 ( .A(n11336), .B(n11424), .ZN(n11337) );
  XNOR2_X1 U15856 ( .A(n11337), .B(n11789), .ZN(n11345) );
  MUX2_X1 U15857 ( .A(n11340), .B(n11339), .S(n11338), .Z(n11939) );
  INV_X1 U15858 ( .A(n11935), .ZN(n11341) );
  AOI21_X1 U15859 ( .B1(n11939), .B2(n11342), .A(n11341), .ZN(n12263) );
  INV_X1 U15860 ( .A(n12263), .ZN(n12161) );
  XNOR2_X1 U15861 ( .A(n11343), .B(n12161), .ZN(n11344) );
  XNOR2_X1 U15862 ( .A(n11345), .B(n11344), .ZN(n11350) );
  XNOR2_X1 U15863 ( .A(n12065), .B(n11396), .ZN(n11347) );
  XNOR2_X1 U15864 ( .A(n12277), .B(n21944), .ZN(n11346) );
  XNOR2_X1 U15865 ( .A(n12276), .B(n12396), .ZN(n12136) );
  INV_X1 U15866 ( .A(n12136), .ZN(n11348) );
  XNOR2_X1 U15867 ( .A(n11349), .B(n25047), .ZN(n11684) );
  AOI21_X1 U15868 ( .B1(n13211), .B2(n13206), .A(n11684), .ZN(n11367) );
  INV_X1 U15869 ( .A(n11350), .ZN(n13004) );
  XNOR2_X1 U15870 ( .A(n12282), .B(n11385), .ZN(n11351) );
  XNOR2_X1 U15871 ( .A(n11351), .B(n11991), .ZN(n11354) );
  XNOR2_X1 U15872 ( .A(n12212), .B(n1920), .ZN(n11352) );
  INV_X1 U15873 ( .A(n12150), .ZN(n12408) );
  XNOR2_X1 U15874 ( .A(n12408), .B(n12286), .ZN(n11781) );
  XNOR2_X1 U15875 ( .A(n11352), .B(n11781), .ZN(n11353) );
  XNOR2_X1 U15876 ( .A(n11353), .B(n11354), .ZN(n13000) );
  NAND2_X1 U15877 ( .A1(n13004), .A2(n13000), .ZN(n11361) );
  INV_X1 U15878 ( .A(n11355), .ZN(n12247) );
  XNOR2_X1 U15879 ( .A(n12247), .B(n11356), .ZN(n11359) );
  XNOR2_X1 U15880 ( .A(n12234), .B(n2033), .ZN(n11357) );
  XNOR2_X1 U15881 ( .A(n11986), .B(n11357), .ZN(n11358) );
  NAND2_X1 U15882 ( .A1(n11361), .A2(n11360), .ZN(n12892) );
  XNOR2_X1 U15883 ( .A(n11581), .B(n12241), .ZN(n12124) );
  XNOR2_X1 U15884 ( .A(n12197), .B(n888), .ZN(n11362) );
  XNOR2_X1 U15885 ( .A(n12124), .B(n11362), .ZN(n11365) );
  XNOR2_X1 U15886 ( .A(n11761), .B(n12378), .ZN(n11800) );
  XNOR2_X1 U15887 ( .A(n12375), .B(n25016), .ZN(n11363) );
  XNOR2_X1 U15888 ( .A(n11800), .B(n11363), .ZN(n11364) );
  OAI21_X1 U15889 ( .B1(n13213), .B2(n13206), .A(n13000), .ZN(n11366) );
  INV_X1 U15890 ( .A(n11411), .ZN(n14290) );
  AOI21_X1 U15891 ( .B1(n13951), .B2(n14294), .A(n14290), .ZN(n11368) );
  NAND2_X1 U15892 ( .A1(n11369), .A2(n11368), .ZN(n14686) );
  XNOR2_X1 U15893 ( .A(n11628), .B(n12129), .ZN(n11375) );
  AND3_X1 U15894 ( .A1(n24913), .A2(n11371), .A3(n2211), .ZN(n11373) );
  AOI21_X1 U15895 ( .B1(n11371), .B2(n24913), .A(n2211), .ZN(n11372) );
  NOR2_X1 U15896 ( .A1(n11373), .A2(n11372), .ZN(n11374) );
  XNOR2_X1 U15897 ( .A(n11375), .B(n11374), .ZN(n11379) );
  XNOR2_X1 U15898 ( .A(n11638), .B(n12306), .ZN(n11377) );
  XNOR2_X1 U15899 ( .A(n11440), .B(n11967), .ZN(n11376) );
  XNOR2_X1 U15900 ( .A(n11376), .B(n11377), .ZN(n11378) );
  XNOR2_X1 U15901 ( .A(n11414), .B(n12364), .ZN(n11380) );
  XNOR2_X1 U15902 ( .A(n11946), .B(n11380), .ZN(n11383) );
  XNOR2_X1 U15903 ( .A(n11735), .B(n860), .ZN(n11381) );
  XNOR2_X1 U15904 ( .A(n12370), .B(n12297), .ZN(n11610) );
  XNOR2_X1 U15905 ( .A(n11610), .B(n11381), .ZN(n11382) );
  INV_X1 U15906 ( .A(n13027), .ZN(n13030) );
  XNOR2_X1 U15907 ( .A(n12414), .B(n853), .ZN(n11384) );
  XNOR2_X1 U15908 ( .A(n11384), .B(n12152), .ZN(n11387) );
  XNOR2_X1 U15909 ( .A(n11385), .B(n12324), .ZN(n11386) );
  XNOR2_X1 U15910 ( .A(n11387), .B(n11386), .ZN(n11389) );
  XNOR2_X1 U15911 ( .A(n11388), .B(n12409), .ZN(n11956) );
  XNOR2_X1 U15913 ( .A(n11717), .B(n12315), .ZN(n11941) );
  XNOR2_X1 U15914 ( .A(n11941), .B(n11614), .ZN(n11393) );
  XNOR2_X1 U15915 ( .A(n11661), .B(n20046), .ZN(n11390) );
  XNOR2_X1 U15916 ( .A(n11391), .B(n11390), .ZN(n11392) );
  XNOR2_X1 U15917 ( .A(n11393), .B(n11392), .ZN(n13023) );
  INV_X1 U15918 ( .A(n12494), .ZN(n11410) );
  XNOR2_X1 U15919 ( .A(n12334), .B(n12067), .ZN(n11394) );
  XNOR2_X1 U15920 ( .A(n11394), .B(n24970), .ZN(n11955) );
  XNOR2_X1 U15921 ( .A(n11795), .B(n16574), .ZN(n11395) );
  XNOR2_X1 U15922 ( .A(n12404), .B(n11395), .ZN(n11398) );
  XNOR2_X1 U15923 ( .A(n11396), .B(n11622), .ZN(n11397) );
  XNOR2_X1 U15924 ( .A(n11398), .B(n11397), .ZN(n11399) );
  XNOR2_X1 U15925 ( .A(n12343), .B(n12375), .ZN(n11604) );
  INV_X1 U15926 ( .A(n11401), .ZN(n12382) );
  XNOR2_X1 U15927 ( .A(n12382), .B(n25016), .ZN(n11402) );
  XNOR2_X1 U15928 ( .A(n11402), .B(n11604), .ZN(n11405) );
  XNOR2_X1 U15929 ( .A(n12344), .B(n12121), .ZN(n11931) );
  XNOR2_X1 U15930 ( .A(n11765), .B(n1757), .ZN(n11403) );
  XNOR2_X1 U15931 ( .A(n11931), .B(n11403), .ZN(n11404) );
  INV_X1 U15932 ( .A(n13028), .ZN(n13024) );
  INV_X1 U15933 ( .A(n13023), .ZN(n12758) );
  OAI21_X1 U15934 ( .B1(n13029), .B2(n13027), .A(n11406), .ZN(n11409) );
  NOR2_X1 U15935 ( .A1(n12784), .A2(n13030), .ZN(n11408) );
  INV_X1 U15936 ( .A(n11406), .ZN(n11407) );
  NOR2_X1 U15938 ( .A1(n13907), .A2(n11411), .ZN(n11453) );
  XNOR2_X1 U15939 ( .A(n12168), .B(n12089), .ZN(n11985) );
  XNOR2_X1 U15940 ( .A(n11985), .B(n11413), .ZN(n11418) );
  XNOR2_X1 U15941 ( .A(n11414), .B(n12362), .ZN(n11416) );
  XNOR2_X1 U15942 ( .A(n25371), .B(n2044), .ZN(n11415) );
  XNOR2_X1 U15943 ( .A(n11416), .B(n11415), .ZN(n11417) );
  XNOR2_X1 U15945 ( .A(n11951), .B(n12108), .ZN(n11419) );
  XNOR2_X1 U15946 ( .A(n11419), .B(n11420), .ZN(n11423) );
  XNOR2_X1 U15947 ( .A(n11689), .B(n2049), .ZN(n11421) );
  XNOR2_X1 U15948 ( .A(n11975), .B(n11421), .ZN(n11422) );
  XNOR2_X1 U15949 ( .A(n11423), .B(n11422), .ZN(n13056) );
  XNOR2_X1 U15951 ( .A(n11425), .B(n11942), .ZN(n11427) );
  XNOR2_X1 U15952 ( .A(n11427), .B(n11426), .ZN(n11430) );
  INV_X1 U15953 ( .A(n12082), .ZN(n11428) );
  XNOR2_X1 U15954 ( .A(n11429), .B(n11428), .ZN(n12013) );
  INV_X1 U15955 ( .A(n13057), .ZN(n13054) );
  XNOR2_X1 U15956 ( .A(n12383), .B(n21046), .ZN(n11431) );
  XNOR2_X1 U15957 ( .A(n11432), .B(n11431), .ZN(n11437) );
  XNOR2_X1 U15958 ( .A(n11433), .B(n11706), .ZN(n11434) );
  XNOR2_X1 U15959 ( .A(n11435), .B(n11434), .ZN(n11436) );
  XNOR2_X1 U15960 ( .A(n12005), .B(n11439), .ZN(n11444) );
  XNOR2_X1 U15961 ( .A(n11457), .B(n11440), .ZN(n11442) );
  INV_X1 U15962 ( .A(n12002), .ZN(n12075) );
  XNOR2_X1 U15963 ( .A(n12075), .B(n2208), .ZN(n11441) );
  XNOR2_X1 U15964 ( .A(n11442), .B(n11441), .ZN(n11443) );
  NOR2_X1 U15965 ( .A1(n303), .A2(n13056), .ZN(n12751) );
  XNOR2_X1 U15966 ( .A(n12147), .B(n11960), .ZN(n11445) );
  XNOR2_X1 U15967 ( .A(n11446), .B(n11445), .ZN(n11450) );
  XNOR2_X1 U15968 ( .A(n11741), .B(n12102), .ZN(n11448) );
  XNOR2_X1 U15969 ( .A(n11448), .B(n11447), .ZN(n11449) );
  XNOR2_X1 U15970 ( .A(n11450), .B(n11449), .ZN(n13052) );
  INV_X1 U15971 ( .A(n13052), .ZN(n13055) );
  AND2_X1 U15972 ( .A1(n13053), .A2(n13055), .ZN(n12485) );
  AOI21_X1 U15973 ( .B1(n12751), .B2(n25085), .A(n12485), .ZN(n11451) );
  NAND2_X1 U15974 ( .A1(n11452), .A2(n11451), .ZN(n14289) );
  INV_X1 U15975 ( .A(n12184), .ZN(n11455) );
  XNOR2_X1 U15976 ( .A(n11455), .B(n12129), .ZN(n11701) );
  XNOR2_X1 U15977 ( .A(n11701), .B(n11456), .ZN(n11461) );
  XNOR2_X1 U15978 ( .A(n11457), .B(n11637), .ZN(n11459) );
  XNOR2_X1 U15979 ( .A(n12356), .B(n912), .ZN(n11458) );
  XNOR2_X1 U15980 ( .A(n11459), .B(n11458), .ZN(n11460) );
  XNOR2_X1 U15981 ( .A(n11461), .B(n11460), .ZN(n12462) );
  INV_X1 U15982 ( .A(n12462), .ZN(n12713) );
  XNOR2_X1 U15985 ( .A(n11812), .B(n11463), .ZN(n11468) );
  XNOR2_X1 U15986 ( .A(n11464), .B(n12201), .ZN(n11466) );
  XNOR2_X1 U15987 ( .A(n24964), .B(n641), .ZN(n11465) );
  XNOR2_X1 U15988 ( .A(n11466), .B(n11465), .ZN(n11467) );
  XNOR2_X2 U15989 ( .A(n11468), .B(n11467), .ZN(n12483) );
  NOR2_X1 U15990 ( .A1(n12713), .A2(n12483), .ZN(n12464) );
  XNOR2_X1 U15991 ( .A(n11469), .B(n11816), .ZN(n11473) );
  XNOR2_X1 U15992 ( .A(n12404), .B(n12189), .ZN(n11471) );
  XNOR2_X1 U15993 ( .A(n11951), .B(n3178), .ZN(n11470) );
  XNOR2_X1 U15994 ( .A(n11471), .B(n11470), .ZN(n11472) );
  XNOR2_X1 U15995 ( .A(n11473), .B(n11472), .ZN(n12715) );
  INV_X1 U15996 ( .A(n12715), .ZN(n13078) );
  NOR2_X1 U15997 ( .A1(n12462), .A2(n13078), .ZN(n11474) );
  NOR2_X1 U15998 ( .A1(n12464), .A2(n11474), .ZN(n11589) );
  INV_X1 U15999 ( .A(n11960), .ZN(n11475) );
  XNOR2_X1 U16000 ( .A(n12144), .B(n11475), .ZN(n11476) );
  XNOR2_X1 U16001 ( .A(n11822), .B(n11476), .ZN(n11480) );
  XNOR2_X1 U16002 ( .A(n12414), .B(n12207), .ZN(n11478) );
  XNOR2_X1 U16003 ( .A(n25087), .B(n24287), .ZN(n11477) );
  XNOR2_X1 U16004 ( .A(n11478), .B(n11477), .ZN(n11479) );
  XNOR2_X1 U16006 ( .A(n11717), .B(n11660), .ZN(n11482) );
  XNOR2_X1 U16007 ( .A(n11482), .B(n11481), .ZN(n11485) );
  XNOR2_X1 U16008 ( .A(n11827), .B(n11483), .ZN(n11484) );
  XNOR2_X1 U16009 ( .A(n11485), .B(n11484), .ZN(n12707) );
  MUX2_X1 U16010 ( .A(n12710), .B(n12707), .S(n12483), .Z(n11592) );
  XNOR2_X1 U16011 ( .A(n25090), .B(n11486), .ZN(n11488) );
  XNOR2_X1 U16012 ( .A(n12370), .B(n3129), .ZN(n11487) );
  XNOR2_X1 U16013 ( .A(n11488), .B(n11487), .ZN(n11491) );
  XNOR2_X1 U16014 ( .A(n11489), .B(n11833), .ZN(n11490) );
  MUX2_X2 U16016 ( .A(n11589), .B(n11592), .S(n24573), .Z(n14362) );
  INV_X1 U16017 ( .A(n11492), .ZN(n11770) );
  XNOR2_X1 U16018 ( .A(n11770), .B(n12186), .ZN(n11493) );
  XNOR2_X1 U16019 ( .A(n11494), .B(n11493), .ZN(n11497) );
  XNOR2_X1 U16020 ( .A(n11627), .B(n836), .ZN(n11495) );
  XNOR2_X1 U16021 ( .A(n11856), .B(n11495), .ZN(n11496) );
  MUX2_X1 U16022 ( .A(n11500), .B(n11499), .S(n11498), .Z(n11503) );
  INV_X1 U16023 ( .A(n11501), .ZN(n11502) );
  NOR2_X1 U16024 ( .A1(n11503), .A2(n11502), .ZN(n11577) );
  XNOR2_X1 U16025 ( .A(n11619), .B(n11577), .ZN(n11505) );
  XNOR2_X1 U16026 ( .A(n12333), .B(n2735), .ZN(n11506) );
  XNOR2_X1 U16027 ( .A(n11868), .B(n11506), .ZN(n11507) );
  XNOR2_X1 U16028 ( .A(n11508), .B(n11507), .ZN(n12469) );
  NOR2_X1 U16029 ( .A1(n13067), .A2(n12469), .ZN(n11541) );
  XNOR2_X1 U16030 ( .A(n11915), .B(n11766), .ZN(n11509) );
  XNOR2_X1 U16031 ( .A(n11510), .B(n11509), .ZN(n11514) );
  XNOR2_X1 U16032 ( .A(n12200), .B(n1827), .ZN(n11511) );
  XNOR2_X1 U16033 ( .A(n11511), .B(n11512), .ZN(n11513) );
  INV_X1 U16034 ( .A(n11515), .ZN(n11517) );
  XNOR2_X1 U16035 ( .A(n24401), .B(n12040), .ZN(n11531) );
  NAND2_X1 U16036 ( .A1(n11520), .A2(n11524), .ZN(n11528) );
  INV_X1 U16037 ( .A(n11518), .ZN(n11521) );
  NAND3_X1 U16038 ( .A1(n11521), .A2(n11520), .A3(n11519), .ZN(n11523) );
  AND2_X1 U16039 ( .A1(n11522), .A2(n11523), .ZN(n11527) );
  NAND3_X1 U16040 ( .A1(n11525), .A2(n1332), .A3(n11524), .ZN(n11526) );
  XNOR2_X1 U16042 ( .A(n12323), .B(n3115), .ZN(n11530) );
  XNOR2_X1 U16043 ( .A(n11531), .B(n11530), .ZN(n11532) );
  INV_X1 U16044 ( .A(n12471), .ZN(n13072) );
  XNOR2_X1 U16045 ( .A(n12234), .B(n1724), .ZN(n11534) );
  XNOR2_X1 U16046 ( .A(n11535), .B(n11534), .ZN(n11540) );
  INV_X1 U16047 ( .A(n11536), .ZN(n11538) );
  XNOR2_X1 U16048 ( .A(n11538), .B(n11537), .ZN(n11539) );
  XNOR2_X1 U16049 ( .A(n11542), .B(n12313), .ZN(n11544) );
  XNOR2_X1 U16050 ( .A(n11544), .B(n11543), .ZN(n11547) );
  XNOR2_X1 U16051 ( .A(n11863), .B(n11545), .ZN(n11546) );
  INV_X1 U16052 ( .A(n12773), .ZN(n13071) );
  NOR2_X1 U16053 ( .A1(n13071), .A2(n12471), .ZN(n11548) );
  NOR3_X1 U16054 ( .A1(n11549), .A2(n13070), .A3(n11548), .ZN(n11550) );
  NOR2_X2 U16055 ( .A1(n11551), .A2(n11550), .ZN(n14361) );
  NAND2_X1 U16056 ( .A1(n14362), .A2(n14361), .ZN(n13711) );
  XNOR2_X1 U16057 ( .A(n11715), .B(n11659), .ZN(n12259) );
  XNOR2_X1 U16058 ( .A(n11789), .B(n12259), .ZN(n11554) );
  XNOR2_X1 U16059 ( .A(n12225), .B(n2215), .ZN(n11552) );
  XNOR2_X1 U16060 ( .A(n12011), .B(n11552), .ZN(n11553) );
  XNOR2_X1 U16061 ( .A(n11554), .B(n11553), .ZN(n13038) );
  INV_X1 U16062 ( .A(n13038), .ZN(n12476) );
  XNOR2_X1 U16063 ( .A(n11555), .B(n12214), .ZN(n11557) );
  XNOR2_X1 U16064 ( .A(n24027), .B(n11653), .ZN(n12284) );
  XNOR2_X1 U16065 ( .A(n11557), .B(n12284), .ZN(n11560) );
  XNOR2_X1 U16066 ( .A(n12040), .B(n869), .ZN(n11558) );
  XNOR2_X1 U16067 ( .A(n11781), .B(n11558), .ZN(n11559) );
  XNOR2_X1 U16068 ( .A(n11560), .B(n11559), .ZN(n13037) );
  INV_X1 U16069 ( .A(n13037), .ZN(n12798) );
  XNOR2_X1 U16072 ( .A(n11563), .B(n12365), .ZN(n12166) );
  XNOR2_X1 U16073 ( .A(n12246), .B(n12166), .ZN(n11567) );
  XNOR2_X1 U16074 ( .A(n11564), .B(n11983), .ZN(n12230) );
  XNOR2_X1 U16075 ( .A(n11908), .B(n887), .ZN(n11565) );
  XNOR2_X1 U16076 ( .A(n12230), .B(n11565), .ZN(n11566) );
  XNOR2_X1 U16077 ( .A(n11879), .B(n12186), .ZN(n11569) );
  XNOR2_X1 U16078 ( .A(n11568), .B(n11640), .ZN(n12268) );
  XNOR2_X1 U16079 ( .A(n11569), .B(n12268), .ZN(n11573) );
  XNOR2_X1 U16080 ( .A(n11570), .B(n11571), .ZN(n11572) );
  XNOR2_X1 U16081 ( .A(n12277), .B(n12396), .ZN(n11792) );
  XNOR2_X1 U16082 ( .A(n11792), .B(n25236), .ZN(n11575) );
  XNOR2_X1 U16083 ( .A(n11672), .B(n11689), .ZN(n12273) );
  XNOR2_X1 U16084 ( .A(n11575), .B(n12273), .ZN(n11579) );
  XNOR2_X1 U16085 ( .A(n11977), .B(n3152), .ZN(n11576) );
  XNOR2_X1 U16086 ( .A(n11577), .B(n11576), .ZN(n11578) );
  XNOR2_X1 U16087 ( .A(n11579), .B(n11578), .ZN(n12800) );
  XNOR2_X1 U16088 ( .A(n12239), .B(n11800), .ZN(n11586) );
  XNOR2_X1 U16089 ( .A(n11581), .B(n11582), .ZN(n11584) );
  XNOR2_X1 U16090 ( .A(n12196), .B(n1874), .ZN(n11583) );
  XNOR2_X1 U16091 ( .A(n11584), .B(n11583), .ZN(n11585) );
  XNOR2_X1 U16092 ( .A(n11586), .B(n11585), .ZN(n12519) );
  INV_X1 U16093 ( .A(n12519), .ZN(n13039) );
  NOR2_X1 U16094 ( .A1(n13039), .A2(n13038), .ZN(n11588) );
  INV_X1 U16095 ( .A(n13041), .ZN(n11587) );
  OAI21_X1 U16096 ( .B1(n11588), .B2(n13044), .A(n11587), .ZN(n11590) );
  INV_X1 U16097 ( .A(n11590), .ZN(n11591) );
  AOI21_X1 U16098 ( .B1(n11592), .B2(n24573), .A(n11591), .ZN(n11593) );
  NAND2_X1 U16099 ( .A1(n11594), .A2(n11593), .ZN(n11601) );
  INV_X1 U16100 ( .A(n11595), .ZN(n11600) );
  INV_X1 U16101 ( .A(n13169), .ZN(n12718) );
  OAI22_X1 U16102 ( .A1(n12716), .A2(n11597), .B1(n12719), .B2(n10502), .ZN(
        n11598) );
  XNOR2_X1 U16103 ( .A(n11914), .B(n1810), .ZN(n11603) );
  XNOR2_X1 U16104 ( .A(n11602), .B(n11603), .ZN(n11606) );
  XNOR2_X1 U16105 ( .A(n11704), .B(n11766), .ZN(n12342) );
  XNOR2_X1 U16106 ( .A(n12342), .B(n11604), .ZN(n11605) );
  XNOR2_X1 U16107 ( .A(n11736), .B(n11607), .ZN(n12292) );
  XNOR2_X1 U16108 ( .A(n11608), .B(n12292), .ZN(n11612) );
  XNOR2_X1 U16109 ( .A(n12249), .B(n22986), .ZN(n11609) );
  XNOR2_X1 U16110 ( .A(n11610), .B(n11609), .ZN(n11611) );
  XNOR2_X1 U16112 ( .A(n12388), .B(n2318), .ZN(n11613) );
  XNOR2_X1 U16113 ( .A(n11613), .B(n12255), .ZN(n11615) );
  XNOR2_X1 U16114 ( .A(n11749), .B(n11616), .ZN(n12312) );
  XNOR2_X1 U16115 ( .A(n12312), .B(n24915), .ZN(n11617) );
  XNOR2_X1 U16116 ( .A(n11618), .B(n11619), .ZN(n12339) );
  XNOR2_X1 U16117 ( .A(n12112), .B(n3131), .ZN(n11620) );
  XNOR2_X1 U16118 ( .A(n11620), .B(n12397), .ZN(n11621) );
  XNOR2_X1 U16119 ( .A(n11621), .B(n12339), .ZN(n11625) );
  XNOR2_X1 U16120 ( .A(n11622), .B(n12275), .ZN(n11623) );
  XNOR2_X1 U16121 ( .A(n12404), .B(n11623), .ZN(n11624) );
  XNOR2_X1 U16122 ( .A(n11699), .B(n11626), .ZN(n11631) );
  XNOR2_X1 U16123 ( .A(n11698), .B(n11627), .ZN(n12307) );
  XNOR2_X1 U16124 ( .A(n11628), .B(n11809), .ZN(n11629) );
  XNOR2_X1 U16125 ( .A(n12307), .B(n11629), .ZN(n11630) );
  XNOR2_X1 U16127 ( .A(n12283), .B(n12324), .ZN(n11632) );
  XNOR2_X1 U16128 ( .A(n11632), .B(n12320), .ZN(n11636) );
  XNOR2_X1 U16129 ( .A(n11897), .B(n12413), .ZN(n11634) );
  XNOR2_X1 U16130 ( .A(n12414), .B(n92), .ZN(n11633) );
  XNOR2_X1 U16131 ( .A(n11634), .B(n11633), .ZN(n11635) );
  XNOR2_X1 U16132 ( .A(n12132), .B(n11639), .ZN(n11644) );
  XNOR2_X1 U16133 ( .A(n11640), .B(n1924), .ZN(n11641) );
  XNOR2_X1 U16134 ( .A(n11642), .B(n11641), .ZN(n11643) );
  XNOR2_X1 U16135 ( .A(n25090), .B(n11735), .ZN(n12165) );
  XNOR2_X1 U16136 ( .A(n11734), .B(n12165), .ZN(n11650) );
  XNOR2_X1 U16137 ( .A(n11646), .B(n2477), .ZN(n11647) );
  XNOR2_X1 U16138 ( .A(n11648), .B(n11647), .ZN(n11649) );
  INV_X1 U16139 ( .A(Key[172]), .ZN(n23271) );
  XNOR2_X1 U16140 ( .A(n12325), .B(n23271), .ZN(n11651) );
  XNOR2_X1 U16141 ( .A(n11651), .B(n12146), .ZN(n11652) );
  XNOR2_X1 U16142 ( .A(n12409), .B(n12102), .ZN(n11743) );
  XNOR2_X1 U16143 ( .A(n11652), .B(n11743), .ZN(n11656) );
  XNOR2_X1 U16144 ( .A(n25087), .B(n11653), .ZN(n11654) );
  XNOR2_X1 U16145 ( .A(n12152), .B(n11654), .ZN(n11655) );
  XNOR2_X1 U16148 ( .A(n12053), .B(n2747), .ZN(n11657) );
  XNOR2_X1 U16149 ( .A(n11658), .B(n11657), .ZN(n11664) );
  XNOR2_X1 U16150 ( .A(n11659), .B(n12082), .ZN(n11662) );
  XNOR2_X1 U16151 ( .A(n11661), .B(n11660), .ZN(n12157) );
  XNOR2_X1 U16152 ( .A(n12157), .B(n11662), .ZN(n11663) );
  XNOR2_X1 U16153 ( .A(n11666), .B(n11665), .ZN(n11669) );
  XNOR2_X1 U16154 ( .A(n11765), .B(n11464), .ZN(n11798) );
  XNOR2_X1 U16155 ( .A(n11838), .B(n1815), .ZN(n11667) );
  XNOR2_X1 U16156 ( .A(n11798), .B(n11667), .ZN(n11668) );
  XNOR2_X1 U16157 ( .A(n11668), .B(n11669), .ZN(n12454) );
  NOR2_X1 U16158 ( .A1(n13063), .A2(n13061), .ZN(n11678) );
  XNOR2_X1 U16159 ( .A(n11795), .B(n1854), .ZN(n11670) );
  XNOR2_X1 U16160 ( .A(n11670), .B(n12334), .ZN(n11671) );
  XNOR2_X1 U16161 ( .A(n12108), .B(n12402), .ZN(n11758) );
  XNOR2_X1 U16162 ( .A(n11671), .B(n11758), .ZN(n11676) );
  INV_X1 U16163 ( .A(n11672), .ZN(n11673) );
  XNOR2_X1 U16164 ( .A(n11673), .B(n25236), .ZN(n11674) );
  XNOR2_X1 U16165 ( .A(n11796), .B(n11674), .ZN(n11675) );
  XNOR2_X1 U16166 ( .A(n11676), .B(n11675), .ZN(n12439) );
  INV_X1 U16167 ( .A(n12439), .ZN(n13163) );
  NAND2_X1 U16168 ( .A1(n13163), .A2(n1353), .ZN(n11677) );
  NAND2_X1 U16169 ( .A1(n13394), .A2(n13568), .ZN(n11679) );
  OR2_X1 U16170 ( .A1(n13712), .A2(n11679), .ZN(n11680) );
  XNOR2_X1 U16171 ( .A(n11682), .B(n15401), .ZN(n14884) );
  NAND2_X1 U16172 ( .A1(n13211), .A2(n11684), .ZN(n12551) );
  NAND3_X1 U16173 ( .A1(n13213), .A2(n11684), .A3(n13004), .ZN(n11683) );
  OAI21_X1 U16174 ( .B1(n12551), .B2(n11360), .A(n11683), .ZN(n11685) );
  INV_X1 U16175 ( .A(n13000), .ZN(n13212) );
  XNOR2_X1 U16176 ( .A(n11686), .B(n23699), .ZN(n11687) );
  XNOR2_X1 U16177 ( .A(n11687), .B(n24969), .ZN(n11688) );
  XNOR2_X1 U16178 ( .A(n12064), .B(n11688), .ZN(n11691) );
  XNOR2_X1 U16179 ( .A(n11689), .B(n11690), .ZN(n11926) );
  XNOR2_X1 U16180 ( .A(n11691), .B(n11926), .ZN(n12613) );
  INV_X1 U16181 ( .A(n11692), .ZN(n11906) );
  XNOR2_X1 U16182 ( .A(n11906), .B(n12030), .ZN(n11697) );
  INV_X1 U16183 ( .A(n11693), .ZN(n11695) );
  XNOR2_X1 U16184 ( .A(n12167), .B(n21742), .ZN(n11694) );
  XNOR2_X1 U16185 ( .A(n11695), .B(n11694), .ZN(n11696) );
  NAND2_X1 U16187 ( .A1(n12613), .A2(n13305), .ZN(n12558) );
  XNOR2_X1 U16188 ( .A(n11698), .B(n5286), .ZN(n11700) );
  INV_X1 U16189 ( .A(n11701), .ZN(n11702) );
  XNOR2_X1 U16190 ( .A(n11703), .B(n12201), .ZN(n12045) );
  XNOR2_X1 U16191 ( .A(n11704), .B(n925), .ZN(n11705) );
  XNOR2_X1 U16192 ( .A(n12096), .B(n12200), .ZN(n11707) );
  XNOR2_X1 U16193 ( .A(n11706), .B(n11707), .ZN(n11918) );
  XNOR2_X1 U16194 ( .A(n11708), .B(n11918), .ZN(n12611) );
  XNOR2_X1 U16196 ( .A(n11959), .B(n2744), .ZN(n11709) );
  XNOR2_X1 U16197 ( .A(n25418), .B(n11709), .ZN(n11713) );
  XNOR2_X1 U16198 ( .A(n11897), .B(n12144), .ZN(n11711) );
  XNOR2_X1 U16199 ( .A(n11711), .B(n11900), .ZN(n11712) );
  OAI21_X1 U16200 ( .B1(n12558), .B2(n12915), .A(n11714), .ZN(n11723) );
  XNOR2_X1 U16201 ( .A(n11715), .B(n12224), .ZN(n11890) );
  XNOR2_X1 U16202 ( .A(n11716), .B(n11890), .ZN(n11721) );
  XNOR2_X1 U16203 ( .A(n11717), .B(n1856), .ZN(n11719) );
  INV_X1 U16204 ( .A(n11718), .ZN(n12058) );
  XNOR2_X1 U16205 ( .A(n11719), .B(n12058), .ZN(n11720) );
  INV_X1 U16206 ( .A(n11724), .ZN(n11726) );
  XNOR2_X1 U16207 ( .A(n11725), .B(n11726), .ZN(n11731) );
  XNOR2_X1 U16208 ( .A(n11771), .B(n11966), .ZN(n11729) );
  INV_X1 U16209 ( .A(n12351), .ZN(n11727) );
  XNOR2_X1 U16210 ( .A(n11727), .B(n768), .ZN(n11728) );
  XNOR2_X1 U16211 ( .A(n11729), .B(n11728), .ZN(n11730) );
  XNOR2_X1 U16213 ( .A(n12362), .B(n24514), .ZN(n11733) );
  XNOR2_X1 U16214 ( .A(n11734), .B(n11733), .ZN(n11740) );
  INV_X1 U16215 ( .A(n21169), .ZN(n22556) );
  XNOR2_X1 U16216 ( .A(n11735), .B(n22556), .ZN(n11738) );
  XNOR2_X1 U16217 ( .A(n11736), .B(n25371), .ZN(n11737) );
  XNOR2_X1 U16218 ( .A(n11738), .B(n11737), .ZN(n11739) );
  XNOR2_X1 U16219 ( .A(n11741), .B(n11960), .ZN(n12416) );
  XNOR2_X1 U16220 ( .A(n12286), .B(n2040), .ZN(n11742) );
  XNOR2_X1 U16221 ( .A(n12416), .B(n11742), .ZN(n11744) );
  INV_X1 U16222 ( .A(n13227), .ZN(n11754) );
  XNOR2_X1 U16223 ( .A(n12053), .B(n11746), .ZN(n11748) );
  XNOR2_X1 U16224 ( .A(n11747), .B(n11748), .ZN(n12395) );
  XNOR2_X1 U16225 ( .A(n11749), .B(n2847), .ZN(n11750) );
  XNOR2_X1 U16226 ( .A(n12257), .B(n12082), .ZN(n11751) );
  XNOR2_X1 U16227 ( .A(n11752), .B(n11751), .ZN(n11753) );
  NOR2_X1 U16228 ( .A1(n13221), .A2(n11755), .ZN(n12920) );
  XNOR2_X1 U16229 ( .A(n11756), .B(n11951), .ZN(n12400) );
  XNOR2_X1 U16230 ( .A(n12277), .B(n23620), .ZN(n11757) );
  XNOR2_X1 U16231 ( .A(n11759), .B(n11758), .ZN(n11760) );
  XNOR2_X1 U16232 ( .A(n11761), .B(n923), .ZN(n11762) );
  XNOR2_X1 U16233 ( .A(n12376), .B(n11762), .ZN(n11763) );
  XNOR2_X1 U16234 ( .A(n11765), .B(n24964), .ZN(n11767) );
  XNOR2_X1 U16235 ( .A(n11767), .B(n11766), .ZN(n11768) );
  INV_X1 U16236 ( .A(n12569), .ZN(n12924) );
  OAI211_X1 U16237 ( .C1(n13223), .C2(n12885), .A(n12924), .B(n13224), .ZN(
        n11769) );
  OAI21_X1 U16238 ( .B1(n13010), .B2(n12920), .A(n11769), .ZN(n13965) );
  XNOR2_X1 U16239 ( .A(n12132), .B(n12074), .ZN(n11775) );
  XNOR2_X1 U16240 ( .A(n11771), .B(n11770), .ZN(n11773) );
  XNOR2_X1 U16241 ( .A(n12355), .B(n1758), .ZN(n11772) );
  XNOR2_X1 U16242 ( .A(n11773), .B(n11772), .ZN(n11774) );
  XNOR2_X1 U16243 ( .A(n12165), .B(n12088), .ZN(n11780) );
  XNOR2_X1 U16244 ( .A(n12296), .B(n12365), .ZN(n11778) );
  XNOR2_X1 U16245 ( .A(n11908), .B(n763), .ZN(n11777) );
  XNOR2_X1 U16246 ( .A(n11778), .B(n11777), .ZN(n11779) );
  INV_X1 U16247 ( .A(n12594), .ZN(n12597) );
  XNOR2_X1 U16248 ( .A(n24980), .B(n12323), .ZN(n11784) );
  XNOR2_X1 U16249 ( .A(n25087), .B(n62), .ZN(n11783) );
  XNOR2_X1 U16250 ( .A(n11784), .B(n11783), .ZN(n11785) );
  XNOR2_X1 U16252 ( .A(n12157), .B(n11787), .ZN(n11791) );
  XNOR2_X1 U16253 ( .A(n12313), .B(n2190), .ZN(n11788) );
  XNOR2_X1 U16254 ( .A(n11789), .B(n11788), .ZN(n11790) );
  XNOR2_X1 U16255 ( .A(n11790), .B(n11791), .ZN(n13288) );
  XNOR2_X1 U16257 ( .A(n12333), .B(n1777), .ZN(n11793) );
  XNOR2_X1 U16258 ( .A(n11792), .B(n11793), .ZN(n11794) );
  XNOR2_X1 U16260 ( .A(n11796), .B(n11795), .ZN(n12141) );
  XNOR2_X1 U16261 ( .A(n12095), .B(n11800), .ZN(n11801) );
  XNOR2_X1 U16262 ( .A(n11802), .B(n11801), .ZN(n12593) );
  BUF_X2 U16263 ( .A(n12593), .Z(n12827) );
  NOR2_X1 U16264 ( .A1(n11804), .A2(n11803), .ZN(n11805) );
  INV_X1 U16265 ( .A(n11805), .ZN(n13884) );
  XNOR2_X1 U16267 ( .A(n12019), .B(n12002), .ZN(n11808) );
  XNOR2_X1 U16268 ( .A(n12357), .B(n1855), .ZN(n11807) );
  XNOR2_X1 U16269 ( .A(n11808), .B(n11807), .ZN(n11811) );
  XNOR2_X1 U16270 ( .A(n12186), .B(n11809), .ZN(n12025) );
  XNOR2_X1 U16271 ( .A(n12306), .B(n12129), .ZN(n11970) );
  XNOR2_X1 U16272 ( .A(n12025), .B(n11970), .ZN(n11810) );
  XNOR2_X1 U16273 ( .A(n11812), .B(n12046), .ZN(n11815) );
  XNOR2_X1 U16274 ( .A(n11931), .B(n11813), .ZN(n11814) );
  XNOR2_X1 U16276 ( .A(n12334), .B(n12138), .ZN(n11817) );
  XNOR2_X1 U16277 ( .A(n11816), .B(n11817), .ZN(n11820) );
  XNOR2_X1 U16278 ( .A(n12108), .B(n23679), .ZN(n11818) );
  XNOR2_X1 U16279 ( .A(n12063), .B(n11818), .ZN(n11819) );
  XNOR2_X1 U16280 ( .A(n12144), .B(n12324), .ZN(n11821) );
  XNOR2_X1 U16281 ( .A(n11822), .B(n11821), .ZN(n11826) );
  XNOR2_X1 U16282 ( .A(n12040), .B(n12102), .ZN(n11824) );
  XNOR2_X1 U16283 ( .A(n12325), .B(n1746), .ZN(n11823) );
  XNOR2_X1 U16284 ( .A(n11824), .B(n11823), .ZN(n11825) );
  XNOR2_X1 U16285 ( .A(n11826), .B(n11825), .ZN(n12935) );
  XNOR2_X1 U16287 ( .A(n12082), .B(n20744), .ZN(n11828) );
  XNOR2_X1 U16288 ( .A(n11827), .B(n11828), .ZN(n11831) );
  INV_X1 U16289 ( .A(n11829), .ZN(n12057) );
  XNOR2_X1 U16290 ( .A(n11941), .B(n12057), .ZN(n11830) );
  INV_X1 U16291 ( .A(n13298), .ZN(n12936) );
  XNOR2_X1 U16292 ( .A(n12089), .B(n1875), .ZN(n11832) );
  XNOR2_X1 U16293 ( .A(n11832), .B(n11946), .ZN(n11835) );
  XNOR2_X1 U16294 ( .A(n11833), .B(n12028), .ZN(n11834) );
  XNOR2_X1 U16295 ( .A(n12377), .B(n25016), .ZN(n11841) );
  XNOR2_X1 U16296 ( .A(n11842), .B(n11841), .ZN(n11843) );
  XNOR2_X1 U16298 ( .A(n12413), .B(n11845), .ZN(n11847) );
  XNOR2_X1 U16299 ( .A(n12323), .B(n2970), .ZN(n11846) );
  INV_X1 U16300 ( .A(n11848), .ZN(n12105) );
  XNOR2_X1 U16301 ( .A(n11849), .B(n12105), .ZN(n11850) );
  XNOR2_X1 U16302 ( .A(n25234), .B(n1870), .ZN(n11853) );
  INV_X1 U16303 ( .A(n11851), .ZN(n11852) );
  XNOR2_X1 U16304 ( .A(n11852), .B(n11853), .ZN(n11855) );
  XNOR2_X1 U16305 ( .A(n12087), .B(n11905), .ZN(n11854) );
  XNOR2_X1 U16308 ( .A(n12073), .B(n11856), .ZN(n11860) );
  XNOR2_X1 U16309 ( .A(n12020), .B(n921), .ZN(n11857) );
  XNOR2_X1 U16310 ( .A(n11858), .B(n11857), .ZN(n11859) );
  INV_X1 U16311 ( .A(n11861), .ZN(n12080) );
  XNOR2_X1 U16312 ( .A(n12388), .B(n2036), .ZN(n11862) );
  XNOR2_X1 U16313 ( .A(n12080), .B(n11862), .ZN(n11865) );
  XNOR2_X1 U16314 ( .A(n11863), .B(n11893), .ZN(n11864) );
  XNOR2_X1 U16315 ( .A(n11865), .B(n11864), .ZN(n12900) );
  NAND2_X1 U16316 ( .A1(n12899), .A2(n12900), .ZN(n11866) );
  NAND3_X1 U16317 ( .A1(n11867), .A2(n5672), .A3(n11866), .ZN(n11875) );
  XNOR2_X1 U16318 ( .A(n11924), .B(n12110), .ZN(n11872) );
  XNOR2_X1 U16319 ( .A(n12397), .B(n1864), .ZN(n11870) );
  INV_X1 U16320 ( .A(n11868), .ZN(n11869) );
  XNOR2_X1 U16321 ( .A(n11870), .B(n11869), .ZN(n11871) );
  NAND3_X1 U16322 ( .A1(n12928), .A2(n12897), .A3(n11873), .ZN(n11874) );
  XNOR2_X1 U16323 ( .A(n12183), .B(n2717), .ZN(n11877) );
  XNOR2_X1 U16324 ( .A(n11878), .B(n11877), .ZN(n11883) );
  XNOR2_X1 U16325 ( .A(n11879), .B(n12019), .ZN(n11881) );
  XNOR2_X1 U16326 ( .A(n11881), .B(n11880), .ZN(n11882) );
  NAND2_X1 U16327 ( .A1(n714), .A2(n11884), .ZN(n11887) );
  NAND2_X1 U16328 ( .A1(n10690), .A2(n11147), .ZN(n11886) );
  MUX2_X1 U16329 ( .A(n11887), .B(n11886), .S(n11885), .Z(n11889) );
  NAND2_X1 U16330 ( .A1(n11889), .A2(n11888), .ZN(n12055) );
  XNOR2_X1 U16331 ( .A(n12055), .B(n12226), .ZN(n11891) );
  XNOR2_X1 U16332 ( .A(n11891), .B(n11890), .ZN(n11896) );
  XNOR2_X1 U16333 ( .A(n11892), .B(n889), .ZN(n11894) );
  XNOR2_X1 U16334 ( .A(n11894), .B(n11893), .ZN(n11895) );
  XNOR2_X1 U16335 ( .A(n11895), .B(n11896), .ZN(n12942) );
  INV_X1 U16336 ( .A(n12101), .ZN(n11898) );
  XNOR2_X1 U16337 ( .A(n12283), .B(n11898), .ZN(n11899) );
  XNOR2_X1 U16338 ( .A(n11899), .B(n11900), .ZN(n11904) );
  XNOR2_X1 U16339 ( .A(n12039), .B(n12286), .ZN(n11902) );
  XNOR2_X1 U16340 ( .A(n12323), .B(n4189), .ZN(n11901) );
  XNOR2_X1 U16341 ( .A(n11902), .B(n11901), .ZN(n11903) );
  INV_X1 U16342 ( .A(n12031), .ZN(n11909) );
  XNOR2_X1 U16343 ( .A(n11909), .B(n22745), .ZN(n11910) );
  XNOR2_X1 U16344 ( .A(n11911), .B(n11910), .ZN(n11912) );
  XNOR2_X2 U16345 ( .A(n5749), .B(n11912), .ZN(n13317) );
  NOR2_X1 U16346 ( .A1(n12945), .A2(n13317), .ZN(n11920) );
  XNOR2_X1 U16347 ( .A(n11916), .B(n11915), .ZN(n11917) );
  MUX2_X1 U16348 ( .A(n11921), .B(n11920), .S(n25499), .Z(n11928) );
  XNOR2_X1 U16349 ( .A(n12277), .B(n23883), .ZN(n11923) );
  INV_X1 U16350 ( .A(n12066), .ZN(n11922) );
  INV_X1 U16352 ( .A(n13318), .ZN(n12580) );
  INV_X1 U16353 ( .A(n12942), .ZN(n13316) );
  OAI22_X1 U16354 ( .A1(n13321), .A2(n12580), .B1(n12687), .B2(n13316), .ZN(
        n11927) );
  XNOR2_X1 U16355 ( .A(n12382), .B(n12241), .ZN(n11930) );
  XNOR2_X1 U16356 ( .A(n24964), .B(n2826), .ZN(n11929) );
  XNOR2_X1 U16357 ( .A(n11930), .B(n11929), .ZN(n11933) );
  XNOR2_X1 U16358 ( .A(n12342), .B(n11931), .ZN(n11932) );
  XNOR2_X1 U16359 ( .A(n11932), .B(n11933), .ZN(n12600) );
  NAND2_X1 U16360 ( .A1(n11935), .A2(n4711), .ZN(n11938) );
  NAND2_X1 U16361 ( .A1(n11939), .A2(n11934), .ZN(n11937) );
  MUX2_X1 U16362 ( .A(n4711), .B(n1495), .S(n11935), .Z(n11936) );
  OAI211_X1 U16363 ( .C1(n11939), .C2(n11938), .A(n11937), .B(n11936), .ZN(
        n11940) );
  XNOR2_X1 U16364 ( .A(n11941), .B(n11940), .ZN(n11945) );
  XNOR2_X1 U16365 ( .A(n12053), .B(n11942), .ZN(n11944) );
  INV_X1 U16366 ( .A(n12312), .ZN(n11943) );
  NOR2_X1 U16367 ( .A1(n12966), .A2(n12963), .ZN(n11974) );
  XNOR2_X1 U16368 ( .A(n12292), .B(n11946), .ZN(n11950) );
  XNOR2_X1 U16369 ( .A(n12364), .B(n25371), .ZN(n11948) );
  XNOR2_X1 U16370 ( .A(n12168), .B(n2039), .ZN(n11947) );
  XNOR2_X1 U16371 ( .A(n11948), .B(n11947), .ZN(n11949) );
  XNOR2_X1 U16372 ( .A(n11950), .B(n11949), .ZN(n11965) );
  XNOR2_X1 U16373 ( .A(n12276), .B(n2058), .ZN(n11952) );
  XNOR2_X1 U16374 ( .A(n11952), .B(n11951), .ZN(n11953) );
  XNOR2_X1 U16375 ( .A(n11953), .B(n12339), .ZN(n11954) );
  XNOR2_X1 U16376 ( .A(n11954), .B(n11955), .ZN(n13275) );
  INV_X1 U16377 ( .A(n11956), .ZN(n11964) );
  XNOR2_X1 U16378 ( .A(n11957), .B(n896), .ZN(n11958) );
  XNOR2_X1 U16379 ( .A(n12282), .B(n11958), .ZN(n11962) );
  XNOR2_X1 U16380 ( .A(n11960), .B(n11959), .ZN(n11961) );
  XNOR2_X1 U16381 ( .A(n11962), .B(n11961), .ZN(n11963) );
  XNOR2_X1 U16382 ( .A(n11966), .B(n12130), .ZN(n11969) );
  INV_X1 U16383 ( .A(n11967), .ZN(n12352) );
  XNOR2_X1 U16384 ( .A(n12352), .B(n2193), .ZN(n11968) );
  XNOR2_X1 U16385 ( .A(n11969), .B(n11968), .ZN(n11973) );
  INV_X1 U16386 ( .A(n11970), .ZN(n11971) );
  XNOR2_X1 U16387 ( .A(n12307), .B(n11971), .ZN(n11972) );
  NOR2_X1 U16388 ( .A1(n24588), .A2(n13945), .ZN(n13890) );
  XNOR2_X1 U16389 ( .A(n12401), .B(n2236), .ZN(n11976) );
  XNOR2_X1 U16390 ( .A(n11975), .B(n11976), .ZN(n11980) );
  INV_X1 U16391 ( .A(n12108), .ZN(n11978) );
  XNOR2_X1 U16392 ( .A(n11977), .B(n11978), .ZN(n11979) );
  XNOR2_X1 U16393 ( .A(n12363), .B(n11983), .ZN(n11984) );
  XNOR2_X1 U16394 ( .A(n11985), .B(n11984), .ZN(n11989) );
  XNOR2_X1 U16395 ( .A(n12362), .B(n876), .ZN(n11987) );
  XNOR2_X1 U16396 ( .A(n11986), .B(n11987), .ZN(n11988) );
  XNOR2_X1 U16398 ( .A(n12102), .B(n2772), .ZN(n11990) );
  XNOR2_X1 U16399 ( .A(n11992), .B(n12410), .ZN(n11993) );
  XNOR2_X1 U16400 ( .A(n11994), .B(n11993), .ZN(n12680) );
  INV_X1 U16401 ( .A(n11995), .ZN(n11997) );
  XNOR2_X1 U16402 ( .A(n11997), .B(n11996), .ZN(n12001) );
  XNOR2_X1 U16403 ( .A(n12196), .B(n2726), .ZN(n11998) );
  XNOR2_X1 U16404 ( .A(n11999), .B(n11998), .ZN(n12000) );
  XNOR2_X1 U16405 ( .A(n12002), .B(n25396), .ZN(n12004) );
  XNOR2_X1 U16406 ( .A(n12005), .B(n12004), .ZN(n12009) );
  XNOR2_X1 U16407 ( .A(n12357), .B(n187), .ZN(n12007) );
  XNOR2_X1 U16408 ( .A(n12356), .B(n12127), .ZN(n12006) );
  XNOR2_X1 U16409 ( .A(n12006), .B(n12007), .ZN(n12008) );
  XNOR2_X1 U16410 ( .A(n12008), .B(n12009), .ZN(n12934) );
  XNOR2_X1 U16411 ( .A(n12010), .B(n12389), .ZN(n12012) );
  XNOR2_X1 U16412 ( .A(n12012), .B(n12011), .ZN(n12015) );
  INV_X1 U16413 ( .A(n12013), .ZN(n12014) );
  NAND2_X1 U16414 ( .A1(n25015), .A2(n13264), .ZN(n12016) );
  AOI21_X1 U16415 ( .B1(n12829), .B2(n12016), .A(n13265), .ZN(n12017) );
  NOR2_X1 U16416 ( .A1(n13890), .A2(n12018), .ZN(n12177) );
  INV_X1 U16417 ( .A(n12019), .ZN(n12022) );
  XNOR2_X1 U16418 ( .A(n12020), .B(n12352), .ZN(n12021) );
  XNOR2_X1 U16419 ( .A(n12022), .B(n12021), .ZN(n12027) );
  XNOR2_X1 U16420 ( .A(n12023), .B(n1726), .ZN(n12024) );
  XNOR2_X1 U16421 ( .A(n12029), .B(n12030), .ZN(n12035) );
  XNOR2_X1 U16422 ( .A(n12031), .B(n12364), .ZN(n12033) );
  XNOR2_X1 U16423 ( .A(n12234), .B(n1804), .ZN(n12032) );
  XNOR2_X1 U16424 ( .A(n12033), .B(n12032), .ZN(n12034) );
  INV_X1 U16425 ( .A(n12324), .ZN(n12036) );
  XNOR2_X1 U16426 ( .A(n12036), .B(n12409), .ZN(n12037) );
  XNOR2_X1 U16427 ( .A(n12038), .B(n12037), .ZN(n12044) );
  XNOR2_X1 U16428 ( .A(n12039), .B(n12212), .ZN(n12042) );
  XNOR2_X1 U16429 ( .A(n12040), .B(n891), .ZN(n12041) );
  XNOR2_X1 U16430 ( .A(n12042), .B(n12041), .ZN(n12043) );
  INV_X1 U16431 ( .A(n12045), .ZN(n12047) );
  XNOR2_X1 U16432 ( .A(n12047), .B(n12046), .ZN(n12052) );
  XNOR2_X1 U16433 ( .A(n12382), .B(n12197), .ZN(n12050) );
  XNOR2_X1 U16434 ( .A(n12048), .B(n1768), .ZN(n12049) );
  XNOR2_X1 U16435 ( .A(n12050), .B(n12049), .ZN(n12051) );
  XNOR2_X1 U16436 ( .A(n12052), .B(n12051), .ZN(n13328) );
  NAND2_X1 U16437 ( .A1(n12684), .A2(n24422), .ZN(n12062) );
  INV_X1 U16438 ( .A(n12053), .ZN(n12054) );
  XNOR2_X1 U16439 ( .A(n12055), .B(n12054), .ZN(n12056) );
  XNOR2_X1 U16440 ( .A(n12056), .B(n12057), .ZN(n12061) );
  XNOR2_X1 U16441 ( .A(n12221), .B(n21703), .ZN(n12059) );
  XNOR2_X1 U16442 ( .A(n12058), .B(n12059), .ZN(n12060) );
  XNOR2_X1 U16443 ( .A(n12060), .B(n12061), .ZN(n12951) );
  INV_X1 U16444 ( .A(n12951), .ZN(n13330) );
  XNOR2_X1 U16445 ( .A(n12064), .B(n12063), .ZN(n12071) );
  XNOR2_X1 U16446 ( .A(n12065), .B(n12066), .ZN(n12069) );
  XNOR2_X1 U16447 ( .A(n12067), .B(n3183), .ZN(n12068) );
  XNOR2_X1 U16448 ( .A(n12069), .B(n12068), .ZN(n12070) );
  NAND2_X1 U16449 ( .A1(n24588), .A2(n14306), .ZN(n12120) );
  XNOR2_X1 U16450 ( .A(n12074), .B(n12073), .ZN(n12079) );
  XNOR2_X1 U16451 ( .A(n12075), .B(n12183), .ZN(n12077) );
  XNOR2_X1 U16452 ( .A(n12128), .B(n21623), .ZN(n12076) );
  XNOR2_X1 U16453 ( .A(n12077), .B(n12076), .ZN(n12078) );
  XNOR2_X1 U16454 ( .A(n12080), .B(n12081), .ZN(n12086) );
  XNOR2_X1 U16455 ( .A(n12082), .B(n12226), .ZN(n12084) );
  XNOR2_X1 U16456 ( .A(n12159), .B(n21711), .ZN(n12083) );
  XNOR2_X1 U16457 ( .A(n12084), .B(n12083), .ZN(n12085) );
  XNOR2_X1 U16458 ( .A(n12086), .B(n12085), .ZN(n12840) );
  INV_X1 U16459 ( .A(n12840), .ZN(n13338) );
  NOR2_X1 U16460 ( .A1(n231), .A2(n13338), .ZN(n12107) );
  XNOR2_X1 U16461 ( .A(n12087), .B(n12088), .ZN(n12093) );
  XNOR2_X1 U16462 ( .A(n24323), .B(n1891), .ZN(n12090) );
  XNOR2_X1 U16463 ( .A(n12091), .B(n12090), .ZN(n12092) );
  XNOR2_X1 U16464 ( .A(n12092), .B(n12093), .ZN(n12576) );
  XNOR2_X1 U16465 ( .A(n12095), .B(n12094), .ZN(n12100) );
  XNOR2_X1 U16466 ( .A(n12122), .B(n1739), .ZN(n12097) );
  XNOR2_X1 U16467 ( .A(n12098), .B(n12097), .ZN(n12099) );
  XNOR2_X1 U16468 ( .A(n12151), .B(n11897), .ZN(n12104) );
  AOI21_X1 U16470 ( .B1(n13335), .B2(n13341), .A(n231), .ZN(n12119) );
  INV_X1 U16471 ( .A(n12839), .ZN(n12118) );
  XNOR2_X1 U16472 ( .A(n12109), .B(n12108), .ZN(n12111) );
  XNOR2_X1 U16473 ( .A(n12110), .B(n12111), .ZN(n12116) );
  XNOR2_X1 U16474 ( .A(n25027), .B(n3089), .ZN(n12113) );
  NAND2_X1 U16475 ( .A1(n231), .A2(n12956), .ZN(n12642) );
  INV_X1 U16476 ( .A(n12642), .ZN(n12117) );
  XNOR2_X1 U16477 ( .A(n12122), .B(n1776), .ZN(n12123) );
  XNOR2_X1 U16478 ( .A(n12124), .B(n12123), .ZN(n12125) );
  XNOR2_X1 U16479 ( .A(n12130), .B(n12129), .ZN(n12131) );
  INV_X1 U16480 ( .A(n12132), .ZN(n12133) );
  INV_X1 U16481 ( .A(n13358), .ZN(n13366) );
  XNOR2_X1 U16482 ( .A(n12134), .B(n21335), .ZN(n12135) );
  XNOR2_X1 U16483 ( .A(n12136), .B(n12135), .ZN(n12140) );
  XNOR2_X1 U16484 ( .A(n24970), .B(n25236), .ZN(n12139) );
  XNOR2_X1 U16485 ( .A(n12140), .B(n12139), .ZN(n12142) );
  XNOR2_X1 U16486 ( .A(n12142), .B(n12141), .ZN(n12625) );
  XNOR2_X1 U16487 ( .A(n12143), .B(n20995), .ZN(n12145) );
  XNOR2_X1 U16488 ( .A(n12145), .B(n12144), .ZN(n12149) );
  XNOR2_X1 U16489 ( .A(n12147), .B(n12146), .ZN(n12148) );
  XNOR2_X1 U16490 ( .A(n12149), .B(n12148), .ZN(n12155) );
  XNOR2_X1 U16491 ( .A(n12151), .B(n25032), .ZN(n12153) );
  XNOR2_X1 U16492 ( .A(n12152), .B(n12153), .ZN(n12154) );
  XNOR2_X2 U16493 ( .A(n12155), .B(n12154), .ZN(n12980) );
  INV_X1 U16494 ( .A(n12980), .ZN(n13359) );
  AOI22_X1 U16495 ( .A1(n24552), .A2(n13366), .B1(n12625), .B2(n13359), .ZN(
        n12175) );
  INV_X1 U16496 ( .A(n12156), .ZN(n12158) );
  XNOR2_X1 U16497 ( .A(n12157), .B(n12158), .ZN(n12164) );
  XNOR2_X1 U16498 ( .A(n12159), .B(n22886), .ZN(n12160) );
  XNOR2_X1 U16499 ( .A(n12160), .B(n12391), .ZN(n12162) );
  XNOR2_X1 U16500 ( .A(n12161), .B(n12162), .ZN(n12163) );
  XNOR2_X1 U16501 ( .A(n12164), .B(n12163), .ZN(n12583) );
  XNOR2_X1 U16503 ( .A(n12165), .B(n12166), .ZN(n12172) );
  XNOR2_X1 U16504 ( .A(n12167), .B(n24323), .ZN(n12170) );
  XNOR2_X1 U16505 ( .A(n12168), .B(n1896), .ZN(n12169) );
  XNOR2_X1 U16506 ( .A(n12170), .B(n12169), .ZN(n12171) );
  NAND2_X1 U16507 ( .A1(n13358), .A2(n12976), .ZN(n12626) );
  INV_X1 U16508 ( .A(n12626), .ZN(n12173) );
  AOI22_X1 U16509 ( .A1(n12173), .A2(n12878), .B1(n13366), .B2(n12980), .ZN(
        n12174) );
  OAI21_X1 U16510 ( .B1(n12175), .B2(n12977), .A(n12174), .ZN(n13453) );
  INV_X1 U16511 ( .A(n13453), .ZN(n13947) );
  MUX2_X2 U16512 ( .A(n12177), .B(n12176), .S(n13947), .Z(n15416) );
  XNOR2_X1 U16513 ( .A(n15416), .B(n14732), .ZN(n14691) );
  INV_X1 U16514 ( .A(n14691), .ZN(n15176) );
  INV_X1 U16515 ( .A(n12178), .ZN(n13093) );
  INV_X1 U16516 ( .A(n14311), .ZN(n13733) );
  XNOR2_X1 U16517 ( .A(n12182), .B(n12181), .ZN(n12188) );
  XNOR2_X1 U16518 ( .A(n12184), .B(n12183), .ZN(n12185) );
  XNOR2_X1 U16519 ( .A(n12186), .B(n12185), .ZN(n12187) );
  INV_X1 U16520 ( .A(n12854), .ZN(n13107) );
  XNOR2_X1 U16521 ( .A(n12334), .B(n12189), .ZN(n12191) );
  XNOR2_X1 U16522 ( .A(n12191), .B(n12190), .ZN(n12195) );
  XNOR2_X1 U16523 ( .A(n12193), .B(n12192), .ZN(n12194) );
  XNOR2_X1 U16524 ( .A(n12195), .B(n12194), .ZN(n13112) );
  INV_X1 U16525 ( .A(n13112), .ZN(n12673) );
  XNOR2_X1 U16526 ( .A(n12197), .B(n12196), .ZN(n12199) );
  XNOR2_X1 U16527 ( .A(n12198), .B(n12199), .ZN(n12205) );
  XNOR2_X1 U16528 ( .A(n12344), .B(n2042), .ZN(n12203) );
  XNOR2_X1 U16529 ( .A(n12203), .B(n12202), .ZN(n12204) );
  NAND2_X1 U16530 ( .A1(n3827), .A2(n12856), .ZN(n12633) );
  XNOR2_X1 U16531 ( .A(n12209), .B(n12208), .ZN(n12211) );
  XNOR2_X1 U16532 ( .A(n12210), .B(n12211), .ZN(n12217) );
  XNOR2_X1 U16533 ( .A(n12214), .B(n12215), .ZN(n12216) );
  XNOR2_X1 U16534 ( .A(n12217), .B(n12216), .ZN(n12672) );
  INV_X1 U16535 ( .A(n12672), .ZN(n13109) );
  XNOR2_X1 U16536 ( .A(n12219), .B(n12220), .ZN(n12223) );
  XNOR2_X1 U16537 ( .A(n12221), .B(n12315), .ZN(n12222) );
  XNOR2_X1 U16538 ( .A(n12223), .B(n12222), .ZN(n12229) );
  XNOR2_X1 U16539 ( .A(n12225), .B(n12224), .ZN(n12227) );
  XNOR2_X1 U16540 ( .A(n24915), .B(n12227), .ZN(n12228) );
  INV_X1 U16541 ( .A(n12230), .ZN(n12232) );
  XNOR2_X1 U16542 ( .A(n12248), .B(n12295), .ZN(n12231) );
  XNOR2_X1 U16543 ( .A(n12232), .B(n12231), .ZN(n12238) );
  XNOR2_X1 U16544 ( .A(n12234), .B(n20284), .ZN(n12235) );
  XNOR2_X1 U16545 ( .A(n12236), .B(n12235), .ZN(n12237) );
  INV_X1 U16546 ( .A(n13110), .ZN(n12674) );
  INV_X1 U16547 ( .A(n12239), .ZN(n12240) );
  XNOR2_X1 U16548 ( .A(n12241), .B(n1767), .ZN(n12243) );
  XNOR2_X1 U16549 ( .A(n12243), .B(n12242), .ZN(n12244) );
  XNOR2_X1 U16550 ( .A(n12245), .B(n12244), .ZN(n12868) );
  XNOR2_X1 U16551 ( .A(n12247), .B(n12246), .ZN(n12254) );
  XNOR2_X1 U16552 ( .A(n12249), .B(n12248), .ZN(n12252) );
  XNOR2_X1 U16553 ( .A(n24323), .B(n1826), .ZN(n12251) );
  XNOR2_X1 U16554 ( .A(n12251), .B(n12252), .ZN(n12253) );
  XNOR2_X1 U16555 ( .A(n12255), .B(n2120), .ZN(n12256) );
  XNOR2_X1 U16556 ( .A(n12256), .B(n12257), .ZN(n12258) );
  XNOR2_X1 U16557 ( .A(n12258), .B(n12259), .ZN(n12265) );
  XNOR2_X1 U16558 ( .A(n12260), .B(n24987), .ZN(n12262) );
  XNOR2_X1 U16559 ( .A(n12263), .B(n12262), .ZN(n12264) );
  XNOR2_X1 U16561 ( .A(n12267), .B(n12266), .ZN(n12271) );
  INV_X1 U16562 ( .A(n12268), .ZN(n12270) );
  NOR2_X1 U16563 ( .A1(n12865), .A2(n12272), .ZN(n12659) );
  XNOR2_X1 U16564 ( .A(n12274), .B(n12273), .ZN(n12281) );
  XNOR2_X1 U16565 ( .A(n12276), .B(n12275), .ZN(n12279) );
  XNOR2_X1 U16566 ( .A(n12277), .B(n5131), .ZN(n12278) );
  XNOR2_X1 U16567 ( .A(n12279), .B(n12278), .ZN(n12280) );
  XNOR2_X1 U16568 ( .A(n12281), .B(n12280), .ZN(n12864) );
  INV_X1 U16569 ( .A(n12864), .ZN(n12503) );
  XNOR2_X1 U16570 ( .A(n12282), .B(n12283), .ZN(n12285) );
  XNOR2_X1 U16571 ( .A(n12285), .B(n12284), .ZN(n12290) );
  XNOR2_X1 U16572 ( .A(n12286), .B(n1789), .ZN(n12287) );
  XNOR2_X1 U16573 ( .A(n12288), .B(n12287), .ZN(n12289) );
  NOR2_X1 U16574 ( .A1(n13114), .A2(n3327), .ZN(n12291) );
  INV_X1 U16575 ( .A(n12292), .ZN(n12294) );
  XNOR2_X1 U16576 ( .A(n12294), .B(n12293), .ZN(n12301) );
  XNOR2_X1 U16577 ( .A(n12295), .B(n12296), .ZN(n12299) );
  XNOR2_X1 U16578 ( .A(n12297), .B(n2882), .ZN(n12298) );
  XNOR2_X1 U16579 ( .A(n12299), .B(n12298), .ZN(n12300) );
  INV_X1 U16580 ( .A(n13123), .ZN(n12874) );
  INV_X1 U16581 ( .A(n12302), .ZN(n12305) );
  INV_X1 U16582 ( .A(n12303), .ZN(n12304) );
  XNOR2_X1 U16583 ( .A(n12304), .B(n12305), .ZN(n12310) );
  XNOR2_X1 U16584 ( .A(n12306), .B(n3084), .ZN(n12308) );
  XNOR2_X1 U16585 ( .A(n12308), .B(n12307), .ZN(n12309) );
  XNOR2_X1 U16587 ( .A(n12312), .B(n12311), .ZN(n12319) );
  XNOR2_X1 U16588 ( .A(n12314), .B(n12313), .ZN(n12317) );
  XNOR2_X1 U16589 ( .A(n12315), .B(n2240), .ZN(n12316) );
  XNOR2_X1 U16590 ( .A(n12317), .B(n12316), .ZN(n12318) );
  XNOR2_X1 U16591 ( .A(n12319), .B(n12318), .ZN(n12349) );
  INV_X1 U16592 ( .A(n12320), .ZN(n12321) );
  XNOR2_X1 U16593 ( .A(n12321), .B(n12322), .ZN(n12329) );
  XNOR2_X1 U16594 ( .A(n12324), .B(n12323), .ZN(n12327) );
  XNOR2_X1 U16595 ( .A(n12325), .B(n1797), .ZN(n12326) );
  XNOR2_X1 U16596 ( .A(n12327), .B(n12326), .ZN(n12328) );
  INV_X1 U16597 ( .A(n13354), .ZN(n12332) );
  NAND2_X1 U16598 ( .A1(n13352), .A2(n13123), .ZN(n13122) );
  INV_X1 U16599 ( .A(n13122), .ZN(n12331) );
  XNOR2_X1 U16600 ( .A(n12334), .B(n12333), .ZN(n12337) );
  XNOR2_X1 U16601 ( .A(n12335), .B(n3073), .ZN(n12336) );
  XNOR2_X1 U16602 ( .A(n12339), .B(n12338), .ZN(n12340) );
  XNOR2_X1 U16603 ( .A(n12343), .B(n11915), .ZN(n12346) );
  XNOR2_X1 U16604 ( .A(n12344), .B(n899), .ZN(n12345) );
  XNOR2_X1 U16605 ( .A(n12346), .B(n12345), .ZN(n12347) );
  INV_X1 U16606 ( .A(n12349), .ZN(n13351) );
  NAND2_X1 U16607 ( .A1(n406), .A2(n13351), .ZN(n12350) );
  XNOR2_X1 U16608 ( .A(n12351), .B(n12352), .ZN(n12353) );
  XNOR2_X1 U16609 ( .A(n12354), .B(n12353), .ZN(n12361) );
  XNOR2_X1 U16610 ( .A(n12356), .B(n12355), .ZN(n12359) );
  XNOR2_X1 U16611 ( .A(n12357), .B(n1833), .ZN(n12358) );
  XNOR2_X1 U16612 ( .A(n12359), .B(n12358), .ZN(n12360) );
  XNOR2_X1 U16613 ( .A(n12362), .B(n12363), .ZN(n12367) );
  XNOR2_X1 U16614 ( .A(n12364), .B(n12365), .ZN(n12366) );
  XNOR2_X1 U16615 ( .A(n12366), .B(n12367), .ZN(n12374) );
  XNOR2_X1 U16616 ( .A(n12370), .B(n4034), .ZN(n12371) );
  XNOR2_X1 U16617 ( .A(n12372), .B(n12371), .ZN(n12373) );
  XNOR2_X1 U16618 ( .A(n12375), .B(n12376), .ZN(n12380) );
  XNOR2_X1 U16619 ( .A(n12378), .B(n12377), .ZN(n12379) );
  XNOR2_X1 U16620 ( .A(n12379), .B(n12380), .ZN(n12387) );
  XNOR2_X1 U16622 ( .A(n24964), .B(n494), .ZN(n12384) );
  XNOR2_X1 U16623 ( .A(n12385), .B(n12384), .ZN(n12386) );
  XNOR2_X1 U16624 ( .A(n12387), .B(n12386), .ZN(n12859) );
  XNOR2_X1 U16625 ( .A(n12388), .B(n2031), .ZN(n12390) );
  XNOR2_X1 U16626 ( .A(n12390), .B(n12389), .ZN(n12393) );
  XNOR2_X1 U16627 ( .A(n12393), .B(n12392), .ZN(n12394) );
  NAND2_X1 U16629 ( .A1(n12859), .A2(n13344), .ZN(n12407) );
  XNOR2_X1 U16630 ( .A(n12396), .B(n23983), .ZN(n12398) );
  XNOR2_X1 U16631 ( .A(n12398), .B(n12397), .ZN(n12399) );
  XNOR2_X1 U16632 ( .A(n12400), .B(n12399), .ZN(n12406) );
  XNOR2_X1 U16633 ( .A(n12402), .B(n12401), .ZN(n12403) );
  XNOR2_X1 U16634 ( .A(n12404), .B(n12403), .ZN(n12405) );
  XNOR2_X1 U16635 ( .A(n12406), .B(n12405), .ZN(n13347) );
  NAND2_X1 U16636 ( .A1(n13347), .A2(n12636), .ZN(n12419) );
  XNOR2_X1 U16637 ( .A(n12408), .B(n2126), .ZN(n12412) );
  XNOR2_X1 U16638 ( .A(n12412), .B(n12411), .ZN(n12418) );
  XNOR2_X1 U16639 ( .A(n12414), .B(n12413), .ZN(n12415) );
  XNOR2_X1 U16640 ( .A(n12416), .B(n12415), .ZN(n12417) );
  AOI21_X1 U16642 ( .B1(n12419), .B2(n13345), .A(n12859), .ZN(n12420) );
  NOR2_X1 U16643 ( .A1(n12421), .A2(n12420), .ZN(n13903) );
  INV_X1 U16644 ( .A(n12422), .ZN(n12424) );
  NOR3_X1 U16645 ( .A1(n13903), .A2(n12424), .A3(n12423), .ZN(n14310) );
  INV_X1 U16646 ( .A(n14310), .ZN(n12425) );
  OAI21_X1 U16647 ( .B1(n13959), .B2(n13958), .A(n12425), .ZN(n12427) );
  INV_X1 U16648 ( .A(n13132), .ZN(n13129) );
  INV_X1 U16649 ( .A(n12498), .ZN(n13131) );
  INV_X1 U16650 ( .A(n12483), .ZN(n12712) );
  INV_X1 U16651 ( .A(n12707), .ZN(n12711) );
  INV_X1 U16652 ( .A(n12710), .ZN(n12431) );
  INV_X1 U16653 ( .A(n12433), .ZN(n13145) );
  NAND3_X1 U16654 ( .A1(n13145), .A2(n12729), .A3(n13144), .ZN(n12438) );
  NAND2_X1 U16655 ( .A1(n13144), .A2(n12455), .ZN(n13146) );
  INV_X1 U16656 ( .A(n13146), .ZN(n12434) );
  NAND2_X1 U16657 ( .A1(n12434), .A2(n12728), .ZN(n12436) );
  NAND3_X1 U16658 ( .A1(n13140), .A2(n12729), .A3(n13143), .ZN(n12435) );
  MUX2_X1 U16659 ( .A(n24601), .B(n13061), .S(n13063), .Z(n12441) );
  NAND3_X1 U16660 ( .A1(n13049), .A2(n12490), .A3(n12535), .ZN(n12442) );
  NOR2_X1 U16661 ( .A1(n14166), .A2(n14168), .ZN(n12445) );
  INV_X1 U16662 ( .A(n12774), .ZN(n13068) );
  NAND2_X1 U16663 ( .A1(n13068), .A2(n12773), .ZN(n12472) );
  NOR2_X1 U16664 ( .A1(n13067), .A2(n12470), .ZN(n12530) );
  INV_X1 U16665 ( .A(n12469), .ZN(n12778) );
  OAI21_X1 U16666 ( .B1(n12530), .B2(n1439), .A(n12778), .ZN(n12446) );
  AND2_X1 U16667 ( .A1(n14165), .A2(n13744), .ZN(n13745) );
  AOI21_X1 U16668 ( .B1(n12718), .B2(n12447), .A(n304), .ZN(n12448) );
  NAND2_X1 U16669 ( .A1(n13745), .A2(n13742), .ZN(n13529) );
  MUX2_X1 U16671 ( .A(n13165), .B(n24930), .S(n24373), .Z(n12453) );
  NAND2_X1 U16672 ( .A1(n13170), .A2(n24930), .ZN(n12452) );
  NAND2_X1 U16673 ( .A1(n13137), .A2(n13144), .ZN(n12458) );
  OAI211_X1 U16674 ( .C1(n13144), .C2(n12455), .A(n13140), .B(n13136), .ZN(
        n12457) );
  NAND3_X1 U16675 ( .A1(n11109), .A2(n13138), .A3(n13143), .ZN(n12456) );
  AOI21_X1 U16676 ( .B1(n1355), .B2(n14049), .A(n14050), .ZN(n12468) );
  NAND2_X1 U16677 ( .A1(n12462), .A2(n12715), .ZN(n12482) );
  OAI21_X1 U16678 ( .B1(n12710), .B2(n12707), .A(n12713), .ZN(n12461) );
  OAI21_X1 U16679 ( .B1(n12712), .B2(n24573), .A(n12710), .ZN(n12463) );
  AOI22_X1 U16680 ( .A1(n12490), .A2(n12534), .B1(n25408), .B2(n13049), .ZN(
        n12466) );
  OAI21_X2 U16681 ( .B1(n12466), .B2(n13048), .A(n12465), .ZN(n14054) );
  AND2_X1 U16682 ( .A1(n14054), .A2(n13521), .ZN(n13611) );
  NAND2_X1 U16683 ( .A1(n14049), .A2(n14048), .ZN(n12820) );
  INV_X1 U16684 ( .A(n12820), .ZN(n12467) );
  XNOR2_X1 U16685 ( .A(n15054), .B(n2005), .ZN(n12518) );
  AND2_X1 U16686 ( .A1(n12774), .A2(n12470), .ZN(n13073) );
  AND2_X1 U16687 ( .A1(n12469), .A2(n12470), .ZN(n12532) );
  AOI21_X1 U16688 ( .B1(n12774), .B2(n12471), .A(n12470), .ZN(n12473) );
  AND2_X1 U16689 ( .A1(n12472), .A2(n12473), .ZN(n12474) );
  INV_X1 U16690 ( .A(n12520), .ZN(n12478) );
  NAND2_X1 U16691 ( .A1(n12478), .A2(n12476), .ZN(n12477) );
  NAND3_X1 U16693 ( .A1(n12799), .A2(n12478), .A3(n13044), .ZN(n12479) );
  NAND2_X1 U16694 ( .A1(n12796), .A2(n12484), .ZN(n12488) );
  NOR2_X1 U16695 ( .A1(n25085), .A2(n409), .ZN(n12486) );
  AOI22_X1 U16696 ( .A1(n3065), .A2(n12486), .B1(n12485), .B2(n25085), .ZN(
        n12487) );
  AOI22_X1 U16697 ( .A1(n14241), .A2(n25209), .B1(n13931), .B2(n13200), .ZN(
        n12497) );
  OAI211_X1 U16698 ( .C1(n12534), .C2(n12535), .A(n25494), .B(n13048), .ZN(
        n12492) );
  NAND3_X1 U16699 ( .A1(n12490), .A2(n12489), .A3(n13051), .ZN(n12491) );
  INV_X1 U16700 ( .A(n14244), .ZN(n12496) );
  NAND2_X1 U16702 ( .A1(n25369), .A2(n12786), .ZN(n12493) );
  AOI22_X1 U16703 ( .A1(n12494), .A2(n13029), .B1(n12493), .B2(n302), .ZN(
        n13635) );
  INV_X1 U16704 ( .A(n13635), .ZN(n14240) );
  NOR2_X1 U16706 ( .A1(n13132), .A2(n13150), .ZN(n12500) );
  NOR2_X1 U16707 ( .A1(n13151), .A2(n12498), .ZN(n12499) );
  NAND2_X1 U16708 ( .A1(n13145), .A2(n13139), .ZN(n12502) );
  NAND2_X1 U16709 ( .A1(n14090), .A2(n13533), .ZN(n12509) );
  AOI22_X1 U16710 ( .A1(n12659), .A2(n12864), .B1(n13119), .B2(n13114), .ZN(
        n13536) );
  NAND3_X1 U16711 ( .A1(n3328), .A2(n12864), .A3(n12660), .ZN(n12504) );
  NAND2_X1 U16712 ( .A1(n5324), .A2(n13092), .ZN(n12650) );
  MUX2_X1 U16713 ( .A(n12506), .B(n10360), .S(n12459), .Z(n12508) );
  NAND2_X1 U16714 ( .A1(n12652), .A2(n12724), .ZN(n12507) );
  AOI21_X1 U16715 ( .B1(n12509), .B2(n12817), .A(n14018), .ZN(n12515) );
  NAND2_X1 U16717 ( .A1(n13102), .A2(n13187), .ZN(n13183) );
  INV_X1 U16718 ( .A(n13187), .ZN(n13103) );
  NAND2_X1 U16719 ( .A1(n13103), .A2(n12656), .ZN(n13191) );
  NAND3_X1 U16720 ( .A1(n13183), .A2(n13185), .A3(n13191), .ZN(n13535) );
  AOI21_X1 U16721 ( .B1(n14085), .B2(n12513), .A(n14090), .ZN(n12514) );
  NOR2_X2 U16722 ( .A1(n12515), .A2(n12514), .ZN(n15056) );
  INV_X1 U16723 ( .A(n15056), .ZN(n12516) );
  XNOR2_X1 U16724 ( .A(n14377), .B(n12516), .ZN(n12517) );
  XNOR2_X1 U16725 ( .A(n12518), .B(n12517), .ZN(n12620) );
  MUX2_X1 U16726 ( .A(n12800), .B(n12523), .S(n13041), .Z(n12522) );
  NOR2_X1 U16727 ( .A1(n13044), .A2(n12523), .ZN(n12521) );
  NAND2_X1 U16728 ( .A1(n12523), .A2(n13040), .ZN(n13045) );
  NOR2_X1 U16731 ( .A1(n12753), .A2(n25085), .ZN(n12528) );
  NOR2_X2 U16732 ( .A1(n12529), .A2(n12528), .ZN(n13840) );
  NAND2_X1 U16733 ( .A1(n12774), .A2(n13071), .ZN(n12531) );
  NOR2_X1 U16734 ( .A1(n13840), .A2(n397), .ZN(n12537) );
  MUX2_X1 U16735 ( .A(n13023), .B(n13028), .S(n12786), .Z(n12538) );
  NAND2_X1 U16736 ( .A1(n12786), .A2(n13028), .ZN(n13025) );
  INV_X1 U16737 ( .A(n13623), .ZN(n12543) );
  AOI22_X1 U16738 ( .A1(n12543), .A2(n13839), .B1(n12542), .B2(n13837), .ZN(
        n12544) );
  NOR2_X1 U16739 ( .A1(n12546), .A2(n13298), .ZN(n12549) );
  NAND2_X1 U16740 ( .A1(n13301), .A2(n12902), .ZN(n12903) );
  NAND2_X1 U16741 ( .A1(n12546), .A2(n12903), .ZN(n13239) );
  NOR2_X1 U16742 ( .A1(n13239), .A2(n405), .ZN(n13853) );
  INV_X1 U16743 ( .A(n13211), .ZN(n13205) );
  OAI21_X1 U16744 ( .B1(n13205), .B2(n13207), .A(n13213), .ZN(n12550) );
  AND2_X1 U16745 ( .A1(n13000), .A2(n13207), .ZN(n13001) );
  NOR2_X1 U16746 ( .A1(n12551), .A2(n13207), .ZN(n12552) );
  NOR2_X2 U16747 ( .A1(n12553), .A2(n12552), .ZN(n12704) );
  INV_X1 U16748 ( .A(n12704), .ZN(n14074) );
  OAI21_X1 U16749 ( .B1(n12611), .B2(n12555), .A(n12914), .ZN(n12554) );
  NAND2_X1 U16750 ( .A1(n24487), .A2(n12554), .ZN(n12557) );
  INV_X1 U16751 ( .A(n13245), .ZN(n12559) );
  NAND3_X1 U16752 ( .A1(n13244), .A2(n13011), .A3(n12559), .ZN(n12562) );
  NAND2_X1 U16753 ( .A1(n12563), .A2(n13246), .ZN(n12564) );
  NAND2_X1 U16756 ( .A1(n13009), .A2(n13222), .ZN(n12568) );
  OAI211_X1 U16757 ( .C1(n24965), .C2(n13009), .A(n24490), .B(n12568), .ZN(
        n12572) );
  OAI21_X1 U16758 ( .B1(n14075), .B2(n14076), .A(n14077), .ZN(n12573) );
  NAND2_X1 U16759 ( .A1(n12573), .A2(n12704), .ZN(n12574) );
  XNOR2_X1 U16760 ( .A(n14857), .B(n15169), .ZN(n15408) );
  NOR2_X1 U16761 ( .A1(n12838), .A2(n13336), .ZN(n12579) );
  NAND2_X1 U16764 ( .A1(n12577), .A2(n12839), .ZN(n12578) );
  INV_X1 U16765 ( .A(n12688), .ZN(n12947) );
  MUX2_X1 U16766 ( .A(n25053), .B(n12980), .S(n12976), .Z(n12586) );
  INV_X1 U16767 ( .A(n24554), .ZN(n13365) );
  AOI21_X1 U16768 ( .B1(n12586), .B2(n13365), .A(n12585), .ZN(n13847) );
  OAI21_X1 U16770 ( .B1(n13108), .B2(n12856), .A(n12672), .ZN(n12587) );
  NOR3_X1 U16771 ( .A1(n13109), .A2(n13112), .A3(n13108), .ZN(n12588) );
  MUX2_X1 U16772 ( .A(n25430), .B(n13123), .S(n13124), .Z(n12590) );
  INV_X1 U16773 ( .A(n14064), .ZN(n13426) );
  NOR2_X1 U16775 ( .A1(n13291), .A2(n12593), .ZN(n12596) );
  AND2_X1 U16778 ( .A1(n12600), .A2(n13272), .ZN(n12965) );
  NAND2_X1 U16779 ( .A1(n13275), .A2(n12695), .ZN(n12602) );
  NAND2_X1 U16780 ( .A1(n12834), .A2(n13274), .ZN(n12601) );
  MUX2_X1 U16781 ( .A(n12602), .B(n12601), .S(n24346), .Z(n12603) );
  INV_X1 U16782 ( .A(n13325), .ZN(n12683) );
  OAI21_X1 U16783 ( .B1(n12955), .B2(n12604), .A(n13329), .ZN(n12605) );
  NAND2_X1 U16784 ( .A1(n14849), .A2(n14852), .ZN(n12617) );
  INV_X1 U16785 ( .A(n12900), .ZN(n13282) );
  AND2_X1 U16787 ( .A1(n12900), .A2(n11873), .ZN(n12925) );
  NAND2_X1 U16788 ( .A1(n12614), .A2(n24572), .ZN(n12616) );
  AND2_X1 U16789 ( .A1(n14059), .A2(n14278), .ZN(n14280) );
  NAND2_X1 U16790 ( .A1(n14280), .A2(n14849), .ZN(n12615) );
  OAI211_X1 U16791 ( .C1(n24572), .C2(n12617), .A(n12616), .B(n12615), .ZN(
        n14721) );
  XNOR2_X1 U16793 ( .A(n14699), .B(n15408), .ZN(n12619) );
  INV_X1 U16794 ( .A(n13350), .ZN(n13125) );
  NAND2_X1 U16795 ( .A1(n5624), .A2(n12349), .ZN(n12622) );
  INV_X1 U16797 ( .A(n12976), .ZN(n13364) );
  INV_X1 U16799 ( .A(n12625), .ZN(n13357) );
  INV_X1 U16800 ( .A(n12865), .ZN(n13117) );
  INV_X1 U16801 ( .A(n12660), .ZN(n13116) );
  OAI21_X1 U16802 ( .B1(n3328), .B2(n13116), .A(n13114), .ZN(n12630) );
  NAND2_X1 U16803 ( .A1(n12854), .A2(n13108), .ZN(n12634) );
  NAND3_X1 U16804 ( .A1(n12673), .A2(n4923), .A3(n13107), .ZN(n12635) );
  NAND2_X1 U16805 ( .A1(n3889), .A2(n3888), .ZN(n12646) );
  NOR2_X1 U16806 ( .A1(n25415), .A2(n25366), .ZN(n12637) );
  INV_X1 U16807 ( .A(n14198), .ZN(n14946) );
  MUX2_X1 U16808 ( .A(n13335), .B(n12956), .S(n13341), .Z(n12644) );
  INV_X1 U16809 ( .A(n12960), .ZN(n12643) );
  NAND2_X1 U16810 ( .A1(n13336), .A2(n12956), .ZN(n12640) );
  NAND2_X1 U16811 ( .A1(n13337), .A2(n12640), .ZN(n12641) );
  NAND2_X1 U16813 ( .A1(n2570), .A2(n2684), .ZN(n12645) );
  OAI21_X1 U16814 ( .B1(n12646), .B2(n14946), .A(n12645), .ZN(n12647) );
  INV_X1 U16815 ( .A(n14988), .ZN(n12679) );
  INV_X1 U16817 ( .A(n14003), .ZN(n13484) );
  INV_X1 U16818 ( .A(n13102), .ZN(n12744) );
  NAND2_X1 U16819 ( .A1(n12744), .A2(n12656), .ZN(n12655) );
  OAI211_X1 U16820 ( .C1(n12744), .C2(n12742), .A(n12655), .B(n12654), .ZN(
        n12658) );
  NAND3_X1 U16821 ( .A1(n13185), .A2(n12656), .A3(n12740), .ZN(n12657) );
  INV_X1 U16822 ( .A(n12668), .ZN(n13486) );
  INV_X1 U16823 ( .A(n12659), .ZN(n12662) );
  NOR2_X1 U16824 ( .A1(n12868), .A2(n12660), .ZN(n12661) );
  INV_X1 U16825 ( .A(n13130), .ZN(n13149) );
  NOR2_X1 U16826 ( .A1(n13129), .A2(n13149), .ZN(n12665) );
  NOR2_X1 U16827 ( .A1(n13131), .A2(n13152), .ZN(n12664) );
  INV_X1 U16828 ( .A(n5754), .ZN(n12667) );
  OAI22_X1 U16829 ( .A1(n13158), .A2(n13150), .B1(n12667), .B2(n13130), .ZN(
        n13660) );
  NAND2_X1 U16830 ( .A1(n14002), .A2(n12669), .ZN(n12670) );
  INV_X1 U16832 ( .A(n13262), .ZN(n12676) );
  MUX2_X1 U16833 ( .A(n13265), .B(n13266), .S(n5361), .Z(n12682) );
  NAND2_X1 U16835 ( .A1(n13329), .A2(n13323), .ZN(n12685) );
  NAND2_X1 U16836 ( .A1(n13788), .A2(n14143), .ZN(n12703) );
  OAI21_X1 U16839 ( .B1(n13316), .B2(n25499), .A(n12945), .ZN(n12689) );
  NOR2_X1 U16840 ( .A1(n12827), .A2(n24476), .ZN(n12691) );
  OAI21_X1 U16841 ( .B1(n12692), .B2(n12691), .A(n12690), .ZN(n12693) );
  INV_X1 U16842 ( .A(n13275), .ZN(n12964) );
  NOR2_X1 U16843 ( .A1(n13785), .A2(n14143), .ZN(n13789) );
  OAI21_X1 U16844 ( .B1(n12897), .B2(n13282), .A(n24988), .ZN(n12699) );
  OAI21_X1 U16845 ( .B1(n13789), .B2(n14142), .A(n24347), .ZN(n12701) );
  XNOR2_X1 U16848 ( .A(n15070), .B(n15185), .ZN(n12783) );
  MUX2_X1 U16849 ( .A(n12721), .B(n12720), .S(n24930), .Z(n12722) );
  NOR2_X1 U16851 ( .A1(n14440), .A2(n24556), .ZN(n13257) );
  OAI211_X1 U16853 ( .C1(n3974), .C2(n13178), .A(n13177), .B(n12724), .ZN(
        n12727) );
  NAND2_X1 U16855 ( .A1(n12728), .A2(n13136), .ZN(n12731) );
  MUX2_X1 U16857 ( .A(n12731), .B(n12730), .S(n13138), .Z(n12732) );
  OAI22_X1 U16858 ( .A1(n24571), .A2(n24713), .B1(n14440), .B2(n14510), .ZN(
        n12739) );
  NAND2_X1 U16859 ( .A1(n12439), .A2(n1353), .ZN(n12738) );
  NAND2_X1 U16860 ( .A1(n25061), .A2(n13061), .ZN(n12736) );
  NAND2_X1 U16861 ( .A1(n12742), .A2(n24640), .ZN(n12743) );
  INV_X1 U16863 ( .A(n13188), .ZN(n12745) );
  AND2_X2 U16864 ( .A1(n12746), .A2(n12745), .ZN(n13693) );
  INV_X1 U16865 ( .A(n13693), .ZN(n14507) );
  NOR2_X1 U16866 ( .A1(n24556), .A2(n14507), .ZN(n13260) );
  XNOR2_X1 U16867 ( .A(n14911), .B(n1896), .ZN(n12781) );
  NAND2_X1 U16868 ( .A1(n14052), .A2(n14054), .ZN(n12749) );
  NAND3_X1 U16869 ( .A1(n13521), .A2(n14054), .A3(n1355), .ZN(n12747) );
  INV_X1 U16870 ( .A(n15184), .ZN(n12780) );
  NOR2_X1 U16871 ( .A1(n12796), .A2(n13053), .ZN(n12750) );
  NOR2_X1 U16872 ( .A1(n12751), .A2(n12750), .ZN(n12755) );
  NAND2_X1 U16873 ( .A1(n13053), .A2(n13057), .ZN(n12752) );
  AND2_X1 U16874 ( .A1(n12753), .A2(n12752), .ZN(n12754) );
  MUX2_X2 U16875 ( .A(n12755), .B(n12754), .S(n25085), .Z(n14178) );
  NAND2_X1 U16876 ( .A1(n12560), .A2(n13011), .ZN(n12756) );
  INV_X1 U16877 ( .A(n13011), .ZN(n13243) );
  OAI21_X1 U16878 ( .B1(n13244), .B2(n13243), .A(n13015), .ZN(n12757) );
  AOI22_X1 U16879 ( .A1(n13242), .A2(n13245), .B1(n13017), .B2(n12757), .ZN(
        n13578) );
  INV_X1 U16880 ( .A(n12761), .ZN(n12760) );
  INV_X1 U16881 ( .A(n12786), .ZN(n12759) );
  NAND3_X1 U16883 ( .A1(n2793), .A2(n12761), .A3(n13027), .ZN(n12762) );
  NAND2_X1 U16884 ( .A1(n24949), .A2(n13792), .ZN(n12771) );
  NOR2_X1 U16885 ( .A1(n4651), .A2(n13215), .ZN(n12764) );
  NAND2_X1 U16886 ( .A1(n12764), .A2(n13220), .ZN(n12766) );
  NAND2_X1 U16887 ( .A1(n12766), .A2(n12765), .ZN(n12770) );
  INV_X1 U16888 ( .A(n13217), .ZN(n12768) );
  INV_X1 U16889 ( .A(n12772), .ZN(n13769) );
  AOI21_X1 U16890 ( .B1(n13797), .B2(n12771), .A(n13769), .ZN(n12779) );
  AOI22_X1 U16891 ( .A1(n13067), .A2(n13066), .B1(n12774), .B2(n12773), .ZN(
        n12777) );
  NAND2_X1 U16892 ( .A1(n12775), .A2(n13068), .ZN(n12776) );
  XNOR2_X1 U16893 ( .A(n14669), .B(n12780), .ZN(n15367) );
  XNOR2_X1 U16894 ( .A(n15367), .B(n12781), .ZN(n12782) );
  XNOR2_X1 U16895 ( .A(n12783), .B(n12782), .ZN(n15822) );
  AND2_X1 U16897 ( .A1(n12787), .A2(n25369), .ZN(n12789) );
  NOR2_X1 U16898 ( .A1(n14327), .A2(n14041), .ZN(n12804) );
  NAND2_X1 U16899 ( .A1(n12800), .A2(n12799), .ZN(n12802) );
  NOR2_X1 U16900 ( .A1(n13045), .A2(n11580), .ZN(n12801) );
  AOI22_X1 U16901 ( .A1(n5230), .A2(n12804), .B1(n14327), .B2(n12803), .ZN(
        n12816) );
  MUX2_X1 U16902 ( .A(n25198), .B(n13011), .S(n12808), .Z(n12805) );
  MUX2_X1 U16904 ( .A(n12810), .B(n12809), .S(n24512), .Z(n12813) );
  NOR3_X1 U16905 ( .A1(n298), .A2(n14330), .A3(n14324), .ZN(n12815) );
  NAND2_X1 U16906 ( .A1(n13741), .A2(n13742), .ZN(n12818) );
  INV_X1 U16907 ( .A(n13742), .ZN(n14169) );
  NAND3_X1 U16908 ( .A1(n13526), .A2(n14169), .A3(n14167), .ZN(n12819) );
  XNOR2_X1 U16909 ( .A(n14900), .B(n1797), .ZN(n12852) );
  NAND2_X1 U16910 ( .A1(n12825), .A2(n13292), .ZN(n13507) );
  NOR2_X1 U16911 ( .A1(n12827), .A2(n13288), .ZN(n12826) );
  NAND2_X1 U16912 ( .A1(n13507), .A2(n13502), .ZN(n13877) );
  INV_X1 U16913 ( .A(n12830), .ZN(n12831) );
  OAI21_X1 U16914 ( .B1(n12832), .B2(n2632), .A(n12831), .ZN(n12833) );
  MUX2_X1 U16915 ( .A(n13278), .B(n13273), .S(n1200), .Z(n12837) );
  AOI22_X1 U16916 ( .A1(n12835), .A2(n13278), .B1(n13274), .B2(n12965), .ZN(
        n12836) );
  INV_X1 U16917 ( .A(n12956), .ZN(n12842) );
  OAI21_X1 U16919 ( .B1(n12840), .B2(n13341), .A(n13335), .ZN(n12841) );
  INV_X1 U16920 ( .A(n14339), .ZN(n14334) );
  NOR2_X1 U16921 ( .A1(n14333), .A2(n14339), .ZN(n14337) );
  NAND2_X1 U16922 ( .A1(n13318), .A2(n12844), .ZN(n12843) );
  INV_X1 U16923 ( .A(n13323), .ZN(n12952) );
  NOR2_X1 U16925 ( .A1(n13325), .A2(n3256), .ZN(n12849) );
  XNOR2_X1 U16929 ( .A(n12852), .B(n15347), .ZN(n12908) );
  NAND3_X1 U16931 ( .A1(n13109), .A2(n4923), .A3(n12856), .ZN(n12857) );
  INV_X1 U16932 ( .A(n13344), .ZN(n12860) );
  NOR2_X1 U16933 ( .A1(n14321), .A2(n13871), .ZN(n14457) );
  INV_X1 U16934 ( .A(n13114), .ZN(n12869) );
  MUX2_X1 U16935 ( .A(n3328), .B(n13116), .S(n12869), .Z(n12867) );
  NOR2_X1 U16936 ( .A1(n12864), .A2(n13113), .ZN(n12866) );
  INV_X1 U16937 ( .A(n14460), .ZN(n12883) );
  NAND2_X1 U16938 ( .A1(n13124), .A2(n13351), .ZN(n12872) );
  NOR2_X1 U16939 ( .A1(n24552), .A2(n12977), .ZN(n12876) );
  INV_X1 U16940 ( .A(n12981), .ZN(n12877) );
  NAND2_X1 U16941 ( .A1(n12877), .A2(n12878), .ZN(n12880) );
  NAND2_X1 U16942 ( .A1(n13366), .A2(n12976), .ZN(n12879) );
  NAND2_X1 U16943 ( .A1(n3401), .A2(n13868), .ZN(n12881) );
  OAI22_X1 U16944 ( .A1(n14459), .A2(n13868), .B1(n12881), .B2(n14321), .ZN(
        n12882) );
  NOR2_X1 U16945 ( .A1(n12884), .A2(n12924), .ZN(n12888) );
  INV_X1 U16946 ( .A(n13223), .ZN(n12919) );
  NAND2_X1 U16948 ( .A1(n13208), .A2(n12891), .ZN(n12896) );
  NOR2_X1 U16949 ( .A1(n5418), .A2(n11360), .ZN(n12894) );
  INV_X1 U16950 ( .A(n13208), .ZN(n12893) );
  NOR2_X1 U16951 ( .A1(n12899), .A2(n13282), .ZN(n12898) );
  AOI21_X1 U16952 ( .B1(n13283), .B2(n12900), .A(n12899), .ZN(n12901) );
  INV_X1 U16953 ( .A(n13806), .ZN(n12905) );
  NOR2_X1 U16954 ( .A1(n3859), .A2(n13305), .ZN(n12904) );
  NOR2_X1 U16955 ( .A1(n12905), .A2(n13513), .ZN(n12906) );
  NOR2_X2 U16956 ( .A1(n12907), .A2(n12906), .ZN(n14936) );
  XNOR2_X1 U16957 ( .A(n14936), .B(n14992), .ZN(n14714) );
  XNOR2_X1 U16958 ( .A(n12908), .B(n14714), .ZN(n12909) );
  AOI21_X1 U16959 ( .B1(n12911), .B2(n24476), .A(n12910), .ZN(n12912) );
  NOR3_X1 U16960 ( .A1(n12824), .A2(n13292), .A3(n13291), .ZN(n12913) );
  OAI21_X1 U16961 ( .B1(n13307), .B2(n13304), .A(n12915), .ZN(n12916) );
  AND2_X1 U16962 ( .A1(n12918), .A2(n13227), .ZN(n12923) );
  NOR2_X1 U16963 ( .A1(n12569), .A2(n13224), .ZN(n12921) );
  OAI21_X1 U16964 ( .B1(n12921), .B2(n12920), .A(n12919), .ZN(n12922) );
  INV_X1 U16965 ( .A(n12925), .ZN(n12926) );
  NAND2_X1 U16966 ( .A1(n12926), .A2(n12928), .ZN(n12930) );
  NAND2_X1 U16970 ( .A1(n12935), .A2(n13298), .ZN(n13236) );
  NAND2_X1 U16972 ( .A1(n25193), .A2(n14130), .ZN(n12939) );
  INV_X1 U16973 ( .A(n13826), .ZN(n12938) );
  AOI21_X1 U16974 ( .B1(n13896), .B2(n12939), .A(n12938), .ZN(n12940) );
  NOR2_X2 U16975 ( .A1(n12941), .A2(n12940), .ZN(n14928) );
  NOR2_X1 U16976 ( .A1(n12942), .A2(n12688), .ZN(n12943) );
  MUX2_X1 U16977 ( .A(n12944), .B(n12943), .S(n13317), .Z(n12950) );
  NOR2_X1 U16979 ( .A1(n12948), .A2(n12947), .ZN(n12949) );
  OAI211_X1 U16980 ( .C1(n13329), .C2(n12952), .A(n12951), .B(n24422), .ZN(
        n12954) );
  NAND3_X1 U16981 ( .A1(n13330), .A2(n13327), .A3(n13323), .ZN(n12953) );
  OR2_X1 U16982 ( .A1(n14208), .A2(n14205), .ZN(n12975) );
  NOR2_X1 U16983 ( .A1(n231), .A2(n12956), .ZN(n12957) );
  NOR3_X1 U16984 ( .A1(n12960), .A2(n12959), .A3(n12958), .ZN(n12961) );
  NAND3_X1 U16985 ( .A1(n13278), .A2(n13272), .A3(n12964), .ZN(n12970) );
  NAND2_X1 U16986 ( .A1(n13273), .A2(n12966), .ZN(n12967) );
  AND4_X2 U16987 ( .A1(n12970), .A2(n12969), .A3(n12968), .A4(n12967), .ZN(
        n13549) );
  NAND2_X1 U16988 ( .A1(n14206), .A2(n13549), .ZN(n12974) );
  AOI21_X1 U16989 ( .B1(n398), .B2(n25415), .A(n13345), .ZN(n12971) );
  MUX2_X1 U16990 ( .A(n12975), .B(n12974), .S(n14123), .Z(n12983) );
  NOR2_X1 U16991 ( .A1(n13357), .A2(n25584), .ZN(n12979) );
  NOR2_X1 U16993 ( .A1(n12981), .A2(n12980), .ZN(n13419) );
  INV_X1 U16994 ( .A(n14208), .ZN(n13422) );
  NAND2_X1 U16995 ( .A1(n12983), .A2(n12982), .ZN(n14466) );
  INV_X1 U16996 ( .A(n14466), .ZN(n15341) );
  XNOR2_X1 U16997 ( .A(n15341), .B(n14928), .ZN(n14677) );
  INV_X1 U16998 ( .A(n14222), .ZN(n14218) );
  NAND2_X1 U16999 ( .A1(n25080), .A2(n12993), .ZN(n13231) );
  INV_X1 U17000 ( .A(n13231), .ZN(n12996) );
  NAND2_X1 U17001 ( .A1(n12996), .A2(n12995), .ZN(n12997) );
  INV_X1 U17002 ( .A(n14219), .ZN(n13032) );
  NAND2_X1 U17003 ( .A1(n13211), .A2(n13000), .ZN(n13003) );
  NAND2_X1 U17004 ( .A1(n13001), .A2(n1335), .ZN(n13002) );
  OAI21_X1 U17005 ( .B1(n13003), .B2(n1335), .A(n13002), .ZN(n13008) );
  OAI22_X1 U17006 ( .A1(n13006), .A2(n11684), .B1(n13005), .B2(n13004), .ZN(
        n13007) );
  INV_X1 U17007 ( .A(n13830), .ZN(n14223) );
  NAND2_X1 U17008 ( .A1(n14223), .A2(n13829), .ZN(n14226) );
  NOR2_X1 U17009 ( .A1(n13011), .A2(n13014), .ZN(n13021) );
  OAI21_X1 U17010 ( .B1(n13013), .B2(n13246), .A(n25199), .ZN(n13020) );
  AOI22_X1 U17011 ( .A1(n13018), .A2(n13017), .B1(n13016), .B2(n13015), .ZN(
        n13019) );
  MUX2_X1 U17012 ( .A(n13022), .B(n14226), .S(n14225), .Z(n13036) );
  INV_X1 U17013 ( .A(n14225), .ZN(n13399) );
  NAND2_X1 U17014 ( .A1(n13399), .A2(n13829), .ZN(n13555) );
  INV_X1 U17015 ( .A(n13555), .ZN(n13034) );
  NAND2_X1 U17016 ( .A1(n13024), .A2(n13023), .ZN(n13026) );
  NOR2_X1 U17017 ( .A1(n13032), .A2(n14221), .ZN(n13033) );
  AOI22_X1 U17018 ( .A1(n13034), .A2(n14222), .B1(n14119), .B2(n13033), .ZN(
        n13035) );
  MUX2_X1 U17019 ( .A(n13039), .B(n13038), .S(n13037), .Z(n13043) );
  NOR2_X1 U17020 ( .A1(n11580), .A2(n13040), .ZN(n13042) );
  NOR2_X1 U17022 ( .A1(n13045), .A2(n13044), .ZN(n13046) );
  AOI21_X1 U17024 ( .B1(n13054), .B2(n13053), .A(n13052), .ZN(n13060) );
  NAND2_X1 U17025 ( .A1(n12526), .A2(n303), .ZN(n13058) );
  NOR2_X1 U17026 ( .A1(n13386), .A2(n24589), .ZN(n13820) );
  NAND2_X1 U17027 ( .A1(n24876), .A2(n13820), .ZN(n13085) );
  INV_X1 U17028 ( .A(n13061), .ZN(n13161) );
  INV_X1 U17029 ( .A(n13385), .ZN(n13644) );
  INV_X1 U17030 ( .A(n13067), .ZN(n13070) );
  NAND2_X1 U17031 ( .A1(n13073), .A2(n13072), .ZN(n13079) );
  NAND3_X1 U17032 ( .A1(n13644), .A2(n24589), .A3(n392), .ZN(n13084) );
  NOR2_X1 U17033 ( .A1(n13074), .A2(n24573), .ZN(n13075) );
  NOR2_X1 U17034 ( .A1(n12709), .A2(n13075), .ZN(n13081) );
  NAND2_X1 U17035 ( .A1(n24589), .A2(n13647), .ZN(n13082) );
  NAND3_X1 U17036 ( .A1(n13559), .A2(n13082), .A3(n24507), .ZN(n13083) );
  XNOR2_X1 U17037 ( .A(n14675), .B(n15210), .ZN(n15383) );
  XNOR2_X1 U17038 ( .A(n14677), .B(n15383), .ZN(n13199) );
  NAND2_X1 U17039 ( .A1(n5526), .A2(n13394), .ZN(n13571) );
  NOR3_X1 U17040 ( .A1(n13087), .A2(n14360), .A3(n13086), .ZN(n13573) );
  NOR2_X1 U17041 ( .A1(n13394), .A2(n13589), .ZN(n13090) );
  NAND2_X1 U17042 ( .A1(n13712), .A2(n13090), .ZN(n14366) );
  OAI211_X1 U17043 ( .C1(n14361), .C2(n13571), .A(n13091), .B(n14366), .ZN(
        n14345) );
  XNOR2_X1 U17044 ( .A(n14345), .B(n3155), .ZN(n13197) );
  NOR2_X1 U17045 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  NOR2_X1 U17048 ( .A1(n13109), .A2(n13108), .ZN(n13111) );
  INV_X1 U17049 ( .A(n13417), .ZN(n14099) );
  MUX2_X1 U17050 ( .A(n13117), .B(n13114), .S(n13113), .Z(n13120) );
  INV_X1 U17051 ( .A(n13115), .ZN(n13118) );
  INV_X1 U17052 ( .A(n14101), .ZN(n14213) );
  NAND2_X1 U17053 ( .A1(n406), .A2(n12349), .ZN(n13121) );
  AOI21_X1 U17054 ( .B1(n13122), .B2(n13121), .A(n13353), .ZN(n13128) );
  NAND2_X1 U17055 ( .A1(n13124), .A2(n13123), .ZN(n13126) );
  OAI21_X1 U17056 ( .B1(n13131), .B2(n13130), .A(n13129), .ZN(n13134) );
  NOR2_X1 U17057 ( .A1(n13150), .A2(n13152), .ZN(n13133) );
  NAND2_X1 U17058 ( .A1(n12433), .A2(n13136), .ZN(n13142) );
  MUX2_X1 U17060 ( .A(n13142), .B(n13141), .S(n13140), .Z(n13193) );
  NAND2_X1 U17061 ( .A1(n13144), .A2(n13143), .ZN(n13147) );
  MUX2_X1 U17062 ( .A(n13147), .B(n13146), .S(n13145), .Z(n13192) );
  NAND3_X1 U17063 ( .A1(n13150), .A2(n13149), .A3(n13148), .ZN(n13155) );
  AND3_X1 U17064 ( .A1(n13155), .A2(n13154), .A3(n13153), .ZN(n13156) );
  OAI21_X1 U17065 ( .B1(n13158), .B2(n13157), .A(n13156), .ZN(n13565) );
  NOR2_X1 U17066 ( .A1(n14106), .A2(n13565), .ZN(n14111) );
  AOI22_X1 U17067 ( .A1(n13168), .A2(n13167), .B1(n13166), .B2(n24373), .ZN(
        n13173) );
  NAND2_X1 U17068 ( .A1(n13175), .A2(n13174), .ZN(n13181) );
  NAND3_X1 U17069 ( .A1(n12459), .A2(n13176), .A3(n13178), .ZN(n13180) );
  NAND3_X1 U17070 ( .A1(n13181), .A2(n13180), .A3(n13179), .ZN(n13583) );
  OAI21_X1 U17071 ( .B1(n13566), .B2(n14105), .A(n14112), .ZN(n13182) );
  OAI21_X1 U17072 ( .B1(n14111), .B2(n14112), .A(n13182), .ZN(n13196) );
  INV_X1 U17073 ( .A(n13183), .ZN(n13186) );
  OAI21_X1 U17074 ( .B1(n13186), .B2(n13185), .A(n24640), .ZN(n13190) );
  NAND3_X1 U17076 ( .A1(n13193), .A2(n13192), .A3(n13582), .ZN(n13194) );
  OAI211_X1 U17077 ( .C1(n14112), .C2(n13582), .A(n13194), .B(n14105), .ZN(
        n13195) );
  NAND2_X1 U17078 ( .A1(n13196), .A2(n13195), .ZN(n14865) );
  XNOR2_X1 U17079 ( .A(n14976), .B(n14865), .ZN(n15028) );
  XNOR2_X1 U17080 ( .A(n13197), .B(n15028), .ZN(n13198) );
  INV_X1 U17081 ( .A(n16597), .ZN(n15890) );
  MUX2_X1 U17082 ( .A(n25209), .B(n14244), .S(n13636), .Z(n13204) );
  OAI21_X1 U17085 ( .B1(n13207), .B2(n13206), .A(n5418), .ZN(n13209) );
  NAND3_X1 U17086 ( .A1(n13213), .A2(n13212), .A3(n11360), .ZN(n13214) );
  NAND2_X1 U17087 ( .A1(n4651), .A2(n13215), .ZN(n13219) );
  NAND2_X1 U17088 ( .A1(n13217), .A2(n12767), .ZN(n13218) );
  AND2_X1 U17089 ( .A1(n13988), .A2(n13981), .ZN(n13241) );
  NAND2_X1 U17090 ( .A1(n13223), .A2(n13222), .ZN(n13226) );
  INV_X1 U17091 ( .A(n13918), .ZN(n13653) );
  NOR2_X1 U17092 ( .A1(n13230), .A2(n13229), .ZN(n13233) );
  MUX2_X2 U17093 ( .A(n13233), .B(n13232), .S(n24750), .Z(n13989) );
  NOR2_X1 U17094 ( .A1(n13653), .A2(n13989), .ZN(n13240) );
  MUX2_X1 U17095 ( .A(n13241), .B(n13240), .S(n13982), .Z(n13251) );
  OAI211_X1 U17096 ( .C1(n13246), .C2(n13245), .A(n13244), .B(n13243), .ZN(
        n13247) );
  MUX2_X1 U17097 ( .A(n13987), .B(n13988), .S(n13981), .Z(n13249) );
  INV_X1 U17098 ( .A(n13989), .ZN(n13652) );
  NOR2_X1 U17099 ( .A1(n13249), .A2(n13652), .ZN(n13250) );
  NOR2_X2 U17100 ( .A1(n13251), .A2(n13250), .ZN(n14703) );
  NAND2_X1 U17102 ( .A1(n13385), .A2(n13818), .ZN(n13822) );
  INV_X1 U17103 ( .A(n13822), .ZN(n13255) );
  INV_X1 U17104 ( .A(n13648), .ZN(n13252) );
  NAND2_X1 U17105 ( .A1(n13252), .A2(n13385), .ZN(n13254) );
  OAI21_X1 U17107 ( .B1(n13693), .B2(n24713), .A(n24715), .ZN(n13259) );
  NAND2_X1 U17108 ( .A1(n13257), .A2(n13693), .ZN(n14513) );
  NOR2_X1 U17109 ( .A1(n14436), .A2(n14439), .ZN(n14511) );
  NAND2_X1 U17110 ( .A1(n14511), .A2(n14510), .ZN(n13258) );
  OAI211_X1 U17111 ( .C1(n13260), .C2(n13259), .A(n14513), .B(n13258), .ZN(
        n13261) );
  XNOR2_X1 U17112 ( .A(n14952), .B(n13261), .ZN(n14287) );
  XNOR2_X1 U17113 ( .A(n15392), .B(n14287), .ZN(n13372) );
  XNOR2_X1 U17114 ( .A(n15062), .B(n1935), .ZN(n13370) );
  NAND2_X1 U17115 ( .A1(n5361), .A2(n13265), .ZN(n13269) );
  MUX2_X1 U17116 ( .A(n13269), .B(n13268), .S(n13267), .Z(n13270) );
  OAI21_X1 U17117 ( .B1(n5361), .B2(n13271), .A(n13270), .ZN(n14252) );
  NAND2_X1 U17118 ( .A1(n13275), .A2(n13272), .ZN(n13277) );
  INV_X1 U17119 ( .A(n14251), .ZN(n14008) );
  NAND2_X1 U17120 ( .A1(n24988), .A2(n12928), .ZN(n13280) );
  NAND2_X1 U17121 ( .A1(n13281), .A2(n13280), .ZN(n13287) );
  INV_X1 U17123 ( .A(n13923), .ZN(n14011) );
  NOR2_X1 U17124 ( .A1(n13291), .A2(n24476), .ZN(n13295) );
  NOR2_X1 U17125 ( .A1(n25466), .A2(n12594), .ZN(n13294) );
  NOR2_X2 U17126 ( .A1(n13297), .A2(n13296), .ZN(n14254) );
  NAND2_X1 U17127 ( .A1(n545), .A2(n13298), .ZN(n13300) );
  OAI22_X1 U17128 ( .A1(n4493), .A2(n13300), .B1(n24220), .B2(n545), .ZN(
        n13302) );
  NAND2_X1 U17129 ( .A1(n14009), .A2(n14251), .ZN(n13703) );
  OAI22_X1 U17130 ( .A1(n13701), .A2(n14011), .B1(n14254), .B2(n13703), .ZN(
        n13315) );
  NAND2_X1 U17131 ( .A1(n14254), .A2(n14009), .ZN(n13313) );
  INV_X1 U17132 ( .A(n14009), .ZN(n14253) );
  NOR2_X1 U17133 ( .A1(n13304), .A2(n13303), .ZN(n13312) );
  OAI211_X1 U17134 ( .C1(n13318), .C2(n13317), .A(n25499), .B(n13316), .ZN(
        n13319) );
  INV_X1 U17135 ( .A(n13319), .ZN(n13320) );
  NOR2_X1 U17136 ( .A1(n13329), .A2(n13323), .ZN(n13324) );
  NAND2_X1 U17137 ( .A1(n5311), .A2(n13324), .ZN(n13334) );
  NAND2_X1 U17138 ( .A1(n13326), .A2(n13329), .ZN(n13333) );
  NAND2_X1 U17139 ( .A1(n5139), .A2(n13327), .ZN(n13332) );
  NAND3_X1 U17140 ( .A1(n13330), .A2(n4634), .A3(n24422), .ZN(n13331) );
  AND2_X1 U17141 ( .A1(n14230), .A2(n13682), .ZN(n13356) );
  NAND2_X1 U17142 ( .A1(n13345), .A2(n25415), .ZN(n13346) );
  NOR2_X1 U17144 ( .A1(n25053), .A2(n13357), .ZN(n13362) );
  NOR2_X1 U17145 ( .A1(n24552), .A2(n13359), .ZN(n13361) );
  NAND3_X1 U17146 ( .A1(n14231), .A2(n25434), .A3(n14233), .ZN(n13368) );
  INV_X1 U17147 ( .A(n14231), .ZN(n14234) );
  NAND3_X1 U17148 ( .A1(n14234), .A2(n13995), .A3(n14233), .ZN(n13367) );
  XNOR2_X1 U17149 ( .A(n15273), .B(n15203), .ZN(n14704) );
  XNOR2_X1 U17150 ( .A(n14704), .B(n13370), .ZN(n13371) );
  XNOR2_X1 U17151 ( .A(n13371), .B(n13372), .ZN(n15821) );
  NOR2_X1 U17152 ( .A1(n24890), .A2(n24080), .ZN(n13373) );
  NAND2_X1 U17153 ( .A1(n13374), .A2(n15888), .ZN(n13375) );
  INV_X1 U17154 ( .A(n14230), .ZN(n13680) );
  NAND3_X1 U17155 ( .A1(n14234), .A2(n25435), .A3(n13680), .ZN(n13377) );
  OAI22_X1 U17156 ( .A1(n25434), .A2(n24402), .B1(n14230), .B2(n13682), .ZN(
        n13929) );
  NAND2_X1 U17157 ( .A1(n13929), .A2(n13997), .ZN(n13376) );
  NOR2_X1 U17158 ( .A1(n13667), .A2(n14005), .ZN(n13378) );
  NAND2_X1 U17159 ( .A1(n13987), .A2(n13981), .ZN(n13921) );
  AND2_X1 U17160 ( .A1(n13988), .A2(n13987), .ZN(n13655) );
  INV_X1 U17161 ( .A(n13981), .ZN(n13379) );
  XNOR2_X1 U17163 ( .A(n14377), .B(n14620), .ZN(n13384) );
  INV_X1 U17164 ( .A(n14252), .ZN(n14256) );
  NOR2_X1 U17165 ( .A1(n14254), .A2(n13924), .ZN(n13702) );
  OAI21_X1 U17166 ( .B1(n13702), .B2(n14253), .A(n14011), .ZN(n13382) );
  INV_X1 U17167 ( .A(n3089), .ZN(n22382) );
  XNOR2_X1 U17168 ( .A(n14694), .B(n22382), .ZN(n13383) );
  XNOR2_X1 U17169 ( .A(n13383), .B(n13384), .ZN(n13393) );
  NAND2_X1 U17170 ( .A1(n13385), .A2(n13647), .ZN(n13561) );
  NAND2_X1 U17171 ( .A1(n25011), .A2(n13386), .ZN(n13560) );
  AND2_X1 U17172 ( .A1(n13818), .A2(n13647), .ZN(n13387) );
  OAI21_X1 U17173 ( .B1(n13387), .B2(n13644), .A(n13646), .ZN(n13388) );
  OAI211_X1 U17174 ( .C1(n13561), .C2(n13824), .A(n13389), .B(n13388), .ZN(
        n15229) );
  NOR2_X1 U17175 ( .A1(n14510), .A2(n13693), .ZN(n13390) );
  OAI22_X1 U17176 ( .A1(n14436), .A2(n14507), .B1(n24556), .B2(n14510), .ZN(
        n13392) );
  NOR2_X1 U17177 ( .A1(n13712), .A2(n13569), .ZN(n13713) );
  NOR2_X1 U17179 ( .A1(n14361), .A2(n13394), .ZN(n13395) );
  INV_X1 U17180 ( .A(n13396), .ZN(n13397) );
  NOR2_X1 U17182 ( .A1(n13829), .A2(n14219), .ZN(n13404) );
  XNOR2_X1 U17183 ( .A(n14952), .B(n24418), .ZN(n13405) );
  NAND3_X1 U17184 ( .A1(n14127), .A2(n1331), .A3(n4844), .ZN(n13409) );
  INV_X1 U17185 ( .A(n14130), .ZN(n13894) );
  NAND3_X1 U17186 ( .A1(n13894), .A2(n13893), .A3(n14127), .ZN(n13408) );
  NAND4_X2 U17187 ( .A1(n13408), .A2(n13410), .A3(n13409), .A4(n13407), .ZN(
        n15396) );
  XNOR2_X1 U17188 ( .A(n15396), .B(n1792), .ZN(n13416) );
  NAND2_X1 U17189 ( .A1(n14106), .A2(n13565), .ZN(n13413) );
  NAND2_X1 U17190 ( .A1(n14107), .A2(n4868), .ZN(n13411) );
  MUX2_X1 U17191 ( .A(n13413), .B(n13411), .S(n5333), .Z(n13415) );
  INV_X1 U17192 ( .A(n13565), .ZN(n13584) );
  AOI21_X1 U17193 ( .B1(n13584), .B2(n14108), .A(n14105), .ZN(n13412) );
  NAND2_X1 U17194 ( .A1(n13413), .A2(n13412), .ZN(n13414) );
  NAND2_X1 U17195 ( .A1(n13415), .A2(n13414), .ZN(n13873) );
  INV_X1 U17196 ( .A(n13873), .ZN(n15199) );
  XNOR2_X1 U17197 ( .A(n13416), .B(n15199), .ZN(n13423) );
  OAI21_X1 U17198 ( .B1(n13417), .B2(n14211), .A(n14213), .ZN(n13418) );
  NOR2_X1 U17199 ( .A1(n14124), .A2(n13419), .ZN(n13420) );
  NAND2_X1 U17200 ( .A1(n13421), .A2(n13420), .ZN(n13548) );
  XNOR2_X1 U17201 ( .A(n14834), .B(n15463), .ZN(n15270) );
  XNOR2_X1 U17202 ( .A(n13423), .B(n15270), .ZN(n13424) );
  INV_X1 U17203 ( .A(n15915), .ZN(n16336) );
  INV_X1 U17204 ( .A(n13845), .ZN(n13844) );
  NOR2_X1 U17205 ( .A1(n14063), .A2(n13844), .ZN(n13425) );
  NAND2_X1 U17206 ( .A1(n13426), .A2(n13425), .ZN(n13431) );
  NAND2_X1 U17207 ( .A1(n13427), .A2(n13845), .ZN(n14069) );
  NOR2_X1 U17208 ( .A1(n13843), .A2(n13845), .ZN(n13428) );
  NAND2_X1 U17209 ( .A1(n14064), .A2(n13428), .ZN(n13429) );
  NAND2_X1 U17210 ( .A1(n13566), .A2(n14108), .ZN(n13436) );
  OAI21_X1 U17211 ( .B1(n5333), .B2(n13566), .A(n13584), .ZN(n13432) );
  NOR2_X1 U17213 ( .A1(n5333), .A2(n14105), .ZN(n13433) );
  NAND2_X1 U17214 ( .A1(n13433), .A2(n13566), .ZN(n13434) );
  INV_X1 U17216 ( .A(n13552), .ZN(n14216) );
  NAND2_X1 U17217 ( .A1(n14216), .A2(n24376), .ZN(n13440) );
  OAI21_X1 U17218 ( .B1(n13417), .B2(n13552), .A(n25445), .ZN(n13438) );
  XNOR2_X1 U17219 ( .A(n15183), .B(n1870), .ZN(n13441) );
  INV_X1 U17220 ( .A(n13982), .ZN(n13922) );
  OAI21_X1 U17221 ( .B1(n13918), .B2(n13989), .A(n13922), .ZN(n13443) );
  INV_X1 U17222 ( .A(n13988), .ZN(n13656) );
  INV_X1 U17223 ( .A(n13917), .ZN(n13986) );
  OAI21_X1 U17224 ( .B1(n13656), .B2(n13981), .A(n13986), .ZN(n13442) );
  NAND3_X1 U17228 ( .A1(n24572), .A2(n24958), .A3(n14852), .ZN(n13446) );
  NAND3_X1 U17229 ( .A1(n14849), .A2(n14850), .A3(n14852), .ZN(n13445) );
  NOR2_X1 U17231 ( .A1(n14271), .A2(n13840), .ZN(n13761) );
  NOR3_X1 U17233 ( .A1(n24368), .A2(n397), .A3(n14268), .ZN(n13449) );
  AOI21_X1 U17234 ( .B1(n3947), .B2(n16336), .A(n290), .ZN(n13547) );
  MUX2_X1 U17241 ( .A(n13459), .B(n13458), .S(n14307), .Z(n13462) );
  XNOR2_X1 U17242 ( .A(n14477), .B(n14676), .ZN(n15290) );
  INV_X1 U17243 ( .A(n14289), .ZN(n14293) );
  NAND3_X1 U17244 ( .A1(n14293), .A2(n13909), .A3(n394), .ZN(n13465) );
  AOI21_X1 U17245 ( .B1(n13909), .B2(n24974), .A(n14294), .ZN(n13463) );
  XNOR2_X1 U17246 ( .A(n14345), .B(n14468), .ZN(n14933) );
  XNOR2_X1 U17247 ( .A(n15290), .B(n14933), .ZN(n13476) );
  NAND2_X1 U17248 ( .A1(n14172), .A2(n14168), .ZN(n13527) );
  NOR2_X1 U17249 ( .A1(n13775), .A2(n13954), .ZN(n13716) );
  AOI22_X1 U17250 ( .A1(n13716), .A2(n14156), .B1(n13467), .B2(n13954), .ZN(
        n13468) );
  OAI21_X2 U17251 ( .B1(n14160), .B2(n13469), .A(n13468), .ZN(n15386) );
  XNOR2_X1 U17252 ( .A(n14979), .B(n15386), .ZN(n13474) );
  AOI22_X1 U17253 ( .A1(n13969), .A2(n13596), .B1(n13470), .B2(n13968), .ZN(
        n13471) );
  INV_X1 U17254 ( .A(n1726), .ZN(n13472) );
  XNOR2_X1 U17255 ( .A(n15488), .B(n13472), .ZN(n13473) );
  XNOR2_X1 U17256 ( .A(n13474), .B(n13473), .ZN(n13475) );
  AND2_X1 U17258 ( .A1(n13785), .A2(n14142), .ZN(n13477) );
  AND2_X1 U17259 ( .A1(n14144), .A2(n14199), .ZN(n13481) );
  INV_X1 U17261 ( .A(n13804), .ZN(n13480) );
  NOR2_X1 U17262 ( .A1(n14200), .A2(n3888), .ZN(n13479) );
  NOR2_X1 U17264 ( .A1(n13792), .A2(n13795), .ZN(n13482) );
  INV_X1 U17265 ( .A(n14178), .ZN(n13580) );
  OAI21_X1 U17266 ( .B1(n13482), .B2(n13580), .A(n14182), .ZN(n13483) );
  XNOR2_X1 U17267 ( .A(n14900), .B(n15190), .ZN(n14940) );
  INV_X1 U17268 ( .A(n14078), .ZN(n14073) );
  OAI21_X1 U17269 ( .B1(n13491), .B2(n13628), .A(n13629), .ZN(n13492) );
  XNOR2_X1 U17270 ( .A(n15191), .B(n15514), .ZN(n13497) );
  OAI211_X1 U17271 ( .C1(n14439), .C2(n13974), .A(n24556), .B(n24713), .ZN(
        n13495) );
  NAND3_X1 U17272 ( .A1(n14440), .A2(n13693), .A3(n13975), .ZN(n13494) );
  AND3_X1 U17273 ( .A1(n13978), .A2(n13495), .A3(n13494), .ZN(n14996) );
  INV_X1 U17274 ( .A(n14996), .ZN(n14549) );
  XNOR2_X1 U17275 ( .A(n14549), .B(n2772), .ZN(n13496) );
  XNOR2_X1 U17276 ( .A(n13497), .B(n13496), .ZN(n13498) );
  NOR2_X1 U17277 ( .A1(n16332), .A2(n25092), .ZN(n13545) );
  INV_X1 U17278 ( .A(n14333), .ZN(n13593) );
  INV_X1 U17279 ( .A(n25196), .ZN(n13501) );
  INV_X1 U17280 ( .A(n13504), .ZN(n13505) );
  OAI211_X1 U17281 ( .C1(n25197), .C2(n14025), .A(n14334), .B(n13508), .ZN(
        n13510) );
  NAND3_X1 U17282 ( .A1(n14336), .A2(n13593), .A3(n14339), .ZN(n13509) );
  XNOR2_X1 U17283 ( .A(n14880), .B(n14815), .ZN(n15281) );
  NOR2_X1 U17284 ( .A1(n13807), .A2(n14149), .ZN(n13512) );
  OAI21_X1 U17285 ( .B1(n13515), .B2(n14153), .A(n13514), .ZN(n13516) );
  NOR2_X1 U17286 ( .A1(n13614), .A2(n1355), .ZN(n13520) );
  NAND2_X1 U17287 ( .A1(n13612), .A2(n13610), .ZN(n13519) );
  NOR2_X1 U17289 ( .A1(n14325), .A2(n14041), .ZN(n13590) );
  OAI21_X1 U17290 ( .B1(n14172), .B2(n13741), .A(n13526), .ZN(n13531) );
  INV_X1 U17291 ( .A(n13527), .ZN(n13530) );
  NAND3_X1 U17292 ( .A1(n13741), .A2(n14164), .A3(n13744), .ZN(n13528) );
  OAI211_X1 U17293 ( .C1(n13531), .C2(n13530), .A(n13529), .B(n13528), .ZN(
        n13532) );
  NAND4_X1 U17294 ( .A1(n13538), .A2(n13537), .A3(n13536), .A4(n13535), .ZN(
        n13539) );
  AOI21_X1 U17295 ( .B1(n13540), .B2(n13539), .A(n14088), .ZN(n13541) );
  XNOR2_X1 U17296 ( .A(n15178), .B(n4711), .ZN(n13543) );
  XNOR2_X1 U17297 ( .A(n14964), .B(n13543), .ZN(n13544) );
  NOR2_X1 U17298 ( .A1(n16331), .A2(n15667), .ZN(n16337) );
  OAI21_X1 U17299 ( .B1(n13545), .B2(n16337), .A(n15915), .ZN(n13546) );
  INV_X1 U17300 ( .A(n13813), .ZN(n13550) );
  NOR2_X1 U17302 ( .A1(n14101), .A2(n4894), .ZN(n13554) );
  OAI21_X1 U17303 ( .B1(n14217), .B2(n13554), .A(n13553), .ZN(n15194) );
  XNOR2_X1 U17304 ( .A(n14993), .B(n15194), .ZN(n15513) );
  OAI211_X1 U17305 ( .C1(n14223), .C2(n13829), .A(n14218), .B(n14219), .ZN(
        n13557) );
  XNOR2_X1 U17307 ( .A(n15444), .B(n173), .ZN(n13558) );
  XNOR2_X1 U17308 ( .A(n15513), .B(n13558), .ZN(n13577) );
  INV_X1 U17309 ( .A(n13561), .ZN(n13564) );
  NAND2_X1 U17310 ( .A1(n13824), .A2(n24589), .ZN(n13563) );
  OAI211_X1 U17311 ( .C1(n13561), .C2(n25011), .A(n13560), .B(n13559), .ZN(
        n13562) );
  INV_X1 U17313 ( .A(n14106), .ZN(n14109) );
  INV_X1 U17314 ( .A(n13581), .ZN(n13567) );
  XNOR2_X1 U17315 ( .A(n14667), .B(n15244), .ZN(n14770) );
  AND2_X1 U17316 ( .A1(n14132), .A2(n13895), .ZN(n13575) );
  NAND3_X1 U17317 ( .A1(n14127), .A2(n14126), .A3(n14132), .ZN(n13574) );
  XNOR2_X1 U17318 ( .A(n14488), .B(n15034), .ZN(n14825) );
  XNOR2_X1 U17319 ( .A(n14825), .B(n14770), .ZN(n13576) );
  INV_X1 U17320 ( .A(n16200), .ZN(n16403) );
  NOR2_X1 U17321 ( .A1(n14178), .A2(n13578), .ZN(n13793) );
  XNOR2_X1 U17322 ( .A(n15165), .B(n729), .ZN(n13585) );
  INV_X1 U17323 ( .A(n14361), .ZN(n13586) );
  INV_X1 U17324 ( .A(n13712), .ZN(n14364) );
  NAND3_X1 U17325 ( .A1(n24995), .A2(n14364), .A3(n3701), .ZN(n13588) );
  NOR2_X1 U17326 ( .A1(n13590), .A2(n14328), .ZN(n13591) );
  INV_X1 U17327 ( .A(n25413), .ZN(n13592) );
  XNOR2_X1 U17328 ( .A(n15230), .B(n13592), .ZN(n14763) );
  INV_X1 U17329 ( .A(n14336), .ZN(n14026) );
  INV_X1 U17330 ( .A(n13877), .ZN(n14340) );
  OAI21_X2 U17331 ( .B1(n13595), .B2(n14026), .A(n13594), .ZN(n15051) );
  XNOR2_X1 U17333 ( .A(n15051), .B(n15430), .ZN(n13605) );
  XNOR2_X1 U17335 ( .A(n13605), .B(n25431), .ZN(n14633) );
  NAND2_X1 U17337 ( .A1(n14017), .A2(n14089), .ZN(n13608) );
  NAND2_X1 U17338 ( .A1(n14054), .A2(n14049), .ZN(n13613) );
  OAI22_X1 U17339 ( .A1(n13614), .A2(n13613), .B1(n14054), .B2(n13612), .ZN(
        n13615) );
  XNOR2_X1 U17340 ( .A(n14755), .B(n15487), .ZN(n15241) );
  NOR2_X1 U17341 ( .A1(n14059), .A2(n14852), .ZN(n13617) );
  NAND2_X1 U17342 ( .A1(n14267), .A2(n14269), .ZN(n13621) );
  OR2_X1 U17343 ( .A1(n13840), .A2(n14269), .ZN(n13620) );
  AOI21_X1 U17345 ( .B1(n13621), .B2(n13620), .A(n123), .ZN(n13625) );
  OAI21_X1 U17346 ( .B1(n13839), .B2(n13623), .A(n13622), .ZN(n13624) );
  INV_X1 U17348 ( .A(n14678), .ZN(n14756) );
  XNOR2_X1 U17349 ( .A(n14756), .B(n14789), .ZN(n13626) );
  XNOR2_X1 U17350 ( .A(n13626), .B(n15241), .ZN(n13642) );
  OAI211_X1 U17351 ( .C1(n14076), .C2(n14078), .A(n13629), .B(n14074), .ZN(
        n13630) );
  XNOR2_X1 U17352 ( .A(n15486), .B(n15436), .ZN(n14649) );
  NAND2_X1 U17353 ( .A1(n14240), .A2(n14244), .ZN(n13634) );
  OAI211_X1 U17354 ( .C1(n13633), .C2(n14244), .A(n4116), .B(n13634), .ZN(
        n13638) );
  XNOR2_X1 U17358 ( .A(n14792), .B(n1865), .ZN(n13640) );
  XNOR2_X1 U17359 ( .A(n14649), .B(n13640), .ZN(n13641) );
  NOR2_X1 U17360 ( .A1(n13989), .A2(n13656), .ZN(n13654) );
  INV_X1 U17361 ( .A(n13655), .ZN(n13658) );
  NAND2_X1 U17362 ( .A1(n13656), .A2(n13981), .ZN(n13657) );
  XNOR2_X1 U17363 ( .A(n14644), .B(n14816), .ZN(n13691) );
  INV_X1 U17364 ( .A(n13659), .ZN(n13666) );
  AOI21_X1 U17365 ( .B1(n13661), .B2(n13662), .A(n13660), .ZN(n13665) );
  NAND2_X1 U17366 ( .A1(n13663), .A2(n13662), .ZN(n13664) );
  INV_X1 U17367 ( .A(n13668), .ZN(n13673) );
  INV_X1 U17368 ( .A(n13669), .ZN(n13672) );
  INV_X1 U17369 ( .A(n13670), .ZN(n13671) );
  NAND3_X1 U17370 ( .A1(n13673), .A2(n13672), .A3(n13671), .ZN(n13674) );
  NAND2_X1 U17371 ( .A1(n14003), .A2(n13676), .ZN(n13677) );
  OAI21_X2 U17372 ( .B1(n13679), .B2(n13678), .A(n13677), .ZN(n15175) );
  NAND2_X1 U17373 ( .A1(n13680), .A2(n13683), .ZN(n13688) );
  NAND2_X1 U17374 ( .A1(n13680), .A2(n13681), .ZN(n13687) );
  NOR2_X1 U17375 ( .A1(n13682), .A2(n13681), .ZN(n13685) );
  INV_X1 U17376 ( .A(n13683), .ZN(n13684) );
  AOI21_X1 U17377 ( .B1(n13685), .B2(n13684), .A(n24402), .ZN(n13686) );
  NAND3_X1 U17378 ( .A1(n13688), .A2(n13687), .A3(n13686), .ZN(n13690) );
  NOR2_X1 U17379 ( .A1(n24556), .A2(n14439), .ZN(n13692) );
  MUX2_X1 U17380 ( .A(n14511), .B(n13692), .S(n14510), .Z(n13696) );
  OAI21_X1 U17383 ( .B1(n14440), .B2(n14509), .A(n14434), .ZN(n13695) );
  NOR2_X1 U17384 ( .A1(n13696), .A2(n13695), .ZN(n13700) );
  XNOR2_X1 U17387 ( .A(n14690), .B(n13700), .ZN(n14781) );
  INV_X1 U17388 ( .A(n14254), .ZN(n14250) );
  NAND3_X1 U17389 ( .A1(n14250), .A2(n14008), .A3(n13923), .ZN(n13706) );
  NAND2_X1 U17390 ( .A1(n13702), .A2(n14251), .ZN(n13705) );
  XNOR2_X1 U17392 ( .A(n24938), .B(n20046), .ZN(n13708) );
  XNOR2_X1 U17393 ( .A(n14781), .B(n13708), .ZN(n13709) );
  AND3_X1 U17394 ( .A1(n14361), .A2(n13712), .A3(n14360), .ZN(n13714) );
  NOR2_X1 U17395 ( .A1(n13714), .A2(n13713), .ZN(n13715) );
  INV_X1 U17396 ( .A(n13716), .ZN(n13955) );
  NAND2_X1 U17397 ( .A1(n14156), .A2(n5080), .ZN(n13717) );
  NAND2_X1 U17398 ( .A1(n13955), .A2(n13717), .ZN(n13721) );
  NAND2_X1 U17399 ( .A1(n13718), .A2(n13776), .ZN(n13720) );
  XNOR2_X1 U17400 ( .A(n14671), .B(n15253), .ZN(n14749) );
  INV_X1 U17401 ( .A(n24973), .ZN(n14292) );
  NAND2_X1 U17402 ( .A1(n14289), .A2(n13907), .ZN(n13723) );
  XNOR2_X1 U17403 ( .A(n15452), .B(n15074), .ZN(n14653) );
  XNOR2_X1 U17404 ( .A(n14653), .B(n14749), .ZN(n13738) );
  AOI21_X1 U17405 ( .B1(n13892), .B2(n14306), .A(n13947), .ZN(n13729) );
  INV_X1 U17406 ( .A(n13892), .ZN(n13728) );
  OAI21_X1 U17407 ( .B1(n13959), .B2(n13900), .A(n13956), .ZN(n13732) );
  NAND2_X1 U17408 ( .A1(n14311), .A2(n14307), .ZN(n13730) );
  NAND2_X1 U17409 ( .A1(n13900), .A2(n4525), .ZN(n14314) );
  OAI21_X1 U17410 ( .B1(n13730), .B2(n13958), .A(n14314), .ZN(n13731) );
  INV_X1 U17411 ( .A(n14168), .ZN(n13743) );
  XNOR2_X1 U17412 ( .A(n14800), .B(n1724), .ZN(n13736) );
  XNOR2_X1 U17413 ( .A(n14389), .B(n13736), .ZN(n13737) );
  INV_X1 U17414 ( .A(n13785), .ZN(n14191) );
  MUX2_X1 U17415 ( .A(n14189), .B(n14141), .S(n14190), .Z(n13739) );
  NOR2_X1 U17416 ( .A1(n25560), .A2(n13739), .ZN(n13740) );
  OAI21_X1 U17417 ( .B1(n14164), .B2(n13741), .A(n14172), .ZN(n13749) );
  NOR2_X1 U17418 ( .A1(n14167), .A2(n13742), .ZN(n13748) );
  NOR2_X1 U17419 ( .A1(n13744), .A2(n13743), .ZN(n13746) );
  AOI22_X1 U17420 ( .A1(n14166), .A2(n13746), .B1(n13745), .B2(n14167), .ZN(
        n13747) );
  XNOR2_X1 U17421 ( .A(n15318), .B(n15219), .ZN(n13756) );
  OR2_X1 U17422 ( .A1(n14035), .A2(n14149), .ZN(n14033) );
  OAI211_X1 U17423 ( .C1(n297), .C2(n14034), .A(n14033), .B(n14153), .ZN(
        n13751) );
  NOR2_X1 U17424 ( .A1(n3889), .A2(n3888), .ZN(n14947) );
  NAND2_X1 U17425 ( .A1(n14947), .A2(n14946), .ZN(n13755) );
  NOR2_X1 U17426 ( .A1(n2570), .A2(n25458), .ZN(n13753) );
  NOR2_X1 U17427 ( .A1(n2684), .A2(n12629), .ZN(n13752) );
  OAI21_X1 U17428 ( .B1(n13753), .B2(n13752), .A(n14198), .ZN(n13754) );
  NAND3_X1 U17429 ( .A1(n13755), .A2(n13754), .A3(n14949), .ZN(n14383) );
  XNOR2_X1 U17430 ( .A(n15464), .B(n14383), .ZN(n14638) );
  XNOR2_X1 U17431 ( .A(n13756), .B(n14638), .ZN(n13784) );
  INV_X1 U17432 ( .A(n13757), .ZN(n13758) );
  NOR3_X1 U17433 ( .A1(n397), .A2(n13759), .A3(n13758), .ZN(n13760) );
  NOR2_X1 U17434 ( .A1(n13839), .A2(n13760), .ZN(n13763) );
  INV_X1 U17435 ( .A(n13761), .ZN(n13762) );
  NAND2_X1 U17436 ( .A1(n13763), .A2(n13762), .ZN(n13767) );
  NOR2_X1 U17437 ( .A1(n14271), .A2(n14274), .ZN(n13765) );
  AOI22_X1 U17438 ( .A1(n13765), .A2(n24368), .B1(n13839), .B2(n13764), .ZN(
        n13766) );
  NAND2_X1 U17439 ( .A1(n13767), .A2(n13766), .ZN(n14516) );
  NOR2_X1 U17440 ( .A1(n14178), .A2(n14182), .ZN(n13770) );
  NOR2_X1 U17441 ( .A1(n13796), .A2(n13792), .ZN(n13768) );
  AOI22_X1 U17442 ( .A1(n13770), .A2(n13769), .B1(n13768), .B2(n14178), .ZN(
        n13772) );
  XNOR2_X1 U17443 ( .A(n14775), .B(n14516), .ZN(n13782) );
  NAND2_X1 U17444 ( .A1(n13775), .A2(n13954), .ZN(n13779) );
  INV_X1 U17445 ( .A(n13776), .ZN(n13777) );
  NAND2_X1 U17446 ( .A1(n13777), .A2(n5080), .ZN(n13778) );
  XNOR2_X1 U17447 ( .A(n25436), .B(n1831), .ZN(n13781) );
  XNOR2_X1 U17448 ( .A(n13782), .B(n13781), .ZN(n13783) );
  XNOR2_X1 U17449 ( .A(n13784), .B(n13783), .ZN(n16202) );
  INV_X1 U17450 ( .A(n16202), .ZN(n16406) );
  NOR2_X1 U17451 ( .A1(n13788), .A2(n14141), .ZN(n13787) );
  NAND2_X1 U17453 ( .A1(n13789), .A2(n13788), .ZN(n13790) );
  NOR2_X1 U17454 ( .A1(n14178), .A2(n24949), .ZN(n13794) );
  MUX2_X1 U17455 ( .A(n13794), .B(n13793), .S(n13792), .Z(n13799) );
  OAI22_X1 U17456 ( .A1(n13797), .A2(n14179), .B1(n14182), .B2(n5755), .ZN(
        n13798) );
  XNOR2_X1 U17457 ( .A(n15484), .B(n1359), .ZN(n13800) );
  XNOR2_X1 U17458 ( .A(n14979), .B(n14678), .ZN(n14534) );
  XNOR2_X1 U17459 ( .A(n13800), .B(n14534), .ZN(n13810) );
  XNOR2_X1 U17460 ( .A(n15386), .B(n921), .ZN(n13808) );
  NAND3_X1 U17461 ( .A1(n14945), .A2(n14199), .A3(n25458), .ZN(n13803) );
  XNOR2_X1 U17462 ( .A(n14977), .B(n25013), .ZN(n14608) );
  XNOR2_X1 U17463 ( .A(n13808), .B(n14608), .ZN(n13809) );
  XNOR2_X1 U17464 ( .A(n13810), .B(n13809), .ZN(n15638) );
  INV_X1 U17465 ( .A(n15638), .ZN(n15973) );
  NOR2_X1 U17466 ( .A1(n3341), .A2(n14205), .ZN(n13812) );
  OAI21_X1 U17467 ( .B1(n13813), .B2(n13812), .A(n13811), .ZN(n13817) );
  AOI21_X1 U17468 ( .B1(n13815), .B2(n14209), .A(n13814), .ZN(n13816) );
  XNOR2_X1 U17469 ( .A(n14671), .B(n15094), .ZN(n13825) );
  NOR2_X1 U17470 ( .A1(n13819), .A2(n13818), .ZN(n13821) );
  OAI21_X1 U17471 ( .B1(n13821), .B2(n13820), .A(n13824), .ZN(n13823) );
  OAI211_X1 U17472 ( .C1(n13824), .C2(n13648), .A(n13823), .B(n13822), .ZN(
        n14737) );
  XNOR2_X1 U17473 ( .A(n14737), .B(n14654), .ZN(n14986) );
  XNOR2_X1 U17474 ( .A(n14986), .B(n13825), .ZN(n13836) );
  NOR2_X1 U17475 ( .A1(n13895), .A2(n1331), .ZN(n13827) );
  XNOR2_X1 U17476 ( .A(n15507), .B(n15183), .ZN(n15368) );
  NOR2_X1 U17477 ( .A1(n13830), .A2(n14219), .ZN(n13828) );
  AND2_X1 U17478 ( .A1(n13830), .A2(n14225), .ZN(n14116) );
  NAND3_X1 U17479 ( .A1(n14222), .A2(n13830), .A3(n14219), .ZN(n13832) );
  OAI211_X2 U17480 ( .C1(n13833), .C2(n14119), .A(n13832), .B(n13831), .ZN(
        n15359) );
  XNOR2_X1 U17481 ( .A(n15359), .B(n2033), .ZN(n13834) );
  XNOR2_X1 U17482 ( .A(n15368), .B(n13834), .ZN(n13835) );
  INV_X1 U17483 ( .A(n16186), .ZN(n16398) );
  NOR2_X1 U17484 ( .A1(n15973), .A2(n16398), .ZN(n13916) );
  NOR2_X1 U17485 ( .A1(n13839), .A2(n14268), .ZN(n13838) );
  AOI21_X1 U17486 ( .B1(n13840), .B2(n13839), .A(n13838), .ZN(n13841) );
  MUX2_X1 U17487 ( .A(n13842), .B(n13841), .S(n14274), .Z(n15002) );
  XNOR2_X1 U17488 ( .A(n1351), .B(n15002), .ZN(n13850) );
  NOR2_X1 U17489 ( .A1(n13627), .A2(n14063), .ZN(n13846) );
  NAND2_X1 U17490 ( .A1(n14069), .A2(n13846), .ZN(n13848) );
  AND2_X1 U17491 ( .A1(n13847), .A2(n14063), .ZN(n14065) );
  XNOR2_X1 U17493 ( .A(n14611), .B(n15178), .ZN(n14965) );
  XNOR2_X1 U17494 ( .A(n14965), .B(n13850), .ZN(n13862) );
  OAI21_X1 U17495 ( .B1(n14075), .B2(n13852), .A(n13851), .ZN(n13857) );
  OAI21_X1 U17496 ( .B1(n13854), .B2(n13853), .A(n12704), .ZN(n13856) );
  AOI21_X1 U17497 ( .B1(n14074), .B2(n14079), .A(n14078), .ZN(n13855) );
  AOI21_X1 U17498 ( .B1(n24572), .B2(n14849), .A(n14852), .ZN(n13858) );
  OAI21_X1 U17499 ( .B1(n24572), .B2(n14416), .A(n13858), .ZN(n13859) );
  XNOR2_X1 U17500 ( .A(n24956), .B(n14558), .ZN(n14614) );
  XNOR2_X1 U17501 ( .A(n14690), .B(n1856), .ZN(n13860) );
  XNOR2_X1 U17502 ( .A(n14614), .B(n13860), .ZN(n13861) );
  XNOR2_X1 U17503 ( .A(n13862), .B(n13861), .ZN(n13940) );
  INV_X1 U17504 ( .A(n13940), .ZN(n16188) );
  NOR2_X1 U17505 ( .A1(n14325), .A2(n14328), .ZN(n14043) );
  OAI21_X1 U17506 ( .B1(n14043), .B2(n13864), .A(n13863), .ZN(n13866) );
  OAI21_X1 U17507 ( .B1(n13864), .B2(n14324), .A(n14328), .ZN(n13865) );
  XNOR2_X1 U17508 ( .A(n13867), .B(n14775), .ZN(n13874) );
  OR2_X1 U17509 ( .A1(n14319), .A2(n13868), .ZN(n13870) );
  NAND3_X1 U17510 ( .A1(n14321), .A2(n13868), .A3(n14320), .ZN(n13869) );
  OAI21_X1 U17511 ( .B1(n14317), .B2(n13870), .A(n13869), .ZN(n13872) );
  XNOR2_X1 U17512 ( .A(n15120), .B(n13873), .ZN(n14955) );
  XNOR2_X1 U17513 ( .A(n13874), .B(n14955), .ZN(n13887) );
  NAND2_X1 U17514 ( .A1(n14340), .A2(n14335), .ZN(n13876) );
  NAND2_X1 U17515 ( .A1(n13877), .A2(n25197), .ZN(n13875) );
  AOI21_X1 U17516 ( .B1(n13876), .B2(n13875), .A(n14333), .ZN(n13882) );
  NOR2_X1 U17517 ( .A1(n25196), .A2(n14339), .ZN(n14028) );
  NAND2_X1 U17518 ( .A1(n13878), .A2(n14336), .ZN(n13879) );
  NAND2_X1 U17519 ( .A1(n13880), .A2(n13879), .ZN(n13881) );
  XNOR2_X1 U17520 ( .A(n25443), .B(n15393), .ZN(n14593) );
  XNOR2_X1 U17521 ( .A(n15019), .B(n14593), .ZN(n13886) );
  XNOR2_X1 U17522 ( .A(n13887), .B(n13886), .ZN(n15637) );
  INV_X1 U17523 ( .A(n15637), .ZN(n16399) );
  NOR2_X1 U17524 ( .A1(n16188), .A2(n16399), .ZN(n13915) );
  OAI21_X1 U17525 ( .B1(n13890), .B2(n3966), .A(n1527), .ZN(n13891) );
  NAND2_X1 U17526 ( .A1(n13894), .A2(n4133), .ZN(n13898) );
  XNOR2_X1 U17528 ( .A(n15326), .B(n24423), .ZN(n14619) );
  AOI21_X1 U17529 ( .B1(n13901), .B2(n13900), .A(n13903), .ZN(n13905) );
  XNOR2_X1 U17531 ( .A(n14973), .B(n14619), .ZN(n13914) );
  XNOR2_X1 U17532 ( .A(n25413), .B(n15229), .ZN(n14543) );
  AOI21_X1 U17533 ( .B1(n24974), .B2(n13907), .A(n14293), .ZN(n13911) );
  INV_X1 U17534 ( .A(n14294), .ZN(n14291) );
  NOR2_X1 U17535 ( .A1(n14294), .A2(n13909), .ZN(n13948) );
  OAI21_X1 U17536 ( .B1(n13911), .B2(n14291), .A(n13910), .ZN(n14719) );
  XNOR2_X1 U17537 ( .A(n14719), .B(n2236), .ZN(n13912) );
  XNOR2_X1 U17538 ( .A(n14543), .B(n13912), .ZN(n13913) );
  MUX2_X1 U17539 ( .A(n13916), .B(n13915), .S(n3630), .Z(n13943) );
  NAND2_X1 U17540 ( .A1(n1846), .A2(n16186), .ZN(n15639) );
  INV_X1 U17541 ( .A(n13985), .ZN(n13920) );
  OAI21_X1 U17542 ( .B1(n13918), .B2(n13922), .A(n13917), .ZN(n13919) );
  NOR2_X1 U17543 ( .A1(n14008), .A2(n13923), .ZN(n14255) );
  NOR2_X1 U17544 ( .A1(n14252), .A2(n14251), .ZN(n13926) );
  NAND2_X1 U17545 ( .A1(n14254), .A2(n13924), .ZN(n13925) );
  OAI22_X1 U17546 ( .A1(n13927), .A2(n14255), .B1(n13926), .B2(n13925), .ZN(
        n15515) );
  XNOR2_X1 U17547 ( .A(n15515), .B(n15350), .ZN(n14600) );
  XNOR2_X1 U17548 ( .A(n14600), .B(n13928), .ZN(n13939) );
  NOR2_X1 U17549 ( .A1(n13995), .A2(n13997), .ZN(n13930) );
  XNOR2_X1 U17550 ( .A(n15112), .B(n14996), .ZN(n13937) );
  NAND3_X1 U17551 ( .A1(n13931), .A2(n13935), .A3(n14244), .ZN(n13934) );
  NOR2_X1 U17552 ( .A1(n25208), .A2(n14244), .ZN(n13933) );
  XNOR2_X1 U17553 ( .A(n14997), .B(n1746), .ZN(n13936) );
  XNOR2_X1 U17554 ( .A(n13937), .B(n13936), .ZN(n13938) );
  AOI21_X1 U17556 ( .B1(n15639), .B2(n13941), .A(n15971), .ZN(n13942) );
  AOI21_X1 U17557 ( .B1(n24588), .B2(n24710), .A(n14306), .ZN(n13946) );
  INV_X1 U17558 ( .A(n13948), .ZN(n13950) );
  NAND2_X1 U17559 ( .A1(n13953), .A2(n14158), .ZN(n13952) );
  XNOR2_X1 U17560 ( .A(n15111), .B(n14579), .ZN(n14429) );
  XNOR2_X1 U17561 ( .A(n14429), .B(n14715), .ZN(n13973) );
  NAND2_X1 U17562 ( .A1(n13957), .A2(n13956), .ZN(n13961) );
  OAI211_X1 U17563 ( .C1(n14311), .C2(n14307), .A(n13959), .B(n13958), .ZN(
        n13960) );
  XNOR2_X1 U17565 ( .A(n15109), .B(n25008), .ZN(n13971) );
  NAND3_X1 U17566 ( .A1(n13968), .A2(n13966), .A3(n13965), .ZN(n13967) );
  XNOR2_X1 U17567 ( .A(n15153), .B(n1754), .ZN(n13970) );
  XNOR2_X1 U17568 ( .A(n13971), .B(n13970), .ZN(n13972) );
  XNOR2_X1 U17573 ( .A(n15088), .B(n15210), .ZN(n14423) );
  INV_X1 U17574 ( .A(n14423), .ZN(n13999) );
  NOR2_X1 U17575 ( .A1(n13988), .A2(n13981), .ZN(n13983) );
  NAND2_X1 U17576 ( .A1(n13986), .A2(n13985), .ZN(n13992) );
  XNOR2_X1 U17577 ( .A(n14788), .B(n15483), .ZN(n14532) );
  XNOR2_X1 U17578 ( .A(n13999), .B(n14532), .ZN(n14016) );
  AOI21_X1 U17579 ( .B1(n299), .B2(n14000), .A(n14003), .ZN(n14001) );
  NOR2_X1 U17580 ( .A1(n14009), .A2(n14251), .ZN(n14010) );
  XNOR2_X1 U17581 ( .A(n14980), .B(n24502), .ZN(n14014) );
  XNOR2_X1 U17582 ( .A(n14792), .B(n1924), .ZN(n14013) );
  XNOR2_X1 U17583 ( .A(n14014), .B(n14013), .ZN(n14015) );
  XNOR2_X1 U17584 ( .A(n14015), .B(n14016), .ZN(n15640) );
  NAND2_X1 U17585 ( .A1(n14022), .A2(n14085), .ZN(n14092) );
  NOR2_X1 U17586 ( .A1(n14018), .A2(n14022), .ZN(n14019) );
  AOI21_X1 U17587 ( .B1(n14020), .B2(n14092), .A(n14019), .ZN(n14024) );
  NOR3_X1 U17588 ( .A1(n14022), .A2(n14089), .A3(n14021), .ZN(n14023) );
  XNOR2_X1 U17589 ( .A(n15184), .B(n15097), .ZN(n14414) );
  AND2_X1 U17590 ( .A1(n14025), .A2(n25197), .ZN(n14027) );
  OAI21_X1 U17591 ( .B1(n14337), .B2(n14027), .A(n14026), .ZN(n14030) );
  NAND2_X1 U17592 ( .A1(n14028), .A2(n14336), .ZN(n14029) );
  NAND2_X1 U17593 ( .A1(n14033), .A2(n14032), .ZN(n14037) );
  NOR2_X1 U17594 ( .A1(n14150), .A2(n14034), .ZN(n14036) );
  XNOR2_X1 U17595 ( .A(n15506), .B(n14846), .ZN(n15150) );
  NOR2_X1 U17596 ( .A1(n14321), .A2(n3401), .ZN(n14038) );
  NOR2_X1 U17597 ( .A1(n14319), .A2(n14458), .ZN(n14039) );
  OAI21_X1 U17598 ( .B1(n14039), .B2(n14320), .A(n14321), .ZN(n14040) );
  NOR2_X1 U17599 ( .A1(n14330), .A2(n14041), .ZN(n14042) );
  XNOR2_X1 U17600 ( .A(n15095), .B(n15298), .ZN(n14046) );
  XNOR2_X1 U17601 ( .A(n14800), .B(n19392), .ZN(n14045) );
  XNOR2_X1 U17602 ( .A(n14046), .B(n14045), .ZN(n14047) );
  NAND2_X1 U17603 ( .A1(n14050), .A2(n14049), .ZN(n14051) );
  NAND2_X1 U17604 ( .A1(n14053), .A2(n14051), .ZN(n14057) );
  NOR2_X1 U17605 ( .A1(n14052), .A2(n14054), .ZN(n14056) );
  XNOR2_X1 U17606 ( .A(n15119), .B(n641), .ZN(n14061) );
  XNOR2_X1 U17607 ( .A(n14061), .B(n15133), .ZN(n14084) );
  INV_X1 U17608 ( .A(n14069), .ZN(n14062) );
  NOR2_X1 U17609 ( .A1(n14062), .A2(n14063), .ZN(n14072) );
  NAND2_X1 U17610 ( .A1(n14064), .A2(n14063), .ZN(n14264) );
  INV_X1 U17611 ( .A(n14065), .ZN(n14066) );
  AOI21_X1 U17613 ( .B1(n13627), .B2(n14067), .A(n300), .ZN(n14068) );
  NAND2_X1 U17614 ( .A1(n14069), .A2(n14068), .ZN(n14070) );
  NAND2_X1 U17616 ( .A1(n14074), .A2(n14073), .ZN(n14082) );
  XNOR2_X1 U17618 ( .A(n15497), .B(n15274), .ZN(n14725) );
  XNOR2_X1 U17619 ( .A(n14084), .B(n14725), .ZN(n14095) );
  XNOR2_X1 U17620 ( .A(n14553), .B(n14516), .ZN(n14093) );
  INV_X1 U17621 ( .A(n14085), .ZN(n14086) );
  NAND2_X1 U17622 ( .A1(n14092), .A2(n14087), .ZN(n14091) );
  XNOR2_X1 U17623 ( .A(n14093), .B(n15321), .ZN(n14094) );
  NAND2_X1 U17624 ( .A1(n4892), .A2(n25445), .ZN(n14097) );
  NOR2_X1 U17625 ( .A1(n14101), .A2(n24376), .ZN(n14102) );
  MUX2_X1 U17626 ( .A(n14107), .B(n14106), .S(n14105), .Z(n14114) );
  NOR2_X1 U17627 ( .A1(n14109), .A2(n14108), .ZN(n14110) );
  NOR2_X1 U17628 ( .A1(n14111), .A2(n14110), .ZN(n14113) );
  XNOR2_X1 U17629 ( .A(n15082), .B(n15401), .ZN(n14403) );
  XNOR2_X1 U17630 ( .A(n14403), .B(n14115), .ZN(n14137) );
  INV_X1 U17631 ( .A(n14116), .ZN(n14117) );
  NAND2_X1 U17632 ( .A1(n14118), .A2(n14117), .ZN(n14120) );
  XNOR2_X1 U17633 ( .A(n15284), .B(n15480), .ZN(n14731) );
  AND2_X1 U17636 ( .A1(n14130), .A2(n1331), .ZN(n14131) );
  XNOR2_X1 U17637 ( .A(n15415), .B(n4164), .ZN(n14135) );
  XNOR2_X1 U17638 ( .A(n14731), .B(n14135), .ZN(n14136) );
  XNOR2_X1 U17639 ( .A(n14137), .B(n14136), .ZN(n15905) );
  NOR2_X1 U17640 ( .A1(n16368), .A2(n15905), .ZN(n15641) );
  INV_X1 U17641 ( .A(n15641), .ZN(n14139) );
  NAND2_X1 U17642 ( .A1(n14139), .A2(n14138), .ZN(n14176) );
  XNOR2_X1 U17643 ( .A(n14858), .B(n3131), .ZN(n14155) );
  NAND2_X1 U17644 ( .A1(n14200), .A2(n3888), .ZN(n14148) );
  OAI21_X1 U17645 ( .B1(n14945), .B2(n14944), .A(n2684), .ZN(n14146) );
  XNOR2_X1 U17646 ( .A(n15526), .B(n15055), .ZN(n14541) );
  XNOR2_X1 U17647 ( .A(n14155), .B(n14541), .ZN(n14175) );
  NAND2_X1 U17648 ( .A1(n14159), .A2(n14158), .ZN(n14161) );
  NAND2_X1 U17649 ( .A1(n14161), .A2(n14160), .ZN(n14162) );
  NAND2_X1 U17650 ( .A1(n14163), .A2(n14162), .ZN(n14897) );
  NAND3_X1 U17651 ( .A1(n14169), .A2(n14168), .A3(n14167), .ZN(n14170) );
  XNOR2_X1 U17652 ( .A(n14809), .B(n14897), .ZN(n15102) );
  XNOR2_X1 U17653 ( .A(n14806), .B(n15169), .ZN(n14173) );
  XNOR2_X1 U17654 ( .A(n14173), .B(n15102), .ZN(n14174) );
  XNOR2_X1 U17655 ( .A(n14892), .B(n15002), .ZN(n14373) );
  MUX2_X1 U17656 ( .A(n24949), .B(n14179), .S(n14178), .Z(n14184) );
  XNOR2_X1 U17657 ( .A(n14185), .B(n14642), .ZN(n14186) );
  NAND2_X1 U17658 ( .A1(n25560), .A2(n25360), .ZN(n14192) );
  NOR2_X1 U17660 ( .A1(n25560), .A2(n14194), .ZN(n14196) );
  NAND2_X1 U17661 ( .A1(n14201), .A2(n14200), .ZN(n14203) );
  OAI21_X1 U17662 ( .B1(n14206), .B2(n14205), .A(n14204), .ZN(n14207) );
  AOI22_X2 U17663 ( .A1(n14210), .A2(n14209), .B1(n14207), .B2(n2378), .ZN(
        n15409) );
  XNOR2_X1 U17664 ( .A(n15409), .B(n14377), .ZN(n14972) );
  OAI21_X1 U17665 ( .B1(n24503), .B2(n13417), .A(n14211), .ZN(n14214) );
  NAND2_X1 U17666 ( .A1(n14214), .A2(n14213), .ZN(n14215) );
  OAI21_X1 U17667 ( .B1(n14217), .B2(n14216), .A(n14215), .ZN(n15164) );
  XNOR2_X1 U17668 ( .A(n15164), .B(n15054), .ZN(n14860) );
  XNOR2_X1 U17669 ( .A(n14860), .B(n14972), .ZN(n14229) );
  XNOR2_X1 U17670 ( .A(n14719), .B(n3073), .ZN(n14227) );
  OAI21_X1 U17671 ( .B1(n14219), .B2(n14218), .A(n14221), .ZN(n14220) );
  NAND3_X1 U17672 ( .A1(n14223), .A2(n14222), .A3(n14221), .ZN(n14224) );
  XNOR2_X1 U17673 ( .A(n14694), .B(n25384), .ZN(n14896) );
  XNOR2_X1 U17674 ( .A(n14896), .B(n14227), .ZN(n14228) );
  XNOR2_X1 U17675 ( .A(n14845), .B(n15369), .ZN(n14239) );
  XNOR2_X1 U17676 ( .A(n14911), .B(n14239), .ZN(n14263) );
  NAND3_X1 U17677 ( .A1(n14241), .A2(n14245), .A3(n14240), .ZN(n14248) );
  NAND3_X1 U17678 ( .A1(n14245), .A2(n13633), .A3(n14244), .ZN(n14246) );
  XNOR2_X1 U17679 ( .A(n14907), .B(n2039), .ZN(n14249) );
  XNOR2_X1 U17680 ( .A(n14737), .B(n14249), .ZN(n14261) );
  OR2_X1 U17682 ( .A1(n14254), .A2(n14253), .ZN(n14258) );
  NAND2_X1 U17683 ( .A1(n14256), .A2(n14255), .ZN(n14257) );
  XNOR2_X1 U17684 ( .A(n14958), .B(n15505), .ZN(n15366) );
  XNOR2_X1 U17685 ( .A(n14261), .B(n15366), .ZN(n14262) );
  XNOR2_X1 U17686 ( .A(n295), .B(n14900), .ZN(n14354) );
  XNOR2_X1 U17687 ( .A(n15033), .B(n15375), .ZN(n14266) );
  XNOR2_X1 U17688 ( .A(n14354), .B(n14266), .ZN(n14286) );
  OAI21_X1 U17689 ( .B1(n14268), .B2(n14267), .A(n397), .ZN(n14273) );
  NAND2_X1 U17690 ( .A1(n14274), .A2(n14269), .ZN(n14270) );
  NOR2_X2 U17692 ( .A1(n14277), .A2(n14276), .ZN(n14902) );
  XNOR2_X1 U17693 ( .A(n14902), .B(n15514), .ZN(n14284) );
  NOR2_X1 U17694 ( .A1(n14850), .A2(n14278), .ZN(n14279) );
  OAI21_X1 U17695 ( .B1(n14849), .B2(n14852), .A(n14279), .ZN(n14282) );
  NAND2_X1 U17696 ( .A1(n14280), .A2(n14415), .ZN(n14281) );
  OAI211_X1 U17697 ( .C1(n24572), .C2(n14415), .A(n14281), .B(n14282), .ZN(
        n15378) );
  XNOR2_X1 U17698 ( .A(n15378), .B(n4189), .ZN(n14283) );
  XNOR2_X1 U17699 ( .A(n14284), .B(n14283), .ZN(n14285) );
  XNOR2_X1 U17700 ( .A(n14285), .B(n14286), .ZN(n14350) );
  INV_X1 U17701 ( .A(n14350), .ZN(n16382) );
  OAI21_X1 U17702 ( .B1(n15656), .B2(n25210), .A(n15990), .ZN(n14352) );
  XNOR2_X1 U17703 ( .A(n14724), .B(n494), .ZN(n14288) );
  XNOR2_X1 U17704 ( .A(n14288), .B(n14287), .ZN(n14316) );
  OAI21_X1 U17705 ( .B1(n394), .B2(n14290), .A(n14289), .ZN(n14297) );
  NAND3_X1 U17707 ( .A1(n14294), .A2(n14293), .A3(n14292), .ZN(n14295) );
  XNOR2_X1 U17708 ( .A(n14634), .B(n15396), .ZN(n15495) );
  NOR2_X1 U17709 ( .A1(n14302), .A2(n1527), .ZN(n14300) );
  NOR2_X1 U17710 ( .A1(n14301), .A2(n13888), .ZN(n14299) );
  AOI22_X1 U17711 ( .A1(n14300), .A2(n13728), .B1(n14299), .B2(n1527), .ZN(
        n14305) );
  NAND2_X1 U17712 ( .A1(n14302), .A2(n14301), .ZN(n14303) );
  INV_X1 U17713 ( .A(n14307), .ZN(n14315) );
  OAI21_X1 U17714 ( .B1(n14310), .B2(n14309), .A(n14308), .ZN(n14313) );
  OAI211_X1 U17715 ( .C1(n14315), .C2(n14314), .A(n14313), .B(n14312), .ZN(
        n15204) );
  XNOR2_X1 U17716 ( .A(n15204), .B(n15275), .ZN(n15398) );
  NOR2_X1 U17717 ( .A1(n14321), .A2(n14320), .ZN(n14322) );
  XNOR2_X1 U17718 ( .A(n15238), .B(n14982), .ZN(n14332) );
  MUX2_X1 U17719 ( .A(n14325), .B(n14327), .S(n14324), .Z(n14326) );
  XNOR2_X1 U17721 ( .A(n14332), .B(n14331), .ZN(n14349) );
  OAI21_X1 U17722 ( .B1(n14335), .B2(n14334), .A(n14333), .ZN(n14343) );
  NAND2_X1 U17723 ( .A1(n14337), .A2(n14336), .ZN(n14342) );
  NAND3_X1 U17724 ( .A1(n14340), .A2(n14339), .A3(n25197), .ZN(n14341) );
  OAI211_X2 U17725 ( .C1(n14344), .C2(n14343), .A(n14342), .B(n14341), .ZN(
        n15387) );
  XNOR2_X1 U17726 ( .A(n14345), .B(n15387), .ZN(n14347) );
  XNOR2_X1 U17727 ( .A(n15488), .B(n449), .ZN(n14346) );
  XNOR2_X1 U17728 ( .A(n14347), .B(n14346), .ZN(n14348) );
  XNOR2_X1 U17729 ( .A(n14348), .B(n14349), .ZN(n15657) );
  OAI21_X1 U17731 ( .B1(n16383), .B2(n16177), .A(n15837), .ZN(n14351) );
  INV_X1 U17732 ( .A(n14354), .ZN(n14356) );
  XNOR2_X1 U17733 ( .A(n24975), .B(n62), .ZN(n14355) );
  XOR2_X1 U17734 ( .A(n14356), .B(n14355), .Z(n14358) );
  XNOR2_X1 U17735 ( .A(n15515), .B(n15444), .ZN(n15113) );
  XNOR2_X1 U17736 ( .A(n15113), .B(n15513), .ZN(n14357) );
  NAND2_X1 U17737 ( .A1(n14359), .A2(n3701), .ZN(n14367) );
  NOR2_X1 U17738 ( .A1(n24995), .A2(n3701), .ZN(n14365) );
  XNOR2_X1 U17739 ( .A(n14368), .B(n15487), .ZN(n14920) );
  XNOR2_X1 U17740 ( .A(n15486), .B(n2193), .ZN(n14369) );
  XNOR2_X1 U17741 ( .A(n14920), .B(n14369), .ZN(n14372) );
  XNOR2_X1 U17742 ( .A(n15436), .B(n15484), .ZN(n15087) );
  XNOR2_X1 U17743 ( .A(n15087), .B(n14370), .ZN(n14371) );
  XNOR2_X1 U17744 ( .A(n24956), .B(n14644), .ZN(n14780) );
  XNOR2_X1 U17745 ( .A(n14780), .B(n14373), .ZN(n14376) );
  XNOR2_X1 U17746 ( .A(n15284), .B(n2881), .ZN(n14374) );
  XNOR2_X1 U17747 ( .A(n14375), .B(n14376), .ZN(n16156) );
  INV_X1 U17748 ( .A(n16156), .ZN(n16154) );
  XNOR2_X1 U17749 ( .A(n25431), .B(n14719), .ZN(n15012) );
  XNOR2_X1 U17750 ( .A(n15012), .B(n15106), .ZN(n14380) );
  XNOR2_X1 U17751 ( .A(n15055), .B(n23883), .ZN(n14378) );
  XNOR2_X1 U17752 ( .A(n14898), .B(n14378), .ZN(n14379) );
  NAND2_X1 U17753 ( .A1(n16122), .A2(n15842), .ZN(n14381) );
  NAND2_X1 U17755 ( .A1(n16156), .A2(n25449), .ZN(n15619) );
  INV_X1 U17756 ( .A(n15619), .ZN(n14388) );
  XNOR2_X1 U17757 ( .A(n14724), .B(n14383), .ZN(n15016) );
  XNOR2_X1 U17758 ( .A(n15393), .B(n15464), .ZN(n15123) );
  XNOR2_X1 U17759 ( .A(n15274), .B(n1768), .ZN(n14385) );
  XNOR2_X1 U17760 ( .A(n15123), .B(n14385), .ZN(n14386) );
  XNOR2_X1 U17761 ( .A(n14387), .B(n14386), .ZN(n16123) );
  INV_X1 U17762 ( .A(n16123), .ZN(n16155) );
  NAND2_X1 U17763 ( .A1(n14388), .A2(n16155), .ZN(n14395) );
  XNOR2_X1 U17764 ( .A(n15298), .B(n21742), .ZN(n14390) );
  XNOR2_X1 U17765 ( .A(n15504), .B(n14390), .ZN(n14393) );
  INV_X1 U17766 ( .A(n15507), .ZN(n14391) );
  XNOR2_X1 U17767 ( .A(n14392), .B(n14393), .ZN(n16125) );
  NAND3_X1 U17768 ( .A1(n24459), .A2(n381), .A3(n16122), .ZN(n14394) );
  INV_X1 U17769 ( .A(n14398), .ZN(n23602) );
  OAI21_X1 U17770 ( .B1(n5487), .B2(n14397), .A(n23602), .ZN(n14400) );
  NAND3_X1 U17771 ( .A1(n5486), .A2(n14398), .A3(n2556), .ZN(n14399) );
  NAND2_X1 U17772 ( .A1(n14400), .A2(n14399), .ZN(n14401) );
  XNOR2_X1 U17773 ( .A(n14402), .B(n14401), .ZN(n14404) );
  XNOR2_X1 U17774 ( .A(n14880), .B(n14642), .ZN(n14891) );
  INV_X1 U17775 ( .A(n16170), .ZN(n16424) );
  XNOR2_X1 U17776 ( .A(n14634), .B(n15200), .ZN(n14406) );
  XNOR2_X1 U17777 ( .A(n15119), .B(n3125), .ZN(n14405) );
  XNOR2_X1 U17778 ( .A(n14406), .B(n14405), .ZN(n14408) );
  XNOR2_X1 U17779 ( .A(n15273), .B(n14591), .ZN(n15201) );
  XNOR2_X1 U17780 ( .A(n15201), .B(n15270), .ZN(n14407) );
  XNOR2_X1 U17781 ( .A(n14408), .B(n14407), .ZN(n16426) );
  INV_X1 U17782 ( .A(n16426), .ZN(n16169) );
  XNOR2_X1 U17783 ( .A(n15170), .B(n15268), .ZN(n14412) );
  INV_X1 U17784 ( .A(n15522), .ZN(n14409) );
  XNOR2_X1 U17785 ( .A(n14409), .B(n15169), .ZN(n14562) );
  XNOR2_X1 U17786 ( .A(n14809), .B(n2137), .ZN(n14410) );
  XNOR2_X1 U17787 ( .A(n14562), .B(n14410), .ZN(n14411) );
  NAND2_X1 U17788 ( .A1(n16169), .A2(n15958), .ZN(n14433) );
  INV_X1 U17789 ( .A(n20284), .ZN(n23523) );
  AOI21_X1 U17790 ( .B1(n14849), .B2(n14416), .A(n14415), .ZN(n14417) );
  OAI21_X1 U17791 ( .B1(n24572), .B2(n14849), .A(n14417), .ZN(n14418) );
  NAND2_X1 U17792 ( .A1(n14419), .A2(n14418), .ZN(n14420) );
  XNOR2_X1 U17793 ( .A(n14799), .B(n14420), .ZN(n15299) );
  XNOR2_X1 U17794 ( .A(n15188), .B(n15299), .ZN(n14421) );
  OAI21_X1 U17795 ( .B1(n16169), .B2(n244), .A(n16427), .ZN(n14427) );
  XNOR2_X1 U17796 ( .A(n14928), .B(n14468), .ZN(n15208) );
  XNOR2_X1 U17797 ( .A(n15290), .B(n15208), .ZN(n14426) );
  XNOR2_X1 U17798 ( .A(n14919), .B(n2795), .ZN(n14424) );
  XNOR2_X1 U17799 ( .A(n14423), .B(n14424), .ZN(n14425) );
  NAND2_X1 U17800 ( .A1(n14427), .A2(n1329), .ZN(n14432) );
  XNOR2_X1 U17801 ( .A(n15190), .B(n859), .ZN(n14428) );
  INV_X1 U17802 ( .A(n16422), .ZN(n15961) );
  NAND3_X1 U17803 ( .A1(n15961), .A2(n707), .A3(n16169), .ZN(n14431) );
  NOR2_X1 U17804 ( .A1(n17283), .A2(n17229), .ZN(n16952) );
  INV_X1 U17805 ( .A(n14434), .ZN(n14438) );
  NOR2_X1 U17806 ( .A1(n14438), .A2(n14437), .ZN(n14441) );
  XNOR2_X1 U17808 ( .A(n15223), .B(n14816), .ZN(n14443) );
  XNOR2_X1 U17809 ( .A(n14442), .B(n15415), .ZN(n14729) );
  XNOR2_X1 U17810 ( .A(n15177), .B(n15416), .ZN(n14444) );
  XNOR2_X1 U17811 ( .A(n15230), .B(n14806), .ZN(n14446) );
  XNOR2_X1 U17812 ( .A(n15168), .B(n15056), .ZN(n14445) );
  XNOR2_X1 U17813 ( .A(n14446), .B(n14445), .ZN(n14450) );
  XNOR2_X1 U17814 ( .A(n14620), .B(n14858), .ZN(n14448) );
  XNOR2_X1 U17815 ( .A(n14857), .B(n2049), .ZN(n14447) );
  XNOR2_X1 U17816 ( .A(n14448), .B(n14447), .ZN(n14449) );
  XNOR2_X1 U17817 ( .A(n14450), .B(n14449), .ZN(n16408) );
  XNOR2_X1 U17818 ( .A(n14800), .B(n21662), .ZN(n14451) );
  XNOR2_X1 U17819 ( .A(n15253), .B(n14669), .ZN(n14452) );
  XNOR2_X1 U17820 ( .A(n14988), .B(n14846), .ZN(n14739) );
  XNOR2_X1 U17821 ( .A(n14739), .B(n15358), .ZN(n15456) );
  XNOR2_X1 U17822 ( .A(n15456), .B(n14453), .ZN(n16414) );
  INV_X1 U17823 ( .A(n16414), .ZN(n16140) );
  XNOR2_X1 U17824 ( .A(n15244), .B(n24287), .ZN(n14454) );
  XNOR2_X1 U17825 ( .A(n25008), .B(n15190), .ZN(n14455) );
  XNOR2_X1 U17826 ( .A(n14456), .B(n14455), .ZN(n14465) );
  INV_X1 U17827 ( .A(n14457), .ZN(n14462) );
  AND2_X1 U17828 ( .A1(n14458), .A2(n14459), .ZN(n14461) );
  XNOR2_X1 U17829 ( .A(n15153), .B(n14463), .ZN(n14464) );
  XNOR2_X1 U17830 ( .A(n15347), .B(n14464), .ZN(n15449) );
  XNOR2_X2 U17831 ( .A(n14465), .B(n15449), .ZN(n16412) );
  NAND2_X1 U17832 ( .A1(n16140), .A2(n16412), .ZN(n15653) );
  INV_X1 U17833 ( .A(n16408), .ZN(n16416) );
  XNOR2_X1 U17834 ( .A(n15138), .B(n14976), .ZN(n14467) );
  XNOR2_X1 U17835 ( .A(n14467), .B(n14466), .ZN(n15441) );
  XNOR2_X1 U17836 ( .A(n14755), .B(n14792), .ZN(n14470) );
  XNOR2_X1 U17837 ( .A(n14468), .B(n836), .ZN(n14469) );
  XNOR2_X1 U17838 ( .A(n15441), .B(n14471), .ZN(n15986) );
  INV_X1 U17839 ( .A(n15986), .ZN(n16409) );
  INV_X1 U17840 ( .A(n16412), .ZN(n14472) );
  XNOR2_X1 U17841 ( .A(n15203), .B(n14516), .ZN(n14831) );
  XNOR2_X1 U17842 ( .A(n15462), .B(n14831), .ZN(n14476) );
  XNOR2_X1 U17843 ( .A(n14703), .B(n15219), .ZN(n14474) );
  XNOR2_X1 U17844 ( .A(n24418), .B(n1874), .ZN(n14473) );
  XNOR2_X1 U17845 ( .A(n14474), .B(n14473), .ZN(n14475) );
  XNOR2_X1 U17846 ( .A(n14476), .B(n14475), .ZN(n16417) );
  INV_X1 U17847 ( .A(n16417), .ZN(n15868) );
  XNOR2_X1 U17848 ( .A(n15238), .B(n15488), .ZN(n15385) );
  XNOR2_X1 U17849 ( .A(n14865), .B(n14792), .ZN(n15293) );
  XNOR2_X1 U17850 ( .A(n15385), .B(n15293), .ZN(n14481) );
  XNOR2_X1 U17851 ( .A(n14977), .B(n14477), .ZN(n14479) );
  XNOR2_X1 U17852 ( .A(n14468), .B(n673), .ZN(n14478) );
  XNOR2_X1 U17853 ( .A(n14479), .B(n14478), .ZN(n14480) );
  XNOR2_X1 U17854 ( .A(n15359), .B(n3164), .ZN(n14482) );
  XNOR2_X1 U17855 ( .A(n14482), .B(n15369), .ZN(n14483) );
  XNOR2_X1 U17856 ( .A(n14483), .B(n14909), .ZN(n14486) );
  INV_X1 U17857 ( .A(n14800), .ZN(n14484) );
  XNOR2_X1 U17858 ( .A(n14484), .B(n14845), .ZN(n15297) );
  XNOR2_X1 U17859 ( .A(n15297), .B(n15188), .ZN(n14485) );
  XNOR2_X1 U17860 ( .A(n15514), .B(n4233), .ZN(n14487) );
  XNOR2_X1 U17861 ( .A(n14487), .B(n15375), .ZN(n14492) );
  INV_X1 U17862 ( .A(n15033), .ZN(n14489) );
  XNOR2_X1 U17863 ( .A(n14488), .B(n14489), .ZN(n15303) );
  XNOR2_X1 U17864 ( .A(n15280), .B(n14494), .ZN(n14498) );
  XNOR2_X1 U17865 ( .A(n15476), .B(n15417), .ZN(n14496) );
  INV_X1 U17866 ( .A(n14558), .ZN(n15333) );
  XNOR2_X1 U17867 ( .A(n15333), .B(n1869), .ZN(n14495) );
  XNOR2_X1 U17868 ( .A(n14495), .B(n14496), .ZN(n14497) );
  XNOR2_X1 U17869 ( .A(n14498), .B(n14497), .ZN(n14499) );
  OAI21_X1 U17870 ( .B1(n15856), .B2(n15611), .A(n16118), .ZN(n14522) );
  INV_X1 U17871 ( .A(n14499), .ZN(n16113) );
  XNOR2_X1 U17873 ( .A(n14694), .B(n2765), .ZN(n15407) );
  XNOR2_X1 U17874 ( .A(n15407), .B(n15267), .ZN(n14504) );
  XNOR2_X1 U17875 ( .A(n15431), .B(n14620), .ZN(n14502) );
  XNOR2_X1 U17876 ( .A(n15326), .B(n3178), .ZN(n14501) );
  XNOR2_X1 U17877 ( .A(n14502), .B(n14501), .ZN(n14503) );
  NAND2_X1 U17878 ( .A1(n16113), .A2(n15857), .ZN(n16680) );
  OAI21_X1 U17879 ( .B1(n16117), .B2(n15856), .A(n16680), .ZN(n14521) );
  INV_X1 U17880 ( .A(n15204), .ZN(n14505) );
  XNOR2_X1 U17881 ( .A(n15463), .B(n14505), .ZN(n14873) );
  MUX2_X1 U17882 ( .A(n14512), .B(n14511), .S(n14510), .Z(n14515) );
  INV_X1 U17883 ( .A(n14513), .ZN(n14514) );
  XNOR2_X1 U17884 ( .A(n15063), .B(n14516), .ZN(n15271) );
  XNOR2_X1 U17885 ( .A(n15271), .B(n14873), .ZN(n14520) );
  XNOR2_X1 U17886 ( .A(n25443), .B(n14591), .ZN(n14518) );
  XNOR2_X1 U17887 ( .A(n15396), .B(n1815), .ZN(n14517) );
  XNOR2_X1 U17888 ( .A(n14518), .B(n14517), .ZN(n14519) );
  OR2_X1 U17891 ( .A1(n16952), .A2(n16753), .ZN(n14590) );
  XNOR2_X1 U17892 ( .A(n15318), .B(n15274), .ZN(n14833) );
  XNOR2_X1 U17893 ( .A(n14775), .B(n923), .ZN(n14523) );
  XNOR2_X1 U17894 ( .A(n14523), .B(n15321), .ZN(n14524) );
  XNOR2_X1 U17895 ( .A(n14524), .B(n14833), .ZN(n14527) );
  XNOR2_X1 U17896 ( .A(n14703), .B(n15497), .ZN(n14525) );
  XNOR2_X1 U17897 ( .A(n14525), .B(n15499), .ZN(n14526) );
  INV_X1 U17898 ( .A(n16389), .ZN(n15848) );
  XNOR2_X1 U17899 ( .A(n14731), .B(n15332), .ZN(n14531) );
  XNOR2_X1 U17900 ( .A(n14690), .B(n1351), .ZN(n14529) );
  XNOR2_X1 U17901 ( .A(n14529), .B(n14528), .ZN(n14530) );
  XNOR2_X1 U17902 ( .A(n15338), .B(n14532), .ZN(n14536) );
  XNOR2_X1 U17903 ( .A(n14675), .B(n1801), .ZN(n14533) );
  XNOR2_X1 U17904 ( .A(n14533), .B(n14534), .ZN(n14535) );
  XNOR2_X1 U17905 ( .A(n15506), .B(n15298), .ZN(n14738) );
  XNOR2_X1 U17906 ( .A(n15074), .B(n15095), .ZN(n15355) );
  XNOR2_X1 U17907 ( .A(n14738), .B(n15355), .ZN(n14540) );
  XNOR2_X1 U17908 ( .A(n14671), .B(n14669), .ZN(n14538) );
  XNOR2_X1 U17909 ( .A(n14654), .B(n860), .ZN(n14537) );
  XNOR2_X1 U17910 ( .A(n14538), .B(n14537), .ZN(n14539) );
  INV_X1 U17912 ( .A(n15980), .ZN(n14546) );
  INV_X1 U17913 ( .A(n14897), .ZN(n14629) );
  XNOR2_X1 U17914 ( .A(n14629), .B(n15051), .ZN(n15324) );
  XNOR2_X1 U17915 ( .A(n15324), .B(n14541), .ZN(n14545) );
  XNOR2_X1 U17916 ( .A(n14857), .B(n23679), .ZN(n14542) );
  XNOR2_X1 U17917 ( .A(n14543), .B(n14542), .ZN(n14544) );
  XNOR2_X1 U17918 ( .A(n14545), .B(n14544), .ZN(n16388) );
  INV_X1 U17919 ( .A(n14715), .ZN(n14548) );
  XNOR2_X1 U17920 ( .A(n14548), .B(n14547), .ZN(n14552) );
  XNOR2_X1 U17921 ( .A(n15034), .B(n15109), .ZN(n15348) );
  XNOR2_X1 U17922 ( .A(n14549), .B(n2050), .ZN(n14550) );
  XNOR2_X1 U17923 ( .A(n15348), .B(n14550), .ZN(n14551) );
  INV_X1 U17924 ( .A(n16393), .ZN(n16163) );
  XNOR2_X1 U17925 ( .A(n15464), .B(n1767), .ZN(n14554) );
  XNOR2_X1 U17926 ( .A(n14553), .B(n14554), .ZN(n14555) );
  XNOR2_X1 U17927 ( .A(n14556), .B(n25426), .ZN(n15218) );
  INV_X1 U17928 ( .A(n16151), .ZN(n14747) );
  INV_X1 U17929 ( .A(n14644), .ZN(n15421) );
  XNOR2_X1 U17930 ( .A(n14642), .B(n15421), .ZN(n14557) );
  XNOR2_X1 U17931 ( .A(n14557), .B(n14965), .ZN(n14561) );
  XNOR2_X1 U17932 ( .A(n15282), .B(n14558), .ZN(n15225) );
  XNOR2_X1 U17933 ( .A(n15401), .B(n2240), .ZN(n14559) );
  XNOR2_X1 U17934 ( .A(n15225), .B(n14559), .ZN(n14560) );
  INV_X1 U17935 ( .A(n14562), .ZN(n14564) );
  XNOR2_X1 U17936 ( .A(n15430), .B(n3190), .ZN(n14563) );
  XNOR2_X1 U17937 ( .A(n14564), .B(n14563), .ZN(n14567) );
  INV_X1 U17938 ( .A(n15409), .ZN(n14565) );
  XNOR2_X1 U17939 ( .A(n14565), .B(n15326), .ZN(n15010) );
  XNOR2_X1 U17940 ( .A(n14973), .B(n15010), .ZN(n14566) );
  NAND2_X1 U17941 ( .A1(n293), .A2(n1762), .ZN(n14586) );
  INV_X1 U17942 ( .A(n14919), .ZN(n14568) );
  XNOR2_X1 U17943 ( .A(n14977), .B(n14568), .ZN(n14569) );
  INV_X1 U17944 ( .A(n14922), .ZN(n14868) );
  XNOR2_X1 U17945 ( .A(n14868), .B(n15386), .ZN(n14929) );
  XNOR2_X1 U17946 ( .A(n14929), .B(n14569), .ZN(n14573) );
  XNOR2_X1 U17947 ( .A(n15387), .B(n15210), .ZN(n14571) );
  XNOR2_X1 U17948 ( .A(n15436), .B(n3133), .ZN(n14570) );
  XNOR2_X1 U17949 ( .A(n14571), .B(n14570), .ZN(n14572) );
  XNOR2_X1 U17950 ( .A(n15094), .B(n15183), .ZN(n14961) );
  XNOR2_X1 U17951 ( .A(n15184), .B(n15452), .ZN(n14574) );
  XNOR2_X1 U17952 ( .A(n14961), .B(n14574), .ZN(n14577) );
  XNOR2_X1 U17953 ( .A(n14958), .B(n15359), .ZN(n15252) );
  XNOR2_X1 U17954 ( .A(n14907), .B(n1891), .ZN(n14575) );
  XNOR2_X1 U17955 ( .A(n15252), .B(n14575), .ZN(n14576) );
  XNOR2_X1 U17958 ( .A(n15378), .B(n15350), .ZN(n15246) );
  XNOR2_X1 U17959 ( .A(n14902), .B(n15444), .ZN(n14581) );
  XNOR2_X1 U17960 ( .A(n14579), .B(n2126), .ZN(n14580) );
  XNOR2_X1 U17961 ( .A(n14581), .B(n14580), .ZN(n14582) );
  NOR2_X1 U17962 ( .A1(n16096), .A2(n16147), .ZN(n14584) );
  INV_X1 U17964 ( .A(n17283), .ZN(n17289) );
  NAND3_X1 U17965 ( .A1(n17289), .A2(n17284), .A3(n17229), .ZN(n14587) );
  NAND4_X1 U17966 ( .A1(n14590), .A2(n14589), .A3(n14588), .A4(n14587), .ZN(
        n17653) );
  XNOR2_X1 U17967 ( .A(n17653), .B(n18146), .ZN(n18323) );
  XNOR2_X1 U17968 ( .A(n15318), .B(n24418), .ZN(n14592) );
  INV_X1 U17969 ( .A(n14594), .ZN(n15187) );
  XNOR2_X1 U17970 ( .A(n15094), .B(n15187), .ZN(n14912) );
  INV_X1 U17971 ( .A(n14912), .ZN(n14598) );
  XNOR2_X1 U17972 ( .A(n15507), .B(n15074), .ZN(n14596) );
  XNOR2_X1 U17973 ( .A(n15359), .B(n2882), .ZN(n14595) );
  XNOR2_X1 U17974 ( .A(n14596), .B(n14595), .ZN(n14597) );
  XNOR2_X1 U17975 ( .A(n14600), .B(n14940), .ZN(n14604) );
  XNOR2_X1 U17976 ( .A(n15112), .B(n15194), .ZN(n14602) );
  XNOR2_X1 U17977 ( .A(n15034), .B(n1789), .ZN(n14601) );
  XNOR2_X1 U17978 ( .A(n14602), .B(n14601), .ZN(n14603) );
  XNOR2_X1 U17979 ( .A(n14604), .B(n14603), .ZN(n15262) );
  INV_X1 U17980 ( .A(n15262), .ZN(n15790) );
  INV_X1 U17981 ( .A(n14789), .ZN(n14605) );
  XNOR2_X1 U17982 ( .A(n14605), .B(n15484), .ZN(n14606) );
  XNOR2_X1 U17983 ( .A(n14606), .B(n14920), .ZN(n14610) );
  XNOR2_X1 U17984 ( .A(n14468), .B(n1952), .ZN(n14607) );
  XNOR2_X1 U17985 ( .A(n14608), .B(n14607), .ZN(n14609) );
  NOR2_X1 U17986 ( .A1(n16043), .A2(n15262), .ZN(n16041) );
  INV_X1 U17987 ( .A(n14611), .ZN(n14889) );
  XNOR2_X1 U17988 ( .A(n14889), .B(n15175), .ZN(n14613) );
  XNOR2_X1 U17989 ( .A(n24937), .B(n22702), .ZN(n14612) );
  XNOR2_X1 U17990 ( .A(n14613), .B(n14612), .ZN(n14617) );
  INV_X1 U17991 ( .A(n14614), .ZN(n14615) );
  XNOR2_X1 U17992 ( .A(n14615), .B(n14964), .ZN(n14616) );
  XNOR2_X1 U17993 ( .A(n14616), .B(n14617), .ZN(n14625) );
  OAI21_X1 U17994 ( .B1(n16041), .B2(n291), .A(n16038), .ZN(n14627) );
  INV_X1 U17995 ( .A(n14898), .ZN(n14618) );
  XNOR2_X1 U17996 ( .A(n14619), .B(n14618), .ZN(n14624) );
  XNOR2_X1 U17997 ( .A(n14620), .B(n15051), .ZN(n14622) );
  XNOR2_X1 U17998 ( .A(n15103), .B(n1863), .ZN(n14621) );
  XNOR2_X1 U17999 ( .A(n14622), .B(n14621), .ZN(n14623) );
  NAND3_X1 U18000 ( .A1(n2251), .A2(n24430), .A3(n15789), .ZN(n14626) );
  XNOR2_X1 U18001 ( .A(n15522), .B(n23983), .ZN(n14628) );
  XNOR2_X1 U18002 ( .A(n14858), .B(n14628), .ZN(n14631) );
  XNOR2_X1 U18003 ( .A(n14629), .B(n24508), .ZN(n15011) );
  INV_X1 U18004 ( .A(n15011), .ZN(n14630) );
  XNOR2_X1 U18005 ( .A(n14631), .B(n14630), .ZN(n14632) );
  XNOR2_X1 U18006 ( .A(n14634), .B(n1776), .ZN(n14635) );
  XNOR2_X1 U18007 ( .A(n14635), .B(n15321), .ZN(n14637) );
  XNOR2_X1 U18008 ( .A(n15133), .B(n15318), .ZN(n14636) );
  XNOR2_X1 U18009 ( .A(n14637), .B(n14636), .ZN(n14641) );
  INV_X1 U18010 ( .A(n14638), .ZN(n14639) );
  XNOR2_X1 U18011 ( .A(n14639), .B(n15499), .ZN(n14640) );
  XNOR2_X1 U18012 ( .A(n14642), .B(n15005), .ZN(n15482) );
  INV_X1 U18013 ( .A(n15332), .ZN(n14643) );
  XNOR2_X1 U18014 ( .A(n14643), .B(n15482), .ZN(n14648) );
  XNOR2_X1 U18015 ( .A(n14644), .B(n15415), .ZN(n14646) );
  XNOR2_X1 U18016 ( .A(n15003), .B(n889), .ZN(n14645) );
  XNOR2_X1 U18017 ( .A(n14646), .B(n14645), .ZN(n14647) );
  XNOR2_X1 U18018 ( .A(n15138), .B(n21623), .ZN(n14650) );
  XNOR2_X1 U18019 ( .A(n14649), .B(n14650), .ZN(n14651) );
  XNOR2_X1 U18020 ( .A(n14651), .B(n14652), .ZN(n14664) );
  INV_X1 U18021 ( .A(n14664), .ZN(n15799) );
  XNOR2_X1 U18022 ( .A(n15071), .B(n15095), .ZN(n14987) );
  XNOR2_X1 U18023 ( .A(n14987), .B(n14653), .ZN(n14657) );
  XNOR2_X1 U18024 ( .A(n14846), .B(n876), .ZN(n14655) );
  XNOR2_X1 U18025 ( .A(n14654), .B(n14907), .ZN(n15503) );
  XNOR2_X1 U18026 ( .A(n14655), .B(n15503), .ZN(n14656) );
  NAND2_X1 U18027 ( .A1(n15799), .A2(n16129), .ZN(n16131) );
  INV_X1 U18028 ( .A(n16129), .ZN(n15800) );
  XNOR2_X1 U18029 ( .A(n14902), .B(n14996), .ZN(n15247) );
  INV_X1 U18030 ( .A(n15247), .ZN(n15512) );
  XNOR2_X1 U18031 ( .A(n15512), .B(n15348), .ZN(n14661) );
  XNOR2_X1 U18032 ( .A(n14993), .B(n15444), .ZN(n14659) );
  XNOR2_X1 U18033 ( .A(n15153), .B(n891), .ZN(n14658) );
  XNOR2_X1 U18034 ( .A(n14659), .B(n14658), .ZN(n14660) );
  INV_X1 U18035 ( .A(n16076), .ZN(n16130) );
  NAND2_X1 U18036 ( .A1(n16131), .A2(n14662), .ZN(n14663) );
  NAND2_X1 U18037 ( .A1(n16077), .A2(n16129), .ZN(n15312) );
  INV_X1 U18038 ( .A(n15312), .ZN(n14665) );
  NAND2_X1 U18039 ( .A1(n14665), .A2(n1365), .ZN(n14666) );
  XNOR2_X1 U18040 ( .A(n15374), .B(n14827), .ZN(n15156) );
  XNOR2_X1 U18041 ( .A(n14667), .B(n14826), .ZN(n15447) );
  XNOR2_X1 U18042 ( .A(n15347), .B(n14936), .ZN(n15195) );
  XNOR2_X1 U18043 ( .A(n15514), .B(n869), .ZN(n14668) );
  INV_X1 U18044 ( .A(n14669), .ZN(n14670) );
  XNOR2_X1 U18045 ( .A(n14670), .B(n14799), .ZN(n15147) );
  XNOR2_X1 U18046 ( .A(n14671), .B(n15097), .ZN(n15454) );
  XNOR2_X1 U18047 ( .A(n15454), .B(n15147), .ZN(n14674) );
  XNOR2_X1 U18048 ( .A(n15505), .B(n22986), .ZN(n14672) );
  XNOR2_X1 U18049 ( .A(n15185), .B(n14672), .ZN(n14673) );
  INV_X1 U18050 ( .A(n14676), .ZN(n14791) );
  XNOR2_X1 U18051 ( .A(n1362), .B(n14791), .ZN(n15139) );
  XNOR2_X1 U18052 ( .A(n14677), .B(n15139), .ZN(n14681) );
  XNOR2_X1 U18053 ( .A(n14678), .B(n15088), .ZN(n15438) );
  XNOR2_X1 U18054 ( .A(n15488), .B(n2211), .ZN(n14679) );
  XNOR2_X1 U18055 ( .A(n15438), .B(n14679), .ZN(n14680) );
  INV_X1 U18056 ( .A(n14686), .ZN(n14684) );
  INV_X1 U18057 ( .A(n14685), .ZN(n14683) );
  INV_X1 U18058 ( .A(n2989), .ZN(n14682) );
  OAI21_X1 U18059 ( .B1(n14684), .B2(n14683), .A(n14682), .ZN(n14688) );
  NAND3_X1 U18060 ( .A1(n14686), .A2(n2989), .A3(n14685), .ZN(n14687) );
  NAND2_X1 U18061 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  XNOR2_X1 U18062 ( .A(n15082), .B(n14690), .ZN(n15420) );
  XNOR2_X1 U18063 ( .A(n15420), .B(n14691), .ZN(n14692) );
  NAND2_X1 U18064 ( .A1(n24532), .A2(n16109), .ZN(n14702) );
  XNOR2_X1 U18065 ( .A(n14694), .B(n14805), .ZN(n14696) );
  XNOR2_X1 U18066 ( .A(n14857), .B(n2100), .ZN(n14695) );
  XNOR2_X1 U18067 ( .A(n14696), .B(n14695), .ZN(n14701) );
  XNOR2_X1 U18068 ( .A(n14697), .B(n14698), .ZN(n15429) );
  XNOR2_X1 U18069 ( .A(n14699), .B(n15429), .ZN(n14700) );
  XNOR2_X1 U18070 ( .A(n14834), .B(n14703), .ZN(n15131) );
  XNOR2_X1 U18071 ( .A(n15131), .B(n14704), .ZN(n14707) );
  XNOR2_X1 U18072 ( .A(n15396), .B(n881), .ZN(n14705) );
  XNOR2_X1 U18073 ( .A(n15461), .B(n14705), .ZN(n14706) );
  NOR2_X1 U18074 ( .A1(n16107), .A2(n15782), .ZN(n14708) );
  INV_X1 U18076 ( .A(n15804), .ZN(n16114) );
  XNOR2_X1 U18078 ( .A(n14755), .B(n14982), .ZN(n15339) );
  XNOR2_X1 U18079 ( .A(n14928), .B(n14788), .ZN(n15291) );
  XNOR2_X1 U18080 ( .A(n15291), .B(n15339), .ZN(n14713) );
  XNOR2_X1 U18081 ( .A(n15483), .B(n24502), .ZN(n14711) );
  XNOR2_X1 U18082 ( .A(n14976), .B(n5286), .ZN(n14710) );
  XNOR2_X1 U18083 ( .A(n14711), .B(n14710), .ZN(n14712) );
  XNOR2_X1 U18084 ( .A(n14715), .B(n14714), .ZN(n14718) );
  XNOR2_X1 U18085 ( .A(n15153), .B(n2040), .ZN(n14716) );
  XNOR2_X1 U18086 ( .A(n15351), .B(n14716), .ZN(n14717) );
  XNOR2_X1 U18087 ( .A(n15230), .B(n14719), .ZN(n15325) );
  XNOR2_X1 U18088 ( .A(n15526), .B(n1777), .ZN(n14720) );
  XNOR2_X1 U18089 ( .A(n15325), .B(n14720), .ZN(n14723) );
  XNOR2_X1 U18090 ( .A(n15427), .B(n15269), .ZN(n14722) );
  XNOR2_X1 U18091 ( .A(n15462), .B(n15126), .ZN(n14728) );
  XNOR2_X1 U18092 ( .A(n15273), .B(n1835), .ZN(n14726) );
  XNOR2_X1 U18093 ( .A(n14726), .B(n14725), .ZN(n14727) );
  XNOR2_X1 U18094 ( .A(n14728), .B(n14727), .ZN(n16080) );
  NAND2_X1 U18095 ( .A1(n16080), .A2(n15584), .ZN(n16082) );
  INV_X1 U18096 ( .A(n14729), .ZN(n14730) );
  XNOR2_X1 U18097 ( .A(n14730), .B(n15331), .ZN(n14736) );
  INV_X1 U18098 ( .A(n14731), .ZN(n14734) );
  XNOR2_X1 U18099 ( .A(n15285), .B(n20744), .ZN(n14733) );
  XNOR2_X1 U18100 ( .A(n14734), .B(n14733), .ZN(n14735) );
  NOR2_X1 U18101 ( .A1(n16100), .A2(n15584), .ZN(n15780) );
  XNOR2_X1 U18102 ( .A(n14737), .B(n15253), .ZN(n15356) );
  XNOR2_X1 U18103 ( .A(n15356), .B(n14738), .ZN(n14742) );
  INV_X1 U18104 ( .A(n14739), .ZN(n14741) );
  XNOR2_X1 U18105 ( .A(n14960), .B(n2745), .ZN(n14740) );
  INV_X1 U18106 ( .A(n17273), .ZN(n17254) );
  INV_X1 U18107 ( .A(n17272), .ZN(n17279) );
  OAI21_X1 U18108 ( .B1(n16151), .B2(n213), .A(n16095), .ZN(n14744) );
  INV_X1 U18112 ( .A(n14749), .ZN(n14750) );
  XNOR2_X1 U18113 ( .A(n15093), .B(n14750), .ZN(n14754) );
  XNOR2_X1 U18114 ( .A(n14988), .B(n15506), .ZN(n14752) );
  XNOR2_X1 U18115 ( .A(n14799), .B(n924), .ZN(n14751) );
  XNOR2_X1 U18116 ( .A(n14752), .B(n14751), .ZN(n14753) );
  XNOR2_X1 U18117 ( .A(n14754), .B(n14753), .ZN(n15938) );
  XNOR2_X1 U18118 ( .A(n14755), .B(n15484), .ZN(n14758) );
  XNOR2_X1 U18119 ( .A(n14756), .B(n14791), .ZN(n14757) );
  XNOR2_X1 U18120 ( .A(n14757), .B(n14758), .ZN(n14762) );
  XNOR2_X1 U18121 ( .A(n15436), .B(n15483), .ZN(n14760) );
  XNOR2_X1 U18122 ( .A(n14976), .B(n2761), .ZN(n14759) );
  XNOR2_X1 U18123 ( .A(n14760), .B(n14759), .ZN(n14761) );
  XNOR2_X2 U18124 ( .A(n14762), .B(n14761), .ZN(n16247) );
  INV_X1 U18125 ( .A(n15526), .ZN(n14764) );
  XNOR2_X1 U18126 ( .A(n14764), .B(n14805), .ZN(n15159) );
  XNOR2_X1 U18127 ( .A(n15056), .B(n2903), .ZN(n14765) );
  XNOR2_X1 U18128 ( .A(n15159), .B(n14765), .ZN(n14766) );
  XNOR2_X1 U18129 ( .A(n14766), .B(n14767), .ZN(n15764) );
  INV_X1 U18130 ( .A(n15764), .ZN(n16018) );
  NAND2_X1 U18131 ( .A1(n16247), .A2(n16018), .ZN(n14787) );
  XNOR2_X1 U18132 ( .A(n14827), .B(n765), .ZN(n14768) );
  XNOR2_X1 U18133 ( .A(n14769), .B(n14768), .ZN(n14772) );
  XNOR2_X1 U18134 ( .A(n15113), .B(n14770), .ZN(n14771) );
  XNOR2_X1 U18137 ( .A(n14834), .B(n15464), .ZN(n14774) );
  XNOR2_X1 U18138 ( .A(n15062), .B(n15219), .ZN(n14773) );
  XNOR2_X1 U18139 ( .A(n14773), .B(n14774), .ZN(n14779) );
  XNOR2_X1 U18140 ( .A(n15393), .B(n2805), .ZN(n14777) );
  XNOR2_X1 U18141 ( .A(n15497), .B(n14775), .ZN(n14776) );
  XNOR2_X1 U18142 ( .A(n14776), .B(n14777), .ZN(n14778) );
  XNOR2_X1 U18143 ( .A(n14779), .B(n14778), .ZN(n15762) );
  XNOR2_X1 U18145 ( .A(n15480), .B(n14815), .ZN(n15141) );
  INV_X1 U18146 ( .A(n14780), .ZN(n15081) );
  XNOR2_X1 U18147 ( .A(n15081), .B(n15141), .ZN(n14784) );
  XNOR2_X1 U18148 ( .A(n15422), .B(n2120), .ZN(n14782) );
  XNOR2_X1 U18149 ( .A(n14782), .B(n14781), .ZN(n14783) );
  XNOR2_X1 U18150 ( .A(n14789), .B(n14788), .ZN(n15029) );
  INV_X1 U18151 ( .A(n15029), .ZN(n14790) );
  XNOR2_X1 U18152 ( .A(n15238), .B(n15341), .ZN(n15209) );
  XNOR2_X1 U18153 ( .A(n14790), .B(n15209), .ZN(n14796) );
  XNOR2_X1 U18154 ( .A(n15088), .B(n14791), .ZN(n14794) );
  XNOR2_X1 U18155 ( .A(n14792), .B(n2717), .ZN(n14793) );
  XNOR2_X1 U18156 ( .A(n14794), .B(n14793), .ZN(n14795) );
  XNOR2_X1 U18157 ( .A(n15097), .B(n15298), .ZN(n14798) );
  XNOR2_X1 U18158 ( .A(n15358), .B(n15369), .ZN(n14797) );
  XNOR2_X1 U18159 ( .A(n14797), .B(n14798), .ZN(n14804) );
  XNOR2_X1 U18160 ( .A(n14799), .B(n15074), .ZN(n14802) );
  XNOR2_X1 U18161 ( .A(n14800), .B(n763), .ZN(n14801) );
  XNOR2_X1 U18162 ( .A(n14802), .B(n14801), .ZN(n14803) );
  XNOR2_X1 U18164 ( .A(n15168), .B(n14805), .ZN(n14808) );
  XNOR2_X1 U18165 ( .A(n14806), .B(n15051), .ZN(n14807) );
  XNOR2_X1 U18166 ( .A(n14808), .B(n14807), .ZN(n14813) );
  XNOR2_X1 U18167 ( .A(n2765), .B(n15055), .ZN(n14811) );
  XNOR2_X1 U18168 ( .A(n14809), .B(n21335), .ZN(n14810) );
  XNOR2_X1 U18169 ( .A(n14811), .B(n14810), .ZN(n14812) );
  NAND2_X1 U18170 ( .A1(n16491), .A2(n16232), .ZN(n14823) );
  INV_X1 U18171 ( .A(n15416), .ZN(n14814) );
  XNOR2_X1 U18172 ( .A(n14814), .B(n14815), .ZN(n14818) );
  XNOR2_X1 U18173 ( .A(n15082), .B(n14816), .ZN(n14817) );
  XNOR2_X1 U18174 ( .A(n14818), .B(n14817), .ZN(n14822) );
  XNOR2_X1 U18175 ( .A(n15174), .B(n15284), .ZN(n14820) );
  XNOR2_X1 U18176 ( .A(n24937), .B(n21703), .ZN(n14819) );
  XNOR2_X1 U18177 ( .A(n14820), .B(n14819), .ZN(n14821) );
  OAI22_X1 U18178 ( .A1(n16229), .A2(n14823), .B1(n16230), .B2(n16232), .ZN(
        n14839) );
  XNOR2_X1 U18179 ( .A(n15347), .B(n15375), .ZN(n14824) );
  XNOR2_X1 U18180 ( .A(n14825), .B(n14824), .ZN(n14830) );
  XNOR2_X1 U18181 ( .A(n24976), .B(n14826), .ZN(n14829) );
  INV_X1 U18182 ( .A(n896), .ZN(n23798) );
  XNOR2_X1 U18183 ( .A(n14827), .B(n23798), .ZN(n14828) );
  INV_X1 U18184 ( .A(n14831), .ZN(n14832) );
  XNOR2_X1 U18185 ( .A(n14832), .B(n14833), .ZN(n14838) );
  XNOR2_X1 U18186 ( .A(n15119), .B(n1739), .ZN(n14836) );
  XNOR2_X1 U18187 ( .A(n14834), .B(n15204), .ZN(n14835) );
  XNOR2_X1 U18188 ( .A(n14836), .B(n14835), .ZN(n14837) );
  XNOR2_X1 U18189 ( .A(n14838), .B(n14837), .ZN(n16231) );
  INV_X1 U18190 ( .A(n14840), .ZN(n14844) );
  XNOR2_X1 U18191 ( .A(n14841), .B(n15446), .ZN(n14843) );
  XNOR2_X1 U18192 ( .A(n15112), .B(n15375), .ZN(n14842) );
  XNOR2_X1 U18193 ( .A(n14845), .B(n15094), .ZN(n14848) );
  XNOR2_X1 U18194 ( .A(n14846), .B(n3062), .ZN(n14847) );
  XNOR2_X1 U18195 ( .A(n14848), .B(n14847), .ZN(n14856) );
  MUX2_X1 U18196 ( .A(n24572), .B(n14850), .S(n14849), .Z(n14853) );
  XNOR2_X1 U18197 ( .A(n15451), .B(n15369), .ZN(n14854) );
  XNOR2_X1 U18198 ( .A(n14854), .B(n15367), .ZN(n14855) );
  XNOR2_X1 U18199 ( .A(n15169), .B(n1864), .ZN(n14859) );
  XNOR2_X1 U18200 ( .A(n15160), .B(n14859), .ZN(n14863) );
  INV_X1 U18201 ( .A(n14860), .ZN(n14861) );
  XNOR2_X1 U18202 ( .A(n15431), .B(n15103), .ZN(n14895) );
  XNOR2_X1 U18203 ( .A(n14861), .B(n14895), .ZN(n14862) );
  NAND2_X1 U18204 ( .A1(n14864), .A2(n16458), .ZN(n14888) );
  XNOR2_X1 U18206 ( .A(n14477), .B(n14865), .ZN(n14866) );
  XNOR2_X1 U18207 ( .A(n14867), .B(n14866), .ZN(n14872) );
  XNOR2_X1 U18208 ( .A(n14868), .B(n24502), .ZN(n14870) );
  XNOR2_X1 U18209 ( .A(n15210), .B(n1855), .ZN(n14869) );
  XNOR2_X1 U18210 ( .A(n14870), .B(n14869), .ZN(n14871) );
  INV_X1 U18211 ( .A(n14873), .ZN(n14874) );
  XNOR2_X1 U18212 ( .A(n14874), .B(n15392), .ZN(n14878) );
  XNOR2_X1 U18213 ( .A(n15063), .B(n15133), .ZN(n14876) );
  XNOR2_X1 U18214 ( .A(n15120), .B(n925), .ZN(n14875) );
  XNOR2_X1 U18215 ( .A(n14876), .B(n14875), .ZN(n14877) );
  XNOR2_X1 U18216 ( .A(n14881), .B(n15415), .ZN(n14883) );
  XNOR2_X1 U18217 ( .A(n14889), .B(n15174), .ZN(n14882) );
  XNOR2_X1 U18218 ( .A(n14883), .B(n14882), .ZN(n14886) );
  INV_X1 U18219 ( .A(n14884), .ZN(n14885) );
  INV_X1 U18220 ( .A(n17608), .ZN(n16940) );
  INV_X1 U18221 ( .A(n15084), .ZN(n14890) );
  XNOR2_X1 U18222 ( .A(n14892), .B(n15175), .ZN(n14894) );
  XNOR2_X1 U18223 ( .A(n15476), .B(n2743), .ZN(n14893) );
  XNOR2_X1 U18224 ( .A(n14895), .B(n14896), .ZN(n14899) );
  XNOR2_X1 U18225 ( .A(n14900), .B(n853), .ZN(n14901) );
  XNOR2_X1 U18226 ( .A(n14902), .B(n15194), .ZN(n14903) );
  INV_X1 U18227 ( .A(n15514), .ZN(n14904) );
  XNOR2_X1 U18228 ( .A(n14906), .B(n14905), .ZN(n14926) );
  INV_X1 U18229 ( .A(n14926), .ZN(n15572) );
  XNOR2_X1 U18230 ( .A(n14907), .B(n887), .ZN(n14908) );
  XNOR2_X1 U18231 ( .A(n14908), .B(n15095), .ZN(n14910) );
  XNOR2_X1 U18232 ( .A(n14909), .B(n14910), .ZN(n14914) );
  XNOR2_X1 U18233 ( .A(n14912), .B(n14911), .ZN(n14913) );
  XNOR2_X1 U18234 ( .A(n14914), .B(n14913), .ZN(n16028) );
  AOI22_X1 U18235 ( .A1(n16274), .A2(n16029), .B1(n15572), .B2(n16028), .ZN(
        n16280) );
  XNOR2_X1 U18236 ( .A(n15463), .B(n15321), .ZN(n14916) );
  XNOR2_X1 U18237 ( .A(n15120), .B(n2241), .ZN(n14917) );
  XNOR2_X1 U18238 ( .A(n14917), .B(n15495), .ZN(n14918) );
  XNOR2_X1 U18239 ( .A(n14477), .B(n14919), .ZN(n14921) );
  XNOR2_X1 U18240 ( .A(n14920), .B(n14921), .ZN(n14925) );
  XNOR2_X1 U18241 ( .A(n14980), .B(n25013), .ZN(n15090) );
  XNOR2_X1 U18242 ( .A(n15488), .B(n1745), .ZN(n14923) );
  XNOR2_X1 U18243 ( .A(n15090), .B(n14923), .ZN(n14924) );
  XNOR2_X1 U18244 ( .A(n14925), .B(n14924), .ZN(n15573) );
  OAI21_X1 U18246 ( .B1(n24403), .B2(n16277), .A(n16028), .ZN(n14927) );
  MUX2_X1 U18247 ( .A(n17607), .B(n16940), .S(n17615), .Z(n15026) );
  XNOR2_X1 U18248 ( .A(n14928), .B(n15387), .ZN(n14931) );
  INV_X1 U18249 ( .A(n14929), .ZN(n14930) );
  XNOR2_X1 U18250 ( .A(n14930), .B(n14931), .ZN(n14935) );
  XNOR2_X1 U18251 ( .A(n15486), .B(n2208), .ZN(n14932) );
  XNOR2_X1 U18252 ( .A(n14933), .B(n14932), .ZN(n14934) );
  XNOR2_X1 U18253 ( .A(n14935), .B(n14934), .ZN(n14970) );
  XNOR2_X1 U18254 ( .A(n15378), .B(n14936), .ZN(n15306) );
  XNOR2_X1 U18255 ( .A(n14937), .B(n15306), .ZN(n14942) );
  INV_X1 U18256 ( .A(n14993), .ZN(n14938) );
  XNOR2_X1 U18257 ( .A(n14938), .B(n3115), .ZN(n14939) );
  XNOR2_X1 U18258 ( .A(n14939), .B(n14940), .ZN(n14941) );
  NOR2_X1 U18260 ( .A1(n16448), .A2(n16447), .ZN(n14963) );
  MUX2_X1 U18262 ( .A(n14948), .B(n14947), .S(n14946), .Z(n14951) );
  XNOR2_X1 U18263 ( .A(n14952), .B(n15494), .ZN(n14953) );
  XNOR2_X1 U18264 ( .A(n15201), .B(n14953), .ZN(n14957) );
  XNOR2_X1 U18265 ( .A(n15275), .B(n1757), .ZN(n14954) );
  XNOR2_X1 U18266 ( .A(n14954), .B(n14955), .ZN(n14956) );
  XNOR2_X1 U18267 ( .A(n14956), .B(n14957), .ZN(n16452) );
  INV_X1 U18268 ( .A(n14958), .ZN(n14959) );
  XNOR2_X1 U18269 ( .A(n14959), .B(n14960), .ZN(n15296) );
  XNOR2_X1 U18270 ( .A(n15071), .B(n3129), .ZN(n14962) );
  AOI22_X1 U18271 ( .A1(n14963), .A2(n16452), .B1(n223), .B2(n16448), .ZN(
        n14975) );
  XNOR2_X1 U18272 ( .A(n14965), .B(n14964), .ZN(n14969) );
  XNOR2_X1 U18273 ( .A(n15282), .B(n15003), .ZN(n14967) );
  XNOR2_X1 U18274 ( .A(n14967), .B(n14966), .ZN(n14968) );
  XNOR2_X1 U18275 ( .A(n15521), .B(n23476), .ZN(n14971) );
  INV_X1 U18276 ( .A(n17409), .ZN(n17255) );
  XNOR2_X1 U18279 ( .A(n15486), .B(n15387), .ZN(n14983) );
  XNOR2_X1 U18280 ( .A(n14983), .B(n1359), .ZN(n14984) );
  INV_X1 U18281 ( .A(n15774), .ZN(n16303) );
  XNOR2_X1 U18282 ( .A(n14986), .B(n14987), .ZN(n14991) );
  XNOR2_X1 U18283 ( .A(n14988), .B(n21204), .ZN(n14989) );
  XNOR2_X1 U18284 ( .A(n15252), .B(n14989), .ZN(n14990) );
  INV_X1 U18285 ( .A(n16022), .ZN(n16224) );
  XNOR2_X1 U18286 ( .A(n14993), .B(n25416), .ZN(n15032) );
  INV_X1 U18287 ( .A(n15032), .ZN(n14995) );
  INV_X1 U18288 ( .A(n15246), .ZN(n14994) );
  XNOR2_X1 U18290 ( .A(n15109), .B(n14996), .ZN(n14999) );
  XNOR2_X1 U18291 ( .A(n14997), .B(n663), .ZN(n14998) );
  XNOR2_X1 U18292 ( .A(n14999), .B(n14998), .ZN(n15000) );
  XNOR2_X1 U18293 ( .A(n15422), .B(n15003), .ZN(n15039) );
  XNOR2_X1 U18294 ( .A(n15039), .B(n15004), .ZN(n15008) );
  XNOR2_X1 U18295 ( .A(n1351), .B(n2747), .ZN(n15006) );
  XNOR2_X1 U18296 ( .A(n15225), .B(n15006), .ZN(n15007) );
  OAI21_X1 U18297 ( .B1(n16224), .B2(n16225), .A(n16226), .ZN(n15024) );
  XNOR2_X1 U18298 ( .A(n15056), .B(n2735), .ZN(n15009) );
  XNOR2_X1 U18299 ( .A(n15010), .B(n15009), .ZN(n15014) );
  XNOR2_X1 U18300 ( .A(n15012), .B(n15011), .ZN(n15013) );
  INV_X1 U18301 ( .A(n16226), .ZN(n15773) );
  XNOR2_X1 U18302 ( .A(n25443), .B(n1810), .ZN(n15015) );
  XNOR2_X1 U18303 ( .A(n15015), .B(n15321), .ZN(n15017) );
  XNOR2_X1 U18304 ( .A(n15017), .B(n15016), .ZN(n15021) );
  XNOR2_X1 U18305 ( .A(n15062), .B(n25426), .ZN(n15018) );
  XNOR2_X1 U18306 ( .A(n15019), .B(n15018), .ZN(n15020) );
  XNOR2_X1 U18307 ( .A(n18251), .B(n18326), .ZN(n17897) );
  XNOR2_X1 U18308 ( .A(n17897), .B(n18323), .ZN(n15555) );
  XNOR2_X1 U18309 ( .A(n15486), .B(n20825), .ZN(n15027) );
  XNOR2_X1 U18310 ( .A(n15028), .B(n15027), .ZN(n15031) );
  XNOR2_X1 U18311 ( .A(n15029), .B(n15438), .ZN(n15030) );
  XNOR2_X1 U18312 ( .A(n15032), .B(n15447), .ZN(n15038) );
  XNOR2_X1 U18313 ( .A(n24976), .B(n15033), .ZN(n15036) );
  XNOR2_X1 U18314 ( .A(n15034), .B(n886), .ZN(n15035) );
  XNOR2_X1 U18315 ( .A(n15036), .B(n15035), .ZN(n15037) );
  XNOR2_X1 U18316 ( .A(n15038), .B(n15037), .ZN(n16341) );
  INV_X1 U18317 ( .A(n16341), .ZN(n16285) );
  XNOR2_X1 U18318 ( .A(n15420), .B(n15039), .ZN(n15050) );
  XNOR2_X1 U18319 ( .A(n24938), .B(n15284), .ZN(n15048) );
  INV_X1 U18320 ( .A(n15044), .ZN(n15042) );
  INV_X1 U18321 ( .A(n15043), .ZN(n15041) );
  OAI21_X1 U18322 ( .B1(n15042), .B2(n15041), .A(n21079), .ZN(n15046) );
  NAND3_X1 U18323 ( .A1(n15044), .A2(n2991), .A3(n15043), .ZN(n15045) );
  NAND2_X1 U18324 ( .A1(n15046), .A2(n15045), .ZN(n15047) );
  XNOR2_X1 U18325 ( .A(n15048), .B(n15047), .ZN(n15049) );
  XNOR2_X1 U18327 ( .A(n15521), .B(n15051), .ZN(n15053) );
  INV_X1 U18328 ( .A(n15429), .ZN(n15052) );
  XNOR2_X1 U18329 ( .A(n15052), .B(n15053), .ZN(n15060) );
  XNOR2_X1 U18330 ( .A(n15054), .B(n2757), .ZN(n15058) );
  XNOR2_X1 U18331 ( .A(n15055), .B(n15056), .ZN(n15057) );
  XNOR2_X1 U18332 ( .A(n15058), .B(n15057), .ZN(n15059) );
  NAND2_X1 U18335 ( .A1(n1654), .A2(n16341), .ZN(n15061) );
  XNOR2_X1 U18336 ( .A(n15494), .B(n15318), .ZN(n15065) );
  XNOR2_X1 U18337 ( .A(n15063), .B(n15062), .ZN(n15064) );
  XNOR2_X1 U18338 ( .A(n15065), .B(n15064), .ZN(n15068) );
  XNOR2_X1 U18339 ( .A(n15274), .B(n688), .ZN(n15066) );
  XNOR2_X1 U18340 ( .A(n15461), .B(n15066), .ZN(n15067) );
  XNOR2_X1 U18341 ( .A(n15067), .B(n15068), .ZN(n16345) );
  NAND3_X1 U18342 ( .A1(n16345), .A2(n25441), .A3(n24539), .ZN(n15080) );
  XNOR2_X1 U18343 ( .A(n15069), .B(n15070), .ZN(n15078) );
  INV_X1 U18344 ( .A(n15071), .ZN(n15073) );
  INV_X1 U18345 ( .A(n15298), .ZN(n15072) );
  XNOR2_X1 U18346 ( .A(n15074), .B(n1826), .ZN(n15075) );
  NAND3_X1 U18348 ( .A1(n16342), .A2(n1122), .A3(n1654), .ZN(n15079) );
  XNOR2_X1 U18349 ( .A(n15081), .B(n15331), .ZN(n15086) );
  XNOR2_X1 U18350 ( .A(n15082), .B(n20609), .ZN(n15083) );
  XNOR2_X1 U18351 ( .A(n15084), .B(n15083), .ZN(n15085) );
  XNOR2_X1 U18352 ( .A(n15087), .B(n15339), .ZN(n15092) );
  XNOR2_X1 U18353 ( .A(n15088), .B(n677), .ZN(n15089) );
  XNOR2_X1 U18354 ( .A(n15090), .B(n15089), .ZN(n15091) );
  XNOR2_X1 U18355 ( .A(n15092), .B(n15091), .ZN(n16355) );
  XNOR2_X1 U18356 ( .A(n15093), .B(n15356), .ZN(n15101) );
  XNOR2_X1 U18357 ( .A(n15094), .B(n2477), .ZN(n15096) );
  INV_X1 U18358 ( .A(n15097), .ZN(n15098) );
  INV_X1 U18359 ( .A(n16359), .ZN(n16293) );
  INV_X1 U18360 ( .A(n15102), .ZN(n15105) );
  XNOR2_X1 U18361 ( .A(n15103), .B(n16574), .ZN(n15104) );
  XNOR2_X1 U18362 ( .A(n15105), .B(n15104), .ZN(n15108) );
  XNOR2_X1 U18363 ( .A(n15325), .B(n15106), .ZN(n15107) );
  NOR2_X1 U18366 ( .A1(n16293), .A2(n3451), .ZN(n15118) );
  XNOR2_X1 U18368 ( .A(n15109), .B(n92), .ZN(n15110) );
  XNOR2_X1 U18369 ( .A(n15110), .B(n15351), .ZN(n15116) );
  XNOR2_X1 U18370 ( .A(n15113), .B(n15114), .ZN(n15115) );
  NOR2_X1 U18371 ( .A1(n16359), .A2(n16360), .ZN(n15117) );
  XNOR2_X1 U18372 ( .A(n15119), .B(n21046), .ZN(n15122) );
  INV_X1 U18373 ( .A(n15120), .ZN(n15121) );
  XNOR2_X1 U18374 ( .A(n15122), .B(n15121), .ZN(n15125) );
  INV_X1 U18375 ( .A(n15123), .ZN(n15124) );
  XNOR2_X1 U18376 ( .A(n15125), .B(n15124), .ZN(n15128) );
  XNOR2_X1 U18377 ( .A(n15319), .B(n15321), .ZN(n15127) );
  XNOR2_X1 U18378 ( .A(n15128), .B(n15127), .ZN(n16357) );
  INV_X1 U18379 ( .A(n16357), .ZN(n15894) );
  NOR2_X1 U18380 ( .A1(n15894), .A2(n24456), .ZN(n15129) );
  NAND2_X1 U18381 ( .A1(n15129), .A2(n16290), .ZN(n15130) );
  INV_X1 U18382 ( .A(n15131), .ZN(n15132) );
  XNOR2_X1 U18383 ( .A(n15132), .B(n15271), .ZN(n15137) );
  XNOR2_X1 U18384 ( .A(n15133), .B(n13873), .ZN(n15135) );
  XNOR2_X1 U18385 ( .A(n15497), .B(n899), .ZN(n15134) );
  XNOR2_X1 U18386 ( .A(n15135), .B(n15134), .ZN(n15136) );
  INV_X1 U18387 ( .A(n15139), .ZN(n15140) );
  XNOR2_X1 U18388 ( .A(n15280), .B(n15141), .ZN(n15145) );
  XNOR2_X1 U18389 ( .A(n15415), .B(n22886), .ZN(n15143) );
  XNOR2_X1 U18390 ( .A(n15178), .B(n24966), .ZN(n15404) );
  XNOR2_X1 U18391 ( .A(n15404), .B(n15143), .ZN(n15144) );
  INV_X1 U18392 ( .A(n16266), .ZN(n15146) );
  MUX2_X1 U18393 ( .A(n16001), .B(n24366), .S(n15146), .Z(n15163) );
  INV_X1 U18394 ( .A(n15147), .ZN(n15148) );
  XNOR2_X1 U18395 ( .A(n15148), .B(n15297), .ZN(n15152) );
  XNOR2_X1 U18396 ( .A(n15183), .B(n1804), .ZN(n15149) );
  XNOR2_X1 U18397 ( .A(n15150), .B(n15149), .ZN(n15151) );
  XNOR2_X1 U18398 ( .A(n15152), .B(n15151), .ZN(n16002) );
  INV_X1 U18399 ( .A(n16002), .ZN(n16269) );
  XNOR2_X1 U18400 ( .A(n15153), .B(n16), .ZN(n15154) );
  XNOR2_X1 U18401 ( .A(n15155), .B(n15154), .ZN(n15158) );
  XNOR2_X1 U18402 ( .A(n15156), .B(n4556), .ZN(n15157) );
  XNOR2_X1 U18403 ( .A(n15410), .B(n2746), .ZN(n15161) );
  MUX2_X1 U18404 ( .A(n17424), .B(n17381), .S(n17379), .Z(n15261) );
  NAND2_X1 U18405 ( .A1(n15573), .A2(n16028), .ZN(n15771) );
  XNOR2_X1 U18407 ( .A(n15165), .B(n2058), .ZN(n15166) );
  XNOR2_X1 U18408 ( .A(n15167), .B(n15166), .ZN(n15173) );
  XNOR2_X1 U18409 ( .A(n15168), .B(n15169), .ZN(n15171) );
  XNOR2_X1 U18410 ( .A(n15170), .B(n15171), .ZN(n15172) );
  XNOR2_X1 U18411 ( .A(n15172), .B(n15173), .ZN(n16008) );
  XNOR2_X1 U18412 ( .A(n15175), .B(n15174), .ZN(n15226) );
  XNOR2_X1 U18413 ( .A(n15176), .B(n15226), .ZN(n15182) );
  XNOR2_X1 U18414 ( .A(n15177), .B(n15401), .ZN(n15180) );
  XNOR2_X1 U18415 ( .A(n15178), .B(n2036), .ZN(n15179) );
  XNOR2_X1 U18416 ( .A(n15180), .B(n15179), .ZN(n15181) );
  NAND2_X1 U18417 ( .A1(n3554), .A2(n16311), .ZN(n16638) );
  INV_X1 U18418 ( .A(n16638), .ZN(n15216) );
  XNOR2_X1 U18419 ( .A(n15185), .B(n15186), .ZN(n15189) );
  XNOR2_X1 U18420 ( .A(n15369), .B(n15187), .ZN(n15251) );
  XNOR2_X1 U18421 ( .A(n15191), .B(n15190), .ZN(n15193) );
  XNOR2_X1 U18422 ( .A(n14579), .B(n2744), .ZN(n15192) );
  XNOR2_X1 U18423 ( .A(n15193), .B(n15192), .ZN(n15197) );
  XNOR2_X1 U18424 ( .A(n15375), .B(n15194), .ZN(n15248) );
  XNOR2_X1 U18425 ( .A(n15248), .B(n15195), .ZN(n15196) );
  XNOR2_X1 U18426 ( .A(n15196), .B(n15197), .ZN(n15556) );
  AND2_X1 U18427 ( .A1(n15767), .A2(n24297), .ZN(n15215) );
  XNOR2_X1 U18428 ( .A(n15200), .B(n15199), .ZN(n15202) );
  XNOR2_X1 U18429 ( .A(n15201), .B(n15202), .ZN(n15207) );
  INV_X1 U18430 ( .A(n15203), .ZN(n15465) );
  XNOR2_X1 U18431 ( .A(n15465), .B(n2726), .ZN(n15205) );
  XNOR2_X1 U18432 ( .A(n25436), .B(n15204), .ZN(n15217) );
  XNOR2_X1 U18433 ( .A(n15205), .B(n15217), .ZN(n15206) );
  XNOR2_X1 U18435 ( .A(n15209), .B(n15208), .ZN(n15214) );
  XNOR2_X1 U18436 ( .A(n15487), .B(n1758), .ZN(n15212) );
  XNOR2_X1 U18437 ( .A(n15386), .B(n15210), .ZN(n15211) );
  XNOR2_X1 U18438 ( .A(n15212), .B(n15211), .ZN(n15213) );
  NAND2_X1 U18439 ( .A1(n16945), .A2(n17424), .ZN(n17378) );
  NAND2_X1 U18440 ( .A1(n16644), .A2(n17378), .ZN(n15260) );
  XNOR2_X1 U18441 ( .A(n15218), .B(n15217), .ZN(n15222) );
  XNOR2_X1 U18442 ( .A(n15219), .B(n2222), .ZN(n15220) );
  XNOR2_X1 U18443 ( .A(n15499), .B(n15220), .ZN(n15221) );
  XNOR2_X1 U18444 ( .A(n15223), .B(n3093), .ZN(n15224) );
  XNOR2_X1 U18445 ( .A(n15482), .B(n15224), .ZN(n15228) );
  XNOR2_X1 U18446 ( .A(n15225), .B(n15226), .ZN(n15227) );
  INV_X1 U18447 ( .A(n15229), .ZN(n15520) );
  XNOR2_X1 U18448 ( .A(n15230), .B(n15520), .ZN(n15233) );
  XNOR2_X1 U18449 ( .A(n2765), .B(n15409), .ZN(n15232) );
  XNOR2_X1 U18450 ( .A(n15233), .B(n15232), .ZN(n15237) );
  XNOR2_X1 U18451 ( .A(n25384), .B(n15326), .ZN(n15235) );
  XNOR2_X1 U18452 ( .A(n15165), .B(n23699), .ZN(n15234) );
  XNOR2_X1 U18453 ( .A(n15235), .B(n15234), .ZN(n15236) );
  INV_X1 U18454 ( .A(n15674), .ZN(n16197) );
  XNOR2_X1 U18455 ( .A(n15387), .B(n768), .ZN(n15240) );
  XNOR2_X1 U18456 ( .A(n15241), .B(n15240), .ZN(n15242) );
  INV_X1 U18457 ( .A(n16324), .ZN(n15742) );
  XNOR2_X1 U18458 ( .A(n15244), .B(n2739), .ZN(n15245) );
  XNOR2_X1 U18459 ( .A(n15246), .B(n15245), .ZN(n15250) );
  XNOR2_X1 U18460 ( .A(n15248), .B(n15247), .ZN(n15249) );
  XNOR2_X1 U18461 ( .A(n15249), .B(n15250), .ZN(n16323) );
  INV_X1 U18462 ( .A(n16323), .ZN(n16193) );
  XNOR2_X1 U18463 ( .A(n15251), .B(n15503), .ZN(n15257) );
  AND2_X1 U18468 ( .A1(n15262), .A2(n16043), .ZN(n15263) );
  OAI21_X1 U18469 ( .B1(n15263), .B2(n15789), .A(n24430), .ZN(n15265) );
  INV_X1 U18470 ( .A(n15270), .ZN(n15272) );
  XNOR2_X1 U18471 ( .A(n15272), .B(n15271), .ZN(n15279) );
  XNOR2_X1 U18472 ( .A(n15273), .B(n888), .ZN(n15277) );
  XNOR2_X1 U18473 ( .A(n25426), .B(n15274), .ZN(n15276) );
  XNOR2_X1 U18474 ( .A(n15277), .B(n15276), .ZN(n15278) );
  XNOR2_X1 U18475 ( .A(n15280), .B(n15281), .ZN(n15289) );
  INV_X1 U18476 ( .A(n15282), .ZN(n15283) );
  XNOR2_X1 U18477 ( .A(n15284), .B(n15283), .ZN(n15287) );
  XNOR2_X1 U18478 ( .A(n15285), .B(n681), .ZN(n15286) );
  XNOR2_X1 U18479 ( .A(n15287), .B(n15286), .ZN(n15288) );
  XNOR2_X1 U18480 ( .A(n15290), .B(n15291), .ZN(n15295) );
  XNOR2_X1 U18481 ( .A(n15387), .B(n1364), .ZN(n15292) );
  XNOR2_X1 U18482 ( .A(n15293), .B(n15292), .ZN(n15294) );
  XNOR2_X1 U18483 ( .A(n15295), .B(n15294), .ZN(n15706) );
  XNOR2_X1 U18484 ( .A(n15296), .B(n15297), .ZN(n15302) );
  XNOR2_X1 U18485 ( .A(n15298), .B(n2044), .ZN(n15300) );
  XNOR2_X1 U18486 ( .A(n15300), .B(n15299), .ZN(n15301) );
  XNOR2_X1 U18487 ( .A(n15302), .B(n15301), .ZN(n15605) );
  NAND3_X1 U18488 ( .A1(n294), .A2(n4541), .A3(n15605), .ZN(n15310) );
  XNOR2_X1 U18489 ( .A(n24975), .B(n3118), .ZN(n15305) );
  XNOR2_X1 U18490 ( .A(n15306), .B(n15305), .ZN(n15307) );
  NOR2_X1 U18491 ( .A1(n17342), .A2(n17241), .ZN(n17202) );
  NAND3_X1 U18493 ( .A1(n15802), .A2(n15799), .A3(n16076), .ZN(n15311) );
  XNOR2_X1 U18494 ( .A(n15316), .B(n2042), .ZN(n15317) );
  XNOR2_X1 U18496 ( .A(n15465), .B(n15497), .ZN(n15322) );
  XNOR2_X1 U18497 ( .A(n15322), .B(n15321), .ZN(n15323) );
  XNOR2_X1 U18498 ( .A(n15324), .B(n15325), .ZN(n15330) );
  XNOR2_X1 U18499 ( .A(n15168), .B(n15326), .ZN(n15328) );
  XNOR2_X1 U18500 ( .A(n15526), .B(n5131), .ZN(n15327) );
  XNOR2_X1 U18501 ( .A(n15328), .B(n15327), .ZN(n15329) );
  XNOR2_X1 U18502 ( .A(n15330), .B(n15329), .ZN(n15696) );
  XNOR2_X1 U18503 ( .A(n15332), .B(n15331), .ZN(n15337) );
  XNOR2_X1 U18504 ( .A(n15416), .B(n25019), .ZN(n15335) );
  XNOR2_X1 U18505 ( .A(n15333), .B(n2031), .ZN(n15334) );
  XNOR2_X1 U18506 ( .A(n15334), .B(n15335), .ZN(n15336) );
  OAI21_X1 U18507 ( .B1(n15695), .B2(n15696), .A(n25238), .ZN(n15952) );
  INV_X1 U18508 ( .A(n25237), .ZN(n16484) );
  INV_X1 U18509 ( .A(n15338), .ZN(n15340) );
  XNOR2_X1 U18510 ( .A(n15340), .B(n15339), .ZN(n15346) );
  XNOR2_X1 U18511 ( .A(n15342), .B(n15341), .ZN(n15344) );
  XNOR2_X1 U18512 ( .A(n15483), .B(n3084), .ZN(n15343) );
  XNOR2_X1 U18513 ( .A(n15344), .B(n15343), .ZN(n15345) );
  XNOR2_X1 U18514 ( .A(n15349), .B(n15348), .ZN(n15354) );
  XNOR2_X1 U18515 ( .A(n15350), .B(n20995), .ZN(n15352) );
  XNOR2_X1 U18516 ( .A(n15354), .B(n15353), .ZN(n16480) );
  XNOR2_X1 U18517 ( .A(n15356), .B(n15355), .ZN(n15363) );
  XNOR2_X1 U18518 ( .A(n15359), .B(n2087), .ZN(n15360) );
  XNOR2_X1 U18519 ( .A(n15361), .B(n15360), .ZN(n15362) );
  XNOR2_X1 U18520 ( .A(n15363), .B(n15362), .ZN(n16481) );
  INV_X1 U18521 ( .A(n15695), .ZN(n15364) );
  NAND3_X1 U18522 ( .A1(n15364), .A2(n16480), .A3(n16481), .ZN(n15365) );
  XNOR2_X1 U18523 ( .A(n15366), .B(n15367), .ZN(n15373) );
  INV_X1 U18524 ( .A(n15368), .ZN(n15371) );
  XNOR2_X1 U18525 ( .A(n15369), .B(n17960), .ZN(n15370) );
  XNOR2_X1 U18526 ( .A(n15371), .B(n15370), .ZN(n15372) );
  XNOR2_X1 U18527 ( .A(n15375), .B(n15514), .ZN(n15376) );
  XNOR2_X1 U18528 ( .A(n15376), .B(n15377), .ZN(n15382) );
  XNOR2_X1 U18529 ( .A(n25501), .B(n14579), .ZN(n15380) );
  XNOR2_X1 U18530 ( .A(n15378), .B(n23271), .ZN(n15379) );
  XNOR2_X1 U18531 ( .A(n15380), .B(n15379), .ZN(n15381) );
  INV_X1 U18532 ( .A(n15383), .ZN(n15384) );
  XNOR2_X1 U18533 ( .A(n15385), .B(n15384), .ZN(n15391) );
  XNOR2_X1 U18534 ( .A(n15484), .B(n15386), .ZN(n15389) );
  XNOR2_X1 U18535 ( .A(n15387), .B(n2034), .ZN(n15388) );
  XNOR2_X1 U18536 ( .A(n15389), .B(n15388), .ZN(n15390) );
  XNOR2_X2 U18537 ( .A(n15391), .B(n15390), .ZN(n16064) );
  INV_X1 U18538 ( .A(n16064), .ZN(n15550) );
  INV_X1 U18539 ( .A(n15392), .ZN(n15395) );
  INV_X1 U18540 ( .A(n15393), .ZN(n15498) );
  XNOR2_X1 U18541 ( .A(n15498), .B(n13873), .ZN(n15394) );
  XNOR2_X1 U18542 ( .A(n15395), .B(n15394), .ZN(n15400) );
  XNOR2_X1 U18543 ( .A(n15396), .B(n1827), .ZN(n15397) );
  XNOR2_X1 U18544 ( .A(n15398), .B(n15397), .ZN(n15399) );
  XNOR2_X1 U18545 ( .A(n15478), .B(n2782), .ZN(n15402) );
  XNOR2_X1 U18546 ( .A(n15405), .B(n15406), .ZN(n15549) );
  XNOR2_X1 U18547 ( .A(n15407), .B(n15408), .ZN(n15414) );
  XNOR2_X1 U18548 ( .A(n15409), .B(n24423), .ZN(n15412) );
  XNOR2_X1 U18549 ( .A(n15412), .B(n15411), .ZN(n15413) );
  XNOR2_X1 U18550 ( .A(n15414), .B(n15413), .ZN(n15548) );
  NOR2_X1 U18551 ( .A1(n17341), .A2(n17346), .ZN(n17235) );
  XNOR2_X1 U18552 ( .A(n15416), .B(n15415), .ZN(n15419) );
  XNOR2_X1 U18553 ( .A(n15417), .B(n2190), .ZN(n15418) );
  XNOR2_X1 U18554 ( .A(n15419), .B(n15418), .ZN(n15426) );
  INV_X1 U18555 ( .A(n15420), .ZN(n15424) );
  XNOR2_X1 U18556 ( .A(n15422), .B(n15421), .ZN(n15423) );
  XNOR2_X1 U18557 ( .A(n15424), .B(n15423), .ZN(n15425) );
  XNOR2_X1 U18558 ( .A(n15425), .B(n15426), .ZN(n15715) );
  INV_X1 U18559 ( .A(n15427), .ZN(n15428) );
  XNOR2_X1 U18560 ( .A(n15428), .B(n15429), .ZN(n15435) );
  XNOR2_X1 U18561 ( .A(n15430), .B(n3183), .ZN(n15433) );
  XNOR2_X1 U18562 ( .A(n15168), .B(n15431), .ZN(n15432) );
  XNOR2_X1 U18563 ( .A(n15433), .B(n15432), .ZN(n15434) );
  XNOR2_X1 U18564 ( .A(n15436), .B(n187), .ZN(n15437) );
  XNOR2_X1 U18565 ( .A(n14477), .B(n15437), .ZN(n15440) );
  INV_X1 U18566 ( .A(n15438), .ZN(n15439) );
  XNOR2_X1 U18567 ( .A(n15440), .B(n15439), .ZN(n15443) );
  INV_X1 U18568 ( .A(n15441), .ZN(n15442) );
  XNOR2_X1 U18569 ( .A(n15444), .B(n2970), .ZN(n15445) );
  XNOR2_X1 U18570 ( .A(n15445), .B(n15446), .ZN(n15448) );
  XNOR2_X1 U18571 ( .A(n15448), .B(n15447), .ZN(n15450) );
  NAND2_X1 U18572 ( .A1(n16474), .A2(n24550), .ZN(n15459) );
  XNOR2_X1 U18573 ( .A(n15451), .B(n1875), .ZN(n15453) );
  XNOR2_X1 U18574 ( .A(n15453), .B(n15452), .ZN(n15455) );
  XNOR2_X1 U18575 ( .A(n15454), .B(n15455), .ZN(n15458) );
  INV_X1 U18576 ( .A(n15456), .ZN(n15457) );
  XNOR2_X1 U18577 ( .A(n15458), .B(n15457), .ZN(n15714) );
  MUX2_X1 U18578 ( .A(n15460), .B(n15459), .S(n16471), .Z(n17237) );
  XNOR2_X1 U18579 ( .A(n15461), .B(n15462), .ZN(n15469) );
  XNOR2_X1 U18580 ( .A(n15464), .B(n15463), .ZN(n15467) );
  XNOR2_X1 U18581 ( .A(n15465), .B(n2826), .ZN(n15466) );
  XNOR2_X1 U18582 ( .A(n15467), .B(n15466), .ZN(n15468) );
  INV_X1 U18583 ( .A(n16473), .ZN(n16476) );
  NOR2_X1 U18584 ( .A1(n16476), .A2(n16472), .ZN(n15471) );
  NAND2_X1 U18585 ( .A1(n17237), .A2(n3872), .ZN(n16780) );
  NOR2_X1 U18586 ( .A1(n17241), .A2(n17346), .ZN(n15472) );
  XNOR2_X1 U18587 ( .A(n18074), .B(n18523), .ZN(n17987) );
  MUX2_X1 U18588 ( .A(n16484), .B(n24981), .S(n15953), .Z(n15475) );
  NOR2_X1 U18589 ( .A1(n25238), .A2(n16480), .ZN(n15474) );
  INV_X1 U18590 ( .A(n16481), .ZN(n15950) );
  INV_X1 U18591 ( .A(n15872), .ZN(n15534) );
  XNOR2_X1 U18592 ( .A(n15476), .B(n2228), .ZN(n15477) );
  INV_X1 U18593 ( .A(n24956), .ZN(n15479) );
  XNOR2_X1 U18594 ( .A(n15479), .B(n25019), .ZN(n15481) );
  XNOR2_X1 U18595 ( .A(n15484), .B(n15483), .ZN(n15485) );
  XNOR2_X1 U18596 ( .A(n15486), .B(n15487), .ZN(n15490) );
  INV_X1 U18597 ( .A(n2990), .ZN(n23239) );
  XNOR2_X1 U18598 ( .A(n15488), .B(n23239), .ZN(n15489) );
  XNOR2_X1 U18599 ( .A(n15490), .B(n15489), .ZN(n15491) );
  XNOR2_X1 U18600 ( .A(n15492), .B(n15491), .ZN(n15710) );
  INV_X1 U18601 ( .A(n15710), .ZN(n16443) );
  XNOR2_X1 U18602 ( .A(n14384), .B(n21423), .ZN(n15493) );
  XNOR2_X1 U18603 ( .A(n15493), .B(n15494), .ZN(n15496) );
  XNOR2_X1 U18604 ( .A(n15496), .B(n15495), .ZN(n15502) );
  XNOR2_X1 U18605 ( .A(n15498), .B(n15497), .ZN(n15500) );
  XNOR2_X1 U18606 ( .A(n15500), .B(n15499), .ZN(n15501) );
  XNOR2_X1 U18607 ( .A(n15502), .B(n15501), .ZN(n16243) );
  INV_X1 U18608 ( .A(n16243), .ZN(n15943) );
  XNOR2_X1 U18609 ( .A(n15505), .B(n15506), .ZN(n15509) );
  XNOR2_X1 U18610 ( .A(n15507), .B(n21553), .ZN(n15508) );
  XNOR2_X1 U18611 ( .A(n15509), .B(n15508), .ZN(n15510) );
  INV_X1 U18612 ( .A(n16437), .ZN(n15945) );
  XNOR2_X1 U18613 ( .A(n15512), .B(n15513), .ZN(n15519) );
  XNOR2_X1 U18614 ( .A(n25501), .B(n812), .ZN(n15516) );
  XNOR2_X1 U18615 ( .A(n15517), .B(n15516), .ZN(n15518) );
  XNOR2_X1 U18616 ( .A(n25431), .B(n15520), .ZN(n15525) );
  XNOR2_X1 U18617 ( .A(n25384), .B(n15523), .ZN(n15524) );
  XNOR2_X1 U18618 ( .A(n15525), .B(n15524), .ZN(n15530) );
  XNOR2_X1 U18619 ( .A(n15526), .B(n14694), .ZN(n15528) );
  XNOR2_X1 U18620 ( .A(n15165), .B(n1854), .ZN(n15527) );
  XNOR2_X1 U18621 ( .A(n15528), .B(n15527), .ZN(n15529) );
  INV_X1 U18622 ( .A(n15707), .ZN(n15946) );
  NOR2_X1 U18624 ( .A1(n15952), .A2(n15695), .ZN(n15871) );
  NOR2_X1 U18625 ( .A1(n16578), .A2(n15871), .ZN(n15533) );
  NAND2_X1 U18626 ( .A1(n16043), .A2(n15790), .ZN(n15537) );
  INV_X1 U18627 ( .A(n16043), .ZN(n15535) );
  AND2_X1 U18628 ( .A1(n15535), .A2(n16042), .ZN(n15788) );
  NAND2_X1 U18630 ( .A1(n16742), .A2(n15538), .ZN(n16653) );
  INV_X1 U18631 ( .A(n16051), .ZN(n16509) );
  NAND2_X1 U18632 ( .A1(n15691), .A2(n16509), .ZN(n15544) );
  NAND2_X1 U18633 ( .A1(n15539), .A2(n16508), .ZN(n15543) );
  MUX2_X1 U18637 ( .A(n17087), .B(n17086), .S(n16578), .Z(n16647) );
  INV_X1 U18638 ( .A(n15548), .ZN(n16062) );
  INV_X1 U18640 ( .A(n15694), .ZN(n15794) );
  OAI211_X1 U18641 ( .C1(n16062), .C2(n15794), .A(n15550), .B(n16067), .ZN(
        n15551) );
  XNOR2_X1 U18642 ( .A(n18351), .B(n869), .ZN(n15553) );
  XNOR2_X1 U18643 ( .A(n17987), .B(n15553), .ZN(n15554) );
  INV_X1 U18646 ( .A(n17335), .ZN(n15563) );
  MUX2_X1 U18647 ( .A(n16225), .B(n16022), .S(n15774), .Z(n15562) );
  INV_X1 U18649 ( .A(n16917), .ZN(n16727) );
  OAI21_X1 U18650 ( .B1(n16974), .B2(n15563), .A(n16727), .ZN(n15578) );
  OAI21_X1 U18651 ( .B1(n15933), .B2(n16230), .A(n15565), .ZN(n15566) );
  INV_X1 U18652 ( .A(n16491), .ZN(n15937) );
  INV_X1 U18653 ( .A(n16016), .ZN(n16251) );
  AOI21_X1 U18654 ( .B1(n16251), .B2(n16247), .A(n2605), .ZN(n15571) );
  NAND2_X1 U18655 ( .A1(n16247), .A2(n25484), .ZN(n15569) );
  MUX2_X1 U18656 ( .A(n15569), .B(n15568), .S(n16016), .Z(n15570) );
  OAI21_X1 U18657 ( .B1(n15571), .B2(n16018), .A(n15570), .ZN(n17334) );
  OAI21_X1 U18658 ( .B1(n16971), .B2(n25412), .A(n16917), .ZN(n15577) );
  NOR2_X1 U18659 ( .A1(n15573), .A2(n16028), .ZN(n15574) );
  AOI21_X1 U18660 ( .B1(n17335), .B2(n376), .A(n17332), .ZN(n15575) );
  INV_X1 U18661 ( .A(n15579), .ZN(n15581) );
  INV_X1 U18662 ( .A(n25409), .ZN(n16084) );
  NAND2_X1 U18663 ( .A1(n16084), .A2(n16105), .ZN(n15580) );
  NAND2_X1 U18664 ( .A1(n15581), .A2(n15580), .ZN(n15586) );
  INV_X1 U18665 ( .A(n15582), .ZN(n15585) );
  NAND2_X1 U18666 ( .A1(n16038), .A2(n24429), .ZN(n15588) );
  NAND3_X1 U18667 ( .A1(n15789), .A2(n15790), .A3(n24430), .ZN(n15587) );
  OAI21_X1 U18668 ( .B1(n24928), .B2(n16107), .A(n25030), .ZN(n15591) );
  INV_X1 U18669 ( .A(n16107), .ZN(n15783) );
  NAND3_X1 U18671 ( .A1(n24826), .A2(n16077), .A3(n15801), .ZN(n15597) );
  NAND3_X1 U18672 ( .A1(n1365), .A2(n16077), .A3(n16076), .ZN(n15596) );
  NAND2_X1 U18674 ( .A1(n16067), .A2(n16060), .ZN(n15599) );
  INV_X1 U18679 ( .A(n17068), .ZN(n16730) );
  XNOR2_X1 U18680 ( .A(n18262), .B(n18240), .ZN(n17906) );
  NOR2_X1 U18681 ( .A1(n15611), .A2(n14499), .ZN(n15614) );
  NOR2_X1 U18682 ( .A1(n15612), .A2(n15857), .ZN(n15613) );
  NAND3_X1 U18683 ( .A1(n15804), .A2(n16118), .A3(n15857), .ZN(n15615) );
  OAI21_X1 U18684 ( .B1(n16680), .B2(n16117), .A(n15615), .ZN(n15616) );
  INV_X1 U18685 ( .A(n24585), .ZN(n15883) );
  NAND2_X1 U18686 ( .A1(n16125), .A2(n15842), .ZN(n15965) );
  NAND2_X1 U18687 ( .A1(n15965), .A2(n16122), .ZN(n15618) );
  AOI22_X1 U18688 ( .A1(n15620), .A2(n15846), .B1(n15619), .B2(n15618), .ZN(
        n17061) );
  INV_X1 U18689 ( .A(n17061), .ZN(n16929) );
  INV_X1 U18691 ( .A(n16388), .ZN(n16162) );
  NOR2_X1 U18692 ( .A1(n16394), .A2(n16162), .ZN(n15847) );
  NOR2_X1 U18693 ( .A1(n16393), .A2(n15849), .ZN(n15622) );
  OAI21_X1 U18694 ( .B1(n15847), .B2(n15622), .A(n15848), .ZN(n15623) );
  AOI21_X1 U18696 ( .B1(n293), .B2(n15625), .A(n16095), .ZN(n15626) );
  NAND2_X1 U18697 ( .A1(n17059), .A2(n15631), .ZN(n16935) );
  INV_X1 U18698 ( .A(n16935), .ZN(n15634) );
  MUX2_X1 U18699 ( .A(n16082), .B(n15632), .S(n16102), .Z(n15633) );
  NAND2_X1 U18700 ( .A1(n15634), .A2(n17054), .ZN(n15636) );
  NOR2_X1 U18701 ( .A1(n16932), .A2(n24585), .ZN(n15880) );
  NAND2_X1 U18702 ( .A1(n15638), .A2(n15970), .ZN(n16187) );
  NAND2_X1 U18703 ( .A1(n17183), .A2(n15641), .ZN(n15644) );
  NAND2_X1 U18704 ( .A1(n15907), .A2(n16367), .ZN(n15642) );
  NAND3_X1 U18705 ( .A1(n17312), .A2(n17596), .A3(n17597), .ZN(n15664) );
  NAND2_X1 U18707 ( .A1(n16422), .A2(n16427), .ZN(n15648) );
  MUX2_X1 U18708 ( .A(n15649), .B(n15648), .S(n16170), .Z(n15650) );
  AOI21_X1 U18709 ( .B1(n25492), .B2(n16412), .A(n16414), .ZN(n15651) );
  NAND2_X1 U18710 ( .A1(n16417), .A2(n16408), .ZN(n15984) );
  MUX2_X1 U18711 ( .A(n15651), .B(n15984), .S(n16413), .Z(n15652) );
  NOR2_X1 U18712 ( .A1(n17305), .A2(n17316), .ZN(n17600) );
  NAND2_X1 U18713 ( .A1(n2968), .A2(n17600), .ZN(n15663) );
  NAND2_X1 U18715 ( .A1(n16382), .A2(n25210), .ZN(n15654) );
  NOR2_X1 U18717 ( .A1(n4046), .A2(n15837), .ZN(n16385) );
  NAND2_X1 U18718 ( .A1(n16385), .A2(n25210), .ZN(n15658) );
  NAND2_X1 U18719 ( .A1(n17598), .A2(n16921), .ZN(n17315) );
  INV_X1 U18720 ( .A(n17315), .ZN(n15661) );
  NAND2_X1 U18721 ( .A1(n17312), .A2(n15661), .ZN(n15662) );
  NAND3_X1 U18722 ( .A1(n17316), .A2(n24542), .A3(n16921), .ZN(n17601) );
  NAND4_X1 U18723 ( .A1(n15664), .A2(n15663), .A3(n15662), .A4(n17601), .ZN(
        n15665) );
  XNOR2_X1 U18724 ( .A(n15665), .B(n17875), .ZN(n18317) );
  INV_X1 U18725 ( .A(n18317), .ZN(n15666) );
  XNOR2_X1 U18726 ( .A(n15666), .B(n17906), .ZN(n15736) );
  INV_X1 U18727 ( .A(n16331), .ZN(n15755) );
  NAND2_X1 U18728 ( .A1(n15755), .A2(n16332), .ZN(n15668) );
  INV_X1 U18729 ( .A(n16595), .ZN(n15887) );
  INV_X1 U18730 ( .A(n16349), .ZN(n15885) );
  AOI21_X1 U18731 ( .B1(n16597), .B2(n15885), .A(n25432), .ZN(n15672) );
  NAND3_X1 U18732 ( .A1(n17326), .A2(n15673), .A3(n4426), .ZN(n15685) );
  OAI22_X1 U18733 ( .A1(n1122), .A2(n16285), .B1(n24539), .B2(n1654), .ZN(
        n16015) );
  NAND2_X1 U18734 ( .A1(n24540), .A2(n25441), .ZN(n16344) );
  NAND2_X1 U18735 ( .A1(n16015), .A2(n16344), .ZN(n15683) );
  NOR2_X1 U18736 ( .A1(n16345), .A2(n25441), .ZN(n15747) );
  INV_X1 U18737 ( .A(n15747), .ZN(n15681) );
  INV_X1 U18738 ( .A(n15679), .ZN(n15680) );
  NAND2_X1 U18739 ( .A1(n15681), .A2(n15680), .ZN(n15682) );
  NAND3_X1 U18740 ( .A1(n15673), .A2(n17319), .A3(n16607), .ZN(n15684) );
  INV_X1 U18741 ( .A(n16242), .ZN(n15944) );
  NOR2_X1 U18742 ( .A1(n16243), .A2(n15946), .ZN(n16441) );
  NAND2_X1 U18743 ( .A1(n16443), .A2(n15946), .ZN(n15686) );
  OAI21_X1 U18744 ( .B1(n16450), .B2(n16447), .A(n223), .ZN(n15687) );
  MUX2_X1 U18745 ( .A(n24550), .B(n16471), .S(n16469), .Z(n15690) );
  AOI21_X1 U18746 ( .B1(n15715), .B2(n16475), .A(n16472), .ZN(n15689) );
  MUX2_X1 U18748 ( .A(n15953), .B(n16483), .S(n16480), .Z(n16485) );
  INV_X1 U18749 ( .A(n15698), .ZN(n16547) );
  AOI21_X1 U18750 ( .B1(n16547), .B2(n16795), .A(n16550), .ZN(n15701) );
  INV_X1 U18751 ( .A(n16549), .ZN(n15699) );
  NAND2_X1 U18752 ( .A1(n15699), .A2(n16795), .ZN(n15700) );
  XNOR2_X1 U18753 ( .A(n18080), .B(n18539), .ZN(n15734) );
  INV_X1 U18754 ( .A(n16465), .ZN(n16460) );
  AOI21_X1 U18755 ( .B1(n5269), .B2(n16221), .A(n16460), .ZN(n15705) );
  INV_X1 U18756 ( .A(n15921), .ZN(n16459) );
  NOR2_X1 U18757 ( .A1(n15707), .A2(n16242), .ZN(n15708) );
  NAND3_X1 U18759 ( .A1(n16438), .A2(n16437), .A3(n16442), .ZN(n15712) );
  NAND2_X1 U18760 ( .A1(n16616), .A2(n17299), .ZN(n17302) );
  NOR2_X1 U18761 ( .A1(n16705), .A2(n17299), .ZN(n15724) );
  INV_X1 U18762 ( .A(n15714), .ZN(n16057) );
  NOR2_X1 U18764 ( .A1(n16616), .A2(n17297), .ZN(n15723) );
  INV_X1 U18765 ( .A(n16480), .ZN(n15951) );
  NOR2_X1 U18766 ( .A1(n15718), .A2(n15717), .ZN(n15722) );
  NOR2_X1 U18767 ( .A1(n15953), .A2(n15950), .ZN(n15719) );
  NAND2_X1 U18768 ( .A1(n15719), .A2(n24981), .ZN(n15720) );
  OAI21_X1 U18769 ( .B1(n15724), .B2(n15723), .A(n16708), .ZN(n15732) );
  INV_X1 U18770 ( .A(n16451), .ZN(n15725) );
  XNOR2_X1 U18772 ( .A(n18382), .B(n21623), .ZN(n15733) );
  XNOR2_X1 U18773 ( .A(n15734), .B(n15733), .ZN(n15735) );
  NOR2_X1 U18774 ( .A1(n19302), .A2(n19307), .ZN(n19130) );
  NOR2_X1 U18775 ( .A1(n15737), .A2(n16551), .ZN(n15741) );
  NOR2_X2 U18777 ( .A1(n15741), .A2(n15740), .ZN(n18188) );
  INV_X1 U18778 ( .A(n16194), .ZN(n15744) );
  NAND2_X1 U18779 ( .A1(n16356), .A2(n16290), .ZN(n16363) );
  OAI22_X1 U18780 ( .A1(n16363), .A2(n25546), .B1(n15748), .B2(n16290), .ZN(
        n15749) );
  OAI22_X1 U18781 ( .A1(n16309), .A2(n15751), .B1(n16012), .B2(n15750), .ZN(
        n15754) );
  NAND2_X1 U18782 ( .A1(n15557), .A2(n3554), .ZN(n15752) );
  INV_X1 U18783 ( .A(n15757), .ZN(n15759) );
  INV_X1 U18784 ( .A(n16267), .ZN(n15758) );
  NAND2_X1 U18785 ( .A1(n16230), .A2(n16232), .ZN(n16490) );
  NAND2_X1 U18786 ( .A1(n16491), .A2(n15564), .ZN(n16489) );
  NOR2_X1 U18787 ( .A1(n16489), .A2(n16232), .ZN(n15760) );
  NOR2_X1 U18791 ( .A1(n16312), .A2(n15556), .ZN(n16315) );
  INV_X1 U18792 ( .A(n16809), .ZN(n17481) );
  NAND2_X1 U18793 ( .A1(n16030), .A2(n16273), .ZN(n15769) );
  MUX2_X1 U18794 ( .A(n15770), .B(n15769), .S(n16274), .Z(n16810) );
  INV_X1 U18795 ( .A(n15771), .ZN(n15772) );
  NAND2_X1 U18796 ( .A1(n15772), .A2(n16029), .ZN(n16808) );
  INV_X1 U18797 ( .A(n17076), .ZN(n16588) );
  NAND3_X1 U18798 ( .A1(n16302), .A2(n16022), .A3(n16023), .ZN(n15775) );
  NAND3_X1 U18799 ( .A1(n16220), .A2(n15921), .A3(n16221), .ZN(n15778) );
  NAND2_X1 U18800 ( .A1(n5269), .A2(n16465), .ZN(n15777) );
  INV_X1 U18801 ( .A(n15780), .ZN(n15781) );
  NOR2_X1 U18802 ( .A1(n15781), .A2(n16102), .ZN(n15787) );
  MUX2_X1 U18803 ( .A(n4678), .B(n15854), .S(n24586), .Z(n15785) );
  NOR2_X1 U18804 ( .A1(n17134), .A2(n3458), .ZN(n15809) );
  NOR2_X1 U18805 ( .A1(n16038), .A2(n24429), .ZN(n15786) );
  AOI22_X1 U18806 ( .A1(n15788), .A2(n24430), .B1(n15786), .B2(n2251), .ZN(
        n16576) );
  INV_X1 U18807 ( .A(n15787), .ZN(n15793) );
  INV_X1 U18808 ( .A(n15788), .ZN(n15792) );
  AOI21_X1 U18809 ( .B1(n291), .B2(n15790), .A(n15789), .ZN(n15791) );
  NAND3_X1 U18810 ( .A1(n16576), .A2(n15793), .A3(n16575), .ZN(n15797) );
  OAI21_X1 U18811 ( .B1(n15798), .B2(n15797), .A(n17131), .ZN(n15808) );
  NAND2_X1 U18812 ( .A1(n25245), .A2(n17130), .ZN(n15803) );
  XNOR2_X1 U18813 ( .A(n18289), .B(n18301), .ZN(n17911) );
  XNOR2_X1 U18814 ( .A(n15810), .B(n17911), .ZN(n15879) );
  NAND2_X1 U18816 ( .A1(n15814), .A2(n16204), .ZN(n15815) );
  NAND2_X1 U18817 ( .A1(n15905), .A2(n17183), .ZN(n16366) );
  NOR2_X1 U18821 ( .A1(n16170), .A2(n244), .ZN(n15819) );
  NOR2_X1 U18823 ( .A1(n15890), .A2(n24587), .ZN(n15823) );
  OAI21_X1 U18824 ( .B1(n15824), .B2(n15823), .A(n24080), .ZN(n15827) );
  INV_X1 U18825 ( .A(n16427), .ZN(n15825) );
  OAI21_X1 U18826 ( .B1(n16422), .B2(n707), .A(n15825), .ZN(n15826) );
  NAND2_X1 U18827 ( .A1(n15826), .A2(n16170), .ZN(n15836) );
  AND4_X1 U18828 ( .A1(n15835), .A2(n16598), .A3(n15827), .A4(n15836), .ZN(
        n15834) );
  NOR2_X1 U18829 ( .A1(n16188), .A2(n15970), .ZN(n15829) );
  NAND2_X1 U18830 ( .A1(n16400), .A2(n15970), .ZN(n15831) );
  NAND3_X1 U18831 ( .A1(n16188), .A2(n15972), .A3(n16397), .ZN(n15830) );
  NAND2_X1 U18832 ( .A1(n15831), .A2(n15830), .ZN(n15832) );
  INV_X1 U18833 ( .A(n17729), .ZN(n17735) );
  NOR2_X1 U18834 ( .A1(n15837), .A2(n16177), .ZN(n15838) );
  NOR3_X1 U18835 ( .A1(n15839), .A2(n4045), .A3(n15838), .ZN(n15840) );
  MUX2_X1 U18837 ( .A(n15844), .B(n24654), .S(n16122), .Z(n15845) );
  INV_X1 U18838 ( .A(n15847), .ZN(n15853) );
  NOR2_X1 U18839 ( .A1(n16391), .A2(n15849), .ZN(n16390) );
  NAND2_X1 U18840 ( .A1(n15848), .A2(n16162), .ZN(n15851) );
  INV_X1 U18841 ( .A(n15849), .ZN(n16392) );
  AOI22_X2 U18842 ( .A1(n15852), .A2(n15853), .B1(n15851), .B2(n15850), .ZN(
        n17118) );
  INV_X1 U18843 ( .A(n17118), .ZN(n17100) );
  INV_X1 U18844 ( .A(n17120), .ZN(n17115) );
  OAI21_X1 U18845 ( .B1(n890), .B2(n17100), .A(n17115), .ZN(n15870) );
  NOR2_X1 U18846 ( .A1(n16114), .A2(n16118), .ZN(n15859) );
  INV_X1 U18850 ( .A(n15625), .ZN(n16148) );
  NAND2_X1 U18851 ( .A1(n16409), .A2(n16412), .ZN(n15865) );
  NAND2_X1 U18852 ( .A1(n15984), .A2(n16414), .ZN(n15867) );
  NOR3_X1 U18853 ( .A1(n17088), .A2(n17086), .A3(n16578), .ZN(n15874) );
  AOI21_X1 U18854 ( .B1(n15875), .B2(n17087), .A(n15874), .ZN(n15876) );
  XNOR2_X1 U18855 ( .A(n18294), .B(n20744), .ZN(n15877) );
  XNOR2_X1 U18856 ( .A(n18305), .B(n15877), .ZN(n15878) );
  NAND2_X1 U18857 ( .A1(n25031), .A2(n16929), .ZN(n15884) );
  AOI21_X1 U18858 ( .B1(n17060), .B2(n17059), .A(n17054), .ZN(n15881) );
  OAI22_X1 U18859 ( .A1(n15881), .A2(n15880), .B1(n15883), .B2(n17060), .ZN(
        n15882) );
  NAND2_X1 U18860 ( .A1(n15885), .A2(n24467), .ZN(n15886) );
  NAND3_X1 U18861 ( .A1(n15888), .A2(n15886), .A3(n15887), .ZN(n15892) );
  NAND3_X1 U18862 ( .A1(n15890), .A2(n25432), .A3(n24467), .ZN(n15891) );
  NAND2_X1 U18863 ( .A1(n15894), .A2(n16360), .ZN(n15898) );
  NAND3_X1 U18864 ( .A1(n24841), .A2(n24456), .A3(n15894), .ZN(n15896) );
  OAI211_X1 U18865 ( .C1(n24919), .C2(n15898), .A(n15897), .B(n15896), .ZN(
        n16770) );
  AOI21_X1 U18866 ( .B1(n16196), .B2(n16328), .A(n15899), .ZN(n15903) );
  NAND2_X1 U18867 ( .A1(n15901), .A2(n15900), .ZN(n15902) );
  NAND3_X1 U18869 ( .A1(n16368), .A2(n15904), .A3(n16204), .ZN(n15911) );
  NOR2_X1 U18870 ( .A1(n16367), .A2(n16206), .ZN(n15906) );
  NAND2_X1 U18871 ( .A1(n15906), .A2(n17180), .ZN(n15909) );
  NAND3_X1 U18872 ( .A1(n15907), .A2(n17183), .A3(n16367), .ZN(n15908) );
  NAND4_X1 U18873 ( .A1(n15911), .A2(n15910), .A3(n15909), .A4(n15908), .ZN(
        n16989) );
  NAND2_X1 U18874 ( .A1(n16406), .A2(n24061), .ZN(n16402) );
  NAND2_X1 U18875 ( .A1(n15646), .A2(n25500), .ZN(n15912) );
  NAND3_X1 U18876 ( .A1(n16406), .A2(n15646), .A3(n16403), .ZN(n15913) );
  MUX2_X1 U18877 ( .A(n25455), .B(n16334), .S(n1123), .Z(n15914) );
  NAND2_X1 U18878 ( .A1(n15914), .A2(n267), .ZN(n15919) );
  NAND2_X1 U18880 ( .A1(n17364), .A2(n25214), .ZN(n15920) );
  INV_X1 U18881 ( .A(n16989), .ZN(n17362) );
  NOR2_X1 U18882 ( .A1(n16220), .A2(n16221), .ZN(n15924) );
  NOR2_X1 U18883 ( .A1(n15921), .A2(n16219), .ZN(n15923) );
  INV_X1 U18884 ( .A(n15922), .ZN(n16462) );
  MUX2_X1 U18885 ( .A(n15924), .B(n15923), .S(n16462), .Z(n15927) );
  OAI22_X1 U18886 ( .A1(n15925), .A2(n16461), .B1(n16216), .B2(n16465), .ZN(
        n15926) );
  NOR2_X2 U18887 ( .A1(n15927), .A2(n15926), .ZN(n17048) );
  MUX2_X1 U18888 ( .A(n16447), .B(n257), .S(n16449), .Z(n15931) );
  NAND2_X1 U18889 ( .A1(n16235), .A2(n16451), .ZN(n15928) );
  MUX2_X1 U18890 ( .A(n15929), .B(n15928), .S(n16449), .Z(n15930) );
  INV_X1 U18891 ( .A(n16231), .ZN(n16494) );
  INV_X1 U18892 ( .A(n16230), .ZN(n16492) );
  MUX2_X1 U18893 ( .A(n15935), .B(n15934), .S(n16492), .Z(n15936) );
  INV_X1 U18894 ( .A(n15938), .ZN(n16252) );
  NOR2_X1 U18895 ( .A1(n16252), .A2(n15762), .ZN(n15939) );
  AOI22_X1 U18896 ( .A1(n15939), .A2(n16016), .B1(n16246), .B2(n16252), .ZN(
        n15942) );
  INV_X1 U18897 ( .A(n17048), .ZN(n16628) );
  OAI211_X1 U18898 ( .C1(n15943), .C2(n15946), .A(n16438), .B(n16242), .ZN(
        n15949) );
  NAND3_X1 U18899 ( .A1(n16442), .A2(n15945), .A3(n15944), .ZN(n15948) );
  MUX2_X1 U18900 ( .A(n15951), .B(n15950), .S(n15953), .Z(n15955) );
  NAND2_X1 U18901 ( .A1(n15952), .A2(n24981), .ZN(n15954) );
  AOI22_X1 U18902 ( .A1(n15956), .A2(n372), .B1(n17049), .B2(n16628), .ZN(
        n15957) );
  NOR2_X1 U18903 ( .A1(n1329), .A2(n16427), .ZN(n15959) );
  MUX2_X1 U18904 ( .A(n15960), .B(n15959), .S(n15958), .Z(n15964) );
  NOR2_X1 U18905 ( .A1(n15962), .A2(n16422), .ZN(n15963) );
  OAI21_X1 U18906 ( .B1(n16156), .B2(n16122), .A(n15965), .ZN(n15966) );
  NAND2_X1 U18907 ( .A1(n15966), .A2(n16155), .ZN(n15969) );
  OAI21_X1 U18908 ( .B1(n24459), .B2(n2996), .A(n16125), .ZN(n15967) );
  NAND2_X1 U18909 ( .A1(n15967), .A2(n16156), .ZN(n15968) );
  AOI21_X1 U18911 ( .B1(n15971), .B2(n16399), .A(n3630), .ZN(n15975) );
  NAND2_X1 U18912 ( .A1(n15973), .A2(n15972), .ZN(n15974) );
  INV_X1 U18913 ( .A(n16391), .ZN(n15978) );
  NAND2_X1 U18914 ( .A1(n15978), .A2(n15977), .ZN(n15983) );
  NAND2_X1 U18915 ( .A1(n16391), .A2(n15849), .ZN(n15979) );
  NAND2_X1 U18916 ( .A1(n15980), .A2(n15979), .ZN(n15981) );
  NAND3_X1 U18917 ( .A1(n16394), .A2(n16162), .A3(n16389), .ZN(n15982) );
  INV_X1 U18918 ( .A(n17042), .ZN(n16998) );
  NAND2_X1 U18919 ( .A1(n16418), .A2(n15984), .ZN(n15989) );
  NAND2_X1 U18920 ( .A1(n16408), .A2(n16412), .ZN(n15985) );
  OAI211_X1 U18921 ( .C1(n16412), .C2(n16409), .A(n16413), .B(n15985), .ZN(
        n15988) );
  NOR2_X1 U18922 ( .A1(n16141), .A2(n16408), .ZN(n15987) );
  INV_X1 U18924 ( .A(n15992), .ZN(n15993) );
  AND2_X1 U18925 ( .A1(n15990), .A2(n25210), .ZN(n15991) );
  NAND2_X1 U18926 ( .A1(n15994), .A2(n16997), .ZN(n15997) );
  OAI21_X1 U18927 ( .B1(n16998), .B2(n374), .A(n15995), .ZN(n15996) );
  XNOR2_X1 U18928 ( .A(n18557), .B(n18312), .ZN(n15999) );
  XNOR2_X1 U18929 ( .A(n15999), .B(n16000), .ZN(n16093) );
  NAND2_X1 U18930 ( .A1(n16001), .A2(n16268), .ZN(n16007) );
  NOR2_X1 U18931 ( .A1(n16002), .A2(n25009), .ZN(n16003) );
  NAND2_X1 U18932 ( .A1(n16266), .A2(n16003), .ZN(n16006) );
  MUX2_X1 U18933 ( .A(n3554), .B(n16309), .S(n15556), .Z(n16013) );
  OAI22_X1 U18934 ( .A1(n16638), .A2(n16010), .B1(n16309), .B2(n16009), .ZN(
        n16011) );
  INV_X1 U18935 ( .A(n25406), .ZN(n16844) );
  OAI21_X1 U18936 ( .B1(n16342), .B2(n16285), .A(n16286), .ZN(n16014) );
  NAND2_X1 U18937 ( .A1(n16247), .A2(n16016), .ZN(n16017) );
  OAI21_X1 U18938 ( .B1(n16253), .B2(n25284), .A(n16017), .ZN(n16019) );
  NAND2_X1 U18939 ( .A1(n16019), .A2(n15762), .ZN(n16020) );
  OAI22_X1 U18940 ( .A1(n16226), .A2(n16023), .B1(n16225), .B2(n16022), .ZN(
        n16228) );
  INV_X1 U18941 ( .A(n16024), .ZN(n16026) );
  NAND2_X1 U18942 ( .A1(n16277), .A2(n16029), .ZN(n16031) );
  INV_X1 U18943 ( .A(n16032), .ZN(n16033) );
  NOR2_X1 U18944 ( .A1(n17067), .A2(n369), .ZN(n16035) );
  OAI21_X1 U18945 ( .B1(n16546), .B2(n17069), .A(n17067), .ZN(n16036) );
  INV_X1 U18946 ( .A(n16546), .ZN(n16612) );
  INV_X1 U18947 ( .A(n16041), .ZN(n16046) );
  NAND2_X1 U18948 ( .A1(n16043), .A2(n16042), .ZN(n16045) );
  INV_X1 U18949 ( .A(n16260), .ZN(n16533) );
  MUX2_X1 U18950 ( .A(n16048), .B(n294), .S(n24352), .Z(n16049) );
  NAND2_X1 U18951 ( .A1(n16049), .A2(n16509), .ZN(n16055) );
  NOR2_X1 U18952 ( .A1(n16050), .A2(n16508), .ZN(n16052) );
  OAI21_X1 U18954 ( .B1(n24551), .B2(n16469), .A(n16057), .ZN(n16058) );
  INV_X1 U18956 ( .A(n16060), .ZN(n16061) );
  NOR2_X1 U18957 ( .A1(n16062), .A2(n16061), .ZN(n16066) );
  MUX2_X1 U18958 ( .A(n16066), .B(n16065), .S(n16064), .Z(n16071) );
  NAND2_X1 U18960 ( .A1(n16129), .A2(n16076), .ZN(n16072) );
  NOR2_X1 U18963 ( .A1(n16077), .A2(n16076), .ZN(n16078) );
  OAI21_X1 U18964 ( .B1(n1365), .B2(n16075), .A(n16078), .ZN(n17157) );
  INV_X1 U18965 ( .A(n17164), .ZN(n16262) );
  INV_X1 U18967 ( .A(n16082), .ZN(n16083) );
  NAND2_X1 U18968 ( .A1(n16083), .A2(n16100), .ZN(n16087) );
  NAND3_X1 U18969 ( .A1(n16085), .A2(n16101), .A3(n16084), .ZN(n16086) );
  OAI21_X1 U18970 ( .B1(n16375), .B2(n25219), .A(n17166), .ZN(n16089) );
  XNOR2_X1 U18971 ( .A(n18375), .B(n23883), .ZN(n16090) );
  XNOR2_X1 U18972 ( .A(n16091), .B(n16090), .ZN(n16092) );
  NOR2_X1 U18973 ( .A1(n15625), .A2(n16096), .ZN(n16094) );
  OAI21_X1 U18974 ( .B1(n16151), .B2(n16095), .A(n16094), .ZN(n16098) );
  NOR2_X1 U18975 ( .A1(n16114), .A2(n16113), .ZN(n16115) );
  NAND2_X1 U18976 ( .A1(n16123), .A2(n25449), .ZN(n16128) );
  INV_X1 U18977 ( .A(n24459), .ZN(n16124) );
  NOR2_X1 U18978 ( .A1(n16155), .A2(n2996), .ZN(n16126) );
  AOI21_X1 U18979 ( .B1(n16130), .B2(n16129), .A(n24826), .ZN(n16132) );
  MUX2_X1 U18980 ( .A(n16134), .B(n16432), .S(n17174), .Z(n16135) );
  INV_X1 U18981 ( .A(n16780), .ZN(n17348) );
  INV_X1 U18982 ( .A(n17342), .ZN(n17242) );
  OAI21_X1 U18984 ( .B1(n16778), .B2(n17346), .A(n16136), .ZN(n16137) );
  NOR2_X1 U18985 ( .A1(n16777), .A2(n16137), .ZN(n16138) );
  XNOR2_X1 U18987 ( .A(n25077), .B(n18277), .ZN(n16215) );
  NOR2_X1 U18989 ( .A1(n16418), .A2(n16141), .ZN(n16411) );
  NOR2_X1 U18990 ( .A1(n16413), .A2(n16417), .ZN(n16142) );
  NOR2_X1 U18991 ( .A1(n16411), .A2(n16142), .ZN(n16143) );
  OAI21_X1 U18992 ( .B1(n16148), .B2(n4418), .A(n16147), .ZN(n16150) );
  AOI22_X1 U18993 ( .A1(n16152), .A2(n16151), .B1(n16150), .B2(n213), .ZN(
        n16660) );
  NOR2_X1 U18994 ( .A1(n17399), .A2(n17031), .ZN(n17397) );
  INV_X1 U18995 ( .A(n17397), .ZN(n16182) );
  NAND2_X1 U18998 ( .A1(n381), .A2(n2996), .ZN(n16157) );
  MUX2_X1 U18999 ( .A(n16158), .B(n16157), .S(n16156), .Z(n16159) );
  INV_X1 U19001 ( .A(n17395), .ZN(n17196) );
  MUX2_X1 U19002 ( .A(n16163), .B(n16162), .S(n16392), .Z(n16168) );
  INV_X1 U19003 ( .A(n16161), .ZN(n16165) );
  AND3_X1 U19004 ( .A1(n16163), .A2(n16391), .A3(n16162), .ZN(n16164) );
  AOI21_X1 U19005 ( .B1(n16165), .B2(n16167), .A(n16164), .ZN(n16166) );
  NAND2_X1 U19006 ( .A1(n16169), .A2(n244), .ZN(n16173) );
  NAND2_X1 U19007 ( .A1(n16383), .A2(n16381), .ZN(n16179) );
  NOR3_X1 U19008 ( .A1(n4046), .A2(n16177), .A3(n16381), .ZN(n16178) );
  NOR2_X1 U19009 ( .A1(n17400), .A2(n17192), .ZN(n17396) );
  NAND2_X1 U19010 ( .A1(n17396), .A2(n17031), .ZN(n16181) );
  NAND2_X1 U19011 ( .A1(n16339), .A2(n16183), .ZN(n16184) );
  NAND2_X1 U19012 ( .A1(n16187), .A2(n16186), .ZN(n16189) );
  NAND2_X1 U19013 ( .A1(n16189), .A2(n16188), .ZN(n16190) );
  INV_X1 U19014 ( .A(n17185), .ZN(n16203) );
  NOR2_X1 U19015 ( .A1(n16192), .A2(n16191), .ZN(n16327) );
  NOR2_X1 U19016 ( .A1(n16324), .A2(n16193), .ZN(n16195) );
  NAND2_X1 U19017 ( .A1(n16203), .A2(n17391), .ZN(n16214) );
  NAND3_X1 U19018 ( .A1(n3544), .A2(n16401), .A3(n25500), .ZN(n16201) );
  MUX2_X1 U19019 ( .A(n16205), .B(n17182), .S(n16204), .Z(n16210) );
  INV_X1 U19020 ( .A(n16366), .ZN(n16209) );
  NOR2_X1 U19021 ( .A1(n17180), .A2(n16206), .ZN(n16208) );
  INV_X1 U19022 ( .A(n17387), .ZN(n17186) );
  NAND2_X1 U19024 ( .A1(n16349), .A2(n16597), .ZN(n16211) );
  NAND2_X1 U19025 ( .A1(n17389), .A2(n17185), .ZN(n16212) );
  XNOR2_X1 U19026 ( .A(n17863), .B(n18549), .ZN(n18342) );
  XNOR2_X1 U19027 ( .A(n18342), .B(n16215), .ZN(n16322) );
  INV_X1 U19028 ( .A(n16216), .ZN(n16218) );
  MUX2_X1 U19029 ( .A(n16218), .B(n16217), .S(n16462), .Z(n16223) );
  NOR2_X2 U19030 ( .A1(n16223), .A2(n16222), .ZN(n17212) );
  OAI21_X1 U19031 ( .B1(n16302), .B2(n16225), .A(n16224), .ZN(n16227) );
  NOR2_X1 U19032 ( .A1(n16231), .A2(n16230), .ZN(n16233) );
  OAI211_X1 U19033 ( .C1(n16235), .C2(n385), .A(n16450), .B(n16447), .ZN(
        n16238) );
  INV_X1 U19034 ( .A(n16447), .ZN(n16236) );
  INV_X1 U19035 ( .A(n17017), .ZN(n16240) );
  OAI22_X1 U19036 ( .A1(n2636), .A2(n16442), .B1(n16443), .B2(n16242), .ZN(
        n16244) );
  NAND2_X1 U19037 ( .A1(n16244), .A2(n16243), .ZN(n16245) );
  NOR2_X1 U19038 ( .A1(n16246), .A2(n15762), .ZN(n16250) );
  XNOR2_X1 U19043 ( .A(n24384), .B(n3164), .ZN(n16320) );
  NAND2_X1 U19044 ( .A1(n16375), .A2(n25219), .ZN(n16532) );
  INV_X1 U19046 ( .A(n25219), .ZN(n17160) );
  INV_X1 U19047 ( .A(n17824), .ZN(n18006) );
  AOI21_X1 U19048 ( .B1(n25009), .B2(n16268), .A(n16266), .ZN(n16271) );
  NAND3_X1 U19050 ( .A1(n16277), .A2(n16276), .A3(n24403), .ZN(n16278) );
  INV_X1 U19051 ( .A(n16345), .ZN(n16281) );
  NOR2_X1 U19052 ( .A1(n16281), .A2(n24540), .ZN(n16283) );
  OAI21_X1 U19053 ( .B1(n16286), .B2(n16285), .A(n24540), .ZN(n16287) );
  NOR2_X1 U19054 ( .A1(n16347), .A2(n16287), .ZN(n16288) );
  INV_X1 U19057 ( .A(n16363), .ZN(n16295) );
  NOR2_X1 U19058 ( .A1(n16293), .A2(n25546), .ZN(n16294) );
  OAI21_X1 U19059 ( .B1(n16295), .B2(n16294), .A(n16357), .ZN(n16296) );
  INV_X1 U19061 ( .A(n16298), .ZN(n16300) );
  NAND2_X1 U19062 ( .A1(n16302), .A2(n16301), .ZN(n16306) );
  MUX2_X1 U19063 ( .A(n16306), .B(n16305), .S(n16304), .Z(n16307) );
  AOI21_X1 U19064 ( .B1(n16311), .B2(n15557), .A(n3554), .ZN(n16310) );
  XNOR2_X1 U19065 ( .A(n18646), .B(n18006), .ZN(n16319) );
  XNOR2_X1 U19066 ( .A(n16320), .B(n16319), .ZN(n16321) );
  XNOR2_X1 U19067 ( .A(n16321), .B(n16322), .ZN(n19132) );
  NOR2_X1 U19068 ( .A1(n25323), .A2(n16324), .ZN(n16326) );
  NOR2_X1 U19069 ( .A1(n16327), .A2(n16326), .ZN(n16329) );
  OAI21_X1 U19070 ( .B1(n3947), .B2(n16332), .A(n25455), .ZN(n16340) );
  NOR2_X2 U19075 ( .A1(n16348), .A2(n16347), .ZN(n17455) );
  INV_X1 U19076 ( .A(n17455), .ZN(n16354) );
  NAND2_X1 U19077 ( .A1(n24890), .A2(n24467), .ZN(n16353) );
  OAI21_X1 U19078 ( .B1(n15822), .B2(n16349), .A(n16595), .ZN(n16351) );
  OAI21_X1 U19079 ( .B1(n16357), .B2(n24456), .A(n16355), .ZN(n16362) );
  MUX2_X1 U19081 ( .A(n16362), .B(n16361), .S(n16360), .Z(n16364) );
  AND2_X1 U19086 ( .A1(n17297), .A2(n17296), .ZN(n16371) );
  NAND2_X1 U19087 ( .A1(n17299), .A2(n17297), .ZN(n16372) );
  XNOR2_X1 U19090 ( .A(n18532), .B(n18610), .ZN(n16380) );
  INV_X1 U19091 ( .A(n16375), .ZN(n16838) );
  NAND3_X1 U19092 ( .A1(n17163), .A2(n17160), .A3(n16838), .ZN(n16377) );
  NAND2_X1 U19093 ( .A1(n16533), .A2(n17166), .ZN(n16376) );
  OAI211_X2 U19094 ( .C1(n16378), .C2(n17164), .A(n16377), .B(n16376), .ZN(
        n18270) );
  XNOR2_X1 U19095 ( .A(n18270), .B(n1951), .ZN(n16379) );
  XNOR2_X1 U19096 ( .A(n16380), .B(n16379), .ZN(n16503) );
  NOR2_X1 U19097 ( .A1(n16383), .A2(n16382), .ZN(n16384) );
  NOR2_X1 U19098 ( .A1(n16385), .A2(n16384), .ZN(n16386) );
  OAI21_X1 U19099 ( .B1(n16390), .B2(n5758), .A(n16389), .ZN(n16396) );
  AOI21_X1 U19100 ( .B1(n16393), .B2(n16392), .A(n16391), .ZN(n16395) );
  INV_X1 U19101 ( .A(n16400), .ZN(n17433) );
  INV_X1 U19102 ( .A(n17439), .ZN(n16828) );
  AOI21_X1 U19103 ( .B1(n16402), .B2(n16401), .A(n16404), .ZN(n16407) );
  NOR2_X1 U19104 ( .A1(n16409), .A2(n16408), .ZN(n16410) );
  NOR2_X1 U19105 ( .A1(n16413), .A2(n16412), .ZN(n16415) );
  NAND2_X1 U19106 ( .A1(n16417), .A2(n16416), .ZN(n16419) );
  NOR2_X1 U19107 ( .A1(n16419), .A2(n16418), .ZN(n16420) );
  INV_X1 U19110 ( .A(n17442), .ZN(n16964) );
  INV_X1 U19111 ( .A(n16432), .ZN(n16433) );
  AOI21_X1 U19112 ( .B1(n17171), .B2(n17522), .A(n16433), .ZN(n16436) );
  XNOR2_X1 U19113 ( .A(n24565), .B(n18335), .ZN(n18101) );
  AOI21_X1 U19114 ( .B1(n16438), .B2(n16437), .A(n16442), .ZN(n16439) );
  NAND2_X1 U19115 ( .A1(n16441), .A2(n16440), .ZN(n16445) );
  MUX2_X1 U19116 ( .A(n385), .B(n16448), .S(n16447), .Z(n16457) );
  NAND2_X1 U19117 ( .A1(n16450), .A2(n16449), .ZN(n16455) );
  NAND2_X1 U19118 ( .A1(n385), .A2(n257), .ZN(n16453) );
  OAI22_X1 U19119 ( .A1(n16455), .A2(n223), .B1(n16453), .B2(n16452), .ZN(
        n16456) );
  INV_X1 U19120 ( .A(n16849), .ZN(n17139) );
  AND2_X1 U19121 ( .A1(n17144), .A2(n17139), .ZN(n16488) );
  NOR2_X1 U19123 ( .A1(n5269), .A2(n16464), .ZN(n16467) );
  OAI21_X1 U19124 ( .B1(n16467), .B2(n16466), .A(n16465), .ZN(n16468) );
  INV_X1 U19125 ( .A(n16984), .ZN(n17140) );
  MUX2_X1 U19126 ( .A(n16471), .B(n24550), .S(n16469), .Z(n16479) );
  OAI21_X1 U19127 ( .B1(n16474), .B2(n16473), .A(n16472), .ZN(n16478) );
  NOR2_X1 U19128 ( .A1(n16476), .A2(n16475), .ZN(n16477) );
  INV_X1 U19129 ( .A(n16851), .ZN(n17137) );
  NOR2_X1 U19130 ( .A1(n17140), .A2(n17137), .ZN(n16487) );
  NAND2_X1 U19131 ( .A1(n16485), .A2(n16484), .ZN(n16515) );
  NAND2_X1 U19132 ( .A1(n16486), .A2(n16515), .ZN(n17141) );
  NAND2_X1 U19134 ( .A1(n16490), .A2(n16489), .ZN(n16495) );
  NAND2_X1 U19135 ( .A1(n17138), .A2(n16984), .ZN(n16691) );
  NAND3_X1 U19136 ( .A1(n16991), .A2(n287), .A3(n16499), .ZN(n16501) );
  OAI21_X1 U19137 ( .B1(n16021), .B2(n17461), .A(n16991), .ZN(n16500) );
  XNOR2_X1 U19138 ( .A(n17581), .B(n18331), .ZN(n17722) );
  XNOR2_X1 U19139 ( .A(n18101), .B(n17722), .ZN(n16502) );
  MUX2_X2 U19140 ( .A(n16505), .B(n16504), .S(n24324), .Z(n20670) );
  OAI21_X1 U19141 ( .B1(n17467), .B2(n25572), .A(n16506), .ZN(n16507) );
  INV_X1 U19142 ( .A(n17041), .ZN(n18700) );
  NAND2_X1 U19143 ( .A1(n16511), .A2(n16510), .ZN(n16512) );
  MUX2_X1 U19144 ( .A(n16512), .B(n17297), .S(n17299), .Z(n16514) );
  XNOR2_X1 U19145 ( .A(n18700), .B(n18214), .ZN(n16521) );
  NAND2_X1 U19146 ( .A1(n16515), .A2(n17138), .ZN(n16517) );
  OAI21_X1 U19147 ( .B1(n16518), .B2(n16517), .A(n16848), .ZN(n16519) );
  XNOR2_X1 U19148 ( .A(n18605), .B(n1797), .ZN(n16520) );
  XNOR2_X1 U19149 ( .A(n16521), .B(n16520), .ZN(n16538) );
  AOI22_X1 U19150 ( .A1(n16523), .A2(n17522), .B1(n16522), .B2(n17175), .ZN(
        n16525) );
  NOR2_X1 U19151 ( .A1(n17522), .A2(n17171), .ZN(n16524) );
  MUX2_X1 U19152 ( .A(n16525), .B(n16863), .S(n16524), .Z(n17900) );
  NOR2_X1 U19153 ( .A1(n16526), .A2(n16980), .ZN(n16530) );
  INV_X1 U19154 ( .A(n16527), .ZN(n17451) );
  NOR2_X1 U19155 ( .A1(n17455), .A2(n17450), .ZN(n16528) );
  INV_X1 U19156 ( .A(n16532), .ZN(n16534) );
  MUX2_X1 U19157 ( .A(n17166), .B(n17163), .S(n25218), .Z(n16535) );
  XNOR2_X1 U19158 ( .A(n18420), .B(n18451), .ZN(n17974) );
  XNOR2_X1 U19159 ( .A(n17974), .B(n18348), .ZN(n16537) );
  XNOR2_X1 U19160 ( .A(n16537), .B(n16538), .ZN(n18749) );
  AOI21_X1 U19161 ( .B1(n17474), .B2(n17473), .A(n17472), .ZN(n16542) );
  OAI22_X1 U19162 ( .A1(n16540), .A2(n17633), .B1(n16901), .B2(n16902), .ZN(
        n16541) );
  NAND2_X1 U19163 ( .A1(n17288), .A2(n17229), .ZN(n17539) );
  NAND2_X1 U19164 ( .A1(n17540), .A2(n17539), .ZN(n16755) );
  NAND2_X1 U19165 ( .A1(n17288), .A2(n17283), .ZN(n16543) );
  AOI21_X1 U19166 ( .B1(n16543), .B2(n17229), .A(n17293), .ZN(n16544) );
  XNOR2_X1 U19167 ( .A(n18659), .B(n17993), .ZN(n18359) );
  INV_X1 U19168 ( .A(n18359), .ZN(n18529) );
  INV_X1 U19169 ( .A(n17919), .ZN(n16555) );
  AOI21_X1 U19170 ( .B1(n16796), .B2(n16794), .A(n5375), .ZN(n16554) );
  NOR2_X1 U19171 ( .A1(n16550), .A2(n16547), .ZN(n16548) );
  NAND2_X1 U19172 ( .A1(n16549), .A2(n16548), .ZN(n16553) );
  XNOR2_X1 U19173 ( .A(n17680), .B(n16555), .ZN(n16937) );
  XNOR2_X1 U19174 ( .A(n18529), .B(n16937), .ZN(n16571) );
  OAI21_X1 U19176 ( .B1(n17216), .B2(n17207), .A(n17015), .ZN(n16558) );
  NAND2_X1 U19177 ( .A1(n16558), .A2(n17212), .ZN(n16559) );
  INV_X1 U19178 ( .A(n18102), .ZN(n17649) );
  XNOR2_X1 U19179 ( .A(n17649), .B(n2145), .ZN(n16569) );
  NAND2_X1 U19180 ( .A1(n16942), .A2(n16940), .ZN(n16564) );
  INV_X1 U19181 ( .A(n16743), .ZN(n16560) );
  AOI21_X1 U19182 ( .B1(n17224), .B2(n17413), .A(n16956), .ZN(n16568) );
  INV_X1 U19183 ( .A(n17419), .ZN(n16565) );
  NAND3_X1 U19185 ( .A1(n16565), .A2(n17227), .A3(n25246), .ZN(n16566) );
  XNOR2_X1 U19187 ( .A(n18269), .B(n18530), .ZN(n18405) );
  XNOR2_X1 U19188 ( .A(n18405), .B(n16569), .ZN(n16570) );
  NAND2_X1 U19190 ( .A1(n18749), .A2(n24421), .ZN(n19562) );
  NOR2_X1 U19192 ( .A1(n16572), .A2(n17120), .ZN(n16573) );
  MUX2_X1 U19193 ( .A(n17134), .B(n25245), .S(n17132), .Z(n16577) );
  OAI21_X1 U19194 ( .B1(n16649), .B2(n17086), .A(n16740), .ZN(n16581) );
  NAND2_X1 U19195 ( .A1(n17086), .A2(n16578), .ZN(n16579) );
  INV_X1 U19196 ( .A(n17086), .ZN(n16648) );
  OAI22_X1 U19197 ( .A1(n17084), .A2(n16579), .B1(n16648), .B2(n371), .ZN(
        n16580) );
  XNOR2_X1 U19198 ( .A(n17970), .B(n17881), .ZN(n18246) );
  XNOR2_X1 U19199 ( .A(n18246), .B(n16582), .ZN(n16601) );
  AOI21_X1 U19200 ( .B1(n16901), .B2(n17472), .A(n17629), .ZN(n16587) );
  NAND2_X1 U19201 ( .A1(n17633), .A2(n16539), .ZN(n16583) );
  OAI21_X1 U19202 ( .B1(n2561), .B2(n17633), .A(n16583), .ZN(n16586) );
  INV_X1 U19203 ( .A(n17472), .ZN(n16584) );
  NAND2_X1 U19204 ( .A1(n16584), .A2(n17633), .ZN(n16585) );
  INV_X1 U19206 ( .A(n17478), .ZN(n17079) );
  NAND2_X1 U19207 ( .A1(n17479), .A2(n17079), .ZN(n16589) );
  AOI21_X1 U19208 ( .B1(n16590), .B2(n16589), .A(n16588), .ZN(n16593) );
  NAND2_X1 U19209 ( .A1(n17481), .A2(n17078), .ZN(n16591) );
  XNOR2_X1 U19211 ( .A(n18685), .B(n18042), .ZN(n16599) );
  INV_X1 U19212 ( .A(n16888), .ZN(n17730) );
  INV_X1 U19213 ( .A(n17734), .ZN(n17731) );
  XNOR2_X1 U19214 ( .A(n16599), .B(n18370), .ZN(n18520) );
  INV_X1 U19215 ( .A(n17334), .ZN(n16973) );
  INV_X1 U19216 ( .A(n16726), .ZN(n16606) );
  INV_X1 U19217 ( .A(n17333), .ZN(n16604) );
  NOR2_X1 U19218 ( .A1(n17335), .A2(n16602), .ZN(n16603) );
  AOI22_X1 U19220 ( .A1(n17599), .A2(n17316), .B1(n17304), .B2(n16921), .ZN(
        n16920) );
  INV_X1 U19221 ( .A(n17316), .ZN(n16715) );
  NOR2_X1 U19222 ( .A1(n17304), .A2(n24542), .ZN(n16714) );
  OAI21_X1 U19223 ( .B1(n3783), .B2(n17316), .A(n16714), .ZN(n16608) );
  OAI21_X1 U19224 ( .B1(n16920), .B2(n16716), .A(n16608), .ZN(n17757) );
  XNOR2_X1 U19225 ( .A(n18220), .B(n18431), .ZN(n16625) );
  INV_X1 U19226 ( .A(n16619), .ZN(n16621) );
  NAND2_X1 U19227 ( .A1(n16622), .A2(n16795), .ZN(n16798) );
  NAND2_X1 U19228 ( .A1(n5762), .A2(n16798), .ZN(n16623) );
  XNOR2_X1 U19229 ( .A(n17476), .B(n1870), .ZN(n16624) );
  XNOR2_X1 U19230 ( .A(n16625), .B(n16624), .ZN(n16626) );
  NAND2_X1 U19231 ( .A1(n19560), .A2(n19559), .ZN(n16666) );
  NOR2_X1 U19232 ( .A1(n17216), .A2(n25201), .ZN(n16878) );
  NOR2_X1 U19233 ( .A1(n17185), .A2(n17179), .ZN(n16627) );
  XNOR2_X1 U19234 ( .A(n17515), .B(n18541), .ZN(n18439) );
  MUX2_X1 U19235 ( .A(n17050), .B(n16628), .S(n17049), .Z(n16634) );
  NAND3_X1 U19236 ( .A1(n16775), .A2(n24570), .A3(n17053), .ZN(n16632) );
  INV_X1 U19237 ( .A(n17049), .ZN(n16629) );
  XNOR2_X1 U19238 ( .A(n18439), .B(n16635), .ZN(n16665) );
  INV_X1 U19239 ( .A(n17381), .ZN(n17422) );
  NOR2_X1 U19240 ( .A1(n17379), .A2(n17422), .ZN(n16637) );
  INV_X1 U19241 ( .A(n17425), .ZN(n17382) );
  NOR2_X1 U19242 ( .A1(n17382), .A2(n5409), .ZN(n16636) );
  MUX2_X1 U19243 ( .A(n16637), .B(n16636), .S(n24330), .Z(n16646) );
  NAND2_X1 U19244 ( .A1(n16639), .A2(n16638), .ZN(n16640) );
  NAND2_X1 U19245 ( .A1(n16641), .A2(n16640), .ZN(n17423) );
  INV_X1 U19246 ( .A(n17423), .ZN(n16642) );
  NAND2_X1 U19247 ( .A1(n17382), .A2(n16642), .ZN(n16643) );
  AOI21_X1 U19248 ( .B1(n16644), .B2(n16643), .A(n5406), .ZN(n16645) );
  NOR2_X2 U19249 ( .A1(n16646), .A2(n16645), .ZN(n18666) );
  INV_X1 U19250 ( .A(n16647), .ZN(n16652) );
  NAND2_X1 U19251 ( .A1(n16650), .A2(n16739), .ZN(n16651) );
  NAND2_X1 U19252 ( .A1(n17132), .A2(n16655), .ZN(n16658) );
  NOR2_X1 U19253 ( .A1(n25227), .A2(n3458), .ZN(n16654) );
  NAND2_X1 U19254 ( .A1(n17134), .A2(n16654), .ZN(n16657) );
  OAI211_X1 U19255 ( .C1(n17134), .C2(n16658), .A(n16657), .B(n16656), .ZN(
        n16910) );
  INV_X1 U19256 ( .A(n16910), .ZN(n16663) );
  NAND2_X1 U19257 ( .A1(n17399), .A2(n17395), .ZN(n16659) );
  NAND2_X1 U19258 ( .A1(n16659), .A2(n17031), .ZN(n17030) );
  NAND2_X1 U19260 ( .A1(n17400), .A2(n17028), .ZN(n16661) );
  XNOR2_X1 U19261 ( .A(n16663), .B(n17840), .ZN(n18381) );
  AOI21_X1 U19262 ( .B1(n19562), .B2(n16666), .A(n19555), .ZN(n16701) );
  NAND2_X1 U19263 ( .A1(n17347), .A2(n17346), .ZN(n16668) );
  NAND3_X1 U19264 ( .A1(n17241), .A2(n17343), .A3(n17236), .ZN(n16667) );
  OAI21_X1 U19265 ( .B1(n16668), .B2(n17348), .A(n16667), .ZN(n17206) );
  NOR2_X2 U19266 ( .A1(n16669), .A2(n17206), .ZN(n18227) );
  OAI21_X1 U19267 ( .B1(n17051), .B2(n17050), .A(n17053), .ZN(n16670) );
  MUX2_X1 U19268 ( .A(n25214), .B(n25058), .S(n17039), .Z(n16988) );
  NOR3_X1 U19269 ( .A1(n16770), .A2(n25058), .A3(n25214), .ZN(n16671) );
  NAND2_X1 U19270 ( .A1(n266), .A2(n17351), .ZN(n16672) );
  NAND2_X1 U19271 ( .A1(n16672), .A2(n17356), .ZN(n16675) );
  NOR2_X1 U19272 ( .A1(n17014), .A2(n17351), .ZN(n16876) );
  OR2_X1 U19273 ( .A1(n16672), .A2(n4004), .ZN(n16674) );
  XNOR2_X1 U19274 ( .A(n18674), .B(n17663), .ZN(n18501) );
  XNOR2_X1 U19275 ( .A(n17679), .B(n18501), .ZN(n16698) );
  NAND2_X1 U19276 ( .A1(n374), .A2(n17368), .ZN(n16676) );
  AND2_X1 U19278 ( .A1(n17573), .A2(n17574), .ZN(n16677) );
  NAND3_X1 U19279 ( .A1(n16682), .A2(n16681), .A3(n16680), .ZN(n16685) );
  INV_X1 U19280 ( .A(n16683), .ZN(n16684) );
  OAI22_X1 U19281 ( .A1(n16685), .A2(n16684), .B1(n17277), .B2(n17273), .ZN(
        n16690) );
  NAND4_X1 U19282 ( .A1(n16687), .A2(n17273), .A3(n16686), .A4(n17276), .ZN(
        n16689) );
  NAND3_X1 U19283 ( .A1(n17279), .A2(n17254), .A3(n17249), .ZN(n16688) );
  AND3_X1 U19285 ( .A1(n17145), .A2(n16985), .A3(n17137), .ZN(n16693) );
  INV_X1 U19286 ( .A(n17664), .ZN(n18116) );
  XNOR2_X1 U19287 ( .A(n18116), .B(n21533), .ZN(n16696) );
  XNOR2_X1 U19288 ( .A(n18390), .B(n16696), .ZN(n16697) );
  NAND2_X1 U19289 ( .A1(n19290), .A2(n19559), .ZN(n16699) );
  AOI21_X1 U19290 ( .B1(n16699), .B2(n19560), .A(n19138), .ZN(n16700) );
  INV_X1 U19291 ( .A(n18678), .ZN(n16713) );
  OAI21_X1 U19292 ( .B1(n17319), .B2(n17320), .A(n17321), .ZN(n16712) );
  XNOR2_X1 U19293 ( .A(n16713), .B(n18633), .ZN(n18303) );
  INV_X1 U19294 ( .A(n18303), .ZN(n17912) );
  XNOR2_X1 U19295 ( .A(n17912), .B(n18226), .ZN(n16738) );
  XNOR2_X1 U19296 ( .A(n18188), .B(n2228), .ZN(n16736) );
  NAND3_X1 U19297 ( .A1(n17332), .A2(n17336), .A3(n17335), .ZN(n16729) );
  NAND2_X1 U19298 ( .A1(n25412), .A2(n17335), .ZN(n16725) );
  XNOR2_X1 U19299 ( .A(n17788), .B(n16736), .ZN(n16737) );
  XNOR2_X1 U19301 ( .A(n18195), .B(n1875), .ZN(n16745) );
  NOR2_X1 U19302 ( .A1(n17086), .A2(n17085), .ZN(n16741) );
  NOR2_X1 U19303 ( .A1(n17615), .A2(n17408), .ZN(n16744) );
  XNOR2_X1 U19304 ( .A(n18432), .B(n18693), .ZN(n17785) );
  XNOR2_X1 U19305 ( .A(n17785), .B(n16745), .ZN(n16761) );
  INV_X1 U19308 ( .A(n17421), .ZN(n16752) );
  NOR2_X1 U19309 ( .A1(n17423), .A2(n17424), .ZN(n16749) );
  OAI21_X1 U19310 ( .B1(n17381), .B2(n17421), .A(n16749), .ZN(n16751) );
  NAND3_X1 U19311 ( .A1(n17425), .A2(n16752), .A3(n17423), .ZN(n16750) );
  OAI211_X1 U19312 ( .C1(n17379), .C2(n16752), .A(n16751), .B(n16750), .ZN(
        n18476) );
  NAND2_X1 U19314 ( .A1(n17289), .A2(n17284), .ZN(n17538) );
  NAND2_X1 U19315 ( .A1(n17541), .A2(n17538), .ZN(n16754) );
  OAI21_X1 U19317 ( .B1(n16755), .B2(n16754), .A(n17544), .ZN(n16759) );
  NAND2_X1 U19318 ( .A1(n17419), .A2(n25433), .ZN(n16756) );
  NAND2_X1 U19319 ( .A1(n17227), .A2(n25246), .ZN(n16757) );
  XNOR2_X1 U19320 ( .A(n16759), .B(n17931), .ZN(n18218) );
  XNOR2_X1 U19321 ( .A(n16761), .B(n16760), .ZN(n19261) );
  NAND2_X1 U19322 ( .A1(n24386), .A2(n19261), .ZN(n19146) );
  INV_X1 U19323 ( .A(n17368), .ZN(n17571) );
  INV_X1 U19324 ( .A(n18233), .ZN(n16768) );
  XNOR2_X1 U19325 ( .A(n16768), .B(n17681), .ZN(n18142) );
  INV_X1 U19326 ( .A(n16770), .ZN(n17040) );
  AOI22_X1 U19328 ( .A1(n17364), .A2(n25058), .B1(n16989), .B2(n16770), .ZN(
        n16771) );
  NAND3_X1 U19331 ( .A1(n16775), .A2(n17049), .A3(n17050), .ZN(n16776) );
  XNOR2_X1 U19332 ( .A(n18660), .B(n18611), .ZN(n18333) );
  XNOR2_X1 U19333 ( .A(n18142), .B(n18333), .ZN(n16786) );
  INV_X1 U19334 ( .A(n16778), .ZN(n16779) );
  INV_X1 U19335 ( .A(n17581), .ZN(n16783) );
  XNOR2_X1 U19336 ( .A(n18103), .B(n16783), .ZN(n18178) );
  XNOR2_X1 U19337 ( .A(n16784), .B(n18178), .ZN(n16785) );
  NAND2_X1 U19339 ( .A1(n17134), .A2(n17132), .ZN(n16787) );
  OAI21_X1 U19340 ( .B1(n17134), .B2(n4684), .A(n16787), .ZN(n16790) );
  INV_X1 U19343 ( .A(n18208), .ZN(n16800) );
  XNOR2_X1 U19345 ( .A(n18602), .B(n16799), .ZN(n18324) );
  INV_X1 U19346 ( .A(n18324), .ZN(n17898) );
  XNOR2_X1 U19347 ( .A(n17898), .B(n16800), .ZN(n16821) );
  MUX2_X1 U19348 ( .A(n17100), .B(n25357), .S(n17114), .Z(n16804) );
  NOR2_X1 U19349 ( .A1(n16802), .A2(n16801), .ZN(n16803) );
  MUX2_X2 U19350 ( .A(n16804), .B(n16803), .S(n2581), .Z(n18446) );
  XNOR2_X1 U19351 ( .A(n18446), .B(n20995), .ZN(n16819) );
  NAND2_X1 U19352 ( .A1(n17081), .A2(n16809), .ZN(n16896) );
  AOI21_X1 U19353 ( .B1(n17481), .B2(n17077), .A(n17078), .ZN(n16807) );
  NAND2_X1 U19354 ( .A1(n24660), .A2(n17478), .ZN(n16806) );
  NAND3_X1 U19356 ( .A1(n16810), .A2(n16809), .A3(n16808), .ZN(n17477) );
  NOR2_X1 U19357 ( .A1(n25429), .A2(n17477), .ZN(n16811) );
  NAND2_X1 U19359 ( .A1(n17729), .A2(n25472), .ZN(n16817) );
  NAND2_X1 U19360 ( .A1(n25472), .A2(n17734), .ZN(n16814) );
  NOR2_X1 U19361 ( .A1(n17728), .A2(n17485), .ZN(n17094) );
  INV_X1 U19362 ( .A(n17094), .ZN(n16813) );
  XNOR2_X1 U19364 ( .A(n18418), .B(n18149), .ZN(n18607) );
  INV_X1 U19365 ( .A(n18607), .ZN(n16818) );
  XNOR2_X1 U19366 ( .A(n16819), .B(n16818), .ZN(n16820) );
  XNOR2_X1 U19367 ( .A(n16821), .B(n16820), .ZN(n17556) );
  NAND3_X1 U19368 ( .A1(n19146), .A2(n16822), .A3(n18919), .ZN(n16887) );
  INV_X1 U19369 ( .A(n17171), .ZN(n17523) );
  MUX2_X1 U19370 ( .A(n16862), .B(n16823), .S(n17174), .Z(n16825) );
  OAI21_X1 U19371 ( .B1(n17170), .B2(n17173), .A(n17523), .ZN(n16824) );
  INV_X1 U19372 ( .A(n17445), .ZN(n17125) );
  INV_X1 U19374 ( .A(n16826), .ZN(n16827) );
  AOI22_X1 U19375 ( .A1(n17125), .A2(n2549), .B1(n16827), .B2(n16964), .ZN(
        n16831) );
  OAI22_X1 U19376 ( .A1(n16831), .A2(n16830), .B1(n1612), .B2(n16829), .ZN(
        n17905) );
  XNOR2_X1 U19377 ( .A(n17839), .B(n17905), .ZN(n18237) );
  INV_X1 U19378 ( .A(n16979), .ZN(n17457) );
  AOI21_X1 U19379 ( .B1(n17455), .B2(n523), .A(n17457), .ZN(n16833) );
  OAI21_X1 U19380 ( .B1(n17163), .B2(n17165), .A(n16836), .ZN(n16837) );
  INV_X1 U19381 ( .A(n16837), .ZN(n16842) );
  NAND2_X1 U19382 ( .A1(n17164), .A2(n17166), .ZN(n16840) );
  MUX2_X1 U19384 ( .A(n16840), .B(n16839), .S(n17163), .Z(n16841) );
  XNOR2_X1 U19385 ( .A(n18124), .B(n18121), .ZN(n16843) );
  XNOR2_X1 U19386 ( .A(n18237), .B(n16843), .ZN(n16858) );
  INV_X1 U19387 ( .A(n16847), .ZN(n16854) );
  AND2_X1 U19388 ( .A1(n17144), .A2(n16985), .ZN(n16850) );
  NAND3_X1 U19389 ( .A1(n17138), .A2(n16851), .A3(n17139), .ZN(n16852) );
  XNOR2_X1 U19391 ( .A(n18435), .B(n18669), .ZN(n16856) );
  XNOR2_X1 U19392 ( .A(n18382), .B(n2208), .ZN(n16855) );
  XNOR2_X1 U19393 ( .A(n16855), .B(n16856), .ZN(n16857) );
  XNOR2_X1 U19394 ( .A(n16858), .B(n16857), .ZN(n19266) );
  NAND2_X1 U19395 ( .A1(n19263), .A2(n19266), .ZN(n16886) );
  INV_X1 U19396 ( .A(n17241), .ZN(n17240) );
  XNOR2_X1 U19397 ( .A(n18308), .B(n3152), .ZN(n16868) );
  NOR3_X1 U19398 ( .A1(n17524), .A2(n17170), .A3(n17175), .ZN(n16861) );
  NOR2_X1 U19399 ( .A1(n16862), .A2(n16861), .ZN(n17525) );
  NOR2_X1 U19400 ( .A1(n17524), .A2(n17171), .ZN(n17177) );
  NOR2_X1 U19401 ( .A1(n16863), .A2(n16112), .ZN(n16864) );
  OAI21_X1 U19402 ( .B1(n17177), .B2(n16864), .A(n17522), .ZN(n16865) );
  NAND2_X1 U19403 ( .A1(n17525), .A2(n16865), .ZN(n16866) );
  XNOR2_X1 U19404 ( .A(n16867), .B(n16868), .ZN(n16884) );
  NOR2_X1 U19405 ( .A1(n25003), .A2(n17192), .ZN(n16870) );
  OAI22_X1 U19407 ( .A1(n16873), .A2(n17389), .B1(n16872), .B2(n17387), .ZN(
        n16874) );
  NAND3_X1 U19408 ( .A1(n367), .A2(n4004), .A3(n25491), .ZN(n16877) );
  NAND2_X1 U19409 ( .A1(n16878), .A2(n24391), .ZN(n16882) );
  INV_X1 U19410 ( .A(n17216), .ZN(n17021) );
  NAND2_X1 U19411 ( .A1(n17021), .A2(n17015), .ZN(n16881) );
  NAND3_X1 U19412 ( .A1(n17216), .A2(n17016), .A3(n17208), .ZN(n16879) );
  XNOR2_X1 U19413 ( .A(n18129), .B(n25194), .ZN(n18629) );
  XNOR2_X1 U19414 ( .A(n18248), .B(n18629), .ZN(n16883) );
  XNOR2_X1 U19415 ( .A(n16883), .B(n16884), .ZN(n18914) );
  NAND3_X2 U19416 ( .A1(n16887), .A2(n16886), .A3(n16885), .ZN(n20669) );
  MUX2_X1 U19419 ( .A(n17485), .B(n17728), .S(n17734), .Z(n16889) );
  NOR2_X1 U19420 ( .A1(n17486), .A2(n24410), .ZN(n17737) );
  MUX2_X1 U19421 ( .A(n16889), .B(n17737), .S(n17729), .Z(n16891) );
  NOR3_X1 U19422 ( .A1(n17728), .A2(n17730), .A3(n17731), .ZN(n16890) );
  NOR2_X1 U19423 ( .A1(n16891), .A2(n16890), .ZN(n18122) );
  XNOR2_X1 U19424 ( .A(n18122), .B(n18239), .ZN(n16906) );
  NOR2_X1 U19425 ( .A1(n17077), .A2(n17078), .ZN(n16894) );
  NOR2_X1 U19426 ( .A1(n16896), .A2(n17076), .ZN(n16899) );
  NAND2_X1 U19427 ( .A1(n1033), .A2(n17629), .ZN(n16905) );
  OAI211_X1 U19428 ( .C1(n17472), .C2(n16905), .A(n16904), .B(n16903), .ZN(
        n18038) );
  XNOR2_X1 U19429 ( .A(n18038), .B(n17595), .ZN(n18667) );
  XNOR2_X1 U19430 ( .A(n16906), .B(n18667), .ZN(n16914) );
  MUX2_X1 U19431 ( .A(n17114), .B(n17118), .S(n17119), .Z(n16907) );
  NAND2_X1 U19432 ( .A1(n16907), .A2(n2580), .ZN(n16909) );
  NOR2_X1 U19433 ( .A1(n17120), .A2(n17119), .ZN(n16908) );
  XNOR2_X1 U19434 ( .A(n18582), .B(n836), .ZN(n16912) );
  XNOR2_X1 U19435 ( .A(n17907), .B(n18539), .ZN(n16911) );
  XNOR2_X1 U19436 ( .A(n16912), .B(n16911), .ZN(n16913) );
  XNOR2_X1 U19437 ( .A(n16913), .B(n16914), .ZN(n19309) );
  INV_X1 U19438 ( .A(n16974), .ZN(n16918) );
  OAI21_X1 U19439 ( .B1(n17336), .B2(n16973), .A(n16971), .ZN(n16916) );
  INV_X1 U19441 ( .A(n16920), .ZN(n16922) );
  NAND2_X1 U19442 ( .A1(n17304), .A2(n24543), .ZN(n17314) );
  XNOR2_X1 U19443 ( .A(n17720), .B(n17582), .ZN(n18657) );
  INV_X1 U19444 ( .A(n18657), .ZN(n18176) );
  OAI21_X1 U19446 ( .B1(n17326), .B2(n17319), .A(n4426), .ZN(n16925) );
  AOI22_X2 U19447 ( .A1(n16926), .A2(n16927), .B1(n16925), .B2(n15673), .ZN(
        n18658) );
  XNOR2_X1 U19448 ( .A(n18658), .B(n18532), .ZN(n18267) );
  INV_X1 U19449 ( .A(n18267), .ZN(n16928) );
  XNOR2_X1 U19450 ( .A(n16928), .B(n18176), .ZN(n16939) );
  OAI22_X1 U19451 ( .A1(n16932), .A2(n25031), .B1(n24585), .B2(n17059), .ZN(
        n16930) );
  NAND2_X1 U19452 ( .A1(n16930), .A2(n16929), .ZN(n16934) );
  INV_X1 U19453 ( .A(n17059), .ZN(n16931) );
  NAND2_X1 U19454 ( .A1(n16932), .A2(n16931), .ZN(n16933) );
  XNOR2_X1 U19455 ( .A(n18067), .B(n923), .ZN(n16936) );
  XOR2_X1 U19456 ( .A(n16937), .B(n16936), .Z(n16938) );
  MUX2_X1 U19457 ( .A(n4487), .B(n17407), .S(n16940), .Z(n16943) );
  NOR3_X1 U19458 ( .A1(n17410), .A2(n17615), .A3(n17255), .ZN(n17611) );
  XNOR2_X1 U19460 ( .A(n16946), .B(n18677), .ZN(n16949) );
  XNOR2_X1 U19461 ( .A(n18227), .B(n16947), .ZN(n16948) );
  XNOR2_X1 U19462 ( .A(n16949), .B(n16948), .ZN(n16960) );
  NAND2_X1 U19463 ( .A1(n16952), .A2(n17230), .ZN(n16953) );
  INV_X1 U19464 ( .A(n17791), .ZN(n16959) );
  NOR2_X1 U19465 ( .A1(n17227), .A2(n25433), .ZN(n17416) );
  NAND3_X1 U19466 ( .A1(n16957), .A2(n16956), .A3(n1230), .ZN(n16958) );
  XNOR2_X1 U19467 ( .A(n16959), .B(n18675), .ZN(n18189) );
  INV_X1 U19468 ( .A(n18189), .ZN(n18089) );
  BUF_X2 U19469 ( .A(n17562), .Z(n18923) );
  NAND2_X1 U19470 ( .A1(n16964), .A2(n16962), .ZN(n16968) );
  INV_X1 U19471 ( .A(n17662), .ZN(n16967) );
  NAND2_X1 U19472 ( .A1(n16963), .A2(n24444), .ZN(n17446) );
  INV_X1 U19473 ( .A(n17446), .ZN(n17127) );
  NOR2_X1 U19474 ( .A1(n17439), .A2(n16964), .ZN(n16965) );
  INV_X1 U19475 ( .A(n17661), .ZN(n16966) );
  OAI21_X1 U19476 ( .B1(n16967), .B2(n16966), .A(n23347), .ZN(n16970) );
  NOR2_X1 U19477 ( .A1(n16974), .A2(n17335), .ZN(n16972) );
  NOR2_X1 U19478 ( .A1(n16972), .A2(n16971), .ZN(n16978) );
  NOR2_X1 U19479 ( .A1(n16973), .A2(n376), .ZN(n16975) );
  OAI21_X1 U19480 ( .B1(n16976), .B2(n16975), .A(n16974), .ZN(n16977) );
  NOR2_X1 U19481 ( .A1(n16979), .A2(n16980), .ZN(n16983) );
  OAI21_X1 U19482 ( .B1(n24942), .B2(n17453), .A(n5072), .ZN(n16982) );
  NAND3_X1 U19483 ( .A1(n24942), .A2(n523), .A3(n17451), .ZN(n16981) );
  XNOR2_X1 U19484 ( .A(n18562), .B(n18172), .ZN(n18687) );
  MUX2_X1 U19485 ( .A(n17141), .B(n17137), .S(n17139), .Z(n16987) );
  OAI21_X1 U19486 ( .B1(n16984), .B2(n17144), .A(n17138), .ZN(n16986) );
  INV_X1 U19487 ( .A(n19313), .ZN(n19317) );
  NAND2_X1 U19488 ( .A1(n19317), .A2(n5371), .ZN(n17010) );
  NOR2_X1 U19489 ( .A1(n25214), .A2(n16989), .ZN(n16990) );
  NAND3_X1 U19490 ( .A1(n16991), .A2(n288), .A3(n287), .ZN(n16992) );
  XNOR2_X1 U19493 ( .A(n24536), .B(n18220), .ZN(n16996) );
  XNOR2_X1 U19494 ( .A(n18692), .B(n16996), .ZN(n17008) );
  NAND2_X1 U19495 ( .A1(n17572), .A2(n16998), .ZN(n16999) );
  NAND3_X1 U19496 ( .A1(n17049), .A2(n17053), .A3(n17050), .ZN(n17001) );
  XNOR2_X1 U19497 ( .A(n18200), .B(n18695), .ZN(n17006) );
  XNOR2_X1 U19498 ( .A(n18006), .B(n2033), .ZN(n17005) );
  XNOR2_X1 U19499 ( .A(n17006), .B(n17005), .ZN(n17007) );
  INV_X1 U19500 ( .A(n19312), .ZN(n17009) );
  MUX2_X1 U19501 ( .A(n17011), .B(n17010), .S(n17009), .Z(n17036) );
  MUX2_X1 U19502 ( .A(n17015), .B(n17212), .S(n25200), .Z(n17022) );
  NAND2_X1 U19503 ( .A1(n17016), .A2(n25201), .ZN(n17018) );
  OAI22_X1 U19504 ( .A1(n17018), .A2(n5512), .B1(n17216), .B2(n17017), .ZN(
        n17019) );
  INV_X1 U19505 ( .A(n17019), .ZN(n17020) );
  OAI21_X1 U19506 ( .B1(n17186), .B2(n3602), .A(n17185), .ZN(n17024) );
  XNOR2_X1 U19507 ( .A(n18325), .B(n18096), .ZN(n18704) );
  OAI211_X1 U19508 ( .C1(n17400), .C2(n25003), .A(n17398), .B(n17198), .ZN(
        n17029) );
  INV_X1 U19509 ( .A(n17399), .ZN(n17193) );
  XNOR2_X1 U19510 ( .A(n18451), .B(n4189), .ZN(n17033) );
  NAND2_X1 U19511 ( .A1(n19311), .A2(n19310), .ZN(n18925) );
  NOR2_X1 U19512 ( .A1(n24567), .A2(n20336), .ZN(n20672) );
  NAND2_X1 U19513 ( .A1(n17364), .A2(n17362), .ZN(n17037) );
  XNOR2_X1 U19514 ( .A(n18023), .B(n17041), .ZN(n18349) );
  AOI21_X1 U19515 ( .B1(n17370), .B2(n17044), .A(n17572), .ZN(n17046) );
  NOR3_X1 U19516 ( .A1(n5522), .A2(n17574), .A3(n3371), .ZN(n17045) );
  OR3_X2 U19517 ( .A1(n17576), .A2(n17046), .A3(n17045), .ZN(n17748) );
  INV_X1 U19518 ( .A(n17748), .ZN(n18252) );
  XNOR2_X1 U19519 ( .A(n18252), .B(n18451), .ZN(n17047) );
  XNOR2_X1 U19520 ( .A(n18349), .B(n17047), .ZN(n17074) );
  NAND2_X1 U19521 ( .A1(n17054), .A2(n17059), .ZN(n17055) );
  NAND2_X1 U19522 ( .A1(n17056), .A2(n17055), .ZN(n17058) );
  NOR2_X1 U19523 ( .A1(n17060), .A2(n17059), .ZN(n17064) );
  NOR2_X1 U19524 ( .A1(n24585), .A2(n24398), .ZN(n17063) );
  XNOR2_X1 U19525 ( .A(n17819), .B(n18350), .ZN(n17072) );
  NAND2_X1 U19526 ( .A1(n17068), .A2(n369), .ZN(n17066) );
  XNOR2_X1 U19527 ( .A(n18599), .B(n92), .ZN(n17071) );
  XNOR2_X1 U19528 ( .A(n17071), .B(n17072), .ZN(n17073) );
  AOI21_X1 U19529 ( .B1(n17480), .B2(n17482), .A(n17076), .ZN(n17083) );
  AOI21_X1 U19530 ( .B1(n17079), .B2(n17078), .A(n17077), .ZN(n17080) );
  NOR2_X1 U19531 ( .A1(n25429), .A2(n17080), .ZN(n17082) );
  XNOR2_X1 U19533 ( .A(n17680), .B(n18483), .ZN(n17953) );
  INV_X1 U19534 ( .A(n17084), .ZN(n17091) );
  XNOR2_X1 U19535 ( .A(n17953), .B(n17092), .ZN(n17113) );
  AOI22_X1 U19536 ( .A1(n17093), .A2(n17484), .B1(n17735), .B2(n17731), .ZN(
        n17097) );
  NAND2_X1 U19537 ( .A1(n17735), .A2(n17094), .ZN(n17096) );
  OR2_X1 U19538 ( .A1(n17690), .A2(n17486), .ZN(n17095) );
  NAND2_X1 U19539 ( .A1(n17120), .A2(n17118), .ZN(n17098) );
  AND3_X1 U19540 ( .A1(n17099), .A2(n17116), .A3(n17098), .ZN(n17106) );
  NAND3_X1 U19543 ( .A1(n17114), .A2(n16572), .A3(n25357), .ZN(n17104) );
  OAI211_X2 U19544 ( .C1(n17106), .C2(n2580), .A(n17105), .B(n17104), .ZN(
        n18032) );
  XNOR2_X1 U19545 ( .A(n18356), .B(n18032), .ZN(n18268) );
  NAND2_X1 U19547 ( .A1(n17132), .A2(n17131), .ZN(n17109) );
  XNOR2_X1 U19548 ( .A(n17832), .B(n1935), .ZN(n17110) );
  NOR2_X1 U19550 ( .A1(n18934), .A2(n17496), .ZN(n17495) );
  OAI211_X1 U19551 ( .C1(n17116), .C2(n17115), .A(n17114), .B(n17118), .ZN(
        n17117) );
  INV_X1 U19552 ( .A(n17117), .ZN(n17124) );
  NOR2_X1 U19553 ( .A1(n17119), .A2(n17118), .ZN(n17121) );
  OAI211_X1 U19555 ( .C1(n17125), .C2(n24444), .A(n17439), .B(n17442), .ZN(
        n17126) );
  OAI21_X1 U19556 ( .B1(n17128), .B2(n17127), .A(n17126), .ZN(n18276) );
  XNOR2_X1 U19557 ( .A(n18276), .B(n17958), .ZN(n17136) );
  OAI211_X1 U19558 ( .C1(n17132), .C2(n17131), .A(n4684), .B(n17130), .ZN(
        n17133) );
  XNOR2_X1 U19559 ( .A(n18341), .B(n1826), .ZN(n17135) );
  XNOR2_X1 U19560 ( .A(n17136), .B(n17135), .ZN(n17154) );
  NOR2_X1 U19561 ( .A1(n17138), .A2(n17137), .ZN(n17143) );
  AOI21_X1 U19562 ( .B1(n17145), .B2(n17140), .A(n17139), .ZN(n17142) );
  NOR2_X1 U19563 ( .A1(n17145), .A2(n17144), .ZN(n17146) );
  NAND2_X1 U19565 ( .A1(n17460), .A2(n17451), .ZN(n17151) );
  NAND2_X1 U19566 ( .A1(n523), .A2(n17450), .ZN(n17148) );
  XNOR2_X1 U19569 ( .A(n18694), .B(n18060), .ZN(n18367) );
  INV_X1 U19570 ( .A(n18367), .ZN(n17693) );
  XNOR2_X1 U19571 ( .A(n17693), .B(n18475), .ZN(n17153) );
  XNOR2_X2 U19572 ( .A(n17153), .B(n17154), .ZN(n19326) );
  NAND3_X1 U19573 ( .A1(n17158), .A2(n17157), .A3(n17156), .ZN(n17162) );
  INV_X1 U19574 ( .A(n17159), .ZN(n17161) );
  NAND3_X1 U19576 ( .A1(n17165), .A2(n17164), .A3(n17163), .ZN(n17168) );
  XNOR2_X1 U19577 ( .A(n25380), .B(n3093), .ZN(n17178) );
  XNOR2_X1 U19579 ( .A(n17178), .B(n17806), .ZN(n17191) );
  AND2_X1 U19580 ( .A1(n3602), .A2(n17184), .ZN(n17188) );
  NOR2_X1 U19581 ( .A1(n17185), .A2(n17391), .ZN(n17187) );
  AOI22_X1 U19582 ( .A1(n17188), .A2(n17389), .B1(n17187), .B2(n3604), .ZN(
        n17189) );
  OAI21_X2 U19583 ( .B1(n17190), .B2(n16203), .A(n17189), .ZN(n18295) );
  XNOR2_X1 U19584 ( .A(n17191), .B(n18387), .ZN(n17222) );
  MUX2_X1 U19585 ( .A(n17198), .B(n17195), .S(n17192), .Z(n17194) );
  AND2_X1 U19586 ( .A1(n17194), .A2(n17193), .ZN(n17201) );
  NAND2_X1 U19587 ( .A1(n4039), .A2(n17400), .ZN(n17199) );
  OAI22_X1 U19588 ( .A1(n17199), .A2(n17198), .B1(n17197), .B2(n17196), .ZN(
        n17200) );
  INV_X1 U19589 ( .A(n17202), .ZN(n17204) );
  NAND2_X1 U19590 ( .A1(n17342), .A2(n17346), .ZN(n17203) );
  AOI21_X1 U19591 ( .B1(n17204), .B2(n17203), .A(n17347), .ZN(n17205) );
  NOR2_X1 U19592 ( .A1(n17206), .A2(n17205), .ZN(n17220) );
  NAND2_X1 U19594 ( .A1(n25201), .A2(n17208), .ZN(n17209) );
  NAND3_X1 U19595 ( .A1(n17210), .A2(n5512), .A3(n17209), .ZN(n17219) );
  NAND3_X1 U19596 ( .A1(n24391), .A2(n17212), .A3(n17211), .ZN(n17218) );
  NAND3_X1 U19597 ( .A1(n17216), .A2(n25201), .A3(n17214), .ZN(n17217) );
  XNOR2_X1 U19598 ( .A(n17220), .B(n18187), .ZN(n18459) );
  XNOR2_X1 U19599 ( .A(n18290), .B(n18459), .ZN(n17221) );
  XNOR2_X1 U19600 ( .A(n17222), .B(n17221), .ZN(n17497) );
  NOR2_X1 U19602 ( .A1(n24583), .A2(n19326), .ZN(n17223) );
  NOR2_X1 U19603 ( .A1(n17495), .A2(n17223), .ZN(n17310) );
  XNOR2_X1 U19604 ( .A(n18261), .B(n18666), .ZN(n18380) );
  MUX2_X1 U19605 ( .A(n17288), .B(n17283), .S(n17229), .Z(n17233) );
  NAND2_X1 U19606 ( .A1(n17283), .A2(n17229), .ZN(n17286) );
  MUX2_X1 U19607 ( .A(n17286), .B(n17231), .S(n17230), .Z(n17232) );
  XNOR2_X1 U19608 ( .A(n18239), .B(n18665), .ZN(n17234) );
  XNOR2_X1 U19609 ( .A(n18380), .B(n17234), .ZN(n17263) );
  INV_X1 U19610 ( .A(n17235), .ZN(n17239) );
  NAND2_X1 U19611 ( .A1(n17239), .A2(n17238), .ZN(n17246) );
  AND2_X1 U19612 ( .A1(n17346), .A2(n17344), .ZN(n17245) );
  MUX2_X1 U19613 ( .A(n17242), .B(n17241), .S(n15314), .Z(n17243) );
  NAND2_X1 U19614 ( .A1(n17347), .A2(n17243), .ZN(n17244) );
  NAND3_X1 U19616 ( .A1(n17275), .A2(n17277), .A3(n17249), .ZN(n17250) );
  NAND3_X1 U19617 ( .A1(n17407), .A2(n17607), .A3(n17408), .ZN(n17256) );
  NOR2_X1 U19618 ( .A1(n4487), .A2(n17257), .ZN(n17258) );
  NOR2_X2 U19619 ( .A1(n17259), .A2(n17258), .ZN(n18489) );
  XNOR2_X1 U19620 ( .A(n18489), .B(n1726), .ZN(n17260) );
  XNOR2_X1 U19621 ( .A(n17261), .B(n17260), .ZN(n17262) );
  XNOR2_X1 U19622 ( .A(n17263), .B(n17262), .ZN(n17264) );
  INV_X1 U19623 ( .A(n17264), .ZN(n18933) );
  NOR2_X1 U19624 ( .A1(n17264), .A2(n17496), .ZN(n19331) );
  INV_X1 U19625 ( .A(n17319), .ZN(n17265) );
  NOR2_X1 U19626 ( .A1(n17267), .A2(n17266), .ZN(n17270) );
  INV_X1 U19627 ( .A(n17326), .ZN(n17323) );
  NOR2_X1 U19628 ( .A1(n17322), .A2(n17323), .ZN(n17268) );
  AND2_X1 U19630 ( .A1(n17273), .A2(n17276), .ZN(n17271) );
  NAND2_X1 U19631 ( .A1(n17272), .A2(n17271), .ZN(n17281) );
  NOR2_X1 U19632 ( .A1(n17277), .A2(n17276), .ZN(n17278) );
  NAND2_X1 U19633 ( .A1(n3855), .A2(n17278), .ZN(n17280) );
  AND2_X1 U19634 ( .A1(n17285), .A2(n17286), .ZN(n17291) );
  XNOR2_X1 U19636 ( .A(n18512), .B(n2058), .ZN(n17294) );
  XNOR2_X1 U19637 ( .A(n17294), .B(n17520), .ZN(n17295) );
  XNOR2_X1 U19638 ( .A(n17295), .B(n18372), .ZN(n17308) );
  INV_X1 U19639 ( .A(n17296), .ZN(n17298) );
  NAND2_X1 U19640 ( .A1(n17298), .A2(n17297), .ZN(n17301) );
  XNOR2_X1 U19642 ( .A(n18465), .B(n25411), .ZN(n17306) );
  XNOR2_X1 U19643 ( .A(n17306), .B(n5300), .ZN(n17307) );
  OAI21_X1 U19644 ( .B1(n19331), .B2(n3034), .A(n24583), .ZN(n17309) );
  INV_X1 U19645 ( .A(n20668), .ZN(n20671) );
  MUX2_X1 U19646 ( .A(n17311), .B(n20672), .S(n20671), .Z(n17494) );
  NOR2_X1 U19647 ( .A1(n20670), .A2(n20335), .ZN(n19709) );
  NAND2_X1 U19648 ( .A1(n17315), .A2(n17314), .ZN(n17317) );
  XNOR2_X1 U19649 ( .A(n18448), .B(n17819), .ZN(n18422) );
  INV_X1 U19650 ( .A(n18447), .ZN(n17327) );
  XNOR2_X1 U19651 ( .A(n17328), .B(n17327), .ZN(n17329) );
  XNOR2_X1 U19652 ( .A(n17329), .B(n18422), .ZN(n17340) );
  NAND2_X1 U19653 ( .A1(n3817), .A2(n17335), .ZN(n17338) );
  XNOR2_X1 U19654 ( .A(n18423), .B(n18599), .ZN(n17506) );
  XNOR2_X1 U19655 ( .A(n17506), .B(n18214), .ZN(n17657) );
  XNOR2_X1 U19656 ( .A(n17340), .B(n17657), .ZN(n18761) );
  AOI21_X1 U19657 ( .B1(n17343), .B2(n17342), .A(n17341), .ZN(n17345) );
  NOR3_X1 U19658 ( .A1(n17348), .A2(n17347), .A3(n17346), .ZN(n17349) );
  NOR2_X1 U19659 ( .A1(n17350), .A2(n17349), .ZN(n17359) );
  NAND2_X1 U19660 ( .A1(n17357), .A2(n17351), .ZN(n17355) );
  NAND2_X1 U19661 ( .A1(n17353), .A2(n25491), .ZN(n17354) );
  OAI211_X1 U19662 ( .C1(n17357), .C2(n17356), .A(n17355), .B(n17354), .ZN(
        n17358) );
  XNOR2_X1 U19663 ( .A(n17359), .B(n18123), .ZN(n17642) );
  XNOR2_X1 U19664 ( .A(n17642), .B(n17360), .ZN(n17377) );
  NOR2_X1 U19665 ( .A1(n17362), .A2(n25215), .ZN(n17365) );
  NOR2_X1 U19666 ( .A1(n17366), .A2(n370), .ZN(n17367) );
  XNOR2_X1 U19667 ( .A(n18491), .B(n18669), .ZN(n17375) );
  NAND2_X1 U19668 ( .A1(n24471), .A2(n17368), .ZN(n17369) );
  NOR2_X1 U19669 ( .A1(n24471), .A2(n17574), .ZN(n17372) );
  NAND2_X1 U19670 ( .A1(n17378), .A2(n17425), .ZN(n17380) );
  MUX2_X1 U19671 ( .A(n17426), .B(n17380), .S(n17379), .Z(n17385) );
  NAND2_X1 U19672 ( .A1(n17423), .A2(n17381), .ZN(n17383) );
  NOR2_X1 U19673 ( .A1(n17383), .A2(n17382), .ZN(n17384) );
  NOR2_X2 U19674 ( .A1(n17385), .A2(n17384), .ZN(n18407) );
  INV_X1 U19675 ( .A(n17389), .ZN(n17388) );
  MUX2_X1 U19676 ( .A(n17391), .B(n17390), .S(n17389), .Z(n17392) );
  XNOR2_X1 U19678 ( .A(n18531), .B(n18102), .ZN(n18232) );
  INV_X1 U19679 ( .A(n18232), .ZN(n17394) );
  XNOR2_X1 U19680 ( .A(n17394), .B(n17648), .ZN(n17405) );
  OAI21_X1 U19681 ( .B1(n17397), .B2(n17396), .A(n17395), .ZN(n17402) );
  XNOR2_X1 U19683 ( .A(n17832), .B(n18484), .ZN(n18404) );
  XNOR2_X1 U19684 ( .A(n18660), .B(n688), .ZN(n17403) );
  XNOR2_X1 U19685 ( .A(n18404), .B(n17403), .ZN(n17404) );
  XNOR2_X2 U19686 ( .A(n17405), .B(n17404), .ZN(n19531) );
  INV_X1 U19687 ( .A(n17881), .ZN(n17406) );
  XNOR2_X1 U19688 ( .A(n18311), .B(n17406), .ZN(n17660) );
  OAI22_X1 U19689 ( .A1(n17410), .A2(n17608), .B1(n17407), .B2(n17607), .ZN(
        n17411) );
  INV_X1 U19690 ( .A(n17408), .ZN(n17612) );
  XNOR2_X1 U19691 ( .A(n18128), .B(n18308), .ZN(n17412) );
  XNOR2_X1 U19692 ( .A(n17660), .B(n17412), .ZN(n17432) );
  NOR2_X1 U19693 ( .A1(n17414), .A2(n17413), .ZN(n17415) );
  INV_X1 U19694 ( .A(n18512), .ZN(n17420) );
  XNOR2_X1 U19695 ( .A(n18466), .B(n17420), .ZN(n17967) );
  NAND3_X1 U19697 ( .A1(n17423), .A2(n17422), .A3(n5409), .ZN(n17428) );
  OAI21_X1 U19698 ( .B1(n17426), .B2(n17425), .A(n17424), .ZN(n17427) );
  INV_X1 U19700 ( .A(n18515), .ZN(n18467) );
  XNOR2_X1 U19701 ( .A(n17967), .B(n17430), .ZN(n17431) );
  XNOR2_X1 U19702 ( .A(n17432), .B(n17431), .ZN(n19145) );
  INV_X1 U19703 ( .A(n19145), .ZN(n19269) );
  NOR2_X1 U19704 ( .A1(n17439), .A2(n24444), .ZN(n17443) );
  NOR2_X1 U19705 ( .A1(n17446), .A2(n17445), .ZN(n17447) );
  XNOR2_X1 U19706 ( .A(n18456), .B(n17806), .ZN(n18415) );
  XNOR2_X1 U19708 ( .A(n18225), .B(n18415), .ZN(n17471) );
  XNOR2_X1 U19709 ( .A(n24488), .B(n18388), .ZN(n17469) );
  XNOR2_X1 U19710 ( .A(n25379), .B(n2036), .ZN(n17468) );
  XNOR2_X1 U19711 ( .A(n17469), .B(n17468), .ZN(n17470) );
  XNOR2_X1 U19712 ( .A(n17471), .B(n17470), .ZN(n18762) );
  AND2_X1 U19713 ( .A1(n19269), .A2(n19534), .ZN(n19533) );
  XNOR2_X1 U19715 ( .A(n18473), .B(n17476), .ZN(n18219) );
  INV_X1 U19716 ( .A(n18219), .ZN(n17489) );
  INV_X1 U19717 ( .A(n17477), .ZN(n17483) );
  AND2_X1 U19718 ( .A1(n25472), .A2(n17485), .ZN(n17688) );
  NAND2_X1 U19719 ( .A1(n17688), .A2(n17687), .ZN(n17487) );
  NAND3_X1 U19720 ( .A1(n17690), .A2(n17686), .A3(n17487), .ZN(n17488) );
  XNOR2_X1 U19721 ( .A(n18365), .B(n17488), .ZN(n18478) );
  XNOR2_X1 U19722 ( .A(n17489), .B(n18478), .ZN(n17493) );
  XNOR2_X1 U19723 ( .A(n17958), .B(n18693), .ZN(n17491) );
  XNOR2_X1 U19724 ( .A(n18341), .B(n21204), .ZN(n17490) );
  XNOR2_X1 U19725 ( .A(n17491), .B(n17490), .ZN(n17492) );
  INV_X1 U19727 ( .A(n20338), .ZN(n20341) );
  NAND2_X1 U19731 ( .A1(n25566), .A2(n19329), .ZN(n17944) );
  AOI21_X1 U19732 ( .B1(n19327), .B2(n17944), .A(n17495), .ZN(n17500) );
  INV_X1 U19733 ( .A(n17496), .ZN(n19328) );
  INV_X1 U19734 ( .A(n17498), .ZN(n17499) );
  AOI21_X1 U19735 ( .B1(n19132), .B2(n18767), .A(n18766), .ZN(n17503) );
  INV_X1 U19736 ( .A(n19132), .ZN(n19303) );
  AND2_X1 U19737 ( .A1(n19303), .A2(n19133), .ZN(n18768) );
  INV_X1 U19738 ( .A(n18768), .ZN(n17502) );
  NAND2_X1 U19739 ( .A1(n19307), .A2(n24324), .ZN(n17501) );
  XNOR2_X1 U19740 ( .A(n17504), .B(n18446), .ZN(n17505) );
  INV_X1 U19741 ( .A(n18420), .ZN(n18022) );
  XNOR2_X1 U19742 ( .A(n18022), .B(n17816), .ZN(n18521) );
  XNOR2_X1 U19743 ( .A(n18521), .B(n17505), .ZN(n17508) );
  XNOR2_X1 U19744 ( .A(n18098), .B(n17506), .ZN(n17507) );
  XNOR2_X1 U19745 ( .A(n17681), .B(n17993), .ZN(n17833) );
  INV_X1 U19746 ( .A(n17833), .ZN(n17509) );
  XNOR2_X1 U19747 ( .A(n17509), .B(n17648), .ZN(n17512) );
  XNOR2_X1 U19748 ( .A(n18103), .B(n2241), .ZN(n17510) );
  XNOR2_X1 U19749 ( .A(n18405), .B(n17510), .ZN(n17511) );
  XNOR2_X1 U19750 ( .A(n17726), .B(n18621), .ZN(n17514) );
  XNOR2_X1 U19751 ( .A(n17839), .B(n18121), .ZN(n17513) );
  XNOR2_X1 U19752 ( .A(n17514), .B(n17513), .ZN(n17519) );
  XNOR2_X1 U19753 ( .A(n17515), .B(n912), .ZN(n17517) );
  XNOR2_X1 U19754 ( .A(n18123), .B(n18541), .ZN(n17516) );
  XNOR2_X1 U19755 ( .A(n17517), .B(n17516), .ZN(n17518) );
  XNOR2_X1 U19756 ( .A(n17519), .B(n17518), .ZN(n18929) );
  NAND2_X1 U19757 ( .A1(n3653), .A2(n18929), .ZN(n17553) );
  XNOR2_X1 U19758 ( .A(n17811), .B(n1854), .ZN(n17521) );
  XNOR2_X1 U19759 ( .A(n18627), .B(n17521), .ZN(n17531) );
  OAI21_X1 U19760 ( .B1(n17524), .B2(n17523), .A(n17522), .ZN(n17526) );
  OAI21_X1 U19761 ( .B1(n17527), .B2(n17526), .A(n17525), .ZN(n17880) );
  XNOR2_X1 U19762 ( .A(n18370), .B(n17880), .ZN(n17529) );
  XNOR2_X1 U19763 ( .A(n18042), .B(n18128), .ZN(n18399) );
  INV_X1 U19764 ( .A(n18399), .ZN(n17528) );
  XNOR2_X1 U19765 ( .A(n17529), .B(n17528), .ZN(n17530) );
  XNOR2_X1 U19766 ( .A(n17530), .B(n17531), .ZN(n19295) );
  XNOR2_X1 U19767 ( .A(n25379), .B(n17532), .ZN(n18635) );
  INV_X1 U19768 ( .A(n18635), .ZN(n18160) );
  XNOR2_X1 U19769 ( .A(n18160), .B(n17533), .ZN(n17537) );
  XNOR2_X1 U19770 ( .A(n17807), .B(n18388), .ZN(n17535) );
  XNOR2_X1 U19771 ( .A(n18190), .B(n2120), .ZN(n17534) );
  XNOR2_X1 U19772 ( .A(n17535), .B(n17534), .ZN(n17536) );
  XNOR2_X2 U19773 ( .A(n17537), .B(n17536), .ZN(n19296) );
  OAI211_X1 U19774 ( .C1(n19297), .C2(n18929), .A(n24457), .B(n19296), .ZN(
        n17551) );
  INV_X1 U19775 ( .A(n18929), .ZN(n18967) );
  NAND3_X1 U19776 ( .A1(n17540), .A2(n17539), .A3(n17538), .ZN(n17543) );
  INV_X1 U19777 ( .A(n17541), .ZN(n17542) );
  XNOR2_X1 U19779 ( .A(n18472), .B(n17757), .ZN(n17827) );
  XNOR2_X1 U19780 ( .A(n18341), .B(n18431), .ZN(n18648) );
  INV_X1 U19781 ( .A(n18648), .ZN(n17545) );
  XNOR2_X1 U19782 ( .A(n17545), .B(n17827), .ZN(n17549) );
  XNOR2_X1 U19783 ( .A(n18365), .B(n3062), .ZN(n17547) );
  XNOR2_X1 U19784 ( .A(n18198), .B(n18429), .ZN(n17546) );
  XNOR2_X1 U19785 ( .A(n17547), .B(n17546), .ZN(n17548) );
  XNOR2_X1 U19786 ( .A(n17549), .B(n17548), .ZN(n18927) );
  INV_X1 U19789 ( .A(n19531), .ZN(n19272) );
  NOR2_X1 U19790 ( .A1(n17559), .A2(n1299), .ZN(n17555) );
  NOR2_X1 U19791 ( .A1(n18919), .A2(n17555), .ZN(n17561) );
  INV_X1 U19792 ( .A(n17556), .ZN(n18756) );
  NAND2_X1 U19794 ( .A1(n17558), .A2(n18756), .ZN(n17560) );
  AND2_X1 U19795 ( .A1(n20322), .A2(n20316), .ZN(n17566) );
  INV_X1 U19796 ( .A(n17562), .ZN(n19315) );
  NAND2_X1 U19797 ( .A1(n18923), .A2(n19313), .ZN(n17563) );
  INV_X1 U19798 ( .A(n19309), .ZN(n18841) );
  NAND2_X1 U19799 ( .A1(n18923), .A2(n24912), .ZN(n19318) );
  XNOR2_X1 U19800 ( .A(n25202), .B(n21273), .ZN(n17952) );
  INV_X1 U19801 ( .A(n18074), .ZN(n18600) );
  XNOR2_X1 U19802 ( .A(n18351), .B(n18600), .ZN(n17569) );
  XNOR2_X1 U19803 ( .A(n18325), .B(n17819), .ZN(n18524) );
  XNOR2_X1 U19804 ( .A(n18524), .B(n17569), .ZN(n17580) );
  INV_X1 U19805 ( .A(n17900), .ZN(n17570) );
  XNOR2_X1 U19806 ( .A(n17570), .B(n23225), .ZN(n17578) );
  NOR2_X1 U19807 ( .A1(n24471), .A2(n17572), .ZN(n17575) );
  XNOR2_X1 U19808 ( .A(n17580), .B(n17579), .ZN(n18735) );
  INV_X1 U19809 ( .A(n18735), .ZN(n19482) );
  XNOR2_X1 U19810 ( .A(n17581), .B(n17919), .ZN(n18360) );
  XNOR2_X1 U19811 ( .A(n17832), .B(n17582), .ZN(n18528) );
  XNOR2_X1 U19812 ( .A(n18360), .B(n18528), .ZN(n17586) );
  XNOR2_X1 U19813 ( .A(n24565), .B(n18610), .ZN(n17584) );
  XNOR2_X1 U19814 ( .A(n18032), .B(n494), .ZN(n17583) );
  XNOR2_X1 U19815 ( .A(n17584), .B(n17583), .ZN(n17585) );
  XNOR2_X1 U19816 ( .A(n17587), .B(n18549), .ZN(n17588) );
  XNOR2_X1 U19817 ( .A(n18646), .B(n18695), .ZN(n18196) );
  XNOR2_X1 U19818 ( .A(n18512), .B(n23699), .ZN(n17589) );
  XNOR2_X1 U19819 ( .A(n17589), .B(n18513), .ZN(n17591) );
  OAI21_X1 U19820 ( .B1(n19482), .B2(n19477), .A(n17594), .ZN(n17896) );
  INV_X1 U19821 ( .A(n17601), .ZN(n17602) );
  XNOR2_X1 U19822 ( .A(n16910), .B(n18382), .ZN(n17604) );
  INV_X1 U19823 ( .A(n18665), .ZN(n17603) );
  XNOR2_X1 U19824 ( .A(n17604), .B(n17603), .ZN(n18040) );
  INV_X1 U19825 ( .A(n18040), .ZN(n17605) );
  XNOR2_X1 U19826 ( .A(n17606), .B(n17605), .ZN(n18730) );
  INV_X1 U19827 ( .A(n18730), .ZN(n18848) );
  NAND2_X1 U19828 ( .A1(n17608), .A2(n17607), .ZN(n17616) );
  NOR2_X1 U19829 ( .A1(n17611), .A2(n17610), .ZN(n17618) );
  NAND2_X1 U19830 ( .A1(n17613), .A2(n17612), .ZN(n17614) );
  NAND3_X1 U19831 ( .A1(n17616), .A2(n17615), .A3(n17614), .ZN(n17617) );
  XNOR2_X1 U19833 ( .A(n17619), .B(n18018), .ZN(n17636) );
  INV_X1 U19834 ( .A(n17620), .ZN(n17621) );
  NOR2_X1 U19835 ( .A1(n17622), .A2(n17621), .ZN(n17627) );
  INV_X1 U19836 ( .A(n17623), .ZN(n17625) );
  NOR2_X1 U19837 ( .A1(n17625), .A2(n17624), .ZN(n17626) );
  AOI21_X1 U19838 ( .B1(n17627), .B2(n17626), .A(n17629), .ZN(n17628) );
  NAND2_X1 U19839 ( .A1(n17628), .A2(n17632), .ZN(n17631) );
  NAND3_X1 U19840 ( .A1(n17633), .A2(n2561), .A3(n17629), .ZN(n17630) );
  OAI211_X1 U19841 ( .C1(n17633), .C2(n17632), .A(n17631), .B(n17630), .ZN(
        n18017) );
  INV_X1 U19842 ( .A(n18017), .ZN(n17634) );
  XOR2_X1 U19843 ( .A(n18157), .B(n17634), .Z(n17635) );
  XNOR2_X1 U19844 ( .A(n17636), .B(n17635), .ZN(n17639) );
  XNOR2_X1 U19845 ( .A(n18188), .B(n24433), .ZN(n17638) );
  NAND2_X1 U19846 ( .A1(n19482), .A2(n17640), .ZN(n17641) );
  XNOR2_X1 U19847 ( .A(n17905), .B(n18541), .ZN(n17981) );
  XNOR2_X1 U19848 ( .A(n17642), .B(n17981), .ZN(n17647) );
  XNOR2_X1 U19849 ( .A(n25000), .B(n17643), .ZN(n17645) );
  XNOR2_X1 U19850 ( .A(n17645), .B(n17644), .ZN(n17646) );
  XNOR2_X1 U19851 ( .A(n18233), .B(n18067), .ZN(n17918) );
  XNOR2_X1 U19852 ( .A(n18335), .B(n1827), .ZN(n17651) );
  XNOR2_X1 U19853 ( .A(n17649), .B(n18530), .ZN(n17650) );
  XNOR2_X1 U19854 ( .A(n17651), .B(n17650), .ZN(n17652) );
  XNOR2_X1 U19855 ( .A(n18149), .B(n2040), .ZN(n17654) );
  XNOR2_X1 U19857 ( .A(n17654), .B(n18601), .ZN(n17656) );
  XNOR2_X1 U19858 ( .A(n18022), .B(n17899), .ZN(n17655) );
  XNOR2_X1 U19859 ( .A(n17656), .B(n17655), .ZN(n17659) );
  INV_X1 U19860 ( .A(n17657), .ZN(n17658) );
  INV_X1 U19861 ( .A(n18312), .ZN(n17709) );
  XNOR2_X1 U19862 ( .A(n17709), .B(n17969), .ZN(n18626) );
  XNOR2_X1 U19863 ( .A(n18637), .B(n17791), .ZN(n17915) );
  XNOR2_X1 U19864 ( .A(n18413), .B(n17915), .ZN(n17668) );
  XNOR2_X1 U19865 ( .A(n25493), .B(n24337), .ZN(n17666) );
  XNOR2_X1 U19866 ( .A(n25380), .B(n889), .ZN(n17665) );
  XNOR2_X1 U19867 ( .A(n17666), .B(n17665), .ZN(n17667) );
  XNOR2_X1 U19869 ( .A(n18341), .B(n18365), .ZN(n17670) );
  XNOR2_X1 U19870 ( .A(n17476), .B(n22986), .ZN(n17669) );
  XNOR2_X1 U19871 ( .A(n17670), .B(n17669), .ZN(n17673) );
  INV_X1 U19872 ( .A(n17863), .ZN(n17671) );
  XNOR2_X1 U19873 ( .A(n17671), .B(n18200), .ZN(n17672) );
  XNOR2_X1 U19874 ( .A(n18429), .B(n17931), .ZN(n17963) );
  NAND2_X1 U19875 ( .A1(n25440), .A2(n19346), .ZN(n17674) );
  XNOR2_X1 U19877 ( .A(n18456), .B(n18636), .ZN(n17851) );
  XNOR2_X1 U19878 ( .A(n17851), .B(n17676), .ZN(n17678) );
  INV_X1 U19879 ( .A(n18387), .ZN(n17677) );
  XNOR2_X1 U19881 ( .A(n17681), .B(n17680), .ZN(n18481) );
  XNOR2_X1 U19884 ( .A(n18481), .B(n17994), .ZN(n17685) );
  XNOR2_X1 U19885 ( .A(n18269), .B(n18335), .ZN(n18616) );
  XNOR2_X1 U19886 ( .A(n18659), .B(n1739), .ZN(n17683) );
  XNOR2_X1 U19887 ( .A(n18616), .B(n17683), .ZN(n17684) );
  OAI22_X1 U19889 ( .A1(n17689), .A2(n17688), .B1(n17687), .B2(n17733), .ZN(
        n17691) );
  XNOR2_X1 U19890 ( .A(n18004), .B(n18472), .ZN(n17692) );
  XNOR2_X1 U19891 ( .A(n17693), .B(n17692), .ZN(n17697) );
  XNOR2_X1 U19892 ( .A(n17863), .B(n18220), .ZN(n17695) );
  XNOR2_X1 U19893 ( .A(n18431), .B(n2087), .ZN(n17694) );
  XNOR2_X1 U19894 ( .A(n17695), .B(n17694), .ZN(n17696) );
  INV_X1 U19896 ( .A(n18349), .ZN(n17699) );
  XNOR2_X1 U19897 ( .A(n18601), .B(n18446), .ZN(n17698) );
  XNOR2_X1 U19898 ( .A(n17699), .B(n17698), .ZN(n17703) );
  XNOR2_X1 U19899 ( .A(n18605), .B(n812), .ZN(n17700) );
  XNOR2_X1 U19900 ( .A(n17701), .B(n17700), .ZN(n17702) );
  NAND2_X1 U19903 ( .A1(n19037), .A2(n19451), .ZN(n17712) );
  XNOR2_X1 U19904 ( .A(n18261), .B(n1855), .ZN(n17705) );
  XNOR2_X1 U19905 ( .A(n17705), .B(n18666), .ZN(n17706) );
  XNOR2_X1 U19906 ( .A(n17706), .B(n18619), .ZN(n17708) );
  XNOR2_X1 U19908 ( .A(n18397), .B(n23620), .ZN(n17710) );
  XNOR2_X1 U19910 ( .A(n18290), .B(n18188), .ZN(n17715) );
  XNOR2_X1 U19911 ( .A(n17911), .B(n17715), .ZN(n17719) );
  XNOR2_X1 U19912 ( .A(n17807), .B(n18633), .ZN(n17717) );
  XNOR2_X1 U19913 ( .A(n17716), .B(n17717), .ZN(n17718) );
  XNOR2_X1 U19914 ( .A(n18270), .B(n18032), .ZN(n18656) );
  INV_X1 U19915 ( .A(n17720), .ZN(n18104) );
  XNOR2_X1 U19916 ( .A(n18104), .B(n641), .ZN(n17721) );
  XNOR2_X1 U19917 ( .A(n18656), .B(n17721), .ZN(n17725) );
  XNOR2_X1 U19918 ( .A(n17993), .B(n18611), .ZN(n17723) );
  XNOR2_X1 U19919 ( .A(n17723), .B(n17722), .ZN(n17724) );
  NOR2_X1 U19920 ( .A1(n19389), .A2(n24451), .ZN(n19109) );
  INV_X1 U19921 ( .A(n19109), .ZN(n19387) );
  XNOR2_X1 U19922 ( .A(n17726), .B(n18665), .ZN(n17727) );
  XNOR2_X1 U19923 ( .A(n18124), .B(n18240), .ZN(n18318) );
  XNOR2_X1 U19924 ( .A(n18318), .B(n17727), .ZN(n17743) );
  MUX2_X1 U19925 ( .A(n17730), .B(n17729), .S(n25472), .Z(n17732) );
  NOR2_X1 U19926 ( .A1(n17732), .A2(n17731), .ZN(n17739) );
  NOR2_X1 U19927 ( .A1(n17734), .A2(n17733), .ZN(n17736) );
  MUX2_X1 U19928 ( .A(n17737), .B(n17736), .S(n17735), .Z(n17738) );
  NOR2_X1 U19929 ( .A1(n17739), .A2(n17738), .ZN(n17740) );
  XNOR2_X1 U19930 ( .A(n18262), .B(n17740), .ZN(n18671) );
  XNOR2_X1 U19931 ( .A(n18382), .B(n3155), .ZN(n17741) );
  XNOR2_X1 U19932 ( .A(n18671), .B(n17741), .ZN(n17742) );
  XNOR2_X1 U19933 ( .A(n17743), .B(n17742), .ZN(n19021) );
  XNOR2_X1 U19934 ( .A(n18172), .B(n18370), .ZN(n17745) );
  XNOR2_X1 U19935 ( .A(n18375), .B(n2746), .ZN(n17744) );
  XNOR2_X1 U19936 ( .A(n17744), .B(n17745), .ZN(n17747) );
  XNOR2_X1 U19937 ( .A(n18557), .B(n18129), .ZN(n18309) );
  XNOR2_X1 U19938 ( .A(n18309), .B(n18683), .ZN(n17746) );
  INV_X1 U19939 ( .A(n19217), .ZN(n19388) );
  OAI22_X1 U19940 ( .A1(n19387), .A2(n17762), .B1(n19389), .B2(n19388), .ZN(
        n17766) );
  NAND2_X1 U19941 ( .A1(n19390), .A2(n17762), .ZN(n17764) );
  XNOR2_X1 U19942 ( .A(n17748), .B(n18351), .ZN(n18024) );
  INV_X1 U19943 ( .A(n18024), .ZN(n17749) );
  XNOR2_X1 U19944 ( .A(n17897), .B(n17749), .ZN(n17754) );
  INV_X1 U19945 ( .A(n17816), .ZN(n17750) );
  XNOR2_X1 U19946 ( .A(n18602), .B(n17750), .ZN(n17752) );
  XNOR2_X1 U19947 ( .A(n18096), .B(n2739), .ZN(n17751) );
  XNOR2_X1 U19948 ( .A(n17752), .B(n17751), .ZN(n17753) );
  INV_X1 U19949 ( .A(n18277), .ZN(n17859) );
  XNOR2_X1 U19951 ( .A(n17755), .B(n17859), .ZN(n17932) );
  INV_X1 U19952 ( .A(n17757), .ZN(n18506) );
  XNOR2_X1 U19953 ( .A(n18197), .B(n18506), .ZN(n17759) );
  XNOR2_X1 U19954 ( .A(n18476), .B(n2477), .ZN(n17758) );
  XNOR2_X1 U19955 ( .A(n17759), .B(n17758), .ZN(n17760) );
  INV_X1 U19958 ( .A(n18146), .ZN(n17768) );
  XNOR2_X1 U19960 ( .A(n18418), .B(n859), .ZN(n17769) );
  XNOR2_X1 U19961 ( .A(n17769), .B(n18447), .ZN(n17770) );
  XNOR2_X1 U19962 ( .A(n17770), .B(n18573), .ZN(n17774) );
  XNOR2_X1 U19963 ( .A(n17772), .B(n17771), .ZN(n17773) );
  XNOR2_X2 U19964 ( .A(n17774), .B(n17773), .ZN(n19376) );
  INV_X1 U19965 ( .A(n18032), .ZN(n17775) );
  XNOR2_X1 U19966 ( .A(n18103), .B(n17775), .ZN(n17776) );
  XNOR2_X1 U19967 ( .A(n24565), .B(n18531), .ZN(n18143) );
  XNOR2_X1 U19968 ( .A(n17776), .B(n18143), .ZN(n17778) );
  XNOR2_X1 U19969 ( .A(n18067), .B(n1768), .ZN(n17777) );
  XNOR2_X1 U19970 ( .A(n18435), .B(n18491), .ZN(n18238) );
  XNOR2_X1 U19971 ( .A(n18579), .B(n18121), .ZN(n17779) );
  XNOR2_X1 U19972 ( .A(n18238), .B(n17779), .ZN(n17782) );
  XNOR2_X1 U19973 ( .A(n18669), .B(n18582), .ZN(n18081) );
  XNOR2_X1 U19974 ( .A(n18665), .B(n1801), .ZN(n17780) );
  XNOR2_X1 U19975 ( .A(n18081), .B(n17780), .ZN(n17781) );
  INV_X1 U19977 ( .A(n19097), .ZN(n18724) );
  XNOR2_X1 U19978 ( .A(n18276), .B(n18549), .ZN(n17783) );
  XNOR2_X1 U19979 ( .A(n18200), .B(n18198), .ZN(n18550) );
  XNOR2_X1 U19980 ( .A(n17783), .B(n18550), .ZN(n17787) );
  XNOR2_X1 U19981 ( .A(n18473), .B(n2039), .ZN(n17784) );
  XNOR2_X1 U19982 ( .A(n17785), .B(n17784), .ZN(n17786) );
  INV_X1 U19983 ( .A(n19370), .ZN(n19364) );
  XNOR2_X1 U19987 ( .A(n17791), .B(n18157), .ZN(n18569) );
  XNOR2_X1 U19988 ( .A(n17792), .B(n18569), .ZN(n17793) );
  NAND3_X1 U19989 ( .A1(n19222), .A2(n19364), .A3(n19371), .ZN(n17802) );
  XNOR2_X1 U19990 ( .A(n18559), .B(n18308), .ZN(n17796) );
  XNOR2_X1 U19991 ( .A(n18310), .B(n17880), .ZN(n17795) );
  XNOR2_X1 U19992 ( .A(n17796), .B(n17795), .ZN(n17800) );
  XNOR2_X1 U19993 ( .A(n25411), .B(n25194), .ZN(n17798) );
  XNOR2_X1 U19994 ( .A(n17798), .B(n17797), .ZN(n17799) );
  XNOR2_X1 U19996 ( .A(n18675), .B(n451), .ZN(n17805) );
  XNOR2_X1 U19998 ( .A(n17807), .B(n17806), .ZN(n17808) );
  XNOR2_X1 U19999 ( .A(n17808), .B(n18294), .ZN(n18503) );
  XNOR2_X1 U20001 ( .A(n18512), .B(n2903), .ZN(n17810) );
  XNOR2_X1 U20002 ( .A(n17810), .B(n18370), .ZN(n17813) );
  XNOR2_X1 U20003 ( .A(n17811), .B(n18172), .ZN(n17812) );
  NAND2_X1 U20004 ( .A1(n19460), .A2(n19457), .ZN(n17887) );
  XNOR2_X1 U20005 ( .A(n17816), .B(n18446), .ZN(n17818) );
  XNOR2_X1 U20006 ( .A(n18350), .B(n17817), .ZN(n18253) );
  XNOR2_X1 U20007 ( .A(n18253), .B(n17818), .ZN(n17823) );
  XNOR2_X1 U20008 ( .A(n18523), .B(n18096), .ZN(n17821) );
  XNOR2_X1 U20009 ( .A(n17821), .B(n17820), .ZN(n17822) );
  XNOR2_X1 U20010 ( .A(n17823), .B(n17822), .ZN(n19456) );
  INV_X1 U20011 ( .A(n18430), .ZN(n17826) );
  XNOR2_X1 U20012 ( .A(n18275), .B(n887), .ZN(n17825) );
  XNOR2_X1 U20013 ( .A(n17826), .B(n17825), .ZN(n17830) );
  INV_X1 U20014 ( .A(n18692), .ZN(n17828) );
  XNOR2_X1 U20015 ( .A(n17828), .B(n17827), .ZN(n17829) );
  INV_X1 U20016 ( .A(n19457), .ZN(n19028) );
  NAND2_X1 U20017 ( .A1(n18976), .A2(n19028), .ZN(n17831) );
  NAND3_X1 U20018 ( .A1(n17887), .A2(n19456), .A3(n17831), .ZN(n17848) );
  XNOR2_X1 U20019 ( .A(n17832), .B(n18658), .ZN(n17834) );
  XNOR2_X1 U20020 ( .A(n17833), .B(n17834), .ZN(n17838) );
  XNOR2_X1 U20021 ( .A(n18104), .B(n18483), .ZN(n17836) );
  XNOR2_X1 U20023 ( .A(n17836), .B(n17835), .ZN(n17837) );
  XNOR2_X1 U20024 ( .A(n17837), .B(n17838), .ZN(n17845) );
  INV_X1 U20025 ( .A(n17845), .ZN(n18979) );
  XNOR2_X1 U20026 ( .A(n17839), .B(n18122), .ZN(n17841) );
  XNOR2_X1 U20027 ( .A(n17841), .B(n18537), .ZN(n17844) );
  XNOR2_X1 U20028 ( .A(n18038), .B(n18489), .ZN(n18259) );
  XNOR2_X1 U20029 ( .A(n18539), .B(n20825), .ZN(n17842) );
  XNOR2_X1 U20030 ( .A(n18259), .B(n17842), .ZN(n17843) );
  XNOR2_X1 U20031 ( .A(n17843), .B(n17844), .ZN(n18977) );
  INV_X1 U20032 ( .A(n18977), .ZN(n19032) );
  NAND3_X1 U20033 ( .A1(n24172), .A2(n18979), .A3(n19032), .ZN(n17847) );
  NAND3_X1 U20034 ( .A1(n19460), .A2(n19457), .A3(n19464), .ZN(n17846) );
  NOR2_X1 U20035 ( .A1(n19887), .A2(n25388), .ZN(n17849) );
  XNOR2_X1 U20036 ( .A(n18190), .B(n681), .ZN(n17850) );
  INV_X1 U20037 ( .A(n18484), .ZN(n17853) );
  XNOR2_X1 U20038 ( .A(n18103), .B(n17853), .ZN(n17854) );
  XNOR2_X1 U20039 ( .A(n17854), .B(n18232), .ZN(n17858) );
  XNOR2_X1 U20040 ( .A(n24568), .B(n18335), .ZN(n17856) );
  XNOR2_X1 U20041 ( .A(n18270), .B(n2042), .ZN(n17855) );
  XNOR2_X1 U20042 ( .A(n17856), .B(n17855), .ZN(n17857) );
  XNOR2_X1 U20043 ( .A(n18004), .B(n17859), .ZN(n17861) );
  XNOR2_X1 U20044 ( .A(n18198), .B(n2882), .ZN(n17860) );
  XNOR2_X1 U20045 ( .A(n17861), .B(n17860), .ZN(n17865) );
  XNOR2_X1 U20046 ( .A(n17862), .B(n17863), .ZN(n18645) );
  XNOR2_X1 U20047 ( .A(n18645), .B(n18219), .ZN(n17864) );
  XNOR2_X1 U20048 ( .A(n17864), .B(n17865), .ZN(n19321) );
  MUX2_X1 U20049 ( .A(n18959), .B(n19470), .S(n19321), .Z(n17886) );
  XNOR2_X1 U20050 ( .A(n18251), .B(n18448), .ZN(n17868) );
  XNOR2_X1 U20051 ( .A(n18418), .B(Key[172]), .ZN(n17866) );
  XNOR2_X1 U20054 ( .A(n18447), .B(n18214), .ZN(n17869) );
  XNOR2_X1 U20055 ( .A(n18098), .B(n17869), .ZN(n17870) );
  XNOR2_X1 U20056 ( .A(n17873), .B(n18121), .ZN(n18580) );
  XNOR2_X1 U20057 ( .A(n18580), .B(n18238), .ZN(n17879) );
  XNOR2_X1 U20058 ( .A(n25000), .B(n4942), .ZN(n17877) );
  XNOR2_X1 U20059 ( .A(n18262), .B(n187), .ZN(n17876) );
  XNOR2_X1 U20060 ( .A(n17877), .B(n17876), .ZN(n17878) );
  XNOR2_X1 U20061 ( .A(n17881), .B(n17880), .ZN(n18560) );
  XNOR2_X1 U20062 ( .A(n18130), .B(n17882), .ZN(n17885) );
  XNOR2_X1 U20063 ( .A(n18515), .B(n25194), .ZN(n18247) );
  XNOR2_X1 U20064 ( .A(n17883), .B(n18247), .ZN(n17884) );
  INV_X1 U20065 ( .A(n19466), .ZN(n18960) );
  INV_X1 U20066 ( .A(n19460), .ZN(n18739) );
  AND2_X1 U20067 ( .A1(n17888), .A2(n17887), .ZN(n17893) );
  NAND2_X1 U20068 ( .A1(n19456), .A2(n18977), .ZN(n19465) );
  NAND2_X1 U20071 ( .A1(n17890), .A2(n19464), .ZN(n17891) );
  OAI21_X2 U20072 ( .B1(n17893), .B2(n17892), .A(n17891), .ZN(n19896) );
  NAND2_X1 U20073 ( .A1(n19697), .A2(n19896), .ZN(n17947) );
  INV_X1 U20074 ( .A(n17947), .ZN(n17950) );
  NOR2_X1 U20075 ( .A1(n18735), .A2(n19477), .ZN(n19480) );
  XNOR2_X1 U20076 ( .A(n17897), .B(n17898), .ZN(n17904) );
  XNOR2_X1 U20077 ( .A(n17900), .B(n17899), .ZN(n17902) );
  XNOR2_X1 U20078 ( .A(n18149), .B(n62), .ZN(n17901) );
  XNOR2_X1 U20079 ( .A(n17902), .B(n17901), .ZN(n17903) );
  XNOR2_X1 U20080 ( .A(n18124), .B(n17905), .ZN(n18623) );
  XNOR2_X1 U20081 ( .A(n18623), .B(n17906), .ZN(n17910) );
  XNOR2_X1 U20082 ( .A(n17907), .B(n673), .ZN(n17908) );
  XNOR2_X1 U20083 ( .A(n17908), .B(n18081), .ZN(n17909) );
  XNOR2_X1 U20084 ( .A(n17909), .B(n17910), .ZN(n19502) );
  XNOR2_X1 U20085 ( .A(n17912), .B(n17911), .ZN(n17917) );
  XNOR2_X1 U20086 ( .A(n24433), .B(n2240), .ZN(n17914) );
  XNOR2_X1 U20087 ( .A(n17915), .B(n17914), .ZN(n17916) );
  INV_X1 U20088 ( .A(n18719), .ZN(n19335) );
  XNOR2_X1 U20089 ( .A(n25006), .B(n17918), .ZN(n17923) );
  XNOR2_X1 U20090 ( .A(n24431), .B(n18331), .ZN(n17921) );
  XNOR2_X1 U20091 ( .A(n18270), .B(n881), .ZN(n17920) );
  XNOR2_X1 U20092 ( .A(n17921), .B(n17920), .ZN(n17922) );
  NOR2_X1 U20093 ( .A1(n18986), .A2(n17924), .ZN(n17940) );
  INV_X1 U20094 ( .A(n18559), .ZN(n17925) );
  XNOR2_X1 U20095 ( .A(n17926), .B(n17925), .ZN(n18058) );
  INV_X1 U20096 ( .A(n18058), .ZN(n17930) );
  XNOR2_X1 U20098 ( .A(n17927), .B(n18374), .ZN(n17928) );
  XNOR2_X1 U20099 ( .A(n17928), .B(n18309), .ZN(n17929) );
  NAND2_X1 U20101 ( .A1(n19335), .A2(n19499), .ZN(n18987) );
  XNOR2_X1 U20102 ( .A(n18476), .B(n17931), .ZN(n18644) );
  XNOR2_X1 U20103 ( .A(n17932), .B(n18644), .ZN(n17937) );
  XNOR2_X1 U20104 ( .A(n24536), .B(n18693), .ZN(n17935) );
  XNOR2_X1 U20105 ( .A(n18200), .B(n860), .ZN(n17934) );
  XNOR2_X1 U20106 ( .A(n17935), .B(n17934), .ZN(n17936) );
  XNOR2_X1 U20107 ( .A(n17937), .B(n17936), .ZN(n19498) );
  NAND2_X1 U20108 ( .A1(n19497), .A2(n25459), .ZN(n17938) );
  OAI21_X1 U20109 ( .B1(n24370), .B2(n19896), .A(n21033), .ZN(n17949) );
  NAND3_X1 U20110 ( .A1(n18970), .A2(n19297), .A3(n18967), .ZN(n17941) );
  MUX2_X1 U20111 ( .A(n17947), .B(n17946), .S(n21038), .Z(n17948) );
  XNOR2_X1 U20112 ( .A(n17951), .B(n17952), .ZN(n18712) );
  XNOR2_X1 U20113 ( .A(n17953), .B(n18404), .ZN(n17957) );
  XNOR2_X1 U20114 ( .A(n18233), .B(n18658), .ZN(n17955) );
  XNOR2_X1 U20115 ( .A(n18530), .B(n21423), .ZN(n17954) );
  XNOR2_X1 U20116 ( .A(n17955), .B(n17954), .ZN(n17956) );
  XNOR2_X1 U20117 ( .A(n18004), .B(n17958), .ZN(n17962) );
  INV_X1 U20118 ( .A(n17959), .ZN(n18548) );
  XNOR2_X1 U20119 ( .A(n18548), .B(n17960), .ZN(n17961) );
  XNOR2_X1 U20120 ( .A(n17962), .B(n17961), .ZN(n17965) );
  XNOR2_X1 U20121 ( .A(n18475), .B(n17963), .ZN(n17964) );
  XNOR2_X1 U20122 ( .A(n17964), .B(n17965), .ZN(n18876) );
  XNOR2_X1 U20123 ( .A(n18465), .B(n23983), .ZN(n17966) );
  XNOR2_X1 U20124 ( .A(n17966), .B(n18562), .ZN(n17968) );
  XNOR2_X1 U20125 ( .A(n17968), .B(n17967), .ZN(n17973) );
  XNOR2_X1 U20126 ( .A(n18042), .B(n17969), .ZN(n17971) );
  XNOR2_X1 U20127 ( .A(n17970), .B(n17971), .ZN(n17972) );
  XNOR2_X1 U20128 ( .A(n17974), .B(n18422), .ZN(n17975) );
  INV_X1 U20129 ( .A(n19092), .ZN(n18819) );
  AOI21_X1 U20130 ( .B1(n18876), .B2(n19094), .A(n18819), .ZN(n17980) );
  XNOR2_X1 U20131 ( .A(n18227), .B(n17663), .ZN(n17976) );
  XNOR2_X1 U20132 ( .A(n17976), .B(n24371), .ZN(n17979) );
  XNOR2_X1 U20133 ( .A(n18637), .B(n2190), .ZN(n17977) );
  XNOR2_X1 U20134 ( .A(n17977), .B(n18415), .ZN(n17978) );
  XNOR2_X1 U20135 ( .A(n17979), .B(n17978), .ZN(n19382) );
  XNOR2_X1 U20136 ( .A(n17981), .B(n17982), .ZN(n17985) );
  XNOR2_X1 U20137 ( .A(n4942), .B(n3084), .ZN(n17983) );
  XNOR2_X1 U20138 ( .A(n18259), .B(n17983), .ZN(n17984) );
  NOR3_X1 U20139 ( .A1(n24335), .A2(n19380), .A3(n19377), .ZN(n17986) );
  INV_X1 U20140 ( .A(n17987), .ZN(n17988) );
  XNOR2_X1 U20141 ( .A(n17988), .B(n18348), .ZN(n17992) );
  XNOR2_X1 U20142 ( .A(n18325), .B(n765), .ZN(n17989) );
  XNOR2_X1 U20143 ( .A(n17989), .B(n17990), .ZN(n17991) );
  XNOR2_X1 U20144 ( .A(n17993), .B(n18610), .ZN(n17995) );
  XNOR2_X1 U20145 ( .A(n17995), .B(n17994), .ZN(n17999) );
  XNOR2_X1 U20146 ( .A(n24431), .B(n17582), .ZN(n17997) );
  XNOR2_X1 U20147 ( .A(n18532), .B(n2726), .ZN(n17996) );
  XNOR2_X1 U20148 ( .A(n17997), .B(n17996), .ZN(n17998) );
  XNOR2_X1 U20150 ( .A(n18466), .B(n23476), .ZN(n18000) );
  XNOR2_X1 U20151 ( .A(n18000), .B(n18370), .ZN(n18001) );
  XNOR2_X1 U20152 ( .A(n18285), .B(n18628), .ZN(n18057) );
  XNOR2_X1 U20153 ( .A(n18057), .B(n18001), .ZN(n18003) );
  XNOR2_X1 U20154 ( .A(n18003), .B(n18002), .ZN(n18817) );
  XNOR2_X1 U20155 ( .A(n18196), .B(n18005), .ZN(n18008) );
  XNOR2_X1 U20156 ( .A(n18060), .B(n18006), .ZN(n18281) );
  XNOR2_X1 U20157 ( .A(n18363), .B(n18281), .ZN(n18007) );
  INV_X1 U20158 ( .A(n19360), .ZN(n18009) );
  INV_X1 U20159 ( .A(n1745), .ZN(n23508) );
  XNOR2_X1 U20160 ( .A(n18261), .B(n23508), .ZN(n18011) );
  XNOR2_X1 U20161 ( .A(n4942), .B(n18539), .ZN(n18010) );
  XNOR2_X1 U20162 ( .A(n18011), .B(n18010), .ZN(n18012) );
  INV_X1 U20163 ( .A(n18295), .ZN(n18014) );
  XNOR2_X1 U20164 ( .A(n18014), .B(n18294), .ZN(n18016) );
  XNOR2_X1 U20165 ( .A(n18456), .B(n2747), .ZN(n18015) );
  XNOR2_X1 U20166 ( .A(n18016), .B(n18015), .ZN(n18020) );
  XNOR2_X1 U20167 ( .A(n18018), .B(n18017), .ZN(n18192) );
  XNOR2_X1 U20168 ( .A(n18192), .B(n18390), .ZN(n18019) );
  INV_X1 U20170 ( .A(n19878), .ZN(n20329) );
  NOR2_X1 U20171 ( .A1(n20554), .A2(n20329), .ZN(n18136) );
  XNOR2_X1 U20172 ( .A(n18022), .B(n18023), .ZN(n18025) );
  XNOR2_X1 U20173 ( .A(n18024), .B(n18025), .ZN(n18030) );
  INV_X1 U20174 ( .A(n18326), .ZN(n18026) );
  XNOR2_X1 U20175 ( .A(n18026), .B(n3115), .ZN(n18027) );
  XNOR2_X1 U20176 ( .A(n18028), .B(n18027), .ZN(n18029) );
  INV_X1 U20177 ( .A(n19595), .ZN(n18037) );
  INV_X1 U20178 ( .A(n18360), .ZN(n18031) );
  XNOR2_X1 U20179 ( .A(n18331), .B(n18658), .ZN(n18587) );
  XNOR2_X1 U20180 ( .A(n18031), .B(n18587), .ZN(n18036) );
  XNOR2_X1 U20181 ( .A(n18032), .B(n18530), .ZN(n18034) );
  XNOR2_X1 U20182 ( .A(n18356), .B(n2805), .ZN(n18033) );
  XNOR2_X1 U20183 ( .A(n18034), .B(n18033), .ZN(n18035) );
  AND2_X1 U20184 ( .A1(n18037), .A2(n19598), .ZN(n19257) );
  XNOR2_X1 U20185 ( .A(n18038), .B(n18240), .ZN(n18584) );
  XNOR2_X1 U20186 ( .A(n18039), .B(n18584), .ZN(n18041) );
  XNOR2_X1 U20187 ( .A(n18042), .B(n3183), .ZN(n18043) );
  XNOR2_X1 U20189 ( .A(n18045), .B(n18429), .ZN(n18047) );
  XNOR2_X1 U20190 ( .A(n18548), .B(n18060), .ZN(n18046) );
  XNOR2_X1 U20191 ( .A(n18047), .B(n18046), .ZN(n18048) );
  XNOR2_X1 U20192 ( .A(n18295), .B(n2847), .ZN(n18050) );
  XNOR2_X1 U20193 ( .A(n18052), .B(n18051), .ZN(n18830) );
  NAND2_X1 U20195 ( .A1(n19597), .A2(n24079), .ZN(n18053) );
  OAI21_X2 U20196 ( .B1(n18054), .B2(n18055), .A(n18053), .ZN(n20330) );
  INV_X1 U20197 ( .A(n20330), .ZN(n20556) );
  XNOR2_X1 U20198 ( .A(n18172), .B(n2735), .ZN(n18056) );
  XNOR2_X1 U20199 ( .A(n18197), .B(n18277), .ZN(n18062) );
  XNOR2_X1 U20200 ( .A(n18060), .B(n18693), .ZN(n18061) );
  XNOR2_X1 U20201 ( .A(n18062), .B(n18061), .ZN(n18066) );
  XNOR2_X1 U20202 ( .A(n18552), .B(n18200), .ZN(n18064) );
  XNOR2_X1 U20203 ( .A(n18432), .B(n21169), .ZN(n18063) );
  XNOR2_X1 U20204 ( .A(n18064), .B(n18063), .ZN(n18065) );
  XNOR2_X1 U20205 ( .A(n18067), .B(n18610), .ZN(n18588) );
  XNOR2_X1 U20206 ( .A(n18104), .B(n18660), .ZN(n18068) );
  XNOR2_X1 U20207 ( .A(n2052), .B(n18068), .ZN(n18072) );
  XNOR2_X1 U20208 ( .A(n24568), .B(n18356), .ZN(n18070) );
  XNOR2_X1 U20209 ( .A(n18270), .B(n2222), .ZN(n18069) );
  XNOR2_X1 U20210 ( .A(n18070), .B(n18069), .ZN(n18071) );
  AND2_X1 U20211 ( .A1(n24483), .A2(n19080), .ZN(n18093) );
  XNOR2_X1 U20212 ( .A(n18073), .B(n18074), .ZN(n18574) );
  INV_X1 U20213 ( .A(n18574), .ZN(n18207) );
  XNOR2_X1 U20214 ( .A(n18251), .B(n18254), .ZN(n18075) );
  XNOR2_X1 U20215 ( .A(n18207), .B(n18075), .ZN(n18079) );
  XNOR2_X1 U20216 ( .A(n18418), .B(n16), .ZN(n18077) );
  XNOR2_X1 U20217 ( .A(n18077), .B(n18076), .ZN(n18078) );
  XNOR2_X1 U20218 ( .A(n18079), .B(n18078), .ZN(n19078) );
  INV_X1 U20219 ( .A(n19078), .ZN(n19592) );
  INV_X1 U20220 ( .A(n19589), .ZN(n18092) );
  INV_X1 U20221 ( .A(n18620), .ZN(n18082) );
  XNOR2_X1 U20222 ( .A(n18082), .B(n18081), .ZN(n18084) );
  XNOR2_X1 U20223 ( .A(n18261), .B(n677), .ZN(n18083) );
  XNOR2_X1 U20224 ( .A(n24488), .B(n2991), .ZN(n18085) );
  AND2_X1 U20226 ( .A1(n19591), .A2(n19077), .ZN(n18806) );
  XNOR2_X1 U20227 ( .A(n18423), .B(n173), .ZN(n18094) );
  XNOR2_X1 U20228 ( .A(n18094), .B(n18602), .ZN(n18095) );
  XNOR2_X1 U20229 ( .A(n18095), .B(n18323), .ZN(n18100) );
  XNOR2_X1 U20230 ( .A(n18096), .B(n18214), .ZN(n18097) );
  XOR2_X1 U20231 ( .A(n18098), .B(n18097), .Z(n18099) );
  XNOR2_X1 U20232 ( .A(n18611), .B(n18407), .ZN(n18482) );
  XNOR2_X1 U20233 ( .A(n18101), .B(n18482), .ZN(n18108) );
  XNOR2_X1 U20234 ( .A(n18103), .B(n18102), .ZN(n18591) );
  INV_X1 U20235 ( .A(n18591), .ZN(n18106) );
  XNOR2_X1 U20236 ( .A(n18104), .B(n3125), .ZN(n18105) );
  XNOR2_X1 U20237 ( .A(n18105), .B(n18106), .ZN(n18107) );
  XNOR2_X1 U20238 ( .A(n18197), .B(n18365), .ZN(n18110) );
  XNOR2_X1 U20239 ( .A(n18110), .B(n18109), .ZN(n18113) );
  INV_X1 U20240 ( .A(n19392), .ZN(n23693) );
  XNOR2_X1 U20241 ( .A(n17476), .B(n23693), .ZN(n18111) );
  XNOR2_X1 U20242 ( .A(n18342), .B(n18111), .ZN(n18112) );
  XNOR2_X1 U20243 ( .A(n18112), .B(n18113), .ZN(n19607) );
  XNOR2_X1 U20247 ( .A(n18116), .B(n18190), .ZN(n18568) );
  XNOR2_X2 U20250 ( .A(n18118), .B(n18119), .ZN(n19233) );
  AOI21_X1 U20251 ( .B1(n19607), .B2(n19112), .A(n19233), .ZN(n18120) );
  XNOR2_X1 U20252 ( .A(n18122), .B(n18121), .ZN(n18184) );
  XNOR2_X1 U20253 ( .A(n18317), .B(n18125), .ZN(n18126) );
  XNOR2_X1 U20254 ( .A(n18127), .B(n18126), .ZN(n19237) );
  XNOR2_X1 U20255 ( .A(n18310), .B(n3089), .ZN(n18132) );
  XNOR2_X1 U20256 ( .A(n18172), .B(n18312), .ZN(n18131) );
  XNOR2_X1 U20257 ( .A(n18132), .B(n18131), .ZN(n18133) );
  AOI21_X1 U20258 ( .B1(n19610), .B2(n24310), .A(n1404), .ZN(n18134) );
  INV_X1 U20259 ( .A(n20328), .ZN(n20089) );
  XNOR2_X1 U20260 ( .A(n18258), .B(n18579), .ZN(n18137) );
  XNOR2_X1 U20261 ( .A(n18538), .B(n18137), .ZN(n18141) );
  INV_X1 U20262 ( .A(n18237), .ZN(n18139) );
  XNOR2_X1 U20263 ( .A(n18621), .B(n2211), .ZN(n18138) );
  XNOR2_X1 U20264 ( .A(n18139), .B(n18138), .ZN(n18140) );
  INV_X1 U20265 ( .A(n18142), .ZN(n18144) );
  XNOR2_X1 U20266 ( .A(n18144), .B(n18143), .ZN(n18145) );
  XNOR2_X1 U20267 ( .A(n18447), .B(n18700), .ZN(n18522) );
  INV_X1 U20268 ( .A(n18522), .ZN(n18148) );
  XNOR2_X1 U20269 ( .A(n18146), .B(n18446), .ZN(n18147) );
  XNOR2_X1 U20270 ( .A(n18149), .B(n18599), .ZN(n18151) );
  XNOR2_X1 U20271 ( .A(n18605), .B(n2126), .ZN(n18150) );
  XNOR2_X1 U20272 ( .A(n18151), .B(n18150), .ZN(n18152) );
  XNOR2_X1 U20273 ( .A(n18248), .B(n18627), .ZN(n18156) );
  XNOR2_X1 U20274 ( .A(n364), .B(n18685), .ZN(n18154) );
  XNOR2_X1 U20275 ( .A(n18154), .B(n18153), .ZN(n18155) );
  XNOR2_X1 U20276 ( .A(n18155), .B(n18156), .ZN(n19579) );
  INV_X1 U20277 ( .A(n19579), .ZN(n19198) );
  XNOR2_X1 U20278 ( .A(n18674), .B(n1869), .ZN(n18158) );
  XNOR2_X1 U20279 ( .A(n18159), .B(n18158), .ZN(n18162) );
  XNOR2_X1 U20280 ( .A(n18160), .B(n18226), .ZN(n18161) );
  XNOR2_X1 U20281 ( .A(n18161), .B(n18162), .ZN(n19199) );
  NAND3_X1 U20282 ( .A1(n3412), .A2(n24481), .A3(n19198), .ZN(n18168) );
  XNOR2_X1 U20283 ( .A(n18473), .B(n18694), .ZN(n18509) );
  XNOR2_X1 U20284 ( .A(n18549), .B(n21742), .ZN(n18163) );
  XNOR2_X1 U20285 ( .A(n18163), .B(n18648), .ZN(n18164) );
  XNOR2_X1 U20286 ( .A(n18164), .B(n18165), .ZN(n18809) );
  INV_X1 U20287 ( .A(n18809), .ZN(n19580) );
  XNOR2_X1 U20289 ( .A(n18465), .B(n2100), .ZN(n18169) );
  XNOR2_X1 U20290 ( .A(n18169), .B(n18559), .ZN(n18170) );
  XNOR2_X1 U20291 ( .A(n18170), .B(n18171), .ZN(n18175) );
  XNOR2_X1 U20292 ( .A(n18173), .B(n18513), .ZN(n18174) );
  XNOR2_X1 U20294 ( .A(n18483), .B(n2826), .ZN(n18177) );
  XNOR2_X1 U20295 ( .A(n18178), .B(n18177), .ZN(n18179) );
  XNOR2_X1 U20296 ( .A(n18582), .B(n18382), .ZN(n18182) );
  XNOR2_X1 U20297 ( .A(n18489), .B(n1364), .ZN(n18181) );
  XNOR2_X1 U20298 ( .A(n18182), .B(n18181), .ZN(n18186) );
  XNOR2_X1 U20299 ( .A(n18183), .B(n18184), .ZN(n18185) );
  XNOR2_X1 U20300 ( .A(n18185), .B(n18186), .ZN(n19518) );
  XNOR2_X1 U20301 ( .A(n18187), .B(n18188), .ZN(n18386) );
  XNOR2_X1 U20302 ( .A(n18386), .B(n18189), .ZN(n18194) );
  XNOR2_X1 U20303 ( .A(n18190), .B(n2782), .ZN(n18191) );
  XNOR2_X1 U20304 ( .A(n18192), .B(n18191), .ZN(n18193) );
  OAI21_X1 U20305 ( .B1(n19518), .B2(n19522), .A(n19279), .ZN(n18205) );
  XNOR2_X1 U20306 ( .A(n25077), .B(n18275), .ZN(n18364) );
  XNOR2_X1 U20307 ( .A(n18364), .B(n18196), .ZN(n18204) );
  INV_X1 U20308 ( .A(n18197), .ZN(n18199) );
  XNOR2_X1 U20309 ( .A(n18199), .B(n18198), .ZN(n18202) );
  XNOR2_X1 U20310 ( .A(n18200), .B(n876), .ZN(n18201) );
  XNOR2_X1 U20311 ( .A(n18202), .B(n18201), .ZN(n18203) );
  XNOR2_X1 U20312 ( .A(n18203), .B(n18204), .ZN(n19284) );
  MUX2_X1 U20313 ( .A(n18206), .B(n18205), .S(n19284), .Z(n19723) );
  XNOR2_X1 U20314 ( .A(n18207), .B(n18704), .ZN(n18211) );
  XNOR2_X1 U20315 ( .A(n18350), .B(n1789), .ZN(n18209) );
  INV_X1 U20316 ( .A(n19720), .ZN(n18212) );
  XNOR2_X1 U20318 ( .A(n18447), .B(n18446), .ZN(n18213) );
  XNOR2_X1 U20319 ( .A(n18213), .B(n18607), .ZN(n18217) );
  XNOR2_X1 U20320 ( .A(n18451), .B(n886), .ZN(n18215) );
  XNOR2_X1 U20321 ( .A(n18576), .B(n18215), .ZN(n18216) );
  INV_X1 U20322 ( .A(n19184), .ZN(n19552) );
  XNOR2_X1 U20323 ( .A(n18219), .B(n18218), .ZN(n18224) );
  XNOR2_X1 U20324 ( .A(n18432), .B(n18220), .ZN(n18222) );
  XNOR2_X1 U20325 ( .A(n24383), .B(n1804), .ZN(n18221) );
  XNOR2_X1 U20326 ( .A(n18222), .B(n18221), .ZN(n18223) );
  XNOR2_X1 U20327 ( .A(n18226), .B(n18225), .ZN(n18231) );
  XNOR2_X1 U20328 ( .A(n18227), .B(n24416), .ZN(n18229) );
  XNOR2_X1 U20329 ( .A(n18229), .B(n18228), .ZN(n18230) );
  XNOR2_X1 U20330 ( .A(n18481), .B(n18232), .ZN(n18236) );
  XNOR2_X1 U20331 ( .A(n18331), .B(n1792), .ZN(n18234) );
  XNOR2_X1 U20332 ( .A(n18612), .B(n18234), .ZN(n18235) );
  XNOR2_X1 U20333 ( .A(n18237), .B(n18238), .ZN(n18244) );
  XNOR2_X1 U20334 ( .A(n18240), .B(n18239), .ZN(n18242) );
  XNOR2_X1 U20335 ( .A(n18242), .B(n18241), .ZN(n18243) );
  XNOR2_X1 U20336 ( .A(n18244), .B(n18243), .ZN(n19402) );
  NAND2_X1 U20337 ( .A1(n19184), .A2(n19402), .ZN(n19719) );
  XNOR2_X1 U20338 ( .A(n18557), .B(n21944), .ZN(n18245) );
  XNOR2_X1 U20339 ( .A(n18246), .B(n18245), .ZN(n18250) );
  XNOR2_X1 U20340 ( .A(n18247), .B(n18248), .ZN(n18249) );
  INV_X1 U20341 ( .A(n20560), .ZN(n20023) );
  XNOR2_X1 U20342 ( .A(n18252), .B(n18251), .ZN(n18703) );
  XNOR2_X1 U20343 ( .A(n18703), .B(n18253), .ZN(n18257) );
  XNOR2_X1 U20344 ( .A(n18254), .B(n2050), .ZN(n18255) );
  XNOR2_X1 U20345 ( .A(n18523), .B(n18605), .ZN(n18425) );
  XNOR2_X1 U20346 ( .A(n18425), .B(n18255), .ZN(n18256) );
  XNOR2_X1 U20347 ( .A(n18258), .B(n18665), .ZN(n18260) );
  XNOR2_X1 U20348 ( .A(n18259), .B(n18260), .ZN(n18266) );
  XNOR2_X1 U20349 ( .A(n18261), .B(n18539), .ZN(n18264) );
  XNOR2_X1 U20350 ( .A(n18262), .B(n3133), .ZN(n18263) );
  XNOR2_X1 U20351 ( .A(n18264), .B(n18263), .ZN(n18265) );
  XNOR2_X1 U20352 ( .A(n18266), .B(n18265), .ZN(n19277) );
  XNOR2_X1 U20353 ( .A(n18268), .B(n18267), .ZN(n18274) );
  XNOR2_X1 U20354 ( .A(n18269), .B(n18483), .ZN(n18272) );
  XNOR2_X1 U20355 ( .A(n18270), .B(n1815), .ZN(n18271) );
  XNOR2_X1 U20356 ( .A(n18272), .B(n18271), .ZN(n18273) );
  OAI21_X1 U20357 ( .B1(n5573), .B2(n1334), .A(n19126), .ZN(n18299) );
  XNOR2_X1 U20358 ( .A(n18548), .B(n18275), .ZN(n18279) );
  XNOR2_X1 U20359 ( .A(n18276), .B(n18277), .ZN(n18691) );
  INV_X1 U20360 ( .A(n18691), .ZN(n18278) );
  XNOR2_X1 U20361 ( .A(n18279), .B(n18278), .ZN(n18282) );
  XNOR2_X1 U20362 ( .A(n18431), .B(n21662), .ZN(n18280) );
  XNOR2_X1 U20363 ( .A(n18287), .B(n18288), .ZN(n18772) );
  XNOR2_X1 U20364 ( .A(n18290), .B(n18289), .ZN(n18680) );
  INV_X1 U20365 ( .A(n18680), .ZN(n18292) );
  XNOR2_X1 U20366 ( .A(n18292), .B(n24371), .ZN(n18298) );
  XNOR2_X1 U20367 ( .A(n18293), .B(n18294), .ZN(n18412) );
  XNOR2_X1 U20368 ( .A(n18295), .B(n2881), .ZN(n18296) );
  XNOR2_X1 U20369 ( .A(n18412), .B(n18296), .ZN(n18297) );
  XNOR2_X1 U20370 ( .A(n18298), .B(n18297), .ZN(n18902) );
  XNOR2_X1 U20371 ( .A(n25380), .B(n21703), .ZN(n18302) );
  XNOR2_X1 U20372 ( .A(n24416), .B(n18302), .ZN(n18304) );
  XNOR2_X1 U20373 ( .A(n18303), .B(n18304), .ZN(n18307) );
  XNOR2_X1 U20374 ( .A(n18305), .B(n18677), .ZN(n18306) );
  XNOR2_X1 U20375 ( .A(n18308), .B(n18513), .ZN(n18684) );
  XNOR2_X1 U20376 ( .A(n18309), .B(n18684), .ZN(n18316) );
  XNOR2_X1 U20377 ( .A(n18310), .B(n5131), .ZN(n18314) );
  XNOR2_X1 U20378 ( .A(n18312), .B(n18311), .ZN(n18313) );
  XNOR2_X1 U20379 ( .A(n18313), .B(n18314), .ZN(n18315) );
  NOR2_X1 U20380 ( .A1(n19191), .A2(n19565), .ZN(n18340) );
  XNOR2_X1 U20381 ( .A(n18318), .B(n18317), .ZN(n18322) );
  XNOR2_X1 U20382 ( .A(n18540), .B(n18621), .ZN(n18320) );
  XNOR2_X1 U20383 ( .A(n18669), .B(n2761), .ZN(n18319) );
  XNOR2_X1 U20384 ( .A(n18320), .B(n18319), .ZN(n18321) );
  XNOR2_X1 U20385 ( .A(n18324), .B(n18323), .ZN(n18330) );
  XNOR2_X1 U20386 ( .A(n18325), .B(n18326), .ZN(n18328) );
  XNOR2_X1 U20387 ( .A(n18599), .B(n1920), .ZN(n18327) );
  XNOR2_X1 U20388 ( .A(n18327), .B(n18328), .ZN(n18329) );
  XNOR2_X1 U20389 ( .A(n24565), .B(n18331), .ZN(n18332) );
  XNOR2_X1 U20390 ( .A(n25006), .B(n18332), .ZN(n18339) );
  XNOR2_X1 U20391 ( .A(n18334), .B(n17582), .ZN(n18337) );
  XNOR2_X1 U20392 ( .A(n18335), .B(n1810), .ZN(n18336) );
  XNOR2_X1 U20393 ( .A(n18337), .B(n18336), .ZN(n18338) );
  XNOR2_X1 U20394 ( .A(n18693), .B(n18341), .ZN(n18343) );
  XNOR2_X1 U20395 ( .A(n18342), .B(n18343), .ZN(n18347) );
  INV_X1 U20396 ( .A(n3129), .ZN(n23825) );
  XNOR2_X1 U20397 ( .A(n18476), .B(n23825), .ZN(n18345) );
  XNOR2_X1 U20398 ( .A(n24384), .B(n18695), .ZN(n18344) );
  XNOR2_X1 U20399 ( .A(n18345), .B(n18344), .ZN(n18346) );
  XNOR2_X1 U20400 ( .A(n18347), .B(n18346), .ZN(n19273) );
  NOR2_X1 U20401 ( .A1(n19566), .A2(n19273), .ZN(n18395) );
  XNOR2_X1 U20403 ( .A(n18349), .B(n18348), .ZN(n18354) );
  XNOR2_X1 U20404 ( .A(n18423), .B(n18350), .ZN(n18453) );
  XNOR2_X1 U20405 ( .A(n18351), .B(n4233), .ZN(n18352) );
  XNOR2_X1 U20406 ( .A(n18453), .B(n18352), .ZN(n18353) );
  INV_X1 U20407 ( .A(n18407), .ZN(n18355) );
  XNOR2_X1 U20408 ( .A(n18355), .B(n18483), .ZN(n18358) );
  XNOR2_X1 U20409 ( .A(n18356), .B(n1776), .ZN(n18357) );
  XNOR2_X1 U20410 ( .A(n18358), .B(n18357), .ZN(n18362) );
  XNOR2_X1 U20411 ( .A(n18359), .B(n18360), .ZN(n18361) );
  XNOR2_X1 U20412 ( .A(n18364), .B(n18363), .ZN(n18369) );
  XNOR2_X1 U20413 ( .A(n18365), .B(n1891), .ZN(n18366) );
  XNOR2_X1 U20414 ( .A(n18367), .B(n18366), .ZN(n18368) );
  XNOR2_X1 U20415 ( .A(n18369), .B(n18368), .ZN(n19176) );
  INV_X1 U20416 ( .A(n19176), .ZN(n18777) );
  XNOR2_X1 U20417 ( .A(n18371), .B(n18370), .ZN(n18373) );
  XNOR2_X1 U20418 ( .A(n18372), .B(n18373), .ZN(n18379) );
  XNOR2_X1 U20419 ( .A(n18374), .B(n23679), .ZN(n18377) );
  XNOR2_X1 U20420 ( .A(n18465), .B(n18375), .ZN(n18376) );
  XNOR2_X1 U20421 ( .A(n18376), .B(n18377), .ZN(n18378) );
  XNOR2_X1 U20422 ( .A(n18380), .B(n18381), .ZN(n18384) );
  XNOR2_X1 U20423 ( .A(n18437), .B(n18382), .ZN(n18383) );
  XNOR2_X1 U20424 ( .A(n18387), .B(n18386), .ZN(n18392) );
  XNOR2_X1 U20425 ( .A(n18388), .B(n2989), .ZN(n18389) );
  XNOR2_X1 U20426 ( .A(n18390), .B(n18389), .ZN(n18391) );
  OAI21_X1 U20427 ( .B1(n25195), .B2(n19176), .A(n19428), .ZN(n18393) );
  NAND2_X1 U20428 ( .A1(n19183), .A2(n18393), .ZN(n18394) );
  NOR2_X1 U20429 ( .A1(n19730), .A2(n19729), .ZN(n18445) );
  XNOR2_X1 U20430 ( .A(n18397), .B(n25194), .ZN(n18398) );
  XNOR2_X1 U20431 ( .A(n18399), .B(n18398), .ZN(n18403) );
  XNOR2_X1 U20432 ( .A(n18512), .B(n2005), .ZN(n18400) );
  XNOR2_X1 U20433 ( .A(n18401), .B(n18400), .ZN(n18402) );
  XNOR2_X1 U20434 ( .A(n18405), .B(n18404), .ZN(n18411) );
  XNOR2_X1 U20435 ( .A(n24568), .B(n18407), .ZN(n18409) );
  XNOR2_X1 U20436 ( .A(n18532), .B(n1874), .ZN(n18408) );
  XNOR2_X1 U20437 ( .A(n18409), .B(n18408), .ZN(n18410) );
  XNOR2_X1 U20438 ( .A(n18412), .B(n18413), .ZN(n18417) );
  XNOR2_X1 U20439 ( .A(n18415), .B(n18414), .ZN(n18416) );
  XNOR2_X1 U20440 ( .A(n18417), .B(n18416), .ZN(n19015) );
  INV_X1 U20441 ( .A(n19015), .ZN(n19164) );
  XNOR2_X1 U20443 ( .A(n18422), .B(n18421), .ZN(n18427) );
  XNOR2_X1 U20444 ( .A(n18423), .B(n1746), .ZN(n18424) );
  XNOR2_X1 U20445 ( .A(n18424), .B(n18425), .ZN(n18426) );
  XNOR2_X1 U20447 ( .A(n18431), .B(n1724), .ZN(n18433) );
  XNOR2_X1 U20448 ( .A(n18432), .B(n18433), .ZN(n18434) );
  NOR2_X1 U20449 ( .A1(n18788), .A2(n24326), .ZN(n18442) );
  XNOR2_X1 U20450 ( .A(n18435), .B(n18539), .ZN(n18436) );
  XNOR2_X1 U20451 ( .A(n18439), .B(n18438), .ZN(n18440) );
  NOR2_X1 U20452 ( .A1(n20094), .A2(n20567), .ZN(n18444) );
  XNOR2_X1 U20453 ( .A(n21559), .B(n21699), .ZN(n18710) );
  XNOR2_X1 U20454 ( .A(n18602), .B(n18446), .ZN(n18450) );
  XNOR2_X1 U20455 ( .A(n18448), .B(n18447), .ZN(n18449) );
  XNOR2_X1 U20456 ( .A(n18450), .B(n18449), .ZN(n18455) );
  XNOR2_X1 U20457 ( .A(n18451), .B(n24287), .ZN(n18452) );
  XNOR2_X1 U20458 ( .A(n18453), .B(n18452), .ZN(n18454) );
  XNOR2_X1 U20459 ( .A(n18454), .B(n18455), .ZN(n19061) );
  INV_X1 U20460 ( .A(n19061), .ZN(n19007) );
  XNOR2_X1 U20461 ( .A(n18458), .B(n18457), .ZN(n18462) );
  XNOR2_X1 U20462 ( .A(n18460), .B(n18459), .ZN(n18461) );
  XNOR2_X1 U20463 ( .A(n18465), .B(n18466), .ZN(n18469) );
  XNOR2_X1 U20464 ( .A(n18467), .B(n2236), .ZN(n18468) );
  XNOR2_X1 U20465 ( .A(n18469), .B(n18468), .ZN(n18470) );
  NAND3_X1 U20466 ( .A1(n19007), .A2(n280), .A3(n1002), .ZN(n18498) );
  XNOR2_X1 U20467 ( .A(n18473), .B(n18472), .ZN(n18474) );
  XNOR2_X1 U20468 ( .A(n18475), .B(n18474), .ZN(n18480) );
  XNOR2_X1 U20469 ( .A(n18476), .B(n20284), .ZN(n18477) );
  XNOR2_X1 U20470 ( .A(n18478), .B(n18477), .ZN(n18479) );
  OR3_X1 U20471 ( .A1(n19061), .A2(n19575), .A3(n1002), .ZN(n18497) );
  XNOR2_X1 U20472 ( .A(n18481), .B(n18482), .ZN(n18488) );
  XNOR2_X1 U20473 ( .A(n18483), .B(n18531), .ZN(n18486) );
  XNOR2_X1 U20474 ( .A(n18484), .B(n1767), .ZN(n18485) );
  XNOR2_X1 U20475 ( .A(n18486), .B(n18485), .ZN(n18487) );
  XNOR2_X1 U20476 ( .A(n18489), .B(n2193), .ZN(n18490) );
  XNOR2_X1 U20477 ( .A(n18493), .B(n18494), .ZN(n19059) );
  OR3_X1 U20478 ( .A1(n19007), .A2(n24982), .A3(n19059), .ZN(n18496) );
  NAND2_X1 U20479 ( .A1(n1443), .A2(n1002), .ZN(n18495) );
  XNOR2_X1 U20481 ( .A(n18499), .B(n22702), .ZN(n18500) );
  XNOR2_X1 U20482 ( .A(n18500), .B(n18677), .ZN(n18502) );
  XNOR2_X1 U20483 ( .A(n18502), .B(n18501), .ZN(n18504) );
  INV_X1 U20484 ( .A(n18505), .ZN(n18511) );
  XNOR2_X1 U20485 ( .A(n18695), .B(n2745), .ZN(n18507) );
  XNOR2_X1 U20486 ( .A(n18507), .B(n18506), .ZN(n18508) );
  XNOR2_X1 U20487 ( .A(n18508), .B(n18509), .ZN(n18510) );
  INV_X1 U20488 ( .A(n3178), .ZN(n22385) );
  XNOR2_X1 U20489 ( .A(n18512), .B(n22385), .ZN(n18514) );
  XNOR2_X1 U20490 ( .A(n18514), .B(n18513), .ZN(n18518) );
  XNOR2_X1 U20491 ( .A(n18516), .B(n18515), .ZN(n18517) );
  XNOR2_X1 U20492 ( .A(n18518), .B(n18517), .ZN(n18519) );
  XNOR2_X1 U20493 ( .A(n18522), .B(n18521), .ZN(n18527) );
  XNOR2_X1 U20494 ( .A(n18523), .B(n891), .ZN(n18525) );
  XNOR2_X1 U20495 ( .A(n18524), .B(n18525), .ZN(n18526) );
  XNOR2_X1 U20497 ( .A(n18529), .B(n18528), .ZN(n18536) );
  XNOR2_X1 U20498 ( .A(n18531), .B(n18530), .ZN(n18534) );
  XNOR2_X1 U20499 ( .A(n18532), .B(n888), .ZN(n18533) );
  XNOR2_X1 U20500 ( .A(n18534), .B(n18533), .ZN(n18535) );
  XNOR2_X1 U20501 ( .A(n18536), .B(n18535), .ZN(n19066) );
  XNOR2_X1 U20502 ( .A(n18538), .B(n18537), .ZN(n18545) );
  XNOR2_X1 U20503 ( .A(n18540), .B(n18539), .ZN(n18543) );
  XNOR2_X1 U20504 ( .A(n18541), .B(n2034), .ZN(n18542) );
  XNOR2_X1 U20505 ( .A(n18543), .B(n18542), .ZN(n18544) );
  XNOR2_X1 U20507 ( .A(n18548), .B(n18549), .ZN(n18551) );
  XNOR2_X1 U20508 ( .A(n18550), .B(n18551), .ZN(n18556) );
  XNOR2_X1 U20509 ( .A(n18552), .B(n17476), .ZN(n18555) );
  INV_X1 U20511 ( .A(n18557), .ZN(n18558) );
  XNOR2_X1 U20512 ( .A(n18559), .B(n18558), .ZN(n18561) );
  XNOR2_X1 U20513 ( .A(n18560), .B(n18561), .ZN(n18566) );
  XNOR2_X1 U20514 ( .A(n364), .B(n18562), .ZN(n18564) );
  XNOR2_X1 U20515 ( .A(n25482), .B(n1864), .ZN(n18563) );
  XNOR2_X1 U20516 ( .A(n18564), .B(n18563), .ZN(n18565) );
  XNOR2_X1 U20517 ( .A(n18568), .B(n18567), .ZN(n18572) );
  XNOR2_X1 U20518 ( .A(n18570), .B(n18569), .ZN(n18571) );
  MUX2_X1 U20519 ( .A(n19084), .B(n19417), .S(n24584), .Z(n18595) );
  XNOR2_X1 U20520 ( .A(n18574), .B(n18573), .ZN(n18578) );
  XNOR2_X1 U20521 ( .A(n18576), .B(n18575), .ZN(n18577) );
  XNOR2_X1 U20522 ( .A(n18582), .B(n1758), .ZN(n18583) );
  XNOR2_X1 U20523 ( .A(n18584), .B(n18583), .ZN(n18585) );
  INV_X1 U20524 ( .A(n19420), .ZN(n19083) );
  AND2_X1 U20525 ( .A1(n19088), .A2(n18586), .ZN(n18594) );
  XNOR2_X1 U20526 ( .A(n18588), .B(n18587), .ZN(n18593) );
  INV_X1 U20527 ( .A(n899), .ZN(n22739) );
  XNOR2_X1 U20528 ( .A(n24565), .B(n22739), .ZN(n18590) );
  XNOR2_X1 U20529 ( .A(n18591), .B(n18590), .ZN(n18592) );
  NAND3_X1 U20530 ( .A1(n18597), .A2(n25195), .A3(n18777), .ZN(n18598) );
  XNOR2_X1 U20531 ( .A(n18600), .B(n18599), .ZN(n18604) );
  XNOR2_X1 U20532 ( .A(n18602), .B(n18601), .ZN(n18603) );
  XNOR2_X1 U20533 ( .A(n18603), .B(n18604), .ZN(n18609) );
  XNOR2_X1 U20534 ( .A(n18605), .B(n2772), .ZN(n18606) );
  XNOR2_X1 U20535 ( .A(n18607), .B(n18606), .ZN(n18608) );
  XNOR2_X1 U20536 ( .A(n18609), .B(n18608), .ZN(n19436) );
  XNOR2_X1 U20537 ( .A(n18611), .B(n18610), .ZN(n18614) );
  XNOR2_X1 U20538 ( .A(n18613), .B(n18614), .ZN(n18618) );
  XNOR2_X1 U20539 ( .A(n18616), .B(n18615), .ZN(n18617) );
  XNOR2_X1 U20540 ( .A(n18620), .B(n18619), .ZN(n18625) );
  XNOR2_X1 U20541 ( .A(n18621), .B(n1924), .ZN(n18622) );
  XNOR2_X1 U20542 ( .A(n18623), .B(n18622), .ZN(n18624) );
  XNOR2_X1 U20543 ( .A(n18627), .B(n18626), .ZN(n18632) );
  XNOR2_X1 U20544 ( .A(n25482), .B(n2757), .ZN(n18630) );
  XNOR2_X1 U20545 ( .A(n18630), .B(n18629), .ZN(n18631) );
  INV_X1 U20546 ( .A(n19438), .ZN(n18642) );
  XNOR2_X1 U20547 ( .A(n18635), .B(n18634), .ZN(n18641) );
  XNOR2_X1 U20548 ( .A(n18637), .B(n25493), .ZN(n18639) );
  XNOR2_X1 U20549 ( .A(n18639), .B(n18638), .ZN(n18640) );
  XNOR2_X1 U20550 ( .A(n18641), .B(n18640), .ZN(n18832) );
  OAI21_X1 U20551 ( .B1(n5007), .B2(n19245), .A(n18643), .ZN(n18655) );
  XNOR2_X1 U20552 ( .A(n18645), .B(n18644), .ZN(n18650) );
  XNOR2_X1 U20553 ( .A(n18646), .B(n20690), .ZN(n18647) );
  XNOR2_X1 U20554 ( .A(n18648), .B(n18647), .ZN(n18649) );
  XNOR2_X1 U20555 ( .A(n18650), .B(n18649), .ZN(n18834) );
  INV_X1 U20556 ( .A(n18834), .ZN(n19081) );
  OAI21_X1 U20557 ( .B1(n19081), .B2(n25260), .A(n18651), .ZN(n18653) );
  NOR2_X1 U20558 ( .A1(n18653), .A2(n19435), .ZN(n18654) );
  NOR2_X1 U20559 ( .A1(n24835), .A2(n20569), .ZN(n18706) );
  XNOR2_X1 U20560 ( .A(n18656), .B(n18657), .ZN(n18664) );
  XNOR2_X1 U20561 ( .A(n18659), .B(n18658), .ZN(n18662) );
  XNOR2_X1 U20562 ( .A(n18660), .B(n1757), .ZN(n18661) );
  XNOR2_X1 U20563 ( .A(n18662), .B(n18661), .ZN(n18663) );
  INV_X1 U20564 ( .A(n18690), .ZN(n19170) );
  XNOR2_X1 U20565 ( .A(n18666), .B(n18665), .ZN(n18668) );
  XNOR2_X1 U20567 ( .A(n18669), .B(n2990), .ZN(n18670) );
  XNOR2_X1 U20568 ( .A(n18671), .B(n18670), .ZN(n18672) );
  XNOR2_X1 U20569 ( .A(n18674), .B(n18675), .ZN(n18676) );
  XNOR2_X1 U20570 ( .A(n18677), .B(n18676), .ZN(n18682) );
  XNOR2_X1 U20571 ( .A(n18678), .B(n2031), .ZN(n18679) );
  XNOR2_X1 U20572 ( .A(n18684), .B(n18683), .ZN(n18689) );
  XNOR2_X1 U20573 ( .A(n18685), .B(n1863), .ZN(n18686) );
  XNOR2_X1 U20574 ( .A(n18687), .B(n18686), .ZN(n18688) );
  XNOR2_X1 U20575 ( .A(n18688), .B(n18689), .ZN(n19406) );
  INV_X1 U20576 ( .A(n19406), .ZN(n19169) );
  XNOR2_X1 U20577 ( .A(n18692), .B(n18691), .ZN(n18699) );
  XNOR2_X1 U20578 ( .A(n18694), .B(n18693), .ZN(n18697) );
  XNOR2_X1 U20579 ( .A(n18695), .B(n2044), .ZN(n18696) );
  XNOR2_X1 U20580 ( .A(n18697), .B(n18696), .ZN(n18698) );
  NOR2_X1 U20582 ( .A1(n20617), .A2(n20615), .ZN(n18705) );
  AOI22_X1 U20583 ( .A1(n18706), .A2(n20614), .B1(n24338), .B2(n18705), .ZN(
        n18708) );
  NAND2_X1 U20584 ( .A1(n24338), .A2(n20623), .ZN(n18707) );
  OAI211_X1 U20585 ( .C1(n20619), .C2(n24338), .A(n18708), .B(n18707), .ZN(
        n20742) );
  XNOR2_X1 U20586 ( .A(n20742), .B(n2190), .ZN(n18709) );
  XNOR2_X1 U20587 ( .A(n18710), .B(n18709), .ZN(n18711) );
  NAND2_X1 U20589 ( .A1(n19357), .A2(n19444), .ZN(n18717) );
  OR3_X1 U20590 ( .A1(n19357), .A2(n19451), .A3(n19452), .ZN(n18716) );
  NAND2_X1 U20591 ( .A1(n25002), .A2(n19446), .ZN(n18714) );
  NAND2_X1 U20592 ( .A1(n18990), .A2(n19445), .ZN(n19351) );
  INV_X1 U20593 ( .A(n19498), .ZN(n18718) );
  NAND3_X1 U20595 ( .A1(n18724), .A2(n19371), .A3(n24361), .ZN(n18725) );
  NAND2_X1 U20596 ( .A1(n19345), .A2(n19346), .ZN(n18728) );
  OAI21_X1 U20597 ( .B1(n19487), .B2(n240), .A(n18727), .ZN(n19208) );
  NAND2_X1 U20598 ( .A1(n19230), .A2(n18729), .ZN(n18743) );
  NAND2_X1 U20599 ( .A1(n18730), .A2(n19477), .ZN(n18733) );
  INV_X1 U20600 ( .A(n19478), .ZN(n18731) );
  NAND2_X1 U20601 ( .A1(n19476), .A2(n18731), .ZN(n18732) );
  MUX2_X1 U20602 ( .A(n18733), .B(n18732), .S(n19482), .Z(n18738) );
  INV_X1 U20603 ( .A(n18734), .ZN(n18974) );
  NOR2_X1 U20604 ( .A1(n18735), .A2(n18974), .ZN(n18736) );
  OAI21_X1 U20605 ( .B1(n18971), .B2(n18736), .A(n19478), .ZN(n18737) );
  NAND3_X1 U20606 ( .A1(n18739), .A2(n18979), .A3(n19028), .ZN(n18740) );
  OAI21_X1 U20608 ( .B1(n20191), .B2(n20185), .A(n25478), .ZN(n18742) );
  XNOR2_X1 U20610 ( .A(n21135), .B(n1745), .ZN(n18746) );
  NAND2_X1 U20611 ( .A1(n20336), .A2(n20669), .ZN(n18744) );
  NAND2_X1 U20612 ( .A1(n18744), .A2(n20668), .ZN(n18745) );
  NAND2_X1 U20613 ( .A1(n19309), .A2(n19311), .ZN(n18921) );
  NAND2_X1 U20614 ( .A1(n18921), .A2(n19313), .ZN(n18748) );
  NOR2_X1 U20615 ( .A1(n19309), .A2(n19312), .ZN(n18747) );
  NOR2_X1 U20616 ( .A1(n3284), .A2(n19555), .ZN(n18750) );
  INV_X1 U20617 ( .A(n19556), .ZN(n19558) );
  MUX2_X1 U20618 ( .A(n18752), .B(n18750), .S(n19558), .Z(n18754) );
  OAI21_X1 U20619 ( .B1(n19560), .B2(n4262), .A(n3284), .ZN(n18751) );
  NOR2_X1 U20620 ( .A1(n18752), .A2(n18751), .ZN(n18753) );
  INV_X1 U20621 ( .A(n19266), .ZN(n18917) );
  NOR2_X1 U20622 ( .A1(n18919), .A2(n18917), .ZN(n18758) );
  NOR2_X1 U20623 ( .A1(n18756), .A2(n24386), .ZN(n18757) );
  NOR2_X1 U20624 ( .A1(n18758), .A2(n18757), .ZN(n18760) );
  MUX2_X1 U20625 ( .A(n19531), .B(n19534), .S(n24393), .Z(n18763) );
  INV_X1 U20626 ( .A(n18762), .ZN(n19530) );
  NAND2_X1 U20627 ( .A1(n19535), .A2(n19532), .ZN(n18764) );
  NOR2_X1 U20629 ( .A1(n24441), .A2(n18767), .ZN(n18770) );
  INV_X1 U20631 ( .A(n18772), .ZN(n19540) );
  AOI22_X1 U20632 ( .A1(n5573), .A2(n19539), .B1(n19540), .B2(n1334), .ZN(
        n18773) );
  MUX2_X1 U20633 ( .A(n19546), .B(n19185), .S(n19548), .Z(n18775) );
  NAND3_X1 U20635 ( .A1(n24758), .A2(n19177), .A3(n19179), .ZN(n18781) );
  AOI21_X1 U20636 ( .B1(n19427), .B2(n19177), .A(n1361), .ZN(n18776) );
  OAI21_X1 U20637 ( .B1(n19183), .B2(n19427), .A(n18776), .ZN(n18780) );
  NOR2_X1 U20638 ( .A1(n18777), .A2(n19428), .ZN(n18778) );
  NAND2_X1 U20639 ( .A1(n19183), .A2(n18778), .ZN(n18779) );
  INV_X1 U20640 ( .A(n19173), .ZN(n19411) );
  AND2_X1 U20641 ( .A1(n19413), .A2(n19406), .ZN(n19172) );
  INV_X1 U20642 ( .A(n19172), .ZN(n18784) );
  NOR2_X1 U20644 ( .A1(n20060), .A2(n25088), .ZN(n19641) );
  NAND2_X1 U20645 ( .A1(n20470), .A2(n19641), .ZN(n18803) );
  INV_X1 U20646 ( .A(n24326), .ZN(n18899) );
  INV_X1 U20647 ( .A(n18788), .ZN(n19396) );
  OAI21_X1 U20648 ( .B1(n18790), .B2(n18899), .A(n18789), .ZN(n18792) );
  NOR2_X1 U20649 ( .A1(n19191), .A2(n1053), .ZN(n18794) );
  NAND2_X1 U20650 ( .A1(n19192), .A2(n19568), .ZN(n18793) );
  INV_X1 U20651 ( .A(n19518), .ZN(n18795) );
  AOI22_X1 U20652 ( .A1(n18897), .A2(n19522), .B1(n19523), .B2(n19521), .ZN(
        n18799) );
  INV_X1 U20653 ( .A(n19284), .ZN(n19519) );
  NAND2_X1 U20654 ( .A1(n19279), .A2(n19519), .ZN(n18797) );
  MUX2_X1 U20655 ( .A(n18797), .B(n18796), .S(n19518), .Z(n18798) );
  OAI21_X1 U20656 ( .B1(n25490), .B2(n19928), .A(n20062), .ZN(n18800) );
  NAND2_X1 U20658 ( .A1(n18800), .A2(n5115), .ZN(n18802) );
  INV_X1 U20659 ( .A(n20060), .ZN(n19121) );
  NAND3_X1 U20660 ( .A1(n20062), .A2(n20055), .A3(n19121), .ZN(n18801) );
  XNOR2_X1 U20661 ( .A(n21084), .B(n21212), .ZN(n21696) );
  NAND2_X1 U20662 ( .A1(n19233), .A2(n19607), .ZN(n19113) );
  NOR2_X1 U20663 ( .A1(n19237), .A2(n19112), .ZN(n18804) );
  NOR2_X1 U20664 ( .A1(n19113), .A2(n18804), .ZN(n18805) );
  INV_X1 U20665 ( .A(n20359), .ZN(n20911) );
  INV_X1 U20666 ( .A(n19591), .ZN(n19250) );
  INV_X1 U20667 ( .A(n18806), .ZN(n18807) );
  INV_X1 U20668 ( .A(n19199), .ZN(n19581) );
  MUX2_X1 U20669 ( .A(n19198), .B(n18809), .S(n19581), .Z(n18811) );
  INV_X1 U20670 ( .A(n19105), .ZN(n19582) );
  INV_X1 U20671 ( .A(n19107), .ZN(n19586) );
  OAI21_X1 U20672 ( .B1(n19582), .B2(n19581), .A(n19202), .ZN(n18810) );
  NOR2_X1 U20673 ( .A1(n24909), .A2(n19021), .ZN(n19108) );
  INV_X1 U20674 ( .A(n19108), .ZN(n18815) );
  OAI21_X1 U20676 ( .B1(n24931), .B2(n19389), .A(n25052), .ZN(n18813) );
  AND2_X1 U20677 ( .A1(n19386), .A2(n19217), .ZN(n19631) );
  INV_X1 U20678 ( .A(n19021), .ZN(n19630) );
  NAND2_X1 U20679 ( .A1(n19631), .A2(n19630), .ZN(n18814) );
  AOI22_X1 U20680 ( .A1(n20911), .A2(n20909), .B1(n20913), .B2(n20491), .ZN(
        n20363) );
  INV_X1 U20681 ( .A(n19041), .ZN(n18816) );
  NAND2_X1 U20682 ( .A1(n18817), .A2(n25392), .ZN(n18818) );
  OAI21_X1 U20685 ( .B1(n19380), .B2(n24452), .A(n18819), .ZN(n18821) );
  NOR2_X1 U20686 ( .A1(n19382), .A2(n18876), .ZN(n19205) );
  NAND3_X1 U20688 ( .A1(n25067), .A2(n24318), .A3(n19094), .ZN(n18820) );
  OAI21_X1 U20689 ( .B1(n18821), .B2(n19205), .A(n18820), .ZN(n18823) );
  NOR2_X1 U20690 ( .A1(n19379), .A2(n19377), .ZN(n18822) );
  NAND2_X1 U20692 ( .A1(n20487), .A2(n20909), .ZN(n18824) );
  NAND2_X1 U20693 ( .A1(n18824), .A2(n347), .ZN(n18825) );
  MUX2_X1 U20695 ( .A(n18826), .B(n19406), .S(n19408), .Z(n18827) );
  INV_X1 U20696 ( .A(n19417), .ZN(n19087) );
  NAND2_X1 U20697 ( .A1(n19419), .A2(n19084), .ZN(n18829) );
  NOR2_X1 U20698 ( .A1(n19166), .A2(n19084), .ZN(n18828) );
  NAND2_X1 U20699 ( .A1(n25423), .A2(n361), .ZN(n18833) );
  INV_X1 U20700 ( .A(n19065), .ZN(n19241) );
  INV_X1 U20701 ( .A(n19066), .ZN(n19615) );
  MUX2_X1 U20702 ( .A(n18837), .B(n18836), .S(n19615), .Z(n18838) );
  INV_X1 U20703 ( .A(n20478), .ZN(n18839) );
  XNOR2_X1 U20705 ( .A(n21572), .B(n25073), .ZN(n20954) );
  INV_X1 U20706 ( .A(n18959), .ZN(n18944) );
  INV_X1 U20708 ( .A(n19470), .ZN(n19322) );
  INV_X1 U20709 ( .A(n19321), .ZN(n19467) );
  AOI21_X1 U20710 ( .B1(n18842), .B2(n18925), .A(n18841), .ZN(n18845) );
  OAI22_X1 U20711 ( .A1(n18923), .A2(n18843), .B1(n19317), .B2(n24912), .ZN(
        n18844) );
  NOR2_X1 U20712 ( .A1(n357), .A2(n19501), .ZN(n18847) );
  INV_X1 U20713 ( .A(n19480), .ZN(n18851) );
  NOR2_X1 U20714 ( .A1(n18974), .A2(n19476), .ZN(n18849) );
  NAND2_X1 U20715 ( .A1(n18971), .A2(n19479), .ZN(n18850) );
  AND2_X1 U20716 ( .A1(n19658), .A2(n20068), .ZN(n19194) );
  AOI21_X1 U20717 ( .B1(n20071), .B2(n19660), .A(n19194), .ZN(n18859) );
  INV_X1 U20718 ( .A(n19329), .ZN(n18935) );
  MUX2_X1 U20719 ( .A(n24583), .B(n25566), .S(n18935), .Z(n18855) );
  NAND2_X1 U20720 ( .A1(n5736), .A2(n18934), .ZN(n18854) );
  AND2_X1 U20721 ( .A1(n19329), .A2(n19328), .ZN(n18938) );
  INV_X1 U20722 ( .A(n19195), .ZN(n19850) );
  NAND2_X1 U20723 ( .A1(n19297), .A2(n24427), .ZN(n18856) );
  NAND3_X1 U20724 ( .A1(n24457), .A2(n19297), .A3(n356), .ZN(n18857) );
  INV_X1 U20725 ( .A(n20068), .ZN(n20073) );
  AOI21_X1 U20726 ( .B1(n19849), .B2(n19658), .A(n20073), .ZN(n18858) );
  XNOR2_X1 U20728 ( .A(n20954), .B(n25222), .ZN(n18860) );
  NAND2_X1 U20730 ( .A1(n18865), .A2(n18864), .ZN(n18866) );
  INV_X1 U20732 ( .A(n19596), .ZN(n18871) );
  OAI21_X1 U20733 ( .B1(n18037), .B2(n19601), .A(n19254), .ZN(n18874) );
  NAND3_X1 U20734 ( .A1(n19071), .A2(n18871), .A3(n19601), .ZN(n18872) );
  NOR2_X1 U20735 ( .A1(n20289), .A2(n19668), .ZN(n18887) );
  OAI22_X1 U20736 ( .A1(n24335), .A2(n24318), .B1(n24452), .B2(n19094), .ZN(
        n19206) );
  NAND2_X1 U20737 ( .A1(n19382), .A2(n18876), .ZN(n19093) );
  MUX2_X1 U20740 ( .A(n19581), .B(n19580), .S(n19198), .Z(n18882) );
  NAND2_X1 U20741 ( .A1(n19105), .A2(n19107), .ZN(n18881) );
  INV_X1 U20742 ( .A(n21009), .ZN(n20530) );
  INV_X1 U20743 ( .A(n21008), .ZN(n20528) );
  INV_X1 U20744 ( .A(n19066), .ZN(n18883) );
  INV_X1 U20745 ( .A(n19067), .ZN(n19614) );
  NAND2_X1 U20746 ( .A1(n18884), .A2(n19239), .ZN(n18885) );
  INV_X1 U20748 ( .A(n19546), .ZN(n18889) );
  INV_X1 U20751 ( .A(n19402), .ZN(n19549) );
  NAND3_X1 U20752 ( .A1(n19552), .A2(n19549), .A3(n19186), .ZN(n18892) );
  NAND3_X1 U20753 ( .A1(n24929), .A2(n18889), .A3(n1711), .ZN(n18891) );
  NAND3_X1 U20754 ( .A1(n24929), .A2(n19185), .A3(n19546), .ZN(n18890) );
  NAND2_X1 U20755 ( .A1(n18894), .A2(n19522), .ZN(n18898) );
  NOR2_X1 U20756 ( .A1(n19526), .A2(n19523), .ZN(n18896) );
  NAND2_X1 U20757 ( .A1(n20126), .A2(n20309), .ZN(n20548) );
  NAND2_X1 U20758 ( .A1(n19540), .A2(n19543), .ZN(n18904) );
  OAI21_X1 U20759 ( .B1(n1334), .B2(n19126), .A(n19275), .ZN(n18903) );
  INV_X1 U20760 ( .A(n19276), .ZN(n18905) );
  NOR2_X1 U20762 ( .A1(n19191), .A2(n363), .ZN(n18908) );
  NAND2_X1 U20763 ( .A1(n19555), .A2(n24421), .ZN(n18912) );
  INV_X1 U20764 ( .A(n19290), .ZN(n19554) );
  NAND3_X1 U20765 ( .A1(n19554), .A2(n19559), .A3(n19555), .ZN(n18911) );
  INV_X1 U20766 ( .A(n20127), .ZN(n20543) );
  NAND3_X1 U20767 ( .A1(n20130), .A2(n20545), .A3(n20543), .ZN(n18913) );
  XNOR2_X1 U20768 ( .A(n21678), .B(n21597), .ZN(n21116) );
  INV_X1 U20769 ( .A(n19263), .ZN(n19150) );
  INV_X1 U20770 ( .A(n18921), .ZN(n18922) );
  NAND3_X1 U20771 ( .A1(n18923), .A2(n5371), .A3(n19313), .ZN(n18924) );
  OAI21_X1 U20772 ( .B1(n18925), .B2(n19312), .A(n18924), .ZN(n18926) );
  INV_X1 U20773 ( .A(n18928), .ZN(n18931) );
  AND2_X1 U20774 ( .A1(n19297), .A2(n18929), .ZN(n19301) );
  INV_X1 U20775 ( .A(n19301), .ZN(n18930) );
  AOI22_X2 U20776 ( .A1(n18968), .A2(n18932), .B1(n18930), .B2(n18931), .ZN(
        n19785) );
  MUX2_X1 U20777 ( .A(n19684), .B(n19984), .S(n19785), .Z(n18942) );
  NOR2_X1 U20778 ( .A1(n18934), .A2(n18933), .ZN(n18937) );
  NOR2_X2 U20779 ( .A1(n18941), .A2(n18940), .ZN(n19987) );
  NOR2_X1 U20780 ( .A1(n18942), .A2(n24979), .ZN(n18955) );
  NOR2_X1 U20781 ( .A1(n19472), .A2(n19467), .ZN(n18943) );
  MUX2_X1 U20782 ( .A(n19466), .B(n18943), .S(n18959), .Z(n18946) );
  INV_X1 U20783 ( .A(n19472), .ZN(n18956) );
  NAND2_X1 U20784 ( .A1(n19984), .A2(n24464), .ZN(n18953) );
  NAND2_X1 U20786 ( .A1(n19303), .A2(n18947), .ZN(n18948) );
  AND2_X1 U20787 ( .A1(n19306), .A2(n18948), .ZN(n18952) );
  NOR2_X1 U20789 ( .A1(n25364), .A2(n19128), .ZN(n18950) );
  AOI22_X1 U20790 ( .A1(n24441), .A2(n18950), .B1(n18949), .B2(n24324), .ZN(
        n18951) );
  OAI22_X1 U20791 ( .A1(n19986), .A2(n18953), .B1(n24315), .B2(n19786), .ZN(
        n18954) );
  NOR2_X1 U20792 ( .A1(n18955), .A2(n18954), .ZN(n20767) );
  NOR2_X1 U20794 ( .A1(n19466), .A2(n19321), .ZN(n18957) );
  AOI21_X1 U20796 ( .B1(n18962), .B2(n18961), .A(n18960), .ZN(n18963) );
  NAND2_X1 U20798 ( .A1(n19296), .A2(n24427), .ZN(n18966) );
  AND2_X1 U20799 ( .A1(n4075), .A2(n18966), .ZN(n18969) );
  NAND2_X1 U20801 ( .A1(n18971), .A2(n19476), .ZN(n18972) );
  INV_X1 U20802 ( .A(n19459), .ZN(n18976) );
  NAND2_X1 U20803 ( .A1(n18976), .A2(n19457), .ZN(n19030) );
  NAND3_X1 U20804 ( .A1(n19030), .A2(n18979), .A3(n18977), .ZN(n18981) );
  OAI21_X1 U20805 ( .B1(n19030), .B2(n19464), .A(n18978), .ZN(n18980) );
  AOI21_X2 U20806 ( .B1(n18980), .B2(n18981), .A(n19029), .ZN(n20019) );
  OAI211_X1 U20807 ( .C1(n25459), .C2(n19501), .A(n358), .B(n19334), .ZN(
        n18988) );
  NAND2_X1 U20808 ( .A1(n19500), .A2(n18983), .ZN(n18984) );
  OAI211_X1 U20809 ( .C1(n18987), .C2(n19501), .A(n18988), .B(n18984), .ZN(
        n18985) );
  NOR2_X1 U20810 ( .A1(n20136), .A2(n20014), .ZN(n18991) );
  NAND2_X1 U20812 ( .A1(n18991), .A2(n19755), .ZN(n20925) );
  XNOR2_X1 U20813 ( .A(n20767), .B(n21523), .ZN(n20439) );
  XNOR2_X1 U20814 ( .A(n21116), .B(n20439), .ZN(n19054) );
  NAND2_X1 U20815 ( .A1(n20317), .A2(n18994), .ZN(n18993) );
  INV_X1 U20816 ( .A(n19889), .ZN(n20320) );
  MUX2_X1 U20818 ( .A(n18993), .B(n18992), .S(n20319), .Z(n18997) );
  AND2_X1 U20819 ( .A1(n19714), .A2(n20316), .ZN(n18995) );
  AOI22_X1 U20820 ( .A1(n19888), .A2(n24917), .B1(n18995), .B2(n341), .ZN(
        n18996) );
  NOR2_X1 U20822 ( .A1(n19417), .A2(n19418), .ZN(n18999) );
  AOI22_X1 U20823 ( .A1(n19000), .A2(n18998), .B1(n24584), .B2(n18999), .ZN(
        n19001) );
  NOR2_X1 U20824 ( .A1(n18385), .A2(n19177), .ZN(n19180) );
  AND2_X1 U20825 ( .A1(n19003), .A2(n19177), .ZN(n19005) );
  OAI211_X1 U20826 ( .C1(n19179), .C2(n19760), .A(n19176), .B(n25195), .ZN(
        n19004) );
  NOR2_X1 U20827 ( .A1(n20536), .A2(n20537), .ZN(n19689) );
  OAI21_X1 U20828 ( .B1(n280), .B2(n354), .A(n1002), .ZN(n19006) );
  INV_X1 U20830 ( .A(n20537), .ZN(n19011) );
  MUX2_X1 U20831 ( .A(n19413), .B(n19407), .S(n19170), .Z(n19010) );
  NAND2_X1 U20832 ( .A1(n19173), .A2(n19413), .ZN(n19009) );
  OAI21_X1 U20833 ( .B1(n20149), .B2(n19011), .A(n20447), .ZN(n19012) );
  MUX2_X1 U20835 ( .A(n18834), .B(n361), .S(n19438), .Z(n19013) );
  NAND2_X1 U20836 ( .A1(n20533), .A2(n20149), .ZN(n19019) );
  NAND2_X1 U20837 ( .A1(n19397), .A2(n19164), .ZN(n19014) );
  NAND2_X1 U20838 ( .A1(n19016), .A2(n19396), .ZN(n19017) );
  INV_X1 U20839 ( .A(n20445), .ZN(n19018) );
  XNOR2_X1 U20840 ( .A(n21679), .B(n21639), .ZN(n21096) );
  NAND2_X1 U20841 ( .A1(n24451), .A2(n19021), .ZN(n19391) );
  NAND2_X1 U20842 ( .A1(n19384), .A2(n25052), .ZN(n19022) );
  OAI21_X1 U20843 ( .B1(n19024), .B2(n19490), .A(n19023), .ZN(n19027) );
  MUX2_X1 U20844 ( .A(n19345), .B(n240), .S(n19488), .Z(n19025) );
  NOR2_X1 U20845 ( .A1(n19025), .A2(n25473), .ZN(n19026) );
  NAND2_X1 U20848 ( .A1(n19452), .A2(n19444), .ZN(n19039) );
  NOR2_X1 U20849 ( .A1(n18816), .A2(n19210), .ZN(n19043) );
  MUX2_X1 U20850 ( .A(n19043), .B(n19042), .S(n24312), .Z(n19046) );
  NAND2_X1 U20851 ( .A1(n19361), .A2(n19210), .ZN(n19044) );
  OAI22_X1 U20852 ( .A1(n19211), .A2(n19044), .B1(n19103), .B2(n24312), .ZN(
        n19045) );
  NAND2_X1 U20853 ( .A1(n19047), .A2(n20297), .ZN(n19048) );
  INV_X1 U20854 ( .A(n2126), .ZN(n19051) );
  XNOR2_X1 U20855 ( .A(n20870), .B(n19051), .ZN(n19052) );
  XNOR2_X1 U20856 ( .A(n21096), .B(n19052), .ZN(n19053) );
  OAI21_X1 U20859 ( .B1(n19615), .B2(n24606), .A(n355), .ZN(n19070) );
  NOR2_X1 U20860 ( .A1(n19065), .A2(n19064), .ZN(n19243) );
  NAND2_X1 U20861 ( .A1(n19243), .A2(n25086), .ZN(n19069) );
  NAND2_X1 U20862 ( .A1(n19067), .A2(n19613), .ZN(n19068) );
  NOR2_X1 U20863 ( .A1(n18037), .A2(n19602), .ZN(n19076) );
  NOR3_X1 U20864 ( .A1(n19071), .A2(n18037), .A3(n19598), .ZN(n19072) );
  NOR2_X1 U20865 ( .A1(n19073), .A2(n19072), .ZN(n19074) );
  NOR2_X1 U20866 ( .A1(n19591), .A2(n19077), .ZN(n19079) );
  INV_X1 U20867 ( .A(n20497), .ZN(n19904) );
  NAND3_X1 U20868 ( .A1(n24887), .A2(n20224), .A3(n20501), .ZN(n19090) );
  NAND3_X1 U20869 ( .A1(n24584), .A2(n19084), .A3(n19083), .ZN(n19086) );
  NAND3_X1 U20870 ( .A1(n19166), .A2(n19420), .A3(n19418), .ZN(n19085) );
  MUX2_X1 U20871 ( .A(n19382), .B(n19381), .S(n19092), .Z(n19096) );
  OAI21_X1 U20872 ( .B1(n19382), .B2(n19094), .A(n19093), .ZN(n19095) );
  AOI22_X1 U20874 ( .A1(n19363), .A2(n19376), .B1(n19098), .B2(n19097), .ZN(
        n19102) );
  NAND2_X1 U20875 ( .A1(n19100), .A2(n25243), .ZN(n19101) );
  NAND3_X1 U20876 ( .A1(n19103), .A2(n18816), .A3(n19359), .ZN(n19104) );
  NOR2_X1 U20877 ( .A1(n19386), .A2(n25052), .ZN(n19110) );
  AOI22_X1 U20878 ( .A1(n20276), .A2(n19924), .B1(n20517), .B2(n20272), .ZN(
        n19117) );
  OAI21_X1 U20879 ( .B1(n19235), .B2(n19237), .A(n19112), .ZN(n19116) );
  OAI21_X1 U20880 ( .B1(n19233), .B2(n19608), .A(n19113), .ZN(n19115) );
  INV_X1 U20881 ( .A(n19233), .ZN(n19606) );
  NOR2_X1 U20882 ( .A1(n18863), .A2(n19606), .ZN(n19114) );
  NAND2_X1 U20883 ( .A1(n20276), .A2(n20272), .ZN(n19118) );
  XNOR2_X1 U20884 ( .A(n21587), .B(n20826), .ZN(n21448) );
  OAI21_X1 U20885 ( .B1(n25388), .B2(n339), .A(n19917), .ZN(n19119) );
  AOI21_X2 U20886 ( .B1(n19120), .B2(n19119), .A(n19916), .ZN(n21686) );
  XNOR2_X1 U20887 ( .A(n21686), .B(n1528), .ZN(n19124) );
  INV_X1 U20888 ( .A(n20062), .ZN(n20472) );
  NAND2_X1 U20889 ( .A1(n20060), .A2(n20055), .ZN(n19122) );
  MUX2_X1 U20890 ( .A(n20472), .B(n19122), .S(n20054), .Z(n19123) );
  AOI21_X1 U20891 ( .B1(n19523), .B2(n19519), .A(n19520), .ZN(n19127) );
  NOR2_X1 U20892 ( .A1(n19133), .A2(n25364), .ZN(n19129) );
  OAI21_X1 U20893 ( .B1(n19130), .B2(n19129), .A(n24324), .ZN(n19137) );
  NAND3_X1 U20894 ( .A1(n19133), .A2(n19132), .A3(n25364), .ZN(n19134) );
  AND2_X1 U20895 ( .A1(n19135), .A2(n19134), .ZN(n19136) );
  AOI21_X1 U20896 ( .B1(n19743), .B2(n25421), .A(n20410), .ZN(n19154) );
  NAND2_X1 U20897 ( .A1(n19290), .A2(n19138), .ZN(n19139) );
  MUX2_X1 U20898 ( .A(n19562), .B(n19139), .S(n4262), .Z(n19144) );
  NOR2_X1 U20899 ( .A1(n19290), .A2(n24421), .ZN(n19142) );
  AOI22_X1 U20900 ( .A1(n19142), .A2(n19141), .B1(n19140), .B2(n3284), .ZN(
        n19143) );
  NOR3_X1 U20901 ( .A1(n4172), .A2(n19537), .A3(n19531), .ZN(n20257) );
  NAND2_X1 U20902 ( .A1(n20255), .A2(n25421), .ZN(n19911) );
  INV_X1 U20903 ( .A(n19911), .ZN(n19152) );
  AOI21_X2 U20905 ( .B1(n19150), .B2(n19149), .A(n19148), .ZN(n20262) );
  NOR2_X1 U20906 ( .A1(n20262), .A2(n20411), .ZN(n19151) );
  OAI21_X1 U20907 ( .B1(n19152), .B2(n19151), .A(n2024), .ZN(n19153) );
  OAI21_X1 U20908 ( .B1(n19154), .B2(n20263), .A(n19153), .ZN(n21228) );
  INV_X1 U20910 ( .A(n19697), .ZN(n20103) );
  INV_X1 U20911 ( .A(n19896), .ZN(n20104) );
  XNOR2_X1 U20912 ( .A(n21228), .B(n21266), .ZN(n19159) );
  NAND2_X1 U20913 ( .A1(n19849), .A2(n19851), .ZN(n20072) );
  NAND2_X1 U20914 ( .A1(n19658), .A2(n19852), .ZN(n19157) );
  MUX2_X1 U20915 ( .A(n20072), .B(n19157), .S(n19850), .Z(n19158) );
  XNOR2_X1 U20916 ( .A(n19159), .B(n21689), .ZN(n19160) );
  NOR2_X1 U20917 ( .A1(n18998), .A2(n19417), .ZN(n19423) );
  NAND2_X1 U20918 ( .A1(n19172), .A2(n19407), .ZN(n19175) );
  NOR2_X1 U20920 ( .A1(n19428), .A2(n19760), .ZN(n19178) );
  AOI22_X1 U20921 ( .A1(n19180), .A2(n19179), .B1(n19178), .B2(n25195), .ZN(
        n19181) );
  INV_X1 U20923 ( .A(n19185), .ZN(n19547) );
  NOR2_X1 U20924 ( .A1(n25057), .A2(n19547), .ZN(n19188) );
  NAND2_X1 U20925 ( .A1(n19402), .A2(n19186), .ZN(n19187) );
  OAI211_X1 U20926 ( .C1(n25223), .C2(n20216), .A(n25347), .B(n20510), .ZN(
        n19190) );
  NOR3_X1 U20927 ( .A1(n25224), .A2(n20510), .A3(n20199), .ZN(n19193) );
  NOR2_X1 U20928 ( .A1(n19194), .A2(n19660), .ZN(n19197) );
  OAI21_X1 U20930 ( .B1(n19195), .B2(n19660), .A(n19659), .ZN(n19196) );
  XNOR2_X1 U20931 ( .A(n20780), .B(n21514), .ZN(n21645) );
  NAND2_X1 U20932 ( .A1(n19584), .A2(n19198), .ZN(n19200) );
  MUX2_X1 U20933 ( .A(n19200), .B(n19586), .S(n24481), .Z(n19201) );
  OAI21_X1 U20934 ( .B1(n19345), .B2(n19346), .A(n2333), .ZN(n19207) );
  NAND2_X1 U20935 ( .A1(n19208), .A2(n5454), .ZN(n19209) );
  AOI21_X1 U20936 ( .B1(n19211), .B2(n19359), .A(n19361), .ZN(n19214) );
  NAND2_X1 U20937 ( .A1(n24940), .A2(n19841), .ZN(n19227) );
  NOR2_X1 U20938 ( .A1(n19219), .A2(n19367), .ZN(n19220) );
  AND2_X1 U20939 ( .A1(n19221), .A2(n19220), .ZN(n19223) );
  OAI211_X2 U20940 ( .C1(n20583), .C2(n20433), .A(n19227), .B(n19226), .ZN(
        n21728) );
  NOR2_X1 U20941 ( .A1(n20183), .A2(n25212), .ZN(n19231) );
  INV_X1 U20943 ( .A(n20182), .ZN(n20041) );
  NAND2_X1 U20944 ( .A1(n19228), .A2(n20041), .ZN(n19229) );
  OAI211_X1 U20945 ( .C1(n19231), .C2(n19662), .A(n19230), .B(n19229), .ZN(
        n21515) );
  XNOR2_X1 U20946 ( .A(n21728), .B(n21515), .ZN(n20842) );
  INV_X1 U20947 ( .A(n20842), .ZN(n19232) );
  XNOR2_X1 U20948 ( .A(n19232), .B(n21645), .ZN(n19342) );
  OAI21_X1 U20949 ( .B1(n19233), .B2(n19607), .A(n19608), .ZN(n19234) );
  NOR2_X1 U20950 ( .A1(n19241), .A2(n25012), .ZN(n19242) );
  NOR2_X1 U20951 ( .A1(n19243), .A2(n19242), .ZN(n19244) );
  NAND3_X1 U20952 ( .A1(n3986), .A2(n25260), .A3(n361), .ZN(n19247) );
  INV_X1 U20953 ( .A(n19576), .ZN(n19249) );
  MUX2_X1 U20954 ( .A(n19592), .B(n2346), .S(n19250), .Z(n19253) );
  NAND2_X1 U20955 ( .A1(n25476), .A2(n20428), .ZN(n19259) );
  NOR2_X1 U20956 ( .A1(n19255), .A2(n19598), .ZN(n19256) );
  AOI22_X1 U20957 ( .A1(n19257), .A2(n24079), .B1(n19597), .B2(n19256), .ZN(
        n19258) );
  NOR2_X1 U20959 ( .A1(n19264), .A2(n19261), .ZN(n19262) );
  NOR2_X1 U20960 ( .A1(n19263), .A2(n19262), .ZN(n19268) );
  NAND2_X1 U20961 ( .A1(n19265), .A2(n19264), .ZN(n19267) );
  NAND3_X1 U20962 ( .A1(n19531), .A2(n19530), .A3(n19270), .ZN(n19271) );
  INV_X1 U20963 ( .A(n19565), .ZN(n19569) );
  NAND2_X1 U20964 ( .A1(n20400), .A2(n20414), .ZN(n19293) );
  NOR2_X1 U20965 ( .A1(n19278), .A2(n19277), .ZN(n19541) );
  NAND2_X1 U20966 ( .A1(n20417), .A2(n20415), .ZN(n19288) );
  INV_X1 U20967 ( .A(n19523), .ZN(n19279) );
  OAI21_X1 U20968 ( .B1(n19282), .B2(n19281), .A(n19521), .ZN(n19287) );
  NAND3_X1 U20969 ( .A1(n19283), .A2(n19518), .A3(n18895), .ZN(n19286) );
  NAND3_X1 U20970 ( .A1(n19526), .A2(n19284), .A3(n19520), .ZN(n19285) );
  MUX2_X1 U20971 ( .A(n3284), .B(n19560), .S(n19556), .Z(n19289) );
  MUX2_X1 U20973 ( .A(n24457), .B(n18927), .S(n19296), .Z(n19299) );
  NOR2_X1 U20974 ( .A1(n19300), .A2(n19296), .ZN(n19298) );
  AOI21_X1 U20975 ( .B1(n19304), .B2(n19303), .A(n24441), .ZN(n19305) );
  NAND3_X1 U20976 ( .A1(n19313), .A2(n264), .A3(n19312), .ZN(n19314) );
  NAND2_X1 U20977 ( .A1(n19315), .A2(n5371), .ZN(n19316) );
  NAND3_X1 U20978 ( .A1(n19318), .A2(n19317), .A3(n19316), .ZN(n19319) );
  NAND2_X1 U20979 ( .A1(n19320), .A2(n19319), .ZN(n20241) );
  INV_X1 U20981 ( .A(n19936), .ZN(n20244) );
  NOR2_X1 U20982 ( .A1(n19329), .A2(n19328), .ZN(n19330) );
  INV_X1 U20983 ( .A(n19937), .ZN(n20243) );
  INV_X1 U20984 ( .A(n19499), .ZN(n19496) );
  OAI21_X1 U20985 ( .B1(n19500), .B2(n357), .A(n19501), .ZN(n19337) );
  NOR2_X1 U20986 ( .A1(n19502), .A2(n19497), .ZN(n19336) );
  NAND3_X1 U20988 ( .A1(n19936), .A2(n20242), .A3(n19939), .ZN(n19339) );
  XNOR2_X1 U20989 ( .A(n21106), .B(n2735), .ZN(n19340) );
  XNOR2_X1 U20990 ( .A(n21121), .B(n19340), .ZN(n19341) );
  NAND2_X1 U20991 ( .A1(n25474), .A2(n19346), .ZN(n20389) );
  NAND2_X1 U20992 ( .A1(n20389), .A2(n20388), .ZN(n19347) );
  OAI21_X1 U20993 ( .B1(n19348), .B2(n20388), .A(n19347), .ZN(n19350) );
  NAND2_X1 U20994 ( .A1(n19349), .A2(n352), .ZN(n20390) );
  NAND2_X1 U20997 ( .A1(n19357), .A2(n19353), .ZN(n19448) );
  INV_X1 U20998 ( .A(n19448), .ZN(n19354) );
  NAND2_X1 U20999 ( .A1(n19354), .A2(n19452), .ZN(n19355) );
  NOR2_X1 U21002 ( .A1(n19364), .A2(n2216), .ZN(n19369) );
  NOR2_X1 U21003 ( .A1(n19366), .A2(n24968), .ZN(n19368) );
  AOI22_X1 U21004 ( .A1(n19376), .A2(n19369), .B1(n19368), .B2(n19367), .ZN(
        n19374) );
  NOR2_X1 U21005 ( .A1(n19371), .A2(n24361), .ZN(n19372) );
  AND3_X1 U21006 ( .A1(n19382), .A2(n19381), .A3(n19380), .ZN(n19383) );
  NAND2_X1 U21007 ( .A1(n19384), .A2(n19389), .ZN(n19385) );
  XNOR2_X1 U21008 ( .A(n1326), .B(n19392), .ZN(n19443) );
  NOR2_X1 U21009 ( .A1(n19396), .A2(n24407), .ZN(n19398) );
  OAI21_X1 U21010 ( .B1(n19402), .B2(n1711), .A(n19719), .ZN(n19405) );
  NAND2_X1 U21011 ( .A1(n19406), .A2(n19412), .ZN(n19410) );
  MUX2_X1 U21012 ( .A(n19410), .B(n19409), .S(n19408), .Z(n19416) );
  NOR2_X1 U21013 ( .A1(n19412), .A2(n19411), .ZN(n19414) );
  OAI21_X1 U21014 ( .B1(n24584), .B2(n19418), .A(n19417), .ZN(n19422) );
  INV_X1 U21015 ( .A(n19761), .ZN(n19431) );
  AOI21_X1 U21016 ( .B1(n19428), .B2(n19760), .A(n19427), .ZN(n19429) );
  OAI21_X1 U21017 ( .B1(n24758), .B2(n19760), .A(n19429), .ZN(n19430) );
  NAND2_X1 U21018 ( .A1(n19431), .A2(n19430), .ZN(n19432) );
  MUX2_X1 U21019 ( .A(n20174), .B(n20586), .S(n19432), .Z(n19442) );
  OAI21_X1 U21020 ( .B1(n19435), .B2(n25423), .A(n19433), .ZN(n19440) );
  XNOR2_X1 U21021 ( .A(n19443), .B(n21505), .ZN(n19514) );
  NAND2_X1 U21029 ( .A1(n19459), .A2(n19464), .ZN(n19461) );
  MUX2_X1 U21030 ( .A(n19462), .B(n19461), .S(n19460), .Z(n19463) );
  NAND2_X1 U21032 ( .A1(n19468), .A2(n19471), .ZN(n19475) );
  OAI21_X1 U21033 ( .B1(n17872), .B2(n19470), .A(n19469), .ZN(n19473) );
  NAND2_X1 U21034 ( .A1(n19473), .A2(n19472), .ZN(n19474) );
  AND2_X2 U21035 ( .A1(n19475), .A2(n19474), .ZN(n20173) );
  MUX2_X1 U21036 ( .A(n20169), .B(n20235), .S(n20173), .Z(n19484) );
  NOR2_X1 U21039 ( .A1(n19484), .A2(n20168), .ZN(n19509) );
  OAI21_X1 U21040 ( .B1(n19490), .B2(n240), .A(n20388), .ZN(n19486) );
  NAND3_X1 U21042 ( .A1(n19490), .A2(n19345), .A3(n19488), .ZN(n19491) );
  OAI211_X1 U21043 ( .C1(n19500), .C2(n19497), .A(n19496), .B(n19495), .ZN(
        n19506) );
  NAND3_X1 U21044 ( .A1(n19500), .A2(n19499), .A3(n25459), .ZN(n19505) );
  NOR2_X1 U21045 ( .A1(n19502), .A2(n19501), .ZN(n19503) );
  NOR2_X1 U21046 ( .A1(n19494), .A2(n19777), .ZN(n19507) );
  INV_X1 U21049 ( .A(n19939), .ZN(n19788) );
  INV_X1 U21050 ( .A(n20242), .ZN(n19513) );
  OAI21_X1 U21051 ( .B1(n19939), .B2(n19936), .A(n19937), .ZN(n19511) );
  OAI21_X1 U21052 ( .B1(n19819), .B2(n19513), .A(n19512), .ZN(n21616) );
  XNOR2_X1 U21053 ( .A(n21659), .B(n21616), .ZN(n20285) );
  XNOR2_X1 U21054 ( .A(n20285), .B(n19514), .ZN(n19624) );
  OR2_X1 U21055 ( .A1(n21068), .A2(n19986), .ZN(n19988) );
  MUX2_X1 U21056 ( .A(n19987), .B(n19785), .S(n19986), .Z(n19516) );
  INV_X1 U21057 ( .A(n19983), .ZN(n19751) );
  NAND2_X1 U21058 ( .A1(n19986), .A2(n19751), .ZN(n19515) );
  INV_X1 U21059 ( .A(n19520), .ZN(n19521) );
  AOI22_X1 U21062 ( .A1(n19532), .A2(n19531), .B1(n19530), .B2(n19529), .ZN(
        n19538) );
  AOI21_X1 U21063 ( .B1(n19535), .B2(n5480), .A(n19533), .ZN(n19536) );
  INV_X1 U21064 ( .A(n24454), .ZN(n19962) );
  MUX2_X1 U21065 ( .A(n19540), .B(n3773), .S(n19539), .Z(n19545) );
  AOI21_X1 U21067 ( .B1(n25057), .B2(n19547), .A(n19546), .ZN(n19553) );
  OAI21_X1 U21069 ( .B1(n19553), .B2(n19552), .A(n19551), .ZN(n20373) );
  MUX2_X1 U21070 ( .A(n19962), .B(n20368), .S(n20369), .Z(n19574) );
  NAND2_X1 U21071 ( .A1(n19554), .A2(n4262), .ZN(n19564) );
  INV_X1 U21072 ( .A(n19555), .ZN(n19557) );
  NOR2_X1 U21073 ( .A1(n19557), .A2(n24421), .ZN(n19563) );
  NAND3_X1 U21074 ( .A1(n19560), .A2(n19559), .A3(n19558), .ZN(n19561) );
  NOR2_X1 U21075 ( .A1(n20370), .A2(n24558), .ZN(n19573) );
  NOR2_X1 U21076 ( .A1(n19569), .A2(n1053), .ZN(n19571) );
  NOR2_X1 U21077 ( .A1(n20368), .A2(n3428), .ZN(n19572) );
  INV_X1 U21078 ( .A(n20961), .ZN(n20450) );
  AOI21_X1 U21079 ( .B1(n19581), .B2(n19580), .A(n19198), .ZN(n19583) );
  MUX2_X1 U21080 ( .A(n19584), .B(n19583), .S(n19582), .Z(n19585) );
  INV_X1 U21081 ( .A(n20451), .ZN(n19942) );
  NAND3_X1 U21082 ( .A1(n19587), .A2(n24483), .A3(n19591), .ZN(n19588) );
  NOR2_X1 U21083 ( .A1(n25001), .A2(n24079), .ZN(n19600) );
  NOR2_X1 U21084 ( .A1(n19597), .A2(n19596), .ZN(n19599) );
  NAND2_X1 U21085 ( .A1(n20960), .A2(n19942), .ZN(n19605) );
  OAI211_X1 U21086 ( .C1(n20450), .C2(n19942), .A(n20377), .B(n19605), .ZN(
        n19621) );
  NOR2_X1 U21087 ( .A1(n19608), .A2(n2644), .ZN(n19609) );
  INV_X1 U21088 ( .A(n19612), .ZN(n19619) );
  NOR2_X1 U21089 ( .A1(n19613), .A2(n19615), .ZN(n19618) );
  OAI21_X1 U21090 ( .B1(n19616), .B2(n19615), .A(n19614), .ZN(n19617) );
  NOR2_X1 U21091 ( .A1(n20377), .A2(n20448), .ZN(n19620) );
  AOI22_X1 U21092 ( .A1(n20158), .A2(n20960), .B1(n19620), .B2(n20451), .ZN(
        n20962) );
  NAND2_X1 U21093 ( .A1(n19621), .A2(n20962), .ZN(n19622) );
  XNOR2_X1 U21094 ( .A(n24305), .B(n19622), .ZN(n20723) );
  XNOR2_X1 U21095 ( .A(n24898), .B(n20723), .ZN(n19623) );
  INV_X1 U21098 ( .A(n19629), .ZN(n19632) );
  OAI21_X1 U21099 ( .B1(n19632), .B2(n19631), .A(n19630), .ZN(n19633) );
  INV_X1 U21100 ( .A(n19636), .ZN(n19634) );
  MUX2_X1 U21101 ( .A(n19634), .B(n20484), .S(n20359), .Z(n19639) );
  NAND2_X1 U21104 ( .A1(n20482), .A2(n19636), .ZN(n19637) );
  NOR2_X1 U21106 ( .A1(n25088), .A2(n19928), .ZN(n19640) );
  INV_X1 U21111 ( .A(n20343), .ZN(n19645) );
  NOR2_X1 U21113 ( .A1(n20281), .A2(n1733), .ZN(n19646) );
  NAND3_X1 U21114 ( .A1(n20345), .A2(n20281), .A3(n20279), .ZN(n19647) );
  NAND4_X2 U21115 ( .A1(n19650), .A2(n19649), .A3(n19648), .A4(n19647), .ZN(
        n21193) );
  XNOR2_X1 U21116 ( .A(n21193), .B(n25265), .ZN(n21715) );
  XNOR2_X1 U21117 ( .A(n21715), .B(n20831), .ZN(n19667) );
  NOR2_X1 U21118 ( .A1(n24567), .A2(n20338), .ZN(n19653) );
  NOR2_X1 U21119 ( .A1(n20669), .A2(n20668), .ZN(n19652) );
  MUX2_X1 U21120 ( .A(n19653), .B(n19652), .S(n20666), .Z(n19656) );
  NOR2_X1 U21121 ( .A1(n20669), .A2(n20336), .ZN(n20349) );
  AND2_X1 U21122 ( .A1(n20666), .A2(n20336), .ZN(n19654) );
  XNOR2_X1 U21125 ( .A(n21306), .B(n24916), .ZN(n19665) );
  INV_X1 U21126 ( .A(n20183), .ZN(n20186) );
  INV_X1 U21127 ( .A(n20181), .ZN(n20038) );
  NAND3_X1 U21128 ( .A1(n20191), .A2(n20041), .A3(n20038), .ZN(n19663) );
  XNOR2_X1 U21129 ( .A(n21311), .B(n869), .ZN(n19664) );
  XNOR2_X1 U21130 ( .A(n19665), .B(n19664), .ZN(n19666) );
  XNOR2_X1 U21131 ( .A(n19667), .B(n19666), .ZN(n22688) );
  INV_X1 U21135 ( .A(n19675), .ZN(n19677) );
  OAI211_X1 U21136 ( .C1(n19675), .C2(n20124), .A(n20130), .B(n19674), .ZN(
        n19676) );
  XNOR2_X1 U21137 ( .A(n21649), .B(n21436), .ZN(n21253) );
  INV_X1 U21138 ( .A(n19991), .ZN(n20135) );
  OAI211_X1 U21139 ( .C1(n20135), .C2(n20014), .A(n1954), .B(n20019), .ZN(
        n19678) );
  XNOR2_X1 U21140 ( .A(n21336), .B(n2058), .ZN(n19679) );
  XNOR2_X1 U21141 ( .A(n21253), .B(n19679), .ZN(n19696) );
  INV_X1 U21142 ( .A(n20301), .ZN(n20008) );
  NAND2_X1 U21143 ( .A1(n20008), .A2(n19976), .ZN(n19682) );
  INV_X1 U21144 ( .A(n19680), .ZN(n19681) );
  INV_X1 U21145 ( .A(n19785), .ZN(n19980) );
  OAI211_X1 U21146 ( .C1(n19784), .C2(n19986), .A(n19984), .B(n19785), .ZN(
        n19683) );
  OAI21_X1 U21147 ( .B1(n19986), .B2(n19750), .A(n19683), .ZN(n19685) );
  NOR2_X1 U21148 ( .A1(n19684), .A2(n19987), .ZN(n21066) );
  XNOR2_X1 U21150 ( .A(n21332), .B(n21997), .ZN(n19694) );
  NAND2_X1 U21151 ( .A1(n20539), .A2(n20147), .ZN(n19690) );
  INV_X1 U21153 ( .A(n20145), .ZN(n19686) );
  NAND2_X1 U21154 ( .A1(n20145), .A2(n20149), .ZN(n20534) );
  NAND2_X1 U21155 ( .A1(n19691), .A2(n19714), .ZN(n19693) );
  XNOR2_X1 U21156 ( .A(n21729), .B(n21582), .ZN(n21200) );
  XNOR2_X1 U21157 ( .A(n19694), .B(n21200), .ZN(n19695) );
  XNOR2_X1 U21158 ( .A(n19696), .B(n19695), .ZN(n22685) );
  OR2_X1 U21159 ( .A1(n22688), .A2(n22685), .ZN(n22352) );
  MUX2_X1 U21160 ( .A(n19896), .B(n21033), .S(n19155), .Z(n19699) );
  NOR2_X1 U21162 ( .A1(n19700), .A2(n19880), .ZN(n19702) );
  MUX2_X1 U21163 ( .A(n3480), .B(n20554), .S(n20328), .Z(n19701) );
  MUX2_X2 U21164 ( .A(n19702), .B(n19701), .S(n20555), .Z(n21258) );
  XNOR2_X1 U21165 ( .A(n21300), .B(n21258), .ZN(n19713) );
  MUX2_X1 U21166 ( .A(n20616), .B(n20571), .S(n20618), .Z(n19706) );
  NAND3_X1 U21167 ( .A1(n19704), .A2(n20614), .A3(n19703), .ZN(n19705) );
  INV_X1 U21168 ( .A(n20669), .ZN(n20337) );
  NAND2_X1 U21169 ( .A1(n20337), .A2(n20668), .ZN(n19707) );
  OAI22_X1 U21170 ( .A1(n19710), .A2(n19709), .B1(n20337), .B2(n20670), .ZN(
        n19711) );
  XNOR2_X1 U21171 ( .A(n21745), .B(n21975), .ZN(n21208) );
  XNOR2_X1 U21172 ( .A(n21208), .B(n19713), .ZN(n19738) );
  INV_X1 U21173 ( .A(n21506), .ZN(n21979) );
  INV_X1 U21174 ( .A(n20111), .ZN(n20118) );
  XNOR2_X1 U21177 ( .A(n21297), .B(n21979), .ZN(n19736) );
  INV_X1 U21178 ( .A(n19719), .ZN(n19722) );
  INV_X1 U21179 ( .A(n19725), .ZN(n19721) );
  AOI21_X1 U21180 ( .B1(n19722), .B2(n19721), .A(n19720), .ZN(n19724) );
  OAI211_X1 U21181 ( .C1(n19726), .C2(n19725), .A(n19724), .B(n19723), .ZN(
        n19728) );
  INV_X1 U21182 ( .A(n19729), .ZN(n19733) );
  INV_X1 U21183 ( .A(n19730), .ZN(n19731) );
  NAND2_X1 U21184 ( .A1(n19733), .A2(n19732), .ZN(n19734) );
  XNOR2_X1 U21185 ( .A(n24491), .B(n2033), .ZN(n19735) );
  XNOR2_X1 U21186 ( .A(n19736), .B(n19735), .ZN(n19737) );
  INV_X1 U21187 ( .A(n21848), .ZN(n21289) );
  NAND2_X1 U21188 ( .A1(n22352), .A2(n21289), .ZN(n19836) );
  INV_X1 U21189 ( .A(n20419), .ZN(n20204) );
  NAND3_X1 U21190 ( .A1(n20422), .A2(n20400), .A3(n5590), .ZN(n19739) );
  INV_X1 U21192 ( .A(n20426), .ZN(n20598) );
  NAND2_X1 U21193 ( .A1(n20427), .A2(n20598), .ZN(n19846) );
  INV_X1 U21194 ( .A(n25442), .ZN(n19749) );
  OAI21_X1 U21195 ( .B1(n20263), .B2(n20262), .A(n20410), .ZN(n19742) );
  NOR2_X1 U21196 ( .A1(n20193), .A2(n20192), .ZN(n19745) );
  NAND2_X1 U21197 ( .A1(n20437), .A2(n19745), .ZN(n19747) );
  NOR2_X1 U21198 ( .A1(n20193), .A2(n20576), .ZN(n20195) );
  NAND2_X1 U21199 ( .A1(n20195), .A2(n24940), .ZN(n19746) );
  XNOR2_X1 U21200 ( .A(n19749), .B(n19748), .ZN(n19769) );
  INV_X1 U21201 ( .A(n19750), .ZN(n21065) );
  NAND2_X1 U21202 ( .A1(n21065), .A2(n25579), .ZN(n19754) );
  OAI21_X1 U21203 ( .B1(n19984), .B2(n19785), .A(n19751), .ZN(n19752) );
  NAND3_X1 U21205 ( .A1(n19754), .A2(n19753), .A3(n21067), .ZN(n21132) );
  NOR2_X1 U21206 ( .A1(n25242), .A2(n20134), .ZN(n19759) );
  XNOR2_X1 U21207 ( .A(n21132), .B(n21245), .ZN(n21328) );
  INV_X1 U21210 ( .A(n20593), .ZN(n20176) );
  OAI21_X1 U21211 ( .B1(n20590), .B2(n20586), .A(n20176), .ZN(n19764) );
  NAND3_X1 U21212 ( .A1(n20589), .A2(n20176), .A3(n3734), .ZN(n19765) );
  OAI211_X2 U21213 ( .C1(n19952), .C2(n20591), .A(n19766), .B(n19765), .ZN(
        n21720) );
  XNOR2_X1 U21214 ( .A(n21720), .B(n450), .ZN(n19767) );
  XNOR2_X1 U21215 ( .A(n21328), .B(n19767), .ZN(n19768) );
  AND2_X1 U21217 ( .A1(n22685), .A2(n21816), .ZN(n22349) );
  INV_X1 U21218 ( .A(n22688), .ZN(n22686) );
  NAND3_X1 U21219 ( .A1(n2688), .A2(n20448), .A3(n20377), .ZN(n19773) );
  XNOR2_X1 U21221 ( .A(n21750), .B(n21608), .ZN(n20708) );
  AND2_X1 U21222 ( .A1(n24461), .A2(n20384), .ZN(n20385) );
  NAND2_X1 U21224 ( .A1(n20459), .A2(n20384), .ZN(n19776) );
  NAND3_X1 U21225 ( .A1(n20234), .A2(n20231), .A3(n25205), .ZN(n19780) );
  OAI21_X1 U21226 ( .B1(n20169), .B2(n20236), .A(n20168), .ZN(n19779) );
  NOR2_X1 U21227 ( .A1(n20173), .A2(n20236), .ZN(n19778) );
  AOI22_X1 U21228 ( .A1(n19780), .A2(n19779), .B1(n20235), .B2(n19778), .ZN(
        n21042) );
  XNOR2_X1 U21229 ( .A(n21267), .B(n21042), .ZN(n21345) );
  XNOR2_X1 U21230 ( .A(n20708), .B(n21345), .ZN(n19796) );
  OAI21_X1 U21231 ( .B1(n20589), .B2(n20590), .A(n20586), .ZN(n19782) );
  NOR2_X1 U21232 ( .A1(n20587), .A2(n20588), .ZN(n19781) );
  AOI22_X2 U21233 ( .A1(n19783), .A2(n19782), .B1(n20174), .B2(n19781), .ZN(
        n21227) );
  INV_X1 U21234 ( .A(n21227), .ZN(n21588) );
  OAI21_X1 U21235 ( .B1(n19785), .B2(n19784), .A(n19984), .ZN(n19787) );
  XNOR2_X1 U21236 ( .A(n21588), .B(n21231), .ZN(n19794) );
  NAND2_X1 U21238 ( .A1(n19788), .A2(n1344), .ZN(n19791) );
  OAI211_X1 U21240 ( .C1(n20243), .C2(n20248), .A(n19789), .B(n19821), .ZN(
        n19790) );
  XNOR2_X1 U21241 ( .A(n21141), .B(n2042), .ZN(n19793) );
  XNOR2_X1 U21242 ( .A(n19794), .B(n19793), .ZN(n19795) );
  INV_X1 U21243 ( .A(n22689), .ZN(n21817) );
  NAND3_X1 U21244 ( .A1(n22686), .A2(n21816), .A3(n21817), .ZN(n19835) );
  AND2_X1 U21245 ( .A1(n3519), .A2(n19924), .ZN(n19798) );
  NAND2_X1 U21247 ( .A1(n20169), .A2(n20231), .ZN(n19802) );
  AOI21_X1 U21248 ( .B1(n19803), .B2(n19802), .A(n20239), .ZN(n19808) );
  NAND2_X1 U21249 ( .A1(n20173), .A2(n20236), .ZN(n19806) );
  INV_X1 U21250 ( .A(n20231), .ZN(n19804) );
  NAND2_X1 U21254 ( .A1(n19809), .A2(n20281), .ZN(n19812) );
  MUX2_X1 U21255 ( .A(n20281), .B(n20343), .S(n20345), .Z(n19810) );
  MUX2_X1 U21256 ( .A(n19810), .B(n1484), .S(n20279), .Z(n19811) );
  OAI21_X1 U21257 ( .B1(n19645), .B2(n19812), .A(n19811), .ZN(n21971) );
  INV_X1 U21258 ( .A(n21971), .ZN(n19813) );
  XNOR2_X1 U21259 ( .A(n21430), .B(n19813), .ZN(n19833) );
  NOR2_X1 U21260 ( .A1(n20507), .A2(n20214), .ZN(n20218) );
  NOR2_X1 U21262 ( .A1(n25224), .A2(n100), .ZN(n19814) );
  OAI21_X2 U21264 ( .B1(n19816), .B2(n20199), .A(n19815), .ZN(n21735) );
  INV_X1 U21265 ( .A(n19817), .ZN(n19820) );
  OAI211_X1 U21266 ( .C1(n20244), .C2(n20242), .A(n24077), .B(n19821), .ZN(
        n19822) );
  XNOR2_X1 U21267 ( .A(n21319), .B(n2228), .ZN(n19823) );
  XNOR2_X1 U21268 ( .A(n19823), .B(n21735), .ZN(n19831) );
  INV_X1 U21269 ( .A(n20268), .ZN(n20496) );
  NAND2_X1 U21270 ( .A1(n20501), .A2(n20496), .ZN(n19827) );
  NAND3_X1 U21272 ( .A1(n20411), .A2(n25420), .A3(n20410), .ZN(n19829) );
  XNOR2_X1 U21273 ( .A(n21561), .B(n21738), .ZN(n21224) );
  INV_X1 U21274 ( .A(n21224), .ZN(n19830) );
  XNOR2_X1 U21275 ( .A(n19830), .B(n19831), .ZN(n19832) );
  NOR2_X1 U21276 ( .A1(n21847), .A2(n21816), .ZN(n22690) );
  NAND2_X1 U21277 ( .A1(n22690), .A2(n21848), .ZN(n19834) );
  OAI211_X2 U21278 ( .C1(n19836), .C2(n22349), .A(n19835), .B(n19834), .ZN(
        n23865) );
  NOR2_X1 U21281 ( .A1(n5208), .A2(n20576), .ZN(n19838) );
  NAND3_X1 U21282 ( .A1(n19843), .A2(n19842), .A3(n19841), .ZN(n19844) );
  XNOR2_X1 U21283 ( .A(n20804), .B(n21974), .ZN(n20722) );
  NOR2_X1 U21284 ( .A1(n20597), .A2(n20427), .ZN(n20602) );
  INV_X1 U21285 ( .A(n20427), .ZN(n20595) );
  NAND2_X1 U21286 ( .A1(n20595), .A2(n20599), .ZN(n19845) );
  NAND2_X1 U21287 ( .A1(n19846), .A2(n19845), .ZN(n19847) );
  XNOR2_X1 U21288 ( .A(n21660), .B(n21616), .ZN(n21003) );
  XNOR2_X1 U21289 ( .A(n21003), .B(n20722), .ZN(n19870) );
  INV_X1 U21290 ( .A(n20071), .ZN(n20074) );
  NOR2_X1 U21292 ( .A1(n20415), .A2(n20400), .ZN(n20416) );
  NOR2_X1 U21293 ( .A1(n20416), .A2(n20414), .ZN(n19861) );
  INV_X1 U21294 ( .A(n20415), .ZN(n20399) );
  NOR2_X1 U21295 ( .A1(n20399), .A2(n20414), .ZN(n19856) );
  NAND2_X1 U21296 ( .A1(n19856), .A2(n1662), .ZN(n19859) );
  NAND2_X1 U21297 ( .A1(n19857), .A2(n4509), .ZN(n19858) );
  XNOR2_X1 U21299 ( .A(n21301), .B(n21136), .ZN(n19868) );
  NAND2_X1 U21300 ( .A1(n25212), .A2(n20039), .ZN(n19863) );
  NAND2_X1 U21301 ( .A1(n25212), .A2(n25478), .ZN(n20043) );
  MUX2_X1 U21302 ( .A(n19863), .B(n20043), .S(n20191), .Z(n19864) );
  XNOR2_X1 U21304 ( .A(n20964), .B(n2044), .ZN(n19867) );
  XNOR2_X1 U21305 ( .A(n19868), .B(n19867), .ZN(n19869) );
  OAI21_X1 U21307 ( .B1(n20572), .B2(n3795), .A(n20571), .ZN(n19874) );
  NAND2_X2 U21308 ( .A1(n19874), .A2(n19873), .ZN(n21399) );
  AOI21_X1 U21309 ( .B1(n20023), .B2(n20562), .A(n20094), .ZN(n19877) );
  XNOR2_X1 U21311 ( .A(n25040), .B(n21399), .ZN(n20816) );
  NAND2_X1 U21312 ( .A1(n20556), .A2(n20557), .ZN(n19879) );
  AND2_X1 U21313 ( .A1(n20091), .A2(n19879), .ZN(n19882) );
  OAI21_X1 U21314 ( .B1(n19880), .B2(n20330), .A(n20328), .ZN(n19881) );
  NAND2_X1 U21315 ( .A1(n19917), .A2(n25262), .ZN(n20114) );
  OAI22_X1 U21316 ( .A1(n25262), .A2(n19883), .B1(n20109), .B2(n19887), .ZN(
        n19884) );
  NAND2_X1 U21317 ( .A1(n19884), .A2(n20118), .ZN(n19886) );
  XNOR2_X1 U21318 ( .A(n21496), .B(n20816), .ZN(n19903) );
  INV_X1 U21322 ( .A(n20102), .ZN(n19895) );
  NAND2_X1 U21323 ( .A1(n19895), .A2(n19896), .ZN(n19913) );
  NAND2_X1 U21324 ( .A1(n20101), .A2(n20100), .ZN(n19894) );
  AOI21_X1 U21325 ( .B1(n19913), .B2(n19894), .A(n19893), .ZN(n19899) );
  NAND2_X1 U21326 ( .A1(n19895), .A2(n24378), .ZN(n19897) );
  AOI21_X1 U21327 ( .B1(n19897), .B2(n19896), .A(n20100), .ZN(n19898) );
  XNOR2_X1 U21328 ( .A(n20697), .B(n21621), .ZN(n19901) );
  XNOR2_X1 U21329 ( .A(n21247), .B(n2193), .ZN(n19900) );
  XNOR2_X1 U21330 ( .A(n19901), .B(n19900), .ZN(n19902) );
  XNOR2_X1 U21331 ( .A(n19903), .B(n19902), .ZN(n22227) );
  INV_X1 U21332 ( .A(n22227), .ZN(n21791) );
  INV_X1 U21333 ( .A(n20501), .ZN(n20226) );
  NOR2_X1 U21334 ( .A1(n20502), .A2(n20225), .ZN(n19907) );
  NOR2_X1 U21335 ( .A1(n343), .A2(n20497), .ZN(n19906) );
  OAI211_X1 U21336 ( .C1(n19904), .C2(n20269), .A(n20226), .B(n24887), .ZN(
        n19905) );
  OAI21_X1 U21337 ( .B1(n19907), .B2(n19906), .A(n19905), .ZN(n21510) );
  NAND2_X1 U21338 ( .A1(n2024), .A2(n345), .ZN(n19909) );
  NAND2_X1 U21339 ( .A1(n19909), .A2(n19910), .ZN(n19912) );
  XNOR2_X1 U21340 ( .A(n21510), .B(n20778), .ZN(n21108) );
  MUX2_X1 U21341 ( .A(n21033), .B(n19913), .S(n21038), .Z(n19914) );
  OAI21_X1 U21342 ( .B1(n19915), .B2(n20099), .A(n19914), .ZN(n21331) );
  OAI21_X1 U21343 ( .B1(n25034), .B2(n20118), .A(n25388), .ZN(n19918) );
  NAND3_X1 U21345 ( .A1(n20117), .A2(n20118), .A3(n25514), .ZN(n19920) );
  XNOR2_X1 U21346 ( .A(n21331), .B(n21647), .ZN(n20568) );
  XNOR2_X1 U21347 ( .A(n21108), .B(n20568), .ZN(n19935) );
  NAND2_X1 U21348 ( .A1(n351), .A2(n20517), .ZN(n19923) );
  NAND2_X1 U21349 ( .A1(n20516), .A2(n19924), .ZN(n19922) );
  NAND2_X1 U21350 ( .A1(n19923), .A2(n19922), .ZN(n20222) );
  INV_X1 U21351 ( .A(n19924), .ZN(n20514) );
  NAND2_X1 U21352 ( .A1(n20276), .A2(n20514), .ZN(n20519) );
  OAI21_X1 U21353 ( .B1(n20272), .B2(n20517), .A(n19925), .ZN(n19926) );
  XNOR2_X1 U21355 ( .A(n20780), .B(n24986), .ZN(n19933) );
  NAND3_X1 U21356 ( .A1(n20468), .A2(n19928), .A3(n25490), .ZN(n19931) );
  NAND2_X1 U21358 ( .A1(n20470), .A2(n20473), .ZN(n19930) );
  NAND3_X1 U21359 ( .A1(n20062), .A2(n25088), .A3(n20055), .ZN(n19929) );
  XNOR2_X1 U21361 ( .A(n20999), .B(n23679), .ZN(n19932) );
  XNOR2_X1 U21362 ( .A(n19933), .B(n19932), .ZN(n19934) );
  INV_X1 U21363 ( .A(n22226), .ZN(n21836) );
  MUX2_X1 U21364 ( .A(n20243), .B(n19939), .S(n19936), .Z(n19941) );
  NOR2_X1 U21365 ( .A1(n19937), .A2(n20242), .ZN(n19938) );
  XNOR2_X1 U21366 ( .A(n25062), .B(n663), .ZN(n19946) );
  INV_X1 U21367 ( .A(n20448), .ZN(n20159) );
  AOI21_X1 U21368 ( .B1(n19948), .B2(n20383), .A(n20460), .ZN(n19947) );
  NAND2_X1 U21369 ( .A1(n20461), .A2(n1327), .ZN(n20163) );
  NAND2_X1 U21370 ( .A1(n19947), .A2(n20163), .ZN(n19950) );
  NAND3_X1 U21371 ( .A1(n20588), .A2(n20593), .A3(n20586), .ZN(n19954) );
  NAND2_X1 U21373 ( .A1(n25205), .A2(n20169), .ZN(n19956) );
  MUX2_X1 U21374 ( .A(n19956), .B(n20234), .S(n20235), .Z(n19961) );
  INV_X1 U21375 ( .A(n20169), .ZN(n20232) );
  NAND2_X1 U21377 ( .A1(n20173), .A2(n20231), .ZN(n19957) );
  OAI22_X1 U21378 ( .A1(n20235), .A2(n19958), .B1(n25205), .B2(n19957), .ZN(
        n19959) );
  INV_X1 U21379 ( .A(n19959), .ZN(n19960) );
  XNOR2_X1 U21380 ( .A(n20767), .B(n20948), .ZN(n19965) );
  NOR2_X1 U21381 ( .A1(n20374), .A2(n20370), .ZN(n19964) );
  XNOR2_X1 U21382 ( .A(n19965), .B(n21115), .ZN(n21642) );
  XNOR2_X1 U21383 ( .A(n19966), .B(n21642), .ZN(n20036) );
  NOR2_X1 U21384 ( .A1(n20312), .A2(n20546), .ZN(n19968) );
  NOR3_X1 U21386 ( .A1(n20126), .A2(n20124), .A3(n20309), .ZN(n19969) );
  NOR2_X2 U21387 ( .A1(n19970), .A2(n19969), .ZN(n21126) );
  OAI22_X1 U21389 ( .A1(n20289), .A2(n19971), .B1(n20131), .B2(n21010), .ZN(
        n19974) );
  XNOR2_X1 U21390 ( .A(n21534), .B(n21126), .ZN(n20812) );
  NAND2_X1 U21391 ( .A1(n20301), .A2(n19976), .ZN(n19977) );
  OAI21_X1 U21392 ( .B1(n19979), .B2(n20141), .A(n19978), .ZN(n21967) );
  XNOR2_X1 U21393 ( .A(n20812), .B(n21967), .ZN(n21083) );
  NOR2_X1 U21396 ( .A1(n19988), .A2(n24979), .ZN(n19989) );
  NOR2_X2 U21397 ( .A1(n19990), .A2(n19989), .ZN(n21318) );
  INV_X1 U21398 ( .A(n20016), .ZN(n19996) );
  OAI21_X1 U21399 ( .B1(n20134), .B2(n20019), .A(n25242), .ZN(n19995) );
  NOR2_X1 U21400 ( .A1(n19991), .A2(n20014), .ZN(n19992) );
  INV_X1 U21401 ( .A(n3158), .ZN(n23500) );
  XNOR2_X1 U21402 ( .A(n20914), .B(n23500), .ZN(n19997) );
  XNOR2_X1 U21403 ( .A(n19997), .B(n21318), .ZN(n20001) );
  NAND2_X1 U21404 ( .A1(n20447), .A2(n20147), .ZN(n20000) );
  NOR2_X1 U21405 ( .A1(n20536), .A2(n20445), .ZN(n20150) );
  NOR2_X1 U21406 ( .A1(n20537), .A2(n19018), .ZN(n19998) );
  AND2_X1 U21407 ( .A1(n20536), .A2(n20149), .ZN(n20148) );
  NAND2_X1 U21408 ( .A1(n20148), .A2(n19018), .ZN(n19999) );
  XNOR2_X1 U21409 ( .A(n20001), .B(n20984), .ZN(n20002) );
  AND2_X1 U21410 ( .A1(n20036), .A2(n24905), .ZN(n22232) );
  INV_X1 U21411 ( .A(n22232), .ZN(n21835) );
  AOI21_X1 U21412 ( .B1(n20478), .B2(n20003), .A(n2168), .ZN(n20004) );
  NOR2_X1 U21414 ( .A1(n20486), .A2(n24275), .ZN(n20005) );
  INV_X1 U21415 ( .A(n20484), .ZN(n20910) );
  AND2_X1 U21416 ( .A1(n20910), .A2(n20909), .ZN(n20080) );
  AOI21_X1 U21417 ( .B1(n20005), .B2(n20360), .A(n20080), .ZN(n20007) );
  NAND3_X1 U21418 ( .A1(n24078), .A2(n20486), .A3(n20911), .ZN(n20006) );
  NOR2_X1 U21419 ( .A1(n20298), .A2(n20142), .ZN(n20010) );
  OAI21_X1 U21420 ( .B1(n20010), .B2(n20009), .A(n20008), .ZN(n20013) );
  INV_X1 U21421 ( .A(n20141), .ZN(n20011) );
  NAND2_X1 U21423 ( .A1(n25242), .A2(n20014), .ZN(n20015) );
  NAND2_X1 U21425 ( .A1(n20135), .A2(n1954), .ZN(n20020) );
  INV_X1 U21426 ( .A(n1792), .ZN(n20021) );
  NAND2_X1 U21427 ( .A1(n275), .A2(n20022), .ZN(n20026) );
  NAND3_X1 U21428 ( .A1(n275), .A2(n20562), .A3(n20560), .ZN(n20024) );
  OAI211_X1 U21429 ( .C1(n25221), .C2(n20026), .A(n20025), .B(n20024), .ZN(
        n20798) );
  NOR2_X1 U21430 ( .A1(n20027), .A2(n3671), .ZN(n20031) );
  NOR2_X1 U21431 ( .A1(n20281), .A2(n19809), .ZN(n20029) );
  NOR2_X1 U21432 ( .A1(n19809), .A2(n1733), .ZN(n20028) );
  AOI22_X1 U21433 ( .A1(n19645), .A2(n20029), .B1(n20028), .B2(n20345), .ZN(
        n20030) );
  OAI21_X1 U21434 ( .B1(n20031), .B2(n20345), .A(n20030), .ZN(n21142) );
  XNOR2_X1 U21435 ( .A(n20798), .B(n21142), .ZN(n20032) );
  XNOR2_X1 U21436 ( .A(n20033), .B(n20032), .ZN(n20034) );
  XNOR2_X1 U21437 ( .A(n20035), .B(n20034), .ZN(n22225) );
  INV_X1 U21438 ( .A(n22225), .ZN(n22235) );
  OAI22_X1 U21439 ( .A1(n21835), .A2(n22228), .B1(n22235), .B2(n22233), .ZN(
        n20037) );
  NOR2_X1 U21440 ( .A1(n20040), .A2(n20042), .ZN(n20045) );
  INV_X1 U21441 ( .A(n20046), .ZN(n22697) );
  NOR2_X1 U21442 ( .A1(n20478), .A2(n20477), .ZN(n20048) );
  INV_X1 U21443 ( .A(n20476), .ZN(n20049) );
  NAND2_X1 U21444 ( .A1(n20353), .A2(n20049), .ZN(n20050) );
  AND3_X1 U21445 ( .A1(n20051), .A2(n20050), .A3(n20477), .ZN(n20052) );
  INV_X1 U21446 ( .A(n25490), .ZN(n20056) );
  OAI21_X1 U21447 ( .B1(n20056), .B2(n20472), .A(n5734), .ZN(n20058) );
  NAND2_X1 U21448 ( .A1(n20058), .A2(n5115), .ZN(n20065) );
  NOR2_X1 U21449 ( .A1(n20054), .A2(n25089), .ZN(n20063) );
  NOR2_X1 U21450 ( .A1(n20060), .A2(n20473), .ZN(n20061) );
  AOI22_X1 U21451 ( .A1(n20063), .A2(n20062), .B1(n20061), .B2(n20470), .ZN(
        n20064) );
  NAND2_X1 U21452 ( .A1(n20065), .A2(n20064), .ZN(n21222) );
  XNOR2_X1 U21453 ( .A(n21704), .B(n21222), .ZN(n20628) );
  OAI21_X1 U21454 ( .B1(n20909), .B2(n20359), .A(n347), .ZN(n20079) );
  NOR2_X1 U21455 ( .A1(n20076), .A2(n347), .ZN(n20078) );
  NOR2_X1 U21456 ( .A1(n20483), .A2(n20486), .ZN(n20077) );
  OAI21_X1 U21458 ( .B1(n20080), .B2(n20079), .A(n20912), .ZN(n20626) );
  XNOR2_X1 U21459 ( .A(n25483), .B(n20626), .ZN(n20081) );
  XNOR2_X1 U21460 ( .A(n21971), .B(n20081), .ZN(n20082) );
  NOR3_X1 U21461 ( .A1(n20616), .A2(n20615), .A3(n20614), .ZN(n20086) );
  AOI21_X1 U21462 ( .B1(n20572), .B2(n20617), .A(n20086), .ZN(n20087) );
  XNOR2_X1 U21463 ( .A(n21521), .B(n21676), .ZN(n21114) );
  INV_X1 U21464 ( .A(n20557), .ZN(n20092) );
  INV_X1 U21466 ( .A(n25221), .ZN(n20566) );
  XNOR2_X1 U21468 ( .A(n21192), .B(n21114), .ZN(n20123) );
  NAND2_X1 U21471 ( .A1(n20104), .A2(n20103), .ZN(n21034) );
  MUX2_X1 U21472 ( .A(n20105), .B(n21034), .S(n21038), .Z(n20106) );
  XNOR2_X1 U21473 ( .A(n21469), .B(n21679), .ZN(n20121) );
  NAND2_X1 U21474 ( .A1(n20111), .A2(n25262), .ZN(n20112) );
  MUX2_X1 U21475 ( .A(n20113), .B(n20112), .S(n25034), .Z(n20119) );
  NAND2_X1 U21476 ( .A1(n339), .A2(n25388), .ZN(n20116) );
  XNOR2_X1 U21477 ( .A(n21601), .B(n2744), .ZN(n20120) );
  XNOR2_X1 U21478 ( .A(n20121), .B(n20120), .ZN(n20122) );
  AND2_X1 U21479 ( .A1(n20546), .A2(n20125), .ZN(n20308) );
  INV_X1 U21480 ( .A(n20308), .ZN(n20129) );
  NAND2_X1 U21481 ( .A1(n20545), .A2(n20127), .ZN(n20128) );
  XNOR2_X1 U21483 ( .A(n21665), .B(n22745), .ZN(n20133) );
  XNOR2_X1 U21484 ( .A(n21209), .B(n20133), .ZN(n20155) );
  MUX2_X1 U21485 ( .A(n20136), .B(n20135), .S(n25242), .Z(n20138) );
  MUX2_X2 U21486 ( .A(n20139), .B(n20138), .S(n20137), .Z(n21980) );
  INV_X1 U21487 ( .A(n20140), .ZN(n20299) );
  XNOR2_X1 U21488 ( .A(n21554), .B(n21980), .ZN(n21030) );
  OAI211_X1 U21489 ( .C1(n20533), .C2(n20447), .A(n20147), .B(n20146), .ZN(
        n20153) );
  NAND2_X1 U21490 ( .A1(n20148), .A2(n20537), .ZN(n20152) );
  NAND2_X1 U21491 ( .A1(n20150), .A2(n20149), .ZN(n20151) );
  XNOR2_X1 U21493 ( .A(n21506), .B(n21138), .ZN(n20898) );
  XNOR2_X1 U21494 ( .A(n21030), .B(n20898), .ZN(n20154) );
  XNOR2_X2 U21495 ( .A(n20155), .B(n20154), .ZN(n22356) );
  MUX2_X1 U21496 ( .A(n22355), .B(n22361), .S(n22356), .Z(n20254) );
  AND2_X1 U21497 ( .A1(n24454), .A2(n20369), .ZN(n20156) );
  NOR2_X1 U21498 ( .A1(n20451), .A2(n20159), .ZN(n20157) );
  INV_X1 U21499 ( .A(n20960), .ZN(n20455) );
  AOI22_X1 U21500 ( .A1(n20157), .A2(n20961), .B1(n20455), .B2(n20451), .ZN(
        n20162) );
  INV_X1 U21501 ( .A(n20158), .ZN(n20160) );
  NAND3_X1 U21502 ( .A1(n20160), .A2(n20159), .A3(n20377), .ZN(n20161) );
  XNOR2_X1 U21503 ( .A(n21577), .B(n1381), .ZN(n21199) );
  INV_X1 U21504 ( .A(n20163), .ZN(n20164) );
  OAI21_X1 U21505 ( .B1(n20395), .B2(n24460), .A(n20164), .ZN(n20167) );
  OAI21_X1 U21506 ( .B1(n20458), .B2(n24461), .A(n20165), .ZN(n20166) );
  AND2_X1 U21507 ( .A1(n20167), .A2(n20166), .ZN(n21578) );
  NOR2_X1 U21508 ( .A1(n20169), .A2(n20231), .ZN(n20237) );
  NAND2_X1 U21509 ( .A1(n20237), .A2(n20173), .ZN(n20172) );
  OAI211_X1 U21510 ( .C1(n20170), .C2(n20236), .A(n20169), .B(n20168), .ZN(
        n20171) );
  XNOR2_X1 U21511 ( .A(n21998), .B(n21578), .ZN(n21061) );
  XNOR2_X1 U21512 ( .A(n21061), .B(n21199), .ZN(n20180) );
  XNOR2_X1 U21513 ( .A(n21997), .B(n23151), .ZN(n20178) );
  NAND2_X1 U21514 ( .A1(n20174), .A2(n20588), .ZN(n20175) );
  NAND3_X1 U21515 ( .A1(n20175), .A2(n20590), .A3(n20586), .ZN(n20177) );
  XNOR2_X1 U21516 ( .A(n25386), .B(n21106), .ZN(n21671) );
  XNOR2_X1 U21517 ( .A(n21671), .B(n20178), .ZN(n20179) );
  XNOR2_X1 U21518 ( .A(n20179), .B(n20180), .ZN(n21838) );
  AOI21_X1 U21519 ( .B1(n20183), .B2(n25211), .A(n25478), .ZN(n20190) );
  OAI21_X1 U21520 ( .B1(n20188), .B2(n20187), .A(n20186), .ZN(n20189) );
  XNOR2_X1 U21521 ( .A(n22007), .B(n21689), .ZN(n21093) );
  NAND2_X1 U21522 ( .A1(n20195), .A2(n20194), .ZN(n20196) );
  XNOR2_X1 U21523 ( .A(n20197), .B(n21093), .ZN(n20213) );
  MUX2_X1 U21526 ( .A(n20200), .B(n20199), .S(n20215), .Z(n20201) );
  INV_X1 U21527 ( .A(n20203), .ZN(n20205) );
  AOI22_X1 U21528 ( .A1(n20205), .A2(n20399), .B1(n5733), .B2(n20204), .ZN(
        n20207) );
  NAND3_X1 U21529 ( .A1(n20415), .A2(n20401), .A3(n20400), .ZN(n20206) );
  NOR2_X1 U21530 ( .A1(n20595), .A2(n20599), .ZN(n20208) );
  OAI21_X1 U21531 ( .B1(n1667), .B2(n20426), .A(n20595), .ZN(n20211) );
  NOR2_X1 U21532 ( .A1(n1667), .A2(n25397), .ZN(n20210) );
  XNOR2_X1 U21533 ( .A(n20212), .B(n21445), .ZN(n20642) );
  MUX2_X1 U21535 ( .A(n21782), .B(n21839), .S(n22361), .Z(n20253) );
  AOI22_X1 U21536 ( .A1(n24327), .A2(n20215), .B1(n20216), .B2(n20214), .ZN(
        n20220) );
  OAI21_X1 U21538 ( .B1(n20276), .B2(n20514), .A(n20516), .ZN(n20221) );
  XNOR2_X1 U21539 ( .A(n21495), .B(n21568), .ZN(n21215) );
  OAI21_X1 U21540 ( .B1(n3016), .B2(n20226), .A(n20268), .ZN(n20227) );
  NAND2_X1 U21542 ( .A1(n20237), .A2(n20236), .ZN(n20238) );
  XNOR2_X1 U21543 ( .A(n21070), .B(n21694), .ZN(n20251) );
  NAND3_X1 U21544 ( .A1(n19936), .A2(n20242), .A3(n20241), .ZN(n20247) );
  XNOR2_X1 U21548 ( .A(n21087), .B(n673), .ZN(n20250) );
  XNOR2_X1 U21549 ( .A(n20251), .B(n20250), .ZN(n20252) );
  OR3_X1 U21550 ( .A1(n20255), .A2(n25420), .A3(n20411), .ZN(n20267) );
  NOR2_X1 U21551 ( .A1(n20256), .A2(n25420), .ZN(n20261) );
  NOR3_X1 U21552 ( .A1(n20259), .A2(n20258), .A3(n20257), .ZN(n20260) );
  NAND2_X1 U21553 ( .A1(n20261), .A2(n20260), .ZN(n20266) );
  NAND3_X1 U21554 ( .A1(n20411), .A2(n20262), .A3(n25421), .ZN(n20265) );
  XNOR2_X1 U21555 ( .A(n21172), .B(n20804), .ZN(n21409) );
  MUX2_X2 U21556 ( .A(n20271), .B(n20270), .S(n20497), .Z(n21501) );
  NAND2_X1 U21557 ( .A1(n20515), .A2(n20272), .ZN(n20273) );
  XNOR2_X1 U21558 ( .A(n21501), .B(n21658), .ZN(n21302) );
  XNOR2_X1 U21559 ( .A(n21409), .B(n21302), .ZN(n20288) );
  NOR2_X1 U21560 ( .A1(n20280), .A2(n20343), .ZN(n20282) );
  XNOR2_X1 U21562 ( .A(n20475), .B(n20284), .ZN(n20286) );
  XNOR2_X1 U21563 ( .A(n20285), .B(n20286), .ZN(n20287) );
  NAND2_X1 U21564 ( .A1(n20289), .A2(n21008), .ZN(n20293) );
  NAND2_X1 U21565 ( .A1(n20290), .A2(n20522), .ZN(n20292) );
  AOI21_X1 U21566 ( .B1(n20293), .B2(n20292), .A(n20291), .ZN(n20294) );
  OAI21_X1 U21568 ( .B1(n20298), .B2(n20297), .A(n20296), .ZN(n20300) );
  XNOR2_X1 U21569 ( .A(n25470), .B(n21985), .ZN(n20307) );
  NAND3_X1 U21570 ( .A1(n3428), .A2(n24558), .A3(n24454), .ZN(n20304) );
  XNOR2_X1 U21572 ( .A(n21569), .B(n5514), .ZN(n20306) );
  XNOR2_X1 U21573 ( .A(n20307), .B(n20306), .ZN(n20315) );
  XNOR2_X1 U21574 ( .A(n21399), .B(n25222), .ZN(n20313) );
  NOR2_X1 U21575 ( .A1(n20308), .A2(n20543), .ZN(n20311) );
  XNOR2_X1 U21576 ( .A(n21324), .B(n21247), .ZN(n20990) );
  XNOR2_X1 U21577 ( .A(n20313), .B(n20990), .ZN(n20314) );
  XNOR2_X1 U21579 ( .A(n21686), .B(n1757), .ZN(n20324) );
  INV_X1 U21583 ( .A(n20554), .ZN(n20333) );
  OAI21_X1 U21584 ( .B1(n20554), .B2(n20555), .A(n20330), .ZN(n20331) );
  NAND2_X1 U21585 ( .A1(n20670), .A2(n20335), .ZN(n20350) );
  NAND3_X1 U21586 ( .A1(n20338), .A2(n20337), .A3(n20336), .ZN(n20339) );
  OAI211_X1 U21587 ( .C1(n20350), .C2(n20341), .A(n20340), .B(n20339), .ZN(
        n21157) );
  XNOR2_X1 U21588 ( .A(n20798), .B(n21157), .ZN(n21420) );
  XNOR2_X1 U21589 ( .A(n21420), .B(n21343), .ZN(n20342) );
  NOR2_X1 U21590 ( .A1(n24414), .A2(n1733), .ZN(n20344) );
  OAI211_X1 U21592 ( .C1(n24414), .C2(n19809), .A(n20345), .B(n1733), .ZN(
        n20347) );
  XNOR2_X1 U21594 ( .A(n20780), .B(n21334), .ZN(n20358) );
  OAI21_X1 U21595 ( .B1(n20353), .B2(n20480), .A(n20352), .ZN(n20357) );
  XNOR2_X1 U21598 ( .A(n21058), .B(n21511), .ZN(n20889) );
  XNOR2_X1 U21599 ( .A(n20358), .B(n20889), .ZN(n20366) );
  OAI211_X1 U21600 ( .C1(n20360), .C2(n20491), .A(n20486), .B(n20359), .ZN(
        n20361) );
  XNOR2_X1 U21602 ( .A(n21996), .B(n21515), .ZN(n21668) );
  XNOR2_X1 U21603 ( .A(n20999), .B(n2757), .ZN(n20364) );
  XNOR2_X1 U21604 ( .A(n21668), .B(n20364), .ZN(n20365) );
  XNOR2_X1 U21605 ( .A(n20366), .B(n20365), .ZN(n22655) );
  NOR2_X1 U21606 ( .A1(n20368), .A2(n24558), .ZN(n20372) );
  NOR2_X2 U21607 ( .A1(n20376), .A2(n20375), .ZN(n21429) );
  OAI21_X1 U21609 ( .B1(n20377), .B2(n20451), .A(n20961), .ZN(n20381) );
  OAI21_X1 U21610 ( .B1(n2688), .B2(n20451), .A(n24357), .ZN(n20379) );
  OAI21_X1 U21611 ( .B1(n20961), .B2(n20448), .A(n20960), .ZN(n20378) );
  NAND2_X1 U21612 ( .A1(n20379), .A2(n20378), .ZN(n20380) );
  XNOR2_X1 U21613 ( .A(n21429), .B(n21633), .ZN(n21317) );
  NAND2_X1 U21614 ( .A1(n20385), .A2(n20459), .ZN(n20397) );
  AND2_X1 U21616 ( .A1(n20388), .A2(n20389), .ZN(n20391) );
  OAI21_X1 U21617 ( .B1(n20392), .B2(n20391), .A(n20390), .ZN(n20393) );
  XNOR2_X1 U21619 ( .A(n21965), .B(n21532), .ZN(n21701) );
  XNOR2_X1 U21620 ( .A(n25495), .B(n21701), .ZN(n20408) );
  MUX2_X1 U21621 ( .A(n20400), .B(n20399), .S(n20422), .Z(n20405) );
  NOR2_X1 U21622 ( .A1(n20415), .A2(n20414), .ZN(n20403) );
  AOI22_X1 U21623 ( .A1(n20403), .A2(n20422), .B1(n20402), .B2(n20419), .ZN(
        n20404) );
  XNOR2_X1 U21625 ( .A(n24353), .B(n2847), .ZN(n20406) );
  XNOR2_X1 U21626 ( .A(n20406), .B(n20984), .ZN(n20407) );
  XNOR2_X1 U21627 ( .A(n21600), .B(n891), .ZN(n20424) );
  NAND2_X1 U21628 ( .A1(n20415), .A2(n20414), .ZN(n20423) );
  NAND2_X1 U21629 ( .A1(n20416), .A2(n20419), .ZN(n20421) );
  XNOR2_X1 U21631 ( .A(n21310), .B(n24936), .ZN(n21415) );
  XNOR2_X1 U21632 ( .A(n21415), .B(n20424), .ZN(n20441) );
  NOR2_X1 U21633 ( .A1(n20427), .A2(n20599), .ZN(n20429) );
  AOI22_X1 U21634 ( .A1(n20597), .A2(n20430), .B1(n20429), .B2(n25397), .ZN(
        n20431) );
  NAND2_X1 U21635 ( .A1(n20432), .A2(n20577), .ZN(n20436) );
  OAI211_X1 U21636 ( .C1(n20438), .C2(n20437), .A(n20436), .B(n20435), .ZN(
        n22014) );
  XNOR2_X1 U21637 ( .A(n21308), .B(n20439), .ZN(n20440) );
  NAND2_X1 U21638 ( .A1(n25075), .A2(n22655), .ZN(n20442) );
  NAND2_X1 U21639 ( .A1(n20443), .A2(n22656), .ZN(n20444) );
  AOI21_X1 U21640 ( .B1(n20537), .B2(n20536), .A(n20445), .ZN(n20446) );
  XNOR2_X1 U21641 ( .A(n21721), .B(n25385), .ZN(n20457) );
  AOI21_X1 U21642 ( .B1(n24354), .B2(n20448), .A(n20450), .ZN(n20456) );
  XNOR2_X1 U21645 ( .A(n21246), .B(n20457), .ZN(n20467) );
  OAI211_X1 U21646 ( .C1(n20461), .C2(n1327), .A(n20460), .B(n20459), .ZN(
        n20463) );
  XNOR2_X1 U21647 ( .A(n21621), .B(n21693), .ZN(n21167) );
  INV_X1 U21648 ( .A(Key[60]), .ZN(n22089) );
  XNOR2_X1 U21649 ( .A(n21167), .B(n20465), .ZN(n20466) );
  XNOR2_X1 U21650 ( .A(n20466), .B(n20467), .ZN(n22770) );
  INV_X1 U21651 ( .A(n22770), .ZN(n22680) );
  NAND2_X1 U21652 ( .A1(n25490), .A2(n20472), .ZN(n20474) );
  XNOR2_X1 U21653 ( .A(n21173), .B(n20475), .ZN(n21551) );
  MUX2_X1 U21654 ( .A(n20477), .B(n20476), .S(n20479), .Z(n20481) );
  XNOR2_X1 U21655 ( .A(n21301), .B(n21040), .ZN(n21406) );
  XNOR2_X1 U21656 ( .A(n21551), .B(n21406), .ZN(n20495) );
  XNOR2_X1 U21657 ( .A(n21745), .B(n3129), .ZN(n20493) );
  NOR2_X1 U21659 ( .A1(n20484), .A2(n20491), .ZN(n20485) );
  INV_X1 U21661 ( .A(n20487), .ZN(n20488) );
  NAND2_X1 U21662 ( .A1(n20488), .A2(n20491), .ZN(n20489) );
  XNOR2_X1 U21663 ( .A(n21027), .B(n20964), .ZN(n21618) );
  XNOR2_X1 U21664 ( .A(n21618), .B(n20493), .ZN(n20494) );
  NOR2_X1 U21666 ( .A1(n3016), .A2(n20501), .ZN(n20499) );
  INV_X1 U21667 ( .A(n21193), .ZN(n20503) );
  XNOR2_X1 U21668 ( .A(n21414), .B(n20503), .ZN(n20505) );
  XNOR2_X1 U21669 ( .A(n21312), .B(n886), .ZN(n20504) );
  OAI22_X1 U21670 ( .A1(n20511), .A2(n20510), .B1(n24327), .B2(n20508), .ZN(
        n20512) );
  XNOR2_X1 U21671 ( .A(n21307), .B(n21675), .ZN(n20769) );
  XNOR2_X1 U21672 ( .A(n20769), .B(n20948), .ZN(n21156) );
  XNOR2_X2 U21673 ( .A(n20521), .B(n21156), .ZN(n22774) );
  MUX2_X1 U21674 ( .A(n22680), .B(n21856), .S(n22774), .Z(n20608) );
  INV_X1 U21675 ( .A(n20522), .ZN(n20525) );
  NAND2_X1 U21676 ( .A1(n20525), .A2(n20523), .ZN(n20527) );
  AOI21_X1 U21678 ( .B1(n20530), .B2(n24581), .A(n20528), .ZN(n20531) );
  NOR2_X1 U21679 ( .A1(n21013), .A2(n20531), .ZN(n21045) );
  OAI211_X1 U21680 ( .C1(n20533), .C2(n19018), .A(n20536), .B(n20532), .ZN(
        n20542) );
  INV_X1 U21681 ( .A(n20534), .ZN(n20535) );
  NAND2_X1 U21682 ( .A1(n20539), .A2(n20535), .ZN(n20541) );
  INV_X1 U21683 ( .A(n20536), .ZN(n20538) );
  NAND3_X1 U21684 ( .A1(n20539), .A2(n20538), .A3(n20537), .ZN(n20540) );
  XNOR2_X1 U21686 ( .A(n21422), .B(n21045), .ZN(n20762) );
  NAND2_X1 U21687 ( .A1(n20544), .A2(n20543), .ZN(n20547) );
  XNOR2_X1 U21688 ( .A(n24485), .B(n21158), .ZN(n21593) );
  XNOR2_X1 U21689 ( .A(n20762), .B(n21593), .ZN(n20553) );
  XNOR2_X1 U21690 ( .A(n21751), .B(n2145), .ZN(n20550) );
  XNOR2_X1 U21691 ( .A(n20551), .B(n20550), .ZN(n20552) );
  XNOR2_X1 U21692 ( .A(n20553), .B(n20552), .ZN(n22769) );
  INV_X1 U21693 ( .A(n22769), .ZN(n22369) );
  AND2_X1 U21694 ( .A1(n20556), .A2(n20555), .ZN(n20558) );
  AND2_X1 U21695 ( .A1(n20561), .A2(n20560), .ZN(n20565) );
  XNOR2_X1 U21696 ( .A(n21182), .B(n21579), .ZN(n20781) );
  XNOR2_X1 U21697 ( .A(n20781), .B(n20568), .ZN(n20575) );
  XNOR2_X1 U21698 ( .A(n21058), .B(n24100), .ZN(n21252) );
  XNOR2_X1 U21699 ( .A(n21729), .B(n2100), .ZN(n20573) );
  XNOR2_X1 U21700 ( .A(n21252), .B(n20573), .ZN(n20574) );
  NAND2_X1 U21702 ( .A1(n22369), .A2(n22679), .ZN(n20606) );
  NAND3_X1 U21703 ( .A1(n20577), .A2(n20576), .A3(n24940), .ZN(n20581) );
  NOR2_X1 U21704 ( .A1(n24940), .A2(n5208), .ZN(n20579) );
  NAND2_X1 U21705 ( .A1(n20583), .A2(n20579), .ZN(n20580) );
  XNOR2_X1 U21706 ( .A(n20914), .B(n21053), .ZN(n21635) );
  INV_X1 U21707 ( .A(n21738), .ZN(n21478) );
  XNOR2_X1 U21708 ( .A(n21478), .B(Key[149]), .ZN(n20584) );
  XNOR2_X1 U21709 ( .A(n21635), .B(n20584), .ZN(n20604) );
  INV_X1 U21710 ( .A(n20585), .ZN(n20594) );
  MUX2_X1 U21711 ( .A(n20588), .B(n20587), .S(n20586), .Z(n20592) );
  OAI21_X1 U21712 ( .B1(n276), .B2(n20595), .A(n20599), .ZN(n20601) );
  NOR3_X1 U21713 ( .A1(n24463), .A2(n20599), .A3(n20598), .ZN(n20600) );
  XNOR2_X1 U21714 ( .A(n21318), .B(n21734), .ZN(n21433) );
  XNOR2_X1 U21715 ( .A(n21562), .B(n21433), .ZN(n20603) );
  MUX2_X1 U21716 ( .A(n20606), .B(n20605), .S(n21856), .Z(n20607) );
  INV_X1 U21718 ( .A(n23859), .ZN(n23839) );
  INV_X1 U21719 ( .A(n20609), .ZN(n20625) );
  XNOR2_X1 U21720 ( .A(n21694), .B(n2795), .ZN(n20610) );
  XNOR2_X1 U21721 ( .A(n21215), .B(n20610), .ZN(n20613) );
  XNOR2_X1 U21722 ( .A(n24996), .B(n25073), .ZN(n20611) );
  XNOR2_X1 U21723 ( .A(n21132), .B(n21135), .ZN(n21725) );
  XNOR2_X1 U21724 ( .A(n20611), .B(n21725), .ZN(n20612) );
  XNOR2_X1 U21725 ( .A(n20612), .B(n20613), .ZN(n21908) );
  INV_X1 U21726 ( .A(n21908), .ZN(n22338) );
  XNOR2_X1 U21727 ( .A(n21319), .B(n21481), .ZN(n21739) );
  NAND2_X1 U21728 ( .A1(n20615), .A2(n20614), .ZN(n20622) );
  MUX2_X1 U21729 ( .A(n20617), .B(n20616), .S(n20615), .Z(n20620) );
  MUX2_X1 U21730 ( .A(n20620), .B(n20619), .S(n7), .Z(n20621) );
  XNOR2_X1 U21732 ( .A(n24353), .B(n21630), .ZN(n20624) );
  XNOR2_X1 U21733 ( .A(n21739), .B(n20624), .ZN(n20630) );
  XNOR2_X1 U21734 ( .A(n20626), .B(n20625), .ZN(n20627) );
  XNOR2_X1 U21735 ( .A(n20628), .B(n20627), .ZN(n20629) );
  XNOR2_X1 U21736 ( .A(n20630), .B(n20629), .ZN(n22137) );
  NOR2_X1 U21737 ( .A1(n22338), .A2(n22137), .ZN(n22336) );
  XNOR2_X1 U21738 ( .A(n21138), .B(n21743), .ZN(n21457) );
  XNOR2_X1 U21739 ( .A(n21505), .B(n876), .ZN(n20631) );
  XNOR2_X1 U21740 ( .A(n20631), .B(n21457), .ZN(n20633) );
  XNOR2_X1 U21741 ( .A(n21259), .B(n21300), .ZN(n20632) );
  XNOR2_X1 U21742 ( .A(n20633), .B(n20632), .ZN(n20635) );
  XNOR2_X1 U21744 ( .A(n21639), .B(n1920), .ZN(n20636) );
  XNOR2_X1 U21745 ( .A(n21192), .B(n20636), .ZN(n20639) );
  XNOR2_X1 U21746 ( .A(n21306), .B(n20870), .ZN(n21716) );
  XNOR2_X1 U21747 ( .A(n21676), .B(n21600), .ZN(n20637) );
  XNOR2_X1 U21748 ( .A(n20637), .B(n21716), .ZN(n20638) );
  AND2_X1 U21749 ( .A1(n22139), .A2(n22338), .ZN(n20649) );
  XNOR2_X1 U21750 ( .A(n20882), .B(n688), .ZN(n20640) );
  XNOR2_X1 U21751 ( .A(n20640), .B(n21541), .ZN(n20641) );
  XNOR2_X1 U21752 ( .A(n20826), .B(n21042), .ZN(n21755) );
  XNOR2_X1 U21753 ( .A(n20641), .B(n21755), .ZN(n20643) );
  XNOR2_X1 U21754 ( .A(n21336), .B(n21058), .ZN(n21584) );
  XNOR2_X1 U21755 ( .A(n21199), .B(n21584), .ZN(n20647) );
  XNOR2_X1 U21756 ( .A(n21514), .B(n21728), .ZN(n20645) );
  XNOR2_X1 U21757 ( .A(n25387), .B(n3073), .ZN(n20644) );
  XNOR2_X1 U21758 ( .A(n20645), .B(n20644), .ZN(n20646) );
  XNOR2_X1 U21759 ( .A(n20647), .B(n20646), .ZN(n22138) );
  AND2_X1 U21760 ( .A1(n22138), .A2(n22338), .ZN(n20648) );
  INV_X1 U21761 ( .A(n22139), .ZN(n22141) );
  NOR2_X1 U21762 ( .A1(n22338), .A2(n22139), .ZN(n20650) );
  XNOR2_X1 U21763 ( .A(n21414), .B(n21678), .ZN(n20651) );
  XNOR2_X1 U21764 ( .A(n21308), .B(n20651), .ZN(n20656) );
  XNOR2_X1 U21765 ( .A(n20948), .B(n21679), .ZN(n20654) );
  INV_X1 U21766 ( .A(n62), .ZN(n20652) );
  XNOR2_X1 U21767 ( .A(n24936), .B(n20652), .ZN(n20653) );
  XNOR2_X1 U21768 ( .A(n20654), .B(n20653), .ZN(n20655) );
  XNOR2_X1 U21770 ( .A(n21996), .B(n21511), .ZN(n21333) );
  XNOR2_X1 U21771 ( .A(n21333), .B(n21184), .ZN(n20660) );
  XNOR2_X1 U21772 ( .A(n24100), .B(n21670), .ZN(n20658) );
  XNOR2_X1 U21773 ( .A(n20999), .B(n2903), .ZN(n20657) );
  XNOR2_X1 U21774 ( .A(n20658), .B(n20657), .ZN(n20659) );
  XNOR2_X1 U21775 ( .A(n20660), .B(n20659), .ZN(n22973) );
  AND2_X1 U21776 ( .A1(n22977), .A2(n3213), .ZN(n20684) );
  XNOR2_X1 U21777 ( .A(n20957), .B(n21696), .ZN(n20664) );
  XNOR2_X1 U21778 ( .A(n21492), .B(n21399), .ZN(n20662) );
  XNOR2_X1 U21779 ( .A(n25377), .B(n912), .ZN(n20661) );
  XNOR2_X1 U21780 ( .A(n20662), .B(n20661), .ZN(n20663) );
  INV_X1 U21781 ( .A(n20665), .ZN(n20675) );
  NAND2_X1 U21782 ( .A1(n20666), .A2(n20669), .ZN(n20667) );
  OAI211_X1 U21783 ( .C1(n20670), .C2(n20669), .A(n20668), .B(n20667), .ZN(
        n20674) );
  NAND2_X1 U21784 ( .A1(n20672), .A2(n20671), .ZN(n20673) );
  NAND3_X1 U21785 ( .A1(n20675), .A2(n20674), .A3(n20673), .ZN(n20676) );
  XNOR2_X1 U21786 ( .A(n20676), .B(n681), .ZN(n20678) );
  XNOR2_X1 U21787 ( .A(n21734), .B(n21699), .ZN(n20677) );
  XNOR2_X1 U21788 ( .A(n20914), .B(n21965), .ZN(n20972) );
  XNOR2_X1 U21789 ( .A(n20804), .B(n21665), .ZN(n20680) );
  XNOR2_X1 U21790 ( .A(n21302), .B(n20680), .ZN(n20683) );
  XNOR2_X1 U21791 ( .A(n21205), .B(n20964), .ZN(n20899) );
  XNOR2_X1 U21792 ( .A(n21040), .B(n1896), .ZN(n20681) );
  XNOR2_X1 U21793 ( .A(n20899), .B(n20681), .ZN(n20682) );
  XNOR2_X2 U21794 ( .A(n20683), .B(n20682), .ZN(n22387) );
  XNOR2_X1 U21795 ( .A(n21689), .B(n21160), .ZN(n20945) );
  XNOR2_X1 U21796 ( .A(n20798), .B(n21228), .ZN(n20736) );
  XNOR2_X1 U21797 ( .A(n20945), .B(n20736), .ZN(n20687) );
  XNOR2_X1 U21798 ( .A(n21422), .B(n1827), .ZN(n20685) );
  XNOR2_X1 U21799 ( .A(n21343), .B(n20685), .ZN(n20686) );
  XNOR2_X1 U21800 ( .A(n20687), .B(n20686), .ZN(n22972) );
  OR2_X1 U21802 ( .A1(n22387), .A2(n22972), .ZN(n22293) );
  OAI21_X1 U21803 ( .B1(n25365), .B2(n21891), .A(n22293), .ZN(n20688) );
  NOR2_X1 U21804 ( .A1(n23218), .A2(n23220), .ZN(n23215) );
  XNOR2_X1 U21805 ( .A(n21301), .B(n21554), .ZN(n21207) );
  XNOR2_X1 U21806 ( .A(n21975), .B(n21258), .ZN(n20689) );
  XNOR2_X1 U21807 ( .A(n21207), .B(n20689), .ZN(n20694) );
  XNOR2_X1 U21808 ( .A(n24491), .B(n21138), .ZN(n20692) );
  INV_X1 U21809 ( .A(n20690), .ZN(n22625) );
  XNOR2_X1 U21810 ( .A(n21172), .B(n22625), .ZN(n20691) );
  XNOR2_X1 U21811 ( .A(n20692), .B(n20691), .ZN(n20693) );
  INV_X1 U21812 ( .A(n2717), .ZN(n22549) );
  XNOR2_X1 U21813 ( .A(n21573), .B(n22549), .ZN(n20696) );
  XNOR2_X1 U21814 ( .A(n21622), .B(n21324), .ZN(n20695) );
  XNOR2_X1 U21815 ( .A(n20696), .B(n20695), .ZN(n20699) );
  XNOR2_X1 U21816 ( .A(n21694), .B(n21720), .ZN(n21460) );
  XNOR2_X1 U21817 ( .A(n20697), .B(n21070), .ZN(n21216) );
  XNOR2_X1 U21818 ( .A(n21216), .B(n21460), .ZN(n20698) );
  XNOR2_X1 U21819 ( .A(n20699), .B(n20698), .ZN(n21934) );
  INV_X1 U21820 ( .A(n21318), .ZN(n20701) );
  XNOR2_X1 U21821 ( .A(n21561), .B(n22702), .ZN(n20702) );
  XNOR2_X1 U21822 ( .A(n20867), .B(n20702), .ZN(n20705) );
  XNOR2_X1 U21823 ( .A(n21735), .B(n21704), .ZN(n21480) );
  INV_X1 U21824 ( .A(n21480), .ZN(n20703) );
  XNOR2_X1 U21825 ( .A(n20703), .B(n21429), .ZN(n20704) );
  XNOR2_X1 U21827 ( .A(n21445), .B(n21227), .ZN(n20707) );
  XNOR2_X1 U21828 ( .A(n21157), .B(n1776), .ZN(n20706) );
  XNOR2_X1 U21829 ( .A(n20707), .B(n20706), .ZN(n20710) );
  XNOR2_X1 U21830 ( .A(n21229), .B(n20708), .ZN(n20709) );
  INV_X1 U21831 ( .A(n21934), .ZN(n22563) );
  XNOR2_X1 U21832 ( .A(n21310), .B(n25265), .ZN(n21153) );
  XNOR2_X1 U21833 ( .A(n20831), .B(n21153), .ZN(n20713) );
  INV_X1 U21834 ( .A(n24287), .ZN(n22767) );
  XNOR2_X1 U21835 ( .A(n21676), .B(n22767), .ZN(n20711) );
  XNOR2_X1 U21836 ( .A(n21601), .B(n21312), .ZN(n21191) );
  XNOR2_X1 U21837 ( .A(n21191), .B(n20711), .ZN(n20712) );
  XNOR2_X2 U21838 ( .A(n20712), .B(n20713), .ZN(n22409) );
  OAI21_X1 U21839 ( .B1(n22406), .B2(n24951), .A(n20714), .ZN(n20721) );
  XNOR2_X1 U21840 ( .A(n21331), .B(n21578), .ZN(n21198) );
  XNOR2_X1 U21841 ( .A(n21253), .B(n21198), .ZN(n20718) );
  XNOR2_X1 U21842 ( .A(n21582), .B(n21334), .ZN(n20716) );
  XNOR2_X1 U21843 ( .A(n25386), .B(n1864), .ZN(n20715) );
  XNOR2_X1 U21844 ( .A(n20716), .B(n20715), .ZN(n20717) );
  XNOR2_X1 U21845 ( .A(n20718), .B(n20717), .ZN(n22407) );
  NAND2_X1 U21846 ( .A1(n24971), .A2(n22407), .ZN(n20719) );
  AOI21_X1 U21847 ( .B1(n22132), .B2(n20719), .A(n22133), .ZN(n20720) );
  INV_X1 U21849 ( .A(n24955), .ZN(n23229) );
  XNOR2_X1 U21850 ( .A(n21454), .B(n20722), .ZN(n20726) );
  XNOR2_X1 U21851 ( .A(n21505), .B(n1826), .ZN(n20724) );
  XNOR2_X1 U21852 ( .A(n20724), .B(n20723), .ZN(n20725) );
  XNOR2_X1 U21853 ( .A(n20725), .B(n20726), .ZN(n21380) );
  XNOR2_X1 U21854 ( .A(n21399), .B(n21212), .ZN(n20729) );
  XNOR2_X1 U21855 ( .A(n20727), .B(n2208), .ZN(n20728) );
  XNOR2_X1 U21856 ( .A(n20728), .B(n20729), .ZN(n20731) );
  XNOR2_X1 U21857 ( .A(n21721), .B(n21087), .ZN(n21461) );
  XNOR2_X1 U21858 ( .A(n21461), .B(n20954), .ZN(n20730) );
  XNOR2_X1 U21859 ( .A(n21514), .B(n21998), .ZN(n20732) );
  XNOR2_X1 U21860 ( .A(n20732), .B(n24985), .ZN(n21110) );
  XNOR2_X1 U21861 ( .A(n20733), .B(n20999), .ZN(n20734) );
  XNOR2_X1 U21862 ( .A(n20734), .B(n21121), .ZN(n20735) );
  XNOR2_X1 U21863 ( .A(n21587), .B(n21541), .ZN(n20737) );
  XNOR2_X1 U21864 ( .A(n20736), .B(n20737), .ZN(n20740) );
  XNOR2_X1 U21865 ( .A(n22007), .B(n21751), .ZN(n21449) );
  XNOR2_X1 U21866 ( .A(n22006), .B(n881), .ZN(n20738) );
  XNOR2_X1 U21867 ( .A(n21449), .B(n20738), .ZN(n20739) );
  XNOR2_X1 U21868 ( .A(n20739), .B(n20740), .ZN(n22455) );
  XNOR2_X1 U21869 ( .A(n20741), .B(n21967), .ZN(n20743) );
  XNOR2_X1 U21870 ( .A(n21559), .B(n20742), .ZN(n20969) );
  XNOR2_X1 U21871 ( .A(n20743), .B(n20969), .ZN(n20746) );
  INV_X1 U21872 ( .A(n20744), .ZN(n23183) );
  XNOR2_X1 U21873 ( .A(n21469), .B(n21713), .ZN(n22012) );
  XNOR2_X1 U21874 ( .A(n22012), .B(n21116), .ZN(n20750) );
  XNOR2_X1 U21875 ( .A(n21193), .B(n24936), .ZN(n20748) );
  XNOR2_X1 U21876 ( .A(n21639), .B(Key[190]), .ZN(n20747) );
  XNOR2_X1 U21877 ( .A(n20748), .B(n20747), .ZN(n20749) );
  NOR2_X1 U21878 ( .A1(n1352), .A2(n22453), .ZN(n22326) );
  NOR2_X1 U21879 ( .A1(n23229), .A2(n23227), .ZN(n20787) );
  XNOR2_X1 U21880 ( .A(n21027), .B(n21297), .ZN(n21005) );
  XNOR2_X1 U21881 ( .A(n21975), .B(n23750), .ZN(n20751) );
  XNOR2_X1 U21882 ( .A(n21005), .B(n20751), .ZN(n20753) );
  XNOR2_X1 U21883 ( .A(n21616), .B(n21040), .ZN(n21262) );
  XNOR2_X1 U21884 ( .A(n21173), .B(n21136), .ZN(n20808) );
  XNOR2_X1 U21885 ( .A(n20808), .B(n21262), .ZN(n20752) );
  XNOR2_X1 U21886 ( .A(n20753), .B(n20752), .ZN(n22134) );
  XNOR2_X1 U21887 ( .A(n21133), .B(n21247), .ZN(n21626) );
  XNOR2_X1 U21888 ( .A(n21245), .B(n21693), .ZN(n20992) );
  XNOR2_X1 U21889 ( .A(n20992), .B(n21626), .ZN(n20757) );
  XNOR2_X1 U21890 ( .A(n21573), .B(n1801), .ZN(n20755) );
  XNOR2_X1 U21891 ( .A(n25377), .B(n25385), .ZN(n20754) );
  XNOR2_X1 U21892 ( .A(n20755), .B(n20754), .ZN(n20756) );
  XNOR2_X1 U21893 ( .A(n20757), .B(n20756), .ZN(n21888) );
  AND2_X1 U21894 ( .A1(n22134), .A2(n22401), .ZN(n20775) );
  XNOR2_X1 U21895 ( .A(n21126), .B(n21273), .ZN(n21632) );
  XNOR2_X1 U21896 ( .A(n21561), .B(n21053), .ZN(n20758) );
  XNOR2_X1 U21897 ( .A(n21632), .B(n20758), .ZN(n20761) );
  XNOR2_X1 U21898 ( .A(n21176), .B(n20982), .ZN(n21316) );
  XNOR2_X1 U21899 ( .A(n21734), .B(n3344), .ZN(n20759) );
  XNOR2_X1 U21900 ( .A(n20759), .B(n21316), .ZN(n20760) );
  XNOR2_X1 U21901 ( .A(n20761), .B(n20760), .ZN(n22397) );
  XNOR2_X1 U21902 ( .A(n21158), .B(n21142), .ZN(n20797) );
  XNOR2_X1 U21903 ( .A(n20762), .B(n20797), .ZN(n20766) );
  XNOR2_X1 U21904 ( .A(n21227), .B(n21266), .ZN(n20764) );
  XNOR2_X1 U21905 ( .A(n21267), .B(n2222), .ZN(n20763) );
  XNOR2_X1 U21906 ( .A(n20764), .B(n20763), .ZN(n20765) );
  XNOR2_X1 U21907 ( .A(n20766), .B(n20765), .ZN(n20776) );
  INV_X1 U21908 ( .A(n20776), .ZN(n22265) );
  NOR2_X1 U21909 ( .A1(n22265), .A2(n22401), .ZN(n20774) );
  INV_X1 U21910 ( .A(n21311), .ZN(n20768) );
  XNOR2_X1 U21911 ( .A(n20768), .B(n20767), .ZN(n21241) );
  XNOR2_X1 U21912 ( .A(n21241), .B(n20769), .ZN(n20773) );
  XNOR2_X1 U21913 ( .A(n21414), .B(n21115), .ZN(n20771) );
  XNOR2_X1 U21914 ( .A(n21596), .B(n765), .ZN(n20770) );
  XNOR2_X1 U21915 ( .A(n20771), .B(n20770), .ZN(n20772) );
  AOI22_X1 U21917 ( .A1(n20775), .A2(n22397), .B1(n20774), .B2(n22398), .ZN(
        n20786) );
  INV_X1 U21918 ( .A(n2049), .ZN(n20777) );
  XNOR2_X1 U21919 ( .A(n20779), .B(n21648), .ZN(n20783) );
  XNOR2_X1 U21920 ( .A(n21332), .B(n20780), .ZN(n21254) );
  XNOR2_X1 U21921 ( .A(n21254), .B(n20781), .ZN(n20782) );
  AOI21_X1 U21922 ( .B1(n25381), .B2(n22400), .A(n22134), .ZN(n20784) );
  OAI21_X1 U21923 ( .B1(n22400), .B2(n21885), .A(n20784), .ZN(n20785) );
  OAI21_X1 U21925 ( .B1(n23215), .B2(n20787), .A(n23231), .ZN(n20824) );
  INV_X1 U21926 ( .A(n1340), .ZN(n23213) );
  XNOR2_X1 U21928 ( .A(n21108), .B(n21668), .ZN(n20791) );
  XNOR2_X1 U21929 ( .A(n21579), .B(n25091), .ZN(n20789) );
  XNOR2_X1 U21930 ( .A(n20999), .B(n3798), .ZN(n20788) );
  XNOR2_X1 U21931 ( .A(n20789), .B(n20788), .ZN(n20790) );
  XNOR2_X1 U21932 ( .A(n20791), .B(n20790), .ZN(n21375) );
  XNOR2_X1 U21934 ( .A(n21307), .B(n24916), .ZN(n20794) );
  XNOR2_X1 U21935 ( .A(n20792), .B(n812), .ZN(n20793) );
  INV_X1 U21936 ( .A(n21523), .ZN(n20927) );
  XNOR2_X1 U21938 ( .A(n20795), .B(n20927), .ZN(n21683) );
  XNOR2_X1 U21939 ( .A(n22005), .B(n21444), .ZN(n21684) );
  XNOR2_X1 U21940 ( .A(n20797), .B(n21684), .ZN(n20802) );
  XNOR2_X1 U21941 ( .A(n20798), .B(n21141), .ZN(n20800) );
  XNOR2_X1 U21942 ( .A(n21686), .B(n2726), .ZN(n20799) );
  XNOR2_X1 U21943 ( .A(n20800), .B(n20799), .ZN(n20801) );
  NOR2_X1 U21945 ( .A1(n1363), .A2(n22459), .ZN(n20803) );
  XNOR2_X1 U21946 ( .A(n20804), .B(n21979), .ZN(n20807) );
  XNOR2_X1 U21947 ( .A(n21658), .B(n20805), .ZN(n20806) );
  XNOR2_X1 U21948 ( .A(n20807), .B(n20806), .ZN(n20810) );
  XNOR2_X1 U21949 ( .A(n21659), .B(n21660), .ZN(n21503) );
  XNOR2_X1 U21950 ( .A(n20808), .B(n21503), .ZN(n20809) );
  XNOR2_X1 U21951 ( .A(n21971), .B(n21701), .ZN(n20813) );
  XNOR2_X1 U21952 ( .A(n21567), .B(n921), .ZN(n20815) );
  XNOR2_X1 U21953 ( .A(n20817), .B(n20816), .ZN(n20819) );
  XNOR2_X2 U21955 ( .A(n20819), .B(n21697), .ZN(n22464) );
  AOI21_X1 U21956 ( .B1(n22462), .B2(n22465), .A(n3908), .ZN(n20821) );
  NAND2_X1 U21957 ( .A1(n21929), .A2(n24367), .ZN(n20820) );
  AOI21_X1 U21958 ( .B1(n23213), .B2(n23219), .A(n20822), .ZN(n20823) );
  INV_X1 U21959 ( .A(n20825), .ZN(n21398) );
  XNOR2_X1 U21960 ( .A(n21449), .B(n22004), .ZN(n20829) );
  XNOR2_X1 U21961 ( .A(n21686), .B(n1835), .ZN(n20827) );
  XNOR2_X1 U21962 ( .A(n20881), .B(n20827), .ZN(n20828) );
  XNOR2_X1 U21963 ( .A(n20829), .B(n20828), .ZN(n20845) );
  INV_X1 U21964 ( .A(n20845), .ZN(n22176) );
  XNOR2_X1 U21965 ( .A(n21193), .B(n21469), .ZN(n20830) );
  XNOR2_X1 U21966 ( .A(n20831), .B(n20830), .ZN(n20835) );
  XNOR2_X1 U21967 ( .A(n21520), .B(n21523), .ZN(n20833) );
  XNOR2_X1 U21968 ( .A(n20870), .B(n859), .ZN(n20832) );
  XNOR2_X1 U21969 ( .A(n20833), .B(n20832), .ZN(n20834) );
  XNOR2_X1 U21970 ( .A(n21087), .B(n21495), .ZN(n21986) );
  XNOR2_X1 U21971 ( .A(n21135), .B(n21622), .ZN(n20860) );
  XNOR2_X1 U21972 ( .A(n21986), .B(n20860), .ZN(n20838) );
  XNOR2_X1 U21973 ( .A(n25222), .B(n1855), .ZN(n20836) );
  XNOR2_X1 U21974 ( .A(n25442), .B(n20836), .ZN(n20837) );
  XNOR2_X2 U21975 ( .A(n20837), .B(n20838), .ZN(n22175) );
  BUF_X2 U21976 ( .A(n22175), .Z(n22200) );
  XNOR2_X1 U21977 ( .A(n21200), .B(n20839), .ZN(n20844) );
  XNOR2_X1 U21978 ( .A(n21998), .B(n20840), .ZN(n20841) );
  XNOR2_X1 U21979 ( .A(n20842), .B(n20841), .ZN(n20843) );
  XNOR2_X1 U21980 ( .A(n20844), .B(n20843), .ZN(n21759) );
  MUX2_X1 U21981 ( .A(n22197), .B(n4360), .S(n23571), .Z(n20846) );
  INV_X1 U21982 ( .A(n21222), .ZN(n21536) );
  XNOR2_X1 U21984 ( .A(n20847), .B(n21970), .ZN(n20850) );
  XNOR2_X1 U21985 ( .A(n21224), .B(n20848), .ZN(n20849) );
  NOR2_X1 U21987 ( .A1(n325), .A2(n22200), .ZN(n20856) );
  XNOR2_X1 U21988 ( .A(n21743), .B(n2477), .ZN(n20851) );
  XNOR2_X1 U21989 ( .A(n20851), .B(n25498), .ZN(n20852) );
  XNOR2_X1 U21990 ( .A(n21208), .B(n20852), .ZN(n20855) );
  XNOR2_X1 U21991 ( .A(n21980), .B(n21258), .ZN(n20853) );
  XNOR2_X1 U21992 ( .A(n20853), .B(n21981), .ZN(n20854) );
  INV_X1 U21993 ( .A(n23619), .ZN(n23637) );
  XNOR2_X1 U21994 ( .A(n1326), .B(n887), .ZN(n20857) );
  XNOR2_X1 U21995 ( .A(n21207), .B(n20857), .ZN(n20859) );
  XNOR2_X1 U21996 ( .A(n21501), .B(n21258), .ZN(n21615) );
  XNOR2_X1 U21997 ( .A(n21551), .B(n21615), .ZN(n20858) );
  XNOR2_X1 U21998 ( .A(n21492), .B(n21567), .ZN(n21326) );
  XNOR2_X1 U21999 ( .A(n21326), .B(n20860), .ZN(n20863) );
  XNOR2_X1 U22000 ( .A(n24996), .B(n187), .ZN(n20861) );
  XNOR2_X1 U22001 ( .A(n21216), .B(n20861), .ZN(n20862) );
  XNOR2_X1 U22003 ( .A(n21481), .B(n20864), .ZN(n20865) );
  XNOR2_X1 U22004 ( .A(n20865), .B(n21633), .ZN(n20866) );
  XNOR2_X1 U22005 ( .A(n20866), .B(n21562), .ZN(n20868) );
  XNOR2_X1 U22006 ( .A(n20868), .B(n20867), .ZN(n22889) );
  INV_X1 U22008 ( .A(n20870), .ZN(n21471) );
  XNOR2_X1 U22009 ( .A(n21471), .B(n21307), .ZN(n20871) );
  XNOR2_X1 U22010 ( .A(n21191), .B(n20871), .ZN(n20880) );
  XNOR2_X1 U22011 ( .A(n21525), .B(n25065), .ZN(n20878) );
  NAND3_X1 U22012 ( .A1(n20872), .A2(n23225), .A3(n20412), .ZN(n20875) );
  NAND3_X1 U22013 ( .A1(n20873), .A2(n1754), .A3(n20876), .ZN(n20874) );
  OAI211_X1 U22014 ( .C1(n1754), .C2(n20876), .A(n20875), .B(n20874), .ZN(
        n20877) );
  XNOR2_X1 U22015 ( .A(n20878), .B(n20877), .ZN(n20879) );
  XNOR2_X1 U22017 ( .A(n21229), .B(n20881), .ZN(n20886) );
  XNOR2_X1 U22018 ( .A(n24485), .B(n1768), .ZN(n20884) );
  XNOR2_X1 U22019 ( .A(n21158), .B(n21606), .ZN(n20883) );
  XNOR2_X1 U22020 ( .A(n20884), .B(n20883), .ZN(n20885) );
  XNOR2_X1 U22021 ( .A(n21649), .B(n23620), .ZN(n20888) );
  XNOR2_X1 U22022 ( .A(n21579), .B(n21728), .ZN(n20887) );
  XNOR2_X1 U22023 ( .A(n20887), .B(n20888), .ZN(n20891) );
  XNOR2_X1 U22024 ( .A(n21198), .B(n20889), .ZN(n20890) );
  XNOR2_X1 U22025 ( .A(n20891), .B(n20890), .ZN(n22728) );
  NOR2_X1 U22026 ( .A1(n22889), .A2(n25375), .ZN(n20894) );
  INV_X1 U22027 ( .A(n23634), .ZN(n20896) );
  INV_X1 U22028 ( .A(n21974), .ZN(n20897) );
  XNOR2_X1 U22029 ( .A(n21550), .B(n20897), .ZN(n21747) );
  XNOR2_X1 U22030 ( .A(n21747), .B(n20898), .ZN(n20902) );
  XNOR2_X1 U22031 ( .A(n25498), .B(n2745), .ZN(n20900) );
  XNOR2_X1 U22032 ( .A(n20900), .B(n20899), .ZN(n20901) );
  XNOR2_X2 U22033 ( .A(n20902), .B(n20901), .ZN(n22159) );
  XNOR2_X1 U22034 ( .A(n21694), .B(n21212), .ZN(n20903) );
  XNOR2_X1 U22035 ( .A(n20904), .B(n449), .ZN(n20905) );
  XNOR2_X1 U22036 ( .A(n20905), .B(n25222), .ZN(n20907) );
  XNOR2_X1 U22037 ( .A(n21568), .B(n21621), .ZN(n20906) );
  XNOR2_X1 U22038 ( .A(n20907), .B(n20906), .ZN(n20908) );
  NOR2_X1 U22039 ( .A1(n22159), .A2(n25485), .ZN(n22212) );
  XNOR2_X1 U22040 ( .A(n21736), .B(n2991), .ZN(n20916) );
  XNOR2_X1 U22041 ( .A(n20914), .B(n21532), .ZN(n20915) );
  XNOR2_X1 U22042 ( .A(n20916), .B(n20915), .ZN(n20917) );
  XNOR2_X1 U22043 ( .A(n21699), .B(n21704), .ZN(n21129) );
  XNOR2_X1 U22044 ( .A(n20917), .B(n21129), .ZN(n20918) );
  XNOR2_X1 U22045 ( .A(n21971), .B(n21967), .ZN(n21538) );
  XNOR2_X1 U22046 ( .A(n21445), .B(n21228), .ZN(n21685) );
  XNOR2_X1 U22047 ( .A(n21686), .B(n21141), .ZN(n21543) );
  XNOR2_X1 U22048 ( .A(n21685), .B(n21543), .ZN(n20922) );
  XNOR2_X1 U22049 ( .A(n21591), .B(n22739), .ZN(n20920) );
  XNOR2_X1 U22050 ( .A(n22006), .B(n21160), .ZN(n20919) );
  XNOR2_X1 U22051 ( .A(n20920), .B(n20919), .ZN(n20921) );
  XNOR2_X1 U22052 ( .A(n20922), .B(n20921), .ZN(n22209) );
  XNOR2_X1 U22053 ( .A(n20948), .B(n21678), .ZN(n20923) );
  XNOR2_X1 U22054 ( .A(n21114), .B(n20923), .ZN(n20931) );
  INV_X1 U22055 ( .A(n21713), .ZN(n20924) );
  XNOR2_X1 U22056 ( .A(n21599), .B(n20924), .ZN(n20929) );
  AOI21_X1 U22057 ( .B1(n20927), .B2(n3115), .A(n20926), .ZN(n20928) );
  XNOR2_X1 U22058 ( .A(n20929), .B(n20928), .ZN(n20930) );
  AOI22_X1 U22059 ( .A1(n22212), .A2(n2315), .B1(n20932), .B2(n25018), .ZN(
        n20942) );
  XNOR2_X1 U22060 ( .A(n21992), .B(n21670), .ZN(n20934) );
  XNOR2_X1 U22061 ( .A(n21997), .B(n21577), .ZN(n20933) );
  XNOR2_X1 U22062 ( .A(n20934), .B(n20933), .ZN(n20939) );
  XNOR2_X1 U22063 ( .A(n21515), .B(n21439), .ZN(n20937) );
  INV_X1 U22064 ( .A(n2236), .ZN(n20935) );
  XNOR2_X1 U22065 ( .A(n21647), .B(n20935), .ZN(n20936) );
  XNOR2_X1 U22066 ( .A(n20937), .B(n20936), .ZN(n20938) );
  XNOR2_X1 U22067 ( .A(n20939), .B(n20938), .ZN(n21766) );
  INV_X1 U22068 ( .A(n22205), .ZN(n22156) );
  OAI21_X1 U22069 ( .B1(n22064), .B2(n22156), .A(n22159), .ZN(n20940) );
  XNOR2_X1 U22071 ( .A(n21587), .B(n21267), .ZN(n20944) );
  XNOR2_X1 U22072 ( .A(n22005), .B(n1815), .ZN(n20943) );
  XNOR2_X1 U22073 ( .A(n20944), .B(n20943), .ZN(n20947) );
  XNOR2_X1 U22074 ( .A(n21142), .B(n21541), .ZN(n21612) );
  XNOR2_X1 U22075 ( .A(n21612), .B(n20945), .ZN(n20946) );
  XNOR2_X1 U22076 ( .A(n20946), .B(n20947), .ZN(n22916) );
  XNOR2_X1 U22077 ( .A(n21115), .B(n20948), .ZN(n20949) );
  XNOR2_X1 U22078 ( .A(n21096), .B(n20949), .ZN(n20953) );
  XNOR2_X1 U22079 ( .A(n22014), .B(n24962), .ZN(n20951) );
  XNOR2_X1 U22080 ( .A(n21311), .B(n1746), .ZN(n20950) );
  XNOR2_X1 U22081 ( .A(n20951), .B(n20950), .ZN(n20952) );
  XNOR2_X1 U22082 ( .A(n20953), .B(n20952), .ZN(n22070) );
  NOR2_X1 U22083 ( .A1(n22916), .A2(n24902), .ZN(n22116) );
  XNOR2_X1 U22084 ( .A(n21084), .B(n21133), .ZN(n20955) );
  XNOR2_X1 U22085 ( .A(n20954), .B(n20955), .ZN(n20959) );
  XNOR2_X1 U22086 ( .A(n21245), .B(n2990), .ZN(n20956) );
  XNOR2_X1 U22087 ( .A(n20957), .B(n20956), .ZN(n20958) );
  XNOR2_X1 U22088 ( .A(n21658), .B(n21452), .ZN(n21977) );
  XNOR2_X1 U22089 ( .A(n21136), .B(n21505), .ZN(n21614) );
  XNOR2_X1 U22090 ( .A(n21977), .B(n21614), .ZN(n20968) );
  XNOR2_X1 U22091 ( .A(n20964), .B(n1804), .ZN(n20965) );
  XNOR2_X1 U22092 ( .A(n20965), .B(n21297), .ZN(n20966) );
  XNOR2_X1 U22093 ( .A(n20966), .B(n24898), .ZN(n20967) );
  NAND2_X1 U22094 ( .A1(n22918), .A2(n22072), .ZN(n22115) );
  XNOR2_X1 U22095 ( .A(n25202), .B(n21126), .ZN(n20970) );
  XNOR2_X1 U22096 ( .A(n20970), .B(n20969), .ZN(n20974) );
  XNOR2_X1 U22097 ( .A(n20982), .B(n2989), .ZN(n20971) );
  XNOR2_X1 U22098 ( .A(n20972), .B(n20971), .ZN(n20973) );
  NAND2_X1 U22100 ( .A1(n22917), .A2(n22072), .ZN(n22169) );
  INV_X1 U22101 ( .A(n22115), .ZN(n20980) );
  INV_X1 U22102 ( .A(Key[38]), .ZN(n20975) );
  XNOR2_X1 U22103 ( .A(n21996), .B(n21514), .ZN(n20976) );
  XNOR2_X1 U22104 ( .A(n21648), .B(n20976), .ZN(n20977) );
  NOR2_X1 U22105 ( .A1(n22166), .A2(n22072), .ZN(n20979) );
  AOI22_X1 U22106 ( .A1(n20981), .A2(n23637), .B1(n23648), .B2(n23649), .ZN(
        n21078) );
  XNOR2_X1 U22107 ( .A(n20983), .B(n20982), .ZN(n20985) );
  XNOR2_X1 U22108 ( .A(n20985), .B(n20984), .ZN(n20988) );
  INV_X1 U22109 ( .A(n21053), .ZN(n20986) );
  XNOR2_X1 U22110 ( .A(n21534), .B(n20986), .ZN(n21706) );
  XNOR2_X1 U22111 ( .A(n21706), .B(n21429), .ZN(n20987) );
  XNOR2_X1 U22112 ( .A(n21070), .B(n21399), .ZN(n20989) );
  XNOR2_X1 U22113 ( .A(n20990), .B(n20989), .ZN(n20994) );
  XNOR2_X1 U22114 ( .A(n20992), .B(n20991), .ZN(n20993) );
  XNOR2_X1 U22116 ( .A(n21415), .B(n21241), .ZN(n20998) );
  INV_X1 U22117 ( .A(n20995), .ZN(n23945) );
  XNOR2_X1 U22118 ( .A(n24899), .B(n23945), .ZN(n20996) );
  XNOR2_X1 U22119 ( .A(n21023), .B(n20996), .ZN(n20997) );
  XNOR2_X1 U22121 ( .A(n21182), .B(n21510), .ZN(n21669) );
  XNOR2_X1 U22122 ( .A(n21254), .B(n21669), .ZN(n21002) );
  XNOR2_X1 U22123 ( .A(n21334), .B(n20999), .ZN(n21392) );
  XNOR2_X1 U22124 ( .A(n21578), .B(n3131), .ZN(n21000) );
  XNOR2_X1 U22125 ( .A(n21392), .B(n21000), .ZN(n21001) );
  XNOR2_X1 U22126 ( .A(n21002), .B(n21001), .ZN(n22923) );
  INV_X1 U22127 ( .A(n22923), .ZN(n22712) );
  XNOR2_X1 U22129 ( .A(n21409), .B(n21003), .ZN(n21007) );
  XNOR2_X1 U22130 ( .A(n21554), .B(n3164), .ZN(n21004) );
  XNOR2_X1 U22131 ( .A(n21005), .B(n21004), .ZN(n21006) );
  INV_X1 U22132 ( .A(n22927), .ZN(n22188) );
  NAND2_X1 U22133 ( .A1(n22926), .A2(n22188), .ZN(n21020) );
  NAND2_X1 U22134 ( .A1(n21009), .A2(n21008), .ZN(n21011) );
  NAND2_X1 U22135 ( .A1(n21011), .A2(n21010), .ZN(n21012) );
  XNOR2_X1 U22136 ( .A(n21043), .B(n21687), .ZN(n21015) );
  XNOR2_X1 U22137 ( .A(n21267), .B(n2241), .ZN(n21014) );
  XNOR2_X1 U22138 ( .A(n21015), .B(n21014), .ZN(n21018) );
  XNOR2_X1 U22139 ( .A(n25400), .B(n21266), .ZN(n21016) );
  XNOR2_X1 U22140 ( .A(n21420), .B(n21016), .ZN(n21017) );
  XNOR2_X1 U22141 ( .A(n21017), .B(n21018), .ZN(n22922) );
  NAND2_X1 U22142 ( .A1(n22923), .A2(n22922), .ZN(n21019) );
  OAI21_X1 U22143 ( .B1(n22926), .B2(n22927), .A(n21019), .ZN(n22711) );
  XNOR2_X1 U22144 ( .A(n25265), .B(n21414), .ZN(n21025) );
  XNOR2_X1 U22145 ( .A(n21025), .B(n21600), .ZN(n21243) );
  XNOR2_X1 U22147 ( .A(n21027), .B(n2882), .ZN(n21028) );
  XNOR2_X1 U22148 ( .A(n21028), .B(n20475), .ZN(n21029) );
  OAI21_X1 U22149 ( .B1(n21033), .B2(n24378), .A(n21031), .ZN(n21037) );
  AOI21_X1 U22150 ( .B1(n21035), .B2(n21034), .A(n21038), .ZN(n21036) );
  AOI21_X1 U22151 ( .B1(n21038), .B2(n21037), .A(n21036), .ZN(n21039) );
  XNOR2_X1 U22152 ( .A(n21041), .B(n21040), .ZN(n21748) );
  INV_X1 U22153 ( .A(n22245), .ZN(n22240) );
  XNOR2_X1 U22154 ( .A(n22007), .B(n21750), .ZN(n21044) );
  XNOR2_X1 U22155 ( .A(n21043), .B(n21042), .ZN(n21589) );
  XNOR2_X1 U22156 ( .A(n21044), .B(n21589), .ZN(n21050) );
  XNOR2_X1 U22157 ( .A(n24485), .B(n21045), .ZN(n21048) );
  XNOR2_X1 U22158 ( .A(n21422), .B(n21046), .ZN(n21047) );
  XNOR2_X1 U22159 ( .A(n21048), .B(n21047), .ZN(n21049) );
  XNOR2_X1 U22160 ( .A(n21050), .B(n21049), .ZN(n22239) );
  INV_X1 U22161 ( .A(n22239), .ZN(n22181) );
  XNOR2_X1 U22162 ( .A(n21477), .B(n21735), .ZN(n21052) );
  XNOR2_X1 U22163 ( .A(n21734), .B(n3093), .ZN(n21051) );
  XNOR2_X1 U22164 ( .A(n21052), .B(n21051), .ZN(n21057) );
  XNOR2_X1 U22165 ( .A(n24353), .B(n21053), .ZN(n21055) );
  INV_X1 U22166 ( .A(n21319), .ZN(n21054) );
  XNOR2_X1 U22167 ( .A(n21055), .B(n21564), .ZN(n21056) );
  OAI22_X1 U22168 ( .A1(n22243), .A2(n22240), .B1(n22181), .B2(n22244), .ZN(
        n21077) );
  XNOR2_X1 U22169 ( .A(n21058), .B(n21182), .ZN(n21060) );
  INV_X1 U22170 ( .A(n21336), .ZN(n21059) );
  XNOR2_X1 U22171 ( .A(n21059), .B(n21436), .ZN(n21726) );
  XNOR2_X1 U22172 ( .A(n21726), .B(n21060), .ZN(n21064) );
  XNOR2_X1 U22173 ( .A(n24100), .B(n2137), .ZN(n21062) );
  XNOR2_X1 U22174 ( .A(n21061), .B(n21062), .ZN(n21063) );
  XNOR2_X1 U22175 ( .A(n21064), .B(n21063), .ZN(n22242) );
  INV_X1 U22176 ( .A(n22242), .ZN(n22180) );
  XNOR2_X1 U22179 ( .A(n21071), .B(n21070), .ZN(n21574) );
  XNOR2_X1 U22180 ( .A(n21574), .B(n21246), .ZN(n21075) );
  XNOR2_X1 U22181 ( .A(n21087), .B(n21720), .ZN(n21073) );
  XNOR2_X1 U22182 ( .A(n21693), .B(n836), .ZN(n21072) );
  XNOR2_X1 U22183 ( .A(n21073), .B(n21072), .ZN(n21074) );
  XNOR2_X1 U22184 ( .A(n21074), .B(n21075), .ZN(n22059) );
  XNOR2_X1 U22186 ( .A(n25202), .B(n21630), .ZN(n21080) );
  XNOR2_X1 U22187 ( .A(n21477), .B(n2318), .ZN(n21081) );
  XNOR2_X1 U22189 ( .A(n25073), .B(n21084), .ZN(n21086) );
  XNOR2_X1 U22190 ( .A(n25040), .B(n21324), .ZN(n21085) );
  XNOR2_X1 U22191 ( .A(n21086), .B(n21085), .ZN(n21090) );
  XNOR2_X1 U22192 ( .A(n21087), .B(n1952), .ZN(n21088) );
  XNOR2_X1 U22193 ( .A(n21496), .B(n21088), .ZN(n21089) );
  INV_X1 U22194 ( .A(n21157), .ZN(n21091) );
  XNOR2_X1 U22195 ( .A(n21091), .B(n3125), .ZN(n21092) );
  XNOR2_X1 U22196 ( .A(n21612), .B(n21093), .ZN(n21094) );
  INV_X1 U22198 ( .A(n23998), .ZN(n22373) );
  XNOR2_X1 U22199 ( .A(n22012), .B(n21096), .ZN(n21100) );
  XNOR2_X1 U22200 ( .A(n21310), .B(n21115), .ZN(n21098) );
  XNOR2_X1 U22201 ( .A(n24899), .B(n2739), .ZN(n21097) );
  XNOR2_X1 U22202 ( .A(n21098), .B(n21097), .ZN(n21099) );
  XNOR2_X1 U22204 ( .A(n21172), .B(n21980), .ZN(n21101) );
  XNOR2_X1 U22205 ( .A(n24898), .B(n21101), .ZN(n21105) );
  XNOR2_X1 U22206 ( .A(n21974), .B(n763), .ZN(n21102) );
  XNOR2_X1 U22207 ( .A(n21102), .B(n21660), .ZN(n21103) );
  XNOR2_X1 U22208 ( .A(n21614), .B(n21103), .ZN(n21104) );
  XNOR2_X1 U22209 ( .A(n21107), .B(n21334), .ZN(n21109) );
  XNOR2_X1 U22210 ( .A(n21108), .B(n21109), .ZN(n21111) );
  AND2_X1 U22211 ( .A1(n24439), .A2(n25414), .ZN(n21112) );
  INV_X1 U22212 ( .A(n23997), .ZN(n21855) );
  OAI21_X1 U22213 ( .B1(n22676), .B2(n21112), .A(n21855), .ZN(n21113) );
  XNOR2_X1 U22214 ( .A(n21114), .B(n21716), .ZN(n21119) );
  XNOR2_X1 U22215 ( .A(n21115), .B(Key[172]), .ZN(n21117) );
  XNOR2_X1 U22216 ( .A(n21116), .B(n21117), .ZN(n21118) );
  XNOR2_X1 U22217 ( .A(n21119), .B(n21118), .ZN(n22667) );
  XNOR2_X1 U22218 ( .A(n21439), .B(n23699), .ZN(n21120) );
  XNOR2_X1 U22219 ( .A(n21120), .B(n21728), .ZN(n21122) );
  XNOR2_X1 U22220 ( .A(n21122), .B(n21121), .ZN(n21125) );
  XNOR2_X1 U22221 ( .A(n21336), .B(n25091), .ZN(n21123) );
  XNOR2_X1 U22222 ( .A(n21648), .B(n21123), .ZN(n21124) );
  OR2_X1 U22224 ( .A1(n22667), .A2(n25023), .ZN(n21147) );
  XNOR2_X1 U22225 ( .A(n21127), .B(n21126), .ZN(n21128) );
  XNOR2_X1 U22226 ( .A(n21739), .B(n21128), .ZN(n21131) );
  XNOR2_X1 U22227 ( .A(n21971), .B(n21129), .ZN(n21130) );
  XNOR2_X1 U22229 ( .A(n21132), .B(n1726), .ZN(n21134) );
  XNOR2_X1 U22231 ( .A(n21136), .B(n21506), .ZN(n21137) );
  XNOR2_X1 U22232 ( .A(n21452), .B(n21300), .ZN(n21556) );
  XNOR2_X1 U22233 ( .A(n21556), .B(n21137), .ZN(n21139) );
  OAI21_X1 U22234 ( .B1(n21147), .B2(n22675), .A(n22365), .ZN(n21149) );
  XNOR2_X1 U22235 ( .A(n21587), .B(n21141), .ZN(n22003) );
  XNOR2_X1 U22236 ( .A(n21685), .B(n22003), .ZN(n21145) );
  XNOR2_X1 U22237 ( .A(n21142), .B(n1739), .ZN(n21143) );
  XNOR2_X1 U22238 ( .A(n21755), .B(n21143), .ZN(n21144) );
  XNOR2_X1 U22239 ( .A(n21145), .B(n21144), .ZN(n22670) );
  INV_X1 U22240 ( .A(n22670), .ZN(n22784) );
  OAI22_X1 U22241 ( .A1(n21147), .A2(n25462), .B1(n22784), .B2(n21146), .ZN(
        n21148) );
  NAND2_X1 U22242 ( .A1(n23074), .A2(n25452), .ZN(n21239) );
  NOR3_X1 U22243 ( .A1(n22462), .A2(n24367), .A3(n25450), .ZN(n21150) );
  NAND2_X1 U22244 ( .A1(n21375), .A2(n22459), .ZN(n21930) );
  XNOR2_X1 U22246 ( .A(n21525), .B(n173), .ZN(n21152) );
  XNOR2_X1 U22247 ( .A(n21152), .B(n21679), .ZN(n21154) );
  XNOR2_X1 U22248 ( .A(n21154), .B(n21153), .ZN(n21155) );
  XNOR2_X1 U22249 ( .A(n21689), .B(n21606), .ZN(n21159) );
  XNOR2_X1 U22250 ( .A(n21157), .B(n21158), .ZN(n21342) );
  XNOR2_X1 U22251 ( .A(n21342), .B(n21159), .ZN(n21165) );
  INV_X1 U22252 ( .A(n1767), .ZN(n21161) );
  XNOR2_X1 U22253 ( .A(n21687), .B(n21161), .ZN(n21162) );
  XNOR2_X1 U22254 ( .A(n21163), .B(n21162), .ZN(n21164) );
  XNOR2_X1 U22255 ( .A(n21084), .B(n21720), .ZN(n21166) );
  XNOR2_X1 U22256 ( .A(n21326), .B(n21166), .ZN(n21168) );
  INV_X1 U22257 ( .A(n3084), .ZN(n23045) );
  XNOR2_X1 U22258 ( .A(n21501), .B(n21169), .ZN(n21170) );
  XNOR2_X1 U22259 ( .A(n21170), .B(n24491), .ZN(n21171) );
  XNOR2_X1 U22260 ( .A(n21171), .B(n21618), .ZN(n21175) );
  XNOR2_X1 U22261 ( .A(n21173), .B(n21172), .ZN(n21298) );
  XNOR2_X1 U22262 ( .A(n21298), .B(n24898), .ZN(n21174) );
  NOR2_X1 U22263 ( .A1(n24042), .A2(n274), .ZN(n21181) );
  XNOR2_X1 U22264 ( .A(n25202), .B(n24896), .ZN(n21177) );
  XNOR2_X1 U22265 ( .A(n25495), .B(n21177), .ZN(n21180) );
  XNOR2_X1 U22266 ( .A(n21735), .B(n1869), .ZN(n21178) );
  XNOR2_X1 U22267 ( .A(n21635), .B(n21178), .ZN(n21179) );
  AOI22_X1 U22268 ( .A1(n21923), .A2(n274), .B1(n21181), .B2(n22448), .ZN(
        n21190) );
  XNOR2_X1 U22269 ( .A(n21182), .B(n21511), .ZN(n21646) );
  XNOR2_X1 U22270 ( .A(n21436), .B(n21579), .ZN(n21183) );
  XNOR2_X1 U22271 ( .A(n21646), .B(n21183), .ZN(n21187) );
  XNOR2_X1 U22272 ( .A(n21334), .B(n3183), .ZN(n21185) );
  XNOR2_X1 U22273 ( .A(n21184), .B(n21185), .ZN(n21186) );
  XNOR2_X1 U22274 ( .A(n21191), .B(n21192), .ZN(n21197) );
  XNOR2_X1 U22275 ( .A(n21596), .B(n21678), .ZN(n21195) );
  XNOR2_X1 U22276 ( .A(n21193), .B(n1797), .ZN(n21194) );
  XNOR2_X1 U22277 ( .A(n21195), .B(n21194), .ZN(n21196) );
  XNOR2_X1 U22278 ( .A(n21199), .B(n21198), .ZN(n21203) );
  XNOR2_X1 U22279 ( .A(n21670), .B(n3152), .ZN(n21201) );
  XNOR2_X1 U22280 ( .A(n21200), .B(n21201), .ZN(n21202) );
  XNOR2_X1 U22282 ( .A(n24305), .B(n21204), .ZN(n21206) );
  XNOR2_X1 U22283 ( .A(n21207), .B(n21206), .ZN(n21211) );
  XNOR2_X2 U22284 ( .A(n21210), .B(n21211), .ZN(n22804) );
  INV_X1 U22285 ( .A(n21212), .ZN(n21213) );
  XNOR2_X1 U22286 ( .A(n21213), .B(n1364), .ZN(n21214) );
  XNOR2_X1 U22287 ( .A(n21215), .B(n21214), .ZN(n21219) );
  XNOR2_X1 U22288 ( .A(n21217), .B(n21216), .ZN(n21218) );
  MUX2_X1 U22290 ( .A(n22798), .B(n22804), .S(n24559), .Z(n21238) );
  XNOR2_X1 U22291 ( .A(n24434), .B(n2881), .ZN(n21220) );
  XNOR2_X1 U22292 ( .A(n21221), .B(n21220), .ZN(n21226) );
  XNOR2_X1 U22293 ( .A(n21318), .B(n21222), .ZN(n21223) );
  XNOR2_X1 U22294 ( .A(n21224), .B(n21223), .ZN(n21225) );
  XNOR2_X2 U22295 ( .A(n21225), .B(n21226), .ZN(n22800) );
  NOR2_X1 U22296 ( .A1(n22804), .A2(n22800), .ZN(n22583) );
  XNOR2_X1 U22297 ( .A(n21227), .B(n21228), .ZN(n21230) );
  XNOR2_X1 U22298 ( .A(n21229), .B(n21230), .ZN(n21235) );
  XNOR2_X1 U22299 ( .A(n21591), .B(n923), .ZN(n21232) );
  XNOR2_X1 U22300 ( .A(n21233), .B(n21232), .ZN(n21234) );
  INV_X1 U22302 ( .A(n22805), .ZN(n21236) );
  NOR2_X1 U22303 ( .A1(n21236), .A2(n22803), .ZN(n21237) );
  INV_X1 U22304 ( .A(n24561), .ZN(n22799) );
  XNOR2_X1 U22305 ( .A(n21640), .B(n2970), .ZN(n21240) );
  XNOR2_X1 U22306 ( .A(n21240), .B(n21520), .ZN(n21242) );
  XNOR2_X1 U22307 ( .A(n21241), .B(n21242), .ZN(n21244) );
  XNOR2_X1 U22308 ( .A(n21245), .B(n21622), .ZN(n21403) );
  XNOR2_X1 U22309 ( .A(n21246), .B(n21403), .ZN(n21251) );
  XNOR2_X1 U22310 ( .A(n21495), .B(n1924), .ZN(n21249) );
  XOR2_X1 U22311 ( .A(n21720), .B(n21247), .Z(n21248) );
  XNOR2_X1 U22312 ( .A(n21249), .B(n21248), .ZN(n21250) );
  XNOR2_X1 U22313 ( .A(n21251), .B(n21250), .ZN(n21265) );
  XNOR2_X1 U22314 ( .A(n21253), .B(n21252), .ZN(n21257) );
  XNOR2_X1 U22315 ( .A(n1381), .B(n2005), .ZN(n21255) );
  XNOR2_X1 U22316 ( .A(n21254), .B(n21255), .ZN(n21256) );
  XNOR2_X1 U22317 ( .A(n21297), .B(n21258), .ZN(n21408) );
  XNOR2_X1 U22318 ( .A(n21260), .B(n21259), .ZN(n21261) );
  XNOR2_X1 U22319 ( .A(n21261), .B(n21408), .ZN(n21264) );
  XNOR2_X1 U22320 ( .A(n21262), .B(n21981), .ZN(n21263) );
  XNOR2_X1 U22321 ( .A(n21264), .B(n21263), .ZN(n22619) );
  INV_X1 U22323 ( .A(n22792), .ZN(n22313) );
  INV_X1 U22324 ( .A(n21265), .ZN(n22612) );
  XNOR2_X1 U22325 ( .A(n21750), .B(n21266), .ZN(n21268) );
  XNOR2_X1 U22326 ( .A(n21608), .B(n21267), .ZN(n21421) );
  XNOR2_X1 U22327 ( .A(n21421), .B(n21268), .ZN(n21272) );
  XNOR2_X1 U22328 ( .A(n21422), .B(n1810), .ZN(n21269) );
  XNOR2_X1 U22329 ( .A(n21270), .B(n21269), .ZN(n21271) );
  XNOR2_X1 U22330 ( .A(n21272), .B(n21271), .ZN(n22791) );
  NAND3_X1 U22331 ( .A1(n22313), .A2(n22612), .A3(n22791), .ZN(n21279) );
  NAND2_X1 U22332 ( .A1(n22619), .A2(n22614), .ZN(n21370) );
  XNOR2_X1 U22333 ( .A(n24353), .B(n21273), .ZN(n21274) );
  XNOR2_X1 U22334 ( .A(n21430), .B(n21274), .ZN(n21278) );
  XNOR2_X1 U22335 ( .A(n21536), .B(n21735), .ZN(n21276) );
  XNOR2_X1 U22336 ( .A(n21734), .B(n2743), .ZN(n21275) );
  XNOR2_X1 U22337 ( .A(n21276), .B(n21275), .ZN(n21277) );
  XNOR2_X1 U22338 ( .A(n21278), .B(n21277), .ZN(n22615) );
  NAND2_X1 U22341 ( .A1(n21282), .A2(n21281), .ZN(n21284) );
  INV_X1 U22342 ( .A(n1789), .ZN(n21283) );
  XNOR2_X1 U22343 ( .A(n21284), .B(n21283), .ZN(Ciphertext[10]) );
  AND2_X1 U22344 ( .A1(n23217), .A2(n23228), .ZN(n21285) );
  AOI22_X1 U22345 ( .A1(n23215), .A2(n23219), .B1(n21285), .B2(n1340), .ZN(
        n21286) );
  INV_X1 U22346 ( .A(n21742), .ZN(n21287) );
  XNOR2_X1 U22347 ( .A(n21288), .B(n21287), .ZN(Ciphertext[39]) );
  INV_X1 U22348 ( .A(n21816), .ZN(n22687) );
  NOR2_X1 U22349 ( .A1(n22685), .A2(n22689), .ZN(n21290) );
  OAI21_X1 U22350 ( .B1(n21856), .B2(n22774), .A(n21292), .ZN(n21293) );
  INV_X1 U22351 ( .A(n22679), .ZN(n22771) );
  NAND2_X1 U22352 ( .A1(n21856), .A2(n22770), .ZN(n22682) );
  OR2_X1 U22353 ( .A1(n22682), .A2(n22370), .ZN(n21294) );
  INV_X1 U22355 ( .A(n21841), .ZN(n21840) );
  NOR2_X1 U22356 ( .A1(n23828), .A2(n891), .ZN(n21351) );
  XNOR2_X1 U22357 ( .A(n21297), .B(n1870), .ZN(n21299) );
  XNOR2_X1 U22358 ( .A(n21299), .B(n21298), .ZN(n21305) );
  XNOR2_X1 U22359 ( .A(n21301), .B(n21300), .ZN(n21303) );
  XNOR2_X1 U22360 ( .A(n21303), .B(n21302), .ZN(n21304) );
  INV_X1 U22362 ( .A(n22220), .ZN(n22216) );
  XNOR2_X1 U22363 ( .A(n21306), .B(n21307), .ZN(n21598) );
  XNOR2_X1 U22364 ( .A(n21308), .B(n21598), .ZN(n21315) );
  XNOR2_X1 U22365 ( .A(n21310), .B(n21309), .ZN(n21313) );
  XNOR2_X1 U22366 ( .A(n21311), .B(n25062), .ZN(n21416) );
  XNOR2_X1 U22367 ( .A(n21416), .B(n21313), .ZN(n21314) );
  XNOR2_X1 U22368 ( .A(n21317), .B(n21316), .ZN(n21323) );
  XNOR2_X1 U22369 ( .A(n21318), .B(n21965), .ZN(n21321) );
  XNOR2_X1 U22370 ( .A(n21319), .B(n2782), .ZN(n21320) );
  XNOR2_X1 U22371 ( .A(n21321), .B(n21320), .ZN(n21322) );
  MUX2_X1 U22373 ( .A(n22216), .B(n22222), .S(n22214), .Z(n21347) );
  XNOR2_X1 U22374 ( .A(n21325), .B(n21324), .ZN(n21400) );
  XNOR2_X1 U22375 ( .A(n21400), .B(n21326), .ZN(n21330) );
  XNOR2_X1 U22376 ( .A(n21985), .B(n2761), .ZN(n21327) );
  XNOR2_X1 U22377 ( .A(n21328), .B(n21327), .ZN(n21329) );
  XNOR2_X1 U22378 ( .A(n21332), .B(n21331), .ZN(n21395) );
  XNOR2_X1 U22379 ( .A(n21395), .B(n21333), .ZN(n21340) );
  XNOR2_X1 U22380 ( .A(n21579), .B(n21334), .ZN(n21338) );
  INV_X1 U22381 ( .A(n21335), .ZN(n23961) );
  XNOR2_X1 U22382 ( .A(n21336), .B(n23961), .ZN(n21337) );
  XNOR2_X1 U22383 ( .A(n21338), .B(n21337), .ZN(n21339) );
  XNOR2_X1 U22384 ( .A(n21340), .B(n21339), .ZN(n22219) );
  NAND2_X1 U22385 ( .A1(n22222), .A2(n22219), .ZN(n21341) );
  INV_X1 U22386 ( .A(n1951), .ZN(n23663) );
  OAI21_X2 U22387 ( .B1(n21347), .B2(n2817), .A(n21346), .ZN(n23827) );
  AND2_X1 U22388 ( .A1(n23827), .A2(n891), .ZN(n21361) );
  INV_X1 U22389 ( .A(n21361), .ZN(n21350) );
  INV_X1 U22390 ( .A(n23828), .ZN(n23834) );
  NAND2_X1 U22391 ( .A1(n23834), .A2(n891), .ZN(n21362) );
  AOI22_X1 U22392 ( .A1(n22231), .A2(n24905), .B1(n22226), .B2(n22225), .ZN(
        n22058) );
  NOR2_X1 U22393 ( .A1(n22058), .A2(n21794), .ZN(n21354) );
  AOI211_X1 U22394 ( .C1(n3231), .C2(n22228), .A(n22226), .B(n22056), .ZN(
        n21353) );
  INV_X1 U22395 ( .A(n23817), .ZN(n23811) );
  OAI22_X1 U22397 ( .A1(n21355), .A2(n23827), .B1(n23811), .B2(n21359), .ZN(
        n21356) );
  NAND2_X1 U22398 ( .A1(n23810), .A2(n23827), .ZN(n21358) );
  NAND2_X1 U22399 ( .A1(n21358), .A2(n24972), .ZN(n23034) );
  INV_X1 U22400 ( .A(n23034), .ZN(n21360) );
  NAND3_X1 U22401 ( .A1(n21360), .A2(n21359), .A3(n23827), .ZN(n21366) );
  NAND2_X1 U22402 ( .A1(n21364), .A2(n23034), .ZN(n21365) );
  INV_X1 U22403 ( .A(n22138), .ZN(n22334) );
  OAI21_X1 U22404 ( .B1(n22337), .B2(n22334), .A(n21368), .ZN(n21367) );
  INV_X1 U22406 ( .A(n22137), .ZN(n22274) );
  INV_X1 U22407 ( .A(n22791), .ZN(n22617) );
  NOR2_X1 U22408 ( .A1(n22789), .A2(n22614), .ZN(n21374) );
  INV_X1 U22409 ( .A(n21370), .ZN(n21373) );
  INV_X1 U22410 ( .A(n22615), .ZN(n22790) );
  OAI211_X1 U22411 ( .C1(n22614), .C2(n22790), .A(n22313), .B(n21371), .ZN(
        n21372) );
  INV_X1 U22413 ( .A(n23153), .ZN(n23138) );
  NOR2_X1 U22414 ( .A1(n1363), .A2(n21375), .ZN(n22328) );
  AND2_X1 U22415 ( .A1(n21375), .A2(n22464), .ZN(n21376) );
  INV_X1 U22416 ( .A(n22592), .ZN(n21921) );
  MUX2_X1 U22417 ( .A(n21921), .B(n2393), .S(n25066), .Z(n21378) );
  INV_X1 U22418 ( .A(n23129), .ZN(n23146) );
  INV_X1 U22419 ( .A(n21380), .ZN(n21918) );
  INV_X1 U22420 ( .A(n22453), .ZN(n21382) );
  NOR2_X1 U22421 ( .A1(n22455), .A2(n1352), .ZN(n21381) );
  AOI21_X1 U22422 ( .B1(n21382), .B2(n22455), .A(n21381), .ZN(n21385) );
  INV_X1 U22423 ( .A(n24311), .ZN(n21383) );
  NOR2_X1 U22424 ( .A1(n22456), .A2(n21383), .ZN(n21384) );
  AND2_X1 U22425 ( .A1(n22799), .A2(n22803), .ZN(n22806) );
  INV_X1 U22426 ( .A(n22800), .ZN(n21386) );
  AOI22_X1 U22427 ( .A1(n22806), .A2(n21386), .B1(n22803), .B2(n24992), .ZN(
        n21390) );
  INV_X1 U22431 ( .A(n2033), .ZN(n21391) );
  XNOR2_X1 U22432 ( .A(n24472), .B(n2746), .ZN(n21393) );
  XNOR2_X1 U22433 ( .A(n21392), .B(n21393), .ZN(n21397) );
  XNOR2_X1 U22434 ( .A(n24100), .B(n21577), .ZN(n21727) );
  XNOR2_X1 U22435 ( .A(n21395), .B(n21727), .ZN(n21396) );
  INV_X1 U22436 ( .A(n23334), .ZN(n21413) );
  XNOR2_X1 U22437 ( .A(n21399), .B(n21398), .ZN(n21401) );
  XNOR2_X1 U22438 ( .A(n21400), .B(n21401), .ZN(n21405) );
  XNOR2_X1 U22439 ( .A(n25377), .B(n21568), .ZN(n21723) );
  XNOR2_X1 U22440 ( .A(n21723), .B(n21403), .ZN(n21404) );
  XNOR2_X1 U22441 ( .A(n21550), .B(n2039), .ZN(n21407) );
  XNOR2_X1 U22442 ( .A(n21407), .B(n21406), .ZN(n21411) );
  XNOR2_X1 U22443 ( .A(n21409), .B(n21408), .ZN(n21410) );
  XNOR2_X1 U22446 ( .A(n21599), .B(n21414), .ZN(n21717) );
  XNOR2_X1 U22447 ( .A(n21415), .B(n21717), .ZN(n21419) );
  XNOR2_X1 U22448 ( .A(n25065), .B(n22635), .ZN(n21417) );
  XNOR2_X1 U22449 ( .A(n21417), .B(n21416), .ZN(n21418) );
  INV_X1 U22450 ( .A(n24342), .ZN(n22501) );
  XNOR2_X1 U22451 ( .A(n21420), .B(n21421), .ZN(n21426) );
  XNOR2_X1 U22452 ( .A(n21591), .B(n21422), .ZN(n21754) );
  INV_X1 U22453 ( .A(n21423), .ZN(n22525) );
  XNOR2_X1 U22454 ( .A(n21754), .B(n21424), .ZN(n21425) );
  INV_X1 U22456 ( .A(n23336), .ZN(n22499) );
  OAI21_X1 U22457 ( .B1(n22855), .B2(n21428), .A(n21427), .ZN(n22431) );
  XNOR2_X1 U22458 ( .A(n21430), .B(n21429), .ZN(n21435) );
  XNOR2_X1 U22459 ( .A(n21433), .B(n21432), .ZN(n21434) );
  XNOR2_X1 U22460 ( .A(n21434), .B(n21435), .ZN(n22852) );
  NAND2_X1 U22461 ( .A1(n22852), .A2(n22932), .ZN(n22498) );
  NOR2_X1 U22462 ( .A1(n24309), .A2(n22498), .ZN(n22432) );
  XNOR2_X1 U22464 ( .A(n21436), .B(n21510), .ZN(n21438) );
  XNOR2_X1 U22465 ( .A(n21728), .B(n21998), .ZN(n21437) );
  XNOR2_X1 U22466 ( .A(n21437), .B(n21438), .ZN(n21443) );
  XNOR2_X1 U22467 ( .A(n21583), .B(n25387), .ZN(n21441) );
  XNOR2_X1 U22468 ( .A(n21729), .B(n21942), .ZN(n21440) );
  XNOR2_X1 U22469 ( .A(n21441), .B(n21440), .ZN(n21442) );
  XNOR2_X1 U22470 ( .A(n25400), .B(n21445), .ZN(n21447) );
  XNOR2_X1 U22471 ( .A(n21750), .B(n2826), .ZN(n21446) );
  XNOR2_X1 U22472 ( .A(n21447), .B(n21446), .ZN(n21451) );
  XNOR2_X1 U22473 ( .A(n21449), .B(n21448), .ZN(n21450) );
  XNOR2_X1 U22474 ( .A(n21452), .B(n21660), .ZN(n21453) );
  XNOR2_X1 U22475 ( .A(n21454), .B(n21453), .ZN(n21459) );
  XNOR2_X1 U22476 ( .A(n24491), .B(n1724), .ZN(n21456) );
  XNOR2_X1 U22477 ( .A(n21457), .B(n21456), .ZN(n21458) );
  XNOR2_X1 U22478 ( .A(n21459), .B(n21458), .ZN(n22128) );
  XNOR2_X1 U22479 ( .A(n21461), .B(n21460), .ZN(n21465) );
  XNOR2_X1 U22480 ( .A(n21463), .B(n21462), .ZN(n21464) );
  XNOR2_X1 U22481 ( .A(n21465), .B(n21464), .ZN(n21467) );
  NAND2_X1 U22482 ( .A1(n22128), .A2(n21467), .ZN(n21466) );
  OAI21_X1 U22483 ( .B1(n22965), .B2(n22962), .A(n21466), .ZN(n22131) );
  INV_X1 U22484 ( .A(n22131), .ZN(n21490) );
  INV_X1 U22485 ( .A(n21466), .ZN(n21468) );
  NOR2_X1 U22486 ( .A1(n21468), .A2(n22969), .ZN(n21489) );
  XNOR2_X1 U22487 ( .A(n21676), .B(n21469), .ZN(n21470) );
  XNOR2_X1 U22488 ( .A(n21715), .B(n21470), .ZN(n21475) );
  XNOR2_X1 U22489 ( .A(n24962), .B(n4233), .ZN(n21473) );
  XNOR2_X1 U22490 ( .A(n21471), .B(n24899), .ZN(n21472) );
  XNOR2_X1 U22491 ( .A(n21472), .B(n21473), .ZN(n21474) );
  INV_X1 U22492 ( .A(n21959), .ZN(n21487) );
  XNOR2_X1 U22493 ( .A(n21479), .B(n21480), .ZN(n21485) );
  XNOR2_X1 U22494 ( .A(n21534), .B(n21559), .ZN(n21483) );
  XNOR2_X1 U22495 ( .A(n21481), .B(n2031), .ZN(n21482) );
  XNOR2_X1 U22496 ( .A(n21483), .B(n21482), .ZN(n21484) );
  NAND2_X1 U22498 ( .A1(n21487), .A2(n21486), .ZN(n21488) );
  INV_X1 U22499 ( .A(n23369), .ZN(n22741) );
  OR2_X1 U22500 ( .A1(n24515), .A2(n22741), .ZN(n21954) );
  XNOR2_X1 U22501 ( .A(n25470), .B(n25073), .ZN(n21627) );
  XNOR2_X1 U22502 ( .A(n21494), .B(n21627), .ZN(n21499) );
  XNOR2_X1 U22503 ( .A(n21495), .B(n23072), .ZN(n21497) );
  XNOR2_X1 U22504 ( .A(n21496), .B(n21497), .ZN(n21498) );
  XNOR2_X1 U22505 ( .A(n21498), .B(n21499), .ZN(n21540) );
  INV_X1 U22506 ( .A(n21540), .ZN(n22947) );
  XNOR2_X1 U22507 ( .A(n21974), .B(n21502), .ZN(n21504) );
  XNOR2_X1 U22508 ( .A(n21503), .B(n21504), .ZN(n21509) );
  XNOR2_X1 U22509 ( .A(n21506), .B(n21505), .ZN(n21507) );
  XNOR2_X1 U22510 ( .A(n21981), .B(n21507), .ZN(n21508) );
  XNOR2_X1 U22511 ( .A(n21509), .B(n21508), .ZN(n21872) );
  INV_X1 U22512 ( .A(n21872), .ZN(n22282) );
  XNOR2_X1 U22513 ( .A(n21510), .B(n1381), .ZN(n21513) );
  XNOR2_X1 U22514 ( .A(n21992), .B(n21511), .ZN(n21512) );
  XNOR2_X1 U22515 ( .A(n21512), .B(n21513), .ZN(n21519) );
  XNOR2_X1 U22517 ( .A(n21514), .B(n24624), .ZN(n21517) );
  XNOR2_X1 U22518 ( .A(n25091), .B(n21515), .ZN(n21516) );
  XNOR2_X1 U22519 ( .A(n21517), .B(n21516), .ZN(n21518) );
  INV_X1 U22520 ( .A(n22946), .ZN(n21530) );
  XNOR2_X1 U22521 ( .A(n21521), .B(n21520), .ZN(n22013) );
  XNOR2_X1 U22522 ( .A(n21523), .B(n21522), .ZN(n21524) );
  XNOR2_X1 U22523 ( .A(n22013), .B(n21524), .ZN(n21529) );
  XNOR2_X1 U22524 ( .A(n21525), .B(n853), .ZN(n21527) );
  XNOR2_X1 U22525 ( .A(n21713), .B(n21639), .ZN(n21526) );
  XNOR2_X1 U22526 ( .A(n21527), .B(n21526), .ZN(n21528) );
  XNOR2_X1 U22527 ( .A(n21532), .B(n21630), .ZN(n21535) );
  XNOR2_X1 U22528 ( .A(n21536), .B(n21633), .ZN(n21537) );
  XNOR2_X1 U22529 ( .A(n21539), .B(n21538), .ZN(n22948) );
  INV_X1 U22530 ( .A(n22948), .ZN(n22424) );
  XNOR2_X1 U22531 ( .A(n21541), .B(n21606), .ZN(n21542) );
  XNOR2_X1 U22532 ( .A(n21544), .B(n21543), .ZN(n21545) );
  OAI21_X1 U22533 ( .B1(n22948), .B2(n21548), .A(n21547), .ZN(n22435) );
  INV_X1 U22534 ( .A(n22435), .ZN(n21549) );
  XNOR2_X1 U22535 ( .A(n21550), .B(n21975), .ZN(n21552) );
  XNOR2_X1 U22536 ( .A(n21551), .B(n21552), .ZN(n21558) );
  INV_X1 U22537 ( .A(n21553), .ZN(n23589) );
  XNOR2_X1 U22538 ( .A(n21554), .B(n23589), .ZN(n21555) );
  XNOR2_X1 U22539 ( .A(n21556), .B(n21555), .ZN(n21557) );
  XNOR2_X1 U22542 ( .A(n21561), .B(n24306), .ZN(n21963) );
  XNOR2_X1 U22543 ( .A(n21562), .B(n21963), .ZN(n21566) );
  XNOR2_X1 U22544 ( .A(n24434), .B(n1856), .ZN(n21563) );
  XNOR2_X1 U22545 ( .A(n21564), .B(n21563), .ZN(n21565) );
  XNOR2_X1 U22546 ( .A(n21568), .B(n25385), .ZN(n21571) );
  XNOR2_X1 U22547 ( .A(n24996), .B(n2211), .ZN(n21570) );
  XNOR2_X1 U22548 ( .A(n21571), .B(n21570), .ZN(n21576) );
  XNOR2_X1 U22549 ( .A(n21572), .B(n21573), .ZN(n21989) );
  XNOR2_X1 U22550 ( .A(n21989), .B(n21574), .ZN(n21575) );
  XNOR2_X1 U22551 ( .A(n21575), .B(n21576), .ZN(n22953) );
  XNOR2_X1 U22553 ( .A(n21577), .B(n22385), .ZN(n21581) );
  XNOR2_X1 U22554 ( .A(n21579), .B(n21578), .ZN(n21580) );
  XNOR2_X1 U22555 ( .A(n21580), .B(n21581), .ZN(n21586) );
  XNOR2_X1 U22556 ( .A(n21582), .B(n21583), .ZN(n21993) );
  XNOR2_X1 U22557 ( .A(n21993), .B(n21584), .ZN(n21585) );
  XNOR2_X1 U22558 ( .A(n21586), .B(n21585), .ZN(n22952) );
  XNOR2_X1 U22559 ( .A(n21588), .B(n21587), .ZN(n21590) );
  XNOR2_X1 U22560 ( .A(n21590), .B(n21589), .ZN(n21595) );
  XNOR2_X1 U22561 ( .A(n21591), .B(n1831), .ZN(n21592) );
  XNOR2_X1 U22562 ( .A(n21593), .B(n21592), .ZN(n21594) );
  XNOR2_X1 U22563 ( .A(n21597), .B(n21596), .ZN(n22016) );
  XNOR2_X1 U22564 ( .A(n22016), .B(n21598), .ZN(n21605) );
  XNOR2_X1 U22565 ( .A(n21599), .B(n21600), .ZN(n21603) );
  XNOR2_X1 U22566 ( .A(n21601), .B(n21861), .ZN(n21602) );
  XNOR2_X1 U22567 ( .A(n21603), .B(n21602), .ZN(n21604) );
  NAND2_X1 U22568 ( .A1(n24885), .A2(n22954), .ZN(n21878) );
  XNOR2_X1 U22569 ( .A(n21687), .B(n21606), .ZN(n21610) );
  INV_X1 U22570 ( .A(n494), .ZN(n21607) );
  XNOR2_X1 U22571 ( .A(n21608), .B(n21607), .ZN(n21609) );
  XNOR2_X1 U22572 ( .A(n21610), .B(n21609), .ZN(n21613) );
  INV_X1 U22573 ( .A(n22027), .ZN(n22829) );
  XNOR2_X1 U22574 ( .A(n21614), .B(n21615), .ZN(n21620) );
  INV_X1 U22575 ( .A(n3062), .ZN(n22875) );
  XNOR2_X1 U22576 ( .A(n21616), .B(n22875), .ZN(n21617) );
  XNOR2_X1 U22577 ( .A(n21618), .B(n21617), .ZN(n21619) );
  XNOR2_X1 U22579 ( .A(n21622), .B(n21621), .ZN(n21625) );
  INV_X1 U22580 ( .A(n21623), .ZN(n23916) );
  XNOR2_X1 U22581 ( .A(n21693), .B(n23916), .ZN(n21624) );
  XNOR2_X1 U22582 ( .A(n21625), .B(n21624), .ZN(n21629) );
  XNOR2_X1 U22583 ( .A(n21626), .B(n21627), .ZN(n21628) );
  XNOR2_X1 U22584 ( .A(n21632), .B(n21631), .ZN(n21637) );
  XNOR2_X1 U22585 ( .A(n21633), .B(n23602), .ZN(n21634) );
  XNOR2_X1 U22586 ( .A(n21635), .B(n21634), .ZN(n21636) );
  INV_X1 U22587 ( .A(n22938), .ZN(n21644) );
  INV_X1 U22588 ( .A(n92), .ZN(n23322) );
  XNOR2_X1 U22589 ( .A(n21525), .B(n23322), .ZN(n21638) );
  XNOR2_X1 U22590 ( .A(n25065), .B(n21639), .ZN(n21641) );
  MUX2_X1 U22592 ( .A(n21644), .B(n25063), .S(n24932), .Z(n21656) );
  XNOR2_X1 U22593 ( .A(n21645), .B(n21646), .ZN(n21652) );
  XNOR2_X1 U22594 ( .A(n21647), .B(n1777), .ZN(n21650) );
  XNOR2_X1 U22595 ( .A(n21651), .B(n21652), .ZN(n22722) );
  INV_X1 U22596 ( .A(n22722), .ZN(n22941) );
  NAND2_X1 U22598 ( .A1(n22832), .A2(n22939), .ZN(n21653) );
  MUX2_X1 U22599 ( .A(n21654), .B(n21653), .S(n22027), .Z(n21655) );
  NAND2_X1 U22600 ( .A1(n23374), .A2(n23379), .ZN(n22430) );
  XNOR2_X1 U22601 ( .A(n25498), .B(n21658), .ZN(n21661) );
  INV_X1 U22602 ( .A(n21662), .ZN(n23763) );
  XNOR2_X1 U22603 ( .A(n21027), .B(n23763), .ZN(n21663) );
  XNOR2_X1 U22604 ( .A(n21664), .B(n24898), .ZN(n21666) );
  XNOR2_X1 U22605 ( .A(n21669), .B(n21668), .ZN(n21674) );
  XNOR2_X1 U22606 ( .A(n21670), .B(n16574), .ZN(n21672) );
  XNOR2_X1 U22607 ( .A(n21671), .B(n21672), .ZN(n21673) );
  XNOR2_X1 U22609 ( .A(n21675), .B(n1789), .ZN(n21677) );
  XNOR2_X1 U22610 ( .A(n21677), .B(n21676), .ZN(n21681) );
  XNOR2_X1 U22611 ( .A(n21679), .B(n21678), .ZN(n21680) );
  XNOR2_X1 U22612 ( .A(n21681), .B(n21680), .ZN(n21682) );
  XNOR2_X1 U22613 ( .A(n21685), .B(n21684), .ZN(n21691) );
  XNOR2_X1 U22614 ( .A(n21686), .B(n5433), .ZN(n21688) );
  XNOR2_X1 U22615 ( .A(n21691), .B(n21690), .ZN(n22483) );
  OAI22_X1 U22617 ( .A1(n21692), .A2(n22901), .B1(n22842), .B2(n25569), .ZN(
        n21710) );
  XNOR2_X1 U22618 ( .A(n21693), .B(n447), .ZN(n21695) );
  NAND2_X1 U22619 ( .A1(n25569), .A2(n22900), .ZN(n21709) );
  XNOR2_X1 U22620 ( .A(n25202), .B(n21699), .ZN(n21702) );
  XNOR2_X1 U22621 ( .A(n21702), .B(n21701), .ZN(n21708) );
  INV_X1 U22622 ( .A(n21703), .ZN(n23330) );
  XNOR2_X1 U22623 ( .A(n21704), .B(n23330), .ZN(n21705) );
  XNOR2_X1 U22624 ( .A(n21706), .B(n21705), .ZN(n21707) );
  XNOR2_X1 U22625 ( .A(n21708), .B(n21707), .ZN(n22905) );
  INV_X1 U22626 ( .A(n22905), .ZN(n22907) );
  INV_X1 U22627 ( .A(n22070), .ZN(n21712) );
  XNOR2_X1 U22629 ( .A(n21713), .B(n3118), .ZN(n21714) );
  XNOR2_X1 U22630 ( .A(n21715), .B(n21714), .ZN(n21719) );
  XNOR2_X1 U22631 ( .A(n21717), .B(n21716), .ZN(n21718) );
  XNOR2_X2 U22632 ( .A(n21718), .B(n21719), .ZN(n23016) );
  XNOR2_X1 U22633 ( .A(n21721), .B(n21720), .ZN(n21722) );
  XNOR2_X1 U22634 ( .A(n20727), .B(n3901), .ZN(n21724) );
  XNOR2_X1 U22635 ( .A(n21726), .B(n21727), .ZN(n21733) );
  XNOR2_X1 U22636 ( .A(n24985), .B(n21728), .ZN(n21731) );
  XNOR2_X1 U22637 ( .A(n21729), .B(n22382), .ZN(n21730) );
  XNOR2_X1 U22638 ( .A(n21731), .B(n21730), .ZN(n21732) );
  XNOR2_X1 U22639 ( .A(n21733), .B(n21732), .ZN(n23458) );
  NAND2_X1 U22640 ( .A1(n23016), .A2(n23458), .ZN(n21741) );
  XNOR2_X1 U22641 ( .A(n21736), .B(n2747), .ZN(n21737) );
  XNOR2_X1 U22642 ( .A(n21738), .B(n21739), .ZN(n21740) );
  MUX2_X1 U22643 ( .A(n22914), .B(n21741), .S(n24877), .Z(n21758) );
  XNOR2_X1 U22644 ( .A(n1326), .B(n21742), .ZN(n21744) );
  XNOR2_X1 U22645 ( .A(n21745), .B(n21744), .ZN(n21746) );
  XNOR2_X1 U22646 ( .A(n21747), .B(n21746), .ZN(n21749) );
  XNOR2_X2 U22647 ( .A(n21749), .B(n21748), .ZN(n23464) );
  INV_X1 U22648 ( .A(n23016), .ZN(n23460) );
  XNOR2_X1 U22649 ( .A(n21751), .B(n21750), .ZN(n21753) );
  XNOR2_X1 U22650 ( .A(n21753), .B(n21752), .ZN(n21757) );
  XNOR2_X1 U22651 ( .A(n21754), .B(n21755), .ZN(n21756) );
  XNOR2_X1 U22652 ( .A(n21756), .B(n21757), .ZN(n23015) );
  NAND2_X1 U22653 ( .A1(n24611), .A2(n23595), .ZN(n22639) );
  INV_X1 U22654 ( .A(n23575), .ZN(n22079) );
  INV_X1 U22655 ( .A(n21759), .ZN(n23576) );
  AOI21_X1 U22656 ( .B1(n22079), .B2(n23576), .A(n22176), .ZN(n21760) );
  INV_X1 U22657 ( .A(n23566), .ZN(n21763) );
  INV_X1 U22658 ( .A(n22922), .ZN(n22107) );
  INV_X1 U22659 ( .A(n22209), .ZN(n21767) );
  OAI21_X1 U22660 ( .B1(n24333), .B2(n22208), .A(n21767), .ZN(n21764) );
  NOR2_X1 U22661 ( .A1(n21765), .A2(n21764), .ZN(n21771) );
  NOR2_X1 U22662 ( .A1(n22159), .A2(n22206), .ZN(n21768) );
  NOR2_X1 U22663 ( .A1(n21768), .A2(n21767), .ZN(n21770) );
  NAND2_X1 U22664 ( .A1(n22159), .A2(n24333), .ZN(n21769) );
  INV_X1 U22665 ( .A(n23596), .ZN(n22633) );
  INV_X1 U22666 ( .A(n22889), .ZN(n22496) );
  AOI22_X1 U22668 ( .A1(n21772), .A2(n22887), .B1(n22729), .B2(n22890), .ZN(
        n21773) );
  NAND3_X1 U22669 ( .A1(n24390), .A2(n22633), .A3(n24901), .ZN(n21776) );
  NOR2_X1 U22670 ( .A1(n24390), .A2(n24397), .ZN(n21947) );
  NAND2_X1 U22671 ( .A1(n21947), .A2(n23596), .ZN(n21775) );
  NAND4_X1 U22672 ( .A1(n22639), .A2(n21777), .A3(n21776), .A4(n21775), .ZN(
        n21779) );
  INV_X1 U22673 ( .A(n1801), .ZN(n21778) );
  XNOR2_X1 U22674 ( .A(n21779), .B(n21778), .ZN(Ciphertext[114]) );
  AOI21_X1 U22676 ( .B1(n24114), .B2(n21838), .A(n21839), .ZN(n21785) );
  NOR2_X1 U22677 ( .A1(n22355), .A2(n22354), .ZN(n21781) );
  NAND2_X1 U22678 ( .A1(n21781), .A2(n22356), .ZN(n21784) );
  NOR2_X1 U22679 ( .A1(n21782), .A2(n21839), .ZN(n21845) );
  NAND2_X1 U22681 ( .A1(n21845), .A2(n25082), .ZN(n21783) );
  INV_X1 U22683 ( .A(n23757), .ZN(n21800) );
  INV_X1 U22686 ( .A(n22244), .ZN(n21815) );
  NOR2_X1 U22689 ( .A1(n21800), .A2(n23769), .ZN(n21795) );
  MUX2_X1 U22690 ( .A(n25461), .B(n22217), .S(n22221), .Z(n21790) );
  NAND2_X1 U22691 ( .A1(n21829), .A2(n22222), .ZN(n21789) );
  NOR2_X1 U22692 ( .A1(n25051), .A2(n24921), .ZN(n23771) );
  NAND2_X1 U22693 ( .A1(n22231), .A2(n22226), .ZN(n21792) );
  NOR2_X1 U22694 ( .A1(n22233), .A2(n22226), .ZN(n21793) );
  OAI21_X1 U22695 ( .B1(n21795), .B2(n23771), .A(n23779), .ZN(n21809) );
  INV_X1 U22696 ( .A(n23752), .ZN(n21798) );
  NAND2_X1 U22697 ( .A1(n22522), .A2(n22255), .ZN(n21797) );
  NAND2_X1 U22699 ( .A1(n22521), .A2(n4373), .ZN(n21796) );
  NAND3_X1 U22700 ( .A1(n21798), .A2(n21797), .A3(n21796), .ZN(n21799) );
  NAND3_X1 U22701 ( .A1(n25051), .A2(n21800), .A3(n21799), .ZN(n21808) );
  NOR2_X1 U22702 ( .A1(n22079), .A2(n22197), .ZN(n21801) );
  NOR2_X1 U22703 ( .A1(n21802), .A2(n21801), .ZN(n21805) );
  NOR2_X1 U22704 ( .A1(n22079), .A2(n24369), .ZN(n21803) );
  NAND2_X1 U22705 ( .A1(n23768), .A2(n24921), .ZN(n21806) );
  NAND3_X1 U22706 ( .A1(n21809), .A2(n21808), .A3(n21807), .ZN(n21811) );
  INV_X1 U22707 ( .A(n1777), .ZN(n21810) );
  XNOR2_X1 U22708 ( .A(n21811), .B(n21810), .ZN(Ciphertext[146]) );
  NOR2_X1 U22709 ( .A1(n22243), .A2(n22239), .ZN(n21814) );
  INV_X1 U22710 ( .A(n22184), .ZN(n21813) );
  NAND2_X1 U22711 ( .A1(n21815), .A2(n22243), .ZN(n23001) );
  NOR2_X1 U22712 ( .A1(n21848), .A2(n21816), .ZN(n22348) );
  NAND3_X1 U22714 ( .A1(n21848), .A2(n22688), .A3(n22685), .ZN(n21820) );
  NAND2_X1 U22715 ( .A1(n21848), .A2(n21817), .ZN(n21818) );
  NOR2_X1 U22716 ( .A1(n24468), .A2(n21841), .ZN(n21824) );
  NOR2_X1 U22717 ( .A1(n332), .A2(n21825), .ZN(n21823) );
  MUX2_X1 U22718 ( .A(n21824), .B(n21823), .S(n21822), .Z(n21827) );
  NAND2_X1 U22719 ( .A1(n24362), .A2(n21841), .ZN(n21826) );
  NOR2_X1 U22721 ( .A1(n22214), .A2(n22221), .ZN(n21832) );
  NAND2_X1 U22722 ( .A1(n22222), .A2(n24918), .ZN(n21831) );
  NAND2_X1 U22723 ( .A1(n22216), .A2(n22221), .ZN(n22218) );
  OAI211_X1 U22724 ( .C1(n21832), .C2(n21831), .A(n22218), .B(n21830), .ZN(
        n23799) );
  NAND3_X1 U22725 ( .A1(n24307), .A2(n24895), .A3(n24920), .ZN(n21833) );
  NAND2_X1 U22726 ( .A1(n22233), .A2(n22225), .ZN(n21834) );
  MUX2_X1 U22729 ( .A(n21845), .B(n22356), .S(n21844), .Z(n23893) );
  NAND2_X1 U22730 ( .A1(n22355), .A2(n22354), .ZN(n21846) );
  AND2_X1 U22731 ( .A1(n22359), .A2(n21846), .ZN(n23892) );
  NOR2_X2 U22732 ( .A1(n23893), .A2(n23892), .ZN(n23904) );
  MUX2_X1 U22733 ( .A(n22689), .B(n22685), .S(n22688), .Z(n21849) );
  MUX2_X2 U22734 ( .A(n21850), .B(n21849), .S(n22687), .Z(n23905) );
  INV_X1 U22737 ( .A(n21866), .ZN(n21851) );
  NAND2_X1 U22738 ( .A1(n21851), .A2(n21861), .ZN(n21870) );
  NAND2_X1 U22739 ( .A1(n22813), .A2(n4469), .ZN(n21852) );
  AOI22_X1 U22741 ( .A1(n25439), .A2(n22677), .B1(n23998), .B2(n25414), .ZN(
        n22598) );
  INV_X1 U22742 ( .A(n23995), .ZN(n22596) );
  OAI21_X1 U22743 ( .B1(n22596), .B2(n24439), .A(n23998), .ZN(n21853) );
  INV_X1 U22744 ( .A(n23994), .ZN(n22678) );
  NAND2_X1 U22745 ( .A1(n21853), .A2(n22678), .ZN(n21854) );
  AOI21_X1 U22746 ( .B1(n23906), .B2(n23889), .A(n23905), .ZN(n21869) );
  AND2_X1 U22747 ( .A1(n21856), .A2(n22679), .ZN(n21858) );
  NOR2_X1 U22748 ( .A1(n22769), .A2(n22770), .ZN(n21857) );
  MUX2_X1 U22749 ( .A(n21858), .B(n21857), .S(n22774), .Z(n23891) );
  NOR2_X1 U22750 ( .A1(n23890), .A2(n16), .ZN(n21860) );
  NAND2_X1 U22751 ( .A1(n23879), .A2(n23889), .ZN(n21859) );
  OAI211_X1 U22752 ( .C1(n23905), .C2(n23879), .A(n21860), .B(n21859), .ZN(
        n21868) );
  NOR2_X1 U22753 ( .A1(n23890), .A2(n23889), .ZN(n21862) );
  AOI21_X1 U22754 ( .B1(n21862), .B2(n23879), .A(n21861), .ZN(n21865) );
  NAND2_X1 U22756 ( .A1(n23909), .A2(n23903), .ZN(n21864) );
  INV_X1 U22759 ( .A(n22852), .ZN(n22933) );
  NAND2_X1 U22761 ( .A1(n22426), .A2(n22947), .ZN(n21874) );
  NAND3_X1 U22762 ( .A1(n22422), .A2(n22420), .A3(n22421), .ZN(n21873) );
  OAI21_X1 U22763 ( .B1(n21874), .B2(n22948), .A(n21873), .ZN(n21877) );
  NAND2_X1 U22765 ( .A1(n23317), .A2(n23326), .ZN(n22629) );
  INV_X1 U22766 ( .A(n21878), .ZN(n21882) );
  OAI21_X1 U22767 ( .B1(n22954), .B2(n22953), .A(n22033), .ZN(n21881) );
  NOR2_X1 U22768 ( .A1(n24885), .A2(n22033), .ZN(n22394) );
  AOI21_X1 U22769 ( .B1(n22394), .B2(n24922), .A(n21879), .ZN(n21880) );
  OAI21_X1 U22770 ( .B1(n21882), .B2(n21881), .A(n21880), .ZN(n23324) );
  INV_X1 U22771 ( .A(n23324), .ZN(n23313) );
  OR2_X1 U22772 ( .A1(n22629), .A2(n23313), .ZN(n21897) );
  INV_X1 U22773 ( .A(n22397), .ZN(n21883) );
  NAND2_X1 U22774 ( .A1(n22398), .A2(n22265), .ZN(n21887) );
  INV_X1 U22775 ( .A(n25381), .ZN(n21884) );
  OAI21_X1 U22776 ( .B1(n21885), .B2(n22397), .A(n21884), .ZN(n21886) );
  NOR2_X1 U22777 ( .A1(n22397), .A2(n22134), .ZN(n22268) );
  INV_X1 U22778 ( .A(n21888), .ZN(n22396) );
  NAND2_X1 U22779 ( .A1(n22968), .A2(n21467), .ZN(n21956) );
  NAND3_X1 U22780 ( .A1(n22962), .A2(n21476), .A3(n22969), .ZN(n21890) );
  NAND2_X1 U22781 ( .A1(n24411), .A2(n22965), .ZN(n21889) );
  NAND3_X1 U22782 ( .A1(n23327), .A2(n23318), .A3(n4108), .ZN(n21896) );
  INV_X1 U22783 ( .A(n22975), .ZN(n21892) );
  NOR2_X1 U22784 ( .A1(n21892), .A2(n24881), .ZN(n21893) );
  NOR3_X1 U22785 ( .A1(n21893), .A2(n22977), .A3(n3213), .ZN(n21894) );
  INV_X1 U22786 ( .A(n2039), .ZN(n21898) );
  XNOR2_X1 U22787 ( .A(n21899), .B(n21898), .ZN(Ciphertext[63]) );
  INV_X1 U22788 ( .A(n23805), .ZN(n23788) );
  NAND2_X1 U22789 ( .A1(n23787), .A2(n21902), .ZN(n21901) );
  OAI211_X1 U22790 ( .C1(n23805), .C2(n21901), .A(Key[33]), .B(n21900), .ZN(
        n21906) );
  INV_X1 U22791 ( .A(Key[33]), .ZN(n21903) );
  NAND2_X1 U22792 ( .A1(n21907), .A2(n21903), .ZN(n21904) );
  OAI211_X1 U22793 ( .C1(n21907), .C2(n21906), .A(n21905), .B(n21904), .ZN(
        Ciphertext[153]) );
  NAND2_X1 U22794 ( .A1(n21909), .A2(n24415), .ZN(n21913) );
  AND2_X1 U22795 ( .A1(n22334), .A2(n22139), .ZN(n22273) );
  NOR2_X1 U22796 ( .A1(n22335), .A2(n21910), .ZN(n22142) );
  NAND2_X1 U22797 ( .A1(n22142), .A2(n22274), .ZN(n21912) );
  NAND3_X1 U22798 ( .A1(n22333), .A2(n22139), .A3(n21910), .ZN(n21911) );
  OR2_X1 U22799 ( .A1(n21914), .A2(n22134), .ZN(n21916) );
  AND2_X1 U22800 ( .A1(n22396), .A2(n22134), .ZN(n22404) );
  NOR2_X1 U22802 ( .A1(n21918), .A2(n24311), .ZN(n21919) );
  AND2_X1 U22803 ( .A1(n25066), .A2(n21921), .ZN(n21922) );
  OAI21_X1 U22805 ( .B1(n24043), .B2(n22448), .A(n274), .ZN(n21926) );
  INV_X1 U22806 ( .A(n22448), .ZN(n21924) );
  OAI21_X1 U22808 ( .B1(n21929), .B2(n22464), .A(n21928), .ZN(n21933) );
  INV_X1 U22809 ( .A(n22562), .ZN(n22341) );
  INV_X1 U22810 ( .A(n22407), .ZN(n22567) );
  NOR2_X1 U22811 ( .A1(n22341), .A2(n22567), .ZN(n21935) );
  NOR2_X1 U22812 ( .A1(n333), .A2(n22409), .ZN(n22411) );
  INV_X1 U22813 ( .A(n22411), .ZN(n21937) );
  INV_X1 U22815 ( .A(n21946), .ZN(n21940) );
  NAND3_X1 U22816 ( .A1(n23595), .A2(n24390), .A3(n1328), .ZN(n21939) );
  OAI211_X1 U22817 ( .C1(n22633), .C2(n21940), .A(n21942), .B(n21939), .ZN(
        n21952) );
  INV_X1 U22818 ( .A(n23592), .ZN(n21941) );
  NAND2_X1 U22819 ( .A1(n24372), .A2(n23566), .ZN(n22634) );
  OR2_X1 U22820 ( .A1(n21943), .A2(n21942), .ZN(n21950) );
  AOI21_X1 U22821 ( .B1(n22633), .B2(n21946), .A(n21945), .ZN(n21948) );
  INV_X1 U22822 ( .A(n21947), .ZN(n22632) );
  OAI211_X1 U22823 ( .C1(n24611), .C2(n22634), .A(n21948), .B(n22632), .ZN(
        n21949) );
  INV_X1 U22824 ( .A(n23374), .ZN(n23370) );
  AOI21_X1 U22825 ( .B1(n24515), .B2(n24911), .A(n24404), .ZN(n21953) );
  NAND2_X1 U22826 ( .A1(n21954), .A2(n21953), .ZN(n21955) );
  NAND2_X1 U22827 ( .A1(n24515), .A2(n22987), .ZN(n22744) );
  OAI21_X1 U22828 ( .B1(n22966), .B2(n22969), .A(n21956), .ZN(n21957) );
  INV_X1 U22829 ( .A(n21957), .ZN(n21962) );
  NAND2_X1 U22830 ( .A1(n22962), .A2(n24411), .ZN(n21958) );
  NOR2_X1 U22831 ( .A1(n334), .A2(n24411), .ZN(n21960) );
  AOI21_X2 U22832 ( .B1(n21962), .B2(n21961), .A(n21960), .ZN(n23396) );
  INV_X1 U22833 ( .A(n23396), .ZN(n22032) );
  INV_X1 U22834 ( .A(n21963), .ZN(n21969) );
  XNOR2_X1 U22835 ( .A(n21965), .B(n21964), .ZN(n21966) );
  XNOR2_X1 U22836 ( .A(n21966), .B(n21967), .ZN(n21968) );
  XNOR2_X1 U22837 ( .A(n21968), .B(n21969), .ZN(n21973) );
  XNOR2_X1 U22838 ( .A(n21971), .B(n21970), .ZN(n21972) );
  XNOR2_X1 U22839 ( .A(n21974), .B(n924), .ZN(n21976) );
  XNOR2_X1 U22840 ( .A(n21976), .B(n21975), .ZN(n21978) );
  XNOR2_X1 U22841 ( .A(n21977), .B(n21978), .ZN(n21984) );
  XNOR2_X1 U22842 ( .A(n21979), .B(n21980), .ZN(n21982) );
  XNOR2_X1 U22843 ( .A(n21982), .B(n21981), .ZN(n21983) );
  XNOR2_X1 U22845 ( .A(n21986), .B(n21987), .ZN(n21991) );
  XNOR2_X1 U22846 ( .A(n20727), .B(n3900), .ZN(n21988) );
  XNOR2_X1 U22847 ( .A(n21989), .B(n21988), .ZN(n21990) );
  XNOR2_X1 U22851 ( .A(n25091), .B(n21996), .ZN(n22000) );
  XNOR2_X1 U22852 ( .A(n21998), .B(n1863), .ZN(n21999) );
  XNOR2_X1 U22853 ( .A(n22000), .B(n21999), .ZN(n22001) );
  XNOR2_X1 U22854 ( .A(n22002), .B(n22001), .ZN(n22836) );
  XNOR2_X1 U22855 ( .A(n22004), .B(n22003), .ZN(n22011) );
  INV_X1 U22856 ( .A(n1874), .ZN(n23922) );
  XNOR2_X1 U22857 ( .A(n22005), .B(n23922), .ZN(n22009) );
  XNOR2_X1 U22858 ( .A(n22007), .B(n22006), .ZN(n22008) );
  XNOR2_X1 U22859 ( .A(n22008), .B(n22009), .ZN(n22010) );
  XNOR2_X1 U22860 ( .A(n22011), .B(n22010), .ZN(n22837) );
  OAI22_X1 U22861 ( .A1(n22838), .A2(n22893), .B1(n22836), .B2(n22837), .ZN(
        n22896) );
  XNOR2_X1 U22862 ( .A(n22012), .B(n22013), .ZN(n22018) );
  INV_X1 U22863 ( .A(n2772), .ZN(n23775) );
  XNOR2_X1 U22864 ( .A(n22014), .B(n23775), .ZN(n22015) );
  XNOR2_X1 U22865 ( .A(n22016), .B(n22015), .ZN(n22017) );
  INV_X1 U22866 ( .A(n22837), .ZN(n22841) );
  OAI21_X1 U22867 ( .B1(n25041), .B2(n22836), .A(n22841), .ZN(n22019) );
  NAND3_X1 U22868 ( .A1(n25382), .A2(n22905), .A3(n22842), .ZN(n22025) );
  INV_X1 U22869 ( .A(n22842), .ZN(n22906) );
  NAND3_X1 U22870 ( .A1(n22906), .A2(n25569), .A3(n22901), .ZN(n22024) );
  NOR2_X1 U22871 ( .A1(n22901), .A2(n22483), .ZN(n22903) );
  NAND2_X1 U22872 ( .A1(n22903), .A2(n22904), .ZN(n22023) );
  NOR2_X1 U22873 ( .A1(n25569), .A2(n22900), .ZN(n22021) );
  NAND2_X1 U22874 ( .A1(n22021), .A2(n22906), .ZN(n22022) );
  INV_X1 U22875 ( .A(n22940), .ZN(n22936) );
  OAI21_X1 U22876 ( .B1(n22936), .B2(n22938), .A(n22832), .ZN(n22030) );
  NOR2_X1 U22877 ( .A1(n22940), .A2(n22722), .ZN(n22029) );
  NAND2_X1 U22878 ( .A1(n22029), .A2(n22939), .ZN(n22028) );
  INV_X1 U22880 ( .A(n24449), .ZN(n22031) );
  AOI22_X1 U22881 ( .A1(n24884), .A2(n22953), .B1(n22952), .B2(n22033), .ZN(
        n22393) );
  NAND3_X1 U22882 ( .A1(n22034), .A2(n24922), .A3(n22954), .ZN(n22035) );
  INV_X1 U22883 ( .A(n23394), .ZN(n22036) );
  NOR3_X1 U22884 ( .A1(n24933), .A2(n22036), .A3(n24465), .ZN(n22040) );
  MUX2_X1 U22885 ( .A(n24341), .B(n22852), .S(n23332), .Z(n22038) );
  MUX2_X1 U22886 ( .A(n23334), .B(n25081), .S(n22501), .Z(n22037) );
  NOR3_X1 U22888 ( .A1(n324), .A2(n23392), .A3(n24465), .ZN(n22039) );
  NOR3_X1 U22889 ( .A1(n22041), .A2(n22040), .A3(n22039), .ZN(n22042) );
  XNOR2_X1 U22890 ( .A(n22042), .B(n677), .ZN(Ciphertext[78]) );
  NAND2_X1 U22891 ( .A1(n22044), .A2(n23805), .ZN(n22048) );
  NOR3_X1 U22892 ( .A1(n22046), .A2(n23002), .A3(n22045), .ZN(n22047) );
  OAI21_X1 U22893 ( .B1(n21829), .B2(n22217), .A(n25461), .ZN(n22054) );
  NAND2_X1 U22894 ( .A1(n22216), .A2(n22214), .ZN(n22050) );
  NAND2_X1 U22895 ( .A1(n22050), .A2(n2817), .ZN(n22052) );
  NOR2_X1 U22898 ( .A1(n22239), .A2(n22059), .ZN(n22060) );
  AOI22_X1 U22899 ( .A1(n22184), .A2(n1336), .B1(n22243), .B2(n22060), .ZN(
        n22061) );
  OAI21_X1 U22900 ( .B1(n22063), .B2(n22062), .A(n22061), .ZN(n23697) );
  INV_X1 U22901 ( .A(n22212), .ZN(n22068) );
  AOI22_X2 U22902 ( .A1(n22067), .A2(n22068), .B1(n22065), .B2(n22066), .ZN(
        n23720) );
  INV_X1 U22903 ( .A(n22916), .ZN(n22170) );
  NOR2_X1 U22905 ( .A1(n24674), .A2(n22166), .ZN(n22071) );
  NOR2_X2 U22909 ( .A1(n22075), .A2(n22074), .ZN(n23712) );
  NOR2_X1 U22910 ( .A1(n23712), .A2(n23720), .ZN(n23724) );
  INV_X1 U22911 ( .A(n3125), .ZN(n22082) );
  AOI21_X1 U22912 ( .B1(n23724), .B2(n22082), .A(n23714), .ZN(n22077) );
  OR2_X1 U22913 ( .A1(n23724), .A2(n22082), .ZN(n22076) );
  OAI211_X1 U22914 ( .C1(n23696), .C2(n22148), .A(n22077), .B(n22076), .ZN(
        n22085) );
  AND2_X1 U22916 ( .A1(n23571), .A2(n22200), .ZN(n22081) );
  NAND4_X1 U22917 ( .A1(n24374), .A2(n22082), .A3(n22148), .A4(n23714), .ZN(
        n22083) );
  INV_X1 U22918 ( .A(n23712), .ZN(n23719) );
  OAI21_X1 U22919 ( .B1(n23723), .B2(n23720), .A(n23721), .ZN(n22086) );
  OAI21_X1 U22920 ( .B1(n23719), .B2(n24381), .A(n22086), .ZN(n22091) );
  NAND2_X1 U22921 ( .A1(n23714), .A2(n22089), .ZN(n22087) );
  AOI21_X1 U22922 ( .B1(n23723), .B2(n24381), .A(n22087), .ZN(n22088) );
  OAI21_X1 U22923 ( .B1(n24374), .B2(n23723), .A(n22088), .ZN(n22090) );
  NAND2_X1 U22925 ( .A1(n22496), .A2(n22093), .ZN(n22099) );
  NOR2_X1 U22926 ( .A1(n22890), .A2(n327), .ZN(n22097) );
  INV_X1 U22927 ( .A(n22887), .ZN(n22494) );
  OAI21_X1 U22928 ( .B1(n25375), .B2(n22494), .A(n22095), .ZN(n22096) );
  NAND2_X1 U22929 ( .A1(n24877), .A2(n23014), .ZN(n22100) );
  AND3_X1 U22931 ( .A1(n22100), .A2(n24364), .A3(n23016), .ZN(n22102) );
  AND2_X1 U22932 ( .A1(n23015), .A2(n23458), .ZN(n22862) );
  AND2_X1 U22933 ( .A1(n23014), .A2(n22862), .ZN(n22101) );
  NOR3_X2 U22934 ( .A1(n22102), .A2(n22863), .A3(n22101), .ZN(n23555) );
  INV_X1 U22935 ( .A(n22893), .ZN(n22834) );
  NAND2_X1 U22936 ( .A1(n22834), .A2(n25438), .ZN(n22897) );
  NAND2_X1 U22937 ( .A1(n22717), .A2(n25041), .ZN(n22103) );
  AOI21_X1 U22938 ( .B1(n22897), .B2(n22103), .A(n22835), .ZN(n22106) );
  NAND2_X1 U22939 ( .A1(n22835), .A2(n22834), .ZN(n22104) );
  AOI21_X1 U22940 ( .B1(n22104), .B2(n22837), .A(n25041), .ZN(n22105) );
  NOR2_X1 U22941 ( .A1(n22106), .A2(n22105), .ZN(n23547) );
  OAI22_X1 U22942 ( .A1(n323), .A2(n23554), .B1(n23555), .B2(n23547), .ZN(
        n22701) );
  INV_X1 U22943 ( .A(n22926), .ZN(n22929) );
  NAND2_X1 U22945 ( .A1(n25479), .A2(n22188), .ZN(n22109) );
  NAND3_X1 U22946 ( .A1(n25070), .A2(n22107), .A3(n22927), .ZN(n22108) );
  AND2_X1 U22947 ( .A1(n24379), .A2(n22927), .ZN(n22110) );
  INV_X1 U22948 ( .A(n22110), .ZN(n22111) );
  AND2_X1 U22949 ( .A1(n25071), .A2(n23555), .ZN(n23551) );
  MUX2_X1 U22950 ( .A(n21712), .B(n22166), .S(n22916), .Z(n22114) );
  INV_X1 U22951 ( .A(n22918), .ZN(n22113) );
  NAND2_X1 U22952 ( .A1(n22114), .A2(n22113), .ZN(n22120) );
  OR2_X1 U22953 ( .A1(n22115), .A2(n22917), .ZN(n22119) );
  INV_X1 U22954 ( .A(n22116), .ZN(n22117) );
  NAND2_X1 U22955 ( .A1(n323), .A2(n23537), .ZN(n22121) );
  AOI22_X1 U22956 ( .A1(n22701), .A2(n23544), .B1(n23551), .B2(n22121), .ZN(
        n22122) );
  XNOR2_X1 U22957 ( .A(n22122), .B(n1767), .ZN(Ciphertext[109]) );
  NOR3_X1 U22958 ( .A1(n22948), .A2(n22426), .A3(n22422), .ZN(n22124) );
  NOR3_X1 U22959 ( .A1(n22282), .A2(n22421), .A3(n22946), .ZN(n22123) );
  NOR2_X1 U22960 ( .A1(n22124), .A2(n22123), .ZN(n22127) );
  AOI21_X1 U22961 ( .B1(n22963), .B2(n22129), .A(n22128), .ZN(n22130) );
  NOR2_X1 U22963 ( .A1(n22536), .A2(n24907), .ZN(n22145) );
  INV_X1 U22964 ( .A(n22134), .ZN(n22261) );
  NAND2_X1 U22966 ( .A1(n22337), .A2(n22138), .ZN(n22140) );
  OAI21_X1 U22967 ( .B1(n5767), .B2(n22337), .A(n22140), .ZN(n22143) );
  AOI21_X1 U22968 ( .B1(n22145), .B2(n24360), .A(n22144), .ZN(n22146) );
  XNOR2_X1 U22969 ( .A(n22146), .B(n2145), .ZN(Ciphertext[49]) );
  NAND3_X1 U22970 ( .A1(n23712), .A2(n24381), .A3(n23716), .ZN(n22149) );
  OAI21_X1 U22973 ( .B1(n22159), .B2(n22156), .A(n22155), .ZN(n22157) );
  INV_X1 U22974 ( .A(n25485), .ZN(n22158) );
  NAND2_X1 U22976 ( .A1(n22218), .A2(n22162), .ZN(n22165) );
  OAI21_X1 U22977 ( .B1(n22222), .B2(n22217), .A(n21829), .ZN(n22163) );
  AND2_X1 U22978 ( .A1(n25461), .A2(n22163), .ZN(n22164) );
  INV_X1 U22980 ( .A(n22166), .ZN(n22919) );
  NOR2_X1 U22981 ( .A1(n22919), .A2(n24902), .ZN(n22168) );
  NAND2_X1 U22982 ( .A1(n22169), .A2(n22168), .ZN(n22172) );
  NAND2_X1 U22983 ( .A1(n23576), .A2(n22175), .ZN(n22173) );
  OAI21_X1 U22984 ( .B1(n23576), .B2(n24396), .A(n22173), .ZN(n22174) );
  INV_X1 U22985 ( .A(n22175), .ZN(n22199) );
  NAND3_X1 U22986 ( .A1(n22199), .A2(n1323), .A3(n4360), .ZN(n22177) );
  NOR2_X1 U22987 ( .A1(n22240), .A2(n22180), .ZN(n22182) );
  OR2_X1 U22988 ( .A1(n1336), .A2(n22244), .ZN(n22185) );
  OAI21_X1 U22991 ( .B1(n23686), .B2(n22186), .A(n23658), .ZN(n22194) );
  INV_X1 U22993 ( .A(n25026), .ZN(n23678) );
  OAI21_X1 U22995 ( .B1(n22926), .B2(n25479), .A(n22188), .ZN(n22191) );
  AOI21_X2 U22996 ( .B1(n22192), .B2(n22191), .A(n22190), .ZN(n23690) );
  INV_X1 U22997 ( .A(n1855), .ZN(n22195) );
  NAND2_X1 U22999 ( .A1(n24396), .A2(n22197), .ZN(n22202) );
  OAI21_X1 U23000 ( .B1(n22199), .B2(n22202), .A(n22198), .ZN(n22204) );
  OAI22_X1 U23001 ( .A1(n24369), .A2(n22202), .B1(n22201), .B2(n22175), .ZN(
        n22203) );
  NAND2_X1 U23003 ( .A1(n22208), .A2(n22206), .ZN(n22207) );
  OAI21_X1 U23004 ( .B1(n22209), .B2(n25018), .A(n22207), .ZN(n22210) );
  NAND2_X1 U23006 ( .A1(n22214), .A2(n22221), .ZN(n22215) );
  OAI22_X1 U23007 ( .A1(n22218), .A2(n24918), .B1(n22216), .B2(n22215), .ZN(
        n22224) );
  MUX2_X1 U23009 ( .A(n23740), .B(n23743), .S(n24064), .Z(n22259) );
  NOR2_X1 U23010 ( .A1(n22226), .A2(n22225), .ZN(n22230) );
  NOR2_X1 U23011 ( .A1(n22228), .A2(n24905), .ZN(n22229) );
  MUX2_X1 U23012 ( .A(n22230), .B(n22229), .S(n22231), .Z(n22238) );
  INV_X1 U23013 ( .A(n22231), .ZN(n22234) );
  AOI21_X1 U23014 ( .B1(n22234), .B2(n22233), .A(n22232), .ZN(n22236) );
  NOR2_X1 U23015 ( .A1(n22236), .A2(n22235), .ZN(n22237) );
  NAND2_X1 U23019 ( .A1(n22240), .A2(n22243), .ZN(n22248) );
  OAI21_X1 U23020 ( .B1(n22243), .B2(n22242), .A(n22241), .ZN(n22247) );
  MUX2_X1 U23021 ( .A(n24063), .B(n23730), .S(n23748), .Z(n22258) );
  NAND2_X1 U23022 ( .A1(n24468), .A2(n22252), .ZN(n22253) );
  XNOR2_X1 U23023 ( .A(n22260), .B(n1864), .ZN(Ciphertext[140]) );
  AOI22_X1 U23024 ( .A1(n22456), .A2(n5224), .B1(n25487), .B2(n22324), .ZN(
        n22272) );
  OAI21_X1 U23025 ( .B1(n22452), .B2(n24496), .A(n1352), .ZN(n22271) );
  OAI21_X1 U23026 ( .B1(n22272), .B2(n24311), .A(n22271), .ZN(n23242) );
  OAI21_X1 U23027 ( .B1(n22338), .B2(n22274), .A(n22273), .ZN(n22277) );
  NAND2_X1 U23028 ( .A1(n21368), .A2(n22275), .ZN(n22276) );
  OAI21_X1 U23030 ( .B1(n24377), .B2(n23242), .A(n22298), .ZN(n22278) );
  XNOR2_X1 U23031 ( .A(n22278), .B(n4668), .ZN(n22297) );
  AND2_X1 U23032 ( .A1(n22946), .A2(n22421), .ZN(n22280) );
  NOR2_X1 U23033 ( .A1(n22426), .A2(n22947), .ZN(n22279) );
  INV_X1 U23034 ( .A(n22421), .ZN(n22281) );
  NAND2_X1 U23035 ( .A1(n22341), .A2(n22409), .ZN(n22285) );
  MUX2_X1 U23036 ( .A(n22566), .B(n22409), .S(n24971), .Z(n22284) );
  AND2_X1 U23037 ( .A1(n22411), .A2(n22567), .ZN(n22286) );
  INV_X1 U23038 ( .A(n22977), .ZN(n22288) );
  NAND2_X1 U23039 ( .A1(n22387), .A2(n22288), .ZN(n22291) );
  INV_X1 U23040 ( .A(n22972), .ZN(n22388) );
  AOI21_X1 U23041 ( .B1(n22977), .B2(n22974), .A(n22388), .ZN(n22290) );
  NOR2_X1 U23042 ( .A1(n24881), .A2(n22975), .ZN(n22289) );
  XNOR2_X1 U23044 ( .A(n23252), .B(n4668), .ZN(n22294) );
  XNOR2_X1 U23045 ( .A(n23251), .B(n4668), .ZN(n22295) );
  NAND2_X1 U23046 ( .A1(n23256), .A2(n22295), .ZN(n22296) );
  INV_X1 U23047 ( .A(n23251), .ZN(n23241) );
  INV_X1 U23048 ( .A(n23242), .ZN(n23249) );
  NAND3_X1 U23049 ( .A1(n23245), .A2(n23241), .A3(n23249), .ZN(n22299) );
  INV_X1 U23050 ( .A(n1870), .ZN(n22301) );
  OR2_X1 U23052 ( .A1(n24933), .A2(n23394), .ZN(n23385) );
  AOI21_X1 U23053 ( .B1(n24880), .B2(n23385), .A(n23392), .ZN(n22306) );
  INV_X1 U23054 ( .A(n24465), .ZN(n22304) );
  NAND3_X1 U23055 ( .A1(n23396), .A2(n23394), .A3(n23392), .ZN(n22303) );
  NOR2_X1 U23056 ( .A1(n22306), .A2(n22305), .ZN(n22307) );
  XNOR2_X1 U23057 ( .A(n22307), .B(n1739), .ZN(Ciphertext[79]) );
  NOR2_X1 U23059 ( .A1(n22309), .A2(n23743), .ZN(n22311) );
  XNOR2_X1 U23061 ( .A(n22312), .B(n62), .ZN(Ciphertext[142]) );
  AND2_X1 U23062 ( .A1(n22615), .A2(n22619), .ZN(n22472) );
  INV_X1 U23063 ( .A(n22472), .ZN(n22316) );
  NOR2_X1 U23064 ( .A1(n22615), .A2(n22612), .ZN(n22788) );
  OAI21_X1 U23065 ( .B1(n22788), .B2(n22617), .A(n22792), .ZN(n22315) );
  NOR2_X1 U23066 ( .A1(n22448), .A2(n274), .ZN(n22321) );
  NAND2_X1 U23067 ( .A1(n25066), .A2(n22592), .ZN(n22320) );
  NOR2_X1 U23068 ( .A1(n22591), .A2(n22318), .ZN(n22319) );
  OAI21_X1 U23069 ( .B1(n22321), .B2(n22320), .A(n22319), .ZN(n23178) );
  NOR2_X1 U23070 ( .A1(n24496), .A2(n22323), .ZN(n22325) );
  MUX2_X1 U23071 ( .A(n23164), .B(n23178), .S(n23177), .Z(n22345) );
  INV_X1 U23072 ( .A(n23177), .ZN(n23168) );
  OR3_X1 U23073 ( .A1(n22462), .A2(n22465), .A3(n22464), .ZN(n22332) );
  INV_X1 U23074 ( .A(n22328), .ZN(n22330) );
  OAI21_X1 U23075 ( .B1(n22511), .B2(n25496), .A(n23165), .ZN(n22340) );
  MUX2_X1 U23076 ( .A(n22338), .B(n4350), .S(n22337), .Z(n22512) );
  NOR2_X1 U23077 ( .A1(n22512), .A2(n22511), .ZN(n22339) );
  OAI22_X1 U23078 ( .A1(n23168), .A2(n23165), .B1(n22340), .B2(n22339), .ZN(
        n22344) );
  INV_X1 U23079 ( .A(n22566), .ZN(n22412) );
  OAI21_X1 U23080 ( .B1(n22409), .B2(n22407), .A(n22341), .ZN(n22342) );
  INV_X1 U23082 ( .A(n2005), .ZN(n22346) );
  XNOR2_X1 U23083 ( .A(n22347), .B(n22346), .ZN(Ciphertext[26]) );
  INV_X1 U23085 ( .A(n22348), .ZN(n22351) );
  NAND2_X1 U23086 ( .A1(n22349), .A2(n22689), .ZN(n22350) );
  INV_X1 U23088 ( .A(n23933), .ZN(n23918) );
  AOI21_X1 U23089 ( .B1(n22356), .B2(n22355), .A(n245), .ZN(n22357) );
  INV_X1 U23090 ( .A(n22357), .ZN(n22362) );
  INV_X1 U23091 ( .A(n23940), .ZN(n23934) );
  INV_X1 U23092 ( .A(n22656), .ZN(n22810) );
  MUX2_X1 U23093 ( .A(n23918), .B(n23934), .S(n23926), .Z(n22381) );
  NAND2_X1 U23094 ( .A1(n22670), .A2(n25023), .ZN(n22364) );
  NAND2_X1 U23095 ( .A1(n24963), .A2(n25023), .ZN(n22366) );
  AOI21_X1 U23096 ( .B1(n22366), .B2(n22670), .A(n22779), .ZN(n22367) );
  OR2_X2 U23097 ( .A1(n22368), .A2(n22367), .ZN(n23924) );
  INV_X1 U23098 ( .A(n23924), .ZN(n23938) );
  MUX2_X1 U23099 ( .A(n22679), .B(n22369), .S(n22774), .Z(n22372) );
  NAND2_X1 U23101 ( .A1(n22376), .A2(n25439), .ZN(n22375) );
  NAND2_X1 U23102 ( .A1(n22373), .A2(n25414), .ZN(n22374) );
  OAI211_X1 U23103 ( .C1(n22376), .C2(n22677), .A(n22375), .B(n22374), .ZN(
        n22378) );
  NAND3_X1 U23104 ( .A1(n23997), .A2(n25439), .A3(n25079), .ZN(n22377) );
  AOI21_X1 U23105 ( .B1(n23939), .B2(n23926), .A(n23924), .ZN(n22379) );
  OAI21_X1 U23106 ( .B1(n24948), .B2(n23937), .A(n22379), .ZN(n22380) );
  OAI21_X1 U23107 ( .B1(n22381), .B2(n23938), .A(n22380), .ZN(n22383) );
  XNOR2_X1 U23108 ( .A(n22383), .B(n22382), .ZN(Ciphertext[176]) );
  XNOR2_X1 U23109 ( .A(n22386), .B(n22385), .ZN(Ciphertext[62]) );
  NOR2_X1 U23111 ( .A1(n22387), .A2(n22975), .ZN(n22391) );
  NOR2_X1 U23112 ( .A1(n22388), .A2(n22977), .ZN(n22390) );
  NOR2_X1 U23113 ( .A1(n22397), .A2(n22396), .ZN(n22399) );
  NOR2_X1 U23114 ( .A1(n22399), .A2(n25381), .ZN(n22403) );
  NOR2_X1 U23117 ( .A1(n1593), .A2(n22407), .ZN(n22408) );
  NOR2_X1 U23118 ( .A1(n22562), .A2(n22409), .ZN(n22410) );
  AOI21_X1 U23119 ( .B1(n22412), .B2(n22411), .A(n22410), .ZN(n22413) );
  NOR2_X1 U23120 ( .A1(n23293), .A2(n23305), .ZN(n22415) );
  MUX2_X1 U23121 ( .A(n22969), .B(n22966), .S(n21476), .Z(n22419) );
  NAND2_X1 U23122 ( .A1(n22962), .A2(n22965), .ZN(n22417) );
  MUX2_X1 U23124 ( .A(n22417), .B(n22416), .S(n22966), .Z(n22418) );
  OAI21_X1 U23125 ( .B1(n22419), .B2(n22962), .A(n22418), .ZN(n23297) );
  INV_X1 U23126 ( .A(n23297), .ZN(n23308) );
  INV_X1 U23129 ( .A(n23285), .ZN(n22509) );
  NAND3_X1 U23130 ( .A1(n22510), .A2(n22509), .A3(n23293), .ZN(n22427) );
  OAI21_X1 U23131 ( .B1(n23309), .B2(n23298), .A(n22427), .ZN(n22429) );
  INV_X1 U23132 ( .A(n2726), .ZN(n22428) );
  XNOR2_X1 U23133 ( .A(n22429), .B(n22428), .ZN(Ciphertext[55]) );
  NOR2_X1 U23134 ( .A1(n23371), .A2(n22987), .ZN(n23375) );
  INV_X1 U23135 ( .A(n22987), .ZN(n23368) );
  INV_X1 U23136 ( .A(n22431), .ZN(n22434) );
  INV_X1 U23137 ( .A(n22432), .ZN(n22433) );
  OAI211_X1 U23138 ( .C1(n22436), .C2(n22435), .A(n22434), .B(n22433), .ZN(
        n22437) );
  OAI21_X1 U23139 ( .B1(n24911), .B2(n24412), .A(n22437), .ZN(n22438) );
  NAND2_X1 U23140 ( .A1(n22438), .A2(n4606), .ZN(n22439) );
  NAND2_X1 U23141 ( .A1(n24906), .A2(n23146), .ZN(n22441) );
  OAI21_X1 U23142 ( .B1(n24906), .B2(n22442), .A(n22441), .ZN(n22446) );
  NOR2_X1 U23143 ( .A1(n23155), .A2(n24473), .ZN(n22443) );
  NAND2_X1 U23144 ( .A1(n22443), .A2(n24325), .ZN(n22444) );
  XNOR2_X1 U23146 ( .A(n22447), .B(n886), .ZN(Ciphertext[22]) );
  MUX2_X1 U23148 ( .A(n25450), .B(n24367), .S(n22459), .Z(n22466) );
  INV_X1 U23149 ( .A(n23125), .ZN(n23094) );
  INV_X1 U23151 ( .A(n25462), .ZN(n22603) );
  NAND3_X1 U23152 ( .A1(n25068), .A2(n22603), .A3(n24963), .ZN(n22471) );
  NOR2_X1 U23154 ( .A1(n24963), .A2(n24607), .ZN(n22468) );
  NAND2_X1 U23155 ( .A1(n22675), .A2(n22780), .ZN(n22469) );
  AOI21_X1 U23156 ( .B1(n24941), .B2(n23094), .A(n5036), .ZN(n22480) );
  NOR2_X1 U23157 ( .A1(n22792), .A2(n22619), .ZN(n22623) );
  NOR2_X1 U23158 ( .A1(n22623), .A2(n22472), .ZN(n22473) );
  INV_X1 U23159 ( .A(n23104), .ZN(n23110) );
  INV_X1 U23161 ( .A(n23112), .ZN(n23122) );
  MUX2_X1 U23162 ( .A(n22475), .B(n22804), .S(n25115), .Z(n22477) );
  NOR2_X1 U23164 ( .A1(n23122), .A2(n24059), .ZN(n22478) );
  OAI21_X1 U23165 ( .B1(n23093), .B2(n22478), .A(n23125), .ZN(n22479) );
  NAND2_X1 U23166 ( .A1(n22482), .A2(n22842), .ZN(n22486) );
  INV_X1 U23167 ( .A(n22900), .ZN(n22847) );
  NOR2_X1 U23168 ( .A1(n22905), .A2(n22904), .ZN(n22721) );
  NAND2_X1 U23169 ( .A1(n22906), .A2(n22721), .ZN(n22485) );
  NAND3_X1 U23170 ( .A1(n22837), .A2(n25041), .A3(n22893), .ZN(n22487) );
  INV_X1 U23171 ( .A(n22835), .ZN(n22894) );
  NOR2_X1 U23172 ( .A1(n22897), .A2(n22894), .ZN(n22488) );
  NOR2_X1 U23173 ( .A1(n3176), .A2(n23458), .ZN(n22490) );
  NAND2_X1 U23174 ( .A1(n23464), .A2(n23016), .ZN(n22492) );
  INV_X1 U23175 ( .A(n23015), .ZN(n22864) );
  AOI21_X1 U23176 ( .B1(n22492), .B2(n22914), .A(n22864), .ZN(n22493) );
  AOI21_X1 U23177 ( .B1(n327), .B2(n22889), .A(n22728), .ZN(n22495) );
  AOI21_X1 U23178 ( .B1(n22496), .B2(n22887), .A(n3837), .ZN(n22497) );
  NAND2_X1 U23179 ( .A1(n23332), .A2(n22932), .ZN(n22856) );
  NAND2_X1 U23180 ( .A1(n22856), .A2(n22498), .ZN(n22504) );
  AND2_X1 U23181 ( .A1(n24342), .A2(n22499), .ZN(n22500) );
  NOR2_X1 U23182 ( .A1(n22855), .A2(n22500), .ZN(n22503) );
  NAND2_X1 U23183 ( .A1(n22501), .A2(n24356), .ZN(n22502) );
  NOR2_X1 U23184 ( .A1(n22938), .A2(n22832), .ZN(n22505) );
  XNOR2_X1 U23185 ( .A(n22507), .B(n16574), .ZN(Ciphertext[92]) );
  NOR2_X1 U23186 ( .A1(n23292), .A2(n23305), .ZN(n22763) );
  NOR2_X1 U23187 ( .A1(n24904), .A2(n22509), .ZN(n23306) );
  INV_X1 U23188 ( .A(n23181), .ZN(n22513) );
  INV_X1 U23189 ( .A(n23165), .ZN(n23179) );
  NAND3_X1 U23190 ( .A1(n22513), .A2(n23166), .A3(n23179), .ZN(n22517) );
  INV_X1 U23191 ( .A(n23166), .ZN(n22551) );
  NAND3_X1 U23192 ( .A1(n25488), .A2(n23164), .A3(n22551), .ZN(n22516) );
  INV_X1 U23193 ( .A(n23178), .ZN(n23167) );
  INV_X1 U23194 ( .A(n23164), .ZN(n23176) );
  NAND3_X1 U23195 ( .A1(n23165), .A2(n23167), .A3(n23176), .ZN(n22515) );
  NAND3_X1 U23196 ( .A1(n23168), .A2(n23164), .A3(n23165), .ZN(n22514) );
  NAND4_X1 U23197 ( .A1(n22517), .A2(n22516), .A3(n22515), .A4(n22514), .ZN(
        n22519) );
  INV_X1 U23198 ( .A(n812), .ZN(n22518) );
  XNOR2_X1 U23199 ( .A(n22519), .B(n22518), .ZN(Ciphertext[28]) );
  INV_X1 U23200 ( .A(n23770), .ZN(n23781) );
  AOI22_X1 U23201 ( .A1(n23778), .A2(n23768), .B1(n23781), .B2(n24921), .ZN(
        n23783) );
  NAND2_X1 U23202 ( .A1(n25051), .A2(n23757), .ZN(n23758) );
  INV_X1 U23203 ( .A(n23758), .ZN(n22523) );
  XNOR2_X1 U23204 ( .A(n22526), .B(n22525), .ZN(Ciphertext[145]) );
  NAND2_X1 U23205 ( .A1(n25042), .A2(n1370), .ZN(n23437) );
  INV_X1 U23206 ( .A(n23865), .ZN(n23853) );
  AOI21_X1 U23207 ( .B1(n22982), .B2(n23857), .A(n23853), .ZN(n22533) );
  NOR3_X1 U23208 ( .A1(n23860), .A2(n23862), .A3(n25399), .ZN(n22532) );
  NOR3_X1 U23209 ( .A1(n23858), .A2(n25399), .A3(n23865), .ZN(n22531) );
  XNOR2_X1 U23210 ( .A(n22534), .B(n1726), .ZN(Ciphertext[162]) );
  INV_X1 U23211 ( .A(n23275), .ZN(n23278) );
  XNOR2_X1 U23212 ( .A(n22538), .B(n2757), .ZN(Ciphertext[50]) );
  INV_X1 U23213 ( .A(n22539), .ZN(n23813) );
  NOR2_X1 U23214 ( .A1(n23813), .A2(n23030), .ZN(n23833) );
  AND2_X1 U23215 ( .A1(n22539), .A2(n23828), .ZN(n23818) );
  NAND2_X1 U23216 ( .A1(n23818), .A2(n25391), .ZN(n22541) );
  INV_X1 U23217 ( .A(n2193), .ZN(n22542) );
  XNOR2_X1 U23218 ( .A(n22543), .B(n22542), .ZN(Ciphertext[156]) );
  NOR2_X1 U23219 ( .A1(n23904), .A2(n21863), .ZN(n22545) );
  INV_X1 U23220 ( .A(n23906), .ZN(n22544) );
  OAI21_X1 U23221 ( .B1(n23888), .B2(n22545), .A(n22544), .ZN(n22548) );
  INV_X1 U23222 ( .A(n23890), .ZN(n22546) );
  XNOR2_X1 U23223 ( .A(n22550), .B(n22549), .ZN(Ciphertext[168]) );
  NAND3_X1 U23224 ( .A1(n23168), .A2(n23176), .A3(n23166), .ZN(n22554) );
  XNOR2_X1 U23225 ( .A(n22557), .B(n22556), .ZN(Ciphertext[27]) );
  INV_X1 U23226 ( .A(n23743), .ZN(n22558) );
  OAI21_X1 U23227 ( .B1(n23740), .B2(n24065), .A(n22558), .ZN(n22559) );
  OAI22_X1 U23228 ( .A1(n23743), .A2(n23740), .B1(n24991), .B2(n23748), .ZN(
        n23735) );
  INV_X1 U23229 ( .A(n23730), .ZN(n23745) );
  AOI22_X1 U23230 ( .A1(n23748), .A2(n22559), .B1(n23735), .B2(n23745), .ZN(
        n22560) );
  XNOR2_X1 U23231 ( .A(n22560), .B(n4164), .ZN(Ciphertext[143]) );
  NAND2_X1 U23232 ( .A1(n24971), .A2(n22563), .ZN(n22565) );
  OAI22_X1 U23233 ( .A1(n22568), .A2(n22567), .B1(n24951), .B2(n22565), .ZN(
        n22570) );
  OAI21_X1 U23234 ( .B1(n22571), .B2(n22570), .A(n22569), .ZN(n22572) );
  NOR2_X1 U23235 ( .A1(n22573), .A2(n22572), .ZN(n22574) );
  NOR2_X1 U23236 ( .A1(n23184), .A2(n22575), .ZN(n23203) );
  MUX2_X1 U23237 ( .A(n22574), .B(n23203), .S(n24334), .Z(n22576) );
  INV_X1 U23238 ( .A(n23200), .ZN(n22824) );
  INV_X1 U23239 ( .A(n23201), .ZN(n22820) );
  INV_X1 U23240 ( .A(n22578), .ZN(n23069) );
  INV_X1 U23242 ( .A(n23064), .ZN(n22580) );
  INV_X1 U23244 ( .A(n22872), .ZN(n22579) );
  OAI21_X1 U23245 ( .B1(n22580), .B2(n23077), .A(n22579), .ZN(n22581) );
  NOR2_X1 U23246 ( .A1(n22803), .A2(n22805), .ZN(n22582) );
  NAND2_X1 U23248 ( .A1(n22585), .A2(n22584), .ZN(n22587) );
  NAND2_X1 U23249 ( .A1(n22798), .A2(n24561), .ZN(n22586) );
  NOR2_X2 U23250 ( .A1(n22589), .A2(n22588), .ZN(n23052) );
  OAI21_X1 U23251 ( .B1(n22591), .B2(n22590), .A(n22448), .ZN(n22595) );
  OAI211_X1 U23252 ( .C1(n23997), .C2(n22677), .A(n24439), .B(n22596), .ZN(
        n22597) );
  OAI21_X1 U23253 ( .B1(n22598), .B2(n22676), .A(n22597), .ZN(n23047) );
  MUX2_X1 U23254 ( .A(n23052), .B(n23040), .S(n23047), .Z(n22624) );
  NAND2_X1 U23255 ( .A1(n24963), .A2(n22779), .ZN(n22600) );
  OAI21_X1 U23256 ( .B1(n22675), .B2(n22779), .A(n22600), .ZN(n22601) );
  INV_X1 U23257 ( .A(n22601), .ZN(n22605) );
  MUX2_X1 U23258 ( .A(n22670), .B(n25022), .S(n24963), .Z(n22602) );
  INV_X1 U23259 ( .A(n22602), .ZN(n22604) );
  INV_X1 U23260 ( .A(n23050), .ZN(n23058) );
  NOR2_X1 U23261 ( .A1(n22813), .A2(n25241), .ZN(n22608) );
  NOR3_X1 U23262 ( .A1(n22813), .A2(n22606), .A3(n25075), .ZN(n22607) );
  AOI21_X1 U23263 ( .B1(n22656), .B2(n22608), .A(n22607), .ZN(n22611) );
  NAND2_X1 U23265 ( .A1(n22792), .A2(n22612), .ZN(n22613) );
  NAND2_X1 U23266 ( .A1(n22613), .A2(n22617), .ZN(n22622) );
  NOR2_X1 U23267 ( .A1(n22615), .A2(n22614), .ZN(n22616) );
  NAND2_X1 U23268 ( .A1(n24953), .A2(n22616), .ZN(n22621) );
  NAND2_X1 U23269 ( .A1(n22619), .A2(n22618), .ZN(n22620) );
  OAI211_X1 U23270 ( .C1(n22623), .C2(n22622), .A(n22620), .B(n22621), .ZN(
        n22698) );
  XNOR2_X1 U23271 ( .A(n22626), .B(n22625), .ZN(Ciphertext[3]) );
  OAI22_X1 U23272 ( .A1(n23318), .A2(n23326), .B1(n23327), .B2(n23320), .ZN(
        n23325) );
  NAND2_X1 U23273 ( .A1(n23318), .A2(n23313), .ZN(n22627) );
  AOI22_X1 U23274 ( .A1(n22629), .A2(n23325), .B1(n22628), .B2(n22627), .ZN(
        n22630) );
  XNOR2_X1 U23275 ( .A(n22630), .B(n2826), .ZN(Ciphertext[61]) );
  NAND2_X1 U23276 ( .A1(n24390), .A2(n23592), .ZN(n22631) );
  AOI21_X1 U23277 ( .B1(n22632), .B2(n22631), .A(n23591), .ZN(n22642) );
  INV_X1 U23278 ( .A(n23594), .ZN(n23565) );
  AND2_X1 U23279 ( .A1(n23592), .A2(n23565), .ZN(n22637) );
  AOI21_X1 U23280 ( .B1(n22637), .B2(n23591), .A(n22635), .ZN(n22636) );
  AOI21_X1 U23281 ( .B1(n21941), .B2(n24389), .A(n2040), .ZN(n22638) );
  INV_X1 U23282 ( .A(n23047), .ZN(n23053) );
  NOR2_X1 U23283 ( .A1(n23052), .A2(n23053), .ZN(n23060) );
  INV_X1 U23284 ( .A(n23052), .ZN(n23042) );
  INV_X1 U23285 ( .A(n23040), .ZN(n23049) );
  OAI21_X1 U23286 ( .B1(n23042), .B2(n23059), .A(n23049), .ZN(n22646) );
  NAND2_X1 U23287 ( .A1(n22643), .A2(n23050), .ZN(n22645) );
  OAI211_X1 U23288 ( .C1(n23060), .C2(n22646), .A(n22645), .B(n22644), .ZN(
        n22647) );
  XNOR2_X1 U23289 ( .A(n22647), .B(n3073), .ZN(Ciphertext[2]) );
  INV_X1 U23291 ( .A(n23252), .ZN(n23236) );
  AOI22_X1 U23292 ( .A1(n22650), .A2(n22649), .B1(n22648), .B2(n23256), .ZN(
        n22651) );
  XNOR2_X1 U23293 ( .A(n22651), .B(n663), .ZN(Ciphertext[46]) );
  MUX2_X1 U23294 ( .A(n23227), .B(n23228), .S(n24955), .Z(n22653) );
  XNOR2_X1 U23296 ( .A(n22654), .B(n1863), .ZN(Ciphertext[38]) );
  NOR2_X1 U23297 ( .A1(n22804), .A2(n22805), .ZN(n22802) );
  AND2_X1 U23298 ( .A1(n22798), .A2(n22803), .ZN(n22661) );
  NOR2_X1 U23300 ( .A1(n22800), .A2(n24559), .ZN(n22663) );
  NAND2_X1 U23301 ( .A1(n22663), .A2(n22804), .ZN(n22664) );
  NAND2_X1 U23302 ( .A1(n22779), .A2(n25462), .ZN(n22674) );
  NAND2_X1 U23303 ( .A1(n24963), .A2(n22782), .ZN(n22669) );
  INV_X1 U23304 ( .A(n22667), .ZN(n22783) );
  NOR2_X1 U23305 ( .A1(n22779), .A2(n25023), .ZN(n22671) );
  INV_X1 U23306 ( .A(n23958), .ZN(n23952) );
  NOR2_X1 U23307 ( .A1(n23969), .A2(n23952), .ZN(n23970) );
  INV_X1 U23308 ( .A(n23970), .ZN(n22696) );
  NAND3_X1 U23309 ( .A1(n22771), .A2(n22680), .A3(n22769), .ZN(n22681) );
  AOI22_X1 U23313 ( .A1(n21848), .A2(n22687), .B1(n22686), .B2(n22685), .ZN(
        n22692) );
  OAI21_X1 U23314 ( .B1(n22690), .B2(n22689), .A(n22688), .ZN(n22691) );
  OAI21_X1 U23315 ( .B1(n22692), .B2(n25395), .A(n22691), .ZN(n23966) );
  NAND2_X1 U23316 ( .A1(n22693), .A2(n23966), .ZN(n22694) );
  AND2_X1 U23317 ( .A1(n23966), .A2(n24910), .ZN(n23953) );
  AOI22_X1 U23318 ( .A1(n25076), .A2(n22694), .B1(n23953), .B2(n25017), .ZN(
        n22695) );
  NAND2_X1 U23319 ( .A1(n23040), .A2(n22698), .ZN(n22699) );
  INV_X1 U23320 ( .A(n23537), .ZN(n23557) );
  OAI21_X1 U23321 ( .B1(n25071), .B2(n23555), .A(n24893), .ZN(n22700) );
  AOI22_X1 U23322 ( .A1(n22701), .A2(n23557), .B1(n23554), .B2(n22700), .ZN(
        n22703) );
  XNOR2_X1 U23323 ( .A(n22703), .B(n22702), .ZN(Ciphertext[113]) );
  INV_X1 U23326 ( .A(n23259), .ZN(n23282) );
  INV_X1 U23327 ( .A(n23281), .ZN(n23267) );
  OR2_X1 U23328 ( .A1(n23277), .A2(n24349), .ZN(n22705) );
  OAI22_X1 U23329 ( .A1(n23282), .A2(n24360), .B1(n23267), .B2(n22705), .ZN(
        n22708) );
  NOR2_X1 U23330 ( .A1(n23277), .A2(n23273), .ZN(n22706) );
  NOR2_X1 U23331 ( .A1(n22708), .A2(n22707), .ZN(n22709) );
  XNOR2_X1 U23332 ( .A(n22709), .B(n673), .ZN(Ciphertext[48]) );
  MUX2_X1 U23333 ( .A(n23546), .B(n23537), .S(n23554), .Z(n22710) );
  INV_X1 U23334 ( .A(n22711), .ZN(n22716) );
  NOR2_X1 U23335 ( .A1(n22712), .A2(n22928), .ZN(n22713) );
  OAI21_X1 U23336 ( .B1(n22713), .B2(n22107), .A(n22926), .ZN(n22714) );
  INV_X1 U23337 ( .A(n23479), .ZN(n23483) );
  MUX2_X1 U23338 ( .A(n22717), .B(n22841), .S(n25041), .Z(n22720) );
  INV_X1 U23339 ( .A(n25041), .ZN(n22718) );
  MUX2_X1 U23340 ( .A(n22718), .B(n22835), .S(n25438), .Z(n22719) );
  NAND2_X1 U23341 ( .A1(n24932), .A2(n22832), .ZN(n22724) );
  INV_X1 U23342 ( .A(n22939), .ZN(n22723) );
  NAND2_X1 U23343 ( .A1(n22938), .A2(n22832), .ZN(n22935) );
  AOI21_X1 U23344 ( .B1(n22935), .B2(n22829), .A(n22723), .ZN(n22725) );
  NOR2_X1 U23346 ( .A1(n23491), .A2(n23481), .ZN(n23495) );
  MUX2_X1 U23348 ( .A(n22889), .B(n22727), .S(n22890), .Z(n22732) );
  NOR2_X1 U23349 ( .A1(n22729), .A2(n22890), .ZN(n22731) );
  NOR2_X1 U23350 ( .A1(n23464), .A2(n23458), .ZN(n22734) );
  INV_X1 U23351 ( .A(n23464), .ZN(n22733) );
  INV_X1 U23352 ( .A(n22911), .ZN(n23462) );
  AND3_X1 U23353 ( .A1(n22864), .A2(n23016), .A3(n23014), .ZN(n23467) );
  AOI21_X1 U23354 ( .B1(n22734), .B2(n23460), .A(n23467), .ZN(n22735) );
  NAND3_X1 U23355 ( .A1(n22736), .A2(n23492), .A3(n24442), .ZN(n22737) );
  XNOR2_X1 U23357 ( .A(n22740), .B(n22739), .ZN(Ciphertext[97]) );
  NAND2_X1 U23358 ( .A1(n22988), .A2(n23374), .ZN(n22743) );
  NAND2_X1 U23359 ( .A1(n22741), .A2(n24515), .ZN(n22989) );
  OAI211_X1 U23360 ( .C1(n22741), .C2(n23368), .A(n23379), .B(n22989), .ZN(
        n22742) );
  XNOR2_X1 U23361 ( .A(n22746), .B(n22745), .ZN(Ciphertext[75]) );
  INV_X1 U23362 ( .A(n23670), .ZN(n22749) );
  INV_X1 U23363 ( .A(n23689), .ZN(n22747) );
  NAND2_X1 U23364 ( .A1(n22747), .A2(n23690), .ZN(n23659) );
  OAI21_X1 U23365 ( .B1(n22749), .B2(n23692), .A(n23659), .ZN(n22750) );
  NAND2_X1 U23366 ( .A1(n23676), .A2(n23690), .ZN(n22748) );
  INV_X1 U23369 ( .A(n22752), .ZN(n23193) );
  NAND2_X1 U23370 ( .A1(n23193), .A2(n23206), .ZN(n22754) );
  NAND2_X1 U23371 ( .A1(n23201), .A2(n23184), .ZN(n22753) );
  OAI21_X1 U23372 ( .B1(n22754), .B2(n23196), .A(n22753), .ZN(n22821) );
  AOI21_X1 U23373 ( .B1(n24334), .B2(n25059), .A(n5769), .ZN(n22756) );
  NAND2_X1 U23374 ( .A1(n5769), .A2(n23206), .ZN(n22755) );
  OAI22_X1 U23375 ( .A1(n22821), .A2(n22756), .B1(n22755), .B2(n23200), .ZN(
        n22757) );
  XNOR2_X1 U23376 ( .A(n22757), .B(n2222), .ZN(Ciphertext[31]) );
  MUX2_X1 U23377 ( .A(n23178), .B(n23164), .S(n25488), .Z(n22759) );
  AOI21_X1 U23378 ( .B1(n23181), .B2(n23179), .A(n23166), .ZN(n22758) );
  OAI22_X1 U23379 ( .A1(n22759), .A2(n22758), .B1(n23181), .B2(n24394), .ZN(
        n22760) );
  XNOR2_X1 U23380 ( .A(n22760), .B(n1952), .ZN(Ciphertext[24]) );
  INV_X1 U23381 ( .A(n24904), .ZN(n23299) );
  BUF_X1 U23382 ( .A(n23285), .Z(n23294) );
  OAI21_X1 U23383 ( .B1(n23293), .B2(n22762), .A(n22761), .ZN(n22766) );
  AND2_X1 U23384 ( .A1(n23297), .A2(n23292), .ZN(n22764) );
  AOI22_X1 U23385 ( .A1(n22763), .A2(n23294), .B1(n22764), .B2(n23303), .ZN(
        n22765) );
  OAI21_X1 U23386 ( .B1(n22766), .B2(n23303), .A(n22765), .ZN(n22768) );
  XNOR2_X1 U23387 ( .A(n22768), .B(n22767), .ZN(Ciphertext[58]) );
  MUX2_X1 U23388 ( .A(n25414), .B(n23998), .S(n24439), .Z(n22776) );
  NAND2_X1 U23391 ( .A1(n25068), .A2(n22780), .ZN(n22786) );
  NAND3_X1 U23392 ( .A1(n22784), .A2(n22783), .A3(n25462), .ZN(n22785) );
  NAND2_X1 U23394 ( .A1(n22788), .A2(n24953), .ZN(n22797) );
  NAND2_X1 U23395 ( .A1(n22790), .A2(n22789), .ZN(n22796) );
  NAND2_X1 U23397 ( .A1(n24006), .A2(n24010), .ZN(n23984) );
  NOR2_X1 U23399 ( .A1(n22800), .A2(n25115), .ZN(n22801) );
  AOI22_X1 U23400 ( .A1(n22802), .A2(n22584), .B1(n22801), .B2(n22804), .ZN(
        n22808) );
  NOR2_X1 U23401 ( .A1(n22804), .A2(n22803), .ZN(n22807) );
  NOR2_X1 U23402 ( .A1(n22810), .A2(n25241), .ZN(n22816) );
  NOR2_X1 U23403 ( .A1(n22812), .A2(n22811), .ZN(n22815) );
  OAI21_X1 U23404 ( .B1(n22813), .B2(n22812), .A(n1477), .ZN(n22814) );
  OAI21_X1 U23407 ( .B1(n22820), .B2(n23202), .A(n24889), .ZN(n22823) );
  INV_X1 U23408 ( .A(n23186), .ZN(n22822) );
  AOI22_X1 U23409 ( .A1(n22824), .A2(n22823), .B1(n22822), .B2(n22821), .ZN(
        n22825) );
  XNOR2_X1 U23410 ( .A(n22825), .B(n1856), .ZN(Ciphertext[35]) );
  INV_X1 U23411 ( .A(n24910), .ZN(n23964) );
  INV_X1 U23412 ( .A(n23967), .ZN(n23947) );
  MUX2_X1 U23413 ( .A(n23964), .B(n23947), .S(n23966), .Z(n22828) );
  NOR2_X1 U23414 ( .A1(n22939), .A2(n22829), .ZN(n22830) );
  MUX2_X1 U23415 ( .A(n22834), .B(n25438), .S(n25041), .Z(n22840) );
  NOR2_X1 U23419 ( .A1(n142), .A2(n25035), .ZN(n22851) );
  INV_X1 U23421 ( .A(n22033), .ZN(n22859) );
  OAI21_X1 U23422 ( .B1(n22958), .B2(n22959), .A(n22859), .ZN(n22860) );
  AND2_X1 U23423 ( .A1(n22860), .A2(n4128), .ZN(n22861) );
  XNOR2_X1 U23425 ( .A(n22867), .B(n2049), .ZN(Ciphertext[86]) );
  INV_X1 U23426 ( .A(n23403), .ZN(n23418) );
  XNOR2_X1 U23427 ( .A(n22870), .B(n1896), .ZN(Ciphertext[87]) );
  NOR2_X1 U23429 ( .A1(n24075), .A2(n23064), .ZN(n23076) );
  NAND3_X1 U23431 ( .A1(n23064), .A2(n23074), .A3(n23066), .ZN(n22873) );
  AOI21_X1 U23434 ( .B1(n25179), .B2(n25452), .A(n23064), .ZN(n22878) );
  NAND2_X1 U23435 ( .A1(n23074), .A2(n23066), .ZN(n22877) );
  AOI22_X1 U23436 ( .A1(n22879), .A2(n23064), .B1(n22878), .B2(n22877), .ZN(
        n22880) );
  XNOR2_X1 U23437 ( .A(n22880), .B(n2746), .ZN(Ciphertext[8]) );
  NAND2_X1 U23438 ( .A1(n23394), .A2(n24933), .ZN(n22881) );
  NAND2_X1 U23439 ( .A1(n22881), .A2(n23396), .ZN(n22883) );
  AND3_X1 U23440 ( .A1(n23394), .A2(n23396), .A3(n23393), .ZN(n22882) );
  NOR2_X1 U23441 ( .A1(n25375), .A2(n22887), .ZN(n22892) );
  NOR2_X1 U23442 ( .A1(n22729), .A2(n22889), .ZN(n22891) );
  MUX2_X1 U23443 ( .A(n22892), .B(n22891), .S(n22890), .Z(n23514) );
  NAND2_X1 U23444 ( .A1(n22894), .A2(n22893), .ZN(n22899) );
  INV_X1 U23445 ( .A(n22895), .ZN(n22898) );
  AOI22_X1 U23446 ( .A1(n22899), .A2(n22898), .B1(n22897), .B2(n22896), .ZN(
        n22915) );
  OR2_X1 U23447 ( .A1(n24380), .A2(n23510), .ZN(n23013) );
  AND2_X1 U23448 ( .A1(n22900), .A2(n22901), .ZN(n22902) );
  NOR2_X1 U23449 ( .A1(n22903), .A2(n22902), .ZN(n22910) );
  OAI21_X1 U23450 ( .B1(n22906), .B2(n22905), .A(n22904), .ZN(n22909) );
  MUX2_X1 U23452 ( .A(n23016), .B(n22911), .S(n23464), .Z(n22913) );
  NAND2_X1 U23453 ( .A1(n23016), .A2(n3176), .ZN(n22912) );
  OR2_X1 U23454 ( .A1(n22914), .A2(n24364), .ZN(n23018) );
  INV_X1 U23455 ( .A(n22915), .ZN(n23530) );
  NAND2_X1 U23456 ( .A1(n23530), .A2(n23529), .ZN(n22921) );
  XNOR2_X1 U23458 ( .A(n22930), .B(n2120), .ZN(Ciphertext[107]) );
  NOR2_X1 U23459 ( .A1(n24309), .A2(n23334), .ZN(n22931) );
  AOI21_X1 U23460 ( .B1(n22936), .B2(n22935), .A(n22934), .ZN(n22943) );
  NAND2_X1 U23462 ( .A1(n23361), .A2(n24492), .ZN(n22979) );
  INV_X1 U23464 ( .A(n22945), .ZN(n22950) );
  NOR2_X1 U23466 ( .A1(n22033), .A2(n22953), .ZN(n22955) );
  MUX2_X1 U23467 ( .A(n22958), .B(n24922), .S(n24884), .Z(n22960) );
  INV_X1 U23468 ( .A(n22962), .ZN(n22963) );
  OAI21_X1 U23469 ( .B1(n22965), .B2(n21476), .A(n22964), .ZN(n22971) );
  OAI22_X1 U23470 ( .A1(n22387), .A2(n22974), .B1(n22977), .B2(n22973), .ZN(
        n22976) );
  AOI22_X2 U23471 ( .A1(n22978), .A2(n22977), .B1(n22976), .B2(n25365), .ZN(
        n23359) );
  XNOR2_X1 U23472 ( .A(n22980), .B(n1768), .ZN(Ciphertext[67]) );
  INV_X1 U23475 ( .A(n22989), .ZN(n22990) );
  AOI22_X1 U23476 ( .A1(n22993), .A2(n22992), .B1(n22991), .B2(n22990), .ZN(
        n22994) );
  XNOR2_X1 U23477 ( .A(n22994), .B(n1792), .ZN(Ciphertext[73]) );
  INV_X1 U23478 ( .A(n23350), .ZN(n23340) );
  NAND3_X1 U23479 ( .A1(n22961), .A2(n24492), .A3(n23359), .ZN(n22995) );
  NAND2_X1 U23480 ( .A1(n23670), .A2(n23692), .ZN(n22997) );
  NOR2_X1 U23481 ( .A1(n22997), .A2(n23658), .ZN(n23000) );
  NOR2_X1 U23482 ( .A1(n22998), .A2(n23692), .ZN(n22999) );
  NAND2_X1 U23483 ( .A1(n23805), .A2(n23786), .ZN(n23005) );
  INV_X1 U23484 ( .A(n24392), .ZN(n23796) );
  OAI21_X1 U23485 ( .B1(n21837), .B2(n23002), .A(n23796), .ZN(n23003) );
  XNOR2_X1 U23486 ( .A(n23006), .B(n2782), .ZN(Ciphertext[155]) );
  AOI21_X1 U23487 ( .B1(n23525), .B2(n24351), .A(n23530), .ZN(n23007) );
  AOI22_X1 U23488 ( .A1(n23009), .A2(n23008), .B1(n23527), .B2(n23007), .ZN(
        n23010) );
  XNOR2_X1 U23489 ( .A(n23010), .B(n2042), .ZN(Ciphertext[103]) );
  INV_X1 U23490 ( .A(n23470), .ZN(n23011) );
  XNOR2_X1 U23491 ( .A(n23012), .B(n2050), .ZN(Ciphertext[100]) );
  NAND2_X1 U23492 ( .A1(n24380), .A2(n23529), .ZN(n23533) );
  OAI21_X1 U23493 ( .B1(n25055), .B2(n23460), .A(n23014), .ZN(n23019) );
  NAND3_X1 U23494 ( .A1(n23016), .A2(n23461), .A3(n3176), .ZN(n23017) );
  OAI211_X1 U23495 ( .C1(n24435), .C2(n23019), .A(n23018), .B(n23017), .ZN(
        n23022) );
  NAND2_X1 U23496 ( .A1(n23022), .A2(n23505), .ZN(n23021) );
  OAI211_X1 U23497 ( .C1(n23527), .C2(n23022), .A(n24351), .B(n23021), .ZN(
        n23023) );
  NAND2_X1 U23498 ( .A1(n23024), .A2(n23023), .ZN(n23025) );
  XNOR2_X1 U23499 ( .A(n23025), .B(n2100), .ZN(Ciphertext[104]) );
  NAND2_X1 U23500 ( .A1(n23939), .A2(n23924), .ZN(n23920) );
  NAND2_X1 U23501 ( .A1(n25084), .A2(n23933), .ZN(n23921) );
  NAND2_X1 U23502 ( .A1(n23920), .A2(n23921), .ZN(n23028) );
  INV_X1 U23503 ( .A(n24948), .ZN(n23027) );
  OAI21_X1 U23504 ( .B1(n23926), .B2(n23918), .A(n25084), .ZN(n23026) );
  AOI22_X1 U23505 ( .A1(n23028), .A2(n23937), .B1(n23027), .B2(n23026), .ZN(
        n23029) );
  XNOR2_X1 U23506 ( .A(n23029), .B(n2989), .ZN(Ciphertext[179]) );
  NOR2_X1 U23507 ( .A1(n23810), .A2(n23817), .ZN(n23830) );
  INV_X1 U23508 ( .A(n23828), .ZN(n23032) );
  AND2_X1 U23509 ( .A1(n23828), .A2(n23030), .ZN(n23031) );
  AOI21_X1 U23510 ( .B1(n23810), .B2(n23032), .A(n23031), .ZN(n23033) );
  XNOR2_X1 U23511 ( .A(n23035), .B(n2058), .ZN(Ciphertext[158]) );
  NOR3_X1 U23512 ( .A1(n23361), .A2(n24492), .A3(n22961), .ZN(n23036) );
  AOI211_X1 U23513 ( .C1(n23361), .C2(n23037), .A(n23355), .B(n23036), .ZN(
        n23038) );
  XNOR2_X1 U23514 ( .A(n23038), .B(n2034), .ZN(Ciphertext[66]) );
  OAI21_X1 U23516 ( .B1(n23039), .B2(n23055), .A(n322), .ZN(n23044) );
  OAI21_X1 U23517 ( .B1(n322), .B2(n23040), .A(n23059), .ZN(n23041) );
  NAND2_X1 U23518 ( .A1(n23042), .A2(n23041), .ZN(n23043) );
  NAND2_X1 U23519 ( .A1(n23044), .A2(n23043), .ZN(n23046) );
  XNOR2_X1 U23520 ( .A(n23046), .B(n23045), .ZN(Ciphertext[0]) );
  AOI22_X1 U23521 ( .A1(n23050), .A2(n23049), .B1(n23048), .B2(n23047), .ZN(
        n23062) );
  OAI21_X1 U23522 ( .B1(n23062), .B2(n23055), .A(n23054), .ZN(n23057) );
  INV_X1 U23523 ( .A(n881), .ZN(n23056) );
  XNOR2_X1 U23524 ( .A(n23057), .B(n23056), .ZN(Ciphertext[1]) );
  OAI21_X1 U23525 ( .B1(n23060), .B2(n23059), .A(n23058), .ZN(n23061) );
  INV_X1 U23526 ( .A(n681), .ZN(n23063) );
  INV_X1 U23527 ( .A(n23074), .ZN(n23079) );
  OAI21_X1 U23528 ( .B1(n23076), .B2(n23079), .A(n25179), .ZN(n23071) );
  NOR2_X1 U23529 ( .A1(n23064), .A2(n23077), .ZN(n23068) );
  NOR2_X1 U23530 ( .A1(n23077), .A2(n25452), .ZN(n23067) );
  AOI22_X1 U23531 ( .A1(n23069), .A2(n23068), .B1(n23067), .B2(n23066), .ZN(
        n23070) );
  XNOR2_X1 U23533 ( .A(n23073), .B(n23072), .ZN(Ciphertext[6]) );
  AOI21_X1 U23534 ( .B1(n25179), .B2(n25024), .A(n23074), .ZN(n23082) );
  NAND2_X1 U23535 ( .A1(n23076), .A2(n22578), .ZN(n23081) );
  NAND3_X1 U23536 ( .A1(n23079), .A2(n25024), .A3(n23077), .ZN(n23080) );
  NOR2_X1 U23537 ( .A1(n23119), .A2(n23120), .ZN(n23085) );
  AOI21_X1 U23538 ( .B1(n23123), .B2(n24941), .A(n23085), .ZN(n23126) );
  OAI211_X1 U23539 ( .C1(n23094), .C2(n24941), .A(n23112), .B(n24993), .ZN(
        n23086) );
  OAI21_X1 U23540 ( .B1(n23126), .B2(n23093), .A(n23086), .ZN(n23088) );
  INV_X1 U23541 ( .A(n2241), .ZN(n23087) );
  XNOR2_X1 U23542 ( .A(n23088), .B(n23087), .ZN(Ciphertext[13]) );
  MUX2_X1 U23543 ( .A(n23112), .B(n23125), .S(n23104), .Z(n23089) );
  NOR2_X1 U23544 ( .A1(n24941), .A2(n5036), .ZN(n23090) );
  NAND2_X1 U23545 ( .A1(n23090), .A2(n23112), .ZN(n23097) );
  NAND2_X1 U23546 ( .A1(n24993), .A2(n23112), .ZN(n23091) );
  NAND2_X1 U23547 ( .A1(n23094), .A2(n23093), .ZN(n23095) );
  NAND3_X1 U23548 ( .A1(n23097), .A2(n23096), .A3(n23095), .ZN(n23099) );
  INV_X1 U23549 ( .A(n2745), .ZN(n23098) );
  XNOR2_X1 U23550 ( .A(n23099), .B(n23098), .ZN(Ciphertext[15]) );
  NAND2_X1 U23551 ( .A1(n23120), .A2(n859), .ZN(n23102) );
  INV_X1 U23552 ( .A(n859), .ZN(n23108) );
  NAND3_X1 U23553 ( .A1(n24059), .A2(n23120), .A3(n23108), .ZN(n23101) );
  NOR2_X1 U23554 ( .A1(n23120), .A2(n859), .ZN(n23113) );
  NAND2_X1 U23555 ( .A1(n23112), .A2(n23113), .ZN(n23100) );
  OAI211_X1 U23556 ( .C1(n24059), .C2(n23102), .A(n23101), .B(n23100), .ZN(
        n23106) );
  NAND3_X1 U23557 ( .A1(n24498), .A2(n859), .A3(n5036), .ZN(n23103) );
  NOR2_X1 U23558 ( .A1(n23103), .A2(n23112), .ZN(n23105) );
  OAI21_X1 U23559 ( .B1(n23106), .B2(n23105), .A(n23104), .ZN(n23118) );
  XNOR2_X1 U23560 ( .A(n23125), .B(n859), .ZN(n23107) );
  NAND3_X1 U23561 ( .A1(n23123), .A2(n24498), .A3(n23107), .ZN(n23117) );
  NOR2_X1 U23562 ( .A1(n24498), .A2(n23108), .ZN(n23109) );
  OAI211_X1 U23563 ( .C1(n23120), .C2(n23112), .A(n23123), .B(n23109), .ZN(
        n23116) );
  NOR2_X1 U23564 ( .A1(n23112), .A2(n24498), .ZN(n23114) );
  NAND2_X1 U23565 ( .A1(n23114), .A2(n23113), .ZN(n23115) );
  NAND4_X1 U23566 ( .A1(n23118), .A2(n23117), .A3(n23116), .A4(n23115), .ZN(
        Ciphertext[16]) );
  INV_X1 U23567 ( .A(n24993), .ZN(n23121) );
  AOI21_X1 U23568 ( .B1(n23122), .B2(n23121), .A(n23120), .ZN(n23124) );
  OAI22_X1 U23569 ( .A1(n23126), .A2(n23125), .B1(n23124), .B2(n23123), .ZN(
        n23128) );
  INV_X1 U23570 ( .A(n3093), .ZN(n23127) );
  XNOR2_X1 U23571 ( .A(n23128), .B(n23127), .ZN(Ciphertext[17]) );
  INV_X1 U23572 ( .A(n23157), .ZN(n23131) );
  INV_X1 U23573 ( .A(n23154), .ZN(n23139) );
  OAI21_X1 U23575 ( .B1(n23133), .B2(n22442), .A(n23132), .ZN(n23134) );
  INV_X1 U23576 ( .A(n23134), .ZN(n23136) );
  OAI21_X1 U23577 ( .B1(n23160), .B2(n23155), .A(n24906), .ZN(n23135) );
  INV_X1 U23578 ( .A(n2761), .ZN(n23137) );
  AND2_X1 U23579 ( .A1(n24473), .A2(n23155), .ZN(n23158) );
  NAND2_X1 U23580 ( .A1(n23158), .A2(n23143), .ZN(n23141) );
  OAI211_X1 U23581 ( .C1(n23146), .C2(n1349), .A(n23139), .B(n23138), .ZN(
        n23140) );
  OAI211_X1 U23582 ( .C1(n24325), .C2(n23143), .A(n23141), .B(n23140), .ZN(
        n23142) );
  XNOR2_X1 U23583 ( .A(n23142), .B(n1528), .ZN(Ciphertext[19]) );
  OAI21_X1 U23584 ( .B1(n22442), .B2(n1349), .A(n23143), .ZN(n23150) );
  NOR2_X1 U23585 ( .A1(n24325), .A2(n24906), .ZN(n23149) );
  NAND3_X1 U23586 ( .A1(n23147), .A2(n23146), .A3(n23145), .ZN(n23148) );
  OAI21_X1 U23587 ( .B1(n23150), .B2(n23149), .A(n23148), .ZN(n23152) );
  XNOR2_X1 U23588 ( .A(n23152), .B(n23151), .ZN(Ciphertext[20]) );
  NAND2_X1 U23589 ( .A1(n23154), .A2(n24473), .ZN(n23156) );
  NAND2_X1 U23590 ( .A1(n23156), .A2(n23155), .ZN(n23159) );
  AOI22_X1 U23591 ( .A1(n24325), .A2(n23159), .B1(n23158), .B2(n1349), .ZN(
        n23162) );
  NAND2_X1 U23592 ( .A1(n23160), .A2(n22442), .ZN(n23161) );
  NAND2_X1 U23593 ( .A1(n23162), .A2(n23161), .ZN(n23163) );
  XNOR2_X1 U23594 ( .A(n23163), .B(n14879), .ZN(Ciphertext[23]) );
  AND2_X1 U23595 ( .A1(n23178), .A2(n23164), .ZN(n23174) );
  NOR2_X1 U23596 ( .A1(n23165), .A2(n23166), .ZN(n23175) );
  AOI21_X1 U23597 ( .B1(n23174), .B2(n23166), .A(n23175), .ZN(n23171) );
  NAND2_X1 U23598 ( .A1(n23181), .A2(n23166), .ZN(n23169) );
  NAND3_X1 U23599 ( .A1(n23169), .A2(n23168), .A3(n23167), .ZN(n23170) );
  NAND2_X1 U23600 ( .A1(n23171), .A2(n23170), .ZN(n23173) );
  INV_X1 U23601 ( .A(n923), .ZN(n23172) );
  XNOR2_X1 U23602 ( .A(n23173), .B(n23172), .ZN(Ciphertext[25]) );
  NOR2_X1 U23603 ( .A1(n23175), .A2(n23174), .ZN(n23182) );
  AOI21_X1 U23604 ( .B1(n23178), .B2(n24394), .A(n23176), .ZN(n23180) );
  NAND2_X1 U23605 ( .A1(n23186), .A2(n23206), .ZN(n23190) );
  NAND3_X1 U23606 ( .A1(n23201), .A2(n23202), .A3(n25059), .ZN(n23189) );
  INV_X1 U23607 ( .A(n24889), .ZN(n23185) );
  OAI21_X1 U23608 ( .B1(n25059), .B2(n24334), .A(n23185), .ZN(n23187) );
  NAND2_X1 U23609 ( .A1(n23187), .A2(n23194), .ZN(n23188) );
  INV_X1 U23610 ( .A(n2903), .ZN(n23207) );
  XNOR2_X1 U23611 ( .A(n23186), .B(n23207), .ZN(n23199) );
  NAND3_X1 U23612 ( .A1(n23194), .A2(n23207), .A3(n23193), .ZN(n23195) );
  NOR2_X1 U23614 ( .A1(n23202), .A2(n23201), .ZN(n23204) );
  INV_X1 U23616 ( .A(n23208), .ZN(n23205) );
  NAND3_X1 U23618 ( .A1(n23208), .A2(n23207), .A3(n23206), .ZN(n23209) );
  AND3_X1 U23619 ( .A1(n23211), .A2(n23210), .A3(n23209), .ZN(Ciphertext[32])
         );
  NOR2_X1 U23620 ( .A1(n23227), .A2(n25367), .ZN(n23212) );
  OAI211_X1 U23621 ( .C1(n23213), .C2(n23219), .A(n24955), .B(n23227), .ZN(
        n23214) );
  OAI21_X1 U23622 ( .B1(n23232), .B2(n23215), .A(n23214), .ZN(n23216) );
  XNOR2_X1 U23623 ( .A(n23216), .B(n5433), .ZN(Ciphertext[37]) );
  MUX2_X1 U23624 ( .A(n1340), .B(n23218), .S(n23217), .Z(n23224) );
  OAI21_X1 U23626 ( .B1(n23224), .B2(n25367), .A(n23223), .ZN(n23226) );
  XNOR2_X1 U23627 ( .A(n23226), .B(n23225), .ZN(Ciphertext[40]) );
  AOI21_X1 U23628 ( .B1(n317), .B2(n23229), .A(n25367), .ZN(n23230) );
  OAI22_X1 U23629 ( .A1(n23232), .A2(n23231), .B1(n23218), .B2(n23230), .ZN(
        n23234) );
  INV_X1 U23630 ( .A(n2036), .ZN(n23233) );
  XNOR2_X1 U23631 ( .A(n23234), .B(n23233), .ZN(Ciphertext[41]) );
  OAI21_X1 U23632 ( .B1(n23235), .B2(n23254), .A(n24377), .ZN(n23238) );
  NAND3_X1 U23633 ( .A1(n23236), .A2(n23241), .A3(n23250), .ZN(n23237) );
  AND2_X1 U23634 ( .A1(n23242), .A2(n23250), .ZN(n23253) );
  NAND2_X1 U23635 ( .A1(n23253), .A2(n23245), .ZN(n23243) );
  OAI211_X1 U23636 ( .C1(n189), .C2(n23245), .A(n23244), .B(n23243), .ZN(
        n23248) );
  INV_X1 U23637 ( .A(n1835), .ZN(n23247) );
  XNOR2_X1 U23638 ( .A(n23248), .B(n23247), .ZN(Ciphertext[43]) );
  AOI21_X1 U23639 ( .B1(n24377), .B2(n23250), .A(n23249), .ZN(n23255) );
  INV_X1 U23640 ( .A(n2190), .ZN(n23257) );
  MUX2_X1 U23641 ( .A(n24349), .B(n23274), .S(n23273), .Z(n23261) );
  AND2_X1 U23642 ( .A1(n23275), .A2(n24349), .ZN(n23258) );
  AOI22_X1 U23643 ( .A1(n23259), .A2(n23281), .B1(n23258), .B2(n24360), .ZN(
        n23260) );
  OAI21_X1 U23644 ( .B1(n23261), .B2(n23281), .A(n23260), .ZN(n23262) );
  XNOR2_X1 U23645 ( .A(n23262), .B(n2964), .ZN(Ciphertext[51]) );
  AND2_X1 U23646 ( .A1(n23277), .A2(n24349), .ZN(n23266) );
  NOR2_X1 U23647 ( .A1(n23275), .A2(n24349), .ZN(n23264) );
  AOI22_X1 U23648 ( .A1(n23267), .A2(n23266), .B1(n23265), .B2(n23264), .ZN(
        n23270) );
  NAND2_X1 U23649 ( .A1(n24907), .A2(n23275), .ZN(n23268) );
  OAI211_X1 U23650 ( .C1(n24360), .C2(n24486), .A(n23281), .B(n23268), .ZN(
        n23269) );
  NAND2_X1 U23651 ( .A1(n23270), .A2(n23269), .ZN(n23272) );
  XNOR2_X1 U23652 ( .A(n23272), .B(n23271), .ZN(Ciphertext[52]) );
  NOR2_X1 U23653 ( .A1(n23274), .A2(n23273), .ZN(n23276) );
  OAI21_X1 U23654 ( .B1(n23276), .B2(n24486), .A(n23281), .ZN(n23280) );
  NAND3_X1 U23655 ( .A1(n23278), .A2(n24907), .A3(n23277), .ZN(n23279) );
  OAI211_X1 U23656 ( .C1(n23282), .C2(n23281), .A(n23280), .B(n23279), .ZN(
        n23284) );
  XNOR2_X1 U23657 ( .A(n23284), .B(n23283), .ZN(Ciphertext[53]) );
  NOR2_X1 U23658 ( .A1(n24903), .A2(n23294), .ZN(n23286) );
  OAI21_X1 U23659 ( .B1(n23298), .B2(n23286), .A(n23308), .ZN(n23289) );
  OAI21_X1 U23660 ( .B1(n23292), .B2(n23308), .A(n23305), .ZN(n23287) );
  NAND2_X1 U23661 ( .A1(n23287), .A2(n23294), .ZN(n23288) );
  INV_X1 U23663 ( .A(n1924), .ZN(n23290) );
  XNOR2_X1 U23664 ( .A(n23291), .B(n23290), .ZN(Ciphertext[54]) );
  NAND2_X1 U23665 ( .A1(n23292), .A2(n23305), .ZN(n23296) );
  MUX2_X1 U23666 ( .A(n23296), .B(n23295), .S(n23294), .Z(n23301) );
  INV_X1 U23667 ( .A(n876), .ZN(n23302) );
  INV_X1 U23668 ( .A(n23303), .ZN(n23304) );
  OAI21_X1 U23669 ( .B1(n23306), .B2(n23305), .A(n23304), .ZN(n23307) );
  OAI21_X1 U23670 ( .B1(n23309), .B2(n23308), .A(n23307), .ZN(n23310) );
  XNOR2_X1 U23671 ( .A(n23310), .B(n3344), .ZN(Ciphertext[59]) );
  OAI21_X1 U23672 ( .B1(n4108), .B2(n23318), .A(n24316), .ZN(n23312) );
  NAND3_X1 U23673 ( .A1(n23313), .A2(n23326), .A3(n23317), .ZN(n23314) );
  INV_X1 U23674 ( .A(n912), .ZN(n23315) );
  XNOR2_X1 U23675 ( .A(n23316), .B(n23315), .ZN(Ciphertext[60]) );
  OAI211_X1 U23676 ( .C1(n23320), .C2(n5659), .A(n23319), .B(n23326), .ZN(
        n23321) );
  XNOR2_X1 U23677 ( .A(n23323), .B(n23322), .ZN(Ciphertext[64]) );
  NAND2_X1 U23678 ( .A1(n23325), .A2(n24316), .ZN(n23329) );
  XNOR2_X1 U23680 ( .A(n23331), .B(n23330), .ZN(Ciphertext[65]) );
  AOI21_X1 U23681 ( .B1(n25081), .B2(n24341), .A(n25004), .ZN(n23339) );
  NAND2_X1 U23682 ( .A1(n24342), .A2(n5421), .ZN(n23337) );
  NOR2_X1 U23683 ( .A1(n23334), .A2(n25081), .ZN(n23335) );
  AOI21_X1 U23684 ( .B1(n23337), .B2(n25081), .A(n23335), .ZN(n23338) );
  OAI21_X1 U23685 ( .B1(n23339), .B2(n23338), .A(n1397), .ZN(n23341) );
  AOI21_X1 U23686 ( .B1(n24492), .B2(n23341), .A(n23340), .ZN(n23346) );
  AOI21_X1 U23687 ( .B1(n24400), .B2(n24492), .A(n23350), .ZN(n23345) );
  NOR2_X1 U23688 ( .A1(n23354), .A2(n22961), .ZN(n23360) );
  NOR2_X1 U23689 ( .A1(n24400), .A2(n23359), .ZN(n23343) );
  OAI21_X1 U23690 ( .B1(n23360), .B2(n23343), .A(n23349), .ZN(n23344) );
  OAI21_X1 U23691 ( .B1(n23346), .B2(n23345), .A(n23344), .ZN(n23348) );
  XNOR2_X1 U23692 ( .A(n23348), .B(n23347), .ZN(Ciphertext[68]) );
  INV_X1 U23695 ( .A(n23359), .ZN(n23353) );
  OAI21_X1 U23696 ( .B1(n24343), .B2(n23353), .A(n23350), .ZN(n23356) );
  XNOR2_X1 U23697 ( .A(n23358), .B(n3115), .ZN(Ciphertext[70]) );
  OAI21_X1 U23698 ( .B1(n23360), .B2(n23359), .A(n23350), .ZN(n23365) );
  INV_X1 U23699 ( .A(n889), .ZN(n23366) );
  XNOR2_X1 U23700 ( .A(n23367), .B(n23366), .ZN(Ciphertext[71]) );
  NAND2_X1 U23701 ( .A1(n23370), .A2(n23368), .ZN(n23378) );
  NAND3_X1 U23702 ( .A1(n23370), .A2(n23371), .A3(n24412), .ZN(n23377) );
  INV_X1 U23703 ( .A(n23371), .ZN(n23373) );
  AOI22_X1 U23704 ( .A1(n23375), .A2(n23374), .B1(n23373), .B2(n23372), .ZN(
        n23376) );
  OAI211_X1 U23705 ( .C1(n23379), .C2(n23378), .A(n23377), .B(n23376), .ZN(
        n23381) );
  INV_X1 U23706 ( .A(n836), .ZN(n23380) );
  XNOR2_X1 U23707 ( .A(n23381), .B(n23380), .ZN(Ciphertext[72]) );
  MUX2_X1 U23708 ( .A(n23396), .B(n23394), .S(n23391), .Z(n23383) );
  MUX2_X1 U23709 ( .A(n24933), .B(n23393), .S(n24880), .Z(n23382) );
  MUX2_X1 U23710 ( .A(n23383), .B(n23382), .S(n23392), .Z(n23384) );
  XNOR2_X1 U23711 ( .A(n23384), .B(n5251), .ZN(Ciphertext[80]) );
  AOI22_X1 U23712 ( .A1(n24880), .A2(n23386), .B1(n23392), .B2(n23394), .ZN(
        n23388) );
  NOR3_X1 U23713 ( .A1(n24449), .A2(n22026), .A3(n23396), .ZN(n23387) );
  AOI21_X1 U23714 ( .B1(n23388), .B2(n23389), .A(n23387), .ZN(n23390) );
  XNOR2_X1 U23715 ( .A(n23390), .B(n1891), .ZN(Ciphertext[81]) );
  MUX2_X1 U23716 ( .A(n24880), .B(n22026), .S(n24449), .Z(n23397) );
  INV_X1 U23718 ( .A(n23410), .ZN(n23417) );
  NAND3_X1 U23719 ( .A1(n906), .A2(n25035), .A3(n24426), .ZN(n23399) );
  INV_X1 U23720 ( .A(n2208), .ZN(n23401) );
  INV_X1 U23721 ( .A(n23416), .ZN(n23402) );
  AOI22_X1 U23722 ( .A1(n23402), .A2(n23417), .B1(n23420), .B2(n23411), .ZN(
        n23422) );
  NAND2_X1 U23723 ( .A1(n24977), .A2(n23398), .ZN(n23404) );
  NAND3_X1 U23724 ( .A1(n23404), .A2(n25035), .A3(n24947), .ZN(n23405) );
  OAI21_X1 U23725 ( .B1(n23422), .B2(n23406), .A(n23405), .ZN(n23408) );
  INV_X1 U23726 ( .A(n1776), .ZN(n23407) );
  XNOR2_X1 U23727 ( .A(n23408), .B(n23407), .ZN(Ciphertext[85]) );
  NAND2_X1 U23728 ( .A1(n23416), .A2(n23410), .ZN(n23413) );
  AOI21_X1 U23729 ( .B1(n23418), .B2(n23417), .A(n23416), .ZN(n23419) );
  OAI22_X1 U23730 ( .A1(n23422), .A2(n24426), .B1(n23420), .B2(n23419), .ZN(
        n23424) );
  INV_X1 U23731 ( .A(n2031), .ZN(n23423) );
  XNOR2_X1 U23732 ( .A(n23424), .B(n23423), .ZN(Ciphertext[89]) );
  NAND3_X1 U23733 ( .A1(n23449), .A2(n22528), .A3(n23443), .ZN(n23429) );
  OAI21_X1 U23734 ( .B1(n23449), .B2(n23425), .A(n23442), .ZN(n23433) );
  NAND2_X1 U23735 ( .A1(n23433), .A2(n22506), .ZN(n23427) );
  NOR2_X1 U23736 ( .A1(n24989), .A2(n1370), .ZN(n23426) );
  NAND2_X1 U23737 ( .A1(n23449), .A2(n23426), .ZN(n23428) );
  NAND4_X1 U23738 ( .A1(n23429), .A2(n23427), .A3(n2211), .A4(n23428), .ZN(
        n23436) );
  INV_X1 U23739 ( .A(n23428), .ZN(n23431) );
  INV_X1 U23740 ( .A(n23429), .ZN(n23430) );
  OAI21_X1 U23741 ( .B1(n23431), .B2(n23430), .A(n23432), .ZN(n23435) );
  NAND3_X1 U23742 ( .A1(n23433), .A2(n23432), .A3(n22506), .ZN(n23434) );
  NAND3_X1 U23743 ( .A1(n23436), .A2(n23435), .A3(n23434), .ZN(Ciphertext[90])
         );
  AOI21_X1 U23744 ( .B1(n23449), .B2(n23425), .A(n23437), .ZN(n23439) );
  NAND3_X1 U23745 ( .A1(n23437), .A2(n22528), .A3(n23443), .ZN(n23438) );
  OAI21_X1 U23746 ( .B1(n23439), .B2(n23453), .A(n23438), .ZN(n23440) );
  XNOR2_X1 U23747 ( .A(n23440), .B(n494), .ZN(Ciphertext[91]) );
  NAND3_X1 U23748 ( .A1(n321), .A2(n23450), .A3(n22528), .ZN(n23446) );
  NAND3_X1 U23749 ( .A1(n23442), .A2(n1370), .A3(n22528), .ZN(n23445) );
  INV_X1 U23750 ( .A(n23449), .ZN(n23452) );
  OAI21_X1 U23751 ( .B1(n23450), .B2(n1370), .A(n321), .ZN(n23451) );
  AOI22_X1 U23752 ( .A1(n23453), .A2(n23452), .B1(n23451), .B2(n22528), .ZN(
        n23454) );
  XNOR2_X1 U23753 ( .A(n23454), .B(n2240), .ZN(Ciphertext[95]) );
  MUX2_X1 U23754 ( .A(n23491), .B(n23481), .S(n23480), .Z(n23456) );
  OAI21_X1 U23755 ( .B1(n23499), .B2(n23494), .A(n24336), .ZN(n23455) );
  AOI21_X1 U23758 ( .B1(n23458), .B2(n23461), .A(n23464), .ZN(n23466) );
  NAND2_X1 U23759 ( .A1(n23460), .A2(n24364), .ZN(n23465) );
  AOI22_X1 U23761 ( .A1(n23466), .A2(n23465), .B1(n25055), .B2(n23463), .ZN(
        n23468) );
  NAND2_X1 U23763 ( .A1(n23483), .A2(n23472), .ZN(n23475) );
  NAND2_X1 U23765 ( .A1(n23011), .A2(n23472), .ZN(n23471) );
  OAI211_X1 U23766 ( .C1(n24442), .C2(n23472), .A(n23471), .B(n24336), .ZN(
        n23473) );
  OAI211_X1 U23767 ( .C1(n23499), .C2(n23475), .A(n23474), .B(n23473), .ZN(
        n23477) );
  XNOR2_X1 U23768 ( .A(n23477), .B(n23476), .ZN(Ciphertext[98]) );
  AND2_X1 U23769 ( .A1(n23479), .A2(n23478), .ZN(n23490) );
  NOR2_X1 U23770 ( .A1(n23480), .A2(n23479), .ZN(n23482) );
  AOI22_X1 U23771 ( .A1(n23490), .A2(n23499), .B1(n23482), .B2(n23481), .ZN(
        n23488) );
  OAI211_X1 U23773 ( .C1(n24442), .C2(n24336), .A(n23485), .B(n23484), .ZN(
        n23487) );
  INV_X1 U23774 ( .A(n2882), .ZN(n23489) );
  INV_X1 U23775 ( .A(n23490), .ZN(n23498) );
  NAND2_X1 U23776 ( .A1(n23493), .A2(n23499), .ZN(n23497) );
  NAND2_X1 U23777 ( .A1(n23495), .A2(n23494), .ZN(n23496) );
  OAI211_X1 U23778 ( .C1(n23499), .C2(n23498), .A(n23497), .B(n23496), .ZN(
        n23501) );
  XNOR2_X1 U23779 ( .A(n23501), .B(n23500), .ZN(Ciphertext[101]) );
  NOR2_X1 U23780 ( .A1(n24351), .A2(n23505), .ZN(n23504) );
  INV_X1 U23781 ( .A(n23527), .ZN(n23503) );
  OAI21_X1 U23782 ( .B1(n23510), .B2(n23505), .A(n24380), .ZN(n23506) );
  OAI21_X1 U23783 ( .B1(n23527), .B2(n24313), .A(n23506), .ZN(n23507) );
  XNOR2_X1 U23784 ( .A(n23509), .B(n23508), .ZN(Ciphertext[102]) );
  NOR2_X1 U23785 ( .A1(n23527), .A2(n23530), .ZN(n23512) );
  NOR2_X1 U23786 ( .A1(n24351), .A2(n23510), .ZN(n23511) );
  NAND2_X1 U23787 ( .A1(n23513), .A2(n23531), .ZN(n23521) );
  NOR2_X1 U23788 ( .A1(n23514), .A2(n24313), .ZN(n23519) );
  NOR3_X1 U23789 ( .A1(n23517), .A2(n23516), .A3(n23515), .ZN(n23518) );
  NAND2_X1 U23790 ( .A1(n23519), .A2(n23518), .ZN(n23520) );
  OAI211_X1 U23791 ( .C1(n23522), .C2(n23531), .A(n23521), .B(n23520), .ZN(
        n23524) );
  XNOR2_X1 U23792 ( .A(n23524), .B(n23523), .ZN(Ciphertext[105]) );
  INV_X1 U23793 ( .A(n24313), .ZN(n23526) );
  NOR3_X1 U23794 ( .A1(n23527), .A2(n23526), .A3(n24351), .ZN(n23528) );
  OR2_X1 U23795 ( .A1(n23530), .A2(n23529), .ZN(n23532) );
  XNOR2_X1 U23796 ( .A(n23534), .B(n2739), .ZN(Ciphertext[106]) );
  NOR2_X1 U23797 ( .A1(n23546), .A2(n23547), .ZN(n23563) );
  INV_X1 U23798 ( .A(n23563), .ZN(n23540) );
  NAND2_X1 U23799 ( .A1(n23537), .A2(n23554), .ZN(n23535) );
  OAI21_X1 U23800 ( .B1(n25071), .B2(n23537), .A(n23535), .ZN(n23536) );
  INV_X1 U23801 ( .A(n23555), .ZN(n23538) );
  NAND3_X1 U23802 ( .A1(n23538), .A2(n25071), .A3(n23537), .ZN(n23539) );
  INV_X1 U23803 ( .A(n1364), .ZN(n23541) );
  XNOR2_X1 U23804 ( .A(n23542), .B(n23541), .ZN(Ciphertext[108]) );
  INV_X1 U23805 ( .A(n23554), .ZN(n23556) );
  OAI21_X1 U23806 ( .B1(n23555), .B2(n24057), .A(n23556), .ZN(n23550) );
  NAND3_X1 U23809 ( .A1(n323), .A2(n23547), .A3(n25071), .ZN(n23548) );
  OAI211_X1 U23810 ( .C1(n23551), .C2(n23550), .A(n23549), .B(n23548), .ZN(
        n23553) );
  INV_X1 U23811 ( .A(n1826), .ZN(n23552) );
  XNOR2_X1 U23812 ( .A(n23553), .B(n23552), .ZN(Ciphertext[111]) );
  OAI21_X1 U23813 ( .B1(n24893), .B2(n23555), .A(n23554), .ZN(n23562) );
  NAND3_X1 U23814 ( .A1(n23557), .A2(n23556), .A3(n323), .ZN(n23561) );
  NAND2_X1 U23815 ( .A1(n23563), .A2(n24057), .ZN(n23560) );
  INV_X1 U23816 ( .A(n1920), .ZN(n23564) );
  NOR2_X1 U23817 ( .A1(n23592), .A2(n23566), .ZN(n23597) );
  INV_X1 U23818 ( .A(n23597), .ZN(n23569) );
  OAI211_X1 U23819 ( .C1(n1328), .C2(n23596), .A(n24389), .B(n23565), .ZN(
        n23568) );
  NAND3_X1 U23820 ( .A1(n23595), .A2(n23566), .A3(n24901), .ZN(n23567) );
  NAND3_X1 U23821 ( .A1(n23569), .A2(n23568), .A3(n23567), .ZN(n23570) );
  XNOR2_X1 U23822 ( .A(n23570), .B(n4589), .ZN(Ciphertext[115]) );
  OR2_X1 U23823 ( .A1(n23573), .A2(n23572), .ZN(n23581) );
  AND2_X1 U23824 ( .A1(n23576), .A2(n23577), .ZN(n23582) );
  NOR4_X1 U23825 ( .A1(n23579), .A2(n23581), .A3(n23578), .A4(n23582), .ZN(
        n23580) );
  NAND2_X1 U23826 ( .A1(n23580), .A2(n23591), .ZN(n23588) );
  OAI21_X1 U23827 ( .B1(n23582), .B2(n23581), .A(n23594), .ZN(n23583) );
  OAI21_X1 U23828 ( .B1(n24389), .B2(n24901), .A(n23583), .ZN(n23585) );
  NAND2_X1 U23829 ( .A1(n23585), .A2(n21941), .ZN(n23587) );
  XNOR2_X1 U23830 ( .A(n23590), .B(n23589), .ZN(Ciphertext[117]) );
  NAND2_X1 U23831 ( .A1(n23591), .A2(n23592), .ZN(n23601) );
  NAND3_X1 U23832 ( .A1(n24611), .A2(n23592), .A3(n24901), .ZN(n23600) );
  NAND3_X1 U23833 ( .A1(n23595), .A2(n23596), .A3(n24901), .ZN(n23599) );
  NAND2_X1 U23834 ( .A1(n23597), .A2(n23596), .ZN(n23598) );
  NAND4_X1 U23835 ( .A1(n23601), .A2(n23600), .A3(n23599), .A4(n23598), .ZN(
        n23603) );
  XNOR2_X1 U23836 ( .A(n23603), .B(n23602), .ZN(Ciphertext[119]) );
  INV_X1 U23837 ( .A(n23650), .ZN(n23627) );
  NAND3_X1 U23838 ( .A1(n23627), .A2(n23647), .A3(n23645), .ZN(n23605) );
  NAND4_X1 U23839 ( .A1(n24320), .A2(n23650), .A3(n20896), .A4(n23637), .ZN(
        n23604) );
  OAI211_X1 U23840 ( .C1(n23606), .C2(n23645), .A(n23605), .B(n23604), .ZN(
        n23608) );
  INV_X1 U23841 ( .A(n2805), .ZN(n23607) );
  XNOR2_X1 U23842 ( .A(n23608), .B(n23607), .ZN(Ciphertext[121]) );
  NAND2_X1 U23843 ( .A1(n23612), .A2(n23620), .ZN(n23609) );
  INV_X1 U23844 ( .A(n23609), .ZN(n23610) );
  OAI211_X1 U23845 ( .C1(n23620), .C2(n24320), .A(n23609), .B(n23653), .ZN(
        n23618) );
  INV_X1 U23846 ( .A(n23647), .ZN(n23651) );
  NAND2_X1 U23847 ( .A1(n23610), .A2(n23651), .ZN(n23616) );
  NOR2_X1 U23848 ( .A1(n23648), .A2(n23620), .ZN(n23611) );
  AOI21_X1 U23849 ( .B1(n23611), .B2(n23647), .A(n23645), .ZN(n23615) );
  INV_X1 U23850 ( .A(n23620), .ZN(n23624) );
  XNOR2_X1 U23851 ( .A(n23650), .B(n23624), .ZN(n23613) );
  OR2_X1 U23852 ( .A1(n23613), .A2(n24320), .ZN(n23614) );
  NAND3_X1 U23853 ( .A1(n23616), .A2(n23615), .A3(n23614), .ZN(n23617) );
  NAND2_X1 U23854 ( .A1(n23618), .A2(n23617), .ZN(n23626) );
  NAND2_X1 U23855 ( .A1(n23619), .A2(n23620), .ZN(n23622) );
  NAND2_X1 U23856 ( .A1(n23634), .A2(n23620), .ZN(n23621) );
  NAND4_X1 U23857 ( .A1(n23622), .A2(n23645), .A3(n23649), .A4(n23621), .ZN(
        n23623) );
  AOI21_X1 U23858 ( .B1(n23652), .B2(n23624), .A(n23623), .ZN(n23625) );
  NOR2_X1 U23859 ( .A1(n23626), .A2(n23625), .ZN(Ciphertext[122]) );
  NAND2_X1 U23860 ( .A1(n23627), .A2(n23645), .ZN(n23638) );
  NOR2_X1 U23861 ( .A1(n23647), .A2(n23648), .ZN(n23628) );
  NAND2_X1 U23862 ( .A1(n23628), .A2(n23645), .ZN(n23632) );
  NAND3_X1 U23863 ( .A1(n23629), .A2(n23637), .A3(n23649), .ZN(n23630) );
  NAND4_X1 U23864 ( .A1(n23631), .A2(n3164), .A3(n23632), .A4(n23630), .ZN(
        n23644) );
  INV_X1 U23866 ( .A(n3164), .ZN(n23639) );
  INV_X1 U23868 ( .A(n23645), .ZN(n23636) );
  NOR2_X1 U23869 ( .A1(n23634), .A2(n3164), .ZN(n23635) );
  NAND4_X1 U23870 ( .A1(n23637), .A2(n23636), .A3(n23635), .A4(n23649), .ZN(
        n23642) );
  NAND4_X1 U23871 ( .A1(n23644), .A2(n23643), .A3(n23642), .A4(n23641), .ZN(
        Ciphertext[123]) );
  NAND2_X1 U23872 ( .A1(n23648), .A2(n23645), .ZN(n23646) );
  OAI211_X1 U23873 ( .C1(n23648), .C2(n23649), .A(n23647), .B(n23646), .ZN(
        n23656) );
  NAND3_X1 U23874 ( .A1(n23651), .A2(n23650), .A3(n23649), .ZN(n23655) );
  NAND2_X1 U23875 ( .A1(n23653), .A2(n23652), .ZN(n23654) );
  INV_X1 U23876 ( .A(n1746), .ZN(n23657) );
  AND2_X1 U23877 ( .A1(n23658), .A2(n25026), .ZN(n23662) );
  NAND2_X1 U23878 ( .A1(n23665), .A2(n23689), .ZN(n23661) );
  AND2_X1 U23879 ( .A1(n23659), .A2(n25026), .ZN(n23660) );
  XNOR2_X1 U23880 ( .A(n23664), .B(n23663), .ZN(Ciphertext[127]) );
  INV_X1 U23881 ( .A(n23679), .ZN(n23666) );
  NOR3_X1 U23882 ( .A1(n23669), .A2(n23668), .A3(n23678), .ZN(n23685) );
  AOI21_X1 U23883 ( .B1(n23671), .B2(n23679), .A(n23670), .ZN(n23675) );
  OR3_X1 U23884 ( .A1(n23672), .A2(n23679), .A3(n23671), .ZN(n23674) );
  NAND2_X1 U23885 ( .A1(n23672), .A2(n23679), .ZN(n23673) );
  NAND3_X1 U23886 ( .A1(n23675), .A2(n23674), .A3(n23673), .ZN(n23684) );
  OR2_X1 U23887 ( .A1(n23692), .A2(n23679), .ZN(n23682) );
  INV_X1 U23888 ( .A(n23690), .ZN(n23677) );
  OAI21_X1 U23890 ( .B1(n23682), .B2(n23681), .A(n23680), .ZN(n23683) );
  INV_X1 U23891 ( .A(n23699), .ZN(n23703) );
  NOR2_X1 U23892 ( .A1(n23714), .A2(n23703), .ZN(n23705) );
  INV_X1 U23893 ( .A(n23705), .ZN(n23695) );
  NAND3_X1 U23894 ( .A1(n5284), .A2(n23716), .A3(n23703), .ZN(n23694) );
  OAI21_X1 U23895 ( .B1(n23696), .B2(n23695), .A(n23694), .ZN(n23711) );
  NOR2_X1 U23896 ( .A1(n23715), .A2(n23699), .ZN(n23698) );
  NAND2_X1 U23897 ( .A1(n23714), .A2(n23703), .ZN(n23701) );
  NAND2_X1 U23898 ( .A1(n23712), .A2(n23699), .ZN(n23700) );
  OAI21_X1 U23899 ( .B1(n23712), .B2(n23701), .A(n23700), .ZN(n23708) );
  NAND2_X1 U23900 ( .A1(n23720), .A2(n23703), .ZN(n23702) );
  OAI21_X1 U23901 ( .B1(n23720), .B2(n23703), .A(n23702), .ZN(n23704) );
  NAND3_X1 U23902 ( .A1(n23704), .A2(n23715), .A3(n23714), .ZN(n23707) );
  OAI211_X1 U23903 ( .C1(n23709), .C2(n23708), .A(n23707), .B(n23706), .ZN(
        n23710) );
  AOI21_X1 U23904 ( .B1(n24374), .B2(n23711), .A(n23710), .ZN(Ciphertext[134])
         );
  INV_X1 U23905 ( .A(n23720), .ZN(n23713) );
  MUX2_X1 U23906 ( .A(n23715), .B(n23713), .S(n23712), .Z(n23718) );
  NAND3_X1 U23907 ( .A1(n23719), .A2(n23715), .A3(n23714), .ZN(n23717) );
  OAI21_X1 U23908 ( .B1(n23721), .B2(n23720), .A(n23719), .ZN(n23722) );
  NAND2_X1 U23909 ( .A1(n23724), .A2(n23723), .ZN(n23725) );
  INV_X1 U23910 ( .A(n1869), .ZN(n23729) );
  MUX2_X1 U23911 ( .A(n23743), .B(n23740), .S(n24065), .Z(n23732) );
  AOI22_X1 U23912 ( .A1(n23732), .A2(n23731), .B1(n24064), .B2(n23745), .ZN(
        n23734) );
  INV_X1 U23913 ( .A(n921), .ZN(n23733) );
  XNOR2_X1 U23914 ( .A(n23734), .B(n23733), .ZN(Ciphertext[138]) );
  OAI211_X1 U23915 ( .C1(n23745), .C2(n997), .A(n24065), .B(n23740), .ZN(
        n23736) );
  NAND2_X1 U23916 ( .A1(n23737), .A2(n23736), .ZN(n23739) );
  INV_X1 U23917 ( .A(n688), .ZN(n23738) );
  XNOR2_X1 U23918 ( .A(n23739), .B(n23738), .ZN(Ciphertext[139]) );
  MUX2_X1 U23919 ( .A(n25460), .B(n24063), .S(n23740), .Z(n23749) );
  NAND3_X1 U23920 ( .A1(n23743), .A2(n24064), .A3(n25460), .ZN(n23747) );
  NAND2_X1 U23921 ( .A1(n23745), .A2(n23744), .ZN(n23746) );
  OAI211_X1 U23922 ( .C1(n23749), .C2(n23748), .A(n23747), .B(n23746), .ZN(
        n23751) );
  XNOR2_X1 U23923 ( .A(n23751), .B(n23750), .ZN(Ciphertext[141]) );
  OAI21_X1 U23924 ( .B1(n23779), .B2(n23769), .A(n23758), .ZN(n23755) );
  NAND2_X1 U23925 ( .A1(n23779), .A2(n23768), .ZN(n23753) );
  OAI21_X1 U23926 ( .B1(n23765), .B2(n23782), .A(n23753), .ZN(n23754) );
  AOI21_X1 U23927 ( .B1(n23782), .B2(n23755), .A(n23754), .ZN(n23756) );
  XNOR2_X1 U23928 ( .A(n23756), .B(n1758), .ZN(Ciphertext[144]) );
  OAI21_X1 U23929 ( .B1(n24921), .B2(n23769), .A(n23781), .ZN(n23761) );
  OR3_X1 U23930 ( .A1(n23779), .A2(n23768), .A3(n24921), .ZN(n23760) );
  OR2_X1 U23931 ( .A1(n23758), .A2(n23782), .ZN(n23759) );
  OAI211_X1 U23932 ( .C1(n23762), .C2(n23761), .A(n23760), .B(n23759), .ZN(
        n23764) );
  XNOR2_X1 U23933 ( .A(n23764), .B(n23763), .ZN(Ciphertext[147]) );
  INV_X1 U23934 ( .A(n23779), .ZN(n23767) );
  INV_X1 U23935 ( .A(n23768), .ZN(n23777) );
  OAI21_X1 U23936 ( .B1(n23774), .B2(n23777), .A(n23773), .ZN(n23776) );
  XNOR2_X1 U23937 ( .A(n23776), .B(n23775), .ZN(Ciphertext[148]) );
  AOI21_X1 U23938 ( .B1(n23779), .B2(n23778), .A(n23777), .ZN(n23780) );
  OAI22_X1 U23939 ( .A1(n23783), .A2(n23782), .B1(n23781), .B2(n23780), .ZN(
        n23785) );
  INV_X1 U23940 ( .A(n2747), .ZN(n23784) );
  XNOR2_X1 U23941 ( .A(n23785), .B(n23784), .ZN(Ciphertext[149]) );
  OAI21_X1 U23942 ( .B1(n21837), .B2(n23789), .A(n23788), .ZN(n23809) );
  AND2_X1 U23943 ( .A1(n24895), .A2(n23798), .ZN(n23793) );
  AOI21_X1 U23944 ( .B1(n23790), .B2(n23798), .A(n23793), .ZN(n23791) );
  OAI21_X1 U23945 ( .B1(n23792), .B2(n23798), .A(n23791), .ZN(n23808) );
  NAND3_X1 U23946 ( .A1(n23796), .A2(n23793), .A3(n24307), .ZN(n23807) );
  NAND3_X1 U23947 ( .A1(n23796), .A2(n21837), .A3(n896), .ZN(n23804) );
  OAI211_X1 U23948 ( .C1(n24895), .C2(n23798), .A(n23796), .B(n24307), .ZN(
        n23803) );
  XNOR2_X1 U23949 ( .A(n24920), .B(n23798), .ZN(n23801) );
  NAND2_X1 U23950 ( .A1(n23801), .A2(n24983), .ZN(n23802) );
  NAND4_X1 U23951 ( .A1(n23805), .A2(n23804), .A3(n23803), .A4(n23802), .ZN(
        n23806) );
  OAI211_X1 U23952 ( .C1(n23809), .C2(n23808), .A(n23807), .B(n23806), .ZN(
        Ciphertext[154]) );
  AND2_X1 U23953 ( .A1(n23810), .A2(n23817), .ZN(n23824) );
  OAI21_X1 U23954 ( .B1(n24972), .B2(n23831), .A(n23824), .ZN(n23815) );
  AND2_X1 U23955 ( .A1(n23811), .A2(n23827), .ZN(n23832) );
  NOR2_X1 U23956 ( .A1(n23828), .A2(n23813), .ZN(n23812) );
  AOI21_X1 U23957 ( .B1(n23832), .B2(n23813), .A(n23812), .ZN(n23814) );
  INV_X1 U23958 ( .A(n641), .ZN(n23816) );
  OAI21_X1 U23959 ( .B1(n23817), .B2(n24972), .A(n23032), .ZN(n23823) );
  NAND2_X1 U23960 ( .A1(n23818), .A2(n23831), .ZN(n23822) );
  NOR2_X1 U23961 ( .A1(n23827), .A2(n24972), .ZN(n23820) );
  INV_X1 U23964 ( .A(n23827), .ZN(n23829) );
  OAI21_X1 U23965 ( .B1(n23830), .B2(n23829), .A(n23828), .ZN(n23837) );
  NAND2_X1 U23966 ( .A1(n23832), .A2(n23831), .ZN(n23836) );
  NAND2_X1 U23967 ( .A1(n23032), .A2(n23833), .ZN(n23835) );
  NAND3_X1 U23968 ( .A1(n23837), .A2(n23836), .A3(n23835), .ZN(n23838) );
  XNOR2_X1 U23969 ( .A(n23838), .B(n3696), .ZN(Ciphertext[161]) );
  INV_X1 U23970 ( .A(n23860), .ZN(n23866) );
  INV_X1 U23971 ( .A(n23857), .ZN(n23864) );
  NAND3_X1 U23972 ( .A1(n25240), .A2(n24428), .A3(n23864), .ZN(n23840) );
  INV_X1 U23973 ( .A(n1810), .ZN(n23841) );
  INV_X1 U23974 ( .A(n3183), .ZN(n23842) );
  NOR2_X1 U23975 ( .A1(n23857), .A2(n23842), .ZN(n23844) );
  AOI21_X1 U23976 ( .B1(n23844), .B2(n23843), .A(n23865), .ZN(n23850) );
  NOR2_X1 U23977 ( .A1(n23862), .A2(n3183), .ZN(n23846) );
  NAND2_X1 U23978 ( .A1(n23857), .A2(n23846), .ZN(n23849) );
  AOI21_X1 U23980 ( .B1(n24469), .B2(n23846), .A(n23853), .ZN(n23847) );
  OAI21_X1 U23982 ( .B1(n23853), .B2(n3183), .A(n24428), .ZN(n23852) );
  AOI211_X1 U23983 ( .C1(n3183), .C2(n23853), .A(n23866), .B(n23852), .ZN(
        n23854) );
  NOR3_X1 U23984 ( .A1(n23856), .A2(n23855), .A3(n23854), .ZN(Ciphertext[164])
         );
  NAND2_X1 U23985 ( .A1(n24469), .A2(n23857), .ZN(n23861) );
  NAND2_X1 U23986 ( .A1(n24428), .A2(n23865), .ZN(n23863) );
  OAI211_X1 U23987 ( .C1(n23866), .C2(n23865), .A(n23864), .B(n23863), .ZN(
        n23867) );
  INV_X1 U23988 ( .A(Key[190]), .ZN(n23868) );
  NOR2_X1 U23990 ( .A1(n23904), .A2(n23890), .ZN(n23907) );
  NAND2_X1 U23991 ( .A1(n23907), .A2(n23889), .ZN(n23871) );
  INV_X1 U23992 ( .A(n1827), .ZN(n23873) );
  XNOR2_X1 U23993 ( .A(n23874), .B(n23873), .ZN(Ciphertext[169]) );
  NAND2_X1 U23994 ( .A1(n23896), .A2(n23883), .ZN(n23875) );
  XNOR2_X1 U23996 ( .A(n23890), .B(n24624), .ZN(n23876) );
  OAI21_X1 U23997 ( .B1(n23876), .B2(n23879), .A(n23902), .ZN(n23877) );
  XNOR2_X1 U23998 ( .A(n23906), .B(n24624), .ZN(n23886) );
  NAND2_X1 U23999 ( .A1(n23905), .A2(n23889), .ZN(n23885) );
  NOR2_X1 U24000 ( .A1(n23905), .A2(n23902), .ZN(n23882) );
  NAND2_X1 U24001 ( .A1(n23903), .A2(n23883), .ZN(n23881) );
  NAND2_X1 U24002 ( .A1(n23888), .A2(n23906), .ZN(n23899) );
  NAND3_X1 U24003 ( .A1(n23890), .A2(n23889), .A3(n23903), .ZN(n23898) );
  NOR2_X1 U24004 ( .A1(n23894), .A2(n23905), .ZN(n23895) );
  OAI21_X1 U24005 ( .B1(n23896), .B2(n23902), .A(n23895), .ZN(n23897) );
  INV_X1 U24007 ( .A(n1724), .ZN(n23900) );
  XNOR2_X1 U24008 ( .A(n23901), .B(n23900), .ZN(Ciphertext[171]) );
  AOI21_X1 U24009 ( .B1(n23906), .B2(n23902), .A(n23905), .ZN(n23908) );
  XNOR2_X1 U24010 ( .A(n23910), .B(n5484), .ZN(Ciphertext[173]) );
  NAND2_X1 U24011 ( .A1(n23911), .A2(n25083), .ZN(n23936) );
  INV_X1 U24012 ( .A(n23937), .ZN(n23912) );
  NAND3_X1 U24013 ( .A1(n23912), .A2(n23926), .A3(n23933), .ZN(n23914) );
  NAND4_X1 U24014 ( .A1(n23915), .A2(n23936), .A3(n23914), .A4(n23913), .ZN(
        n23917) );
  XNOR2_X1 U24015 ( .A(n23917), .B(n23916), .ZN(Ciphertext[174]) );
  OAI211_X1 U24016 ( .C1(n23937), .C2(n23924), .A(n23926), .B(n23918), .ZN(
        n23919) );
  OAI211_X1 U24017 ( .C1(n23924), .C2(n23921), .A(n23920), .B(n23919), .ZN(
        n23923) );
  XNOR2_X1 U24018 ( .A(n23923), .B(n23922), .ZN(Ciphertext[175]) );
  NAND2_X1 U24019 ( .A1(n23937), .A2(n23924), .ZN(n23930) );
  NAND3_X1 U24020 ( .A1(n23934), .A2(n23926), .A3(n23938), .ZN(n23929) );
  NAND2_X1 U24021 ( .A1(n23924), .A2(n23933), .ZN(n23925) );
  OAI21_X1 U24022 ( .B1(n23926), .B2(n23933), .A(n23925), .ZN(n23927) );
  INV_X1 U24025 ( .A(n887), .ZN(n23931) );
  AOI21_X1 U24027 ( .B1(n23934), .B2(n23933), .A(n23939), .ZN(n23935) );
  NAND2_X1 U24028 ( .A1(n23936), .A2(n23935), .ZN(n23944) );
  NAND3_X1 U24029 ( .A1(n24948), .A2(n23938), .A3(n23937), .ZN(n23943) );
  NAND2_X1 U24030 ( .A1(n23941), .A2(n25083), .ZN(n23942) );
  NAND3_X1 U24031 ( .A1(n23944), .A2(n23943), .A3(n23942), .ZN(n23946) );
  XNOR2_X1 U24032 ( .A(n23946), .B(n23945), .ZN(Ciphertext[178]) );
  OAI21_X1 U24033 ( .B1(n23970), .B2(n23966), .A(n23967), .ZN(n23951) );
  OR2_X1 U24034 ( .A1(n23969), .A2(n25017), .ZN(n23948) );
  INV_X1 U24035 ( .A(n23949), .ZN(n23950) );
  NAND2_X1 U24036 ( .A1(n23969), .A2(n23952), .ZN(n23955) );
  OR2_X1 U24037 ( .A1(n23967), .A2(n24910), .ZN(n23963) );
  INV_X1 U24038 ( .A(n23963), .ZN(n23954) );
  XNOR2_X1 U24039 ( .A(n23956), .B(n4023), .ZN(Ciphertext[181]) );
  MUX2_X1 U24040 ( .A(n23966), .B(n24910), .S(n23967), .Z(n23960) );
  MUX2_X1 U24041 ( .A(n23960), .B(n23959), .S(n23969), .Z(n23962) );
  XNOR2_X1 U24042 ( .A(n23962), .B(n23961), .ZN(Ciphertext[182]) );
  INV_X1 U24043 ( .A(n23969), .ZN(n23965) );
  NOR2_X1 U24044 ( .A1(n23967), .A2(n23966), .ZN(n23968) );
  AOI22_X1 U24045 ( .A1(n25076), .A2(n23970), .B1(n23969), .B2(n23968), .ZN(
        n23971) );
  INV_X1 U24046 ( .A(n2044), .ZN(n23973) );
  NAND2_X1 U24047 ( .A1(n23982), .A2(n24012), .ZN(n23974) );
  INV_X1 U24048 ( .A(n24011), .ZN(n23978) );
  NOR2_X1 U24049 ( .A1(n23982), .A2(n24011), .ZN(n23975) );
  AND2_X1 U24050 ( .A1(n24011), .A2(n24012), .ZN(n24015) );
  INV_X1 U24051 ( .A(n1757), .ZN(n23976) );
  XNOR2_X1 U24052 ( .A(n23977), .B(n23976), .ZN(Ciphertext[187]) );
  OR2_X1 U24053 ( .A1(n23978), .A2(n23984), .ZN(n23988) );
  OAI21_X1 U24054 ( .B1(n23979), .B2(n24008), .A(n23988), .ZN(n23992) );
  INV_X1 U24055 ( .A(n24448), .ZN(n24005) );
  NAND3_X1 U24056 ( .A1(n24005), .A2(n24012), .A3(n24954), .ZN(n23980) );
  OAI211_X1 U24057 ( .C1(n24440), .C2(n23981), .A(n23983), .B(n23980), .ZN(
        n23991) );
  NOR3_X1 U24058 ( .A1(n24440), .A2(n24448), .A3(n24954), .ZN(n23985) );
  OAI21_X1 U24059 ( .B1(n24008), .B2(n23987), .A(n23986), .ZN(n23990) );
  OAI211_X1 U24060 ( .C1(n23992), .C2(n23991), .A(n23990), .B(n23989), .ZN(
        Ciphertext[188]) );
  INV_X1 U24061 ( .A(n23993), .ZN(n24014) );
  NAND2_X1 U24062 ( .A1(n24014), .A2(n24954), .ZN(n24018) );
  NOR2_X1 U24063 ( .A1(n22677), .A2(n25439), .ZN(n24003) );
  NAND2_X1 U24064 ( .A1(n23997), .A2(n24003), .ZN(n24001) );
  NAND3_X1 U24065 ( .A1(n22677), .A2(n24439), .A3(n23998), .ZN(n24000) );
  OAI211_X1 U24066 ( .C1(n24003), .C2(n24002), .A(n24001), .B(n24000), .ZN(
        n24004) );
  OAI21_X1 U24067 ( .B1(n24011), .B2(n24004), .A(n24448), .ZN(n24007) );
  INV_X1 U24068 ( .A(n860), .ZN(n24009) );
  NAND2_X1 U24069 ( .A1(n24011), .A2(n24010), .ZN(n24013) );
  NAND2_X1 U24070 ( .A1(n24013), .A2(n24012), .ZN(n24016) );
  AOI22_X1 U24071 ( .A1(n24440), .A2(n24016), .B1(n24015), .B2(n24014), .ZN(
        n24017) );
  OAI21_X1 U24072 ( .B1(n24440), .B2(n24018), .A(n24017), .ZN(n24020) );
  XNOR2_X1 U24073 ( .A(n24020), .B(n3208), .ZN(Ciphertext[191]) );
  XNOR2_X2 U1497 ( .A(n12301), .B(n12300), .ZN(n13123) );
  XNOR2_X2 U515 ( .A(n11273), .B(n11272), .ZN(n13013) );
  MUX2_X2 U2461 ( .A(n9278), .B(n9277), .S(n24511), .Z(n10836) );
  OR2_X1 U120 ( .A1(n11031), .A2(n10772), .ZN(n10779) );
  BUF_X1 U1453 ( .A(n14970), .Z(n16448) );
  MUX2_X2 U2570 ( .A(n6285), .B(n6284), .S(n7801), .Z(n9155) );
  NAND3_X2 U7653 ( .A1(n2433), .A2(n9478), .A3(n9479), .ZN(n12396) );
  XNOR2_X2 U2351 ( .A(n11814), .B(n11815), .ZN(n13234) );
  OAI211_X2 U13628 ( .C1(n7965), .C2(n7966), .A(n7964), .B(n7963), .ZN(n8961)
         );
  BUF_X1 U1505 ( .A(n10632), .Z(n10819) );
  NAND2_X1 U477 ( .A1(n4465), .A2(n4461), .ZN(n11414) );
  NAND4_X2 U1529 ( .A1(n7398), .A2(n7396), .A3(n7397), .A4(n7395), .ZN(n8860)
         );
  NAND3_X2 U1994 ( .A1(n16620), .A2(n2942), .A3(n16623), .ZN(n17476) );
  NAND3_X2 U2623 ( .A1(n4370), .A2(n6951), .A3(n5528), .ZN(n7474) );
  NOR2_X2 U157 ( .A1(n24341), .A2(n23334), .ZN(n22855) );
  OAI211_X1 U4942 ( .C1(n3889), .C2(n13804), .A(n13803), .B(n13802), .ZN(
        n14922) );
  AND4_X2 U81 ( .A1(n10598), .A2(n10597), .A3(n10600), .A4(n10599), .ZN(n11628) );
  OAI211_X2 U1816 ( .C1(n1662), .C2(n19293), .A(n19292), .B(n19291), .ZN(
        n21670) );
  XNOR2_X1 U580 ( .A(n8110), .B(n8111), .ZN(n9943) );
  OAI21_X2 U5199 ( .B1(n4512), .B2(n6937), .A(n4511), .ZN(n3362) );
  AND2_X2 U2013 ( .A1(n2937), .A2(n3068), .ZN(n17663) );
  XNOR2_X2 U1943 ( .A(n17857), .B(n17858), .ZN(n19470) );
  AND3_X2 U55 ( .A1(n13085), .A2(n13084), .A3(n13083), .ZN(n15210) );
  BUF_X1 U1443 ( .A(n15873), .Z(n17087) );
  NOR2_X2 U22814 ( .A1(n23196), .A2(n22752), .ZN(n23200) );
  NAND4_X2 U1525 ( .A1(n6586), .A2(n6584), .A3(n1088), .A4(n6585), .ZN(n8634)
         );
  BUF_X1 U1441 ( .A(n16516), .Z(n17145) );
  NAND4_X2 U1528 ( .A1(n7366), .A2(n7368), .A3(n7367), .A4(n7369), .ZN(n5614)
         );
  NAND4_X2 U1805 ( .A1(n1661), .A2(n1664), .A3(n19739), .A4(n1660), .ZN(n21721) );
  OAI211_X2 U2457 ( .C1(n9570), .C2(n5739), .A(n9569), .B(n9568), .ZN(n10901)
         );
  INV_X1 U1053 ( .A(n396), .ZN(n14077) );
  NOR2_X2 U1823 ( .A1(n20513), .A2(n20512), .ZN(n21307) );
  BUF_X1 U2685 ( .A(n5915), .Z(n6162) );
  INV_X1 U5273 ( .A(n8244), .ZN(n8698) );
  NAND2_X2 U1500 ( .A1(n541), .A2(n10938), .ZN(n12389) );
  BUF_X2 U2698 ( .A(n6071), .Z(n6658) );
  XNOR2_X1 U1176 ( .A(n8344), .B(n8343), .ZN(n10100) );
  NAND2_X2 U2613 ( .A1(n1643), .A2(n3444), .ZN(n7735) );
  OAI21_X2 U1110 ( .B1(n10290), .B2(n10291), .A(n4732), .ZN(n11966) );
  XNOR2_X2 U1462 ( .A(n14504), .B(n14503), .ZN(n15857) );
  XNOR2_X1 U245 ( .A(Key[96]), .B(Plaintext[96]), .ZN(n7032) );
  CLKBUF_X1 U1350 ( .A(Key[146]), .Z(n23620) );
  CLKBUF_X1 U1605 ( .A(Key[4]), .Z(n869) );
  CLKBUF_X1 U2752 ( .A(Key[156]), .Z(n20825) );
  CLKBUF_X1 U102 ( .A(Key[184]), .Z(n92) );
  CLKBUF_X1 U253 ( .A(Key[150]), .Z(n1855) );
  CLKBUF_X1 U1662 ( .A(Key[93]), .Z(n2033) );
  CLKBUF_X1 U2738 ( .A(Key[97]), .Z(n923) );
  CLKBUF_X1 U2742 ( .A(Key[101]), .Z(n20744) );
  CLKBUF_X1 U99 ( .A(Key[168]), .Z(n673) );
  CLKBUF_X1 U100 ( .A(Key[74]), .Z(n2757) );
  XNOR2_X1 U2745 ( .A(Key[144]), .B(Plaintext[144]), .ZN(n6373) );
  CLKBUF_X1 U101 ( .A(Key[29]), .Z(n2747) );
  XNOR2_X1 U12400 ( .A(n5954), .B(Key[172]), .ZN(n6490) );
  CLKBUF_X1 U2692 ( .A(n5916), .Z(n7097) );
  INV_X1 U4560 ( .A(n6651), .ZN(n6894) );
  AND2_X1 U447 ( .A1(n70), .A2(n6943), .ZN(n3050) );
  NAND3_X1 U179 ( .A1(n6031), .A2(n6032), .A3(n6030), .ZN(n7257) );
  AND2_X1 U191 ( .A1(n2800), .A2(n6813), .ZN(n4) );
  OR2_X1 U2642 ( .A1(n2824), .A2(n6258), .ZN(n7798) );
  OAI21_X1 U4853 ( .B1(n7513), .B2(n1690), .A(n7512), .ZN(n9058) );
  NAND3_X1 U698 ( .A1(n6045), .A2(n6044), .A3(n120), .ZN(n9181) );
  INV_X1 U892 ( .A(n8475), .ZN(n9194) );
  XNOR2_X1 U8463 ( .A(n2785), .B(n8670), .ZN(n9664) );
  XNOR2_X1 U3190 ( .A(n9112), .B(n9113), .ZN(n10064) );
  INV_X1 U407 ( .A(n10006), .ZN(n9652) );
  BUF_X1 U321 ( .A(n9550), .Z(n10048) );
  BUF_X1 U826 ( .A(n8744), .Z(n10070) );
  BUF_X1 U2497 ( .A(n9820), .Z(n10141) );
  XNOR2_X1 U2481 ( .A(n8984), .B(n8983), .ZN(n9639) );
  OR2_X1 U788 ( .A1(n2565), .A2(n2585), .ZN(n9378) );
  NOR2_X1 U555 ( .A1(n9323), .A2(n9322), .ZN(n10470) );
  AND2_X1 U4346 ( .A1(n5272), .A2(n5276), .ZN(n5271) );
  AND2_X1 U543 ( .A1(n3863), .A2(n3864), .ZN(n11215) );
  OAI211_X1 U14889 ( .C1(n9643), .C2(n24332), .A(n9642), .B(n9641), .ZN(n11207) );
  NAND2_X1 U1126 ( .A1(n1168), .A2(n9224), .ZN(n11122) );
  INV_X1 U6672 ( .A(n11149), .ZN(n4998) );
  INV_X1 U2425 ( .A(n10800), .ZN(n411) );
  INV_X1 U746 ( .A(n10375), .ZN(n10587) );
  NAND3_X1 U7432 ( .A1(n4211), .A2(n8426), .A3(n4213), .ZN(n11464) );
  AOI22_X1 U1173 ( .A1(n11095), .A2(n11094), .B1(n95), .B2(n11093), .ZN(n11556) );
  CLKBUF_X1 U2360 ( .A(n11776), .Z(n12296) );
  XNOR2_X1 U16560 ( .A(n12265), .B(n12264), .ZN(n12660) );
  XNOR2_X1 U16306 ( .A(n11855), .B(n11854), .ZN(n11873) );
  BUF_X1 U16776 ( .A(n12594), .Z(n13292) );
  XNOR2_X1 U2346 ( .A(n11250), .B(n11249), .ZN(n13216) );
  XNOR2_X1 U662 ( .A(n4931), .B(n11979), .ZN(n111) );
  INV_X1 U405 ( .A(n13291), .ZN(n12910) );
  MUX2_X1 U11267 ( .A(n13064), .B(n13063), .S(n12440), .Z(n5113) );
  AND2_X1 U692 ( .A1(n1316), .A2(n1315), .ZN(n13421) );
  NAND3_X1 U2250 ( .A1(n5544), .A2(n5543), .A3(n12502), .ZN(n13533) );
  AND2_X1 U1136 ( .A1(n1553), .A2(n1554), .ZN(n13892) );
  XNOR2_X1 U232 ( .A(n14960), .B(n15358), .ZN(n15185) );
  XNOR2_X1 U2170 ( .A(n14583), .B(n14582), .ZN(n16096) );
  XNOR2_X1 U2140 ( .A(n13973), .B(n13972), .ZN(n16206) );
  XNOR2_X1 U2162 ( .A(n15007), .B(n15008), .ZN(n16226) );
  INV_X1 U1454 ( .A(n14970), .ZN(n16450) );
  OAI211_X1 U3394 ( .C1(n16424), .C2(n14433), .A(n14432), .B(n14431), .ZN(
        n17229) );
  AND2_X1 U742 ( .A1(n17158), .A2(n17156), .ZN(n16260) );
  AND2_X1 U605 ( .A1(n3424), .A2(n15785), .ZN(n17130) );
  BUF_X1 U19045 ( .A(n16260), .Z(n17163) );
  AND2_X1 U5008 ( .A1(n16375), .A2(n16533), .ZN(n2430) );
  XNOR2_X1 U20506 ( .A(n18545), .B(n18544), .ZN(n19613) );
  MUX2_X1 U972 ( .A(n18811), .B(n18810), .S(n3412), .Z(n20913) );
  INV_X1 U21038 ( .A(n25204), .ZN(n20168) );
  AND3_X1 U968 ( .A1(n1290), .A2(n1288), .A3(n1287), .ZN(n20003) );
  AND2_X1 U785 ( .A1(n1503), .A2(n1504), .ZN(n1327) );
  AOI21_X1 U1884 ( .B1(n19236), .B2(n18869), .A(n18805), .ZN(n20359) );
  INV_X1 U5086 ( .A(n19777), .ZN(n20236) );
  NAND2_X1 U7598 ( .A1(n2198), .A2(n18885), .ZN(n20290) );
  NAND2_X1 U4769 ( .A1(n3962), .A2(n3963), .ZN(n21751) );
  OAI22_X1 U151 ( .A1(n1627), .A2(n5227), .B1(n5226), .B2(n22159), .ZN(n23543)
         );
  OR2_X1 U23461 ( .A1(n22943), .A2(n22942), .ZN(n23349) );
  NOR2_X1 U23762 ( .A1(n23468), .A2(n23467), .ZN(n23472) );
  NOR2_X1 U23160 ( .A1(n23110), .A2(n24498), .ZN(n23093) );
  CLKBUF_X1 U241 ( .A(Key[115]), .Z(n688) );
  INV_X1 U12158 ( .A(n6751), .ZN(n6675) );
  INV_X1 U1607 ( .A(n6871), .ZN(n314) );
  INV_X1 U12148 ( .A(n5800), .ZN(n6965) );
  INV_X1 U2606 ( .A(n8511), .ZN(n7250) );
  AND2_X1 U749 ( .A1(n6160), .A2(n6159), .ZN(n8475) );
  NOR2_X1 U14491 ( .A1(n9064), .A2(n9244), .ZN(n10052) );
  BUF_X1 U1494 ( .A(n11287), .Z(n13246) );
  BUF_X1 U1490 ( .A(n1324), .Z(n13178) );
  NAND2_X2 U1085 ( .A1(n13538), .A2(n13535), .ZN(n14022) );
  INV_X1 U4662 ( .A(n13614), .ZN(n14058) );
  INV_X2 U6155 ( .A(n1516), .ZN(n17629) );
  INV_X1 U1946 ( .A(n4748), .ZN(n19501) );
  NOR2_X1 U11312 ( .A1(n18734), .A2(n19477), .ZN(n18971) );
  INV_X1 U146 ( .A(n22093), .ZN(n22890) );
  INV_X1 U1368 ( .A(n22389), .ZN(n22974) );
  BUF_X1 U1486 ( .A(n11965), .Z(n12695) );
  NAND2_X2 U1185 ( .A1(n7753), .A2(n2623), .ZN(n9057) );
  AOI21_X1 U5577 ( .B1(n16922), .B2(n3783), .A(n3782), .ZN(n17720) );
  NOR2_X2 U10755 ( .A1(n9215), .A2(n9216), .ZN(n4590) );
  AND2_X1 U3 ( .A1(n3035), .A2(n21916), .ZN(n24334) );
  XNOR2_X1 U12 ( .A(n15078), .B(n24303), .ZN(n1122) );
  NAND3_X2 U95 ( .A1(n2512), .A2(n24099), .A3(n5586), .ZN(n20125) );
  BUF_X1 U97 ( .A(n22915), .Z(n23510) );
  INV_X1 U114 ( .A(n15696), .ZN(n16483) );
  XNOR2_X1 U138 ( .A(n13906), .B(n15103), .ZN(n14973) );
  INV_X1 U182 ( .A(n15857), .ZN(n16120) );
  BUF_X2 U229 ( .A(n10135), .Z(n24026) );
  XNOR2_X1 U230 ( .A(n9153), .B(n9152), .ZN(n10135) );
  OAI21_X2 U233 ( .B1(n20602), .B2(n20601), .A(n5363), .ZN(n21734) );
  OAI211_X1 U288 ( .C1(n16074), .C2(n15802), .A(n3639), .B(n3637), .ZN(n17107)
         );
  NAND4_X2 U303 ( .A1(n5488), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n7418)
         );
  AND2_X2 U317 ( .A1(n3977), .A2(n3976), .ZN(n18693) );
  XNOR2_X1 U328 ( .A(Key[158]), .B(Plaintext[158]), .ZN(n6919) );
  BUF_X1 U334 ( .A(n18817), .Z(n19103) );
  AND2_X2 U339 ( .A1(n10004), .A2(n10003), .ZN(n11012) );
  OAI21_X2 U344 ( .B1(n3839), .B2(n6058), .A(n3838), .ZN(n8022) );
  XNOR2_X2 U353 ( .A(n5895), .B(Key[52]), .ZN(n6697) );
  NOR2_X1 U381 ( .A1(n20721), .A2(n20720), .ZN(n23217) );
  OAI211_X2 U396 ( .C1(n9247), .C2(n10054), .A(n9246), .B(n5004), .ZN(n10858)
         );
  XNOR2_X2 U399 ( .A(n19342), .B(n19341), .ZN(n22252) );
  XNOR2_X2 U427 ( .A(n11572), .B(n11573), .ZN(n13041) );
  XNOR2_X2 U430 ( .A(n11480), .B(n11479), .ZN(n12710) );
  XNOR2_X1 U444 ( .A(n11490), .B(n11491), .ZN(n13077) );
  XNOR2_X1 U470 ( .A(n21175), .B(n21174), .ZN(n22593) );
  XNOR2_X2 U497 ( .A(n11539), .B(n11540), .ZN(n12470) );
  AOI22_X2 U507 ( .A1(n12700), .A2(n12699), .B1(n12698), .B2(n25191), .ZN(
        n14190) );
  AND2_X2 U512 ( .A1(n5719), .A2(n5720), .ZN(n7771) );
  OAI211_X2 U522 ( .C1(n22929), .C2(n5768), .A(n1396), .B(n5687), .ZN(n23505)
         );
  OAI21_X2 U567 ( .B1(n19866), .B2(n19865), .A(n19864), .ZN(n20964) );
  OAI211_X1 U581 ( .C1(n6728), .C2(n6727), .A(n6726), .B(n6725), .ZN(n263) );
  XNOR2_X1 U614 ( .A(n5783), .B(Key[93]), .ZN(n6236) );
  NOR2_X1 U632 ( .A1(n12599), .A2(n12598), .ZN(n14851) );
  NAND4_X2 U644 ( .A1(n7275), .A2(n7274), .A3(n7273), .A4(n7272), .ZN(n8875)
         );
  XNOR2_X1 U676 ( .A(n3504), .B(n3505), .ZN(n9898) );
  AND2_X2 U696 ( .A1(n18741), .A2(n18740), .ZN(n20191) );
  XNOR2_X2 U708 ( .A(n3473), .B(n11945), .ZN(n13274) );
  OAI211_X2 U744 ( .C1(n7898), .C2(n7233), .A(n5235), .B(n5236), .ZN(n8612) );
  NOR2_X2 U748 ( .A1(n7921), .A2(n8078), .ZN(n9189) );
  BUF_X2 U750 ( .A(n8901), .Z(n24056) );
  OAI22_X1 U758 ( .A1(n7047), .A2(n7827), .B1(n7513), .B2(n7048), .ZN(n8901)
         );
  OAI21_X2 U775 ( .B1(n20323), .B2(n20322), .A(n20321), .ZN(n24485) );
  NOR2_X1 U825 ( .A1(n22477), .A2(n22476), .ZN(n23119) );
  OAI21_X2 U841 ( .B1(n11120), .B2(n11119), .A(n11118), .ZN(n11715) );
  XNOR2_X1 U846 ( .A(n13606), .B(n14633), .ZN(n16405) );
  BUF_X1 U852 ( .A(n23742), .Z(n24064) );
  BUF_X1 U854 ( .A(n23742), .Z(n24065) );
  BUF_X1 U888 ( .A(n6534), .Z(n24067) );
  XNOR2_X1 U909 ( .A(n5865), .B(Key[26]), .ZN(n6534) );
  XNOR2_X2 U910 ( .A(Key[9]), .B(Plaintext[9]), .ZN(n6498) );
  NAND3_X2 U958 ( .A1(n10857), .A2(n3502), .A3(n24251), .ZN(n12391) );
  OAI211_X2 U987 ( .C1(n11156), .C2(n11155), .A(n11154), .B(n11153), .ZN(
        n11977) );
  OAI21_X2 U1009 ( .B1(n6443), .B2(n6442), .A(n6441), .ZN(n2404) );
  AOI22_X1 U1035 ( .A1(n6390), .A2(n6391), .B1(n6388), .B2(n6389), .ZN(n7850)
         );
  XNOR2_X2 U1050 ( .A(n16600), .B(n16601), .ZN(n19560) );
  NAND4_X2 U1074 ( .A1(n4404), .A2(n4403), .A3(n4402), .A4(n18850), .ZN(n20068) );
  OAI211_X2 U1117 ( .C1(n7776), .C2(n7775), .A(n7773), .B(n7774), .ZN(n9106)
         );
  NOR2_X2 U1156 ( .A1(n13675), .A2(n13669), .ZN(n14003) );
  AOI22_X2 U1170 ( .A1(n6085), .A2(n6767), .B1(n6084), .B2(n314), .ZN(n7757)
         );
  XNOR2_X2 U1174 ( .A(n20656), .B(n20655), .ZN(n22977) );
  NOR2_X2 U1177 ( .A1(n10324), .A2(n10323), .ZN(n12189) );
  BUF_X1 U1200 ( .A(n9450), .Z(n24511) );
  OR2_X1 U1202 ( .A1(n6277), .A2(n440), .ZN(n24277) );
  CLKBUF_X1 U1205 ( .A(Key[82]), .Z(n24287) );
  INV_X1 U1225 ( .A(n23411), .ZN(n24074) );
  AND2_X1 U1237 ( .A1(n4947), .A2(n4949), .ZN(n24351) );
  AND3_X1 U1241 ( .A1(n3087), .A2(n4102), .A3(n4099), .ZN(n23220) );
  INV_X1 U1250 ( .A(n23077), .ZN(n24075) );
  AND3_X1 U1251 ( .A1(n24242), .A2(n747), .A3(n3939), .ZN(n23125) );
  OR2_X1 U1252 ( .A1(n21827), .A2(n3890), .ZN(n24307) );
  OR3_X1 U1257 ( .A1(n22212), .A2(n22211), .A3(n22210), .ZN(n22213) );
  AND2_X1 U1259 ( .A1(n24115), .A2(n24113), .ZN(n22046) );
  OAI211_X1 U1276 ( .C1(n20564), .C2(n25221), .A(n4009), .B(n19734), .ZN(
        n24491) );
  NOR2_X1 U1285 ( .A1(n20078), .A2(n20077), .ZN(n20912) );
  OR2_X1 U1294 ( .A1(n19988), .A2(n24315), .ZN(n24154) );
  INV_X1 U1295 ( .A(n20381), .ZN(n24128) );
  AOI21_X1 U1302 ( .B1(n20232), .B2(n25205), .A(n20231), .ZN(n20240) );
  INV_X1 U1309 ( .A(n20615), .ZN(n24076) );
  INV_X1 U1311 ( .A(n20360), .ZN(n24078) );
  BUF_X1 U1312 ( .A(n20618), .Z(n24338) );
  AND3_X1 U1315 ( .A1(n19447), .A2(n19448), .A3(n24136), .ZN(n20169) );
  INV_X1 U1325 ( .A(n3989), .ZN(n19036) );
  XNOR2_X1 U1333 ( .A(n18566), .B(n18565), .ZN(n19417) );
  INV_X1 U1362 ( .A(n19071), .ZN(n24079) );
  XNOR2_X1 U1379 ( .A(n18249), .B(n18250), .ZN(n19546) );
  INV_X1 U1384 ( .A(n372), .ZN(n16775) );
  INV_X1 U1395 ( .A(n17014), .ZN(n367) );
  OR2_X1 U1422 ( .A1(n5024), .A2(n14839), .ZN(n24149) );
  INV_X1 U1445 ( .A(n1122), .ZN(n16286) );
  OR2_X1 U1446 ( .A1(n15549), .A2(n25446), .ZN(n16068) );
  INV_X1 U1452 ( .A(n16352), .ZN(n24080) );
  AND2_X1 U1516 ( .A1(n1203), .A2(n1204), .ZN(n24259) );
  NAND2_X1 U1517 ( .A1(n2774), .A2(n12544), .ZN(n15169) );
  NOR2_X1 U1537 ( .A1(n24503), .A2(n14099), .ZN(n24181) );
  INV_X1 U1538 ( .A(n177), .ZN(n14083) );
  AND2_X1 U1539 ( .A1(n13969), .A2(n13966), .ZN(n13599) );
  AND2_X1 U1542 ( .A1(n14065), .A2(n14064), .ZN(n24135) );
  OR2_X1 U1609 ( .A1(n13854), .A2(n13853), .ZN(n177) );
  AOI21_X1 U1690 ( .B1(n3935), .B2(n12653), .A(n12724), .ZN(n13670) );
  AND2_X1 U1693 ( .A1(n13056), .A2(n12795), .ZN(n12526) );
  INV_X1 U1695 ( .A(n11993), .ZN(n24241) );
  XNOR2_X1 U1704 ( .A(n11313), .B(n11312), .ZN(n12995) );
  INV_X1 U1710 ( .A(n11263), .ZN(n12225) );
  INV_X1 U1771 ( .A(n11149), .ZN(n24286) );
  INV_X1 U1811 ( .A(n11209), .ZN(n24082) );
  AND2_X1 U1821 ( .A1(n11130), .A2(n10714), .ZN(n24164) );
  NOR2_X1 U1852 ( .A1(n9467), .A2(n9466), .ZN(n24345) );
  OR2_X1 U1890 ( .A1(n24534), .A2(n9991), .ZN(n9659) );
  INV_X1 U1911 ( .A(n9898), .ZN(n24083) );
  INV_X1 U1915 ( .A(n9934), .ZN(n24084) );
  XNOR2_X1 U1916 ( .A(n6222), .B(n6221), .ZN(n9461) );
  INV_X1 U1917 ( .A(n9842), .ZN(n24085) );
  INV_X1 U1933 ( .A(n10147), .ZN(n24087) );
  OR2_X1 U1968 ( .A1(n7721), .A2(n24072), .ZN(n7727) );
  OR2_X1 U2069 ( .A1(n6923), .A2(n1175), .ZN(n24147) );
  OR2_X1 U2081 ( .A1(n6940), .A2(n5908), .ZN(n6943) );
  INV_X1 U2085 ( .A(n6969), .ZN(n24089) );
  OR2_X1 U2086 ( .A1(n6390), .A2(n6976), .ZN(n24262) );
  BUF_X1 U2088 ( .A(n5795), .Z(n6619) );
  OR2_X1 U2128 ( .A1(n6373), .A2(n5824), .ZN(n24177) );
  INV_X1 U2134 ( .A(n6112), .ZN(n24125) );
  BUF_X1 U2139 ( .A(n6368), .Z(n6997) );
  AND2_X1 U2211 ( .A1(n6123), .A2(n6838), .ZN(n24255) );
  INV_X1 U2316 ( .A(n7762), .ZN(n7648) );
  OR2_X1 U2334 ( .A1(n7899), .A2(n24103), .ZN(n2758) );
  BUF_X1 U2338 ( .A(n7294), .Z(n8015) );
  OR2_X1 U2341 ( .A1(n7765), .A2(n7648), .ZN(n24119) );
  XNOR2_X1 U2350 ( .A(n8333), .B(n8069), .ZN(n8865) );
  CLKBUF_X1 U2376 ( .A(n9496), .Z(n10089) );
  INV_X1 U2388 ( .A(n11302), .ZN(n95) );
  AND2_X1 U2417 ( .A1(n24345), .A2(n10887), .ZN(n24141) );
  OAI211_X1 U2437 ( .C1(n8804), .C2(n9973), .A(n8803), .B(n24225), .ZN(n11518)
         );
  OAI21_X1 U2460 ( .B1(n1871), .B2(n9691), .A(n9690), .ZN(n1357) );
  INV_X1 U2473 ( .A(n9367), .ZN(n9825) );
  CLKBUF_X1 U2478 ( .A(n10533), .Z(n11145) );
  OR2_X1 U2510 ( .A1(n10767), .A2(n10889), .ZN(n4654) );
  MUX2_X1 U2539 ( .A(n10228), .B(n10227), .S(n10789), .Z(n10231) );
  OR2_X1 U2587 ( .A1(n13234), .A2(n12935), .ZN(n148) );
  NOR2_X1 U2604 ( .A1(n13014), .A2(n13013), .ZN(n13248) );
  OR2_X1 U2656 ( .A1(n14190), .A2(n24347), .ZN(n24186) );
  XNOR2_X1 U2660 ( .A(n11994), .B(n24241), .ZN(n24443) );
  AND2_X1 U2686 ( .A1(n4925), .A2(n4924), .ZN(n5472) );
  AND2_X1 U2695 ( .A1(n14252), .A2(n14251), .ZN(n24301) );
  XNOR2_X1 U2719 ( .A(n3862), .B(n3861), .ZN(n24487) );
  OAI211_X1 U2778 ( .C1(n12532), .C2(n12531), .A(n3315), .B(n3314), .ZN(n14269) );
  OR2_X1 U2788 ( .A1(n13563), .A2(n13564), .ZN(n24121) );
  OR2_X1 U2809 ( .A1(n13773), .A2(n13774), .ZN(n82) );
  NAND3_X1 U2821 ( .A1(n598), .A2(n4907), .A3(n597), .ZN(n14311) );
  OR2_X1 U2826 ( .A1(n13436), .A2(n14106), .ZN(n24519) );
  AOI21_X1 U2841 ( .B1(n13849), .B2(n13848), .A(n24135), .ZN(n14611) );
  NAND2_X1 U2855 ( .A1(n13816), .A2(n13817), .ZN(n15094) );
  XNOR2_X1 U2866 ( .A(n15095), .B(n15098), .ZN(n12) );
  OAI211_X1 U2875 ( .C1(n12703), .C2(n13785), .A(n12702), .B(n12701), .ZN(
        n15358) );
  INV_X1 U2876 ( .A(n1867), .ZN(n15321) );
  AND2_X1 U2886 ( .A1(n24170), .A2(n1261), .ZN(n24169) );
  OAI21_X1 U2932 ( .B1(n24249), .B2(n15625), .A(n24248), .ZN(n15627) );
  OR2_X1 U2933 ( .A1(n16064), .A2(n16060), .ZN(n24227) );
  BUF_X1 U2950 ( .A(n4897), .Z(n16508) );
  OR2_X1 U2958 ( .A1(n17161), .A2(n17162), .ZN(n24250) );
  AND2_X2 U3017 ( .A1(n995), .A2(n646), .ZN(n17335) );
  OAI21_X1 U3021 ( .B1(n2233), .B2(n2234), .A(n5406), .ZN(n4743) );
  AND2_X1 U3023 ( .A1(n17357), .A2(n16877), .ZN(n118) );
  BUF_X1 U3033 ( .A(n18832), .Z(n24478) );
  XNOR2_X1 U3044 ( .A(n39), .B(n16037), .ZN(n17814) );
  CLKBUF_X1 U3045 ( .A(n19370), .Z(n24361) );
  OR2_X1 U3090 ( .A1(n19451), .A2(n19452), .ZN(n24137) );
  AOI21_X1 U3107 ( .B1(n4436), .B2(n18917), .A(n19146), .ZN(n19148) );
  OR2_X1 U3114 ( .A1(n19522), .A2(n19523), .ZN(n24252) );
  INV_X1 U3119 ( .A(n19031), .ZN(n19029) );
  OR2_X1 U3125 ( .A1(n1506), .A2(n19210), .ZN(n160) );
  AOI22_X1 U3129 ( .A1(n1307), .A2(n1306), .B1(n19423), .B2(n19167), .ZN(n1305) );
  NOR2_X1 U3167 ( .A1(n24078), .A2(n20913), .ZN(n20482) );
  OR2_X1 U3191 ( .A1(n20514), .A2(n20517), .ZN(n22) );
  NOR2_X1 U3202 ( .A1(n4287), .A2(n18938), .ZN(n18940) );
  BUF_X1 U3218 ( .A(n20346), .Z(n24414) );
  AOI22_X1 U3223 ( .A1(n20569), .A2(n20617), .B1(n20614), .B2(n20618), .ZN(
        n20327) );
  OR2_X1 U3227 ( .A1(n20452), .A2(n20960), .ZN(n24189) );
  INV_X1 U3231 ( .A(n20022), .ZN(n20567) );
  AND2_X1 U3234 ( .A1(n20341), .A2(n19709), .ZN(n20665) );
  INV_X1 U3237 ( .A(n22361), .ZN(n24114) );
  OR2_X1 U3246 ( .A1(n22792), .A2(n2397), .ZN(n4080) );
  OR2_X1 U3248 ( .A1(n22946), .A2(n2674), .ZN(n2673) );
  OR2_X1 U3260 ( .A1(n24877), .A2(n23014), .ZN(n23463) );
  OR2_X1 U3299 ( .A1(n2987), .A2(n21825), .ZN(n580) );
  OR2_X1 U3304 ( .A1(n22578), .A2(n24075), .ZN(n24278) );
  CLKBUF_X1 U3327 ( .A(Key[183]), .Z(n2745) );
  OAI211_X1 U3344 ( .C1(n22959), .C2(n1259), .A(n1258), .B(n1257), .ZN(n23379)
         );
  OR2_X1 U3347 ( .A1(n23544), .A2(n23537), .ZN(n23549) );
  CLKBUF_X1 U3354 ( .A(Key[185]), .Z(n22702) );
  XNOR2_X1 U3359 ( .A(Key[25]), .B(Plaintext[25]), .ZN(n6533) );
  AND2_X1 U3365 ( .A1(n6827), .A2(n6598), .ZN(n24090) );
  INV_X1 U3371 ( .A(n20578), .ZN(n24194) );
  INV_X1 U3373 ( .A(n3926), .ZN(n24257) );
  AND2_X1 U3410 ( .A1(n6959), .A2(n6703), .ZN(n24091) );
  INV_X1 U3418 ( .A(n3469), .ZN(n24103) );
  XOR2_X1 U3422 ( .A(n9056), .B(n9055), .Z(n24092) );
  INV_X1 U3425 ( .A(n10406), .ZN(n24118) );
  NAND3_X1 U3426 ( .A1(n9346), .A2(n9600), .A3(n9599), .ZN(n24093) );
  OR2_X1 U3427 ( .A1(n13045), .A2(n13038), .ZN(n24094) );
  INV_X1 U3431 ( .A(n12935), .ZN(n24220) );
  AND2_X1 U3449 ( .A1(n1969), .A2(n1967), .ZN(n24095) );
  OR2_X1 U3460 ( .A1(n13235), .A2(n13234), .ZN(n24096) );
  AND2_X1 U3465 ( .A1(n14419), .A2(n2863), .ZN(n24097) );
  INV_X1 U3468 ( .A(n16247), .ZN(n24162) );
  XNOR2_X1 U3485 ( .A(n14576), .B(n14577), .ZN(n16147) );
  INV_X1 U3512 ( .A(n16147), .ZN(n24249) );
  XOR2_X1 U3527 ( .A(n14624), .B(n14623), .Z(n24098) );
  INV_X1 U3551 ( .A(n19456), .ZN(n24172) );
  XNOR2_X1 U3587 ( .A(n17871), .B(n17870), .ZN(n17872) );
  INV_X1 U3594 ( .A(n20491), .ZN(n24275) );
  AND3_X1 U3600 ( .A1(n87), .A2(n3032), .A3(n3794), .ZN(n24100) );
  OR2_X1 U3603 ( .A1(n20960), .A2(n24354), .ZN(n24101) );
  NAND2_X1 U3612 ( .A1(n7232), .A2(n7230), .ZN(n7899) );
  OAI211_X1 U3615 ( .C1(n421), .C2(n9836), .A(n4302), .B(n10098), .ZN(n24104)
         );
  NAND2_X1 U3673 ( .A1(n356), .A2(n18927), .ZN(n18928) );
  OAI22_X1 U3688 ( .A1(n16069), .A2(n15694), .B1(n16068), .B2(n16067), .ZN(
        n16070) );
  NAND2_X1 U3697 ( .A1(n16063), .A2(n16062), .ZN(n16069) );
  NAND3_X2 U3726 ( .A1(n2981), .A2(n24107), .A3(n24106), .ZN(n23554) );
  NAND2_X1 U3727 ( .A1(n22096), .A2(n22890), .ZN(n24106) );
  NAND2_X1 U3738 ( .A1(n22097), .A2(n22729), .ZN(n24107) );
  NAND2_X1 U3739 ( .A1(n5291), .A2(n7054), .ZN(n5294) );
  XNOR2_X1 U3795 ( .A(n15422), .B(n24108), .ZN(n12451) );
  XNOR2_X1 U3834 ( .A(n14892), .B(n3158), .ZN(n24108) );
  NAND3_X1 U3853 ( .A1(n20567), .A2(n20094), .A3(n20560), .ZN(n24109) );
  OAI21_X1 U3890 ( .B1(n19213), .B2(n25392), .A(n24110), .ZN(n3811) );
  NAND3_X1 U3894 ( .A1(n1212), .A2(n24312), .A3(n19361), .ZN(n24110) );
  NAND2_X1 U3928 ( .A1(n16133), .A2(n16074), .ZN(n17159) );
  NAND2_X1 U3966 ( .A1(n19446), .A2(n18990), .ZN(n3989) );
  NAND2_X1 U3967 ( .A1(n13628), .A2(n177), .ZN(n176) );
  OR2_X1 U4003 ( .A1(n16186), .A2(n15970), .ZN(n13941) );
  XNOR2_X1 U4062 ( .A(n24112), .B(n455), .ZN(Ciphertext[4]) );
  NAND2_X1 U4084 ( .A1(n1925), .A2(n1926), .ZN(n6614) );
  NAND2_X1 U4106 ( .A1(n245), .A2(n24114), .ZN(n24113) );
  AOI21_X1 U4108 ( .B1(n22361), .B2(n22356), .A(n21839), .ZN(n24115) );
  INV_X1 U4125 ( .A(n4520), .ZN(n10926) );
  NAND2_X1 U4146 ( .A1(n10994), .A2(n10993), .ZN(n4520) );
  NOR2_X1 U4168 ( .A1(n17451), .A2(n523), .ZN(n17456) );
  NOR2_X2 U4169 ( .A1(n1900), .A2(n5335), .ZN(n12404) );
  OR2_X1 U4187 ( .A1(n9387), .A2(n9959), .ZN(n2875) );
  NAND3_X1 U4191 ( .A1(n4936), .A2(n10730), .A3(n10480), .ZN(n2831) );
  NAND3_X1 U4192 ( .A1(n16756), .A2(n16957), .A3(n17414), .ZN(n16758) );
  NAND3_X2 U4198 ( .A1(n24119), .A2(n24120), .A3(n7308), .ZN(n8799) );
  NAND2_X1 U4201 ( .A1(n2848), .A2(n7306), .ZN(n24120) );
  XNOR2_X1 U4205 ( .A(n5215), .B(n15174), .ZN(n14494) );
  AOI22_X2 U4207 ( .A1(n178), .A2(n14203), .B1(n14202), .B2(n14944), .ZN(
        n15174) );
  NAND3_X1 U4242 ( .A1(n4774), .A2(n16532), .A3(n17164), .ZN(n16265) );
  AOI22_X1 U4257 ( .A1(n16052), .A2(n16051), .B1(n16053), .B2(n16508), .ZN(
        n16054) );
  BUF_X1 U4267 ( .A(n14100), .Z(n24375) );
  BUF_X1 U4283 ( .A(n23479), .Z(n24336) );
  NAND2_X1 U4286 ( .A1(n13562), .A2(n24121), .ZN(n14667) );
  NAND3_X1 U4301 ( .A1(n23896), .A2(n23906), .A3(n23903), .ZN(n23872) );
  NAND3_X1 U4318 ( .A1(n24124), .A2(n24123), .A3(n6608), .ZN(n7767) );
  NAND3_X1 U4338 ( .A1(n6110), .A2(n6606), .A3(n6611), .ZN(n24123) );
  NAND2_X1 U4413 ( .A1(n24125), .A2(n6610), .ZN(n24124) );
  NAND3_X1 U4502 ( .A1(n14271), .A2(n14274), .A3(n13840), .ZN(n13622) );
  OR2_X1 U4525 ( .A1(n16243), .A2(n15707), .ZN(n16241) );
  AND2_X1 U4545 ( .A1(n648), .A2(n16064), .ZN(n24233) );
  NAND3_X1 U4551 ( .A1(n24326), .A2(n19395), .A3(n19393), .ZN(n1458) );
  NAND3_X1 U4641 ( .A1(n20507), .A2(n20216), .A3(n25223), .ZN(n1808) );
  AND2_X1 U4747 ( .A1(n7985), .A2(n7984), .ZN(n24197) );
  NAND2_X1 U4824 ( .A1(n24101), .A2(n24128), .ZN(n24127) );
  NAND3_X1 U4878 ( .A1(n17441), .A2(n17442), .A3(n2549), .ZN(n139) );
  XNOR2_X1 U4884 ( .A(n24131), .B(n24130), .ZN(Ciphertext[131]) );
  INV_X1 U4898 ( .A(n2228), .ZN(n24130) );
  NAND2_X1 U4926 ( .A1(n24133), .A2(n24132), .ZN(n24131) );
  NAND2_X1 U4953 ( .A1(n22748), .A2(n22749), .ZN(n24132) );
  NAND2_X1 U5025 ( .A1(n22750), .A2(n25405), .ZN(n24133) );
  NAND2_X1 U5087 ( .A1(n8023), .A2(n7531), .ZN(n4708) );
  OAI21_X2 U5092 ( .B1(n14072), .B2(n24134), .A(n14070), .ZN(n15497) );
  NAND2_X1 U5115 ( .A1(n14066), .A2(n14264), .ZN(n24134) );
  NAND3_X1 U5130 ( .A1(n4106), .A2(n4053), .A3(n6925), .ZN(n3311) );
  NAND2_X1 U5178 ( .A1(n7514), .A2(n7973), .ZN(n2177) );
  NAND3_X1 U5196 ( .A1(n9133), .A2(n9132), .A3(n9951), .ZN(n1092) );
  NAND2_X1 U5205 ( .A1(n9947), .A2(n9389), .ZN(n9133) );
  NAND3_X1 U5213 ( .A1(n1879), .A2(n7854), .A3(n1880), .ZN(n6419) );
  OR2_X1 U5344 ( .A1(n20449), .A2(n20450), .ZN(n24188) );
  NAND2_X1 U5390 ( .A1(n16177), .A2(n15657), .ZN(n15992) );
  NAND3_X1 U5399 ( .A1(n19449), .A2(n25002), .A3(n24137), .ZN(n24136) );
  NAND2_X1 U5404 ( .A1(n19018), .A2(n20537), .ZN(n19688) );
  NAND3_X1 U5441 ( .A1(n2386), .A2(n10212), .A3(n10886), .ZN(n10214) );
  NAND3_X2 U5470 ( .A1(n1735), .A2(n1734), .A3(n6402), .ZN(n7721) );
  NAND2_X1 U5499 ( .A1(n19918), .A2(n19917), .ZN(n24138) );
  OR2_X1 U5579 ( .A1(n17087), .A2(n16578), .ZN(n2813) );
  NAND2_X1 U5605 ( .A1(n424), .A2(n24139), .ZN(n8572) );
  AND2_X1 U5609 ( .A1(n8571), .A2(n9782), .ZN(n24139) );
  OAI21_X1 U5614 ( .B1(n10544), .B2(n2389), .A(n24140), .ZN(n10545) );
  NAND2_X1 U5635 ( .A1(n2386), .A2(n24141), .ZN(n24140) );
  OAI211_X2 U5722 ( .C1(n16782), .C2(n16859), .A(n24143), .B(n3002), .ZN(
        n18103) );
  NAND2_X1 U5734 ( .A1(n16779), .A2(n16780), .ZN(n24143) );
  OAI211_X1 U5757 ( .C1(n9600), .C2(n24084), .A(n9205), .B(n25217), .ZN(n24144) );
  NAND3_X1 U5878 ( .A1(n391), .A2(n14291), .A3(n13909), .ZN(n24146) );
  NAND3_X1 U5890 ( .A1(n6199), .A2(n6922), .A3(n24147), .ZN(n7294) );
  NAND2_X1 U5956 ( .A1(n9626), .A2(n10046), .ZN(n24148) );
  NAND2_X2 U5970 ( .A1(n5023), .A2(n24149), .ZN(n17607) );
  NAND2_X1 U6031 ( .A1(n24153), .A2(n24150), .ZN(n13457) );
  NAND2_X1 U6134 ( .A1(n24152), .A2(n24151), .ZN(n24150) );
  NOR2_X1 U6136 ( .A1(n13947), .A2(n14306), .ZN(n24151) );
  INV_X1 U6196 ( .A(n13892), .ZN(n24152) );
  NAND2_X1 U6281 ( .A1(n12838), .A2(n12839), .ZN(n3010) );
  NAND3_X1 U6372 ( .A1(n19446), .A2(n19444), .A3(n19445), .ZN(n19447) );
  NAND2_X1 U6404 ( .A1(n883), .A2(n884), .ZN(n24155) );
  INV_X1 U6486 ( .A(n7114), .ZN(n5318) );
  NAND2_X1 U6502 ( .A1(n7762), .A2(n7647), .ZN(n7114) );
  NAND2_X1 U6544 ( .A1(n23875), .A2(n24158), .ZN(n23878) );
  OR2_X1 U6545 ( .A1(n23904), .A2(n23883), .ZN(n24158) );
  NAND2_X1 U6556 ( .A1(n24159), .A2(n19465), .ZN(n17890) );
  NAND2_X1 U6569 ( .A1(n19032), .A2(n19460), .ZN(n24159) );
  AOI22_X1 U6575 ( .A1(n19814), .A2(n20507), .B1(n20510), .B2(n20218), .ZN(
        n19815) );
  OAI21_X1 U6584 ( .B1(n22184), .B2(n1336), .A(n24160), .ZN(n2296) );
  NAND2_X1 U6659 ( .A1(n1336), .A2(n22239), .ZN(n24160) );
  NAND2_X1 U6706 ( .A1(n24161), .A2(n9575), .ZN(n11845) );
  NAND3_X1 U6711 ( .A1(n24167), .A2(n24166), .A3(n2388), .ZN(n24161) );
  INV_X1 U6728 ( .A(n16252), .ZN(n24163) );
  NAND2_X1 U6750 ( .A1(n10840), .A2(n24164), .ZN(n10717) );
  AND2_X2 U6787 ( .A1(n788), .A2(n2282), .ZN(n18388) );
  NAND3_X1 U6818 ( .A1(n17366), .A2(n17363), .A3(n17364), .ZN(n2452) );
  INV_X1 U6907 ( .A(n24383), .ZN(n17755) );
  NAND3_X1 U6914 ( .A1(n2790), .A2(n16259), .A3(n2789), .ZN(n24383) );
  NAND2_X1 U6915 ( .A1(n10884), .A2(n10302), .ZN(n24166) );
  INV_X1 U6930 ( .A(n10884), .ZN(n24168) );
  NAND2_X1 U6943 ( .A1(n2008), .A2(n5907), .ZN(n2007) );
  NAND2_X1 U7002 ( .A1(n16122), .A2(n16155), .ZN(n16158) );
  NAND2_X1 U7012 ( .A1(n9368), .A2(n9398), .ZN(n9367) );
  INV_X1 U7037 ( .A(n17277), .ZN(n24300) );
  INV_X1 U7076 ( .A(n15611), .ZN(n24170) );
  AOI21_X2 U7134 ( .B1(n13442), .B2(n13443), .A(n755), .ZN(n15505) );
  INV_X1 U7167 ( .A(n523), .ZN(n17460) );
  NAND2_X1 U7170 ( .A1(n3451), .A2(n16359), .ZN(n16361) );
  NAND2_X1 U7255 ( .A1(n24597), .A2(n7312), .ZN(n24198) );
  NAND2_X1 U7260 ( .A1(n7582), .A2(n7584), .ZN(n7312) );
  OR2_X1 U7263 ( .A1(n17463), .A2(n16846), .ZN(n17465) );
  NAND2_X1 U7268 ( .A1(n24243), .A2(n24244), .ZN(n18975) );
  NAND2_X1 U7293 ( .A1(n508), .A2(n13953), .ZN(n14159) );
  NAND2_X1 U7303 ( .A1(n11216), .A2(n10623), .ZN(n10620) );
  NAND2_X1 U7368 ( .A1(n24178), .A2(n24177), .ZN(n6790) );
  NAND2_X1 U7380 ( .A1(n6374), .A2(n6375), .ZN(n24178) );
  XNOR2_X1 U7513 ( .A(n24179), .B(n18050), .ZN(n18052) );
  XNOR2_X1 U7515 ( .A(n18567), .B(n17663), .ZN(n24179) );
  NAND2_X1 U7524 ( .A1(n14097), .A2(n24180), .ZN(n14103) );
  NAND2_X1 U7553 ( .A1(n24182), .A2(n24181), .ZN(n24180) );
  INV_X1 U7567 ( .A(n4894), .ZN(n24182) );
  NAND2_X1 U7585 ( .A1(n2909), .A2(n2907), .ZN(n24183) );
  NAND2_X1 U7597 ( .A1(n16619), .A2(n16620), .ZN(n16552) );
  OAI21_X1 U7601 ( .B1(n15694), .B2(n25446), .A(n16060), .ZN(n648) );
  NAND2_X1 U7646 ( .A1(n3456), .A2(n22221), .ZN(n24184) );
  NAND2_X1 U7692 ( .A1(n15562), .A2(n24506), .ZN(n24185) );
  NAND2_X1 U7694 ( .A1(n19752), .A2(n19987), .ZN(n21067) );
  NAND2_X1 U7731 ( .A1(n16344), .A2(n24187), .ZN(n16346) );
  NAND2_X1 U7816 ( .A1(n16341), .A2(n16342), .ZN(n24187) );
  AOI22_X2 U7853 ( .A1(n10204), .A2(n10451), .B1(n9375), .B2(n4505), .ZN(
        n12249) );
  NAND3_X1 U7868 ( .A1(n2082), .A2(n7826), .A3(n2081), .ZN(n2080) );
  NAND2_X1 U7882 ( .A1(n249), .A2(n6848), .ZN(n7028) );
  NAND2_X1 U7897 ( .A1(n24191), .A2(n24190), .ZN(n18964) );
  NAND2_X1 U7899 ( .A1(n18957), .A2(n19471), .ZN(n24190) );
  NAND2_X1 U7936 ( .A1(n18958), .A2(n18945), .ZN(n24191) );
  XNOR2_X1 U7965 ( .A(n24192), .B(n18239), .ZN(n18493) );
  NAND2_X1 U7967 ( .A1(n12960), .A2(n13339), .ZN(n12577) );
  OAI21_X1 U8020 ( .B1(n20194), .B2(n24194), .A(n24193), .ZN(n20582) );
  NAND2_X1 U8022 ( .A1(n20194), .A2(n20576), .ZN(n24193) );
  NAND3_X1 U8063 ( .A1(n690), .A2(n14101), .A3(n689), .ZN(n672) );
  NAND2_X1 U8142 ( .A1(n5464), .A2(n2090), .ZN(n24195) );
  NAND3_X1 U8143 ( .A1(n17287), .A2(n17289), .A3(n17288), .ZN(n24196) );
  NAND2_X1 U8159 ( .A1(n7826), .A2(n24197), .ZN(n7831) );
  NAND3_X1 U8223 ( .A1(n7018), .A2(n24200), .A3(n24199), .ZN(n7965) );
  NAND3_X1 U8237 ( .A1(n7015), .A2(n7016), .A3(n7014), .ZN(n24199) );
  NAND2_X1 U8239 ( .A1(n24090), .A2(n6824), .ZN(n24200) );
  OAI211_X1 U8241 ( .C1(n15535), .C2(n16038), .A(n1718), .B(n24098), .ZN(
        n17158) );
  NAND2_X1 U8257 ( .A1(n9435), .A2(n9634), .ZN(n10038) );
  NAND2_X1 U8275 ( .A1(n24202), .A2(n16708), .ZN(n16374) );
  NAND2_X1 U8276 ( .A1(n16372), .A2(n16616), .ZN(n24202) );
  NAND2_X1 U8281 ( .A1(n16170), .A2(n16426), .ZN(n706) );
  INV_X1 U8298 ( .A(n7926), .ZN(n24203) );
  NAND2_X1 U8309 ( .A1(n6555), .A2(n6554), .ZN(n7926) );
  NOR2_X1 U8336 ( .A1(n24012), .A2(n24011), .ZN(n24204) );
  OAI21_X1 U8387 ( .B1(n7607), .B2(n7608), .A(n7606), .ZN(n24205) );
  NOR2_X1 U8472 ( .A1(n4541), .A2(n24352), .ZN(n15541) );
  NAND2_X1 U8488 ( .A1(n20125), .A2(n20547), .ZN(n5638) );
  NAND2_X1 U8505 ( .A1(n266), .A2(n4004), .ZN(n16316) );
  XNOR2_X1 U8522 ( .A(n20792), .B(n21713), .ZN(n19955) );
  OAI22_X1 U8548 ( .A1(n11086), .A2(n11085), .B1(n11084), .B2(n418), .ZN(n1263) );
  NAND2_X1 U8559 ( .A1(n5559), .A2(n10890), .ZN(n11086) );
  OAI211_X1 U8568 ( .C1(n9340), .C2(n10156), .A(n3988), .B(n10154), .ZN(n10336) );
  OAI211_X1 U8587 ( .C1(n1251), .C2(n19460), .A(n24209), .B(n19465), .ZN(
        n18741) );
  NAND2_X1 U8598 ( .A1(n1251), .A2(n18979), .ZN(n24209) );
  NAND3_X1 U8617 ( .A1(n19470), .A2(n18959), .A3(n18960), .ZN(n5099) );
  XNOR2_X1 U8619 ( .A(n21572), .B(n21135), .ZN(n21463) );
  AND2_X2 U8625 ( .A1(n24211), .A2(n24210), .ZN(n21135) );
  NAND2_X1 U8636 ( .A1(n18743), .A2(n20183), .ZN(n24210) );
  NAND2_X1 U8643 ( .A1(n18742), .A2(n19862), .ZN(n24211) );
  OR2_X1 U8647 ( .A1(n10148), .A2(n25207), .ZN(n9522) );
  NAND3_X1 U8651 ( .A1(n9746), .A2(n24535), .A3(n25121), .ZN(n24212) );
  AND3_X2 U8652 ( .A1(n24214), .A2(n3728), .A3(n24213), .ZN(n11914) );
  INV_X1 U8671 ( .A(n8032), .ZN(n24214) );
  NAND3_X1 U8703 ( .A1(n10292), .A2(n10840), .A3(n10293), .ZN(n10294) );
  NAND2_X1 U8771 ( .A1(n11098), .A2(n11097), .ZN(n24215) );
  NAND2_X1 U8772 ( .A1(n102), .A2(n9490), .ZN(n10914) );
  NAND2_X1 U8809 ( .A1(n16485), .A2(n25238), .ZN(n15698) );
  OR2_X1 U8834 ( .A1(n6135), .A2(n1798), .ZN(n2448) );
  NAND3_X1 U8898 ( .A1(n1594), .A2(n9282), .A3(n2953), .ZN(n9283) );
  NAND2_X1 U8899 ( .A1(n2248), .A2(n2249), .ZN(n19698) );
  BUF_X1 U8925 ( .A(n17421), .Z(n24330) );
  AOI22_X1 U8926 ( .A1(n23847), .A2(n24218), .B1(n23850), .B2(n23849), .ZN(
        n23856) );
  NAND3_X1 U8959 ( .A1(n23851), .A2(n25240), .A3(n3183), .ZN(n24218) );
  NAND2_X1 U8961 ( .A1(n24096), .A2(n24219), .ZN(n34) );
  AOI21_X1 U8972 ( .B1(n4499), .B2(n13234), .A(n24220), .ZN(n24219) );
  NOR2_X1 U9054 ( .A1(n25393), .A2(n24221), .ZN(n1886) );
  NAND2_X1 U9055 ( .A1(n24222), .A2(n9772), .ZN(n24221) );
  INV_X1 U9087 ( .A(n10109), .ZN(n24222) );
  OAI211_X1 U9108 ( .C1(n11122), .C2(n11123), .A(n24223), .B(n11121), .ZN(
        n10462) );
  INV_X1 U9122 ( .A(n10850), .ZN(n24223) );
  NOR2_X2 U9153 ( .A1(n2994), .A2(n9230), .ZN(n10850) );
  AND2_X2 U9231 ( .A1(n24525), .A2(n3153), .ZN(n7217) );
  NAND2_X1 U9242 ( .A1(n14154), .A2(n2775), .ZN(n1025) );
  NAND2_X1 U9287 ( .A1(n7346), .A2(n7349), .ZN(n24224) );
  INV_X1 U9298 ( .A(n17197), .ZN(n16869) );
  NAND2_X1 U9310 ( .A1(n17399), .A2(n17198), .ZN(n17197) );
  NAND2_X1 U9327 ( .A1(n9615), .A2(n9757), .ZN(n24225) );
  INV_X1 U9338 ( .A(n6575), .ZN(n443) );
  NAND2_X1 U9348 ( .A1(n24089), .A2(n6575), .ZN(n4973) );
  NAND3_X1 U9357 ( .A1(n5596), .A2(n4054), .A3(n24226), .ZN(n17341) );
  NAND3_X1 U9379 ( .A1(n613), .A2(n16062), .A3(n24227), .ZN(n24226) );
  NAND2_X1 U9418 ( .A1(n16780), .A2(n17241), .ZN(n24229) );
  NAND2_X1 U9440 ( .A1(n3661), .A2(n3662), .ZN(n3660) );
  OAI21_X1 U9570 ( .B1(n16141), .B2(n24231), .A(n24230), .ZN(n16144) );
  NAND2_X1 U9584 ( .A1(n16141), .A2(n16412), .ZN(n24230) );
  INV_X1 U9591 ( .A(n16140), .ZN(n24231) );
  NAND2_X1 U9612 ( .A1(n19550), .A2(n19549), .ZN(n19551) );
  OAI22_X1 U9660 ( .A1(n19546), .A2(n19185), .B1(n24929), .B2(n19186), .ZN(
        n19550) );
  AOI21_X2 U9673 ( .B1(n649), .B2(n15694), .A(n24233), .ZN(n16550) );
  NAND2_X1 U9717 ( .A1(n24234), .A2(n6762), .ZN(n6763) );
  NAND2_X1 U9738 ( .A1(n1454), .A2(n7460), .ZN(n24234) );
  NAND2_X1 U9816 ( .A1(n3219), .A2(n5678), .ZN(n11310) );
  NAND2_X1 U9818 ( .A1(n3220), .A2(n24168), .ZN(n3219) );
  NAND2_X2 U9833 ( .A1(n10773), .A2(n10776), .ZN(n11101) );
  NAND2_X1 U9836 ( .A1(n9494), .A2(n10020), .ZN(n10773) );
  AND3_X2 U9858 ( .A1(n22470), .A2(n22471), .A3(n22469), .ZN(n23120) );
  NAND2_X1 U9865 ( .A1(n24238), .A2(n24236), .ZN(n22850) );
  NOR2_X1 U9890 ( .A1(n22901), .A2(n22900), .ZN(n24237) );
  INV_X1 U9927 ( .A(n22842), .ZN(n24239) );
  INV_X1 U9943 ( .A(n16782), .ZN(n16777) );
  NAND2_X1 U9965 ( .A1(n17346), .A2(n17341), .ZN(n16782) );
  NAND2_X1 U9975 ( .A1(n3213), .A2(n22972), .ZN(n21891) );
  NAND3_X1 U9984 ( .A1(n10207), .A2(n10206), .A3(n10434), .ZN(n11263) );
  NAND2_X1 U10081 ( .A1(n24240), .A2(n10836), .ZN(n547) );
  NAND2_X1 U10085 ( .A1(n10276), .A2(n10275), .ZN(n24240) );
  NAND3_X1 U10141 ( .A1(n13065), .A2(n13162), .A3(n12736), .ZN(n2859) );
  XNOR2_X1 U10150 ( .A(n1821), .B(n11991), .ZN(n11994) );
  OR2_X1 U10173 ( .A1(n2464), .A2(n18809), .ZN(n18166) );
  NAND2_X1 U10174 ( .A1(n16775), .A2(n17048), .ZN(n1908) );
  NAND2_X1 U10197 ( .A1(n22466), .A2(n3938), .ZN(n24242) );
  XNOR2_X2 U10211 ( .A(n20809), .B(n20810), .ZN(n22462) );
  NAND2_X1 U10233 ( .A1(n16923), .A2(n16924), .ZN(n16926) );
  NAND2_X1 U10235 ( .A1(n17320), .A2(n17321), .ZN(n16924) );
  NAND2_X1 U10288 ( .A1(n7009), .A2(n7006), .ZN(n5982) );
  NAND2_X1 U10298 ( .A1(n19482), .A2(n19477), .ZN(n24243) );
  NAND2_X1 U10326 ( .A1(n19478), .A2(n24803), .ZN(n24244) );
  NAND2_X2 U10463 ( .A1(n2840), .A2(n12605), .ZN(n14852) );
  NAND3_X2 U10464 ( .A1(n3463), .A2(n5640), .A3(n5642), .ZN(n14858) );
  NAND2_X1 U10495 ( .A1(n4350), .A2(n22336), .ZN(n4349) );
  MUX2_X2 U10515 ( .A(n15813), .B(n15812), .S(n24061), .Z(n17729) );
  NAND3_X1 U10517 ( .A1(n17001), .A2(n17002), .A3(n17003), .ZN(n17004) );
  NAND2_X1 U10524 ( .A1(n2613), .A2(n17048), .ZN(n17003) );
  NAND3_X1 U10530 ( .A1(n15949), .A2(n15948), .A3(n15947), .ZN(n17050) );
  NAND3_X1 U10532 ( .A1(n24246), .A2(n6298), .A3(n6174), .ZN(n6212) );
  NAND2_X1 U10562 ( .A1(n6209), .A2(n6296), .ZN(n24246) );
  NAND2_X1 U10574 ( .A1(n1730), .A2(n1729), .ZN(n24247) );
  INV_X1 U10578 ( .A(n23235), .ZN(n5081) );
  AOI22_X1 U10600 ( .A1(n23245), .A2(n23235), .B1(n23250), .B2(n23249), .ZN(
        n22650) );
  NAND3_X1 U10606 ( .A1(n10840), .A2(n5101), .A3(n10470), .ZN(n10472) );
  NAND2_X1 U10618 ( .A1(n6864), .A2(n7148), .ZN(n6865) );
  NAND2_X1 U10619 ( .A1(n4365), .A2(n4366), .ZN(n6864) );
  NAND2_X1 U10634 ( .A1(n15625), .A2(n16096), .ZN(n24248) );
  NAND2_X1 U10639 ( .A1(n17160), .A2(n24250), .ZN(n17169) );
  NAND3_X1 U10670 ( .A1(n10740), .A2(n10854), .A3(n10858), .ZN(n24251) );
  NAND2_X1 U10696 ( .A1(n16777), .A2(n17342), .ZN(n1883) );
  OAI22_X1 U10715 ( .A1(n19525), .A2(n19526), .B1(n19521), .B2(n24252), .ZN(
        n19527) );
  NAND2_X1 U10737 ( .A1(n6533), .A2(n24253), .ZN(n6264) );
  INV_X1 U10769 ( .A(n6530), .ZN(n24253) );
  INV_X1 U10778 ( .A(n4199), .ZN(n24254) );
  NOR2_X1 U10842 ( .A1(n7776), .A2(n7526), .ZN(n2807) );
  AOI21_X2 U10859 ( .B1(n6125), .B2(n6124), .A(n24255), .ZN(n7776) );
  AND2_X1 U10882 ( .A1(n9435), .A2(n9433), .ZN(n9712) );
  OAI211_X1 U10914 ( .C1(n6702), .C2(n6553), .A(n24256), .B(n6960), .ZN(n7930)
         );
  NAND2_X1 U10917 ( .A1(n6702), .A2(n24257), .ZN(n24256) );
  NAND3_X1 U10931 ( .A1(n10095), .A2(n10098), .A3(n10099), .ZN(n10101) );
  XNOR2_X1 U10935 ( .A(n11424), .B(n2989), .ZN(n11425) );
  NAND2_X1 U10962 ( .A1(n14157), .A2(n13955), .ZN(n3303) );
  OR2_X1 U10969 ( .A1(n12901), .A2(n12928), .ZN(n24258) );
  NAND2_X1 U10980 ( .A1(n10134), .A2(n24026), .ZN(n10145) );
  OAI211_X2 U10981 ( .C1(n10562), .C2(n10561), .A(n10560), .B(n4540), .ZN(
        n12200) );
  NAND2_X1 U11025 ( .A1(n806), .A2(n7962), .ZN(n5163) );
  NAND2_X1 U11043 ( .A1(n24260), .A2(n2972), .ZN(n8635) );
  NAND2_X1 U11088 ( .A1(n6924), .A2(n1176), .ZN(n2355) );
  NAND2_X1 U11091 ( .A1(n9233), .A2(n9234), .ZN(n3705) );
  NAND2_X1 U11100 ( .A1(n12827), .A2(n24476), .ZN(n2915) );
  OAI211_X1 U11112 ( .C1(n21870), .C2(n21869), .A(n24261), .B(n21868), .ZN(
        Ciphertext[172]) );
  OAI211_X1 U11121 ( .C1(n21869), .C2(n21866), .A(n21865), .B(n21864), .ZN(
        n24261) );
  NAND2_X1 U11148 ( .A1(n416), .A2(n11038), .ZN(n9130) );
  NAND2_X1 U11155 ( .A1(n24262), .A2(n6067), .ZN(n6068) );
  OAI22_X1 U11156 ( .A1(n22933), .A2(n22853), .B1(n22498), .B2(n25004), .ZN(
        n21871) );
  NAND2_X1 U11157 ( .A1(n23336), .A2(n23334), .ZN(n22853) );
  NAND2_X1 U11259 ( .A1(n9935), .A2(n9938), .ZN(n24264) );
  NAND2_X1 U11260 ( .A1(n9936), .A2(n24511), .ZN(n24265) );
  NOR2_X2 U11272 ( .A1(n16724), .A2(n16723), .ZN(n2667) );
  NAND2_X1 U11290 ( .A1(n16721), .A2(n16931), .ZN(n24267) );
  NAND3_X1 U11317 ( .A1(n22669), .A2(n22670), .A3(n22668), .ZN(n22673) );
  NAND2_X1 U11437 ( .A1(n7590), .A2(n7464), .ZN(n7460) );
  OR2_X2 U11451 ( .A1(n5942), .A2(n5941), .ZN(n7590) );
  XNOR2_X1 U11551 ( .A(n24270), .B(n8761), .ZN(Ciphertext[82]) );
  NAND2_X1 U11678 ( .A1(n19305), .A2(n19306), .ZN(n24272) );
  NAND2_X1 U11682 ( .A1(n19304), .A2(n19133), .ZN(n19306) );
  NAND2_X1 U11737 ( .A1(n24273), .A2(n24091), .ZN(n6708) );
  NAND2_X1 U11786 ( .A1(n6702), .A2(n6705), .ZN(n24273) );
  NAND3_X1 U11810 ( .A1(n6911), .A2(n6916), .A3(n6286), .ZN(n6288) );
  OR2_X1 U11847 ( .A1(n14052), .A2(n12821), .ZN(n12822) );
  NOR2_X1 U11848 ( .A1(n25059), .A2(n23206), .ZN(n4230) );
  NAND3_X1 U11958 ( .A1(n6064), .A2(n6061), .A3(n6731), .ZN(n2401) );
  NAND2_X1 U12016 ( .A1(n20482), .A2(n24275), .ZN(n24274) );
  NAND3_X1 U12084 ( .A1(n6028), .A2(n6278), .A3(n25398), .ZN(n24276) );
  AND2_X1 U12088 ( .A1(n25210), .A2(n16381), .ZN(n692) );
  NAND2_X1 U12101 ( .A1(n25179), .A2(n22578), .ZN(n24279) );
  INV_X1 U12122 ( .A(n1797), .ZN(n24280) );
  NAND2_X1 U12188 ( .A1(n24283), .A2(n4804), .ZN(n4800) );
  NAND2_X1 U12251 ( .A1(n7057), .A2(n7738), .ZN(n24283) );
  NAND2_X1 U12261 ( .A1(n24285), .A2(n24284), .ZN(n9720) );
  NAND2_X1 U12272 ( .A1(n11149), .A2(n24479), .ZN(n24284) );
  NAND2_X1 U12337 ( .A1(n10690), .A2(n24286), .ZN(n24285) );
  NAND3_X2 U12448 ( .A1(n24291), .A2(n24288), .A3(n210), .ZN(n21306) );
  NAND2_X1 U12599 ( .A1(n1936), .A2(n20071), .ZN(n24291) );
  NAND2_X1 U12664 ( .A1(n16241), .A2(n24293), .ZN(n24292) );
  INV_X1 U12716 ( .A(n16440), .ZN(n24293) );
  NAND2_X1 U12721 ( .A1(n15945), .A2(n16440), .ZN(n24294) );
  INV_X1 U12815 ( .A(n6596), .ZN(n6597) );
  NAND2_X1 U12865 ( .A1(n6823), .A2(n6827), .ZN(n6596) );
  NAND2_X1 U12866 ( .A1(n9131), .A2(n9130), .ZN(n24295) );
  BUF_X1 U12869 ( .A(n1363), .Z(n24367) );
  XOR2_X1 U12897 ( .A(n112), .B(n15075), .Z(n24303) );
  NAND3_X1 U12899 ( .A1(n6607), .A2(n6609), .A3(n6610), .ZN(n4018) );
  NAND2_X1 U12915 ( .A1(n19208), .A2(n19024), .ZN(n835) );
  OAI21_X1 U12952 ( .B1(n13356), .B2(n13993), .A(n24296), .ZN(n13369) );
  NAND2_X1 U12953 ( .A1(n13993), .A2(n795), .ZN(n24296) );
  NOR2_X2 U13053 ( .A1(n635), .A2(n15559), .ZN(n16974) );
  NAND2_X1 U13054 ( .A1(n5698), .A2(n6323), .ZN(n5696) );
  NAND2_X1 U13136 ( .A1(n1577), .A2(n25064), .ZN(n9815) );
  INV_X1 U13217 ( .A(n3554), .ZN(n24297) );
  NAND3_X1 U13305 ( .A1(n17252), .A2(n17254), .A3(n24300), .ZN(n24299) );
  NAND2_X1 U13306 ( .A1(n2644), .A2(n19608), .ZN(n2643) );
  NAND2_X1 U13448 ( .A1(n328), .A2(n21794), .ZN(n5075) );
  NAND2_X1 U13473 ( .A1(n148), .A2(n546), .ZN(n11836) );
  NAND2_X1 U13657 ( .A1(n17051), .A2(n372), .ZN(n3643) );
  NAND2_X1 U13659 ( .A1(n14250), .A2(n24301), .ZN(n14260) );
  NAND3_X1 U13674 ( .A1(n19388), .A2(n19389), .A3(n19390), .ZN(n191) );
  NAND3_X1 U13812 ( .A1(n1062), .A2(n14090), .A3(n13607), .ZN(n1061) );
  NAND2_X1 U13816 ( .A1(n24302), .A2(n14059), .ZN(n12614) );
  NAND2_X1 U13817 ( .A1(n14278), .A2(n14850), .ZN(n24302) );
  NAND3_X1 U14125 ( .A1(n9429), .A2(n9984), .A3(n9982), .ZN(n471) );
  NAND2_X1 U14397 ( .A1(n10427), .A2(n3100), .ZN(n10430) );
  NAND2_X1 U14481 ( .A1(n1180), .A2(n10243), .ZN(n10427) );
  NAND2_X1 U14583 ( .A1(n1859), .A2(n1860), .ZN(n12639) );
  NAND3_X1 U14584 ( .A1(n794), .A2(n10055), .A3(n10056), .ZN(n11062) );
  NAND2_X1 U14637 ( .A1(n1122), .A2(n25441), .ZN(n987) );
  OAI211_X1 U14660 ( .C1(n9927), .C2(n9346), .A(n24304), .B(n9604), .ZN(n4730)
         );
  NAND2_X1 U14672 ( .A1(n9927), .A2(n24084), .ZN(n24304) );
  NAND2_X1 U14692 ( .A1(n20388), .A2(n19345), .ZN(n3165) );
  XOR2_X1 U14717 ( .A(n18098), .B(n18351), .Z(n18208) );
  AOI21_X1 U14718 ( .B1(n24317), .B2(n22950), .A(n22949), .ZN(n24343) );
  OR2_X1 U14793 ( .A1(n11114), .A2(n11112), .ZN(n9343) );
  OR2_X1 U14807 ( .A1(n24911), .A2(n22744), .ZN(n2199) );
  AOI21_X1 U14899 ( .B1(n20370), .B2(n19574), .A(n2016), .ZN(n21205) );
  NAND3_X1 U15014 ( .A1(n3483), .A2(n3481), .A3(n3477), .ZN(n24306) );
  XOR2_X1 U15070 ( .A(n21477), .B(n21222), .Z(n21970) );
  XNOR2_X1 U15071 ( .A(n21973), .B(n21972), .ZN(n22835) );
  CLKBUF_X1 U15079 ( .A(n23342), .Z(n24400) );
  CLKBUF_X1 U15081 ( .A(n22395), .Z(n24321) );
  XNOR2_X2 U15098 ( .A(n19870), .B(n19869), .ZN(n22231) );
  OAI21_X1 U15131 ( .B1(n16531), .B2(n16530), .A(n16529), .ZN(n18420) );
  INV_X1 U15182 ( .A(n23332), .ZN(n24309) );
  XOR2_X1 U15204 ( .A(n18418), .B(n18420), .Z(n18421) );
  INV_X1 U15206 ( .A(n4139), .ZN(n24310) );
  INV_X1 U15289 ( .A(n4139), .ZN(n19235) );
  XNOR2_X1 U15327 ( .A(n20746), .B(n20745), .ZN(n24311) );
  XNOR2_X1 U15328 ( .A(n18020), .B(n18019), .ZN(n24312) );
  AOI21_X1 U15366 ( .B1(n22910), .B2(n22909), .A(n22908), .ZN(n24313) );
  XNOR2_X1 U15405 ( .A(n18019), .B(n18020), .ZN(n19359) );
  AOI21_X1 U15458 ( .B1(n22910), .B2(n22909), .A(n22908), .ZN(n23529) );
  OR2_X1 U15580 ( .A1(n18941), .A2(n18940), .ZN(n24315) );
  OAI21_X1 U15708 ( .B1(n21882), .B2(n21881), .A(n21880), .ZN(n24316) );
  XOR2_X1 U15716 ( .A(n8183), .B(n8713), .Z(n8186) );
  OR2_X1 U15786 ( .A1(n22279), .A2(n22280), .ZN(n24317) );
  XNOR2_X1 U15944 ( .A(n20603), .B(n20604), .ZN(n5378) );
  XNOR2_X1 U15950 ( .A(n8290), .B(n8289), .ZN(n9806) );
  OAI21_X1 U16005 ( .B1(n25374), .B2(n18770), .A(n18769), .ZN(n20277) );
  XOR2_X1 U16015 ( .A(n17957), .B(n17956), .Z(n24318) );
  OR2_X1 U16212 ( .A1(n19673), .A2(n19672), .ZN(n24319) );
  CLKBUF_X1 U16256 ( .A(n23612), .Z(n24320) );
  MUX2_X1 U16275 ( .A(n19985), .B(n19986), .S(n2098), .Z(n19990) );
  INV_X1 U16286 ( .A(n3198), .ZN(n20194) );
  AND2_X1 U16397 ( .A1(n2674), .A2(n22946), .ZN(n24322) );
  XOR2_X1 U16670 ( .A(n8622), .B(n8058), .Z(n7042) );
  AND2_X1 U16729 ( .A1(n5678), .A2(n3219), .ZN(n24323) );
  XNOR2_X1 U16730 ( .A(n16502), .B(n16503), .ZN(n24324) );
  XNOR2_X1 U16763 ( .A(n16502), .B(n16503), .ZN(n19128) );
  AOI21_X1 U16837 ( .B1(n15725), .B2(n16457), .A(n16456), .ZN(n16849) );
  XNOR2_X1 U16846 ( .A(n4810), .B(n18505), .ZN(n24326) );
  NAND3_X1 U16882 ( .A1(n5501), .A2(n1458), .A3(n4363), .ZN(n24327) );
  XNOR2_X1 U17046 ( .A(n18505), .B(n4810), .ZN(n19397) );
  XOR2_X1 U17143 ( .A(n12364), .B(n12089), .Z(n24328) );
  XNOR2_X1 U17212 ( .A(n17376), .B(n17377), .ZN(n24329) );
  XNOR2_X1 U17215 ( .A(n17376), .B(n17377), .ZN(n19537) );
  OAI211_X1 U17225 ( .C1(n16196), .C2(n15901), .A(n5408), .B(n5407), .ZN(
        n17421) );
  BUF_X2 U17230 ( .A(n18596), .Z(n19177) );
  XNOR2_X1 U17235 ( .A(n8993), .B(n8992), .ZN(n24332) );
  NOR2_X1 U17237 ( .A1(n22431), .A2(n22432), .ZN(n24515) );
  BUF_X1 U17306 ( .A(n22205), .Z(n24333) );
  XNOR2_X1 U17312 ( .A(n20908), .B(n5503), .ZN(n22205) );
  NOR2_X2 U17332 ( .A1(n23514), .A2(n23517), .ZN(n23527) );
  XNOR2_X1 U17344 ( .A(n17975), .B(n5326), .ZN(n24335) );
  XNOR2_X1 U17492 ( .A(n17975), .B(n5326), .ZN(n19092) );
  XNOR2_X1 U17530 ( .A(n18403), .B(n18402), .ZN(n18788) );
  OR2_X1 U17555 ( .A1(n17886), .A2(n19471), .ZN(n3749) );
  AOI21_X1 U17612 ( .B1(n16695), .B2(n16694), .A(n16693), .ZN(n24337) );
  AOI21_X1 U17615 ( .B1(n16695), .B2(n16694), .A(n16693), .ZN(n17664) );
  NOR2_X1 U17706 ( .A1(n24933), .A2(n23394), .ZN(n24339) );
  NAND2_X1 U17956 ( .A1(n3863), .A2(n3864), .ZN(n24340) );
  BUF_X1 U18077 ( .A(n20904), .Z(n20727) );
  XNOR2_X1 U18109 ( .A(n21419), .B(n21418), .ZN(n24341) );
  XNOR2_X1 U18110 ( .A(n21419), .B(n21418), .ZN(n24342) );
  AOI21_X1 U18135 ( .B1(n24317), .B2(n22950), .A(n22949), .ZN(n23354) );
  OR2_X2 U18347 ( .A1(n4397), .A2(n4398), .ZN(n23714) );
  XNOR2_X1 U18364 ( .A(n18572), .B(n18571), .ZN(n19166) );
  XNOR2_X1 U18629 ( .A(n14493), .B(n4875), .ZN(n15280) );
  OAI211_X1 U18635 ( .C1(n12697), .C2(n13278), .A(n17), .B(n12696), .ZN(n24347) );
  XNOR2_X1 U18639 ( .A(n11972), .B(n11973), .ZN(n13278) );
  OAI211_X1 U18644 ( .C1(n12697), .C2(n13278), .A(n17), .B(n12696), .ZN(n14189) );
  AOI21_X1 U18714 ( .B1(n22131), .B2(n22968), .A(n22130), .ZN(n23263) );
  OR2_X1 U18776 ( .A1(n24075), .A2(n23064), .ZN(n24350) );
  XOR2_X1 U18815 ( .A(n15302), .B(n15301), .Z(n24352) );
  OR2_X1 U18962 ( .A1(n19593), .A2(n4479), .ZN(n24354) );
  INV_X2 U18997 ( .A(n23640), .ZN(n23649) );
  AND2_X2 U19039 ( .A1(n1007), .A2(n1006), .ZN(n23640) );
  INV_X1 U19073 ( .A(n22933), .ZN(n24356) );
  INV_X1 U19074 ( .A(n20960), .ZN(n24357) );
  XNOR2_X1 U19083 ( .A(n21525), .B(n22014), .ZN(n21308) );
  AND2_X1 U19088 ( .A1(n22853), .A2(n5421), .ZN(n602) );
  INV_X1 U19089 ( .A(n23265), .ZN(n24360) );
  XNOR2_X1 U19175 ( .A(n19624), .B(n19623), .ZN(n24362) );
  XNOR2_X1 U19189 ( .A(n19624), .B(n19623), .ZN(n21825) );
  BUF_X1 U19219 ( .A(n20102), .Z(n24370) );
  XOR2_X1 U19306 ( .A(n21733), .B(n21732), .Z(n24364) );
  XNOR2_X1 U19341 ( .A(n1103), .B(n1102), .ZN(n24366) );
  XNOR2_X1 U19342 ( .A(n1103), .B(n1102), .ZN(n16004) );
  XNOR2_X1 U19373 ( .A(n20796), .B(n21683), .ZN(n1363) );
  OR2_X1 U19390 ( .A1(n12529), .A2(n12528), .ZN(n24368) );
  XNOR2_X1 U19406 ( .A(n20850), .B(n20849), .ZN(n24369) );
  XNOR2_X1 U19445 ( .A(n20850), .B(n20849), .ZN(n23574) );
  OAI21_X2 U19575 ( .B1(n21657), .B2(n21656), .A(n21655), .ZN(n23374) );
  BUF_X1 U19707 ( .A(n18291), .Z(n24371) );
  INV_X1 U19726 ( .A(n23592), .ZN(n24372) );
  XNOR2_X1 U19728 ( .A(n10421), .B(n10420), .ZN(n24373) );
  XNOR2_X1 U19907 ( .A(n10421), .B(n10420), .ZN(n13169) );
  BUF_X1 U19950 ( .A(n23727), .Z(n24374) );
  INV_X1 U19986 ( .A(n12510), .ZN(n13185) );
  NAND3_X1 U20069 ( .A1(n13106), .A2(n13105), .A3(n13104), .ZN(n14100) );
  NAND2_X1 U20169 ( .A1(n22269), .A2(n2833), .ZN(n23251) );
  NAND3_X1 U20194 ( .A1(n5099), .A2(n3749), .A3(n3747), .ZN(n24378) );
  XNOR2_X2 U20244 ( .A(n21667), .B(n21666), .ZN(n22842) );
  XNOR2_X1 U20288 ( .A(n21002), .B(n21001), .ZN(n24379) );
  NOR2_X1 U20293 ( .A1(n23514), .A2(n23517), .ZN(n24380) );
  INV_X1 U20442 ( .A(n23697), .ZN(n24381) );
  INV_X1 U20607 ( .A(n23697), .ZN(n23721) );
  NAND3_X1 U20683 ( .A1(n2789), .A2(n2790), .A3(n16259), .ZN(n24384) );
  NAND2_X1 U20687 ( .A1(n15633), .A2(n3592), .ZN(n24385) );
  XNOR2_X1 U20785 ( .A(n16738), .B(n16737), .ZN(n24386) );
  XNOR2_X1 U20795 ( .A(n14796), .B(n14795), .ZN(n24387) );
  XNOR2_X1 U20811 ( .A(n14796), .B(n14795), .ZN(n2607) );
  NOR2_X1 U20922 ( .A1(n23579), .A2(n23578), .ZN(n24389) );
  NOR2_X1 U21000 ( .A1(n23579), .A2(n23578), .ZN(n24390) );
  INV_X1 U21023 ( .A(n2306), .ZN(n10685) );
  OR2_X1 U21024 ( .A1(n16256), .A2(n16255), .ZN(n24391) );
  NAND2_X1 U21025 ( .A1(n4434), .A2(n23001), .ZN(n24392) );
  XNOR2_X1 U21026 ( .A(n17493), .B(n17492), .ZN(n24393) );
  OAI21_X1 U21060 ( .B1(n22327), .B2(n22326), .A(n3682), .ZN(n24394) );
  XNOR2_X1 U21061 ( .A(n17493), .B(n17492), .ZN(n19270) );
  OAI21_X1 U21068 ( .B1(n22327), .B2(n22326), .A(n3682), .ZN(n23177) );
  INV_X1 U21096 ( .A(n1147), .ZN(n24395) );
  NOR2_X1 U21152 ( .A1(n21761), .A2(n23573), .ZN(n24397) );
  NOR2_X1 U21204 ( .A1(n21761), .A2(n23573), .ZN(n23566) );
  INV_X1 U21237 ( .A(n24386), .ZN(n24399) );
  OAI211_X1 U21261 ( .C1(n22960), .C2(n22959), .A(n4127), .B(n4126), .ZN(
        n23342) );
  OAI211_X1 U21263 ( .C1(n10958), .C2(n10699), .A(n10957), .B(n10956), .ZN(
        n24401) );
  OAI211_X1 U21279 ( .C1(n10958), .C2(n10699), .A(n10957), .B(n10956), .ZN(
        n11957) );
  AOI22_X1 U21303 ( .A1(n13354), .A2(n13353), .B1(n5588), .B2(n25430), .ZN(
        n13996) );
  XOR2_X1 U21306 ( .A(n14925), .B(n14924), .Z(n24403) );
  NOR2_X1 U21344 ( .A1(n21710), .A2(n695), .ZN(n24404) );
  NOR2_X1 U21372 ( .A1(n21710), .A2(n695), .ZN(n22987) );
  XNOR2_X1 U21413 ( .A(Key[44]), .B(Plaintext[44]), .ZN(n24405) );
  XNOR2_X1 U21541 ( .A(n18411), .B(n18410), .ZN(n24407) );
  AND2_X2 U21578 ( .A1(n24408), .A2(n24409), .ZN(n23064) );
  NOR2_X1 U21580 ( .A1(n21150), .A2(n570), .ZN(n24408) );
  OR2_X1 U21608 ( .A1(n21932), .A2(n22465), .ZN(n24409) );
  XNOR2_X1 U21624 ( .A(n18411), .B(n18410), .ZN(n19395) );
  NAND2_X1 U21643 ( .A1(n15835), .A2(n15836), .ZN(n24410) );
  XNOR2_X1 U21644 ( .A(n21475), .B(n21474), .ZN(n24411) );
  OAI21_X1 U21658 ( .B1(n21490), .B2(n21489), .A(n21488), .ZN(n24412) );
  XNOR2_X1 U21743 ( .A(n21475), .B(n21474), .ZN(n22967) );
  OAI21_X1 U21769 ( .B1(n21490), .B2(n21489), .A(n21488), .ZN(n23369) );
  XNOR2_X1 U21848 ( .A(n20635), .B(n20634), .ZN(n24415) );
  XNOR2_X1 U21986 ( .A(n20635), .B(n20634), .ZN(n22335) );
  BUF_X1 U22203 ( .A(n18301), .Z(n24416) );
  OAI211_X1 U22228 ( .C1(n16590), .C2(n17076), .A(n2374), .B(n2373), .ZN(
        n18301) );
  OAI21_X1 U22289 ( .B1(n13404), .B2(n13403), .A(n13402), .ZN(n24418) );
  OAI21_X1 U22445 ( .B1(n13404), .B2(n13403), .A(n13402), .ZN(n14591) );
  CLKBUF_X1 U22463 ( .A(n11005), .Z(n24420) );
  XNOR2_X1 U22698 ( .A(n16570), .B(n16571), .ZN(n24421) );
  XNOR2_X1 U22720 ( .A(n16571), .B(n16570), .ZN(n19556) );
  INV_X1 U22727 ( .A(n13328), .ZN(n24422) );
  NAND2_X1 U22757 ( .A1(n13891), .A2(n1819), .ZN(n24423) );
  XNOR2_X1 U22758 ( .A(n17800), .B(n17799), .ZN(n24424) );
  XNOR2_X1 U22896 ( .A(n17800), .B(n17799), .ZN(n19366) );
  AOI21_X1 U22930 ( .B1(n22841), .B2(n22840), .A(n22839), .ZN(n23398) );
  XOR2_X1 U22962 ( .A(n17549), .B(n17548), .Z(n24427) );
  INV_X1 U22965 ( .A(n23843), .ZN(n24428) );
  XNOR2_X1 U23005 ( .A(n14624), .B(n14623), .ZN(n24429) );
  XNOR2_X1 U23008 ( .A(n14624), .B(n14623), .ZN(n24430) );
  BUF_X1 U23163 ( .A(n17919), .Z(n24431) );
  AOI22_X1 U23290 ( .A1(n3306), .A2(n16546), .B1(n723), .B2(n283), .ZN(n17919)
         );
  OAI211_X1 U23368 ( .C1(n17275), .C2(n16690), .A(n16689), .B(n16688), .ZN(
        n24433) );
  OAI211_X1 U23393 ( .C1(n17275), .C2(n16690), .A(n16689), .B(n16688), .ZN(
        n17913) );
  NAND2_X1 U23405 ( .A1(n20912), .A2(n815), .ZN(n24434) );
  NOR2_X1 U23406 ( .A1(n23462), .A2(n22733), .ZN(n24435) );
  AOI21_X2 U23430 ( .B1(n6633), .B2(n6632), .A(n6631), .ZN(n7788) );
  OR2_X1 U23433 ( .A1(n16483), .A2(n25238), .ZN(n757) );
  XNOR2_X1 U23451 ( .A(n21100), .B(n21099), .ZN(n24439) );
  MUX2_X1 U23463 ( .A(n22777), .B(n22776), .S(n22677), .Z(n24440) );
  XNOR2_X1 U23465 ( .A(n21099), .B(n21100), .ZN(n23999) );
  XNOR2_X1 U23717 ( .A(n15555), .B(n15554), .ZN(n24441) );
  XNOR2_X1 U23760 ( .A(n15555), .B(n15554), .ZN(n19302) );
  INV_X1 U23772 ( .A(n2710), .ZN(n24442) );
  OAI21_X1 U23807 ( .B1(n16395), .B2(n16394), .A(n16396), .ZN(n24444) );
  OAI21_X1 U23808 ( .B1(n16395), .B2(n16394), .A(n16396), .ZN(n17438) );
  OAI21_X1 U23979 ( .B1(n7936), .B2(n7935), .A(n7934), .ZN(n24445) );
  XNOR2_X1 U23981 ( .A(n9056), .B(n9055), .ZN(n24446) );
  OAI21_X1 U23989 ( .B1(n7936), .B2(n7935), .A(n7934), .ZN(n9195) );
  OAI211_X1 U24074 ( .C1(n22787), .C2(n24406), .A(n22786), .B(n22785), .ZN(
        n24448) );
  OAI211_X1 U24075 ( .C1(n22787), .C2(n24406), .A(n22786), .B(n22785), .ZN(
        n24010) );
  BUF_X1 U24076 ( .A(n23391), .Z(n24449) );
  OAI211_X1 U24077 ( .C1(n22030), .C2(n22029), .A(n5771), .B(n22028), .ZN(
        n23391) );
  XNOR2_X1 U24080 ( .A(n17724), .B(n17725), .ZN(n24451) );
  XOR2_X1 U24081 ( .A(n17964), .B(n17965), .Z(n24452) );
  XNOR2_X1 U24082 ( .A(n22006), .B(n21444), .ZN(n24453) );
  OAI21_X1 U24084 ( .B1(n19538), .B2(n24329), .A(n19536), .ZN(n24454) );
  XNOR2_X1 U24085 ( .A(n17530), .B(n17531), .ZN(n24457) );
  XNOR2_X1 U24086 ( .A(n15108), .B(n15107), .ZN(n16356) );
  XNOR2_X1 U24087 ( .A(n14371), .B(n14372), .ZN(n24458) );
  XNOR2_X1 U24088 ( .A(n14371), .B(n14372), .ZN(n24459) );
  OAI211_X1 U24089 ( .C1(n24926), .C2(n24582), .A(n19356), .B(n19355), .ZN(
        n24460) );
  OAI211_X1 U24090 ( .C1(n24926), .C2(n24582), .A(n19356), .B(n19355), .ZN(
        n24461) );
  OAI211_X1 U24091 ( .C1(n24926), .C2(n24582), .A(n19356), .B(n19355), .ZN(
        n20394) );
  CLKBUF_X1 U24092 ( .A(n13488), .Z(n24462) );
  INV_X1 U24093 ( .A(n20597), .ZN(n24463) );
  XNOR2_X1 U24094 ( .A(n14620), .B(n14721), .ZN(n15170) );
  NOR2_X1 U24095 ( .A1(n156), .A2(n18946), .ZN(n24464) );
  NOR2_X1 U24096 ( .A1(n156), .A2(n18946), .ZN(n19983) );
  NAND4_X1 U24097 ( .A1(n22024), .A2(n22022), .A3(n22023), .A4(n22025), .ZN(
        n24465) );
  NAND4_X1 U24098 ( .A1(n22024), .A2(n22022), .A3(n22023), .A4(n22025), .ZN(
        n23393) );
  XOR2_X1 U24099 ( .A(Key[6]), .B(Plaintext[6]), .Z(n24466) );
  XNOR2_X1 U24100 ( .A(n12619), .B(n12620), .ZN(n24467) );
  XNOR2_X1 U24101 ( .A(n12619), .B(n12620), .ZN(n16352) );
  XNOR2_X1 U24102 ( .A(n19161), .B(n19160), .ZN(n24468) );
  NOR2_X1 U24103 ( .A1(n19626), .A2(n19625), .ZN(n23858) );
  NOR2_X1 U24104 ( .A1(n2730), .A2(n8225), .ZN(n24470) );
  OAI21_X1 U24105 ( .B1(n15976), .B2(n15975), .A(n15974), .ZN(n24471) );
  OAI21_X1 U24107 ( .B1(n15976), .B2(n15975), .A(n15974), .ZN(n17573) );
  OR2_X1 U24108 ( .A1(n4846), .A2(n16357), .ZN(n18) );
  MUX2_X2 U24109 ( .A(n22136), .B(n22135), .S(n22401), .Z(n23281) );
  NOR2_X1 U24110 ( .A1(n19673), .A2(n19672), .ZN(n24472) );
  NOR2_X1 U24112 ( .A1(n19673), .A2(n19672), .ZN(n21649) );
  OAI21_X1 U24113 ( .B1(n21374), .B2(n21373), .A(n21372), .ZN(n23153) );
  OAI21_X1 U24114 ( .B1(n6880), .B2(n6879), .A(n1888), .ZN(n24474) );
  OAI21_X1 U24115 ( .B1(n6880), .B2(n6879), .A(n1888), .ZN(n24475) );
  OAI21_X1 U24116 ( .B1(n6880), .B2(n6879), .A(n1888), .ZN(n7948) );
  INV_X1 U24117 ( .A(n24931), .ZN(n24477) );
  XNOR2_X1 U24118 ( .A(n17761), .B(n17760), .ZN(n19386) );
  OAI211_X1 U24119 ( .C1(n2079), .C2(n9687), .A(n9685), .B(n9686), .ZN(n24479)
         );
  OAI211_X1 U24120 ( .C1(n2079), .C2(n9687), .A(n9685), .B(n9686), .ZN(n24480)
         );
  INV_X1 U24121 ( .A(n19581), .ZN(n24481) );
  OAI211_X1 U24122 ( .C1(n2079), .C2(n9687), .A(n9685), .B(n9686), .ZN(n11152)
         );
  XNOR2_X1 U24123 ( .A(n15222), .B(n15221), .ZN(n24482) );
  XNOR2_X1 U24124 ( .A(n18072), .B(n18071), .ZN(n24483) );
  XNOR2_X1 U24125 ( .A(n18072), .B(n18071), .ZN(n19590) );
  OR2_X1 U24126 ( .A1(n22222), .A2(n24484), .ZN(n1237) );
  OR2_X1 U24127 ( .A1(n22220), .A2(n22219), .ZN(n24484) );
  OAI21_X1 U24129 ( .B1(n20323), .B2(n20322), .A(n20321), .ZN(n20882) );
  OAI211_X1 U24130 ( .C1(n16709), .C2(n16708), .A(n16707), .B(n2057), .ZN(
        n24488) );
  OAI211_X1 U24132 ( .C1(n16709), .C2(n16708), .A(n16707), .B(n2057), .ZN(
        n18678) );
  XNOR2_X1 U24133 ( .A(n11731), .B(n11730), .ZN(n24490) );
  XNOR2_X1 U24134 ( .A(n11731), .B(n11730), .ZN(n13221) );
  OAI211_X1 U24135 ( .C1(n20564), .C2(n25221), .A(n4009), .B(n19734), .ZN(
        n21455) );
  NAND2_X1 U24136 ( .A1(n24493), .A2(n24494), .ZN(n23357) );
  OR3_X1 U24137 ( .A1(n22961), .A2(n24492), .A3(n23359), .ZN(n24493) );
  OR3_X1 U24138 ( .A1(n23361), .A2(n23350), .A3(n23349), .ZN(n24494) );
  XNOR2_X1 U24139 ( .A(n15227), .B(n15228), .ZN(n16191) );
  XOR2_X1 U24144 ( .A(n10300), .B(n10299), .Z(n24499) );
  XNOR2_X1 U24145 ( .A(n5780), .B(Key[95]), .ZN(n24500) );
  XNOR2_X1 U24146 ( .A(n5780), .B(Key[95]), .ZN(n24501) );
  OAI211_X1 U24147 ( .C1(n14012), .C2(n14011), .A(n856), .B(n855), .ZN(n24502)
         );
  XNOR2_X1 U24148 ( .A(n5780), .B(Key[95]), .ZN(n6715) );
  OAI211_X1 U24149 ( .C1(n14012), .C2(n14011), .A(n856), .B(n855), .ZN(n15138)
         );
  XNOR2_X1 U24153 ( .A(n8547), .B(n8546), .ZN(n24505) );
  XNOR2_X1 U24154 ( .A(n15014), .B(n15013), .ZN(n24506) );
  XNOR2_X1 U24155 ( .A(n8547), .B(n8546), .ZN(n9781) );
  OAI211_X1 U24156 ( .C1(n13711), .C2(n13394), .A(n11681), .B(n11680), .ZN(
        n15401) );
  BUF_X1 U24158 ( .A(n15229), .Z(n24508) );
  AOI22_X2 U24159 ( .A1(n4601), .A2(n3727), .B1(n19017), .B2(n19393), .ZN(
        n20445) );
  XNOR2_X1 U24160 ( .A(Key[156]), .B(Plaintext[156]), .ZN(n24509) );
  XNOR2_X1 U24161 ( .A(n11231), .B(n11230), .ZN(n24512) );
  XNOR2_X1 U24162 ( .A(n11231), .B(n11230), .ZN(n24513) );
  XNOR2_X1 U24163 ( .A(n8027), .B(n8028), .ZN(n9450) );
  AND4_X1 U24164 ( .A1(n10442), .A2(n2766), .A3(n10440), .A4(n10441), .ZN(
        n24514) );
  NOR2_X1 U24165 ( .A1(n22431), .A2(n22432), .ZN(n23371) );
  XNOR2_X2 U24166 ( .A(n10449), .B(n10450), .ZN(n4766) );
  XNOR2_X1 U24168 ( .A(n17222), .B(n17221), .ZN(n24516) );
  NOR2_X1 U24170 ( .A1(n22802), .A2(n22659), .ZN(n24517) );
  AND2_X1 U24171 ( .A1(n2978), .A2(n22664), .ZN(n24518) );
  NAND2_X1 U24172 ( .A1(n23363), .A2(n23362), .ZN(n23364) );
  NAND2_X1 U24173 ( .A1(n1802), .A2(n1803), .ZN(n22839) );
  NAND3_X1 U24174 ( .A1(n24520), .A2(n13434), .A3(n24519), .ZN(n14654) );
  NAND2_X1 U24175 ( .A1(n13432), .A2(n14106), .ZN(n24520) );
  NAND2_X1 U24176 ( .A1(n24521), .A2(n10486), .ZN(n9608) );
  NAND2_X1 U24178 ( .A1(n12687), .A2(n24522), .ZN(n13322) );
  NAND2_X1 U24179 ( .A1(n12945), .A2(n12942), .ZN(n24522) );
  NAND2_X1 U24182 ( .A1(n281), .A2(n17012), .ZN(n17357) );
  OR2_X1 U24183 ( .A1(n6369), .A2(n6071), .ZN(n7003) );
  NAND3_X1 U24184 ( .A1(n5389), .A2(n5390), .A3(n7628), .ZN(n5388) );
  NAND2_X1 U24185 ( .A1(n11101), .A2(n10914), .ZN(n11031) );
  NAND3_X1 U24186 ( .A1(n5312), .A2(n5311), .A3(n5313), .ZN(n5310) );
  AOI22_X1 U24187 ( .A1(n6200), .A2(n6909), .B1(n6201), .B2(n6774), .ZN(n2784)
         );
  NAND2_X1 U24190 ( .A1(n6436), .A2(n25325), .ZN(n24525) );
  NAND2_X1 U24191 ( .A1(n620), .A2(n4844), .ZN(n619) );
  AND2_X1 U24192 ( .A1(n10630), .A2(n10789), .ZN(n24526) );
  OR2_X1 U24193 ( .A1(n12807), .A2(n12808), .ZN(n24527) );
  OR2_X1 U24195 ( .A1(n16128), .A2(n16154), .ZN(n24528) );
  BUF_X1 U24196 ( .A(n17463), .Z(n288) );
  AND2_X1 U24198 ( .A1(n17016), .A2(n17212), .ZN(n24529) );
  INV_X1 U24199 ( .A(n19357), .ZN(n19037) );
  NAND3_X1 U24201 ( .A1(n4017), .A2(n20567), .A3(n20562), .ZN(n24530) );
  NOR2_X1 U24202 ( .A1(n3428), .A2(n349), .ZN(n24531) );
  XNOR2_X2 U8837 ( .A(n3506), .B(n8104), .ZN(n9899) );
  OAI21_X2 U2447 ( .B1(n10157), .B2(n9854), .A(n9350), .ZN(n1499) );
  NAND2_X2 U658 ( .A1(n6185), .A2(n6186), .ZN(n7647) );
  AND3_X2 U1944 ( .A1(n7117), .A2(n5689), .A3(n5691), .ZN(n8616) );
  XNOR2_X2 U2159 ( .A(n15372), .B(n15373), .ZN(n16060) );
  BUF_X2 U3222 ( .A(n19155), .Z(n21038) );
  AOI21_X2 U1152 ( .B1(n22512), .B2(n25496), .A(n22511), .ZN(n23181) );
  NAND4_X2 U2369 ( .A1(n10864), .A2(n10866), .A3(n10865), .A4(n10863), .ZN(
        n12096) );
  OR2_X2 U8717 ( .A1(n9546), .A2(n9545), .ZN(n10445) );
  XNOR2_X2 U1330 ( .A(n12014), .B(n12015), .ZN(n13264) );
  BUF_X1 U2047 ( .A(n16849), .Z(n16985) );
  AND2_X2 U1841 ( .A1(n5473), .A2(n5476), .ZN(n20255) );
  NAND3_X2 U7009 ( .A1(n5750), .A2(n1930), .A3(n1395), .ZN(n14919) );
  BUF_X2 U15937 ( .A(n11411), .Z(n13909) );
  XNOR2_X2 U12115 ( .A(Key[77]), .B(Plaintext[77]), .ZN(n6051) );
  AOI21_X2 U6823 ( .B1(n9720), .B2(n9719), .A(n204), .ZN(n11967) );
  AND2_X2 U3690 ( .A1(n893), .A2(n1572), .ZN(n13785) );
  NAND4_X2 U80 ( .A1(n10797), .A2(n10796), .A3(n10795), .A4(n10794), .ZN(
        n12401) );
  AOI22_X2 U1447 ( .A1(n15690), .A2(n16472), .B1(n15688), .B2(n15689), .ZN(
        n16551) );
  XNOR2_X2 U1521 ( .A(n8101), .B(n8100), .ZN(n2294) );
  BUF_X1 U224 ( .A(n10135), .Z(n24025) );
  BUF_X2 U14020 ( .A(n9348), .Z(n10162) );
  NOR2_X2 U1056 ( .A1(n15872), .A2(n15871), .ZN(n17084) );
  INV_X2 U144 ( .A(n16121), .ZN(n16122) );
  BUF_X1 U2151 ( .A(n5992), .Z(n6824) );
  AND3_X2 U192 ( .A1(n2124), .A2(n3770), .A3(n3768), .ZN(n2602) );
  MUX2_X2 U1684 ( .A(n22605), .B(n22604), .S(n22603), .Z(n23050) );
  BUF_X1 U820 ( .A(n23119), .Z(n24059) );
  AND2_X2 U7560 ( .A1(n4888), .A2(n17358), .ZN(n18123) );
  NAND4_X2 U807 ( .A1(n5602), .A2(n5601), .A3(n7737), .A4(n5600), .ZN(n8690)
         );
  INV_X1 U200 ( .A(n10861), .ZN(n10190) );
  NOR2_X1 U2472 ( .A1(n307), .A2(n9692), .ZN(n9880) );
  NAND2_X2 U4749 ( .A1(n20380), .A2(n24127), .ZN(n21633) );
  BUF_X1 U2297 ( .A(n12433), .Z(n13137) );
  BUF_X2 U16266 ( .A(n11805), .Z(n13968) );
  NAND2_X2 U9360 ( .A1(n16190), .A2(n3222), .ZN(n17185) );
  OAI211_X2 U1423 ( .C1(n16675), .C2(n16876), .A(n16674), .B(n16673), .ZN(
        n18674) );
  NAND2_X2 U336 ( .A1(n2897), .A2(n2896), .ZN(n8699) );
  AND2_X2 U988 ( .A1(n15918), .A2(n15919), .ZN(n17364) );
  BUF_X1 U1918 ( .A(n18749), .Z(n19138) );
  OAI21_X2 U416 ( .B1(n9262), .B2(n9858), .A(n9261), .ZN(n10737) );
  NAND4_X2 U2208 ( .A1(n870), .A2(n14248), .A3(n14247), .A4(n14246), .ZN(
        n14907) );
  INV_X2 U1929 ( .A(n4667), .ZN(n19476) );
  OAI211_X2 U1503 ( .C1(n3575), .C2(n10905), .A(n4343), .B(n3574), .ZN(n12159)
         );
  XNOR2_X2 U17911 ( .A(n14540), .B(n14539), .ZN(n16391) );
  AOI21_X2 U14876 ( .B1(n20370), .B2(n19574), .A(n2016), .ZN(n24305) );
  XNOR2_X1 U2163 ( .A(n14991), .B(n14990), .ZN(n16022) );
  BUF_X2 U2512 ( .A(n9495), .Z(n10090) );
  INV_X1 U5891 ( .A(n19494), .ZN(n20235) );
  OR2_X2 U403 ( .A1(n15754), .A2(n15753), .ZN(n16902) );
  XNOR2_X2 U15697 ( .A(n11182), .B(n11183), .ZN(n12455) );
  BUF_X2 U1864 ( .A(n19851), .Z(n19660) );
  AOI22_X2 U19440 ( .A1(n16919), .A2(n16918), .B1(n16917), .B2(n16916), .ZN(
        n17582) );
  AND2_X1 U12025 ( .A1(n25197), .A2(n14335), .ZN(n14344) );
  NAND3_X2 U6931 ( .A1(n7343), .A2(n7344), .A3(n1999), .ZN(n8964) );
  XNOR2_X1 U3491 ( .A(n15256), .B(n15257), .ZN(n2610) );
  NAND3_X2 U10956 ( .A1(n4156), .A2(n10621), .A3(n3724), .ZN(n11424) );
  XNOR2_X1 U2927 ( .A(n15108), .B(n15107), .ZN(n24456) );
  AND2_X2 U1987 ( .A1(n567), .A2(n566), .ZN(n18334) );
  OAI211_X2 U13340 ( .C1(n7445), .C2(n7375), .A(n7374), .B(n7373), .ZN(n9182)
         );
  AND2_X2 U1420 ( .A1(n3784), .A2(n2641), .ZN(n18128) );
  INV_X1 U19856 ( .A(n17653), .ZN(n18601) );
  XNOR2_X2 U1787 ( .A(n20967), .B(n20968), .ZN(n22918) );
  NOR2_X1 U22755 ( .A1(n25239), .A2(n23890), .ZN(n23909) );
  INV_X1 U19259 ( .A(n16660), .ZN(n17198) );
  OAI21_X1 U18758 ( .B1(n15709), .B2(n15708), .A(n2636), .ZN(n15713) );
  XNOR2_X1 U12417 ( .A(Key[178]), .B(Plaintext[178]), .ZN(n6467) );
  XNOR2_X1 U12357 ( .A(Key[188]), .B(Plaintext[188]), .ZN(n6452) );
  XNOR2_X1 U12478 ( .A(Key[97]), .B(Plaintext[97]), .ZN(n6588) );
  CLKBUF_X1 U1656 ( .A(Key[3]), .Z(n21169) );
  XNOR2_X1 U2735 ( .A(Key[20]), .B(Plaintext[20]), .ZN(n6165) );
  CLKBUF_X1 U1210 ( .A(Key[117]), .Z(n1870) );
  CLKBUF_X1 U348 ( .A(Key[89]), .Z(n3093) );
  XNOR2_X1 U12472 ( .A(Key[115]), .B(Plaintext[115]), .ZN(n7021) );
  XNOR2_X1 U4341 ( .A(Key[100]), .B(Plaintext[100]), .ZN(n7035) );
  CLKBUF_X1 U1352 ( .A(Key[14]), .Z(n21335) );
  CLKBUF_X1 U1601 ( .A(Key[161]), .Z(n2031) );
  XNOR2_X1 U2739 ( .A(Key[139]), .B(Plaintext[139]), .ZN(n6794) );
  XNOR2_X1 U12168 ( .A(Key[78]), .B(Plaintext[78]), .ZN(n6396) );
  CLKBUF_X1 U1208 ( .A(Key[100]), .Z(n16) );
  CLKBUF_X1 U1566 ( .A(Key[142]), .Z(n2040) );
  CLKBUF_X1 U1583 ( .A(Key[15]), .Z(n21742) );
  CLKBUF_X1 U2755 ( .A(Key[116]), .Z(n23983) );
  XNOR2_X1 U12146 ( .A(Key[62]), .B(Plaintext[62]), .ZN(n6969) );
  CLKBUF_X1 U2724 ( .A(Key[63]), .Z(n1896) );
  CLKBUF_X1 U1664 ( .A(Key[37]), .Z(n641) );
  CLKBUF_X1 U1203 ( .A(Key[137]), .Z(n21703) );
  CLKBUF_X1 U1581 ( .A(Key[158]), .Z(n23699) );
  XNOR2_X1 U12210 ( .A(Key[140]), .B(Plaintext[140]), .ZN(n6076) );
  XNOR2_X1 U5902 ( .A(Key[148]), .B(Plaintext[148]), .ZN(n6905) );
  CLKBUF_X1 U1600 ( .A(Key[0]), .Z(n836) );
  BUF_X1 U1551 ( .A(n6081), .Z(n6876) );
  XNOR2_X1 U12497 ( .A(n6023), .B(Key[17]), .ZN(n6275) );
  XNOR2_X1 U2713 ( .A(n495), .B(Key[65]), .ZN(n6570) );
  XNOR2_X1 U1076 ( .A(n5993), .B(Key[103]), .ZN(n6827) );
  XNOR2_X1 U12364 ( .A(n5931), .B(Key[191]), .ZN(n6187) );
  OAI211_X1 U16816 ( .C1(n7002), .C2(n7003), .A(n7001), .B(n7000), .ZN(n7962)
         );
  OR2_X1 U880 ( .A1(n873), .A2(n6361), .ZN(n8367) );
  AOI22_X1 U924 ( .A1(n6902), .A2(n6475), .B1(n6476), .B2(n6905), .ZN(n8074)
         );
  OR2_X1 U2659 ( .A1(n5922), .A2(n5923), .ZN(n7351) );
  AND3_X1 U109 ( .A1(n2737), .A2(n5086), .A3(n2736), .ZN(n1345) );
  OR2_X1 U2631 ( .A1(n6831), .A2(n6830), .ZN(n7984) );
  NAND3_X1 U121 ( .A1(n4682), .A2(n4681), .A3(n6527), .ZN(n7211) );
  NAND3_X1 U10292 ( .A1(n6231), .A2(n4122), .A3(n4121), .ZN(n7642) );
  NAND3_X1 U7185 ( .A1(n2032), .A2(n6914), .A3(n6913), .ZN(n7942) );
  OR2_X1 U2652 ( .A1(n6118), .A2(n6117), .ZN(n7527) );
  INV_X1 U13005 ( .A(n7829), .ZN(n7048) );
  NAND3_X1 U3608 ( .A1(n6562), .A2(n6563), .A3(n6561), .ZN(n7444) );
  OR2_X1 U165 ( .A1(n4994), .A2(n436), .ZN(n7669) );
  OR2_X1 U2580 ( .A1(n7279), .A2(n8511), .ZN(n7254) );
  OR2_X1 U4426 ( .A1(n7540), .A2(n432), .ZN(n7547) );
  OR2_X1 U2578 ( .A1(n7845), .A2(n8374), .ZN(n9176) );
  NAND2_X1 U2564 ( .A1(n6863), .A2(n6862), .ZN(n9167) );
  NAND2_X1 U213 ( .A1(n6854), .A2(n6855), .ZN(n8687) );
  OAI21_X1 U9413 ( .B1(n4483), .B2(n3272), .A(n3363), .ZN(n8238) );
  OAI21_X1 U2563 ( .B1(n5861), .B2(n5860), .A(n5859), .ZN(n8666) );
  AND2_X1 U2550 ( .A1(n569), .A2(n533), .ZN(n5344) );
  NAND2_X1 U633 ( .A1(n1040), .A2(n1037), .ZN(n8874) );
  OR2_X1 U2554 ( .A1(n7712), .A2(n7711), .ZN(n8468) );
  INV_X1 U2547 ( .A(n5344), .ZN(n9139) );
  XNOR2_X1 U4439 ( .A(n8448), .B(n8983), .ZN(n9788) );
  XNOR2_X1 U1094 ( .A(n7876), .B(n7875), .ZN(n9939) );
  XNOR2_X1 U14331 ( .A(n8811), .B(n8810), .ZN(n10020) );
  XNOR2_X1 U2422 ( .A(n7744), .B(n7743), .ZN(n9925) );
  XNOR2_X1 U2530 ( .A(n9085), .B(n1385), .ZN(n4096) );
  BUF_X1 U1243 ( .A(n9859), .Z(n239) );
  XNOR2_X1 U4583 ( .A(n7906), .B(n7907), .ZN(n9449) );
  CLKBUF_X1 U11973 ( .A(n8141), .Z(n9961) );
  BUF_X1 U1044 ( .A(n9328), .Z(n9774) );
  XNOR2_X1 U11116 ( .A(n8380), .B(n8379), .ZN(n10094) );
  INV_X1 U14663 ( .A(n9297), .ZN(n10093) );
  MUX2_X1 U2504 ( .A(n9858), .B(n9280), .S(n239), .Z(n10516) );
  NOR2_X1 U2506 ( .A1(n9959), .A2(n9950), .ZN(n9392) );
  OAI211_X1 U2451 ( .C1(n10049), .C2(n10048), .A(n4068), .B(n1403), .ZN(n11067) );
  NAND2_X1 U10787 ( .A1(n10516), .A2(n10517), .ZN(n10275) );
  AND2_X1 U4872 ( .A1(n9392), .A2(n9951), .ZN(n10256) );
  AND4_X1 U1097 ( .A1(n9457), .A2(n9566), .A3(n957), .A4(n955), .ZN(n10887) );
  OR2_X1 U2465 ( .A1(n9298), .A2(n9498), .ZN(n2501) );
  NOR2_X1 U189 ( .A1(n10174), .A2(n10173), .ZN(n10398) );
  MUX2_X1 U9075 ( .A(n9701), .B(n9240), .S(n9700), .Z(n11149) );
  NAND3_X1 U91 ( .A1(n9371), .A2(n9369), .A3(n9370), .ZN(n10451) );
  NAND3_X1 U1509 ( .A1(n4207), .A2(n9508), .A3(n4210), .ZN(n939) );
  NAND4_X1 U417 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n11741) );
  NAND4_X1 U8420 ( .A1(n2766), .A2(n10440), .A3(n10442), .A4(n10441), .ZN(
        n11908) );
  OR2_X1 U1501 ( .A1(n10330), .A2(n10329), .ZN(n12134) );
  XNOR2_X1 U2556 ( .A(n11246), .B(n11245), .ZN(n13217) );
  XNOR2_X1 U11889 ( .A(n12254), .B(n12253), .ZN(n12272) );
  CLKBUF_X1 U2315 ( .A(n12600), .Z(n12966) );
  BUF_X1 U2312 ( .A(n11755), .Z(n13222) );
  INV_X1 U402 ( .A(n12674), .ZN(n4923) );
  AND2_X1 U530 ( .A1(n11350), .A2(n13213), .ZN(n13208) );
  OR2_X1 U4477 ( .A1(n13306), .A2(n13307), .ZN(n13310) );
  NOR2_X1 U2701 ( .A1(n13093), .A2(n12650), .ZN(n13669) );
  NAND3_X1 U645 ( .A1(n4867), .A2(n5012), .A3(n5010), .ZN(n14112) );
  AOI22_X1 U2284 ( .A1(n13239), .A2(n13238), .B1(n13237), .B2(n4493), .ZN(
        n13982) );
  MUX2_X1 U16926 ( .A(n12849), .B(n12848), .S(n301), .Z(n13504) );
  INV_X1 U2827 ( .A(n13775), .ZN(n14160) );
  AND3_X1 U2904 ( .A1(n12567), .A2(n12566), .A3(n5747), .ZN(n14076) );
  MUX2_X1 U17122 ( .A(n13287), .B(n13286), .S(n25191), .Z(n13923) );
  NAND2_X1 U2813 ( .A1(n13193), .A2(n13192), .ZN(n14106) );
  NAND2_X1 U815 ( .A1(n779), .A2(n12988), .ZN(n14222) );
  AND2_X1 U2246 ( .A1(n622), .A2(n624), .ZN(n13895) );
  OR2_X1 U340 ( .A1(n14126), .A2(n14129), .ZN(n13826) );
  NAND3_X1 U674 ( .A1(n2155), .A2(n985), .A3(n984), .ZN(n15298) );
  NAND2_X1 U2204 ( .A1(n14040), .A2(n5058), .ZN(n15095) );
  AND3_X1 U58 ( .A1(n3368), .A2(n3369), .A3(n3367), .ZN(n14815) );
  NAND2_X1 U337 ( .A1(n48), .A2(n4598), .ZN(n15183) );
  AND2_X1 U10812 ( .A1(n183), .A2(n185), .ZN(n15422) );
  XNOR2_X1 U1510 ( .A(n15505), .B(n24097), .ZN(n14909) );
  INV_X1 U18278 ( .A(n14977), .ZN(n15342) );
  BUF_X1 U2136 ( .A(n14926), .Z(n16277) );
  XNOR2_X1 U2175 ( .A(n15308), .B(n15307), .ZN(n16048) );
  XNOR2_X1 U853 ( .A(n15101), .B(n15100), .ZN(n16359) );
  BUF_X1 U141 ( .A(n14664), .Z(n16077) );
  BUF_X1 U2144 ( .A(n14625), .Z(n15789) );
  XNOR2_X1 U2135 ( .A(n3707), .B(n14918), .ZN(n16030) );
  BUF_X1 U1154 ( .A(n16149), .Z(n213) );
  NOR2_X1 U4495 ( .A1(n16025), .A2(n15773), .ZN(n16602) );
  AND2_X1 U2070 ( .A1(n14974), .A2(n14975), .ZN(n17409) );
  OAI211_X1 U1448 ( .C1(n4091), .C2(n16273), .A(n15771), .B(n4090), .ZN(n17425) );
  NOR2_X1 U1439 ( .A1(n13943), .A2(n13942), .ZN(n17419) );
  NAND3_X1 U8933 ( .A1(n3009), .A2(n3008), .A3(n15982), .ZN(n17042) );
  NAND3_X1 U2056 ( .A1(n4939), .A2(n14666), .A3(n4938), .ZN(n17276) );
  NAND2_X1 U1018 ( .A1(n16575), .A2(n16576), .ZN(n17132) );
  BUF_X1 U479 ( .A(n16561), .Z(n17615) );
  BUF_X1 U21220 ( .A(n17061), .Z(n24398) );
  INV_X1 U5527 ( .A(n16963), .ZN(n1612) );
  AND2_X1 U73 ( .A1(n5167), .A2(n15936), .ZN(n372) );
  AND2_X1 U913 ( .A1(n17159), .A2(n17157), .ZN(n17164) );
  NOR2_X1 U5526 ( .A1(n1612), .A2(n17438), .ZN(n16830) );
  OAI22_X1 U7156 ( .A1(n16430), .A2(n1612), .B1(n17128), .B2(n17445), .ZN(
        n18589) );
  AND2_X1 U2828 ( .A1(n492), .A2(n491), .ZN(n18397) );
  NAND3_X1 U482 ( .A1(n2055), .A2(n5707), .A3(n2054), .ZN(n18466) );
  NAND2_X1 U24079 ( .A1(n17004), .A2(n2614), .ZN(n18695) );
  NAND2_X1 U234 ( .A1(n16614), .A2(n16613), .ZN(n18220) );
  AOI21_X1 U19778 ( .B1(n17544), .B2(n17543), .A(n17542), .ZN(n18472) );
  AND4_X1 U1996 ( .A1(n2510), .A2(n17281), .A3(n17282), .A4(n17280), .ZN(
        n17520) );
  OR2_X1 U19532 ( .A1(n17083), .A2(n17082), .ZN(n18483) );
  XNOR2_X1 U1976 ( .A(n2041), .B(n18585), .ZN(n19420) );
  XNOR2_X1 U695 ( .A(n15735), .B(n15736), .ZN(n19307) );
  XNOR2_X1 U1971 ( .A(n18316), .B(n18315), .ZN(n19565) );
  XNOR2_X1 U9356 ( .A(n16092), .B(n16093), .ZN(n19304) );
  XNOR2_X1 U1965 ( .A(n18224), .B(n18223), .ZN(n19185) );
  INV_X1 U11239 ( .A(n19365), .ZN(n19371) );
  CLKBUF_X1 U35 ( .A(n18830), .Z(n19602) );
  BUF_X1 U23995 ( .A(n2540), .Z(n24447) );
  AOI22_X1 U4319 ( .A1(n19206), .A2(n19379), .B1(n19205), .B2(n19204), .ZN(
        n20192) );
  OAI211_X1 U7838 ( .C1(n19563), .C2(n19564), .A(n19562), .B(n19561), .ZN(
        n20367) );
  NAND4_X1 U20480 ( .A1(n18498), .A2(n18497), .A3(n18496), .A4(n18495), .ZN(
        n20571) );
  INV_X1 U11269 ( .A(n20470), .ZN(n5115) );
  NAND4_X1 U11207 ( .A1(n18893), .A2(n18890), .A3(n18892), .A4(n18891), .ZN(
        n20549) );
  OR2_X1 U21066 ( .A1(n19542), .A2(n19541), .ZN(n19544) );
  AOI21_X1 U5610 ( .B1(n4289), .B2(n18933), .A(n4288), .ZN(n19155) );
  NAND2_X1 U1023 ( .A1(n19008), .A2(n4425), .ZN(n20149) );
  INV_X1 U20909 ( .A(n19155), .ZN(n20101) );
  AND3_X1 U1394 ( .A1(n19062), .A2(n1132), .A3(n1131), .ZN(n20498) );
  NAND2_X1 U1866 ( .A1(n19040), .A2(n5234), .ZN(n20301) );
  NAND2_X1 U8900 ( .A1(n24217), .A2(n17941), .ZN(n1591) );
  AND3_X1 U17232 ( .A1(n19506), .A2(n19505), .A3(n19504), .ZN(n19777) );
  OR2_X1 U5651 ( .A1(n20546), .A2(n20125), .ZN(n19675) );
  AND3_X1 U664 ( .A1(n18802), .A2(n18803), .A3(n18801), .ZN(n21212) );
  AND3_X1 U21360 ( .A1(n19931), .A2(n19930), .A3(n19929), .ZN(n20999) );
  NOR3_X1 U21246 ( .A1(n351), .A2(n19799), .A3(n19798), .ZN(n19800) );
  AND3_X1 U21685 ( .A1(n20542), .A2(n20541), .A3(n20540), .ZN(n21422) );
  OAI21_X1 U12080 ( .B1(n20548), .B2(n19677), .A(n19676), .ZN(n21436) );
  OAI21_X1 U4331 ( .B1(n20131), .B2(n3833), .A(n3831), .ZN(n21550) );
  NAND2_X1 U7110 ( .A1(n1995), .A2(n20201), .ZN(n21445) );
  NAND2_X1 U1812 ( .A1(n19961), .A2(n19960), .ZN(n20948) );
  OAI211_X1 U21618 ( .C1(n20398), .C2(n350), .A(n20397), .B(n20396), .ZN(
        n21965) );
  OAI211_X1 U11735 ( .C1(n20549), .C2(n20548), .A(n5638), .B(n5637), .ZN(
        n21158) );
  NAND2_X1 U3336 ( .A1(n742), .A2(n19822), .ZN(n21319) );
  NAND2_X1 U2999 ( .A1(n2104), .A2(n587), .ZN(n21301) );
  NAND3_X1 U1801 ( .A1(n20144), .A2(n5444), .A3(n5443), .ZN(n21554) );
  NOR2_X1 U1271 ( .A1(n20053), .A2(n20052), .ZN(n21704) );
  XNOR2_X1 U598 ( .A(n21546), .B(n21545), .ZN(n22421) );
  XNOR2_X1 U1778 ( .A(n21187), .B(n21186), .ZN(n22592) );
  BUF_X1 U21103 ( .A(n23575), .Z(n24396) );
  XNOR2_X1 U1263 ( .A(n21485), .B(n21484), .ZN(n22968) );
  XNOR2_X1 U738 ( .A(n21131), .B(n21130), .ZN(n22675) );
  BUF_X1 U584 ( .A(n21888), .Z(n22401) );
  OR2_X1 U3384 ( .A1(n772), .A2(n4371), .ZN(n23265) );
  AOI21_X1 U45 ( .B1(n21936), .B2(n21937), .A(n22562), .ZN(n22571) );
  NOR2_X1 U23016 ( .A1(n22238), .A2(n22237), .ZN(n23730) );
  AND2_X1 U1036 ( .A1(n1587), .A2(n1585), .ZN(n23273) );
  NAND2_X1 U20246 ( .A1(n22213), .A2(n2314), .ZN(n23743) );
  AND2_X1 U912 ( .A1(n21113), .A2(n2595), .ZN(n23074) );
  AND3_X1 U8694 ( .A1(n2901), .A2(n3024), .A3(n3309), .ZN(n23303) );
  OR2_X1 U243 ( .A1(n22045), .A2(n22046), .ZN(n22043) );
  NAND3_X1 U1721 ( .A1(n4283), .A2(n1417), .A3(n4282), .ZN(n23906) );
  CLKBUF_X1 U1567 ( .A(Key[25]), .Z(n21423) );
  CLKBUF_X1 U1608 ( .A(Key[189]), .Z(n21553) );
  XNOR2_X1 U12393 ( .A(n5950), .B(Key[170]), .ZN(n6489) );
  NAND2_X1 U2644 ( .A1(n4756), .A2(n5906), .ZN(n8511) );
  AOI21_X1 U5258 ( .B1(n7143), .B2(n7142), .A(n2780), .ZN(n8168) );
  AOI22_X1 U12832 ( .A1(n6864), .A2(n6466), .B1(n7216), .B2(n6465), .ZN(n9147)
         );
  NOR2_X1 U11965 ( .A1(n24944), .A2(n9463), .ZN(n9351) );
  OAI211_X1 U2456 ( .C1(n10146), .C2(n10145), .A(n10144), .B(n10143), .ZN(
        n10654) );
  NAND4_X1 U3368 ( .A1(n9030), .A2(n9031), .A3(n9029), .A4(n9032), .ZN(n11039)
         );
  BUF_X1 U1197 ( .A(n10192), .Z(n10829) );
  BUF_X1 U1239 ( .A(n11518), .Z(n11525) );
  NAND2_X1 U2377 ( .A1(n11202), .A2(n3011), .ZN(n12023) );
  XNOR2_X1 U1495 ( .A(n12348), .B(n12347), .ZN(n13124) );
  OAI211_X1 U2258 ( .C1(n13065), .C2(n5112), .A(n3710), .B(n2859), .ZN(n13974)
         );
  INV_X1 U1456 ( .A(n16008), .ZN(n3554) );
  BUF_X1 U1261 ( .A(n16428), .Z(n244) );
  INV_X1 U1467 ( .A(n15706), .ZN(n294) );
  INV_X1 U2079 ( .A(n16516), .ZN(n17138) );
  NAND2_X1 U7825 ( .A1(n16020), .A2(n2344), .ZN(n16991) );
  OR2_X1 U2039 ( .A1(n25200), .A2(n17208), .ZN(n17017) );
  MUX2_X1 U9019 ( .A(n17318), .B(n17317), .S(n17316), .Z(n18448) );
  XNOR2_X1 U591 ( .A(n17957), .B(n17956), .ZN(n19380) );
  AOI22_X1 U3972 ( .A1(n19249), .A2(n19248), .B1(n3620), .B2(n1098), .ZN(
        n20426) );
  CLKBUF_X1 U1846 ( .A(n19494), .Z(n20239) );
  INV_X1 U4791 ( .A(n23996), .ZN(n22677) );
  INV_X1 U4780 ( .A(n23014), .ZN(n23461) );
  AND3_X2 U207 ( .A1(n3140), .A2(n20067), .A3(n19158), .ZN(n21689) );
  BUF_X1 U24128 ( .A(n23275), .Z(n24486) );
  NAND4_X2 U7546 ( .A1(n2169), .A2(n19746), .A3(n19747), .A4(n1452), .ZN(
        n21622) );
  OR2_X2 U7505 ( .A1(n4123), .A2(n2153), .ZN(n14221) );
  OR2_X2 U1096 ( .A1(n16318), .A2(n16317), .ZN(n18646) );
  OAI21_X2 U608 ( .B1(n1409), .B2(n2890), .A(n5384), .ZN(n18429) );
  NAND2_X2 U19060 ( .A1(n16297), .A2(n16296), .ZN(n17356) );
  AND2_X2 U1692 ( .A1(n21920), .A2(n211), .ZN(n23196) );
  NAND3_X2 U3442 ( .A1(n4974), .A2(n16958), .A3(n4502), .ZN(n18675) );
  BUF_X2 U6860 ( .A(n9345), .Z(n9927) );
  XNOR2_X2 U653 ( .A(n7837), .B(n7836), .ZN(n9603) );
  AND2_X2 U1196 ( .A1(n2392), .A2(n2390), .ZN(n10302) );
  NOR2_X2 U586 ( .A1(n5340), .A2(n10256), .ZN(n10734) );
  AND2_X2 U833 ( .A1(n4798), .A2(n4797), .ZN(n14319) );
  XNOR2_X2 U9496 ( .A(n17697), .B(n17696), .ZN(n19445) );
  AND2_X2 U1007 ( .A1(n4638), .A2(n4618), .ZN(n13792) );
  AND3_X2 U11342 ( .A1(n5185), .A2(n5186), .A3(n19829), .ZN(n21738) );
  AND2_X2 U1046 ( .A1(n16682), .A2(n16680), .ZN(n17277) );
  OAI21_X2 U176 ( .B1(n3818), .B2(n16606), .A(n16605), .ZN(n18694) );
  OR2_X2 U713 ( .A1(n4501), .A2(n4500), .ZN(n12147) );
  BUF_X2 U6328 ( .A(n18982), .Z(n20014) );
  AND3_X2 U24197 ( .A1(n1913), .A2(n963), .A3(n1911), .ZN(n17293) );
  AND2_X2 U8787 ( .A1(n15698), .A2(n16549), .ZN(n2587) );
  AND2_X2 U502 ( .A1(n4255), .A2(n4253), .ZN(n11058) );
  MUX2_X2 U19344 ( .A(n16793), .B(n16792), .S(n1516), .Z(n18602) );
  INV_X2 U401 ( .A(n11084), .ZN(n3119) );
  NOR2_X2 U14582 ( .A1(n3337), .A2(n12639), .ZN(n14198) );
  NAND2_X2 U1029 ( .A1(n17036), .A2(n18925), .ZN(n20336) );
  OAI21_X2 U930 ( .B1(n20334), .B2(n20333), .A(n20332), .ZN(n22005) );
  BUF_X2 U980 ( .A(n15986), .Z(n16141) );
  OAI211_X2 U345 ( .C1(n8332), .C2(n10169), .A(n4212), .B(n2548), .ZN(n10596)
         );
  NAND2_X2 U246 ( .A1(n21), .A2(n20), .ZN(n13829) );
  OR2_X2 U10252 ( .A1(n4089), .A2(n10636), .ZN(n12167) );
  AND3_X2 U1129 ( .A1(n867), .A2(n1857), .A3(n1858), .ZN(n11045) );
  NOR2_X2 U2974 ( .A1(n575), .A2(n16580), .ZN(n17881) );
  BUF_X2 U1280 ( .A(n6849), .Z(n250) );
  NAND4_X2 U9456 ( .A1(n3318), .A2(n3319), .A3(n15744), .A4(n16198), .ZN(
        n17391) );
  NAND2_X2 U570 ( .A1(n10231), .A2(n10230), .ZN(n11704) );
  NOR2_X2 U691 ( .A1(n14951), .A2(n14950), .ZN(n15494) );
  OR2_X2 U536 ( .A1(n5382), .A2(n5381), .ZN(n12357) );
  NAND2_X2 U1686 ( .A1(n4944), .A2(n4943), .ZN(n14267) );
  XNOR2_X2 U1164 ( .A(n15400), .B(n15399), .ZN(n15694) );
  AND3_X2 U1277 ( .A1(n12997), .A2(n12999), .A3(n12998), .ZN(n14219) );
  BUF_X2 U643 ( .A(n18719), .Z(n19497) );
  BUF_X1 U2502 ( .A(n7183), .Z(n9949) );
  AND2_X2 U2666 ( .A1(n6485), .A2(n6484), .ZN(n7638) );
  XNOR2_X2 U511 ( .A(n8390), .B(n8389), .ZN(n10161) );
  BUF_X1 U2407 ( .A(n9769), .Z(n10364) );
  NOR2_X2 U963 ( .A1(n16421), .A2(n16420), .ZN(n17445) );
  AND3_X1 U2304 ( .A1(n2737), .A2(n5086), .A3(n2736), .ZN(n1985) );
  BUF_X1 U4580 ( .A(n9134), .Z(n9953) );
  NOR2_X1 U6054 ( .A1(n9461), .A2(n9459), .ZN(n1470) );
  AND2_X1 U4438 ( .A1(n9786), .A2(n10082), .ZN(n9789) );
  AOI21_X1 U2386 ( .B1(n10236), .B2(n10237), .A(n10235), .ZN(n11076) );
  OAI211_X1 U717 ( .C1(n9444), .C2(n9443), .A(n9442), .B(n9441), .ZN(n12275)
         );
  BUF_X1 U2305 ( .A(n12625), .Z(n12878) );
  NAND3_X1 U323 ( .A1(n13557), .A2(n13556), .A3(n13555), .ZN(n15444) );
  XNOR2_X1 U762 ( .A(n14531), .B(n14530), .ZN(n16394) );
  BUF_X2 U595 ( .A(n16765), .Z(n17574) );
  OR3_X1 U21239 ( .A1(n20244), .A2(n20241), .A3(n19937), .ZN(n19789) );
  OAI21_X2 U994 ( .B1(n20666), .B2(n19712), .A(n19711), .ZN(n21745) );
  OAI21_X2 U3876 ( .B1(n20481), .B2(n20480), .A(n1022), .ZN(n21040) );
  BUF_X1 U1754 ( .A(n21540), .Z(n22422) );
  OAI21_X1 U1 ( .B1(n21374), .B2(n21373), .A(n21372), .ZN(n24473) );
  NAND2_X1 U2 ( .A1(n1074), .A2(n21890), .ZN(n23311) );
  BUF_X1 U4 ( .A(n22128), .Z(n22966) );
  BUF_X2 U7 ( .A(n19953), .Z(n20591) );
  NOR2_X1 U13 ( .A1(n1014), .A2(n1010), .ZN(n20338) );
  XNOR2_X1 U27 ( .A(n1387), .B(n18556), .ZN(n19084) );
  MUX2_X1 U32 ( .A(n15261), .B(n15260), .S(n24330), .Z(n18074) );
  NAND3_X1 U34 ( .A1(n14030), .A2(n14029), .A3(n76), .ZN(n15506) );
  NAND4_X1 U37 ( .A1(n2302), .A2(n2303), .A3(n2301), .A4(n13723), .ZN(n15452)
         );
  NOR2_X1 U43 ( .A1(n13625), .A2(n13624), .ZN(n14678) );
  NOR2_X1 U48 ( .A1(n8663), .A2(n8662), .ZN(n25016) );
  XNOR2_X2 U82 ( .A(n21643), .B(n21642), .ZN(n22939) );
  OR2_X2 U105 ( .A1(n17451), .A2(n17455), .ZN(n3982) );
  BUF_X2 U122 ( .A(n16284), .Z(n24540) );
  AND3_X2 U134 ( .A1(n24647), .A2(n24646), .A3(n19357), .ZN(n17714) );
  AND3_X2 U143 ( .A1(n24767), .A2(n9663), .A3(n1943), .ZN(n10630) );
  BUF_X2 U155 ( .A(n9992), .Z(n24534) );
  BUF_X1 U169 ( .A(n15922), .Z(n16464) );
  OR2_X2 U175 ( .A1(n7569), .A2(n2026), .ZN(n9191) );
  AND2_X2 U184 ( .A1(n2117), .A2(n2116), .ZN(n24974) );
  AND2_X2 U186 ( .A1(n4706), .A2(n4708), .ZN(n8352) );
  BUF_X1 U222 ( .A(n12226), .Z(n24915) );
  AND3_X2 U250 ( .A1(n4886), .A2(n1202), .A3(n4887), .ZN(n4004) );
  NAND3_X2 U273 ( .A1(n24697), .A2(n1400), .A3(n4014), .ZN(n2242) );
  OR2_X2 U275 ( .A1(n18754), .A2(n18753), .ZN(n19809) );
  INV_X1 U290 ( .A(n19166), .ZN(n24584) );
  OAI21_X1 U292 ( .B1(n20405), .B2(n20419), .A(n20404), .ZN(n20585) );
  INV_X1 U293 ( .A(n22953), .ZN(n22959) );
  XNOR2_X2 U310 ( .A(n8048), .B(n8047), .ZN(n9864) );
  OAI211_X2 U318 ( .C1(n12538), .C2(n1636), .A(n1634), .B(n1633), .ZN(n14268)
         );
  OR2_X2 U320 ( .A1(n24259), .A2(n13516), .ZN(n15476) );
  XOR2_X1 U341 ( .A(n14693), .B(n14692), .Z(n24532) );
  NOR2_X2 U349 ( .A1(n16234), .A2(n1096), .ZN(n17216) );
  NOR2_X2 U351 ( .A1(n16944), .A2(n17611), .ZN(n18677) );
  NAND3_X1 U355 ( .A1(n20497), .A2(n24887), .A3(n20496), .ZN(n24533) );
  NOR2_X2 U367 ( .A1(n21827), .A2(n3890), .ZN(n21837) );
  BUF_X2 U370 ( .A(n19041), .Z(n19361) );
  INV_X2 U372 ( .A(n5692), .ZN(n15375) );
  CLKBUF_X1 U379 ( .A(n9992), .Z(n24535) );
  XNOR2_X1 U387 ( .A(n8894), .B(n8895), .ZN(n9992) );
  XNOR2_X2 U410 ( .A(n8284), .B(n8283), .ZN(n10113) );
  XNOR2_X2 U437 ( .A(n8166), .B(n8165), .ZN(n9564) );
  OR2_X2 U450 ( .A1(n16071), .A2(n16070), .ZN(n17165) );
  NAND2_X2 U454 ( .A1(n20088), .A2(n20087), .ZN(n21676) );
  BUF_X1 U457 ( .A(n9127), .Z(n10062) );
  CLKBUF_X1 U467 ( .A(n16393), .Z(n24537) );
  XNOR2_X1 U476 ( .A(n14536), .B(n14535), .ZN(n16393) );
  XNOR2_X1 U498 ( .A(n15050), .B(n15049), .ZN(n16284) );
  NAND3_X2 U501 ( .A1(n4642), .A2(n6382), .A3(n4641), .ZN(n8370) );
  BUF_X1 U509 ( .A(n17313), .Z(n24542) );
  OAI211_X1 U517 ( .C1(n15660), .C2(n15659), .A(n5502), .B(n15658), .ZN(n17313) );
  XNOR2_X1 U540 ( .A(n20314), .B(n20315), .ZN(n22809) );
  OAI211_X2 U544 ( .C1(n20240), .C2(n20239), .A(n20238), .B(n4750), .ZN(n21070) );
  OAI211_X2 U554 ( .C1(n19861), .C2(n19860), .A(n19859), .B(n19858), .ZN(
        n21136) );
  XNOR2_X2 U557 ( .A(n18048), .B(n18049), .ZN(n19596) );
  XNOR2_X2 U558 ( .A(n4583), .B(n4581), .ZN(n16334) );
  BUF_X2 U562 ( .A(n19878), .Z(n20555) );
  AND2_X2 U583 ( .A1(n5308), .A2(n5307), .ZN(n16037) );
  AND2_X2 U590 ( .A1(n5271), .A2(n5274), .ZN(n11201) );
  NAND2_X2 U615 ( .A1(n3226), .A2(n3228), .ZN(n23805) );
  XNOR2_X2 U621 ( .A(n14784), .B(n14783), .ZN(n16246) );
  AND3_X2 U623 ( .A1(n2144), .A2(n4817), .A3(n4818), .ZN(n17816) );
  XNOR2_X1 U626 ( .A(n8092), .B(n8091), .ZN(n9874) );
  OAI21_X2 U627 ( .B1(n16370), .B2(n17460), .A(n16369), .ZN(n18610) );
  BUF_X1 U629 ( .A(n16470), .Z(n24551) );
  XNOR2_X1 U636 ( .A(n15450), .B(n15449), .ZN(n16470) );
  MUX2_X2 U638 ( .A(n12790), .B(n12789), .S(n13027), .Z(n13864) );
  OAI211_X2 U642 ( .C1(n19996), .C2(n19995), .A(n19994), .B(n19993), .ZN(
        n20914) );
  AND4_X2 U657 ( .A1(n2687), .A2(n19773), .A3(n19772), .A4(n2685), .ZN(n21608)
         );
  XNOR2_X1 U673 ( .A(n2415), .B(n2416), .ZN(n21829) );
  OAI21_X2 U678 ( .B1(n18829), .B2(n19087), .A(n4194), .ZN(n20353) );
  NOR2_X2 U681 ( .A1(n19808), .A2(n19807), .ZN(n20982) );
  XNOR2_X2 U682 ( .A(n8338), .B(n8337), .ZN(n9837) );
  AND2_X2 U683 ( .A1(n972), .A2(n971), .ZN(n23810) );
  XNOR2_X2 U686 ( .A(n14661), .B(n14660), .ZN(n16076) );
  BUF_X1 U741 ( .A(n13360), .Z(n24554) );
  XNOR2_X1 U766 ( .A(n12126), .B(n12125), .ZN(n13360) );
  NAND2_X2 U780 ( .A1(n1751), .A2(n9202), .ZN(n10584) );
  NOR2_X2 U783 ( .A1(n10653), .A2(n10652), .ZN(n12146) );
  XNOR2_X2 U794 ( .A(n8196), .B(n8195), .ZN(n10148) );
  OAI211_X2 U808 ( .C1(n20582), .C2(n20583), .A(n20581), .B(n20580), .ZN(
        n21053) );
  NOR2_X2 U816 ( .A1(n3800), .A2(n9667), .ZN(n10789) );
  NOR2_X1 U840 ( .A1(n12723), .A2(n12722), .ZN(n14435) );
  AOI22_X2 U872 ( .A1(n4713), .A2(n20349), .B1(n20351), .B2(n20350), .ZN(
        n21058) );
  XNOR2_X2 U901 ( .A(n11988), .B(n11989), .ZN(n13267) );
  NOR2_X2 U902 ( .A1(n1866), .A2(n12779), .ZN(n14669) );
  XNOR2_X2 U905 ( .A(n8642), .B(n8641), .ZN(n10104) );
  AND3_X2 U911 ( .A1(n9835), .A2(n9833), .A3(n9834), .ZN(n10548) );
  NOR2_X2 U922 ( .A1(n15903), .A2(n15902), .ZN(n17039) );
  OAI22_X2 U923 ( .A1(n990), .A2(n14017), .B1(n13534), .B2(n13607), .ZN(n15033) );
  XNOR2_X2 U926 ( .A(n21443), .B(n21442), .ZN(n22965) );
  XNOR2_X2 U941 ( .A(n20495), .B(n20494), .ZN(n21856) );
  CLKBUF_X1 U955 ( .A(n24510), .Z(n24561) );
  XNOR2_X1 U956 ( .A(n21218), .B(n21219), .ZN(n24510) );
  XNOR2_X2 U957 ( .A(n15346), .B(n15345), .ZN(n15953) );
  AND2_X2 U962 ( .A1(n1947), .A2(n1946), .ZN(n16795) );
  XNOR2_X2 U966 ( .A(n11850), .B(n1384), .ZN(n12899) );
  AOI21_X2 U1038 ( .B1(n16180), .B2(n16179), .A(n16178), .ZN(n17400) );
  NAND2_X2 U1060 ( .A1(n5092), .A2(n5091), .ZN(n21505) );
  INV_X1 U1065 ( .A(n12902), .ZN(n4499) );
  NOR2_X1 U1089 ( .A1(n17556), .A2(n4436), .ZN(n19263) );
  OAI211_X2 U1092 ( .C1(n7602), .C2(n7603), .A(n3007), .B(n3006), .ZN(n8446)
         );
  NOR2_X2 U1093 ( .A1(n16593), .A2(n24699), .ZN(n18685) );
  NOR2_X2 U1095 ( .A1(n17448), .A2(n17447), .ZN(n18456) );
  OAI211_X2 U1102 ( .C1(n2638), .C2(n2636), .A(n2637), .B(n2635), .ZN(n5376)
         );
  NOR2_X1 U1103 ( .A1(n13112), .A2(n13110), .ZN(n12853) );
  AND2_X1 U1159 ( .A1(n20941), .A2(n20942), .ZN(n23612) );
  INV_X1 U1161 ( .A(n20670), .ZN(n24567) );
  INV_X1 U1167 ( .A(n17364), .ZN(n24569) );
  INV_X1 U1171 ( .A(n17051), .ZN(n24570) );
  OR2_X1 U1181 ( .A1(n16902), .A2(n2562), .ZN(n45) );
  XNOR2_X1 U1187 ( .A(n14552), .B(n14551), .ZN(n15849) );
  INV_X1 U1194 ( .A(n14435), .ZN(n24571) );
  XNOR2_X1 U1201 ( .A(n11882), .B(n11883), .ZN(n4241) );
  BUF_X2 U1204 ( .A(n13077), .Z(n24573) );
  INV_X1 U1213 ( .A(n11112), .ZN(n24574) );
  OR2_X1 U1217 ( .A1(n262), .A2(n9281), .ZN(n25174) );
  OAI211_X1 U1224 ( .C1(n7152), .C2(n7217), .A(n7150), .B(n7149), .ZN(n8627)
         );
  INV_X1 U1226 ( .A(n7864), .ZN(n24576) );
  NAND3_X1 U1228 ( .A1(n25184), .A2(n6501), .A3(n6502), .ZN(n8527) );
  INV_X1 U1231 ( .A(n7734), .ZN(n24578) );
  CLKBUF_X1 U1242 ( .A(Key[113]), .Z(n2036) );
  CLKBUF_X1 U1258 ( .A(Key[166]), .Z(n62) );
  INV_X1 U1265 ( .A(n6975), .ZN(n24579) );
  CLKBUF_X1 U1267 ( .A(Key[107]), .Z(n2228) );
  OR2_X1 U1268 ( .A1(n23483), .A2(n23499), .ZN(n24874) );
  OR2_X1 U1270 ( .A1(n23979), .A2(n24440), .ZN(n24873) );
  OR2_X1 U1282 ( .A1(n23030), .A2(n22539), .ZN(n21352) );
  AND2_X1 U1286 ( .A1(n23052), .A2(n23047), .ZN(n23039) );
  INV_X1 U1288 ( .A(n23219), .ZN(n23231) );
  CLKBUF_X1 U1290 ( .A(n23799), .Z(n24920) );
  AOI21_X1 U1291 ( .B1(n25050), .B2(n22165), .A(n22164), .ZN(n25026) );
  OR2_X1 U1293 ( .A1(n23297), .A2(n22395), .ZN(n22510) );
  INV_X1 U1298 ( .A(n1075), .ZN(n23320) );
  OR2_X1 U1299 ( .A1(n23817), .A2(n891), .ZN(n21355) );
  AND3_X1 U1317 ( .A1(n1068), .A2(n1905), .A3(n1065), .ZN(n23420) );
  OR2_X1 U1361 ( .A1(n21894), .A2(n1076), .ZN(n1075) );
  AND2_X1 U1366 ( .A1(n25138), .A2(n2038), .ZN(n23129) );
  AOI21_X1 U1367 ( .B1(n21927), .B2(n21926), .A(n21925), .ZN(n24889) );
  MUX2_X1 U1369 ( .A(n22038), .B(n22037), .S(n603), .Z(n24880) );
  MUX2_X1 U1374 ( .A(n22372), .B(n22371), .S(n22680), .Z(n24948) );
  NOR2_X1 U1376 ( .A1(n21923), .A2(n21922), .ZN(n21927) );
  AND2_X1 U1381 ( .A1(n24673), .A2(n24672), .ZN(n22074) );
  OAI211_X1 U1385 ( .C1(n4098), .C2(n3213), .A(n22977), .B(n24724), .ZN(n2901)
         );
  INV_X1 U1391 ( .A(n22282), .ZN(n24631) );
  INV_X1 U1399 ( .A(n22677), .ZN(n24869) );
  XNOR2_X1 U1400 ( .A(n21203), .B(n21202), .ZN(n22798) );
  XNOR2_X1 U1402 ( .A(n20575), .B(n20574), .ZN(n22679) );
  XNOR2_X1 U1413 ( .A(n20802), .B(n20801), .ZN(n22459) );
  BUF_X2 U1415 ( .A(n21665), .Z(n24898) );
  NAND3_X1 U1421 ( .A1(n24138), .A2(n5123), .A3(n19920), .ZN(n21647) );
  AND2_X1 U1436 ( .A1(n3903), .A2(n25028), .ZN(n21273) );
  OR2_X1 U1512 ( .A1(n19674), .A2(n20124), .ZN(n5262) );
  NOR2_X1 U1520 ( .A1(n19849), .A2(n19658), .ZN(n19659) );
  NOR2_X1 U1522 ( .A1(n20224), .A2(n20498), .ZN(n24682) );
  NAND2_X1 U1547 ( .A1(n24733), .A2(n18905), .ZN(n20546) );
  AND2_X1 U1554 ( .A1(n100), .A2(n20507), .ZN(n24644) );
  AND2_X1 U1561 ( .A1(n20557), .A2(n3480), .ZN(n24749) );
  INV_X1 U1614 ( .A(n20523), .ZN(n20131) );
  OR2_X1 U1681 ( .A1(n19889), .A2(n20319), .ZN(n2180) );
  INV_X1 U1689 ( .A(n20290), .ZN(n24581) );
  OAI21_X1 U1691 ( .B1(n24638), .B2(n19028), .A(n24637), .ZN(n4067) );
  NAND2_X1 U1700 ( .A1(n3508), .A2(n18879), .ZN(n20523) );
  OR2_X1 U1709 ( .A1(n20169), .A2(n20173), .ZN(n19958) );
  INV_X1 U1712 ( .A(n25034), .ZN(n24829) );
  OR2_X1 U1727 ( .A1(n18787), .A2(n18786), .ZN(n20473) );
  AND2_X1 U1743 ( .A1(n25158), .A2(n25157), .ZN(n20510) );
  AND3_X1 U1748 ( .A1(n17803), .A2(n17802), .A3(n17801), .ZN(n20111) );
  AND2_X1 U1762 ( .A1(n18976), .A2(n19460), .ZN(n24638) );
  NAND3_X1 U1763 ( .A1(n25105), .A2(n2304), .A3(n18716), .ZN(n20042) );
  INV_X1 U1765 ( .A(n24172), .ZN(n24637) );
  INV_X1 U1768 ( .A(n19037), .ZN(n24582) );
  INV_X1 U1789 ( .A(n25002), .ZN(n24809) );
  OR2_X1 U1807 ( .A1(n19548), .A2(n24929), .ZN(n24717) );
  INV_X1 U1817 ( .A(n16737), .ZN(n24719) );
  INV_X1 U1862 ( .A(n17497), .ZN(n24583) );
  XNOR2_X1 U1863 ( .A(n18555), .B(n24769), .ZN(n1387) );
  NAND2_X1 U1875 ( .A1(n2829), .A2(n24615), .ZN(n18523) );
  MUX2_X1 U1885 ( .A(n17301), .B(n17300), .S(n17299), .Z(n17303) );
  AND2_X1 U1914 ( .A1(n17141), .A2(n1653), .ZN(n24688) );
  NOR2_X1 U1927 ( .A1(n16255), .A2(n16256), .ZN(n17016) );
  AND2_X1 U1930 ( .A1(n17293), .A2(n17283), .ZN(n24775) );
  INV_X1 U1937 ( .A(n17249), .ZN(n17252) );
  INV_X1 U1952 ( .A(n17081), .ZN(n16895) );
  OAI21_X1 U1967 ( .B1(n16280), .B2(n25180), .A(n16278), .ZN(n17352) );
  OR2_X1 U1970 ( .A1(n15931), .A2(n16450), .ZN(n25116) );
  NAND2_X1 U1986 ( .A1(n16364), .A2(n16363), .ZN(n523) );
  OAI21_X1 U1997 ( .B1(n16293), .B2(n24842), .A(n24841), .ZN(n16297) );
  AND2_X1 U2019 ( .A1(n257), .A2(n16447), .ZN(n24774) );
  XOR2_X1 U2036 ( .A(n15092), .B(n15091), .Z(n24919) );
  INV_X1 U2037 ( .A(n15782), .ZN(n24586) );
  INV_X1 U2045 ( .A(n15821), .ZN(n24587) );
  MUX2_X2 U2053 ( .A(n14184), .B(n14183), .S(n14182), .Z(n14642) );
  OAI21_X1 U2055 ( .B1(n13721), .B2(n13720), .A(n13719), .ZN(n15253) );
  XNOR2_X1 U2063 ( .A(n14703), .B(n14553), .ZN(n15392) );
  NAND2_X1 U2077 ( .A1(n13698), .A2(n2741), .ZN(n14690) );
  NAND3_X1 U2123 ( .A1(n13919), .A2(n13920), .A3(n760), .ZN(n15350) );
  NAND3_X1 U2155 ( .A1(n24776), .A2(n2151), .A3(n2150), .ZN(n15054) );
  OR2_X1 U2187 ( .A1(n13675), .A2(n13674), .ZN(n24691) );
  INV_X1 U2197 ( .A(n13888), .ZN(n24710) );
  BUF_X1 U2201 ( .A(n12850), .Z(n14335) );
  AND3_X1 U2202 ( .A1(n2906), .A2(n24094), .A3(n2905), .ZN(n13839) );
  AND3_X1 U2212 ( .A1(n5724), .A2(n12762), .A3(n5723), .ZN(n24949) );
  INV_X1 U2220 ( .A(n14059), .ZN(n24785) );
  NAND2_X1 U2233 ( .A1(n498), .A2(n24854), .ZN(n14158) );
  OR3_X1 U2257 ( .A1(n11319), .A2(n13230), .A3(n25080), .ZN(n11331) );
  INV_X1 U2319 ( .A(n14166), .ZN(n24773) );
  INV_X1 U2331 ( .A(n3876), .ZN(n24617) );
  AND2_X1 U2364 ( .A1(n13282), .A2(n24988), .ZN(n12931) );
  XNOR2_X1 U2373 ( .A(n12115), .B(n12116), .ZN(n12956) );
  INV_X1 U2423 ( .A(n11689), .ZN(n24778) );
  NAND3_X1 U2442 ( .A1(n24761), .A2(n9343), .A3(n24760), .ZN(n25090) );
  OR2_X1 U2486 ( .A1(n10725), .A2(n11116), .ZN(n24760) );
  INV_X1 U2508 ( .A(n10914), .ZN(n24753) );
  OAI21_X1 U2529 ( .B1(n10285), .B2(n10875), .A(n11117), .ZN(n24761) );
  OR2_X1 U2533 ( .A1(n11066), .A2(n11068), .ZN(n25103) );
  NOR2_X1 U2544 ( .A1(n11518), .A2(n11519), .ZN(n10918) );
  OR2_X1 U2552 ( .A1(n10753), .A2(n10451), .ZN(n25156) );
  INV_X1 U2568 ( .A(n11171), .ZN(n24591) );
  NAND4_X1 U2573 ( .A1(n8575), .A2(n8572), .A3(n8574), .A4(n8573), .ZN(n24957)
         );
  NAND2_X1 U2630 ( .A1(n9819), .A2(n655), .ZN(n10951) );
  NOR2_X1 U2634 ( .A1(n9624), .A2(n3674), .ZN(n4871) );
  OR2_X1 U2699 ( .A1(n7670), .A2(n7671), .ZN(n25152) );
  OR2_X1 U2716 ( .A1(n7596), .A2(n24772), .ZN(n3007) );
  INV_X1 U2720 ( .A(n7688), .ZN(n7148) );
  AND3_X1 U2771 ( .A1(n25186), .A2(n6453), .A3(n6452), .ZN(n7691) );
  OR2_X1 U2776 ( .A1(n873), .A2(n6361), .ZN(n24878) );
  BUF_X1 U2792 ( .A(n6577), .Z(n6752) );
  CLKBUF_X1 U2798 ( .A(Key[106]), .Z(n173) );
  OR2_X1 U2808 ( .A1(n6504), .A2(n6503), .ZN(n25184) );
  AND3_X1 U2819 ( .A1(n5001), .A2(n5002), .A3(n6734), .ZN(n6868) );
  OR2_X1 U2825 ( .A1(n6335), .A2(n6332), .ZN(n6440) );
  OR2_X1 U2836 ( .A1(n6244), .A2(n6119), .ZN(n6840) );
  AND2_X1 U2837 ( .A1(n6069), .A2(n6971), .ZN(n24810) );
  INV_X1 U2850 ( .A(n6480), .ZN(n6290) );
  CLKBUF_X1 U2864 ( .A(n6845), .Z(n7027) );
  CLKBUF_X1 U2878 ( .A(n6133), .Z(n6543) );
  INV_X1 U2885 ( .A(n7758), .ZN(n432) );
  OR2_X2 U2888 ( .A1(n6927), .A2(n6928), .ZN(n7947) );
  AND2_X1 U2891 ( .A1(n9066), .A2(n9067), .ZN(n8221) );
  MUX2_X1 U2894 ( .A(n7995), .B(n7994), .S(n7993), .Z(n7996) );
  AOI21_X1 U2911 ( .B1(n24599), .B2(n10169), .A(n9814), .ZN(n25187) );
  OR2_X1 U2928 ( .A1(n7059), .A2(n7809), .ZN(n25117) );
  XNOR2_X1 U2931 ( .A(n8632), .B(n8631), .ZN(n9773) );
  XNOR2_X1 U2934 ( .A(n8331), .B(n8330), .ZN(n10166) );
  INV_X1 U2969 ( .A(n24944), .ZN(n24853) );
  XNOR2_X1 U3011 ( .A(n7571), .B(n7570), .ZN(n1595) );
  BUF_X1 U3018 ( .A(n9859), .Z(n238) );
  OR2_X1 U3026 ( .A1(n9961), .A2(n9468), .ZN(n24804) );
  AOI22_X1 U3040 ( .A1(n9422), .A2(n9421), .B1(n9751), .B2(n9420), .ZN(n9432)
         );
  NOR2_X1 U3055 ( .A1(n24575), .A2(n10082), .ZN(n25163) );
  OR2_X1 U3056 ( .A1(n9362), .A2(n9363), .ZN(n25148) );
  XNOR2_X1 U3065 ( .A(n8002), .B(n8001), .ZN(n9905) );
  OAI21_X1 U3088 ( .B1(n262), .B2(n24927), .A(n24804), .ZN(n1186) );
  OAI21_X1 U3108 ( .B1(n9920), .B2(n24844), .A(n24843), .ZN(n7044) );
  OR2_X1 U3110 ( .A1(n24526), .A2(n10477), .ZN(n24799) );
  OR2_X1 U3124 ( .A1(n10910), .A2(n24753), .ZN(n24817) );
  INV_X1 U3128 ( .A(n12121), .ZN(n25166) );
  OR2_X1 U3136 ( .A1(n10958), .A2(n10703), .ZN(n3244) );
  OR2_X1 U3138 ( .A1(n10428), .A2(n10651), .ZN(n10429) );
  OR2_X1 U3161 ( .A1(n10368), .A2(n10369), .ZN(n25134) );
  XNOR2_X1 U3178 ( .A(n12141), .B(n12114), .ZN(n24634) );
  BUF_X1 U3193 ( .A(n12611), .Z(n12612) );
  OR2_X1 U3198 ( .A1(n13108), .A2(n12674), .ZN(n3829) );
  CLKBUF_X1 U3203 ( .A(n12583), .Z(n13363) );
  XNOR2_X1 U3206 ( .A(n11389), .B(n11956), .ZN(n12786) );
  AOI22_X1 U3214 ( .A1(n12798), .A2(n12476), .B1(n13041), .B2(n13040), .ZN(
        n12763) );
  OR2_X1 U3215 ( .A1(n12793), .A2(n24750), .ZN(n12566) );
  NOR2_X1 U3219 ( .A1(n12744), .A2(n13101), .ZN(n13188) );
  AND2_X1 U3243 ( .A1(n13341), .A2(n12840), .ZN(n12960) );
  NAND3_X1 U3261 ( .A1(n5724), .A2(n12762), .A3(n5723), .ZN(n13795) );
  INV_X1 U3264 ( .A(n231), .ZN(n12958) );
  OR2_X1 U3278 ( .A1(n12879), .A2(n12878), .ZN(n2888) );
  AND2_X1 U3285 ( .A1(n297), .A2(n3717), .ZN(n1027) );
  AND2_X1 U3287 ( .A1(n14079), .A2(n14078), .ZN(n25099) );
  INV_X1 U3293 ( .A(n13636), .ZN(n24679) );
  OR2_X1 U3294 ( .A1(n24745), .A2(n24347), .ZN(n24744) );
  OR2_X1 U3310 ( .A1(n13284), .A2(n25191), .ZN(n12929) );
  AND2_X1 U3311 ( .A1(n14083), .A2(n14073), .ZN(n24815) );
  OR2_X1 U3312 ( .A1(n13515), .A2(n297), .ZN(n3536) );
  OR2_X1 U3322 ( .A1(n14243), .A2(n4116), .ZN(n13639) );
  OR2_X1 U3328 ( .A1(n13896), .A2(n13895), .ZN(n13897) );
  OR2_X1 U3330 ( .A1(n14058), .A2(n12468), .ZN(n24776) );
  XNOR2_X1 U3337 ( .A(n14919), .B(n14865), .ZN(n14331) );
  OR2_X1 U3351 ( .A1(n13944), .A2(n14302), .ZN(n1400) );
  OR2_X1 U3390 ( .A1(n15612), .A2(n15611), .ZN(n15860) );
  INV_X1 U3393 ( .A(n24551), .ZN(n24822) );
  XNOR2_X1 U3395 ( .A(n13836), .B(n13835), .ZN(n16186) );
  INV_X1 U3402 ( .A(n1365), .ZN(n15801) );
  OR2_X1 U3403 ( .A1(n16390), .A2(n15977), .ZN(n15852) );
  AND2_X1 U3417 ( .A1(n24919), .A2(n16360), .ZN(n24842) );
  OR2_X1 U3423 ( .A1(n15938), .A2(n16016), .ZN(n16254) );
  XNOR2_X1 U3436 ( .A(n14520), .B(n14519), .ZN(n15804) );
  MUX2_X1 U3437 ( .A(n15600), .B(n15599), .S(n16063), .Z(n15601) );
  OR2_X1 U3470 ( .A1(n3406), .A2(n16230), .ZN(n5023) );
  INV_X1 U3475 ( .A(n381), .ZN(n24655) );
  INV_X1 U3479 ( .A(n1261), .ZN(n24797) );
  OR2_X1 U3489 ( .A1(n17276), .A2(n17273), .ZN(n16746) );
  OR2_X1 U3492 ( .A1(n15266), .A2(n2253), .ZN(n2250) );
  OR2_X1 U3493 ( .A1(n17277), .A2(n17249), .ZN(n1624) );
  OR2_X1 U3494 ( .A1(n16809), .A2(n17478), .ZN(n2372) );
  OR2_X1 U3498 ( .A1(n16702), .A2(n16618), .ZN(n751) );
  AOI22_X1 U3499 ( .A1(n17144), .A2(n16691), .B1(n16985), .B2(n24688), .ZN(
        n16695) );
  OR2_X1 U3506 ( .A1(n16753), .A2(n17293), .ZN(n17544) );
  INV_X1 U3523 ( .A(n16902), .ZN(n2561) );
  AND2_X1 U3545 ( .A1(n17326), .A2(n17319), .ZN(n1409) );
  OAI21_X1 U3550 ( .B1(n17152), .B2(n17151), .A(n17150), .ZN(n18060) );
  XNOR2_X1 U3568 ( .A(n18532), .B(n4023), .ZN(n17835) );
  INV_X1 U3575 ( .A(n17677), .ZN(n24662) );
  OR2_X1 U3577 ( .A1(n24759), .A2(n24457), .ZN(n647) );
  OR2_X1 U3578 ( .A1(n18816), .A2(n19359), .ZN(n19213) );
  AND2_X1 U3591 ( .A1(n19057), .A2(n988), .ZN(n524) );
  BUF_X1 U3599 ( .A(n19485), .Z(n240) );
  BUF_X1 U3604 ( .A(n17556), .Z(n18919) );
  INV_X1 U3616 ( .A(n18830), .ZN(n19597) );
  INV_X1 U3636 ( .A(n19436), .ZN(n19435) );
  INV_X1 U3640 ( .A(n18493), .ZN(n24728) );
  INV_X1 U3645 ( .A(n20615), .ZN(n24835) );
  XNOR2_X1 U3648 ( .A(n17074), .B(n17073), .ZN(n4291) );
  CLKBUF_X1 U3653 ( .A(n19065), .Z(n19239) );
  OR2_X1 U3658 ( .A1(n18909), .A2(n19570), .ZN(n24099) );
  AND2_X1 U3676 ( .A1(n19491), .A2(n19492), .ZN(n25131) );
  OR2_X1 U3683 ( .A1(n19094), .A2(n25067), .ZN(n19378) );
  INV_X1 U3684 ( .A(n988), .ZN(n280) );
  AOI22_X1 U3695 ( .A1(n19421), .A2(n19166), .B1(n19417), .B2(n19420), .ZN(
        n4580) );
  INV_X1 U3773 ( .A(n1155), .ZN(n3016) );
  OR2_X1 U3775 ( .A1(n19403), .A2(n19186), .ZN(n18893) );
  NAND2_X1 U3791 ( .A1(n18737), .A2(n18738), .ZN(n20183) );
  INV_X1 U3832 ( .A(n19904), .ZN(n24681) );
  OR2_X1 U3838 ( .A1(n19875), .A2(n20022), .ZN(n20564) );
  NAND2_X1 U3855 ( .A1(n1613), .A2(n4176), .ZN(n1326) );
  XNOR2_X1 U3860 ( .A(n22005), .B(n21606), .ZN(n21343) );
  AND2_X1 U3872 ( .A1(n22483), .A2(n22901), .ZN(n24718) );
  OAI21_X1 U3881 ( .B1(n20363), .B2(n24078), .A(n18825), .ZN(n21572) );
  INV_X1 U3944 ( .A(n3213), .ZN(n25123) );
  AND2_X1 U3945 ( .A1(n22239), .A2(n22241), .ZN(n24666) );
  AND2_X1 U3969 ( .A1(n22454), .A2(n22323), .ZN(n22452) );
  OR2_X1 U3975 ( .A1(n24415), .A2(n22138), .ZN(n2828) );
  OR2_X1 U3976 ( .A1(n24881), .A2(n22387), .ZN(n24724) );
  AOI21_X1 U4034 ( .B1(n4062), .B2(n1679), .A(n22113), .ZN(n23578) );
  AND2_X1 U4036 ( .A1(n3895), .A2(n21822), .ZN(n24698) );
  NAND3_X1 U4038 ( .A1(n22277), .A2(n22276), .A3(n1507), .ZN(n23250) );
  AOI21_X1 U4041 ( .B1(n25050), .B2(n22165), .A(n22164), .ZN(n23692) );
  NOR2_X1 U4048 ( .A1(n23723), .A2(n23714), .ZN(n23696) );
  OAI21_X1 U4058 ( .B1(n24322), .B2(n22281), .A(n24631), .ZN(n3718) );
  CLKBUF_X1 U4117 ( .A(n23478), .Z(n23494) );
  OR2_X1 U4134 ( .A1(n22637), .A2(n23595), .ZN(n24668) );
  OR2_X1 U4136 ( .A1(n23930), .A2(n24948), .ZN(n24831) );
  CLKBUF_X1 U4139 ( .A(Key[46]), .Z(n886) );
  CLKBUF_X1 U4181 ( .A(Key[94]), .Z(n3115) );
  CLKBUF_X1 U4184 ( .A(Key[79]), .Z(n2042) );
  CLKBUF_X1 U4189 ( .A(Key[32]), .Z(n2100) );
  CLKBUF_X1 U4208 ( .A(Key[149]), .Z(n21711) );
  OAI211_X1 U4231 ( .C1(n21763), .C2(n22639), .A(n22638), .B(n24668), .ZN(
        n4782) );
  INV_X1 U4249 ( .A(n2215), .ZN(n5484) );
  OR2_X1 U4281 ( .A1(n25572), .A2(n288), .ZN(n24594) );
  AND2_X1 U4305 ( .A1(n7865), .A2(n24576), .ZN(n24595) );
  INV_X1 U4313 ( .A(n7896), .ZN(n24861) );
  INV_X1 U4317 ( .A(n7600), .ZN(n24772) );
  OR2_X1 U4321 ( .A1(n7879), .A2(n7882), .ZN(n24596) );
  NOR2_X1 U4334 ( .A1(n7581), .A2(n7882), .ZN(n24597) );
  AND2_X1 U4339 ( .A1(n7313), .A2(n7883), .ZN(n7881) );
  XOR2_X1 U4366 ( .A(n9035), .B(n5014), .Z(n24598) );
  XOR2_X1 U4370 ( .A(n8326), .B(n5619), .Z(n24599) );
  XOR2_X1 U4402 ( .A(n9141), .B(n1869), .Z(n24600) );
  INV_X1 U4409 ( .A(n11004), .ZN(n24622) );
  XNOR2_X1 U4421 ( .A(n11019), .B(n11018), .ZN(n12656) );
  INV_X1 U4442 ( .A(n12656), .ZN(n24640) );
  OAI21_X1 U4464 ( .B1(n4061), .B2(n3343), .A(n3342), .ZN(n13931) );
  INV_X1 U4468 ( .A(n13931), .ZN(n25128) );
  NOR2_X1 U4483 ( .A1(n14247), .A2(n13935), .ZN(n24602) );
  INV_X1 U4494 ( .A(n12995), .ZN(n24750) );
  XNOR2_X1 U4498 ( .A(n11327), .B(n11326), .ZN(n12791) );
  INV_X1 U4510 ( .A(n13975), .ZN(n24713) );
  OR2_X1 U4557 ( .A1(n14747), .A2(n15625), .ZN(n24603) );
  AND2_X1 U4595 ( .A1(n16796), .A2(n16550), .ZN(n24604) );
  INV_X1 U4640 ( .A(n16809), .ZN(n24660) );
  INV_X1 U4682 ( .A(n19477), .ZN(n24803) );
  OR2_X1 U4696 ( .A1(n19478), .A2(n5070), .ZN(n24605) );
  INV_X1 U4704 ( .A(n19353), .ZN(n19444) );
  XOR2_X1 U4716 ( .A(n18511), .B(n18510), .Z(n24606) );
  INV_X1 U4771 ( .A(n20346), .ZN(n20281) );
  INV_X1 U4792 ( .A(n22804), .ZN(n25160) );
  XNOR2_X1 U4796 ( .A(n20974), .B(n20973), .ZN(n22917) );
  INV_X1 U4822 ( .A(n22917), .ZN(n24674) );
  XOR2_X1 U4846 ( .A(n21125), .B(n21124), .Z(n24607) );
  NAND2_X1 U4862 ( .A1(n21838), .A2(n22354), .ZN(n24608) );
  AND2_X1 U4879 ( .A1(n4112), .A2(n24334), .ZN(n24609) );
  OR2_X1 U4930 ( .A1(n2671), .A2(n22422), .ZN(n24610) );
  OR2_X1 U4940 ( .A1(n23579), .A2(n23578), .ZN(n24611) );
  OR2_X1 U4951 ( .A1(n23196), .A2(n23195), .ZN(n24612) );
  OR2_X1 U4962 ( .A1(n23904), .A2(n607), .ZN(n24613) );
  NAND2_X1 U5011 ( .A1(n16702), .A2(n16703), .ZN(n16709) );
  NAND2_X1 U5050 ( .A1(n16443), .A2(n16242), .ZN(n1095) );
  XNOR2_X2 U5071 ( .A(n15519), .B(n15518), .ZN(n16242) );
  OR2_X1 U5123 ( .A1(n15473), .A2(n17202), .ZN(n24615) );
  NAND2_X1 U5219 ( .A1(n7992), .A2(n7993), .ZN(n7501) );
  NAND2_X1 U5249 ( .A1(n12854), .A2(n13112), .ZN(n12206) );
  AND3_X2 U5253 ( .A1(n24618), .A2(n24848), .A3(n9924), .ZN(n10799) );
  NAND2_X1 U5304 ( .A1(n24847), .A2(n9920), .ZN(n24618) );
  NOR2_X1 U5384 ( .A1(n24604), .A2(n5375), .ZN(n15703) );
  BUF_X1 U5396 ( .A(n22217), .Z(n24918) );
  NAND2_X1 U5398 ( .A1(n24729), .A2(n22729), .ZN(n2364) );
  XNOR2_X2 U5428 ( .A(n20858), .B(n20859), .ZN(n22729) );
  NAND2_X1 U5432 ( .A1(n15044), .A2(n15043), .ZN(n14493) );
  NAND3_X1 U5436 ( .A1(n13780), .A2(n14160), .A3(n13954), .ZN(n15043) );
  NAND3_X1 U5452 ( .A1(n19221), .A2(n5461), .A3(n25010), .ZN(n5442) );
  NAND2_X1 U5455 ( .A1(n19371), .A2(n24424), .ZN(n19221) );
  XNOR2_X2 U5464 ( .A(n24619), .B(n15405), .ZN(n15656) );
  XNOR2_X1 U5471 ( .A(n14186), .B(n4834), .ZN(n24619) );
  NAND2_X1 U5472 ( .A1(n24330), .A2(n17422), .ZN(n17429) );
  NOR2_X1 U5489 ( .A1(n595), .A2(n24620), .ZN(n22870) );
  NAND2_X1 U5500 ( .A1(n3025), .A2(n1738), .ZN(n24620) );
  INV_X1 U5508 ( .A(n24621), .ZN(n24174) );
  OAI21_X1 U5515 ( .B1(n16854), .B2(n368), .A(n16852), .ZN(n24621) );
  NAND2_X1 U5530 ( .A1(n113), .A2(n20041), .ZN(n19866) );
  NAND3_X1 U5546 ( .A1(n10369), .A2(n10364), .A3(n24622), .ZN(n24213) );
  NAND2_X1 U5564 ( .A1(n897), .A2(n24623), .ZN(n8368) );
  NAND3_X1 U5565 ( .A1(n3110), .A2(n3111), .A3(n3109), .ZN(n24623) );
  INV_X1 U5623 ( .A(n23883), .ZN(n24624) );
  NAND2_X1 U5642 ( .A1(n23879), .A2(n24624), .ZN(n107) );
  OAI21_X1 U5707 ( .B1(n3805), .B2(n22687), .A(n3804), .ZN(n24625) );
  NAND3_X1 U5725 ( .A1(n24626), .A2(n23539), .A3(n23540), .ZN(n23542) );
  NAND2_X1 U5750 ( .A1(n23536), .A2(n24057), .ZN(n24626) );
  AOI21_X1 U5758 ( .B1(n23155), .B2(n22446), .A(n24627), .ZN(n22447) );
  NAND2_X1 U5780 ( .A1(n10622), .A2(n11214), .ZN(n24628) );
  NAND2_X1 U5786 ( .A1(n2018), .A2(n2017), .ZN(n2016) );
  MUX2_X1 U5790 ( .A(n23410), .B(n23416), .S(n23403), .Z(n22866) );
  NOR2_X1 U5795 ( .A1(n22849), .A2(n22850), .ZN(n23403) );
  NAND2_X1 U5809 ( .A1(n24264), .A2(n24265), .ZN(n24629) );
  XNOR2_X1 U5873 ( .A(n24630), .B(n23816), .ZN(Ciphertext[157]) );
  NAND3_X1 U5887 ( .A1(n536), .A2(n22541), .A3(n22540), .ZN(n22543) );
  AOI21_X1 U5915 ( .B1(n19980), .B2(n19983), .A(n24315), .ZN(n19985) );
  NAND3_X1 U5954 ( .A1(n19819), .A2(n19820), .A3(n19818), .ZN(n742) );
  NAND2_X1 U6014 ( .A1(n24552), .A2(n12976), .ZN(n12981) );
  NAND2_X1 U6048 ( .A1(n24865), .A2(n2581), .ZN(n24632) );
  NAND3_X1 U6090 ( .A1(n776), .A2(n22125), .A3(n22421), .ZN(n22126) );
  AOI21_X2 U6139 ( .B1(n20895), .B2(n2364), .A(n20894), .ZN(n23647) );
  NAND3_X1 U6166 ( .A1(n17252), .A2(n17279), .A3(n17273), .ZN(n14748) );
  NAND3_X1 U6171 ( .A1(n24571), .A2(n14510), .A3(n24713), .ZN(n24712) );
  NAND2_X1 U6191 ( .A1(n25383), .A2(n19573), .ZN(n2018) );
  NAND2_X2 U6252 ( .A1(n24633), .A2(n12857), .ZN(n14321) );
  NAND3_X2 U6310 ( .A1(n17291), .A2(n24196), .A3(n24635), .ZN(n18512) );
  NAND3_X1 U6322 ( .A1(n3539), .A2(n4424), .A3(n24636), .ZN(n3538) );
  NAND2_X1 U6325 ( .A1(n296), .A2(n14031), .ZN(n24636) );
  NAND3_X1 U6331 ( .A1(n23787), .A2(n2476), .A3(n21902), .ZN(n2475) );
  NAND2_X1 U6351 ( .A1(n24641), .A2(n24640), .ZN(n24639) );
  NAND2_X1 U6353 ( .A1(n12742), .A2(n12740), .ZN(n24641) );
  NAND2_X1 U6382 ( .A1(n12511), .A2(n12656), .ZN(n24642) );
  XNOR2_X1 U6389 ( .A(n24643), .B(n22195), .ZN(Ciphertext[126]) );
  NAND3_X1 U6402 ( .A1(n22194), .A2(n22193), .A3(n22998), .ZN(n24643) );
  NOR2_X1 U6410 ( .A1(n24644), .A2(n25345), .ZN(n98) );
  AND2_X1 U6411 ( .A1(n17192), .A2(n4039), .ZN(n24650) );
  NAND2_X1 U6479 ( .A1(n19449), .A2(n25002), .ZN(n24646) );
  NAND2_X1 U6481 ( .A1(n19444), .A2(n19445), .ZN(n24647) );
  BUF_X2 U6555 ( .A(n22593), .Z(n24043) );
  AND2_X2 U6558 ( .A1(n22595), .A2(n22594), .ZN(n23040) );
  NAND2_X1 U6559 ( .A1(n5018), .A2(n24650), .ZN(n5017) );
  NAND2_X1 U6570 ( .A1(n17196), .A2(n17031), .ZN(n5018) );
  NAND2_X1 U6598 ( .A1(n24595), .A2(n4536), .ZN(n24652) );
  NAND2_X1 U6607 ( .A1(n16159), .A2(n24653), .ZN(n17395) );
  NAND3_X1 U6623 ( .A1(n24656), .A2(n24655), .A3(n24654), .ZN(n24653) );
  NAND2_X1 U6638 ( .A1(n16154), .A2(n24458), .ZN(n24654) );
  NAND2_X1 U6663 ( .A1(n16122), .A2(n16124), .ZN(n24656) );
  NAND2_X1 U6690 ( .A1(n5152), .A2(n24657), .ZN(n20961) );
  OAI21_X1 U6715 ( .B1(n5155), .B2(n19576), .A(n24658), .ZN(n24657) );
  INV_X1 U6717 ( .A(n25072), .ZN(n24658) );
  OAI211_X2 U6737 ( .C1(n5391), .C2(n3760), .A(n10379), .B(n24659), .ZN(n12151) );
  NAND2_X1 U6760 ( .A1(n991), .A2(n416), .ZN(n24659) );
  NAND2_X1 U6771 ( .A1(n24660), .A2(n17081), .ZN(n17480) );
  NAND2_X1 U6788 ( .A1(n3908), .A2(n22329), .ZN(n3907) );
  NAND3_X1 U6810 ( .A1(n23139), .A2(n23131), .A3(n24473), .ZN(n23132) );
  AND4_X2 U6825 ( .A1(n24790), .A2(n3660), .A3(n3772), .A4(n3665), .ZN(n20415)
         );
  NAND2_X1 U6826 ( .A1(n7349), .A2(n7348), .ZN(n7279) );
  XNOR2_X1 U6837 ( .A(n24661), .B(n23137), .ZN(Ciphertext[18]) );
  NAND2_X1 U6846 ( .A1(n23136), .A2(n23135), .ZN(n24661) );
  XNOR2_X1 U6852 ( .A(n797), .B(n24662), .ZN(n18990) );
  NAND3_X1 U6881 ( .A1(n3165), .A2(n17674), .A3(n5280), .ZN(n17675) );
  NAND2_X1 U6893 ( .A1(n24785), .A2(n14278), .ZN(n24664) );
  OR2_X2 U6895 ( .A1(n24665), .A2(n16811), .ZN(n18418) );
  AOI22_X1 U6900 ( .A1(n16807), .A2(n16896), .B1(n16806), .B2(n17078), .ZN(
        n24665) );
  OR2_X1 U6901 ( .A1(n4066), .A2(n20140), .ZN(n5445) );
  AOI21_X2 U6903 ( .B1(n4550), .B2(n19589), .A(n4549), .ZN(n20909) );
  NAND3_X1 U6909 ( .A1(n4434), .A2(n23799), .A3(n23001), .ZN(n23786) );
  NAND2_X1 U6916 ( .A1(n22243), .A2(n24666), .ZN(n2885) );
  XNOR2_X2 U6925 ( .A(n24667), .B(n5369), .ZN(n18959) );
  XNOR2_X1 U6929 ( .A(n17852), .B(n18225), .ZN(n24667) );
  NAND2_X2 U6955 ( .A1(n1958), .A2(n1960), .ZN(n7349) );
  NAND3_X1 U7024 ( .A1(n9952), .A2(n9953), .A3(n9951), .ZN(n9954) );
  INV_X1 U7035 ( .A(n7157), .ZN(n7363) );
  NAND2_X1 U7038 ( .A1(n7629), .A2(n7155), .ZN(n7157) );
  NAND3_X1 U7043 ( .A1(n21763), .A2(n24611), .A3(n24901), .ZN(n21943) );
  NAND2_X1 U7052 ( .A1(n10364), .A2(n10369), .ZN(n2751) );
  NAND2_X1 U7067 ( .A1(n19318), .A2(n4874), .ZN(n17564) );
  NAND2_X1 U7082 ( .A1(n13107), .A2(n13661), .ZN(n24669) );
  NAND2_X1 U7090 ( .A1(n24671), .A2(n24670), .ZN(n13698) );
  NAND2_X1 U7091 ( .A1(n13932), .A2(n14241), .ZN(n24670) );
  NAND2_X1 U7121 ( .A1(n13697), .A2(n4116), .ZN(n24671) );
  NAND2_X1 U7129 ( .A1(n13633), .A2(n13935), .ZN(n13697) );
  AOI21_X1 U7147 ( .B1(n22917), .B2(n22918), .A(n22072), .ZN(n24672) );
  NAND2_X1 U7149 ( .A1(n24674), .A2(n21712), .ZN(n24673) );
  OAI22_X1 U7155 ( .A1(n25240), .A2(n24675), .B1(n24428), .B2(n24469), .ZN(
        n22983) );
  INV_X1 U7166 ( .A(n23865), .ZN(n24675) );
  NOR2_X2 U7176 ( .A1(n12647), .A2(n24677), .ZN(n14988) );
  NAND2_X1 U7191 ( .A1(n3885), .A2(n3884), .ZN(n24677) );
  AOI21_X2 U7192 ( .B1(n13639), .B2(n13638), .A(n24678), .ZN(n14792) );
  NOR2_X1 U7194 ( .A1(n13697), .A2(n24679), .ZN(n24678) );
  OR2_X1 U7201 ( .A1(n25247), .A2(n14053), .ZN(n2756) );
  INV_X1 U7206 ( .A(n14553), .ZN(n15200) );
  NOR2_X2 U7230 ( .A1(n24680), .A2(n24602), .ZN(n14553) );
  OAI21_X1 U7252 ( .B1(n13204), .B2(n4116), .A(n13202), .ZN(n24680) );
  NAND2_X1 U7259 ( .A1(n4407), .A2(n4406), .ZN(n24270) );
  NAND2_X1 U7262 ( .A1(n23392), .A2(n24465), .ZN(n4412) );
  NAND2_X1 U7273 ( .A1(n17401), .A2(n17402), .ZN(n18484) );
  AOI22_X2 U7276 ( .A1(n19828), .A2(n19827), .B1(n24682), .B2(n24681), .ZN(
        n21561) );
  NOR2_X1 U7280 ( .A1(n17016), .A2(n17208), .ZN(n16257) );
  NAND3_X1 U7295 ( .A1(n16253), .A2(n24684), .A3(n24683), .ZN(n2093) );
  NAND2_X1 U7301 ( .A1(n25389), .A2(n16016), .ZN(n24683) );
  OR2_X1 U7307 ( .A1(n16016), .A2(n16247), .ZN(n24684) );
  NAND2_X1 U7326 ( .A1(n15869), .A2(n17114), .ZN(n24685) );
  NAND2_X1 U7328 ( .A1(n19093), .A2(n18877), .ZN(n24721) );
  NAND2_X1 U7331 ( .A1(n24687), .A2(n24686), .ZN(n2638) );
  NAND2_X1 U7344 ( .A1(n15945), .A2(n16443), .ZN(n24686) );
  NAND2_X1 U7348 ( .A1(n15944), .A2(n16437), .ZN(n24687) );
  NAND3_X1 U7373 ( .A1(n25154), .A2(n24596), .A3(n7584), .ZN(n1779) );
  NAND3_X1 U7375 ( .A1(n10190), .A2(n10859), .A3(n10860), .ZN(n10864) );
  NAND2_X1 U7376 ( .A1(n24689), .A2(n25189), .ZN(n9342) );
  NAND2_X1 U7378 ( .A1(n25187), .A2(n25188), .ZN(n24689) );
  NAND2_X1 U7384 ( .A1(n7688), .A2(n7217), .ZN(n7216) );
  NOR2_X2 U7419 ( .A1(n18822), .A2(n18823), .ZN(n20484) );
  OAI21_X1 U7434 ( .B1(n3563), .B2(n14000), .A(n24691), .ZN(n13678) );
  XNOR2_X1 U7445 ( .A(n17969), .B(n2137), .ZN(n17927) );
  OAI21_X1 U7458 ( .B1(n23886), .B2(n23885), .A(n24692), .ZN(n23887) );
  NAND3_X1 U7479 ( .A1(n24765), .A2(n24610), .A3(n3713), .ZN(n23285) );
  OAI21_X1 U7525 ( .B1(n22982), .B2(n23860), .A(n24694), .ZN(n22985) );
  NAND3_X1 U7570 ( .A1(n24675), .A2(n23857), .A3(n23862), .ZN(n24694) );
  OR2_X1 U7633 ( .A1(n13946), .A2(n13947), .ZN(n24697) );
  AOI21_X2 U7635 ( .B1(n24698), .B2(n3896), .A(n21842), .ZN(n23890) );
  INV_X1 U7642 ( .A(n10918), .ZN(n1940) );
  OAI21_X1 U7656 ( .B1(n16591), .B2(n17076), .A(n16892), .ZN(n24699) );
  NAND2_X1 U7688 ( .A1(n974), .A2(n975), .ZN(n976) );
  OR2_X1 U7696 ( .A1(n19075), .A2(n19076), .ZN(n24700) );
  OAI21_X2 U7697 ( .B1(n13595), .B2(n14337), .A(n24701), .ZN(n15347) );
  OAI211_X1 U7717 ( .C1(n23909), .C2(n23908), .A(n24613), .B(n24702), .ZN(
        n23910) );
  NAND2_X1 U7718 ( .A1(n23907), .A2(n23906), .ZN(n24702) );
  NAND2_X1 U7719 ( .A1(n24703), .A2(n24012), .ZN(n24281) );
  OAI21_X1 U7723 ( .B1(n23982), .B2(n24008), .A(n23984), .ZN(n24703) );
  OAI22_X1 U7794 ( .A1(n20469), .A2(n5115), .B1(n5114), .B2(n20473), .ZN(
        n24704) );
  AND2_X1 U7803 ( .A1(n21847), .A2(n21816), .ZN(n22353) );
  NAND3_X1 U7842 ( .A1(n24706), .A2(n20418), .A3(n25108), .ZN(n20420) );
  NAND2_X1 U7845 ( .A1(n4509), .A2(n20401), .ZN(n24706) );
  OAI21_X1 U7846 ( .B1(n25022), .B2(n22667), .A(n24707), .ZN(n22787) );
  NAND2_X1 U7851 ( .A1(n25022), .A2(n22782), .ZN(n24707) );
  NAND3_X2 U7854 ( .A1(n15713), .A2(n15711), .A3(n15712), .ZN(n17299) );
  NAND2_X1 U7855 ( .A1(n7044), .A2(n3730), .ZN(n551) );
  OAI211_X2 U7864 ( .C1(n10705), .C2(n2754), .A(n10704), .B(n24709), .ZN(n1568) );
  NAND2_X1 U7875 ( .A1(n10700), .A2(n10701), .ZN(n24709) );
  NAND3_X1 U7889 ( .A1(n24711), .A2(n14306), .A3(n24710), .ZN(n24153) );
  INV_X1 U7891 ( .A(n24588), .ZN(n24711) );
  NAND2_X1 U7907 ( .A1(n24714), .A2(n24712), .ZN(n13980) );
  NAND2_X1 U7924 ( .A1(n5752), .A2(n24715), .ZN(n24714) );
  INV_X1 U7934 ( .A(n14510), .ZN(n24715) );
  NAND2_X1 U7960 ( .A1(n5052), .A2(n16844), .ZN(n16845) );
  NAND2_X1 U7969 ( .A1(n19479), .A2(n19480), .ZN(n24716) );
  NAND2_X1 U7981 ( .A1(n16147), .A2(n16096), .ZN(n16145) );
  NAND2_X1 U7988 ( .A1(n19719), .A2(n24717), .ZN(n18774) );
  NAND2_X1 U8036 ( .A1(n24278), .A2(n24279), .ZN(n22879) );
  NAND2_X1 U8044 ( .A1(n20546), .A2(n20127), .ZN(n19674) );
  NAND2_X1 U8058 ( .A1(n16556), .A2(n16557), .ZN(n4450) );
  NAND2_X1 U8097 ( .A1(n23714), .A2(n23723), .ZN(n23728) );
  OAI21_X2 U8113 ( .B1(n22055), .B2(n22054), .A(n22053), .ZN(n23723) );
  AND2_X2 U8115 ( .A1(n19209), .A2(n3106), .ZN(n20576) );
  NAND2_X1 U8124 ( .A1(n25382), .A2(n24718), .ZN(n22846) );
  NOR2_X1 U8213 ( .A1(n24720), .A2(n17449), .ZN(n17150) );
  NAND3_X1 U8220 ( .A1(n6077), .A2(n6076), .A3(n6883), .ZN(n2786) );
  NOR2_X1 U8229 ( .A1(n17148), .A2(n17455), .ZN(n24720) );
  NAND2_X1 U8240 ( .A1(n4730), .A2(n4731), .ZN(n10753) );
  NAND2_X1 U8248 ( .A1(n24721), .A2(n24335), .ZN(n18879) );
  NAND2_X1 U8268 ( .A1(n20131), .A2(n20522), .ZN(n19971) );
  NOR2_X1 U8284 ( .A1(n22849), .A2(n22850), .ZN(n25035) );
  OAI21_X1 U8285 ( .B1(n22848), .B2(n22847), .A(n22846), .ZN(n22849) );
  NAND2_X1 U8306 ( .A1(n20066), .A2(n20071), .ZN(n24722) );
  NAND2_X1 U8310 ( .A1(n5759), .A2(n16676), .ZN(n16678) );
  NOR2_X1 U8313 ( .A1(n16824), .A2(n16862), .ZN(n807) );
  NOR2_X1 U8314 ( .A1(n282), .A2(n16112), .ZN(n16862) );
  AND2_X2 U8331 ( .A1(n24723), .A2(n5997), .ZN(n7609) );
  NAND2_X1 U8339 ( .A1(n3167), .A2(n5996), .ZN(n24723) );
  NAND2_X1 U8343 ( .A1(n1978), .A2(n1977), .ZN(n19875) );
  OR2_X1 U8350 ( .A1(n10884), .A2(n10885), .ZN(n24167) );
  XNOR2_X2 U8356 ( .A(n21698), .B(n21697), .ZN(n22904) );
  NAND3_X2 U8357 ( .A1(n24269), .A2(n4572), .A3(n4573), .ZN(n18261) );
  NAND2_X1 U8369 ( .A1(n2660), .A2(n2708), .ZN(n2710) );
  NAND2_X1 U8372 ( .A1(n24725), .A2(n642), .ZN(n12465) );
  NAND2_X1 U8375 ( .A1(n401), .A2(n12533), .ZN(n24725) );
  NAND2_X1 U8376 ( .A1(n3046), .A2(n20211), .ZN(n3045) );
  NAND2_X1 U8395 ( .A1(n24726), .A2(n18299), .ZN(n1716) );
  NAND2_X1 U8418 ( .A1(n3752), .A2(n3751), .ZN(n24726) );
  NAND2_X1 U8427 ( .A1(n9468), .A2(n1595), .ZN(n3291) );
  NAND2_X1 U8440 ( .A1(n24442), .A2(n23481), .ZN(n2997) );
  NAND2_X1 U8446 ( .A1(n2168), .A2(n20478), .ZN(n20356) );
  AND3_X2 U8454 ( .A1(n4768), .A2(n4769), .A3(n4770), .ZN(n14789) );
  OAI21_X1 U8455 ( .B1(n24172), .B2(n19464), .A(n24727), .ZN(n19462) );
  NAND2_X1 U8459 ( .A1(n19464), .A2(n19457), .ZN(n24727) );
  XNOR2_X1 U8465 ( .A(n18494), .B(n24728), .ZN(n25072) );
  NOR2_X1 U8469 ( .A1(n22889), .A2(n22093), .ZN(n24729) );
  NAND2_X1 U8477 ( .A1(n20136), .A2(n20134), .ZN(n20016) );
  NAND2_X1 U8483 ( .A1(n25248), .A2(n13303), .ZN(n3847) );
  NAND3_X1 U8487 ( .A1(n4714), .A2(n5428), .A3(n24730), .ZN(n17592) );
  NAND3_X1 U8493 ( .A1(n16572), .A2(n17115), .A3(n890), .ZN(n24730) );
  XOR2_X1 U8542 ( .A(n24383), .B(n924), .Z(n24769) );
  NAND2_X1 U8567 ( .A1(n1355), .A2(n14048), .ZN(n14053) );
  NAND2_X1 U8577 ( .A1(n14141), .A2(n14189), .ZN(n14188) );
  NAND3_X1 U8578 ( .A1(n291), .A2(n24098), .A3(n16043), .ZN(n1897) );
  NAND2_X1 U8580 ( .A1(n10399), .A2(n10659), .ZN(n10315) );
  BUF_X1 U8583 ( .A(n20036), .Z(n22056) );
  AOI21_X1 U8600 ( .B1(n2253), .B2(n15789), .A(n24098), .ZN(n15536) );
  NAND2_X1 U8618 ( .A1(n16706), .A2(n16705), .ZN(n16707) );
  NAND2_X1 U8632 ( .A1(n20242), .A2(n19937), .ZN(n19821) );
  AOI21_X2 U8648 ( .B1(n19338), .B2(n19337), .A(n19336), .ZN(n20242) );
  NAND2_X1 U8663 ( .A1(n548), .A2(n549), .ZN(n24733) );
  NAND2_X1 U8687 ( .A1(n24184), .A2(n22052), .ZN(n22053) );
  NAND2_X1 U8695 ( .A1(n24734), .A2(n14305), .ZN(n15275) );
  NOR2_X1 U8726 ( .A1(n1526), .A2(n1450), .ZN(n24734) );
  NAND2_X1 U8729 ( .A1(n24735), .A2(n11174), .ZN(n11179) );
  NAND2_X1 U8731 ( .A1(n11170), .A2(n24736), .ZN(n24735) );
  INV_X1 U8774 ( .A(n11168), .ZN(n24736) );
  XNOR2_X1 U8776 ( .A(n24737), .B(n11924), .ZN(n861) );
  XNOR2_X1 U8803 ( .A(n11923), .B(n11922), .ZN(n24737) );
  NAND2_X1 U8816 ( .A1(n4514), .A2(n1619), .ZN(n4513) );
  OAI21_X1 U8870 ( .B1(n20069), .B2(n20072), .A(n24738), .ZN(n19854) );
  NAND3_X1 U8882 ( .A1(n19852), .A2(n19660), .A3(n20068), .ZN(n24738) );
  INV_X1 U8915 ( .A(n10103), .ZN(n24740) );
  NAND2_X1 U8918 ( .A1(n524), .A2(n354), .ZN(n1132) );
  NAND2_X1 U8930 ( .A1(n15621), .A2(n24537), .ZN(n24741) );
  NAND2_X1 U8932 ( .A1(n19091), .A2(n19904), .ZN(n2916) );
  NAND2_X2 U8960 ( .A1(n12714), .A2(n24742), .ZN(n14439) );
  OAI21_X1 U8967 ( .B1(n12708), .B2(n12709), .A(n13078), .ZN(n24742) );
  NAND2_X1 U8968 ( .A1(n24743), .A2(n16497), .ZN(n17581) );
  OAI21_X1 U8969 ( .B1(n16487), .B2(n16488), .A(n368), .ZN(n24743) );
  NAND2_X1 U8984 ( .A1(n24746), .A2(n24744), .ZN(n5330) );
  NAND2_X1 U8988 ( .A1(n13785), .A2(n14190), .ZN(n24745) );
  NAND2_X1 U8989 ( .A1(n13787), .A2(n24347), .ZN(n24746) );
  NAND2_X1 U8992 ( .A1(n4946), .A2(n12539), .ZN(n12984) );
  NAND2_X1 U9012 ( .A1(n16138), .A2(n24747), .ZN(n18195) );
  NAND2_X1 U9018 ( .A1(n16780), .A2(n25256), .ZN(n24747) );
  AOI21_X1 U9028 ( .B1(n20328), .B2(n20329), .A(n24749), .ZN(n20334) );
  NAND2_X1 U9032 ( .A1(n11328), .A2(n12791), .ZN(n12793) );
  NAND2_X1 U9037 ( .A1(n2883), .A2(n3257), .ZN(n8506) );
  AOI22_X1 U9041 ( .A1(n17449), .A2(n16980), .B1(n16979), .B2(n17455), .ZN(
        n16369) );
  NAND2_X1 U9076 ( .A1(n24751), .A2(n1806), .ZN(n2198) );
  OAI21_X1 U9080 ( .B1(n19239), .B2(n24606), .A(n19614), .ZN(n24751) );
  NAND2_X1 U9094 ( .A1(n7002), .A2(n7003), .ZN(n4150) );
  NAND2_X1 U9097 ( .A1(n3860), .A2(n4788), .ZN(n14059) );
  NAND2_X1 U9098 ( .A1(n24752), .A2(n5379), .ZN(n5382) );
  NAND3_X1 U9099 ( .A1(n4281), .A2(n4143), .A3(n24753), .ZN(n24752) );
  XNOR2_X1 U9113 ( .A(n24754), .B(n21553), .ZN(n18045) );
  NAND3_X1 U9133 ( .A1(n2790), .A2(n16259), .A3(n2789), .ZN(n24754) );
  NAND2_X2 U9148 ( .A1(n24755), .A2(n13492), .ZN(n15514) );
  NAND2_X1 U9152 ( .A1(n24815), .A2(n25036), .ZN(n24755) );
  NAND3_X1 U9164 ( .A1(n18385), .A2(n24757), .A3(n24756), .ZN(n4792) );
  NAND2_X1 U9195 ( .A1(n25195), .A2(n19176), .ZN(n24756) );
  NAND2_X1 U9196 ( .A1(n19177), .A2(n18777), .ZN(n24757) );
  INV_X1 U9203 ( .A(n19183), .ZN(n24758) );
  NAND2_X1 U9204 ( .A1(n19297), .A2(n19296), .ZN(n24759) );
  XNOR2_X1 U9208 ( .A(n15238), .B(n1362), .ZN(n14867) );
  NOR2_X2 U9211 ( .A1(n14323), .A2(n654), .ZN(n15238) );
  NAND2_X1 U9217 ( .A1(n17296), .A2(n1535), .ZN(n17300) );
  NAND2_X1 U9219 ( .A1(n24855), .A2(n15704), .ZN(n1535) );
  NAND3_X1 U9257 ( .A1(n6261), .A2(n6259), .A3(n6260), .ZN(n6263) );
  NAND2_X1 U9264 ( .A1(n24764), .A2(n24763), .ZN(n15740) );
  NAND3_X1 U9268 ( .A1(n2587), .A2(n16795), .A3(n16550), .ZN(n24763) );
  NAND2_X1 U9336 ( .A1(n15739), .A2(n4554), .ZN(n24764) );
  NAND2_X1 U9341 ( .A1(n22424), .A2(n22945), .ZN(n24765) );
  NAND2_X1 U9384 ( .A1(n9661), .A2(n422), .ZN(n24767) );
  OR3_X1 U9385 ( .A1(n13234), .A2(n12902), .A3(n12935), .ZN(n2545) );
  OAI21_X2 U9402 ( .B1(n16586), .B2(n16587), .A(n16585), .ZN(n18042) );
  NAND3_X1 U9417 ( .A1(n21767), .A2(n25018), .A3(n22156), .ZN(n24768) );
  NAND2_X1 U9424 ( .A1(n22270), .A2(n22453), .ZN(n22451) );
  NAND2_X1 U9471 ( .A1(n2806), .A2(n2004), .ZN(n2175) );
  NAND2_X1 U9490 ( .A1(n98), .A2(n101), .ZN(n1995) );
  NAND3_X1 U9509 ( .A1(n24770), .A2(n17253), .A3(n17250), .ZN(n720) );
  NAND2_X1 U9513 ( .A1(n17247), .A2(n17248), .ZN(n24770) );
  NOR2_X1 U9536 ( .A1(n13265), .A2(n13267), .ZN(n24805) );
  NAND3_X1 U9567 ( .A1(n647), .A2(n4076), .A3(n17942), .ZN(n24217) );
  OAI211_X1 U9595 ( .C1(n7752), .C2(n2640), .A(n7751), .B(n24771), .ZN(n7753)
         );
  NAND2_X1 U9624 ( .A1(n8014), .A2(n7749), .ZN(n24771) );
  NAND2_X1 U9627 ( .A1(n24801), .A2(n24603), .ZN(n17249) );
  NAND2_X1 U9644 ( .A1(n7341), .A2(n7602), .ZN(n7596) );
  NAND3_X1 U9670 ( .A1(n6459), .A2(n6456), .A3(n6454), .ZN(n6032) );
  XNOR2_X2 U9676 ( .A(n14491), .B(n14492), .ZN(n15611) );
  NAND3_X1 U9678 ( .A1(n13743), .A2(n13744), .A3(n24773), .ZN(n2071) );
  NAND2_X1 U9682 ( .A1(n15726), .A2(n24774), .ZN(n15727) );
  INV_X1 U9708 ( .A(n19446), .ZN(n17711) );
  NAND2_X1 U9720 ( .A1(n19645), .A2(n20027), .ZN(n19649) );
  NAND2_X1 U9725 ( .A1(n10137), .A2(n10138), .ZN(n9174) );
  NAND3_X1 U9726 ( .A1(n6812), .A2(n6367), .A3(n6815), .ZN(n6813) );
  NAND2_X1 U9731 ( .A1(n6367), .A2(n6368), .ZN(n6812) );
  NAND2_X1 U9739 ( .A1(n17230), .A2(n24775), .ZN(n14588) );
  NAND2_X1 U9740 ( .A1(n22947), .A2(n2674), .ZN(n22125) );
  NAND2_X1 U9751 ( .A1(n10584), .A2(n10583), .ZN(n10370) );
  INV_X1 U9752 ( .A(n9460), .ZN(n24844) );
  NAND2_X1 U9756 ( .A1(n16299), .A2(n24506), .ZN(n24777) );
  NAND3_X1 U9758 ( .A1(n17186), .A2(n17025), .A3(n3602), .ZN(n16213) );
  NAND2_X1 U9774 ( .A1(n22888), .A2(n22887), .ZN(n22727) );
  INV_X1 U9790 ( .A(n11622), .ZN(n12335) );
  XNOR2_X1 U9793 ( .A(n11622), .B(n24778), .ZN(n11181) );
  NOR2_X2 U9797 ( .A1(n10340), .A2(n10339), .ZN(n11622) );
  NAND2_X1 U9799 ( .A1(n24779), .A2(n6986), .ZN(n5636) );
  NAND2_X1 U9801 ( .A1(n2646), .A2(n6639), .ZN(n24779) );
  XNOR2_X1 U9805 ( .A(n17806), .B(n20046), .ZN(n17619) );
  OAI22_X2 U9806 ( .A1(n4414), .A2(n4413), .B1(n17176), .B2(n17177), .ZN(
        n17806) );
  XNOR2_X1 U9815 ( .A(n24780), .B(n23825), .ZN(Ciphertext[159]) );
  OAI211_X1 U9831 ( .C1(n23823), .C2(n23824), .A(n23822), .B(n23821), .ZN(
        n24780) );
  AND2_X2 U9832 ( .A1(n24782), .A2(n24781), .ZN(n23650) );
  OAI211_X2 U9869 ( .C1(n16568), .C2(n17227), .A(n16566), .B(n24783), .ZN(
        n18530) );
  NAND3_X1 U9883 ( .A1(n16565), .A2(n17225), .A3(n17224), .ZN(n24783) );
  NAND2_X1 U9893 ( .A1(n939), .A2(n11032), .ZN(n3467) );
  NAND3_X1 U9918 ( .A1(n13975), .A2(n14439), .A3(n24571), .ZN(n14434) );
  NAND3_X1 U9919 ( .A1(n24784), .A2(n8512), .A3(n24224), .ZN(n24851) );
  NAND2_X1 U9928 ( .A1(n1279), .A2(n8511), .ZN(n24784) );
  NAND2_X1 U9976 ( .A1(n1108), .A2(n19786), .ZN(n3214) );
  NAND2_X1 U9982 ( .A1(n19986), .A2(n19784), .ZN(n19786) );
  INV_X1 U9989 ( .A(n21352), .ZN(n21363) );
  INV_X1 U10000 ( .A(n14278), .ZN(n4767) );
  NAND3_X2 U10004 ( .A1(n5156), .A2(n1970), .A3(n12609), .ZN(n14278) );
  NAND3_X1 U10005 ( .A1(n23947), .A2(n24910), .A3(n23952), .ZN(n463) );
  XNOR2_X2 U10012 ( .A(n8678), .B(n8679), .ZN(n9981) );
  NAND2_X1 U10025 ( .A1(n21390), .A2(n21389), .ZN(n23155) );
  NAND2_X1 U10056 ( .A1(n23065), .A2(n23066), .ZN(n22872) );
  NAND2_X1 U10059 ( .A1(n14198), .A2(n3888), .ZN(n13804) );
  NAND2_X2 U10063 ( .A1(n5402), .A2(n12631), .ZN(n3888) );
  OR2_X1 U10070 ( .A1(n18979), .A2(n19456), .ZN(n19031) );
  NAND2_X1 U10072 ( .A1(n14708), .A2(n24928), .ZN(n16686) );
  OR2_X1 U10075 ( .A1(n19097), .A2(n2216), .ZN(n18726) );
  NAND2_X1 U10079 ( .A1(n2643), .A2(n18865), .ZN(n19236) );
  NAND2_X1 U10082 ( .A1(n15859), .A2(n16120), .ZN(n24786) );
  NAND2_X1 U10097 ( .A1(n15858), .A2(n15857), .ZN(n24787) );
  INV_X1 U10098 ( .A(n24864), .ZN(n24788) );
  NAND2_X1 U10110 ( .A1(n13526), .A2(n13466), .ZN(n3331) );
  XNOR2_X1 U10133 ( .A(n24789), .B(n4761), .ZN(Ciphertext[7]) );
  NAND3_X1 U10224 ( .A1(n1210), .A2(n24087), .A3(n10148), .ZN(n2732) );
  NAND3_X1 U10225 ( .A1(n21361), .A2(n318), .A3(n23828), .ZN(n1934) );
  NAND2_X1 U10253 ( .A1(n2396), .A2(n22313), .ZN(n22314) );
  NAND2_X1 U10270 ( .A1(n279), .A2(n19541), .ZN(n24790) );
  OAI211_X1 U10286 ( .C1(n3868), .C2(n11214), .A(n233), .B(n24791), .ZN(n543)
         );
  NAND2_X1 U10289 ( .A1(n11214), .A2(n11215), .ZN(n24791) );
  NAND2_X1 U10296 ( .A1(n1340), .A2(n23219), .ZN(n23222) );
  NAND2_X1 U10327 ( .A1(n20785), .A2(n20786), .ZN(n23219) );
  NAND2_X1 U10333 ( .A1(n9943), .A2(n9945), .ZN(n9287) );
  XNOR2_X2 U10347 ( .A(n8123), .B(n8122), .ZN(n9945) );
  NAND2_X1 U10404 ( .A1(n18951), .A2(n3215), .ZN(n19784) );
  NAND3_X1 U10405 ( .A1(n17762), .A2(n24477), .A3(n19389), .ZN(n17763) );
  XNOR2_X1 U10433 ( .A(n24794), .B(n1854), .ZN(Ciphertext[56]) );
  NOR2_X2 U10448 ( .A1(n17765), .A2(n17766), .ZN(n20109) );
  NAND2_X1 U10449 ( .A1(n16769), .A2(n24569), .ZN(n24863) );
  NAND2_X1 U10451 ( .A1(n22969), .A2(n22968), .ZN(n22416) );
  NAND2_X1 U10462 ( .A1(n25120), .A2(n25119), .ZN(n24795) );
  OAI211_X1 U10533 ( .C1(n16120), .C2(n15611), .A(n24797), .B(n24796), .ZN(
        n5178) );
  NAND2_X1 U10573 ( .A1(n16120), .A2(n16118), .ZN(n24796) );
  NAND3_X1 U10576 ( .A1(n366), .A2(n2566), .A3(n24798), .ZN(n1035) );
  NAND2_X1 U10577 ( .A1(n4284), .A2(n4285), .ZN(n24798) );
  NAND2_X1 U10582 ( .A1(n24800), .A2(n24799), .ZN(n11892) );
  NAND2_X1 U10590 ( .A1(n10479), .A2(n10628), .ZN(n24800) );
  INV_X1 U10602 ( .A(n9990), .ZN(n25121) );
  MUX2_X1 U10612 ( .A(n19132), .B(n19304), .S(n19133), .Z(n16504) );
  NAND2_X1 U10623 ( .A1(n2733), .A2(n7324), .ZN(n1254) );
  NAND2_X1 U10631 ( .A1(n14745), .A2(n14744), .ZN(n24801) );
  OAI21_X1 U10642 ( .B1(n19476), .B2(n24803), .A(n24802), .ZN(n19483) );
  NAND2_X1 U10668 ( .A1(n19476), .A2(n18734), .ZN(n24802) );
  NAND2_X1 U10710 ( .A1(n19641), .A2(n5115), .ZN(n19642) );
  NAND3_X1 U10735 ( .A1(n3974), .A2(n10360), .A3(n12506), .ZN(n3633) );
  OAI21_X1 U10766 ( .B1(n25183), .B2(n20846), .A(n1156), .ZN(n23619) );
  NAND2_X1 U10807 ( .A1(n12832), .A2(n24805), .ZN(n5645) );
  NAND2_X1 U10826 ( .A1(n4066), .A2(n20140), .ZN(n4615) );
  NAND2_X2 U10845 ( .A1(n4245), .A2(n4067), .ZN(n4066) );
  NAND2_X1 U10863 ( .A1(n13336), .A2(n231), .ZN(n12839) );
  XNOR2_X2 U10909 ( .A(n10299), .B(n10300), .ZN(n12506) );
  XNOR2_X1 U10930 ( .A(n12303), .B(n12269), .ZN(n10300) );
  NAND2_X1 U10936 ( .A1(n17284), .A2(n17288), .ZN(n16753) );
  OAI21_X1 U10945 ( .B1(n17124), .B2(n17123), .A(n24806), .ZN(n4661) );
  INV_X1 U10960 ( .A(n17824), .ZN(n24806) );
  OAI211_X1 U10963 ( .C1(n19352), .C2(n24809), .A(n19451), .B(n24808), .ZN(
        n24807) );
  NAND2_X1 U10984 ( .A1(n19352), .A2(n19357), .ZN(n24808) );
  NOR2_X1 U10986 ( .A1(n6068), .A2(n24810), .ZN(n7278) );
  NAND3_X1 U11013 ( .A1(n9660), .A2(n9659), .A3(n9745), .ZN(n1943) );
  NAND2_X1 U11021 ( .A1(n3737), .A2(n23851), .ZN(n3739) );
  NAND2_X1 U11022 ( .A1(n1566), .A2(n24811), .ZN(n25107) );
  NAND2_X1 U11027 ( .A1(n12612), .A2(n25248), .ZN(n24811) );
  NAND2_X1 U11068 ( .A1(n23328), .A2(n23329), .ZN(n23331) );
  NAND2_X1 U11115 ( .A1(n1261), .A2(n15612), .ZN(n15861) );
  AND2_X1 U11128 ( .A1(n1147), .A2(n6690), .ZN(n1148) );
  OR2_X1 U11146 ( .A1(n13028), .A2(n302), .ZN(n2794) );
  NAND2_X1 U11162 ( .A1(n4445), .A2(n11974), .ZN(n24812) );
  NAND2_X1 U11170 ( .A1(n19478), .A2(n4667), .ZN(n17594) );
  XNOR2_X2 U11171 ( .A(n10), .B(n17591), .ZN(n19478) );
  OAI211_X2 U11184 ( .C1(n16982), .C2(n16983), .A(n16981), .B(n3982), .ZN(
        n18172) );
  NAND2_X1 U11185 ( .A1(n24813), .A2(n17551), .ZN(n17552) );
  OAI21_X1 U11188 ( .B1(n18927), .B2(n18967), .A(n356), .ZN(n24813) );
  NAND2_X1 U11198 ( .A1(n24169), .A2(n24171), .ZN(n3122) );
  NAND2_X1 U11205 ( .A1(n1689), .A2(n5101), .ZN(n2967) );
  NAND2_X1 U11208 ( .A1(n9231), .A2(n25457), .ZN(n5688) );
  NAND2_X1 U11209 ( .A1(n25103), .A2(n11065), .ZN(n11075) );
  XNOR2_X1 U11215 ( .A(n9143), .B(n24600), .ZN(n1466) );
  NAND2_X1 U11240 ( .A1(n20320), .A2(n20322), .ZN(n18992) );
  OAI21_X1 U11250 ( .B1(n10633), .B2(n11210), .A(n24814), .ZN(n4089) );
  NAND3_X1 U11257 ( .A1(n11210), .A2(n11338), .A3(n24082), .ZN(n24814) );
  NAND2_X1 U11299 ( .A1(n24495), .A2(n8839), .ZN(n10015) );
  NAND3_X2 U11314 ( .A1(n4650), .A2(n13464), .A3(n13465), .ZN(n14468) );
  OR2_X1 U11351 ( .A1(n15705), .A2(n16464), .ZN(n24855) );
  NAND3_X2 U11352 ( .A1(n24817), .A2(n24816), .A3(n9509), .ZN(n11396) );
  NAND3_X1 U11353 ( .A1(n4142), .A2(n5380), .A3(n11032), .ZN(n24816) );
  OAI21_X1 U11376 ( .B1(n20243), .B2(n20244), .A(n20242), .ZN(n24818) );
  NAND3_X2 U11385 ( .A1(n24819), .A2(n1113), .A3(n1114), .ZN(n17086) );
  NAND2_X1 U11411 ( .A1(n24821), .A2(n24820), .ZN(n24819) );
  NAND2_X1 U11462 ( .A1(n16469), .A2(n24551), .ZN(n24820) );
  AOI21_X1 U11481 ( .B1(n15546), .B2(n24822), .A(n383), .ZN(n24821) );
  NAND3_X2 U11491 ( .A1(n9728), .A2(n24824), .A3(n24823), .ZN(n11158) );
  NAND2_X1 U11495 ( .A1(n9726), .A2(n2922), .ZN(n24823) );
  NAND2_X1 U11506 ( .A1(n9725), .A2(n25043), .ZN(n24824) );
  NAND2_X1 U11516 ( .A1(n24826), .A2(n1365), .ZN(n24825) );
  XNOR2_X2 U11518 ( .A(n14632), .B(n14633), .ZN(n1365) );
  INV_X1 U11529 ( .A(n16073), .ZN(n24826) );
  OAI22_X2 U11549 ( .A1(n279), .A2(n19544), .B1(n19543), .B2(n19545), .ZN(
        n20368) );
  OAI21_X1 U11557 ( .B1(n5709), .B2(n13581), .A(n14107), .ZN(n24827) );
  OAI21_X1 U11567 ( .B1(n25388), .B2(n24829), .A(n24828), .ZN(n19717) );
  NAND2_X1 U11568 ( .A1(n25388), .A2(n339), .ZN(n24828) );
  NAND2_X1 U11587 ( .A1(n14150), .A2(n3717), .ZN(n14154) );
  NAND3_X2 U11589 ( .A1(n4860), .A2(n24258), .A3(n4964), .ZN(n3717) );
  NAND2_X1 U11593 ( .A1(n25480), .A2(n6480), .ZN(n6926) );
  NOR2_X1 U11617 ( .A1(n19850), .A2(n19660), .ZN(n20066) );
  NAND2_X1 U11665 ( .A1(n13188), .A2(n13187), .ZN(n13189) );
  XNOR2_X1 U11672 ( .A(n24830), .B(n23931), .ZN(Ciphertext[177]) );
  NAND3_X1 U11685 ( .A1(n24831), .A2(n23928), .A3(n23929), .ZN(n24830) );
  NAND2_X1 U11730 ( .A1(n24833), .A2(n4309), .ZN(n22507) );
  OAI21_X1 U11754 ( .B1(n4311), .B2(n5306), .A(n23425), .ZN(n24833) );
  NAND2_X1 U11757 ( .A1(n24834), .A2(n20616), .ZN(n20326) );
  NAND2_X1 U11779 ( .A1(n20084), .A2(n24835), .ZN(n24834) );
  NAND2_X1 U11783 ( .A1(n20571), .A2(n20614), .ZN(n20084) );
  NOR2_X2 U11795 ( .A1(n4577), .A2(n24836), .ZN(n11385) );
  AOI21_X1 U11821 ( .B1(n9580), .B2(n9581), .A(n11116), .ZN(n24836) );
  NAND2_X1 U11822 ( .A1(n513), .A2(n19662), .ZN(n2339) );
  NAND2_X1 U11826 ( .A1(n23469), .A2(n23499), .ZN(n23474) );
  NAND2_X1 U11828 ( .A1(n24837), .A2(n2713), .ZN(n22026) );
  NAND2_X1 U11833 ( .A1(n22019), .A2(n25438), .ZN(n24837) );
  OAI21_X1 U11838 ( .B1(n324), .B2(n4411), .A(n24838), .ZN(n4407) );
  NAND2_X1 U11841 ( .A1(n4412), .A2(n324), .ZN(n24838) );
  AND3_X2 U11853 ( .A1(n5240), .A2(n5241), .A3(n16797), .ZN(n16799) );
  NAND2_X1 U11868 ( .A1(n20269), .A2(n1155), .ZN(n1154) );
  OAI211_X1 U11871 ( .C1(n9503), .C2(n10104), .A(n24839), .B(n8644), .ZN(n9332) );
  NAND2_X1 U11874 ( .A1(n9503), .A2(n9775), .ZN(n24839) );
  INV_X1 U11938 ( .A(n16290), .ZN(n24841) );
  NAND2_X1 U11959 ( .A1(n9920), .A2(n9461), .ZN(n24843) );
  OAI211_X2 U11979 ( .C1(n20098), .C2(n20566), .A(n24109), .B(n24845), .ZN(
        n21520) );
  NAND3_X1 U12001 ( .A1(n24846), .A2(n3914), .A3(n3912), .ZN(n24112) );
  NAND3_X1 U12005 ( .A1(n3910), .A2(n3909), .A3(n23058), .ZN(n24846) );
  INV_X1 U12007 ( .A(n9921), .ZN(n24847) );
  OR2_X1 U12021 ( .A1(n9922), .A2(n9920), .ZN(n24848) );
  OAI21_X1 U12024 ( .B1(n16063), .B2(n16064), .A(n24849), .ZN(n15602) );
  NAND2_X1 U12028 ( .A1(n16064), .A2(n25446), .ZN(n24849) );
  OAI211_X2 U12033 ( .C1(n7107), .C2(n7250), .A(n24851), .B(n7106), .ZN(n8280)
         );
  NAND2_X1 U12051 ( .A1(n25211), .A2(n20042), .ZN(n19230) );
  NOR2_X1 U12083 ( .A1(n5800), .A2(n6964), .ZN(n6672) );
  OAI211_X1 U12099 ( .C1(n9919), .C2(n9354), .A(n24852), .B(n9355), .ZN(n9357)
         );
  NAND2_X1 U12100 ( .A1(n9919), .A2(n24853), .ZN(n24852) );
  OAI21_X1 U12108 ( .B1(n10199), .B2(n10200), .A(n13092), .ZN(n24854) );
  NAND2_X1 U12129 ( .A1(n10694), .A2(n11499), .ZN(n10331) );
  NAND2_X1 U12147 ( .A1(n23905), .A2(n21863), .ZN(n607) );
  NAND2_X1 U12170 ( .A1(n14000), .A2(n12668), .ZN(n14002) );
  NAND3_X1 U12276 ( .A1(n244), .A2(n707), .A3(n16427), .ZN(n17435) );
  NAND2_X1 U12277 ( .A1(n11211), .A2(n11342), .ZN(n24856) );
  NAND2_X1 U12280 ( .A1(n2071), .A2(n24857), .ZN(n14800) );
  NAND2_X1 U12465 ( .A1(n13734), .A2(n4979), .ZN(n24857) );
  NOR2_X2 U12492 ( .A1(n24858), .A2(n13980), .ZN(n15088) );
  OAI22_X1 U12512 ( .A1(n13977), .A2(n14439), .B1(n13978), .B2(n24713), .ZN(
        n24858) );
  OAI21_X1 U12535 ( .B1(n10020), .B2(n9730), .A(n24859), .ZN(n5372) );
  NAND2_X1 U12541 ( .A1(n9491), .A2(n10019), .ZN(n24859) );
  NOR2_X1 U12546 ( .A1(n16183), .A2(n25455), .ZN(n15916) );
  NAND2_X1 U12601 ( .A1(n15915), .A2(n15667), .ZN(n16183) );
  OAI21_X1 U12636 ( .B1(n7897), .B2(n24861), .A(n24860), .ZN(n7903) );
  NAND2_X1 U12684 ( .A1(n7897), .A2(n7898), .ZN(n24860) );
  NAND3_X1 U12701 ( .A1(n22812), .A2(n22656), .A3(n22813), .ZN(n2527) );
  NAND2_X1 U12739 ( .A1(n6394), .A2(n4178), .ZN(n4177) );
  NAND2_X1 U12770 ( .A1(n24862), .A2(n24354), .ZN(n2685) );
  INV_X1 U12773 ( .A(n20452), .ZN(n24862) );
  NAND2_X1 U12807 ( .A1(n1590), .A2(n20451), .ZN(n20452) );
  NAND3_X2 U12808 ( .A1(n3416), .A2(n3417), .A3(n3415), .ZN(n12306) );
  AOI21_X1 U12831 ( .B1(n15860), .B2(n15861), .A(n16113), .ZN(n24864) );
  NAND2_X1 U12847 ( .A1(n9936), .A2(n2971), .ZN(n2947) );
  NOR2_X1 U12900 ( .A1(n16572), .A2(n2580), .ZN(n24865) );
  OAI21_X1 U12983 ( .B1(n20669), .B2(n24567), .A(n24866), .ZN(n17311) );
  NAND2_X1 U12994 ( .A1(n20669), .A2(n20335), .ZN(n24866) );
  NAND2_X1 U13004 ( .A1(n24868), .A2(n24867), .ZN(n24019) );
  NAND2_X1 U13144 ( .A1(n22776), .A2(n22677), .ZN(n24867) );
  NAND2_X1 U13167 ( .A1(n22777), .A2(n24869), .ZN(n24868) );
  NAND2_X1 U13168 ( .A1(n2618), .A2(n2617), .ZN(n22777) );
  NAND2_X1 U13170 ( .A1(n10491), .A2(n11207), .ZN(n1225) );
  OAI21_X1 U13184 ( .B1(n20586), .B2(n3734), .A(n24870), .ZN(n5094) );
  NAND2_X1 U13185 ( .A1(n20586), .A2(n20593), .ZN(n24870) );
  XNOR2_X1 U13191 ( .A(n10719), .B(n24871), .ZN(n10745) );
  XNOR2_X1 U13192 ( .A(n24969), .B(n11295), .ZN(n24871) );
  XNOR2_X1 U13218 ( .A(n24872), .B(n18087), .ZN(n18090) );
  XNOR2_X1 U13245 ( .A(n18086), .B(n18085), .ZN(n24872) );
  NAND3_X1 U13303 ( .A1(n24281), .A2(n25181), .A3(n24873), .ZN(n25145) );
  NAND3_X1 U13441 ( .A1(n24875), .A2(n22737), .A3(n24874), .ZN(n22740) );
  NAND2_X1 U13456 ( .A1(n23495), .A2(n23483), .ZN(n24875) );
  NAND2_X1 U13468 ( .A1(n5063), .A2(n3442), .ZN(n12449) );
  NAND2_X1 U13480 ( .A1(n2539), .A2(n2997), .ZN(n2538) );
  BUF_X1 U13518 ( .A(n22939), .Z(n25063) );
  INV_X1 U13529 ( .A(n7733), .ZN(n25151) );
  OR2_X1 U13535 ( .A1(n13047), .A2(n13046), .ZN(n24876) );
  MUX2_X1 U13572 ( .A(n13043), .B(n13042), .S(n13041), .Z(n13047) );
  OR2_X1 U13600 ( .A1(n23632), .A2(n3164), .ZN(n23643) );
  XNOR2_X1 U13728 ( .A(n801), .B(n21740), .ZN(n24877) );
  XNOR2_X1 U13839 ( .A(n801), .B(n21740), .ZN(n22911) );
  OR2_X1 U13842 ( .A1(n15804), .A2(n15857), .ZN(n24171) );
  INV_X1 U13907 ( .A(n23420), .ZN(n142) );
  XNOR2_X1 U13937 ( .A(n20664), .B(n20663), .ZN(n24881) );
  XNOR2_X1 U13952 ( .A(n20664), .B(n20663), .ZN(n22389) );
  XNOR2_X1 U14046 ( .A(n24882), .B(n21993), .ZN(n22002) );
  XOR2_X1 U14151 ( .A(n1381), .B(n24986), .Z(n24882) );
  OR3_X1 U14229 ( .A1(n25474), .A2(n19345), .A3(n5280), .ZN(n5455) );
  XNOR2_X1 U14238 ( .A(n18140), .B(n18141), .ZN(n19107) );
  BUF_X1 U14261 ( .A(n23543), .Z(n24057) );
  OR2_X1 U14367 ( .A1(n20598), .A2(n20427), .ZN(n24883) );
  XNOR2_X1 U14532 ( .A(n21558), .B(n21557), .ZN(n24884) );
  XNOR2_X1 U14540 ( .A(n21558), .B(n21557), .ZN(n24885) );
  NAND2_X1 U14541 ( .A1(n835), .A2(n2854), .ZN(n20039) );
  NAND3_X1 U14561 ( .A1(n17458), .A2(n17459), .A3(n522), .ZN(n24886) );
  CLKBUF_X1 U14585 ( .A(n3016), .Z(n24887) );
  NAND3_X1 U14603 ( .A1(n17458), .A2(n17459), .A3(n522), .ZN(n18499) );
  AND2_X1 U14671 ( .A1(n16614), .A2(n16613), .ZN(n24888) );
  AOI21_X1 U14683 ( .B1(n21927), .B2(n21926), .A(n21925), .ZN(n23184) );
  XNOR2_X1 U14686 ( .A(n13371), .B(n13372), .ZN(n24890) );
  NAND2_X2 U14695 ( .A1(n19001), .A2(n2927), .ZN(n20536) );
  NOR2_X1 U14696 ( .A1(n24891), .A2(n24892), .ZN(n5768) );
  AND2_X1 U14697 ( .A1(n22922), .A2(n25070), .ZN(n24891) );
  NOR2_X1 U14704 ( .A1(n24379), .A2(n22922), .ZN(n24892) );
  XOR2_X1 U14705 ( .A(n18458), .B(n18568), .Z(n18118) );
  AND2_X1 U14706 ( .A1(n23146), .A2(n1349), .ZN(n23160) );
  OR2_X1 U14707 ( .A1(n22106), .A2(n22105), .ZN(n24893) );
  NAND4_X2 U14711 ( .A1(n21821), .A2(n21820), .A3(n21819), .A4(n21818), .ZN(
        n24895) );
  INV_X1 U14901 ( .A(n12583), .ZN(n12977) );
  NAND3_X1 U14928 ( .A1(n2363), .A2(n2362), .A3(n2360), .ZN(n24896) );
  NAND3_X1 U14939 ( .A1(n2363), .A2(n2362), .A3(n2360), .ZN(n21176) );
  OR2_X1 U14973 ( .A1(n24897), .A2(n20395), .ZN(n2425) );
  OR2_X1 U15011 ( .A1(n1327), .A2(n20384), .ZN(n24897) );
  NAND2_X1 U15128 ( .A1(n3563), .A2(n13485), .ZN(n4382) );
  NAND2_X1 U15155 ( .A1(n24155), .A2(n24154), .ZN(n21665) );
  OAI211_X1 U15173 ( .C1(n19945), .C2(n20960), .A(n19943), .B(n71), .ZN(n24899) );
  OAI211_X1 U15195 ( .C1(n19945), .C2(n20960), .A(n19943), .B(n71), .ZN(n21522) );
  XNOR2_X1 U15225 ( .A(n21083), .B(n21082), .ZN(n23997) );
  NOR2_X1 U15248 ( .A1(n19626), .A2(n19625), .ZN(n24469) );
  NAND2_X1 U15290 ( .A1(n21773), .A2(n2513), .ZN(n24901) );
  NAND2_X1 U15296 ( .A1(n21773), .A2(n2513), .ZN(n23594) );
  XNOR2_X1 U15300 ( .A(n20953), .B(n20952), .ZN(n24902) );
  NOR2_X1 U15306 ( .A1(n22405), .A2(n22404), .ZN(n24903) );
  NOR2_X1 U15315 ( .A1(n22405), .A2(n22404), .ZN(n24904) );
  XNOR2_X1 U15411 ( .A(n19903), .B(n19902), .ZN(n24905) );
  AND3_X1 U15429 ( .A1(n23805), .A2(n22043), .A3(n21828), .ZN(n21907) );
  NAND2_X1 U15464 ( .A1(n21377), .A2(n3080), .ZN(n24906) );
  NAND2_X1 U15535 ( .A1(n1587), .A2(n1585), .ZN(n24907) );
  XNOR2_X1 U15538 ( .A(n17754), .B(n17753), .ZN(n24908) );
  XNOR2_X1 U15546 ( .A(n17754), .B(n17753), .ZN(n24909) );
  NAND2_X1 U15565 ( .A1(n4633), .A2(n21549), .ZN(n24911) );
  NAND2_X1 U15620 ( .A1(n4633), .A2(n21549), .ZN(n23372) );
  INV_X1 U15621 ( .A(n23066), .ZN(n25179) );
  XNOR2_X1 U15678 ( .A(n17035), .B(n17034), .ZN(n19310) );
  INV_X1 U15690 ( .A(n11191), .ZN(n24913) );
  AOI22_X1 U15694 ( .A1(n10271), .A2(n11185), .B1(n11184), .B2(n10731), .ZN(
        n11370) );
  AND3_X1 U15695 ( .A1(n22277), .A2(n22276), .A3(n1507), .ZN(n24914) );
  NOR3_X1 U15714 ( .A1(n20349), .A2(n19654), .A3(n20670), .ZN(n19655) );
  NOR2_X1 U15806 ( .A1(n19656), .A2(n19655), .ZN(n24916) );
  NOR2_X1 U15813 ( .A1(n19656), .A2(n19655), .ZN(n21521) );
  CLKBUF_X1 U15831 ( .A(Key[98]), .Z(n2735) );
  XOR2_X1 U15839 ( .A(n10880), .B(n11602), .Z(n10882) );
  AND2_X1 U15912 ( .A1(n22800), .A2(n22799), .ZN(n25161) );
  OR2_X1 U15984 ( .A1(n17500), .A2(n17499), .ZN(n24917) );
  OAI211_X1 U16147 ( .C1(n22356), .C2(n21785), .A(n21784), .B(n21783), .ZN(
        n24921) );
  OAI211_X1 U16259 ( .C1(n22356), .C2(n21785), .A(n21784), .B(n21783), .ZN(
        n23757) );
  XOR2_X1 U16297 ( .A(n21586), .B(n21585), .Z(n24922) );
  AND3_X1 U16307 ( .A1(n22679), .A2(n22774), .A3(n5377), .ZN(n24923) );
  NAND2_X1 U16351 ( .A1(n22682), .A2(n22681), .ZN(n24924) );
  INV_X1 U16502 ( .A(n20264), .ZN(n20410) );
  AND2_X1 U16716 ( .A1(n19446), .A2(n19351), .ZN(n24926) );
  XOR2_X1 U16755 ( .A(n7472), .B(n7473), .Z(n24927) );
  XNOR2_X1 U16762 ( .A(n14693), .B(n14692), .ZN(n24928) );
  XNOR2_X1 U16769 ( .A(n18216), .B(n18217), .ZN(n24929) );
  XNOR2_X1 U16831 ( .A(n18216), .B(n18217), .ZN(n19184) );
  BUF_X2 U16847 ( .A(n23869), .Z(n23902) );
  XNOR2_X1 U16850 ( .A(n10565), .B(n10566), .ZN(n24930) );
  XOR2_X1 U16852 ( .A(n17761), .B(n17760), .Z(n24931) );
  XNOR2_X1 U16854 ( .A(n10565), .B(n10566), .ZN(n12719) );
  XNOR2_X1 U16856 ( .A(n21620), .B(n21619), .ZN(n24932) );
  BUF_X1 U16862 ( .A(n23391), .Z(n24933) );
  XNOR2_X1 U16903 ( .A(n21620), .B(n21619), .ZN(n22940) );
  OR3_X1 U16924 ( .A1(n24470), .A2(n10935), .A3(n10505), .ZN(n10598) );
  AOI21_X1 U16928 ( .B1(n23890), .B2(n23904), .A(n25239), .ZN(n21866) );
  INV_X1 U16930 ( .A(n16597), .ZN(n24935) );
  NAND2_X1 U16967 ( .A1(n3465), .A2(n3932), .ZN(n24936) );
  NAND2_X1 U16968 ( .A1(n3465), .A2(n3932), .ZN(n20792) );
  NAND4_X1 U16969 ( .A1(n13706), .A2(n13704), .A3(n13705), .A4(n13707), .ZN(
        n24937) );
  NAND4_X1 U16971 ( .A1(n13706), .A2(n13704), .A3(n13705), .A4(n13707), .ZN(
        n24938) );
  NAND4_X1 U17021 ( .A1(n13706), .A2(n13704), .A3(n13705), .A4(n13707), .ZN(
        n15040) );
  INV_X1 U17023 ( .A(n20414), .ZN(n25108) );
  AND2_X1 U17083 ( .A1(n3810), .A2(n3809), .ZN(n20578) );
  NAND2_X1 U17084 ( .A1(n5583), .A2(n5582), .ZN(n24941) );
  AND2_X1 U17101 ( .A1(n14), .A2(n25165), .ZN(n24942) );
  CLKBUF_X1 U17106 ( .A(n4052), .Z(n24943) );
  XOR2_X1 U17226 ( .A(n6222), .B(n6221), .Z(n24944) );
  NOR2_X1 U17238 ( .A1(n7214), .A2(n7213), .ZN(n24946) );
  NOR2_X1 U17239 ( .A1(n7214), .A2(n7213), .ZN(n8781) );
  BUF_X1 U17240 ( .A(n23410), .Z(n24947) );
  OR2_X1 U17260 ( .A1(n21148), .A2(n21149), .ZN(n25024) );
  MUX2_X1 U17288 ( .A(n22372), .B(n22371), .S(n22680), .Z(n23939) );
  OAI211_X1 U17336 ( .C1(n18726), .C2(n19376), .A(n18725), .B(n4317), .ZN(
        n20181) );
  INV_X1 U17347 ( .A(n20126), .ZN(n25101) );
  INV_X1 U17355 ( .A(n9874), .ZN(n307) );
  NOR2_X1 U17357 ( .A1(n20136), .A2(n20019), .ZN(n24950) );
  XNOR2_X1 U17381 ( .A(n20705), .B(n20704), .ZN(n24951) );
  XNOR2_X1 U17382 ( .A(n20705), .B(n20704), .ZN(n22566) );
  INV_X1 U17385 ( .A(n23120), .ZN(n24952) );
  OR2_X2 U17386 ( .A1(n19899), .A2(n19898), .ZN(n21621) );
  XOR2_X1 U17391 ( .A(n21264), .B(n21263), .Z(n24953) );
  NAND3_X1 U17452 ( .A1(n22795), .A2(n22797), .A3(n22796), .ZN(n24954) );
  NAND3_X1 U17527 ( .A1(n22795), .A2(n22797), .A3(n22796), .ZN(n24006) );
  NOR2_X1 U17569 ( .A1(n20721), .A2(n20720), .ZN(n24955) );
  OAI21_X1 U17570 ( .B1(n5620), .B2(n14415), .A(n13859), .ZN(n24956) );
  OAI21_X1 U17571 ( .B1(n5620), .B2(n14415), .A(n13859), .ZN(n15478) );
  NAND4_X1 U17572 ( .A1(n8575), .A2(n8572), .A3(n8574), .A4(n8573), .ZN(n11169) );
  INV_X1 U17634 ( .A(n14849), .ZN(n24958) );
  XNOR2_X1 U17635 ( .A(n7241), .B(n7240), .ZN(n24959) );
  XNOR2_X1 U17720 ( .A(n7241), .B(n7240), .ZN(n2585) );
  XNOR2_X1 U17754 ( .A(n13641), .B(n13642), .ZN(n24960) );
  XNOR2_X1 U17872 ( .A(n18305), .B(n24961), .ZN(n18119) );
  XOR2_X1 U17889 ( .A(n18675), .B(n1856), .Z(n24961) );
  AOI21_X1 U17890 ( .B1(n19671), .B2(n18887), .A(n18886), .ZN(n24962) );
  XNOR2_X1 U17963 ( .A(n21118), .B(n21119), .ZN(n24963) );
  AOI21_X1 U18075 ( .B1(n19671), .B2(n18887), .A(n18886), .ZN(n21597) );
  OAI21_X2 U18111 ( .B1(n12497), .B2(n12496), .A(n12495), .ZN(n14377) );
  NAND4_X1 U18136 ( .A1(n10266), .A2(n10265), .A3(n10267), .A4(n10264), .ZN(
        n24964) );
  XNOR2_X1 U18205 ( .A(n667), .B(n11763), .ZN(n24965) );
  NAND4_X1 U18245 ( .A1(n10266), .A2(n10265), .A3(n10267), .A4(n10264), .ZN(
        n12383) );
  XNOR2_X1 U18289 ( .A(n667), .B(n11763), .ZN(n12569) );
  AND2_X1 U18326 ( .A1(n14685), .A2(n14686), .ZN(n24966) );
  XNOR2_X1 U18365 ( .A(n11972), .B(n11973), .ZN(n24346) );
  NAND3_X1 U18367 ( .A1(n4352), .A2(n3476), .A3(n4349), .ZN(n24967) );
  XNOR2_X1 U18466 ( .A(n17793), .B(n17794), .ZN(n24968) );
  NOR2_X1 U18634 ( .A1(n1169), .A2(n10723), .ZN(n24969) );
  NOR2_X1 U18636 ( .A1(n1169), .A2(n10723), .ZN(n24970) );
  NOR2_X1 U18645 ( .A1(n1169), .A2(n10723), .ZN(n12138) );
  XNOR2_X1 U18670 ( .A(n20694), .B(n20693), .ZN(n24971) );
  XNOR2_X1 U18673 ( .A(n20694), .B(n20693), .ZN(n22564) );
  AND2_X1 U18675 ( .A1(n2117), .A2(n2116), .ZN(n24973) );
  NAND2_X1 U18690 ( .A1(n4015), .A2(n1836), .ZN(n24975) );
  INV_X1 U18747 ( .A(n23411), .ZN(n24977) );
  INV_X1 U18771 ( .A(n23411), .ZN(n24978) );
  OAI211_X1 U18836 ( .C1(n9279), .C2(n9649), .A(n9648), .B(n9647), .ZN(n24980)
         );
  INV_X1 U18847 ( .A(n15696), .ZN(n24981) );
  OAI211_X1 U18848 ( .C1(n9279), .C2(n9649), .A(n9648), .B(n9647), .ZN(n11782)
         );
  XNOR2_X1 U18849 ( .A(n18488), .B(n18487), .ZN(n24982) );
  NAND2_X1 U18868 ( .A1(n4434), .A2(n23001), .ZN(n24983) );
  XNOR2_X1 U18879 ( .A(n18488), .B(n18487), .ZN(n19057) );
  XOR2_X1 U18953 ( .A(n8425), .B(n8424), .Z(n24984) );
  OAI21_X1 U18959 ( .B1(n200), .B2(n19927), .A(n19926), .ZN(n24985) );
  OAI21_X1 U18961 ( .B1(n200), .B2(n19927), .A(n19926), .ZN(n24986) );
  OAI21_X1 U18986 ( .B1(n200), .B2(n19927), .A(n19926), .ZN(n21992) );
  OAI21_X1 U18988 ( .B1(n22856), .B2(n22855), .A(n22854), .ZN(n23410) );
  INV_X1 U18996 ( .A(n12218), .ZN(n24987) );
  AND3_X1 U19000 ( .A1(n10214), .A2(n10213), .A3(n4327), .ZN(n12261) );
  NOR2_X1 U19023 ( .A1(n3411), .A2(n22803), .ZN(n25159) );
  XNOR2_X1 U19040 ( .A(n11844), .B(n11843), .ZN(n24988) );
  OR2_X1 U19041 ( .A1(n22489), .A2(n22488), .ZN(n24989) );
  XNOR2_X1 U19049 ( .A(n11844), .B(n11843), .ZN(n13279) );
  INV_X1 U19055 ( .A(n11242), .ZN(n12152) );
  XOR2_X1 U19080 ( .A(n25396), .B(n11289), .Z(n24990) );
  INV_X1 U19082 ( .A(n997), .ZN(n24991) );
  INV_X1 U19084 ( .A(n24559), .ZN(n25115) );
  CLKBUF_X1 U19085 ( .A(n22805), .Z(n24992) );
  NOR2_X1 U19133 ( .A1(n22477), .A2(n22476), .ZN(n24993) );
  XNOR2_X1 U19184 ( .A(n21235), .B(n21234), .ZN(n22805) );
  INV_X1 U19186 ( .A(n6529), .ZN(n24994) );
  INV_X1 U19205 ( .A(n13088), .ZN(n24995) );
  CLKBUF_X1 U19210 ( .A(n6060), .Z(n6734) );
  XOR2_X1 U19277 ( .A(n18484), .B(n18356), .Z(n17994) );
  NAND4_X1 U19284 ( .A1(n20305), .A2(n5764), .A3(n20304), .A4(n20303), .ZN(
        n24996) );
  NAND4_X1 U19307 ( .A1(n20305), .A2(n5764), .A3(n20304), .A4(n20303), .ZN(
        n21569) );
  OAI211_X1 U19313 ( .C1(n22179), .C2(n24369), .A(n22177), .B(n22178), .ZN(
        n2305) );
  NAND2_X1 U19316 ( .A1(n10395), .A2(n10394), .ZN(n24999) );
  NAND3_X1 U19327 ( .A1(n1269), .A2(n15635), .A3(n15636), .ZN(n25000) );
  BUF_X1 U19338 ( .A(n19595), .Z(n25001) );
  XNOR2_X1 U19355 ( .A(n18029), .B(n18030), .ZN(n19595) );
  XNOR2_X1 U19363 ( .A(n797), .B(n17677), .ZN(n25002) );
  OAI21_X1 U19417 ( .B1(n16168), .B2(n16167), .A(n16166), .ZN(n25003) );
  OAI21_X1 U19418 ( .B1(n16168), .B2(n16167), .A(n16166), .ZN(n17195) );
  XOR2_X1 U19459 ( .A(n8844), .B(n8577), .Z(n8582) );
  BUF_X1 U19491 ( .A(n23332), .Z(n25004) );
  XNOR2_X1 U19492 ( .A(n21410), .B(n21411), .ZN(n23332) );
  XOR2_X1 U19564 ( .A(n8767), .B(n8768), .Z(n25005) );
  XNOR2_X1 U19567 ( .A(n18660), .B(n18611), .ZN(n25006) );
  XNOR2_X1 U19568 ( .A(n5255), .B(n8441), .ZN(n7146) );
  XOR2_X1 U19615 ( .A(n8811), .B(n8810), .Z(n25007) );
  AOI22_X1 U19641 ( .A1(n13570), .A2(n13571), .B1(n13572), .B2(n13573), .ZN(
        n25008) );
  XNOR2_X1 U19682 ( .A(n15157), .B(n15158), .ZN(n25009) );
  AOI22_X1 U19696 ( .A1(n13570), .A2(n13571), .B1(n13572), .B2(n13573), .ZN(
        n14488) );
  XNOR2_X1 U19787 ( .A(n15157), .B(n15158), .ZN(n16267) );
  INV_X1 U19788 ( .A(n2216), .ZN(n25010) );
  XNOR2_X1 U19793 ( .A(n17778), .B(n2029), .ZN(n4114) );
  INV_X1 U19832 ( .A(n20036), .ZN(n22233) );
  BUF_X1 U19880 ( .A(n13643), .Z(n25011) );
  OAI211_X1 U19882 ( .C1(n13060), .C2(n3065), .A(n13059), .B(n13058), .ZN(
        n13643) );
  XNOR2_X1 U19883 ( .A(n18511), .B(n18510), .ZN(n25012) );
  OAI211_X1 U19888 ( .C1(n3889), .C2(n13804), .A(n13803), .B(n13802), .ZN(
        n25013) );
  XNOR2_X1 U19895 ( .A(n14641), .B(n14640), .ZN(n15802) );
  XNOR2_X1 U19902 ( .A(n5864), .B(Key[24]), .ZN(n25014) );
  CLKBUF_X1 U19909 ( .A(n12607), .Z(n25015) );
  OAI211_X1 U19956 ( .C1(n22675), .C2(n22674), .A(n22673), .B(n22672), .ZN(
        n25017) );
  NOR2_X1 U19957 ( .A1(n8663), .A2(n8662), .ZN(n11840) );
  OAI211_X1 U19995 ( .C1(n25208), .C2(n25128), .A(n14240), .B(n25127), .ZN(
        n2741) );
  XNOR2_X1 U19997 ( .A(n20931), .B(n20930), .ZN(n25018) );
  XNOR2_X1 U20000 ( .A(n20931), .B(n20930), .ZN(n22208) );
  OAI211_X1 U20022 ( .C1(n14125), .C2(n3851), .A(n3849), .B(n3850), .ZN(n25019) );
  OAI211_X1 U20097 ( .C1(n14125), .C2(n3851), .A(n3849), .B(n3850), .ZN(n15480) );
  XNOR2_X1 U20100 ( .A(n9035), .B(n5014), .ZN(n25020) );
  INV_X1 U20149 ( .A(n15164), .ZN(n2765) );
  XOR2_X1 U20188 ( .A(n8110), .B(n8111), .Z(n25021) );
  XNOR2_X1 U20225 ( .A(n21125), .B(n21124), .ZN(n25022) );
  XNOR2_X1 U20245 ( .A(n21125), .B(n21124), .ZN(n25023) );
  AOI21_X1 U20248 ( .B1(n5517), .B2(n5519), .A(n4871), .ZN(n11209) );
  OAI211_X1 U20249 ( .C1(n10818), .C2(n10817), .A(n3594), .B(n3595), .ZN(
        n25027) );
  OAI211_X1 U20496 ( .C1(n10818), .C2(n10817), .A(n3594), .B(n3595), .ZN(
        n12112) );
  NOR2_X1 U20510 ( .A1(n25029), .A2(n17568), .ZN(n25028) );
  AND2_X1 U20588 ( .A1(n17566), .A2(n20317), .ZN(n25029) );
  OAI21_X2 U20634 ( .B1(n18970), .B2(n17553), .A(n17552), .ZN(n19889) );
  XNOR2_X1 U20643 ( .A(n14700), .B(n14701), .ZN(n25030) );
  INV_X1 U20657 ( .A(n15631), .ZN(n25031) );
  XNOR2_X1 U20675 ( .A(n14700), .B(n14701), .ZN(n15782) );
  NOR3_X1 U20684 ( .A1(n14058), .A2(n13521), .A3(n14054), .ZN(n13522) );
  XNOR2_X1 U20694 ( .A(n10640), .B(n10639), .ZN(n25033) );
  OR2_X1 U20704 ( .A1(n17714), .A2(n17713), .ZN(n25034) );
  XOR2_X1 U20731 ( .A(n11798), .B(n11799), .Z(n11802) );
  AOI22_X1 U20738 ( .A1(n14074), .A2(n14078), .B1(n13852), .B2(n14077), .ZN(
        n25036) );
  AOI22_X1 U20739 ( .A1(n14074), .A2(n14078), .B1(n13852), .B2(n14077), .ZN(
        n13491) );
  AND3_X1 U20747 ( .A1(n24277), .A2(n24276), .A3(n6029), .ZN(n25037) );
  INV_X1 U20749 ( .A(n16602), .ZN(n25038) );
  NAND2_X1 U20761 ( .A1(n16604), .A2(n25038), .ZN(n25039) );
  OAI21_X1 U20817 ( .B1(n19877), .B2(n25221), .A(n19876), .ZN(n25040) );
  OAI21_X1 U20846 ( .B1(n19877), .B2(n25221), .A(n19876), .ZN(n21133) );
  NOR2_X1 U20919 ( .A1(n22489), .A2(n22488), .ZN(n25042) );
  NOR2_X1 U20987 ( .A1(n22489), .A2(n22488), .ZN(n23441) );
  XNOR2_X1 U20995 ( .A(n8608), .B(n8607), .ZN(n25043) );
  XNOR2_X1 U20996 ( .A(n8608), .B(n8607), .ZN(n10007) );
  XNOR2_X1 U21022 ( .A(n5991), .B(Key[104]), .ZN(n25044) );
  XNOR2_X1 U21027 ( .A(n5991), .B(Key[104]), .ZN(n25045) );
  XNOR2_X1 U21028 ( .A(n5991), .B(Key[104]), .ZN(n6602) );
  XNOR2_X1 U21037 ( .A(n8326), .B(n5619), .ZN(n25046) );
  INV_X1 U21041 ( .A(n4931), .ZN(n25047) );
  XOR2_X1 U21048 ( .A(n12260), .B(n12221), .Z(n25048) );
  XOR2_X1 U21102 ( .A(n11327), .B(n11326), .Z(n25049) );
  CLKBUF_X1 U21105 ( .A(n22214), .Z(n25050) );
  OAI21_X1 U21108 ( .B1(n21790), .B2(n22222), .A(n2734), .ZN(n25051) );
  XNOR2_X1 U21112 ( .A(n21323), .B(n21322), .ZN(n22214) );
  OAI21_X1 U21123 ( .B1(n21790), .B2(n22222), .A(n2734), .ZN(n23770) );
  XNOR2_X1 U21124 ( .A(n17746), .B(n17747), .ZN(n25052) );
  XNOR2_X1 U21134 ( .A(n17746), .B(n17747), .ZN(n19217) );
  XNOR2_X1 U21149 ( .A(n3205), .B(n3204), .ZN(n25053) );
  INV_X1 U21176 ( .A(n3662), .ZN(n25054) );
  XNOR2_X1 U21209 ( .A(n3205), .B(n3204), .ZN(n13358) );
  CLKBUF_X1 U21223 ( .A(n23441), .Z(n23450) );
  CLKBUF_X1 U21251 ( .A(n23464), .Z(n25055) );
  XNOR2_X1 U21252 ( .A(n13576), .B(n13577), .ZN(n16200) );
  XNOR2_X1 U21271 ( .A(n18231), .B(n18230), .ZN(n25057) );
  XNOR2_X1 U21280 ( .A(n18231), .B(n18230), .ZN(n19548) );
  NOR2_X1 U21291 ( .A1(n22571), .A2(n21938), .ZN(n25059) );
  NOR2_X1 U21298 ( .A1(n22571), .A2(n21938), .ZN(n23186) );
  MUX2_X1 U21357 ( .A(n19380), .B(n17980), .S(n19378), .Z(n3518) );
  XNOR2_X1 U21376 ( .A(n11656), .B(n11655), .ZN(n25061) );
  OAI211_X1 U21388 ( .C1(n24077), .C2(n19941), .A(n2946), .B(n679), .ZN(n25062) );
  OAI211_X1 U21394 ( .C1(n24077), .C2(n19941), .A(n2946), .B(n679), .ZN(n21312) );
  XNOR2_X2 U21395 ( .A(n11636), .B(n11635), .ZN(n12490) );
  XNOR2_X1 U21424 ( .A(n8300), .B(n8299), .ZN(n25064) );
  OAI211_X1 U21467 ( .C1(n19639), .C2(n347), .A(n19638), .B(n19637), .ZN(
        n25065) );
  OAI211_X1 U21534 ( .C1(n19639), .C2(n347), .A(n19638), .B(n19637), .ZN(
        n21640) );
  XNOR2_X1 U21537 ( .A(n21155), .B(n21156), .ZN(n25066) );
  XNOR2_X1 U21545 ( .A(n21155), .B(n21156), .ZN(n22317) );
  XOR2_X1 U21546 ( .A(n17979), .B(n17978), .Z(n25067) );
  XOR2_X1 U21547 ( .A(n21131), .B(n21130), .Z(n25068) );
  XNOR2_X1 U21571 ( .A(n8156), .B(n8155), .ZN(n25069) );
  XNOR2_X1 U21581 ( .A(n8156), .B(n8155), .ZN(n9885) );
  OR2_X1 U21582 ( .A1(n23155), .A2(n23154), .ZN(n23147) );
  XNOR2_X1 U21596 ( .A(n20998), .B(n20997), .ZN(n25070) );
  XNOR2_X1 U21615 ( .A(n20998), .B(n20997), .ZN(n22928) );
  NOR2_X1 U21660 ( .A1(n840), .A2(n22112), .ZN(n23546) );
  OAI21_X1 U21826 ( .B1(n9840), .B2(n10099), .A(n9839), .ZN(n25074) );
  XNOR2_X1 U21924 ( .A(n20441), .B(n20440), .ZN(n25075) );
  INV_X1 U21927 ( .A(n878), .ZN(n25076) );
  XNOR2_X1 U21937 ( .A(n20441), .B(n20440), .ZN(n22657) );
  OAI21_X1 U21944 ( .B1(n4470), .B2(n4469), .A(n481), .ZN(n23972) );
  XOR2_X1 U22007 ( .A(n20891), .B(n20890), .Z(n25078) );
  XNOR2_X2 U22099 ( .A(n10392), .B(n11284), .ZN(n12652) );
  XNOR2_X1 U22120 ( .A(n21089), .B(n21090), .ZN(n25079) );
  XNOR2_X1 U22146 ( .A(n21089), .B(n21090), .ZN(n23996) );
  XOR2_X1 U22185 ( .A(n4996), .B(n4995), .Z(n25080) );
  XNOR2_X1 U22188 ( .A(n21426), .B(n21425), .ZN(n25081) );
  XNOR2_X1 U22197 ( .A(n21426), .B(n21425), .ZN(n23336) );
  XOR2_X1 U22223 ( .A(n20083), .B(n20082), .Z(n25082) );
  AOI21_X1 U22245 ( .B1(n782), .B2(n22362), .A(n1249), .ZN(n25083) );
  AOI21_X1 U22281 ( .B1(n782), .B2(n22362), .A(n1249), .ZN(n25084) );
  AOI21_X1 U22301 ( .B1(n782), .B2(n22362), .A(n1249), .ZN(n23940) );
  INV_X1 U22340 ( .A(n18883), .ZN(n25086) );
  XNOR2_X1 U22354 ( .A(n11418), .B(n11417), .ZN(n12795) );
  OAI211_X1 U22372 ( .C1(n10610), .C2(n9610), .A(n9609), .B(n9608), .ZN(n25087) );
  NOR2_X1 U22396 ( .A1(n18787), .A2(n18786), .ZN(n25088) );
  NOR2_X1 U22405 ( .A1(n18787), .A2(n18786), .ZN(n25089) );
  OAI211_X1 U22412 ( .C1(n10610), .C2(n9610), .A(n9609), .B(n9608), .ZN(n12143) );
  NOR2_X1 U22428 ( .A1(n19685), .A2(n21066), .ZN(n25091) );
  NOR2_X1 U22429 ( .A1(n19685), .A2(n21066), .ZN(n21997) );
  XNOR2_X1 U22430 ( .A(n13476), .B(n13475), .ZN(n25092) );
  NAND4_X2 U22444 ( .A1(n4780), .A2(n19844), .A3(n25094), .A4(n25093), .ZN(
        n21974) );
  NAND2_X1 U22455 ( .A1(n1205), .A2(n3198), .ZN(n25093) );
  NAND2_X1 U22516 ( .A1(n1206), .A2(n24194), .ZN(n25094) );
  NAND3_X1 U22540 ( .A1(n4116), .A2(n13935), .A3(n13200), .ZN(n13202) );
  NAND3_X1 U22578 ( .A1(n10142), .A2(n9821), .A3(n24026), .ZN(n9822) );
  NAND2_X1 U22628 ( .A1(n9918), .A2(n9462), .ZN(n9912) );
  AND2_X1 U22675 ( .A1(n5376), .A2(n16795), .ZN(n4553) );
  NOR2_X1 U22680 ( .A1(n12767), .A2(n13217), .ZN(n12809) );
  XNOR2_X2 U22682 ( .A(n11236), .B(n11235), .ZN(n12767) );
  NAND2_X1 U22713 ( .A1(n25095), .A2(n1170), .ZN(n1169) );
  NAND2_X1 U22728 ( .A1(n1167), .A2(n1166), .ZN(n25095) );
  NAND2_X1 U22736 ( .A1(n24927), .A2(n9965), .ZN(n1602) );
  AOI21_X1 U22760 ( .B1(n6608), .B2(n6112), .A(n6714), .ZN(n5786) );
  NAND2_X1 U22804 ( .A1(n6232), .A2(n6715), .ZN(n6608) );
  NAND2_X1 U22807 ( .A1(n5033), .A2(n1491), .ZN(n5028) );
  NAND3_X1 U22848 ( .A1(n5035), .A2(n24941), .A3(n5037), .ZN(n5033) );
  OR2_X1 U22849 ( .A1(n5800), .A2(n6575), .ZN(n4755) );
  OAI21_X1 U22850 ( .B1(n25097), .B2(n13266), .A(n25096), .ZN(n12681) );
  NAND2_X1 U22879 ( .A1(n13266), .A2(n13264), .ZN(n25096) );
  INV_X1 U22887 ( .A(n24443), .ZN(n25097) );
  NAND2_X1 U22908 ( .A1(n12705), .A2(n25098), .ZN(n14960) );
  NAND2_X1 U22924 ( .A1(n25099), .A2(n177), .ZN(n25098) );
  INV_X1 U22971 ( .A(n16351), .ZN(n25100) );
  NAND2_X1 U22975 ( .A1(n16350), .A2(n25100), .ZN(n25165) );
  NAND3_X1 U22979 ( .A1(n19675), .A2(n25102), .A3(n25101), .ZN(n4570) );
  NAND2_X1 U23002 ( .A1(n20130), .A2(n20546), .ZN(n25102) );
  NAND2_X1 U23017 ( .A1(n13518), .A2(n1355), .ZN(n13610) );
  NOR2_X2 U23018 ( .A1(n2706), .A2(n25104), .ZN(n20460) );
  OAI22_X1 U23029 ( .A1(n19385), .A2(n24908), .B1(n19391), .B2(n5196), .ZN(
        n25104) );
  XNOR2_X1 U23043 ( .A(n20700), .B(n20701), .ZN(n20867) );
  NAND3_X1 U23058 ( .A1(n17735), .A2(n17730), .A3(n17486), .ZN(n16815) );
  NAND3_X1 U23060 ( .A1(n16746), .A2(n17279), .A3(n17277), .ZN(n16747) );
  NAND3_X1 U23084 ( .A1(n18714), .A2(n19351), .A3(n19451), .ZN(n25105) );
  NAND2_X1 U23100 ( .A1(n5162), .A2(n7237), .ZN(n8980) );
  NAND3_X1 U23110 ( .A1(n1984), .A2(n5163), .A3(n1345), .ZN(n5162) );
  NAND2_X1 U23123 ( .A1(n25106), .A2(n17164), .ZN(n687) );
  INV_X1 U23127 ( .A(n16836), .ZN(n25106) );
  NAND2_X1 U23128 ( .A1(n4775), .A2(n17165), .ZN(n16836) );
  AOI22_X2 U23145 ( .A1(n3547), .A2(n16172), .B1(n16174), .B2(n16173), .ZN(
        n17192) );
  NAND2_X1 U23150 ( .A1(n25107), .A2(n13307), .ZN(n1564) );
  NAND2_X1 U23153 ( .A1(n16056), .A2(n4972), .ZN(n16059) );
  NAND2_X1 U23241 ( .A1(n25110), .A2(n25109), .ZN(n11224) );
  NAND2_X1 U23243 ( .A1(n11222), .A2(n13137), .ZN(n25109) );
  NAND2_X1 U23247 ( .A1(n25112), .A2(n25111), .ZN(n25110) );
  INV_X1 U23295 ( .A(n13137), .ZN(n25111) );
  NAND2_X1 U23299 ( .A1(n11142), .A2(n12437), .ZN(n25112) );
  NAND3_X1 U23310 ( .A1(n19558), .A2(n19555), .A3(n3284), .ZN(n4261) );
  NAND2_X1 U23345 ( .A1(n25114), .A2(n25113), .ZN(n22589) );
  NAND2_X1 U23347 ( .A1(n22582), .A2(n24561), .ZN(n25113) );
  NAND2_X1 U23356 ( .A1(n22583), .A2(n25115), .ZN(n25114) );
  NAND3_X1 U23367 ( .A1(n5250), .A2(n6904), .A3(n5249), .ZN(n5248) );
  NAND3_X2 U23398 ( .A1(n7058), .A2(n25118), .A3(n25117), .ZN(n9044) );
  NAND2_X1 U23416 ( .A1(n3248), .A2(n7809), .ZN(n25118) );
  NAND2_X1 U23417 ( .A1(n21829), .A2(n22219), .ZN(n22162) );
  NAND2_X1 U23418 ( .A1(n2788), .A2(n6968), .ZN(n7065) );
  NAND3_X1 U23420 ( .A1(n13950), .A2(n3069), .A3(n13949), .ZN(n1836) );
  NAND3_X1 U23424 ( .A1(n24195), .A2(n15628), .A3(n15629), .ZN(n15631) );
  NAND2_X1 U23428 ( .A1(n25005), .A2(n9977), .ZN(n9416) );
  NAND2_X1 U23432 ( .A1(n25250), .A2(n10556), .ZN(n10657) );
  NAND2_X1 U23457 ( .A1(n9745), .A2(n9990), .ZN(n25119) );
  AOI21_X1 U23473 ( .B1(n25121), .B2(n24534), .A(n9991), .ZN(n25120) );
  AOI21_X1 U23474 ( .B1(n9351), .B2(n9460), .A(n1470), .ZN(n9358) );
  NAND2_X1 U23515 ( .A1(n118), .A2(n119), .ZN(n18129) );
  NAND3_X1 U23613 ( .A1(n13325), .A2(n12952), .A3(n13329), .ZN(n12847) );
  AND3_X2 U23625 ( .A1(n5501), .A2(n4363), .A3(n1458), .ZN(n20507) );
  NAND2_X1 U23679 ( .A1(n22292), .A2(n25122), .ZN(n23252) );
  NAND2_X1 U23693 ( .A1(n25124), .A2(n25123), .ZN(n25122) );
  INV_X1 U23764 ( .A(n22293), .ZN(n25124) );
  NAND2_X1 U23865 ( .A1(n25126), .A2(n25125), .ZN(n20283) );
  NAND2_X1 U23867 ( .A1(n20282), .A2(n20281), .ZN(n25125) );
  NAND2_X1 U23962 ( .A1(n4460), .A2(n24414), .ZN(n25126) );
  NAND2_X1 U23963 ( .A1(n25208), .A2(n14244), .ZN(n25127) );
  NAND2_X1 U24024 ( .A1(n5760), .A2(n17122), .ZN(n25129) );
  NAND2_X1 U24078 ( .A1(n19486), .A2(n25440), .ZN(n25130) );
  OAI21_X1 U24111 ( .B1(n19806), .B2(n20235), .A(n25132), .ZN(n19807) );
  NAND3_X1 U24131 ( .A1(n19804), .A2(n25205), .A3(n20170), .ZN(n25132) );
  XNOR2_X1 U24143 ( .A(n22014), .B(n21522), .ZN(n20795) );
  NAND2_X1 U24167 ( .A1(n14510), .A2(n14439), .ZN(n13978) );
  MUX2_X1 U24177 ( .A(n4273), .B(n22655), .S(n25075), .Z(n22658) );
  NAND2_X1 U24181 ( .A1(n7528), .A2(n7527), .ZN(n25133) );
  NAND2_X1 U24204 ( .A1(n3934), .A2(n10364), .ZN(n25135) );
  NAND2_X1 U24205 ( .A1(n9595), .A2(n10129), .ZN(n7440) );
  OAI22_X1 U24206 ( .A1(n10254), .A2(n24959), .B1(n5057), .B2(n9211), .ZN(
        n9595) );
  OR2_X1 U24207 ( .A1(n12433), .A2(n12455), .ZN(n12730) );
  XNOR2_X1 U24209 ( .A(n8206), .B(n8753), .ZN(n25136) );
  XNOR2_X1 U24210 ( .A(n8204), .B(n8205), .ZN(n25137) );
  NAND3_X1 U24211 ( .A1(n22233), .A2(n3231), .A3(n22235), .ZN(n1164) );
  AOI22_X2 U24212 ( .A1(n6167), .A2(n127), .B1(n6166), .B2(n6542), .ZN(n7761)
         );
  INV_X1 U24213 ( .A(n17330), .ZN(n15559) );
  NAND2_X1 U24214 ( .A1(n3553), .A2(n16309), .ZN(n17330) );
  XNOR2_X1 U24217 ( .A(n18198), .B(n18476), .ZN(n18109) );
  NAND3_X2 U24218 ( .A1(n16747), .A2(n16764), .A3(n24299), .ZN(n18198) );
  NAND2_X1 U24219 ( .A1(n21367), .A2(n4350), .ZN(n25138) );
  AND3_X2 U24220 ( .A1(n3188), .A2(n5843), .A3(n5842), .ZN(n7313) );
  NAND2_X1 U24221 ( .A1(n11678), .A2(n11677), .ZN(n24165) );
  NAND3_X1 U24222 ( .A1(n15557), .A2(n24297), .A3(n16012), .ZN(n634) );
  NAND2_X1 U24223 ( .A1(n1152), .A2(n25139), .ZN(n1150) );
  XNOR2_X1 U24225 ( .A(n17804), .B(n17805), .ZN(n25140) );
  NAND2_X1 U24226 ( .A1(n11170), .A2(n11169), .ZN(n10313) );
  NAND3_X1 U24227 ( .A1(n17242), .A2(n17346), .A3(n17241), .ZN(n16136) );
  NAND2_X1 U24229 ( .A1(n22883), .A2(n24879), .ZN(n25141) );
  INV_X1 U24230 ( .A(n22882), .ZN(n25142) );
  AND3_X2 U24231 ( .A1(n1262), .A2(n1264), .A3(n5558), .ZN(n12214) );
  NAND2_X1 U24232 ( .A1(n25143), .A2(n5478), .ZN(n5477) );
  NAND2_X1 U24233 ( .A1(n5480), .A2(n19270), .ZN(n25143) );
  NAND2_X1 U24234 ( .A1(n10616), .A2(n10412), .ZN(n24521) );
  NAND3_X1 U24235 ( .A1(n25144), .A2(n4852), .A3(n4851), .ZN(n20360) );
  NAND2_X1 U24236 ( .A1(n4314), .A2(n1212), .ZN(n25144) );
  XNOR2_X1 U24237 ( .A(n25145), .B(n24280), .ZN(Ciphertext[190]) );
  NAND3_X1 U24238 ( .A1(n262), .A2(n24927), .A3(n9281), .ZN(n25146) );
  NAND2_X1 U24239 ( .A1(n25147), .A2(n9505), .ZN(n11032) );
  XNOR2_X1 U24241 ( .A(n15350), .B(n15190), .ZN(n14490) );
  NAND2_X1 U24242 ( .A1(n9361), .A2(n25148), .ZN(n10757) );
  NAND2_X1 U24243 ( .A1(n24237), .A2(n22842), .ZN(n24236) );
  OAI21_X2 U24245 ( .B1(n15627), .B2(n16097), .A(n25149), .ZN(n17059) );
  NAND2_X1 U24246 ( .A1(n15864), .A2(n15626), .ZN(n25149) );
  NAND3_X1 U24247 ( .A1(n1548), .A2(n2462), .A3(n2463), .ZN(n19924) );
  OR2_X1 U24250 ( .A1(n17439), .A2(n16962), .ZN(n2550) );
  OAI21_X1 U24251 ( .B1(n7735), .B2(n25151), .A(n25150), .ZN(n6251) );
  NAND2_X1 U24252 ( .A1(n7735), .A2(n7642), .ZN(n25150) );
  NAND3_X1 U24253 ( .A1(n14381), .A2(n14382), .A3(n16154), .ZN(n14396) );
  NAND3_X2 U24254 ( .A1(n25152), .A2(n7669), .A3(n7668), .ZN(n8673) );
  NOR2_X2 U24255 ( .A1(n13457), .A2(n25153), .ZN(n14477) );
  OAI22_X1 U24256 ( .A1(n13454), .A2(n24711), .B1(n13889), .B2(n24710), .ZN(
        n25153) );
  NAND2_X1 U24257 ( .A1(n7222), .A2(n7474), .ZN(n1531) );
  NAND2_X1 U24258 ( .A1(n3362), .A2(n7421), .ZN(n7222) );
  NAND2_X1 U24259 ( .A1(n6050), .A2(n6630), .ZN(n6750) );
  XNOR2_X2 U24260 ( .A(Key[75]), .B(Plaintext[75]), .ZN(n6630) );
  XNOR2_X1 U24261 ( .A(n18628), .B(n16037), .ZN(n16091) );
  NAND2_X1 U24263 ( .A1(n20142), .A2(n4066), .ZN(n20141) );
  NAND2_X1 U24264 ( .A1(n7460), .A2(n268), .ZN(n7467) );
  NAND2_X1 U24265 ( .A1(n10903), .A2(n10445), .ZN(n10443) );
  NAND2_X1 U24266 ( .A1(n10904), .A2(n10746), .ZN(n10903) );
  NAND2_X1 U24267 ( .A1(n10654), .A2(n10660), .ZN(n10399) );
  NOR2_X1 U24268 ( .A1(n13234), .A2(n13298), .ZN(n1445) );
  INV_X1 U24269 ( .A(n7881), .ZN(n25154) );
  NAND2_X1 U24270 ( .A1(n8013), .A2(n8012), .ZN(n8019) );
  NAND2_X1 U24271 ( .A1(n2376), .A2(n2679), .ZN(n2394) );
  NAND2_X1 U24272 ( .A1(n25156), .A2(n25155), .ZN(n10455) );
  NAND2_X1 U24273 ( .A1(n10756), .A2(n10451), .ZN(n25155) );
  NAND2_X1 U24274 ( .A1(n20510), .A2(n20215), .ZN(n20508) );
  NAND2_X1 U24275 ( .A1(n19188), .A2(n19187), .ZN(n25157) );
  NAND2_X1 U24276 ( .A1(n19189), .A2(n19550), .ZN(n25158) );
  NAND2_X1 U24277 ( .A1(n24051), .A2(n6232), .ZN(n6607) );
  AOI21_X1 U24278 ( .B1(n25161), .B2(n25160), .A(n25159), .ZN(n21389) );
  NAND2_X1 U24279 ( .A1(n11178), .A2(n11175), .ZN(n10939) );
  NAND2_X1 U24280 ( .A1(n17040), .A2(n17364), .ZN(n25162) );
  NAND2_X1 U24281 ( .A1(n2469), .A2(n2470), .ZN(n2468) );
  INV_X1 U24283 ( .A(n10088), .ZN(n25164) );
  NAND2_X1 U24284 ( .A1(n14), .A2(n25165), .ZN(n16980) );
  NAND2_X1 U24285 ( .A1(n15992), .A2(n15654), .ZN(n15660) );
  XNOR2_X1 U24286 ( .A(n25166), .B(n12375), .ZN(n11463) );
  NAND2_X2 U24287 ( .A1(n10765), .A2(n734), .ZN(n12375) );
  NAND2_X1 U24288 ( .A1(n11301), .A2(n11298), .ZN(n10435) );
  NAND2_X1 U24289 ( .A1(n6906), .A2(n6905), .ZN(n6787) );
  OAI21_X1 U24290 ( .B1(n1340), .B2(n25168), .A(n25167), .ZN(n22654) );
  NAND2_X1 U24291 ( .A1(n22652), .A2(n1340), .ZN(n25167) );
  INV_X1 U24292 ( .A(n22653), .ZN(n25168) );
  NOR2_X1 U24293 ( .A1(n22311), .A2(n25169), .ZN(n22312) );
  NAND2_X1 U24294 ( .A1(n3095), .A2(n3097), .ZN(n25169) );
  NAND2_X1 U24295 ( .A1(n25172), .A2(n25170), .ZN(n20392) );
  NAND2_X1 U24296 ( .A1(n352), .A2(n19345), .ZN(n25170) );
  NAND2_X1 U24297 ( .A1(n20387), .A2(n25440), .ZN(n25172) );
  NAND2_X1 U24299 ( .A1(n25173), .A2(n392), .ZN(n599) );
  NAND2_X1 U24300 ( .A1(n1), .A2(n3), .ZN(n25173) );
  NAND2_X1 U24301 ( .A1(n665), .A2(n25174), .ZN(n608) );
  NAND3_X2 U24303 ( .A1(n952), .A2(n951), .A3(n18857), .ZN(n19849) );
  NAND2_X1 U24304 ( .A1(n25175), .A2(n593), .ZN(n22405) );
  NAND3_X1 U24306 ( .A1(n24239), .A2(n22905), .A3(n22904), .ZN(n24238) );
  OR2_X2 U24307 ( .A1(n13668), .A2(n13670), .ZN(n14000) );
  NAND3_X1 U24308 ( .A1(n16727), .A2(n16726), .A3(n16725), .ZN(n16728) );
  NAND2_X1 U24309 ( .A1(n22464), .A2(n22462), .ZN(n21932) );
  OR2_X1 U24311 ( .A1(n14122), .A2(n13811), .ZN(n3849) );
  NAND2_X1 U24312 ( .A1(n14123), .A2(n14208), .ZN(n14122) );
  NAND3_X1 U24313 ( .A1(n1231), .A2(n5705), .A3(n5707), .ZN(n24269) );
  NAND2_X1 U24314 ( .A1(n25176), .A2(n576), .ZN(n19604) );
  NAND2_X1 U24315 ( .A1(n19600), .A2(n19601), .ZN(n25176) );
  NAND3_X1 U24317 ( .A1(n23079), .A2(n25178), .A3(n25177), .ZN(n21281) );
  NAND2_X1 U24318 ( .A1(n23066), .A2(n22578), .ZN(n25177) );
  NAND2_X1 U24319 ( .A1(n25179), .A2(n23064), .ZN(n25178) );
  NAND3_X1 U24320 ( .A1(n3037), .A2(n23188), .A3(n23189), .ZN(n3036) );
  NAND2_X1 U24321 ( .A1(n19361), .A2(n19211), .ZN(n1266) );
  NOR2_X1 U24322 ( .A1(n16273), .A2(n16274), .ZN(n25180) );
  NAND2_X1 U24323 ( .A1(n24204), .A2(n24019), .ZN(n25181) );
  NAND2_X1 U24324 ( .A1(n6538), .A2(n6530), .ZN(n6130) );
  OR3_X1 U24325 ( .A1(n10682), .A2(n2306), .A3(n9769), .ZN(n8031) );
  OAI211_X1 U24326 ( .C1(n4232), .C2(n4234), .A(n25182), .B(n4231), .ZN(
        Ciphertext[34]) );
  NAND2_X1 U24327 ( .A1(n4229), .A2(n4236), .ZN(n25182) );
  NAND2_X1 U24328 ( .A1(n1158), .A2(n1146), .ZN(n25183) );
  NAND2_X1 U24329 ( .A1(n1890), .A2(n25469), .ZN(n18785) );
  NAND2_X1 U24331 ( .A1(n4694), .A2(n6051), .ZN(n25185) );
  NAND2_X1 U24332 ( .A1(n6449), .A2(n6450), .ZN(n25186) );
  NAND2_X1 U24333 ( .A1(n25), .A2(n25064), .ZN(n25188) );
  NAND2_X1 U24334 ( .A1(n10172), .A2(n9814), .ZN(n25189) );
  INV_X1 U24338 ( .A(n11873), .ZN(n25191) );
  NAND2_X1 U24339 ( .A1(n12899), .A2(n24988), .ZN(n13284) );
  OAI21_X1 U24340 ( .B1(n1331), .B2(n14127), .A(n25192), .ZN(n14134) );
  NAND2_X1 U24341 ( .A1(n1331), .A2(n25193), .ZN(n25192) );
  INV_X1 U24342 ( .A(n14126), .ZN(n25193) );
  XNOR2_X1 U24343 ( .A(n8311), .B(n8312), .ZN(n10168) );
  XNOR2_X2 U24344 ( .A(n7472), .B(n7473), .ZN(n9468) );
  NAND4_X2 U10040 ( .A1(n3870), .A2(n3867), .A3(n10238), .A4(n3869), .ZN(
        n11582) );
  OR2_X2 U3424 ( .A1(n2962), .A2(n2963), .ZN(n10891) );
  NAND3_X2 U2253 ( .A1(n3524), .A2(n4992), .A3(n3523), .ZN(n13614) );
  OAI211_X2 U20847 ( .C1(n20235), .C2(n20173), .A(n20172), .B(n20171), .ZN(
        n21998) );
  BUF_X2 U1019 ( .A(n7850), .Z(n24072) );
  NAND4_X2 U786 ( .A1(n2534), .A2(n2533), .A3(n5917), .A4(n7104), .ZN(n7350)
         );
  BUF_X1 U1457 ( .A(n16423), .Z(n1329) );
  BUF_X2 U3043 ( .A(n9365), .Z(n10146) );
  INV_X2 U1115 ( .A(n5522), .ZN(n3374) );
  NAND2_X2 U3445 ( .A1(n2136), .A2(n2135), .ZN(n21332) );
  NAND3_X2 U6597 ( .A1(n2622), .A2(n6215), .A3(n6214), .ZN(n8935) );
  NAND2_X2 U1209 ( .A1(n24183), .A2(n2399), .ZN(n11301) );
  AND3_X2 U8646 ( .A1(n4743), .A2(n1416), .A3(n4742), .ZN(n3703) );
  NAND2_X2 U2551 ( .A1(n4803), .A2(n4799), .ZN(n8691) );
  AND2_X2 U8824 ( .A1(n10257), .A2(n10259), .ZN(n10728) );
  NAND2_X2 U3015 ( .A1(n594), .A2(n19617), .ZN(n20448) );
  OAI211_X2 U2385 ( .C1(n10679), .C2(n2984), .A(n4815), .B(n1401), .ZN(n11717)
         );
  BUF_X1 U18822 ( .A(n19987), .Z(n24979) );
  BUF_X1 U2113 ( .A(n15714), .Z(n16471) );
  NAND3_X2 U24194 ( .A1(n2250), .A2(n14627), .A3(n14626), .ZN(n17273) );
  BUF_X1 U24157 ( .A(n13386), .Z(n24507) );
  XNOR2_X2 U1819 ( .A(n15878), .B(n15879), .ZN(n19133) );
  XNOR2_X2 U1750 ( .A(n20978), .B(n20977), .ZN(n22166) );
  AND2_X2 U755 ( .A1(n4415), .A2(n13489), .ZN(n15191) );
  OAI211_X2 U1232 ( .C1(n14586), .C2(n14747), .A(n1675), .B(n1674), .ZN(n2285)
         );
  BUF_X2 U1647 ( .A(n14100), .Z(n24376) );
  XNOR2_X2 U506 ( .A(n12329), .B(n12328), .ZN(n13350) );
  AND2_X2 U1004 ( .A1(n22414), .A2(n22413), .ZN(n23305) );
  NOR2_X2 U1989 ( .A1(n17124), .A2(n17123), .ZN(n17958) );
  NAND4_X2 U9301 ( .A1(n13430), .A2(n13431), .A3(n14069), .A4(n13429), .ZN(
        n14799) );
  CLKBUF_X3 U1839 ( .A(n17567), .Z(n20322) );
  NAND2_X2 U1879 ( .A1(n18799), .A2(n18798), .ZN(n20062) );
  NOR2_X2 U1953 ( .A1(n16979), .A2(n17450), .ZN(n17449) );
  AND2_X2 U17681 ( .A1(n1305), .A2(n1308), .ZN(n20174) );
  MUX2_X2 U709 ( .A(n7979), .B(n7978), .S(n7977), .Z(n8069) );
  AND2_X2 U1877 ( .A1(n3683), .A2(n1476), .ZN(n18310) );
  BUF_X1 U21457 ( .A(n21140), .Z(n24406) );
  XNOR2_X2 U12294 ( .A(n5880), .B(Key[34]), .ZN(n6952) );
  MUX2_X2 U1215 ( .A(n8712), .B(n8711), .S(n9985), .Z(n11529) );
  AND3_X2 U185 ( .A1(n3136), .A2(n3137), .A3(n3135), .ZN(n22578) );
  OAI21_X2 U21731 ( .B1(n20623), .B2(n20622), .A(n20621), .ZN(n21630) );
  AND3_X2 U10086 ( .A1(n8139), .A2(n8138), .A3(n8137), .ZN(n10993) );
  NAND4_X2 U576 ( .A1(n7547), .A2(n7544), .A3(n7546), .A4(n7545), .ZN(n9075)
         );
  BUF_X1 U510 ( .A(n17313), .Z(n24543) );
  AND2_X2 U1191 ( .A1(n3085), .A2(n4824), .ZN(n15044) );
  OR2_X2 U675 ( .A1(n9303), .A2(n9304), .ZN(n10713) );
  XNOR2_X2 U1189 ( .A(n14862), .B(n14863), .ZN(n16219) );
  INV_X2 U2404 ( .A(n10952), .ZN(n2754) );
  AND3_X2 U21492 ( .A1(n20153), .A2(n20152), .A3(n20151), .ZN(n21138) );
  OAI22_X2 U17263 ( .A1(n13481), .A2(n13480), .B1(n13479), .B2(n13801), .ZN(
        n14827) );
  NAND3_X2 U6023 ( .A1(n16909), .A2(n24632), .A3(n2583), .ZN(n18582) );
  BUF_X1 U3618 ( .A(n18761), .Z(n19532) );
  AND3_X2 U824 ( .A1(n17848), .A2(n17847), .A3(n17846), .ZN(n19887) );
  AND3_X2 U149 ( .A1(n17218), .A2(n17219), .A3(n17217), .ZN(n18187) );
  OAI211_X2 U160 ( .C1(n17609), .C2(n16564), .A(n16563), .B(n16562), .ZN(
        n18269) );
  OAI211_X2 U2006 ( .C1(n17054), .C2(n16935), .A(n16934), .B(n16933), .ZN(
        n18067) );
  XNOR2_X1 U22322 ( .A(n11919), .B(n11918), .ZN(n12688) );
  AND2_X2 U1708 ( .A1(n25130), .A2(n25131), .ZN(n20231) );
  OAI211_X2 U985 ( .C1(n16299), .C2(n15024), .A(n15022), .B(n24777), .ZN(
        n17408) );
  OR2_X2 U721 ( .A1(n5868), .A2(n5869), .ZN(n7232) );
  OAI22_X2 U2213 ( .A1(n13599), .A2(n5520), .B1(n13962), .B2(n13598), .ZN(
        n15430) );
  BUF_X1 U2681 ( .A(n6770), .Z(n6909) );
  AND4_X2 U2025 ( .A1(n1701), .A2(n1703), .A3(n1702), .A4(n1705), .ZN(n18157)
         );
  OR2_X2 U488 ( .A1(n19027), .A2(n19026), .ZN(n20142) );
  BUF_X1 U3586 ( .A(n19310), .Z(n24912) );
  NAND2_X2 U23390 ( .A1(n15930), .A2(n25116), .ZN(n17051) );
  MUX2_X2 U593 ( .A(n11021), .B(n11020), .S(n24640), .Z(n13775) );
  NAND3_X2 U1988 ( .A1(n3396), .A2(n5225), .A3(n3395), .ZN(n18375) );
  NOR2_X2 U3659 ( .A1(n21354), .A2(n21353), .ZN(n23817) );
  AND3_X2 U3582 ( .A1(n9254), .A2(n9252), .A3(n9253), .ZN(n10861) );
  AND3_X2 U1064 ( .A1(n19892), .A2(n3541), .A3(n3540), .ZN(n20697) );
  AND2_X2 U2100 ( .A1(n15633), .A2(n3592), .ZN(n17054) );
  XNOR2_X1 U5036 ( .A(n1759), .B(n17815), .ZN(n19457) );
  XNOR2_X2 U2142 ( .A(n14175), .B(n14174), .ZN(n17183) );
  NAND2_X2 U9454 ( .A1(n2158), .A2(n12603), .ZN(n14849) );
  OAI21_X2 U2073 ( .B1(n16315), .B2(n16314), .A(n16313), .ZN(n17351) );
  XNOR2_X2 U2327 ( .A(n11514), .B(n11513), .ZN(n12774) );
  OR3_X2 U1147 ( .A1(n20068), .A2(n19849), .A3(n19660), .ZN(n210) );
  NAND2_X2 U2005 ( .A1(n15876), .A2(n4614), .ZN(n18294) );
  OR2_X2 U2058 ( .A1(n6283), .A2(n6282), .ZN(n7801) );
  BUF_X1 U851 ( .A(n23742), .Z(n24063) );
  NAND2_X2 U2922 ( .A1(n25133), .A2(n7530), .ZN(n8790) );
  NOR2_X2 U1434 ( .A1(n17437), .A2(n3000), .ZN(n17439) );
  AND3_X2 U1810 ( .A1(n2365), .A2(n2371), .A3(n2366), .ZN(n21599) );
  NAND3_X2 U505 ( .A1(n7411), .A2(n4277), .A3(n4278), .ZN(n9015) );
  AND3_X2 U606 ( .A1(n19287), .A2(n19285), .A3(n19286), .ZN(n20401) );
  MUX2_X2 U2087 ( .A(n16144), .B(n16143), .S(n16416), .Z(n17399) );
  BUF_X1 U2293 ( .A(n12560), .Z(n13015) );
  OR2_X2 U14 ( .A1(n19790), .A2(n5338), .ZN(n21141) );
  AND2_X2 U1870 ( .A1(n18898), .A2(n2844), .ZN(n20126) );
  AND3_X2 U5897 ( .A1(n24148), .A2(n9631), .A3(n9630), .ZN(n11342) );
  BUF_X2 U12061 ( .A(n19353), .Z(n19451) );
  XNOR2_X1 U523 ( .A(n4504), .B(n14844), .ZN(n16221) );
  XNOR2_X1 U2349 ( .A(n11663), .B(n11664), .ZN(n13061) );
  AOI21_X1 U2161 ( .B1(n6735), .B2(n6736), .A(n6734), .ZN(n6867) );
  NAND2_X2 U1685 ( .A1(n493), .A2(n3454), .ZN(n13521) );
  NAND2_X2 U6643 ( .A1(n13471), .A2(n1770), .ZN(n15488) );
  AND2_X2 U19056 ( .A1(n19056), .A2(n19057), .ZN(n19576) );
  AND2_X2 U18623 ( .A1(n203), .A2(n530), .ZN(n12122) );
  BUF_X2 U300 ( .A(n13360), .Z(n24552) );
  INV_X1 U1214 ( .A(n10767), .ZN(n11085) );
  NAND3_X2 U7603 ( .A1(n5489), .A2(n7586), .A3(n5490), .ZN(n8782) );
  AND3_X2 U556 ( .A1(n15942), .A2(n3437), .A3(n2771), .ZN(n17053) );
  BUF_X1 U21354 ( .A(n11519), .Z(n25060) );
  NAND3_X2 U7665 ( .A1(n2224), .A2(n7127), .A3(n3898), .ZN(n8755) );
  BUF_X2 U1072 ( .A(n12510), .Z(n12742) );
  BUF_X1 U495 ( .A(n16284), .Z(n24539) );
  NOR2_X2 U1984 ( .A1(n4565), .A2(n4562), .ZN(n18579) );
  AND2_X2 U492 ( .A1(n1115), .A2(n15551), .ZN(n16649) );
  XNOR2_X2 U2538 ( .A(n9014), .B(n9013), .ZN(n10027) );
  NAND4_X2 U1469 ( .A1(n5564), .A2(n5563), .A3(n5565), .A4(n20925), .ZN(n21523) );
  NAND2_X2 U2582 ( .A1(n2080), .A2(n7988), .ZN(n9158) );
  NAND4_X2 U472 ( .A1(n5206), .A2(n5209), .A3(n20196), .A4(n5205), .ZN(n21043)
         );
  XNOR2_X1 U4779 ( .A(n20886), .B(n20885), .ZN(n22887) );
  XNOR2_X1 U804 ( .A(Key[54]), .B(Plaintext[54]), .ZN(n6975) );
  CLKBUF_X1 U13601 ( .A(Key[99]), .Z(n3164) );
  CLKBUF_X1 U789 ( .A(Key[35]), .Z(n4711) );
  CLKBUF_X1 U1597 ( .A(Key[157]), .Z(n1776) );
  CLKBUF_X1 U1247 ( .A(Key[28]), .Z(n2050) );
  CLKBUF_X1 U1633 ( .A(Key[152]), .Z(n2903) );
  XNOR2_X1 U12248 ( .A(Key[153]), .B(Plaintext[153]), .ZN(n6874) );
  XNOR2_X1 U1063 ( .A(Key[114]), .B(Plaintext[114]), .ZN(n7026) );
  XNOR2_X1 U4226 ( .A(Key[165]), .B(Plaintext[165]), .ZN(n6775) );
  CLKBUF_X1 U1240 ( .A(Key[2]), .Z(n23883) );
  XNOR2_X1 U936 ( .A(n5968), .B(Key[175]), .ZN(n6426) );
  INV_X1 U12566 ( .A(n6905), .ZN(n6089) );
  OR2_X1 U426 ( .A1(n6987), .A2(n6119), .ZN(n6642) );
  XNOR2_X1 U792 ( .A(n5789), .B(Key[88]), .ZN(n6622) );
  XNOR2_X1 U1131 ( .A(n5877), .B(Key[30]), .ZN(n6529) );
  XNOR2_X1 U12308 ( .A(n5886), .B(Key[40]), .ZN(n6683) );
  XNOR2_X1 U1249 ( .A(n5892), .B(Key[48]), .ZN(n6556) );
  XNOR2_X1 U12384 ( .A(n5944), .B(Key[181]), .ZN(n6297) );
  XNOR2_X1 U152 ( .A(n5962), .B(Key[164]), .ZN(n6292) );
  XNOR2_X1 U354 ( .A(n6025), .B(Key[15]), .ZN(n6519) );
  BUF_X1 U2680 ( .A(n5835), .Z(n6793) );
  OR2_X1 U9169 ( .A1(n4696), .A2(n5774), .ZN(n6053) );
  INV_X1 U282 ( .A(n5794), .ZN(n6722) );
  INV_X1 U1235 ( .A(n1698), .ZN(n5451) );
  OR2_X1 U4806 ( .A1(n6198), .A2(n6292), .ZN(n6922) );
  OR2_X1 U5174 ( .A1(n6519), .A2(n6179), .ZN(n6518) );
  OAI21_X1 U2632 ( .B1(n2496), .B2(n6578), .A(n2495), .ZN(n7533) );
  OAI211_X1 U343 ( .C1(n3763), .C2(n6940), .A(n4826), .B(n6681), .ZN(n7358) );
  AND3_X1 U2748 ( .A1(n773), .A2(n6462), .A3(n6461), .ZN(n7688) );
  OR2_X1 U6515 ( .A1(n6300), .A2(n6299), .ZN(n7862) );
  NAND2_X1 U2662 ( .A1(n5977), .A2(n5978), .ZN(n7890) );
  OR2_X1 U7342 ( .A1(n5270), .A2(n6472), .ZN(n7917) );
  OAI21_X1 U268 ( .B1(n6278), .B2(n6279), .A(n791), .ZN(n7166) );
  NAND2_X1 U921 ( .A1(n2149), .A2(n2025), .ZN(n8219) );
  INV_X1 U88 ( .A(n7638), .ZN(n7918) );
  OR2_X1 U952 ( .A1(n6417), .A2(n6416), .ZN(n7857) );
  NAND2_X1 U2031 ( .A1(n77), .A2(n703), .ZN(n7255) );
  NAND2_X1 U3087 ( .A1(n6981), .A2(n6980), .ZN(n7477) );
  NOR2_X1 U2629 ( .A1(n5648), .A2(n2836), .ZN(n7973) );
  OR2_X1 U112 ( .A1(n6022), .A2(n2166), .ZN(n7595) );
  MUX2_X1 U12707 ( .A(n6270), .B(n6269), .S(n6136), .Z(n7800) );
  INV_X1 U2649 ( .A(n7351), .ZN(n7346) );
  INV_X1 U1017 ( .A(n7883), .ZN(n7582) );
  AND2_X1 U566 ( .A1(n6851), .A2(n6850), .ZN(n7983) );
  INV_X1 U1230 ( .A(n8367), .ZN(n24577) );
  AND2_X1 U1100 ( .A1(n6149), .A2(n6148), .ZN(n7619) );
  OR2_X1 U2643 ( .A1(n2784), .A2(n6202), .ZN(n8012) );
  NAND2_X1 U2635 ( .A1(n1750), .A2(n4321), .ZN(n7230) );
  NAND3_X1 U480 ( .A1(n2786), .A2(n6079), .A3(n6080), .ZN(n7292) );
  OR2_X1 U1099 ( .A1(n7087), .A2(n7211), .ZN(n7663) );
  BUF_X1 U773 ( .A(n7211), .Z(n8528) );
  INV_X1 U13063 ( .A(n7065), .ZN(n7952) );
  OR2_X1 U5194 ( .A1(n5468), .A2(n7349), .ZN(n7107) );
  AND3_X1 U8484 ( .A1(n5329), .A2(n7417), .A3(n7416), .ZN(n8119) );
  OR3_X1 U2566 ( .A1(n3259), .A2(n4206), .A3(n7533), .ZN(n2883) );
  OAI211_X1 U228 ( .C1(n7289), .C2(n7288), .A(n7287), .B(n7286), .ZN(n8798) );
  AND2_X1 U2559 ( .A1(n3345), .A2(n6495), .ZN(n8960) );
  OAI211_X1 U4007 ( .C1(n1124), .C2(n199), .A(n2092), .B(n5050), .ZN(n8928) );
  AOI22_X1 U13406 ( .A1(n7470), .A2(n7884), .B1(n7469), .B2(n7313), .ZN(n9045)
         );
  OAI211_X1 U1037 ( .C1(n7122), .C2(n7338), .A(n1904), .B(n7121), .ZN(n5179)
         );
  OAI211_X1 U2639 ( .C1(n7903), .C2(n7902), .A(n7899), .B(n7900), .ZN(n8796)
         );
  OAI211_X1 U6640 ( .C1(n6098), .C2(n7755), .A(n2521), .B(n1769), .ZN(n8674)
         );
  AND2_X1 U986 ( .A1(n7407), .A2(n7408), .ZN(n8476) );
  OR2_X1 U652 ( .A1(n7270), .A2(n7269), .ZN(n8989) );
  AND2_X1 U491 ( .A1(n7679), .A2(n7678), .ZN(n8116) );
  OAI21_X1 U409 ( .B1(n7321), .B2(n7320), .A(n2768), .ZN(n8959) );
  OAI21_X1 U197 ( .B1(n5204), .B2(n2522), .A(n5203), .ZN(n5014) );
  BUF_X1 U622 ( .A(n8627), .Z(n24547) );
  OAI21_X1 U6214 ( .B1(n7337), .B2(n7464), .A(n6763), .ZN(n9140) );
  NAND3_X1 U1951 ( .A1(n3082), .A2(n24205), .A3(n3083), .ZN(n8682) );
  OAI21_X1 U21801 ( .B1(n5116), .B2(n7952), .A(n2490), .ZN(n24413) );
  NAND4_X1 U7618 ( .A1(n7871), .A2(n7872), .A3(n7870), .A4(n7869), .ZN(n9179)
         );
  AND2_X1 U2553 ( .A1(n5548), .A2(n5547), .ZN(n9011) );
  XNOR2_X1 U13964 ( .A(n8345), .B(n8970), .ZN(n8725) );
  AND3_X1 U103 ( .A1(n5053), .A2(n5055), .A3(n6010), .ZN(n8951) );
  NAND2_X1 U2789 ( .A1(n472), .A2(n7194), .ZN(n8772) );
  OAI211_X1 U6484 ( .C1(n6319), .C2(n4536), .A(n24652), .B(n24648), .ZN(n8945)
         );
  NAND2_X1 U1079 ( .A1(n7072), .A2(n3814), .ZN(n8923) );
  XNOR2_X1 U1118 ( .A(n3307), .B(n8272), .ZN(n9805) );
  XNOR2_X1 U2527 ( .A(n8743), .B(n8742), .ZN(n9231) );
  BUF_X1 U2433 ( .A(n9893), .Z(n227) );
  XNOR2_X1 U2513 ( .A(n8957), .B(n8958), .ZN(n10044) );
  XNOR2_X1 U14249 ( .A(n8695), .B(n8694), .ZN(n9980) );
  BUF_X1 U625 ( .A(n9874), .Z(n24549) );
  BUF_X1 U823 ( .A(n9856), .Z(n9558) );
  XNOR2_X1 U289 ( .A(n1906), .B(n8665), .ZN(n10082) );
  BUF_X1 U534 ( .A(n9454), .Z(n9887) );
  BUF_X1 U1306 ( .A(n9962), .Z(n262) );
  MUX2_X1 U10264 ( .A(n9063), .B(n5004), .S(n10053), .Z(n9088) );
  OAI21_X1 U14990 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n10971) );
  NAND2_X1 U2625 ( .A1(n9540), .A2(n4594), .ZN(n10751) );
  AND2_X1 U474 ( .A1(n8144), .A2(n8143), .ZN(n10405) );
  OAI21_X1 U15059 ( .B1(n10076), .B2(n10075), .A(n10074), .ZN(n11063) );
  NAND3_X1 U23311 ( .A1(n9283), .A2(n9284), .A3(n25146), .ZN(n2243) );
  OAI211_X1 U2445 ( .C1(n9880), .C2(n9879), .A(n9878), .B(n9877), .ZN(n10968)
         );
  OAI21_X1 U494 ( .B1(n9265), .B2(n9899), .A(n9264), .ZN(n10736) );
  BUF_X1 U2535 ( .A(n8934), .Z(n11524) );
  OAI21_X1 U1838 ( .B1(n2564), .B2(n3134), .A(n9213), .ZN(n10590) );
  OAI22_X1 U1112 ( .A1(n8030), .A2(n9937), .B1(n8029), .B2(n24511), .ZN(n10682) );
  AND3_X1 U787 ( .A1(n9785), .A2(n9784), .A3(n9783), .ZN(n11009) );
  MUX2_X1 U13694 ( .A(n8064), .B(n8063), .S(n25464), .Z(n10406) );
  OAI211_X1 U2450 ( .C1(n4586), .C2(n10120), .A(n5356), .B(n9340), .ZN(n11113)
         );
  NAND3_X1 U140 ( .A1(n24795), .A2(n4832), .A3(n24212), .ZN(n10552) );
  NAND3_X1 U3244 ( .A1(n9593), .A2(n698), .A3(n9594), .ZN(n10486) );
  NOR2_X1 U449 ( .A1(n9467), .A2(n9466), .ZN(n10538) );
  OAI21_X1 U553 ( .B1(n9235), .B2(n10070), .A(n3705), .ZN(n10846) );
  AND2_X1 U1165 ( .A1(n1346), .A2(n1347), .ZN(n11196) );
  OR2_X1 U307 ( .A1(n3261), .A2(n3262), .ZN(n11171) );
  NOR2_X1 U24106 ( .A1(n2730), .A2(n8225), .ZN(n10594) );
  NAND2_X1 U1830 ( .A1(n10086), .A2(n2835), .ZN(n11214) );
  AND3_X1 U89 ( .A1(n9902), .A2(n9901), .A3(n9900), .ZN(n10969) );
  NAND2_X1 U7787 ( .A1(n7440), .A2(n7439), .ZN(n2306) );
  AOI21_X1 U314 ( .B1(n5517), .B2(n5519), .A(n4871), .ZN(n25025) );
  INV_X1 U630 ( .A(n11058), .ZN(n11054) );
  INV_X1 U3103 ( .A(n10538), .ZN(n2388) );
  BUF_X1 U516 ( .A(n9892), .Z(n10606) );
  OR2_X1 U1770 ( .A1(n10961), .A2(n10534), .ZN(n10690) );
  OAI211_X1 U776 ( .C1(n10836), .C2(n10829), .A(n10194), .B(n10193), .ZN(
        n12255) );
  OR2_X1 U884 ( .A1(n10619), .A2(n10618), .ZN(n10627) );
  OAI211_X1 U585 ( .C1(n10735), .C2(n10734), .A(n10733), .B(n10732), .ZN(
        n12137) );
  OAI211_X1 U2387 ( .C1(n10473), .C2(n10840), .A(n10472), .B(n10471), .ZN(
        n12286) );
  NAND3_X1 U2394 ( .A1(n5059), .A2(n5061), .A3(n5062), .ZN(n11659) );
  AOI21_X1 U10632 ( .B1(n11002), .B2(n11067), .A(n11001), .ZN(n12369) );
  OAI21_X1 U3847 ( .B1(n991), .B2(n10946), .A(n10945), .ZN(n12226) );
  NAND2_X1 U126 ( .A1(n4357), .A2(n10750), .ZN(n12048) );
  OR2_X1 U15348 ( .A1(n10511), .A2(n10510), .ZN(n11672) );
  OAI211_X1 U16041 ( .C1(n11529), .C2(n11528), .A(n11527), .B(n11526), .ZN(
        n12323) );
  NAND2_X1 U2476 ( .A1(n10377), .A2(n10376), .ZN(n12324) );
  AOI22_X1 U2555 ( .A1(n11035), .A2(n939), .B1(n11034), .B2(n11033), .ZN(
        n11561) );
  OAI211_X1 U352 ( .C1(n1358), .C2(n11166), .A(n11165), .B(n11164), .ZN(n12065) );
  MUX2_X1 U8576 ( .A(n9910), .B(n9911), .S(n10497), .Z(n12355) );
  NAND2_X1 U10203 ( .A1(n4051), .A2(n4048), .ZN(n12102) );
  NAND3_X1 U2371 ( .A1(n2831), .A2(n10483), .A3(n2830), .ZN(n12224) );
  AND2_X1 U1502 ( .A1(n2763), .A2(n2762), .ZN(n11607) );
  NAND2_X1 U1735 ( .A1(n9243), .A2(n9242), .ZN(n12089) );
  BUF_X1 U1006 ( .A(n12101), .Z(n11897) );
  CLKBUF_X1 U20691 ( .A(n12150), .Z(n25032) );
  NAND2_X1 U6942 ( .A1(n3312), .A2(n10390), .ZN(n12040) );
  NOR2_X1 U2365 ( .A1(n11308), .A2(n11307), .ZN(n11796) );
  AND2_X1 U9473 ( .A1(n3447), .A2(n3446), .ZN(n11295) );
  BUF_X2 U238 ( .A(n11556), .Z(n24027) );
  XNOR2_X1 U464 ( .A(n9409), .B(n9408), .ZN(n12648) );
  XNOR2_X1 U965 ( .A(n11257), .B(n11256), .ZN(n13012) );
  XOR2_X1 U1706 ( .A(n11790), .B(n11791), .Z(n24476) );
  XNOR2_X1 U2401 ( .A(n11794), .B(n24634), .ZN(n12824) );
  XNOR2_X1 U7302 ( .A(n12172), .B(n12171), .ZN(n12976) );
  INV_X1 U77 ( .A(n11287), .ZN(n13014) );
  XNOR2_X1 U16111 ( .A(n11612), .B(n11611), .ZN(n12535) );
  XNOR2_X1 U940 ( .A(n12100), .B(n12099), .ZN(n13341) );
  NOR2_X1 U4623 ( .A1(n12478), .A2(n13041), .ZN(n1646) );
  OR2_X1 U973 ( .A1(n12597), .A2(n13291), .ZN(n13289) );
  AOI22_X1 U4284 ( .A1(n24443), .A2(n13264), .B1(n5361), .B2(n13267), .ZN(
        n12832) );
  NOR2_X1 U10365 ( .A1(n304), .A2(n24930), .ZN(n13171) );
  OR2_X1 U2595 ( .A1(n399), .A2(n13341), .ZN(n13337) );
  OAI211_X1 U8050 ( .C1(n2543), .C2(n13235), .A(n2545), .B(n1374), .ZN(n13807)
         );
  OAI22_X1 U2264 ( .A1(n12441), .A2(n5112), .B1(n5113), .B2(n12737), .ZN(
        n14166) );
  OR2_X1 U359 ( .A1(n11685), .A2(n5538), .ZN(n13966) );
  MUX2_X1 U16834 ( .A(n12682), .B(n12681), .S(n13267), .Z(n13788) );
  AND3_X1 U1055 ( .A1(n12564), .A2(n12562), .A3(n12561), .ZN(n396) );
  NAND3_X1 U569 ( .A1(n12480), .A2(n12481), .A3(n12479), .ZN(n14242) );
  AOI22_X1 U5418 ( .A1(n12892), .A2(n11367), .B1(n11366), .B2(n13211), .ZN(
        n11411) );
  OR2_X1 U326 ( .A1(n4548), .A2(n4547), .ZN(n13981) );
  AND3_X1 U9030 ( .A1(n11331), .A2(n5748), .A3(n11330), .ZN(n13951) );
  AND3_X1 U1481 ( .A1(n12954), .A2(n12953), .A3(n2472), .ZN(n14205) );
  OR2_X1 U330 ( .A1(n12474), .A2(n12475), .ZN(n4116) );
  BUF_X1 U64 ( .A(n13996), .Z(n24402) );
  BUF_X1 U2269 ( .A(n13635), .Z(n13935) );
  NAND2_X1 U10615 ( .A1(n4448), .A2(n4443), .ZN(n14301) );
  OAI21_X1 U255 ( .B1(n4447), .B2(n4446), .A(n24812), .ZN(n13888) );
  NAND3_X1 U4471 ( .A1(n1828), .A2(n2715), .A3(n1393), .ZN(n14009) );
  INV_X1 U159 ( .A(n13965), .ZN(n13962) );
  NAND3_X1 U3420 ( .A1(n2888), .A2(n2889), .A3(n12880), .ZN(n14320) );
  AND2_X1 U10334 ( .A1(n12487), .A2(n12488), .ZN(n14245) );
  NOR2_X1 U17162 ( .A1(n13989), .A2(n13982), .ZN(n13985) );
  BUF_X2 U119 ( .A(n14851), .Z(n24572) );
  INV_X1 U1329 ( .A(n13744), .ZN(n13526) );
  NAND2_X1 U212 ( .A1(n11224), .A2(n2929), .ZN(n14156) );
  AND2_X1 U2222 ( .A1(n13444), .A2(n14060), .ZN(n14419) );
  AOI21_X1 U373 ( .B1(n4129), .B2(n4131), .A(n13827), .ZN(n15507) );
  NAND2_X1 U3364 ( .A1(n5708), .A2(n24827), .ZN(n15165) );
  AOI22_X1 U1052 ( .A1(n13855), .A2(n13856), .B1(n13857), .B2(n14078), .ZN(
        n14558) );
  NAND2_X1 U1533 ( .A1(n1966), .A2(n24095), .ZN(n15483) );
  NAND2_X1 U65 ( .A1(n59), .A2(n684), .ZN(n14993) );
  OAI211_X1 U2192 ( .C1(n2658), .C2(n13255), .A(n13254), .B(n2657), .ZN(n14952) );
  NOR2_X1 U235 ( .A1(n13314), .A2(n13315), .ZN(n15273) );
  NAND3_X1 U6904 ( .A1(n2503), .A2(n2507), .A3(n2502), .ZN(n15177) );
  NAND3_X1 U486 ( .A1(n13897), .A2(n13899), .A3(n13898), .ZN(n15326) );
  AND2_X1 U5467 ( .A1(n4593), .A2(n4592), .ZN(n14500) );
  AND2_X1 U2186 ( .A1(n13992), .A2(n1112), .ZN(n14788) );
  AND3_X1 U8318 ( .A1(n13369), .A2(n13368), .A3(n13367), .ZN(n15203) );
  AND2_X1 U9707 ( .A1(n3538), .A2(n3536), .ZN(n14977) );
  NAND3_X1 U3879 ( .A1(n13751), .A2(n1026), .A3(n1025), .ZN(n15464) );
  XNOR2_X1 U18277 ( .A(n14976), .B(n912), .ZN(n14978) );
  XNOR2_X1 U33 ( .A(n14422), .B(n14421), .ZN(n16427) );
  XNOR2_X1 U597 ( .A(n14771), .B(n14772), .ZN(n16016) );
  XNOR2_X1 U2164 ( .A(n14228), .B(n14229), .ZN(n16176) );
  XNOR2_X1 U18163 ( .A(n14804), .B(n14803), .ZN(n16491) );
  INV_X1 U17181 ( .A(n15019), .ZN(n15499) );
  XNOR2_X1 U374 ( .A(n15337), .B(n15336), .ZN(n15697) );
  XNOR2_X1 U2176 ( .A(n15214), .B(n15213), .ZN(n16312) );
  XNOR2_X1 U9437 ( .A(n3308), .B(n14047), .ZN(n16367) );
  XNOR2_X1 U1461 ( .A(n13738), .B(n13737), .ZN(n15646) );
  XNOR2_X1 U2127 ( .A(n4204), .B(n4205), .ZN(n2253) );
  BUF_X1 U2146 ( .A(n15707), .Z(n16442) );
  XNOR2_X1 U2173 ( .A(n15288), .B(n15289), .ZN(n16051) );
  BUF_X1 U1086 ( .A(n14350), .Z(n16177) );
  INV_X1 U283 ( .A(n15545), .ZN(n16469) );
  XNOR2_X1 U1253 ( .A(n14736), .B(n14735), .ZN(n16102) );
  XNOR2_X1 U11601 ( .A(n5494), .B(n15323), .ZN(n15695) );
  INV_X1 U1450 ( .A(n3779), .ZN(n3544) );
  XNOR2_X1 U18434 ( .A(n15206), .B(n15207), .ZN(n15557) );
  BUF_X1 U446 ( .A(n15637), .Z(n15972) );
  MUX2_X1 U2097 ( .A(n15475), .B(n15474), .S(n15950), .Z(n15872) );
  AND2_X1 U1961 ( .A1(n17436), .A2(n16429), .ZN(n17442) );
  AND4_X1 U1323 ( .A1(n15598), .A2(n15597), .A3(n15595), .A4(n15596), .ZN(
        n1139) );
  AND3_X1 U2078 ( .A1(n16446), .A2(n16444), .A3(n16445), .ZN(n1653) );
  AND2_X1 U4506 ( .A1(n5581), .A2(n15650), .ZN(n17305) );
  AND2_X1 U42 ( .A1(n16810), .A2(n16808), .ZN(n17076) );
  NAND2_X1 U46 ( .A1(n1791), .A2(n1832), .ZN(n17389) );
  AND3_X1 U8230 ( .A1(n2648), .A2(n2649), .A3(n2650), .ZN(n17336) );
  NOR2_X1 U4689 ( .A1(n15744), .A2(n16328), .ZN(n17624) );
  NAND2_X1 U378 ( .A1(n1245), .A2(n4575), .ZN(n17304) );
  AND2_X1 U10488 ( .A1(n4420), .A2(n4416), .ZN(n17114) );
  OR2_X1 U870 ( .A1(n3576), .A2(n15589), .ZN(n16731) );
  NAND2_X1 U688 ( .A1(n15601), .A2(n1673), .ZN(n16546) );
  AND2_X1 U2057 ( .A1(n15683), .A2(n15682), .ZN(n17319) );
  BUF_X2 U274 ( .A(n17062), .Z(n24585) );
  MUX2_X1 U19554 ( .A(n17122), .B(n17121), .S(n17120), .Z(n17123) );
  OR2_X1 U83 ( .A1(n16288), .A2(n2701), .ZN(n17014) );
  NAND2_X1 U769 ( .A1(n3005), .A2(n3003), .ZN(n18200) );
  NAND3_X1 U2000 ( .A1(n1133), .A2(n17070), .A3(n1070), .ZN(n18599) );
  AND3_X1 U3556 ( .A1(n24594), .A2(n16992), .A3(n16993), .ZN(n17959) );
  INV_X1 U1163 ( .A(n3706), .ZN(n24568) );
  OR2_X1 U6441 ( .A1(n1625), .A2(n1623), .ZN(n17681) );
  BUF_X1 U441 ( .A(n17933), .Z(n24536) );
  NAND2_X1 U1383 ( .A1(n24174), .A2(n16853), .ZN(n18669) );
  BUF_X1 U1083 ( .A(n18589), .Z(n24565) );
  OAI21_X1 U11658 ( .B1(n16615), .B2(n16514), .A(n5555), .ZN(n18214) );
  NAND3_X1 U429 ( .A1(n16900), .A2(n4613), .A3(n4612), .ZN(n18540) );
  XNOR2_X1 U19959 ( .A(n18098), .B(n17768), .ZN(n18573) );
  AND2_X1 U710 ( .A1(n1253), .A2(n1252), .ZN(n17819) );
  XNOR2_X1 U388 ( .A(n17930), .B(n17929), .ZN(n19499) );
  BUF_X1 U1932 ( .A(n4748), .Z(n3296) );
  XNOR2_X1 U211 ( .A(n17885), .B(n17884), .ZN(n19466) );
  XNOR2_X1 U425 ( .A(n670), .B(n18148), .ZN(n19105) );
  XNOR2_X1 U19901 ( .A(n17703), .B(n17702), .ZN(n19357) );
  CLKBUF_X1 U1958 ( .A(n18914), .Z(n17559) );
  XNOR2_X1 U1956 ( .A(n17879), .B(n17878), .ZN(n19472) );
  XNOR2_X1 U11003 ( .A(n18013), .B(n18012), .ZN(n19210) );
  BUF_X1 U1318 ( .A(n19015), .Z(n19393) );
  XNOR2_X1 U903 ( .A(n4086), .B(n1408), .ZN(n19255) );
  BUF_X1 U154 ( .A(n18690), .Z(n19412) );
  OR2_X1 U16146 ( .A1(n19412), .A2(n19413), .ZN(n18783) );
  MUX2_X1 U5855 ( .A(n18775), .B(n18774), .S(n19186), .Z(n20470) );
  AND3_X1 U1146 ( .A1(n18167), .A2(n18168), .A3(n1426), .ZN(n3480) );
  NAND4_X1 U1872 ( .A1(n19089), .A2(n3668), .A3(n19085), .A4(n19086), .ZN(
        n20268) );
  AND2_X1 U1878 ( .A1(n19137), .A2(n19136), .ZN(n20264) );
  NAND3_X1 U11719 ( .A1(n19175), .A2(n19174), .A3(n5617), .ZN(n20216) );
  OAI211_X1 U8158 ( .C1(n4580), .C2(n19167), .A(n4579), .B(n4578), .ZN(n20217)
         );
  AND3_X1 U25 ( .A1(n115), .A2(n18790), .A3(n114), .ZN(n20590) );
  OAI211_X1 U7103 ( .C1(n1990), .C2(n19406), .A(n18783), .B(n1987), .ZN(n20617) );
  NAND2_X1 U24200 ( .A1(n1000), .A2(n1003), .ZN(n20480) );
  AND2_X1 U4115 ( .A1(n19224), .A2(n5681), .ZN(n20193) );
  OAI21_X1 U201 ( .B1(n18093), .B2(n18092), .A(n18091), .ZN(n20557) );
  NOR2_X1 U20797 ( .A1(n18964), .A2(n18963), .ZN(n19991) );
  BUF_X1 U6 ( .A(n20484), .Z(n20486) );
  NAND2_X1 U1144 ( .A1(n1822), .A2(n519), .ZN(n20309) );
  NAND2_X1 U1571 ( .A1(n19350), .A2(n20390), .ZN(n20395) );
  OR2_X1 U1392 ( .A1(n17940), .A2(n17939), .ZN(n17943) );
  BUF_X2 U1388 ( .A(n17943), .Z(n20100) );
  AOI22_X1 U20958 ( .A1(n19740), .A2(n25397), .B1(n19259), .B2(n20425), .ZN(
        n19260) );
  AND3_X1 U15 ( .A1(n3430), .A2(n5541), .A3(n3429), .ZN(n1381) );
  AND3_X1 U13641 ( .A1(n3466), .A2(n3732), .A3(n19954), .ZN(n3465) );
  OAI21_X1 U1828 ( .B1(n19657), .B2(n19197), .A(n19196), .ZN(n20780) );
  OR2_X1 U17356 ( .A1(n20017), .A2(n24950), .ZN(n3041) );
  AND3_X1 U7106 ( .A1(n1992), .A2(n1993), .A3(n1991), .ZN(n21596) );
  OAI21_X1 U1827 ( .B1(n1521), .B2(n200), .A(n19118), .ZN(n20826) );
  MUX2_X1 U21385 ( .A(n19968), .B(n19967), .S(n20127), .Z(n19970) );
  NAND2_X1 U22667 ( .A1(n20876), .A2(n20873), .ZN(n21600) );
  NAND2_X1 U20821 ( .A1(n18996), .A2(n18997), .ZN(n21679) );
  NOR2_X1 U21567 ( .A1(n20295), .A2(n20294), .ZN(n21492) );
  BUF_X1 U1274 ( .A(n20585), .Z(n24353) );
  AND3_X1 U8563 ( .A1(n20119), .A2(n2874), .A3(n2873), .ZN(n21601) );
  NOR2_X1 U1806 ( .A1(n21013), .A2(n21012), .ZN(n21687) );
  AND3_X1 U11 ( .A1(n19824), .A2(n2916), .A3(n19090), .ZN(n21587) );
  XNOR2_X1 U1776 ( .A(n20342), .B(n4169), .ZN(n4273) );
  XNOR2_X1 U1407 ( .A(n19935), .B(n19934), .ZN(n22226) );
  XNOR2_X1 U568 ( .A(n19795), .B(n19796), .ZN(n22689) );
  BUF_X1 U8061 ( .A(n21872), .Z(n22426) );
  BUF_X1 U1755 ( .A(n20845), .Z(n23571) );
  BUF_X2 U947 ( .A(n24510), .Z(n24559) );
  NOR2_X1 U19358 ( .A1(n21791), .A2(n22231), .ZN(n21794) );
  NOR2_X1 U5748 ( .A1(n22176), .A2(n24396), .ZN(n21802) );
  XNOR2_X1 U1740 ( .A(n21256), .B(n21257), .ZN(n2397) );
  NOR2_X1 U1002 ( .A1(n4437), .A2(n22244), .ZN(n22184) );
  MUX2_X1 U1715 ( .A(n22183), .B(n22182), .S(n22181), .Z(n23672) );
  OR2_X1 U362 ( .A1(n996), .A2(n998), .ZN(n997) );
  OAI211_X1 U19984 ( .C1(n4362), .C2(n22200), .A(n4361), .B(n4359), .ZN(n23727) );
  MUX2_X1 U7250 ( .A(n22474), .B(n22473), .S(n22612), .Z(n23104) );
  AOI21_X1 U1724 ( .B1(n21804), .B2(n21805), .A(n21803), .ZN(n23768) );
  INV_X1 U254 ( .A(n23911), .ZN(n23926) );
  AND2_X1 U3335 ( .A1(n2296), .A2(n2297), .ZN(n23645) );
  BUF_X1 U1234 ( .A(n23129), .Z(n23143) );
  NOR2_X1 U22990 ( .A1(n23672), .A2(n23671), .ZN(n23658) );
  BUF_X2 U1707 ( .A(n21863), .Z(n23879) );
  NAND2_X1 U24347 ( .A1(n1799), .A2(n22865), .ZN(n23411) );
  NOR2_X1 U976 ( .A1(n840), .A2(n22112), .ZN(n25071) );
  NAND2_X1 U8867 ( .A1(n23650), .A2(n23612), .ZN(n1619) );
  OR2_X1 U4793 ( .A1(n5090), .A2(n24334), .ZN(n4235) );
  MUX2_X1 U23081 ( .A(n22345), .B(n22344), .S(n23166), .Z(n22347) );
  CLKBUF_X1 U1342 ( .A(Key[182]), .Z(n2058) );
  BUF_X1 U2718 ( .A(Key[175]), .Z(n1831) );
  BUF_X1 U1346 ( .A(Key[48]), .Z(n768) );
  BUF_X2 U1348 ( .A(Key[136]), .Z(n859) );
  CLKBUF_X1 U793 ( .A(Key[40]), .Z(n1920) );
  BUF_X1 U1595 ( .A(Key[105]), .Z(n1875) );
  NAND2_X1 U8283 ( .A1(n24203), .A2(n7930), .ZN(n7445) );
  BUF_X1 U6046 ( .A(n7065), .Z(n7476) );
  INV_X1 U1335 ( .A(n7662), .ZN(n269) );
  INV_X1 U8027 ( .A(n7757), .ZN(n2522) );
  NOR2_X2 U322 ( .A1(n7747), .A2(n2402), .ZN(n3588) );
  OAI21_X1 U125 ( .B1(n7998), .B2(n7997), .A(n7996), .ZN(n8779) );
  NAND3_X1 U2565 ( .A1(n2554), .A2(n2553), .A3(n2551), .ZN(n8818) );
  INV_X1 U13808 ( .A(n9886), .ZN(n9563) );
  INV_X2 U6161 ( .A(n9694), .ZN(n4993) );
  INV_X2 U1223 ( .A(n9788), .ZN(n24575) );
  INV_X2 U1221 ( .A(n9786), .ZN(n10088) );
  NAND4_X1 U2452 ( .A1(n8887), .A2(n8886), .A3(n9436), .A4(n8888), .ZN(n8934)
         );
  NAND2_X1 U168 ( .A1(n9088), .A2(n9087), .ZN(n10571) );
  XNOR2_X1 U533 ( .A(n10270), .B(n10269), .ZN(n12459) );
  NOR2_X1 U8208 ( .A1(n13266), .A2(n13264), .ZN(n12830) );
  AOI21_X1 U1482 ( .B1(n13322), .B2(n13321), .A(n13320), .ZN(n14230) );
  OAI211_X1 U1134 ( .C1(n13051), .C2(n25408), .A(n12492), .B(n12491), .ZN(
        n14244) );
  INV_X1 U1643 ( .A(n14852), .ZN(n14415) );
  CLKBUF_X1 U2227 ( .A(n12772), .Z(n14179) );
  OAI211_X1 U665 ( .C1(n13575), .C2(n13826), .A(n13896), .B(n13574), .ZN(
        n15034) );
  AND2_X1 U2189 ( .A1(n5252), .A2(n5253), .ZN(n13906) );
  OR2_X1 U23574 ( .A1(n13881), .A2(n13882), .ZN(n15393) );
  BUF_X1 U53 ( .A(n14499), .Z(n16118) );
  AND3_X1 U18820 ( .A1(n15818), .A2(n16366), .A3(n15817), .ZN(n17485) );
  MUX2_X1 U11872 ( .A(n16790), .B(n16789), .S(n17131), .Z(n18098) );
  INV_X1 U14863 ( .A(n2333), .ZN(n20388) );
  CLKBUF_X1 U1920 ( .A(n18762), .Z(n19534) );
  NAND2_X1 U3472 ( .A1(n19101), .A2(n19102), .ZN(n20517) );
  NAND2_X1 U10572 ( .A1(n3470), .A2(n24247), .ZN(n20422) );
  NAND3_X1 U1284 ( .A1(n171), .A2(n20229), .A3(n170), .ZN(n21694) );
  INV_X1 U299 ( .A(n21467), .ZN(n22969) );
  BUF_X1 U1756 ( .A(n21380), .Z(n22456) );
  NAND3_X1 U1296 ( .A1(n535), .A2(n21294), .A3(n534), .ZN(n24972) );
  NAND2_X1 U620 ( .A1(n22378), .A2(n22377), .ZN(n23937) );
  NAND2_X1 U4072 ( .A1(n3035), .A2(n21916), .ZN(n23206) );
  NOR2_X1 U1157 ( .A1(n22405), .A2(n22404), .ZN(n23293) );
  AND3_X2 U1098 ( .A1(n13511), .A2(n13510), .A3(n13509), .ZN(n14880) );
  MUX2_X2 U319 ( .A(n6962), .B(n6961), .S(n6960), .Z(n7423) );
  BUF_X2 U2494 ( .A(n9918), .Z(n9355) );
  AND2_X2 U2011 ( .A1(n6482), .A2(n839), .ZN(n512) );
  BUF_X2 U518 ( .A(n7941), .Z(n9276) );
  BUF_X2 U24 ( .A(n18730), .Z(n19479) );
  AND3_X2 U2359 ( .A1(n201), .A2(n9293), .A3(n547), .ZN(n12365) );
  OR2_X2 U672 ( .A1(n7690), .A2(n7692), .ZN(n8315) );
  AOI21_X2 U204 ( .B1(n10132), .B2(n10133), .A(n10131), .ZN(n10559) );
  NAND2_X2 U8827 ( .A1(n6205), .A2(n5450), .ZN(n8014) );
  AND3_X2 U10047 ( .A1(n3874), .A2(n3875), .A3(n3873), .ZN(n13417) );
  NAND3_X2 U684 ( .A1(n7394), .A2(n2893), .A3(n7393), .ZN(n8375) );
  OR2_X2 U360 ( .A1(n6433), .A2(n6432), .ZN(n8316) );
  XNOR2_X2 U1266 ( .A(n7780), .B(n7779), .ZN(n9934) );
  AND3_X2 U828 ( .A1(n9413), .A2(n9412), .A3(n2778), .ZN(n11084) );
  OAI21_X2 U1175 ( .B1(n17021), .B2(n17022), .A(n17020), .ZN(n18325) );
  NAND2_X2 U266 ( .A1(n9258), .A2(n10047), .ZN(n10740) );
  OR2_X2 U13297 ( .A1(n7301), .A2(n7300), .ZN(n8147) );
  BUF_X2 U2141 ( .A(n15549), .Z(n16063) );
  NOR2_X2 U2242 ( .A1(n300), .A2(n14063), .ZN(n3533) );
  NAND3_X2 U6701 ( .A1(n24276), .A2(n24277), .A3(n6029), .ZN(n7602) );
  NAND2_X2 U865 ( .A1(n3431), .A2(n3433), .ZN(n18350) );
  OR2_X2 U2655 ( .A1(n6249), .A2(n6248), .ZN(n7734) );
  OR2_X2 U2590 ( .A1(n24578), .A2(n7735), .ZN(n7645) );
  AND2_X2 U3031 ( .A1(n9762), .A2(n9620), .ZN(n9760) );
  OR2_X2 U1077 ( .A1(n16407), .A2(n802), .ZN(n16962) );
  AND3_X2 U1049 ( .A1(n5695), .A2(n2061), .A3(n6181), .ZN(n7762) );
  BUF_X2 U2028 ( .A(n15774), .Z(n16302) );
  AND2_X2 U1995 ( .A1(n3392), .A2(n3390), .ZN(n17970) );
  BUF_X2 U607 ( .A(n6236), .Z(n24051) );
  NAND2_X2 U1979 ( .A1(n16977), .A2(n4246), .ZN(n18562) );
  OR2_X2 U20750 ( .A1(n25039), .A2(n17335), .ZN(n3818) );
  OR2_X2 U12974 ( .A1(n6761), .A2(n6760), .ZN(n8427) );
  XNOR2_X2 U23694 ( .A(n11400), .B(n11399), .ZN(n12785) );
  OAI211_X2 U1222 ( .C1(n1510), .C2(n1512), .A(n1511), .B(n16350), .ZN(n17734)
         );
  XNOR2_X2 U1109 ( .A(n8260), .B(n8259), .ZN(n10176) );
  BUF_X1 U603 ( .A(n6236), .Z(n24050) );
  NAND4_X2 U720 ( .A1(n5986), .A2(n2593), .A3(n5987), .A4(n5988), .ZN(n7323)
         );
  NAND3_X2 U4455 ( .A1(n16238), .A2(n16237), .A3(n16239), .ZN(n17208) );
  BUF_X2 U1127 ( .A(n11217), .Z(n233) );
  OR2_X2 U2277 ( .A1(n3631), .A2(n3632), .ZN(n14089) );
  OR2_X2 U117 ( .A1(n5820), .A2(n5821), .ZN(n7585) );
  AND4_X2 U1025 ( .A1(n3079), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n11268)
         );
  AND2_X2 U414 ( .A1(n6056), .A2(n6055), .ZN(n8021) );
  MUX2_X2 U8534 ( .A(n18595), .B(n18594), .S(n19419), .Z(n20618) );
  NOR2_X2 U23264 ( .A1(n23050), .A2(n23040), .ZN(n23055) );
  XNOR2_X2 U572 ( .A(Key[128]), .B(Plaintext[128]), .ZN(n6072) );
  AND2_X2 U217 ( .A1(n7249), .A2(n7248), .ZN(n8460) );
  OAI211_X2 U19699 ( .C1(n5406), .C2(n17429), .A(n17428), .B(n17427), .ZN(
        n18515) );
  OR2_X2 U2463 ( .A1(n9843), .A2(n24085), .ZN(n9340) );
  NAND2_X2 U386 ( .A1(n19143), .A2(n19144), .ZN(n20411) );
  AND3_X2 U2443 ( .A1(n9396), .A2(n9395), .A3(n9394), .ZN(n10730) );
  XNOR2_X2 U1218 ( .A(Key[0]), .B(Plaintext[0]), .ZN(n6455) );
  NAND2_X2 U242 ( .A1(n40), .A2(n1232), .ZN(n17413) );
  NAND3_X2 U8893 ( .A1(n24740), .A2(n10101), .A3(n4258), .ZN(n11216) );
  NOR2_X2 U1045 ( .A1(n14515), .A2(n14514), .ZN(n15063) );
  NOR2_X2 U532 ( .A1(n1286), .A2(n1285), .ZN(n16859) );
  OR2_X2 U10626 ( .A1(n7624), .A2(n7623), .ZN(n8458) );
  BUF_X2 U707 ( .A(n6267), .Z(n6164) );
  BUF_X2 U843 ( .A(n16405), .Z(n24061) );
  BUF_X2 U1303 ( .A(n9255), .Z(n260) );
  BUF_X2 U2291 ( .A(n12576), .Z(n13336) );
  NOR2_X2 U1513 ( .A1(n10209), .A2(n10208), .ZN(n10884) );
  XNOR2_X2 U12150 ( .A(Key[60]), .B(Plaintext[60]), .ZN(n6964) );
  NAND2_X2 U648 ( .A1(n3628), .A2(n3629), .ZN(n17312) );
  AND2_X2 U2558 ( .A1(n24629), .A2(n9940), .ZN(n10800) );
  NOR2_X2 U11897 ( .A1(n13047), .A2(n13046), .ZN(n13824) );
  NAND2_X2 U2736 ( .A1(n25185), .A2(n4697), .ZN(n7573) );
  NAND2_X2 U2348 ( .A1(n5816), .A2(n3365), .ZN(n8596) );
  MUX2_X2 U264 ( .A(n16387), .B(n16386), .S(n15655), .Z(n16963) );
  BUF_X2 U1411 ( .A(n18812), .Z(n19384) );
  MUX2_X2 U15557 ( .A(n10909), .B(n10908), .S(n10907), .Z(n12183) );
  OR2_X2 U428 ( .A1(n7927), .A2(n7928), .ZN(n5607) );
  XNOR2_X2 U934 ( .A(n5844), .B(Key[160]), .ZN(n6912) );
  OR2_X2 U948 ( .A1(n7050), .A2(n7051), .ZN(n8457) );
  AND3_X2 U39 ( .A1(n16263), .A2(n16265), .A3(n16264), .ZN(n17824) );
  OAI21_X2 U3105 ( .B1(n14256), .B2(n13927), .A(n13382), .ZN(n14694) );
  CLKBUF_X3 U315 ( .A(n14304), .Z(n24588) );
  INV_X2 U11400 ( .A(n6375), .ZN(n6906) );
  OR2_X2 U5430 ( .A1(n13984), .A2(n13922), .ZN(n1899) );
  BUF_X2 U2781 ( .A(n6534), .Z(n24592) );
  BUF_X1 U461 ( .A(n9481), .Z(n10008) );
  INV_X1 U1514 ( .A(n10079), .ZN(n9507) );
  NAND3_X1 U9716 ( .A1(n9607), .A2(n9605), .A3(n9606), .ZN(n10613) );
  OR2_X1 U1788 ( .A1(n9826), .A2(n9825), .ZN(n10952) );
  BUF_X2 U219 ( .A(n10534), .Z(n11151) );
  AND3_X1 U279 ( .A1(n31), .A2(n1893), .A3(n1894), .ZN(n13569) );
  NAND3_X1 U964 ( .A1(n13630), .A2(n13631), .A3(n176), .ZN(n15436) );
  XNOR2_X1 U18259 ( .A(n14942), .B(n14941), .ZN(n16447) );
  AND2_X1 U8921 ( .A1(n24741), .A2(n15623), .ZN(n16932) );
  AOI21_X2 U11851 ( .B1(n16013), .B2(n16012), .A(n16011), .ZN(n16021) );
  NAND2_X1 U1888 ( .A1(n1120), .A2(n1121), .ZN(n20055) );
  AND3_X1 U1861 ( .A1(n18780), .A2(n18781), .A3(n18779), .ZN(n20060) );
  BUF_X2 U9 ( .A(n14435), .Z(n24556) );
  MUX2_X1 U21 ( .A(n10402), .B(n10401), .S(n25250), .Z(n11640) );
  BUF_X2 U23 ( .A(n10147), .Z(n25206) );
  INV_X2 U29 ( .A(n1629), .ZN(n25242) );
  XNOR2_X2 U31 ( .A(n18430), .B(n18429), .ZN(n18505) );
  OR2_X2 U38 ( .A1(n19661), .A2(n19850), .ZN(n24288) );
  NAND2_X2 U44 ( .A1(n25290), .A2(n18988), .ZN(n20136) );
  BUF_X2 U47 ( .A(n20249), .Z(n24077) );
  AND2_X2 U68 ( .A1(n1556), .A2(n209), .ZN(n20345) );
  BUF_X2 U71 ( .A(n10245), .Z(n10648) );
  OR2_X2 U72 ( .A1(n1983), .A2(n16219), .ZN(n15925) );
  OAI21_X2 U75 ( .B1(n8320), .B2(n2404), .A(n1463), .ZN(n8551) );
  BUF_X2 U79 ( .A(n22809), .Z(n25241) );
  OAI211_X1 U84 ( .C1(n20184), .C2(n20186), .A(n19663), .B(n2339), .ZN(n21311)
         );
  NAND3_X1 U87 ( .A1(n20490), .A2(n24274), .A3(n20489), .ZN(n21027) );
  AOI211_X1 U92 ( .C1(n21289), .C2(n22686), .A(n5770), .B(n21817), .ZN(n21291)
         );
  INV_X1 U113 ( .A(n13643), .ZN(n24589) );
  NAND2_X1 U128 ( .A1(n16308), .A2(n16307), .ZN(n17012) );
  BUF_X1 U131 ( .A(n15905), .Z(n15904) );
  INV_X1 U132 ( .A(n15905), .ZN(n17180) );
  AOI22_X1 U136 ( .A1(n3127), .A2(n20562), .B1(n20093), .B2(n25221), .ZN(
        n19876) );
  OAI211_X1 U150 ( .C1(n13614), .C2(n25247), .A(n12823), .B(n12822), .ZN(
        n14900) );
  NOR2_X1 U153 ( .A1(n13788), .A2(n13785), .ZN(n14140) );
  BUF_X2 U161 ( .A(n9931), .Z(n25217) );
  OAI211_X2 U173 ( .C1(n3119), .C2(n10222), .A(n10766), .B(n10221), .ZN(n12313) );
  BUF_X1 U177 ( .A(n13012), .Z(n25198) );
  OAI21_X2 U203 ( .B1(n300), .B2(n12592), .A(n25549), .ZN(n15168) );
  AOI21_X2 U206 ( .B1(n14103), .B2(n4877), .A(n4876), .ZN(n25394) );
  NOR2_X2 U225 ( .A1(n15832), .A2(n151), .ZN(n25472) );
  AND3_X2 U231 ( .A1(n24788), .A2(n24787), .A3(n24786), .ZN(n16572) );
  AND3_X2 U236 ( .A1(n638), .A2(n16632), .A3(n16631), .ZN(n25390) );
  OAI211_X2 U237 ( .C1(n17169), .C2(n2430), .A(n17168), .B(n514), .ZN(n25380)
         );
  XNOR2_X2 U251 ( .A(n20642), .B(n20213), .ZN(n21839) );
  NAND4_X2 U256 ( .A1(n15727), .A2(n15730), .A3(n15728), .A4(n15729), .ZN(
        n17296) );
  OAI21_X2 U258 ( .B1(n22732), .B2(n22731), .A(n22730), .ZN(n23478) );
  BUF_X2 U262 ( .A(n18396), .Z(n25194) );
  NAND4_X1 U271 ( .A1(n16880), .A2(n16881), .A3(n16882), .A4(n16879), .ZN(
        n18396) );
  OAI211_X2 U276 ( .C1(n1409), .C2(n16712), .A(n27), .B(n26), .ZN(n18633) );
  OAI21_X2 U277 ( .B1(n2349), .B2(n2352), .A(n2348), .ZN(n5971) );
  AND4_X2 U278 ( .A1(n5424), .A2(n5425), .A3(n24533), .A4(n5423), .ZN(n21414)
         );
  XNOR2_X2 U297 ( .A(Key[71]), .B(Plaintext[71]), .ZN(n6578) );
  NAND4_X2 U305 ( .A1(n3991), .A2(n3992), .A3(n15684), .A4(n15685), .ZN(n18080) );
  AOI21_X2 U308 ( .B1(n1268), .B2(n12662), .A(n1267), .ZN(n13488) );
  BUF_X2 U309 ( .A(n16405), .Z(n24062) );
  NAND3_X2 U311 ( .A1(n2758), .A2(n2759), .A3(n5901), .ZN(n8412) );
  MUX2_X2 U324 ( .A(n22170), .B(n22071), .S(n21712), .Z(n22075) );
  NAND3_X2 U327 ( .A1(n6043), .A2(n6042), .A3(n6041), .ZN(n7597) );
  OR2_X2 U342 ( .A1(n7632), .A2(n7631), .ZN(n8706) );
  XNOR2_X2 U350 ( .A(Plaintext[64]), .B(Key[64]), .ZN(n6575) );
  MUX2_X2 U358 ( .A(n6349), .B(n6348), .S(n6347), .Z(n7809) );
  XNOR2_X2 U365 ( .A(Key[79]), .B(Plaintext[79]), .ZN(n6732) );
  XNOR2_X2 U366 ( .A(n8254), .B(n8253), .ZN(n10186) );
  XNOR2_X2 U371 ( .A(n21566), .B(n21565), .ZN(n22958) );
  OAI21_X2 U389 ( .B1(n6672), .B2(n6671), .A(n6670), .ZN(n7991) );
  NAND2_X2 U390 ( .A1(n2858), .A2(n3056), .ZN(n8754) );
  OR2_X2 U394 ( .A1(n28), .A2(n6786), .ZN(n7977) );
  XNOR2_X2 U395 ( .A(n5862), .B(Key[28]), .ZN(n6532) );
  BUF_X2 U397 ( .A(n13305), .Z(n13307) );
  XNOR2_X2 U406 ( .A(n11697), .B(n11696), .ZN(n13305) );
  BUF_X2 U408 ( .A(n19762), .Z(n25195) );
  XNOR2_X1 U424 ( .A(n18391), .B(n18392), .ZN(n19762) );
  CLKBUF_X1 U434 ( .A(n14338), .Z(n25196) );
  BUF_X2 U435 ( .A(n14338), .Z(n25197) );
  NOR2_X1 U440 ( .A1(n13503), .A2(n13504), .ZN(n14338) );
  XNOR2_X2 U448 ( .A(n5870), .B(Key[46]), .ZN(n6956) );
  XNOR2_X2 U456 ( .A(n9006), .B(n9005), .ZN(n10026) );
  AOI22_X2 U460 ( .A1(n11454), .A2(n24973), .B1(n14289), .B2(n11453), .ZN(
        n14685) );
  NAND2_X2 U463 ( .A1(n24807), .A2(n818), .ZN(n20134) );
  OR2_X2 U465 ( .A1(n9561), .A2(n25307), .ZN(n10907) );
  BUF_X1 U473 ( .A(n13012), .Z(n25199) );
  XNOR2_X2 U504 ( .A(n17708), .B(n18493), .ZN(n19452) );
  BUF_X2 U513 ( .A(n6414), .Z(n6695) );
  BUF_X2 U514 ( .A(n11350), .Z(n13206) );
  XNOR2_X2 U519 ( .A(n13914), .B(n13913), .ZN(n16397) );
  XNOR2_X2 U525 ( .A(n5872), .B(Key[55]), .ZN(n6690) );
  NAND2_X2 U526 ( .A1(n6614), .A2(n6613), .ZN(n7781) );
  XNOR2_X2 U537 ( .A(n2408), .B(n2407), .ZN(n223) );
  MUX2_X2 U547 ( .A(n19096), .B(n19095), .S(n19380), .Z(n20515) );
  OAI21_X2 U552 ( .B1(n4741), .B2(n13227), .A(n3351), .ZN(n13918) );
  OAI211_X2 U563 ( .C1(n14298), .C2(n14297), .A(n14295), .B(n24146), .ZN(
        n14634) );
  BUF_X1 U565 ( .A(n17215), .Z(n25200) );
  BUF_X2 U571 ( .A(n17215), .Z(n25201) );
  AOI22_X1 U578 ( .A1(n16227), .A2(n16226), .B1(n16228), .B2(n16304), .ZN(
        n17215) );
  CLKBUF_X3 U579 ( .A(n21700), .Z(n25202) );
  NOR2_X1 U582 ( .A1(n17494), .A2(n20665), .ZN(n21700) );
  BUF_X2 U609 ( .A(n11063), .Z(n25203) );
  AND2_X2 U611 ( .A1(n25467), .A2(n25468), .ZN(n18611) );
  OAI211_X2 U624 ( .C1(n7915), .C2(n8076), .A(n7160), .B(n7159), .ZN(n9082) );
  OAI211_X2 U628 ( .C1(n22316), .C2(n22612), .A(n22315), .B(n22314), .ZN(
        n23164) );
  AND2_X2 U635 ( .A1(n2448), .A2(n6540), .ZN(n7384) );
  NOR2_X2 U637 ( .A1(n12949), .A2(n12950), .ZN(n14208) );
  NAND2_X2 U639 ( .A1(n10629), .A2(n25306), .ZN(n11735) );
  AND3_X2 U650 ( .A1(n1435), .A2(n1378), .A3(n4609), .ZN(n1370) );
  NAND4_X2 U655 ( .A1(n7253), .A2(n7254), .A3(n7251), .A4(n7252), .ZN(n8542)
         );
  OAI22_X2 U661 ( .A1(n4807), .A2(n3736), .B1(n4806), .B2(n3735), .ZN(n17275)
         );
  AND2_X2 U667 ( .A1(n683), .A2(n682), .ZN(n4807) );
  AOI22_X1 U669 ( .A1(n9385), .A2(n10185), .B1(n8262), .B2(n8261), .ZN(n10505)
         );
  OR2_X2 U697 ( .A1(n5491), .A2(n3834), .ZN(n21981) );
  AND2_X2 U715 ( .A1(n1665), .A2(n25318), .ZN(n21573) );
  OAI211_X1 U722 ( .C1(n23200), .C2(n23199), .A(n24609), .B(n24612), .ZN(
        n23211) );
  AND2_X2 U728 ( .A1(n473), .A2(n474), .ZN(n18275) );
  NAND2_X2 U731 ( .A1(n13961), .A2(n13960), .ZN(n15109) );
  XNOR2_X2 U732 ( .A(Key[8]), .B(Plaintext[8]), .ZN(n6034) );
  AND2_X2 U734 ( .A1(n3757), .A2(n24295), .ZN(n11401) );
  NOR2_X2 U736 ( .A1(n953), .A2(n954), .ZN(n10886) );
  NOR2_X2 U739 ( .A1(n13616), .A2(n13615), .ZN(n14755) );
  CLKBUF_X1 U740 ( .A(n20233), .Z(n25204) );
  BUF_X2 U752 ( .A(n20233), .Z(n25205) );
  OAI211_X1 U753 ( .C1(n19483), .C2(n19482), .A(n24605), .B(n24716), .ZN(
        n20233) );
  BUF_X1 U754 ( .A(n10147), .Z(n25207) );
  XNOR2_X1 U761 ( .A(n25137), .B(n25136), .ZN(n10147) );
  AND2_X2 U764 ( .A1(n4673), .A2(n4674), .ZN(n4672) );
  AND2_X2 U771 ( .A1(n1318), .A2(n1317), .ZN(n10870) );
  NAND2_X2 U795 ( .A1(n22920), .A2(n23018), .ZN(n23531) );
  MUX2_X2 U803 ( .A(n22913), .B(n22912), .S(n23461), .Z(n22920) );
  NAND2_X2 U809 ( .A1(n10981), .A2(n10980), .ZN(n12410) );
  AND3_X4 U812 ( .A1(n5259), .A2(n5258), .A3(n5260), .ZN(n23112) );
  XNOR2_X2 U819 ( .A(n11963), .B(n11964), .ZN(n12834) );
  OR2_X2 U821 ( .A1(n16701), .A2(n16700), .ZN(n20335) );
  AND2_X2 U822 ( .A1(n1532), .A2(n5273), .ZN(n10793) );
  CLKBUF_X1 U827 ( .A(n14242), .Z(n25208) );
  BUF_X1 U835 ( .A(n14242), .Z(n25209) );
  AOI22_X2 U836 ( .A1(n15578), .A2(n15577), .B1(n15576), .B2(n15575), .ZN(
        n18240) );
  BUF_X2 U842 ( .A(n6062), .Z(n6733) );
  OR2_X2 U844 ( .A1(n18654), .A2(n18655), .ZN(n20616) );
  XNOR2_X2 U845 ( .A(n16664), .B(n16665), .ZN(n19555) );
  XNOR2_X2 U847 ( .A(n5851), .B(Key[154]), .ZN(n6767) );
  OAI211_X2 U857 ( .C1(n7344), .C2(n7256), .A(n7260), .B(n7259), .ZN(n8345) );
  XNOR2_X2 U858 ( .A(Key[176]), .B(Plaintext[176]), .ZN(n5966) );
  XNOR2_X2 U859 ( .A(n5874), .B(Key[58]), .ZN(n6976) );
  NAND2_X2 U860 ( .A1(n3173), .A2(n6646), .ZN(n7364) );
  BUF_X2 U866 ( .A(n12795), .Z(n25085) );
  OAI211_X2 U871 ( .C1(n2413), .C2(n9848), .A(n9847), .B(n9846), .ZN(n10698)
         );
  AOI21_X2 U873 ( .B1(n17269), .B2(n17270), .A(n17268), .ZN(n18285) );
  NAND3_X2 U878 ( .A1(n13608), .A2(n1061), .A3(n1060), .ZN(n15487) );
  XNOR2_X2 U885 ( .A(Key[159]), .B(Plaintext[159]), .ZN(n6915) );
  AND2_X1 U894 ( .A1(n13108), .A2(n12856), .ZN(n13661) );
  XNOR2_X2 U895 ( .A(n12229), .B(n12228), .ZN(n13108) );
  AND3_X2 U897 ( .A1(n5353), .A2(n5352), .A3(n5354), .ZN(n11116) );
  BUF_X1 U904 ( .A(n19105), .Z(n24344) );
  XNOR2_X2 U914 ( .A(n3670), .B(n3669), .ZN(n16268) );
  NAND2_X2 U915 ( .A1(n16860), .A2(n24229), .ZN(n18308) );
  MUX2_X2 U917 ( .A(n10578), .B(n10577), .S(n11175), .Z(n11638) );
  AND3_X2 U918 ( .A1(n3244), .A2(n5108), .A3(n3243), .ZN(n11637) );
  OAI211_X2 U919 ( .C1(n15669), .C2(n16334), .A(n2286), .B(n1444), .ZN(n16927)
         );
  XNOR2_X2 U925 ( .A(n15511), .B(n15510), .ZN(n16437) );
  OAI211_X2 U927 ( .C1(n5630), .C2(n5628), .A(n5629), .B(n5627), .ZN(n11619)
         );
  OAI211_X2 U928 ( .C1(n6754), .C2(n5808), .A(n5807), .B(n5806), .ZN(n7579) );
  XNOR2_X2 U931 ( .A(n21095), .B(n21094), .ZN(n23998) );
  XNOR2_X2 U937 ( .A(n11497), .B(n11496), .ZN(n13067) );
  OR2_X2 U938 ( .A1(n962), .A2(n958), .ZN(n3428) );
  NAND3_X2 U939 ( .A1(n3054), .A2(n17133), .A3(n3053), .ZN(n18341) );
  NAND2_X2 U946 ( .A1(n10998), .A2(n10999), .ZN(n11907) );
  NAND2_X2 U951 ( .A1(n3918), .A2(n109), .ZN(n20597) );
  XNOR2_X2 U960 ( .A(n15030), .B(n15031), .ZN(n16342) );
  XNOR2_X2 U961 ( .A(n5782), .B(Key[94]), .ZN(n6233) );
  XNOR2_X2 U969 ( .A(n6004), .B(Key[101]), .ZN(n625) );
  NAND2_X2 U970 ( .A1(n15652), .A2(n726), .ZN(n17316) );
  XNOR2_X2 U971 ( .A(n5159), .B(n5160), .ZN(n19446) );
  NAND3_X2 U975 ( .A1(n25134), .A2(n25135), .A3(n10366), .ZN(n11960) );
  BUF_X1 U1008 ( .A(n16176), .Z(n25210) );
  MUX2_X2 U1012 ( .A(n9381), .B(n10255), .S(n10128), .Z(n10729) );
  BUF_X1 U1014 ( .A(n20182), .Z(n25211) );
  BUF_X1 U1020 ( .A(n20182), .Z(n25212) );
  OAI21_X1 U1021 ( .B1(n358), .B2(n18723), .A(n18722), .ZN(n20182) );
  XNOR2_X2 U1026 ( .A(n12418), .B(n12417), .ZN(n13345) );
  OR2_X2 U1030 ( .A1(n15722), .A2(n15721), .ZN(n16708) );
  CLKBUF_X1 U1033 ( .A(n17361), .Z(n25213) );
  BUF_X1 U1051 ( .A(n17361), .Z(n25214) );
  BUF_X1 U1057 ( .A(n17361), .Z(n25215) );
  OAI211_X1 U1058 ( .C1(n3544), .C2(n16402), .A(n15913), .B(n24792), .ZN(
        n17361) );
  NAND2_X2 U1067 ( .A1(n12693), .A2(n5021), .ZN(n14141) );
  NOR2_X2 U1068 ( .A1(n17500), .A2(n17499), .ZN(n18994) );
  AOI21_X2 U1070 ( .B1(n13866), .B2(n13865), .A(n2225), .ZN(n14724) );
  XNOR2_X2 U1073 ( .A(n5790), .B(Key[86]), .ZN(n5796) );
  XNOR2_X2 U1078 ( .A(n11720), .B(n11721), .ZN(n12555) );
  AOI22_X1 U1080 ( .A1(n9579), .A2(n9578), .B1(n9577), .B2(n10904), .ZN(n12150) );
  XNOR2_X2 U1081 ( .A(n11430), .B(n12013), .ZN(n13057) );
  OAI21_X2 U1084 ( .B1(n18882), .B2(n24344), .A(n1547), .ZN(n20522) );
  OAI21_X2 U1101 ( .B1(n1282), .B2(n1281), .A(n1280), .ZN(n8613) );
  XNOR2_X2 U1113 ( .A(n21637), .B(n21636), .ZN(n22938) );
  BUF_X2 U1138 ( .A(n16388), .Z(n15977) );
  XNOR2_X2 U1139 ( .A(n5839), .B(Key[138]), .ZN(n6078) );
  CLKBUF_X1 U1143 ( .A(n9931), .Z(n25216) );
  XNOR2_X1 U1148 ( .A(n7614), .B(n7613), .ZN(n9931) );
  CLKBUF_X1 U1150 ( .A(n17167), .Z(n25218) );
  BUF_X2 U1158 ( .A(n17167), .Z(n25219) );
  AOI22_X1 U1160 ( .A1(n16059), .A2(n16473), .B1(n16058), .B2(n16474), .ZN(
        n17167) );
  XNOR2_X2 U1162 ( .A(n7310), .B(n7311), .ZN(n9211) );
  NAND2_X2 U1172 ( .A1(n2841), .A2(n6399), .ZN(n7563) );
  CLKBUF_X1 U1178 ( .A(n20095), .Z(n25220) );
  CLKBUF_X3 U1179 ( .A(n20095), .Z(n25221) );
  NOR2_X1 U1180 ( .A1(n19730), .A2(n18395), .ZN(n20095) );
  XNOR2_X2 U1183 ( .A(n11625), .B(n11624), .ZN(n12534) );
  XNOR2_X2 U1184 ( .A(Key[157]), .B(Plaintext[157]), .ZN(n6918) );
  XNOR2_X2 U1186 ( .A(n5990), .B(Key[105]), .ZN(n6823) );
  XNOR2_X2 U1192 ( .A(n2113), .B(n14316), .ZN(n16381) );
  BUF_X2 U1193 ( .A(n21493), .Z(n25222) );
  OAI22_X1 U1195 ( .A1(n18859), .A2(n19850), .B1(n20071), .B2(n18858), .ZN(
        n21493) );
  XNOR2_X2 U1206 ( .A(n10745), .B(n10744), .ZN(n13150) );
  XNOR2_X2 U1207 ( .A(n20123), .B(n20122), .ZN(n22361) );
  XNOR2_X2 U1219 ( .A(n12374), .B(n12373), .ZN(n12636) );
  NAND3_X2 U1220 ( .A1(n24215), .A2(n11103), .A3(n11104), .ZN(n12212) );
  NAND2_X2 U1238 ( .A1(n3088), .A2(n4561), .ZN(n10772) );
  XNOR2_X2 U1245 ( .A(n11383), .B(n11382), .ZN(n13027) );
  NOR2_X2 U1246 ( .A1(n2385), .A2(n10454), .ZN(n12209) );
  AOI21_X2 U1254 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n10970) );
  OR2_X2 U1255 ( .A1(n14024), .A2(n14023), .ZN(n15097) );
  AND4_X2 U1260 ( .A1(n10697), .A2(n10695), .A3(n10696), .A4(n3209), .ZN(
        n11661) );
  XNOR2_X2 U1269 ( .A(n8097), .B(n8096), .ZN(n9027) );
  OAI21_X2 U1278 ( .B1(n17245), .B2(n17246), .A(n17244), .ZN(n18621) );
  AND2_X2 U1283 ( .A1(n14441), .A2(n1446), .ZN(n15223) );
  XNOR2_X2 U1287 ( .A(Key[107]), .B(Plaintext[107]), .ZN(n5992) );
  INV_X1 U1292 ( .A(n13578), .ZN(n14182) );
  NOR2_X2 U1300 ( .A1(n13542), .A2(n13541), .ZN(n15178) );
  XNOR2_X2 U1301 ( .A(n21405), .B(n21404), .ZN(n22932) );
  BUF_X1 U1307 ( .A(n20217), .Z(n25223) );
  CLKBUF_X1 U1308 ( .A(n20217), .Z(n25224) );
  XNOR2_X2 U1313 ( .A(Key[109]), .B(Plaintext[109]), .ZN(n6244) );
  BUF_X1 U1320 ( .A(n17108), .Z(n25225) );
  BUF_X1 U1321 ( .A(n17108), .Z(n25226) );
  CLKBUF_X1 U1324 ( .A(n17108), .Z(n25227) );
  AOI21_X1 U1326 ( .B1(n4338), .B2(n15805), .A(n4337), .ZN(n17108) );
  OAI211_X2 U1331 ( .C1(n14198), .C2(n14148), .A(n14147), .B(n3678), .ZN(
        n15526) );
  OAI211_X2 U1339 ( .C1(n13484), .C2(n12678), .A(n12677), .B(n12676), .ZN(
        n14845) );
  OAI21_X2 U1358 ( .B1(n5934), .B2(n5935), .A(n5933), .ZN(n7464) );
  BUF_X2 U1372 ( .A(n9045), .Z(n25228) );
  BUF_X1 U1373 ( .A(n10736), .Z(n25229) );
  BUF_X2 U1380 ( .A(n10736), .Z(n25230) );
  XNOR2_X2 U1382 ( .A(n16738), .B(n24719), .ZN(n19264) );
  CLKBUF_X1 U1396 ( .A(n10953), .Z(n25231) );
  BUF_X1 U1416 ( .A(n10953), .Z(n25232) );
  CLKBUF_X1 U1427 ( .A(n10953), .Z(n25233) );
  XNOR2_X2 U1438 ( .A(n11859), .B(n11860), .ZN(n12928) );
  XNOR2_X2 U1444 ( .A(n5961), .B(Key[163]), .ZN(n6480) );
  XNOR2_X2 U1460 ( .A(n11871), .B(n11872), .ZN(n12897) );
  OAI21_X2 U1470 ( .B1(n12832), .B2(n5644), .A(n5643), .ZN(n4844) );
  OAI21_X2 U1479 ( .B1(n6994), .B2(n6995), .A(n6993), .ZN(n7961) );
  XNOR2_X2 U1484 ( .A(n7206), .B(n7207), .ZN(n9388) );
  OAI21_X2 U1498 ( .B1(n20363), .B2(n20362), .A(n20361), .ZN(n21996) );
  XNOR2_X2 U1508 ( .A(n25140), .B(n18503), .ZN(n19460) );
  OAI21_X2 U1515 ( .B1(n4898), .B2(n4896), .A(n16511), .ZN(n16616) );
  AND2_X2 U1527 ( .A1(n4900), .A2(n617), .ZN(n16511) );
  XNOR2_X2 U1541 ( .A(n14872), .B(n14871), .ZN(n16220) );
  XNOR2_X2 U1544 ( .A(n111), .B(n11980), .ZN(n13265) );
  NOR2_X2 U1546 ( .A1(n16874), .A2(n16875), .ZN(n17969) );
  XNOR2_X2 U1553 ( .A(n11405), .B(n11404), .ZN(n13028) );
  XNOR2_X2 U1564 ( .A(n15382), .B(n15381), .ZN(n16067) );
  OAI211_X2 U1612 ( .C1(n12749), .C2(n14058), .A(n12748), .B(n12747), .ZN(
        n15184) );
  NOR2_X2 U1621 ( .A1(n22943), .A2(n22942), .ZN(n24492) );
  OAI21_X2 U1638 ( .B1(n15671), .B2(n5706), .A(n13375), .ZN(n17414) );
  BUF_X2 U1657 ( .A(n12369), .Z(n25234) );
  XNOR2_X2 U1688 ( .A(n12078), .B(n12079), .ZN(n231) );
  XNOR2_X2 U1697 ( .A(n6002), .B(Key[118]), .ZN(n6848) );
  XNOR2_X2 U1698 ( .A(n5303), .B(n5301), .ZN(n19313) );
  OAI21_X2 U1717 ( .B1(n9392), .B2(n1093), .A(n1092), .ZN(n10583) );
  BUF_X2 U1718 ( .A(n8945), .Z(n25235) );
  OAI21_X2 U1722 ( .B1(n3729), .B2(n3730), .A(n551), .ZN(n10369) );
  XNOR2_X2 U1739 ( .A(n1576), .B(Key[59]), .ZN(n1147) );
  BUF_X2 U1775 ( .A(n12137), .Z(n25236) );
  AND3_X2 U1783 ( .A1(n1216), .A2(n1215), .A3(n1220), .ZN(n11440) );
  AOI21_X2 U1804 ( .B1(n7245), .B2(n7186), .A(n1736), .ZN(n9107) );
  XNOR2_X2 U1808 ( .A(n8885), .B(n8884), .ZN(n9433) );
  NAND2_X2 U1809 ( .A1(n20189), .A2(n1487), .ZN(n22007) );
  CLKBUF_X1 U1813 ( .A(n15697), .Z(n25237) );
  BUF_X2 U1818 ( .A(n15697), .Z(n25238) );
  CLKBUF_X1 U1822 ( .A(n23251), .Z(n24377) );
  NAND2_X1 U1848 ( .A1(n21758), .A2(n2690), .ZN(n23595) );
  BUF_X1 U1855 ( .A(n23470), .Z(n23481) );
  OAI211_X1 U1874 ( .C1(n21913), .C2(n22273), .A(n21912), .B(n21911), .ZN(
        n22575) );
  NOR2_X1 U1881 ( .A1(n22204), .A2(n22203), .ZN(n23740) );
  INV_X1 U1882 ( .A(n20561), .ZN(n20562) );
  AOI22_X1 U1889 ( .A1(n16834), .A2(n3981), .B1(n3982), .B2(n16833), .ZN(
        n18124) );
  BUF_X1 U1910 ( .A(n17107), .Z(n25245) );
  INV_X1 U1919 ( .A(n12535), .ZN(n13051) );
  BUF_X1 U1959 ( .A(n9432), .Z(n10890) );
  OR2_X1 U1983 ( .A1(n434), .A2(n25251), .ZN(n7675) );
  INV_X1 U1990 ( .A(n8219), .ZN(n7812) );
  BUF_X1 U1991 ( .A(n8074), .Z(n25253) );
  NAND3_X1 U1999 ( .A1(n1764), .A2(n6816), .A3(n5830), .ZN(n7581) );
  INV_X1 U2007 ( .A(n6699), .ZN(n2008) );
  BUF_X2 U2018 ( .A(Key[45]), .Z(n22986) );
  AND2_X1 U2024 ( .A1(n25550), .A2(n23277), .ZN(n23259) );
  INV_X1 U2052 ( .A(n23905), .ZN(n25239) );
  OAI211_X1 U2054 ( .C1(n22179), .C2(n24369), .A(n22177), .B(n22178), .ZN(
        n24998) );
  AND3_X1 U2076 ( .A1(n22120), .A2(n22119), .A3(n22118), .ZN(n23537) );
  INV_X1 U2082 ( .A(n23858), .ZN(n25240) );
  OR2_X1 U2084 ( .A1(n23201), .A2(n22575), .ZN(n5769) );
  AND3_X1 U2090 ( .A1(n22486), .A2(n4648), .A3(n22485), .ZN(n22528) );
  AND2_X1 U2102 ( .A1(n25299), .A2(n25298), .ZN(n21786) );
  OR2_X1 U2111 ( .A1(n22752), .A2(n211), .ZN(n22569) );
  OR2_X1 U2120 ( .A1(n24924), .A2(n24923), .ZN(n24910) );
  AND2_X1 U2137 ( .A1(n22689), .A2(n22685), .ZN(n25275) );
  INV_X1 U2143 ( .A(n22235), .ZN(n25553) );
  AND2_X1 U2152 ( .A1(n22242), .A2(n22243), .ZN(n22063) );
  AND2_X1 U2188 ( .A1(n22208), .A2(n22064), .ZN(n22066) );
  XNOR2_X1 U2193 ( .A(n25334), .B(n20739), .ZN(n24496) );
  INV_X1 U2196 ( .A(n20740), .ZN(n25334) );
  XNOR2_X1 U2198 ( .A(n21674), .B(n21673), .ZN(n22900) );
  AND3_X1 U2199 ( .A1(n25556), .A2(n20013), .A3(n25555), .ZN(n21160) );
  NOR2_X1 U2200 ( .A1(n20295), .A2(n20294), .ZN(n25470) );
  NAND2_X1 U2247 ( .A1(n5466), .A2(n19123), .ZN(n21541) );
  OAI21_X1 U2265 ( .B1(n20004), .B2(n2864), .A(n1420), .ZN(n25400) );
  NAND3_X1 U2274 ( .A1(n25316), .A2(n20347), .A3(n25315), .ZN(n21334) );
  OR2_X1 U2303 ( .A1(n20328), .A2(n19878), .ZN(n20091) );
  AND2_X1 U2308 ( .A1(n19714), .A2(n20317), .ZN(n19888) );
  NOR2_X1 U2313 ( .A1(n55), .A2(n21008), .ZN(n19668) );
  INV_X1 U2323 ( .A(n21068), .ZN(n25579) );
  OR2_X1 U2325 ( .A1(n20174), .A2(n20588), .ZN(n19952) );
  AND2_X1 U2330 ( .A1(n18212), .A2(n19723), .ZN(n20561) );
  AND2_X1 U2332 ( .A1(n3810), .A2(n3809), .ZN(n24940) );
  OR2_X1 U2344 ( .A1(n18845), .A2(n18844), .ZN(n19851) );
  AOI21_X1 U2367 ( .B1(n19760), .B2(n25540), .A(n25539), .ZN(n2662) );
  INV_X1 U2368 ( .A(n19376), .ZN(n25243) );
  AND2_X1 U2411 ( .A1(n19097), .A2(n4114), .ZN(n19363) );
  INV_X1 U2421 ( .A(n19598), .ZN(n25244) );
  NAND3_X1 U2429 ( .A1(n5103), .A2(n644), .A3(n208), .ZN(n18423) );
  AND2_X1 U2459 ( .A1(n5295), .A2(n16559), .ZN(n18102) );
  NAND2_X1 U2503 ( .A1(n17232), .A2(n1339), .ZN(n18665) );
  OAI211_X1 U2523 ( .C1(n3602), .C2(n16214), .A(n16213), .B(n16212), .ZN(
        n18549) );
  AND2_X1 U2525 ( .A1(n25524), .A2(n16556), .ZN(n2790) );
  INV_X1 U2549 ( .A(n17464), .ZN(n25572) );
  AND3_X1 U2576 ( .A1(n15586), .A2(n25280), .A3(n25279), .ZN(n17069) );
  OR2_X1 U2597 ( .A1(n4624), .A2(n15691), .ZN(n25575) );
  NOR2_X1 U2645 ( .A1(n15693), .A2(n25259), .ZN(n25576) );
  AOI22_X1 U2657 ( .A1(n14352), .A2(n16381), .B1(n15659), .B2(n14351), .ZN(
        n25433) );
  INV_X1 U2675 ( .A(n16303), .ZN(n25272) );
  INV_X1 U2679 ( .A(n16955), .ZN(n25246) );
  AND2_X1 U2683 ( .A1(n16102), .A2(n25586), .ZN(n25585) );
  CLKBUF_X1 U2694 ( .A(n15986), .Z(n25492) );
  OR2_X1 U2704 ( .A1(n4600), .A2(n14101), .ZN(n2002) );
  AND2_X1 U2708 ( .A1(n25570), .A2(n4497), .ZN(n13969) );
  NAND3_X1 U2747 ( .A1(n2436), .A2(n2438), .A3(n25592), .ZN(n14150) );
  INV_X1 U2774 ( .A(n14054), .ZN(n25247) );
  OAI21_X1 U2785 ( .B1(n13661), .B2(n13663), .A(n13662), .ZN(n13485) );
  OR2_X1 U2787 ( .A1(n12733), .A2(n12728), .ZN(n137) );
  OR2_X1 U2801 ( .A1(n12206), .A2(n24617), .ZN(n13662) );
  XNOR2_X1 U2820 ( .A(n11656), .B(n25541), .ZN(n24601) );
  INV_X1 U2830 ( .A(n12914), .ZN(n25248) );
  AND2_X1 U2867 ( .A1(n24856), .A2(n5516), .ZN(n25396) );
  BUF_X2 U2879 ( .A(n12368), .Z(n25371) );
  AND2_X1 U2895 ( .A1(n9333), .A2(n9332), .ZN(n11112) );
  INV_X1 U2908 ( .A(n11128), .ZN(n25249) );
  INV_X1 U2909 ( .A(n11117), .ZN(n10868) );
  AND3_X1 U2943 ( .A1(n711), .A2(n471), .A3(n25341), .ZN(n11046) );
  OAI21_X1 U2956 ( .B1(n10043), .B2(n10042), .A(n10041), .ZN(n11069) );
  BUF_X2 U2976 ( .A(n10336), .Z(n25250) );
  AND3_X1 U2980 ( .A1(n24104), .A2(n5741), .A3(n5334), .ZN(n11117) );
  OR2_X1 U2982 ( .A1(n9281), .A2(n8141), .ZN(n9203) );
  XNOR2_X1 U2987 ( .A(n8822), .B(n8823), .ZN(n9729) );
  AND2_X1 U3001 ( .A1(n25538), .A2(n7219), .ZN(n8336) );
  NAND2_X1 U3012 ( .A1(n25319), .A2(n2217), .ZN(n7813) );
  BUF_X2 U3013 ( .A(n263), .Z(n25251) );
  OR2_X1 U3039 ( .A1(n6366), .A2(n6365), .ZN(n25527) );
  AOI21_X1 U3041 ( .B1(n6879), .B2(n2976), .A(n2045), .ZN(n7449) );
  INV_X1 U3051 ( .A(n7581), .ZN(n7879) );
  INV_X1 U3069 ( .A(n7771), .ZN(n25252) );
  INV_X1 U3072 ( .A(n6686), .ZN(n6977) );
  BUF_X2 U3113 ( .A(n6919), .Z(n24037) );
  XNOR2_X1 U3116 ( .A(n5873), .B(Key[56]), .ZN(n6686) );
  OR2_X1 U3118 ( .A1(n6301), .A2(n6489), .ZN(n6305) );
  XNOR2_X1 U3126 ( .A(Key[35]), .B(Plaintext[35]), .ZN(n25437) );
  AND2_X1 U3137 ( .A1(n6010), .A2(n7609), .ZN(n25277) );
  OR2_X1 U3141 ( .A1(n6398), .A2(n6730), .ZN(n2841) );
  BUF_X1 U3158 ( .A(n6122), .Z(n6990) );
  BUF_X1 U3211 ( .A(n7327), .Z(n248) );
  OR2_X1 U3228 ( .A1(n6551), .A2(n6860), .ZN(n25305) );
  OR2_X1 U3266 ( .A1(n7862), .A2(n7864), .ZN(n25535) );
  OAI211_X1 U3270 ( .C1(n6070), .C2(n1975), .A(n1974), .B(n1973), .ZN(n8604)
         );
  OR2_X1 U3315 ( .A1(n9603), .A2(n9599), .ZN(n9930) );
  BUF_X1 U3329 ( .A(n10018), .Z(n24495) );
  BUF_X1 U3345 ( .A(n9997), .Z(n246) );
  CLKBUF_X1 U3350 ( .A(n9898), .Z(n24054) );
  INV_X1 U3379 ( .A(n714), .ZN(n10306) );
  AND3_X1 U3387 ( .A1(n9326), .A2(n10082), .A3(n10079), .ZN(n10871) );
  OR2_X1 U3389 ( .A1(n9986), .A2(n9985), .ZN(n25341) );
  NAND3_X1 U3392 ( .A1(n9552), .A2(n1399), .A3(n9551), .ZN(n10746) );
  INV_X1 U3399 ( .A(n10371), .ZN(n25507) );
  OAI211_X1 U3400 ( .C1(n7839), .C2(n9346), .A(n848), .B(n847), .ZN(n11005) );
  OR2_X1 U3411 ( .A1(n11112), .A2(n11117), .ZN(n10725) );
  INV_X1 U3459 ( .A(n10728), .ZN(n10481) );
  AND2_X1 U3466 ( .A1(n10574), .A2(n11038), .ZN(n991) );
  NOR2_X1 U3469 ( .A1(n408), .A2(n13057), .ZN(n25551) );
  XNOR2_X1 U3482 ( .A(n12104), .B(n25257), .ZN(n4568) );
  XNOR2_X1 U3486 ( .A(n11637), .B(n11638), .ZN(n12132) );
  XNOR2_X1 U3518 ( .A(n11713), .B(n11712), .ZN(n12914) );
  OR2_X1 U3564 ( .A1(n13056), .A2(n12795), .ZN(n25336) );
  INV_X1 U3579 ( .A(n11655), .ZN(n25541) );
  OAI211_X1 U3590 ( .C1(n13365), .C2(n12980), .A(n13366), .B(n25301), .ZN(
        n1316) );
  BUF_X1 U3593 ( .A(n13039), .Z(n12799) );
  XNOR2_X1 U3605 ( .A(n11904), .B(n11903), .ZN(n12945) );
  AND2_X1 U3613 ( .A1(n14194), .A2(n25360), .ZN(n13478) );
  OR2_X1 U3620 ( .A1(n1579), .A2(n3755), .ZN(n25537) );
  OR2_X1 U3661 ( .A1(n14082), .A2(n14083), .ZN(n25504) );
  AND2_X1 U3663 ( .A1(n14419), .A2(n628), .ZN(n15451) );
  NAND2_X1 U3689 ( .A1(n13715), .A2(n25321), .ZN(n14671) );
  OR2_X1 U3705 ( .A1(n16101), .A2(n16100), .ZN(n15579) );
  CLKBUF_X1 U3745 ( .A(n16008), .Z(n25410) );
  XNOR2_X1 U3749 ( .A(n25518), .B(n15168), .ZN(n14699) );
  AND2_X1 U3790 ( .A1(n1365), .A2(n15802), .ZN(n25294) );
  INV_X1 U3807 ( .A(n16462), .ZN(n25596) );
  CLKBUF_X1 U3808 ( .A(n15470), .Z(n15546) );
  BUF_X1 U3817 ( .A(n16451), .Z(n257) );
  CLKBUF_X1 U3821 ( .A(n16470), .Z(n24550) );
  OR2_X1 U3825 ( .A1(n16422), .A2(n15958), .ZN(n25591) );
  INV_X1 U3846 ( .A(n940), .ZN(n16404) );
  AND2_X1 U3850 ( .A1(n213), .A2(n25510), .ZN(n25509) );
  OR2_X1 U3851 ( .A1(n17207), .A2(n17015), .ZN(n5510) );
  OR2_X1 U3865 ( .A1(n15546), .A2(n383), .ZN(n16056) );
  CLKBUF_X1 U3886 ( .A(n15656), .Z(n15659) );
  OAI21_X1 U3889 ( .B1(n16193), .B2(n25447), .A(n25323), .ZN(n5414) );
  AND2_X1 U3917 ( .A1(n25213), .A2(n16989), .ZN(n16769) );
  OAI21_X1 U3930 ( .B1(n16280), .B2(n4092), .A(n5336), .ZN(n16561) );
  CLKBUF_X1 U3935 ( .A(n17352), .Z(n25491) );
  OAI211_X1 U3993 ( .C1(n4972), .C2(n16472), .A(n16056), .B(n25356), .ZN(
        n17297) );
  OR2_X1 U4017 ( .A1(n376), .A2(n16917), .ZN(n15576) );
  OR2_X1 U4060 ( .A1(n16634), .A2(n24570), .ZN(n638) );
  AND2_X1 U4065 ( .A1(n19472), .A2(n19470), .ZN(n18958) );
  AND3_X1 U4112 ( .A1(n5136), .A2(n1437), .A3(n3993), .ZN(n18435) );
  INV_X1 U4120 ( .A(n4647), .ZN(n19106) );
  INV_X1 U4128 ( .A(n1361), .ZN(n25540) );
  BUF_X1 U4142 ( .A(n17496), .Z(n19327) );
  OR2_X1 U4199 ( .A1(n3470), .A2(n4436), .ZN(n5237) );
  NOR2_X1 U4204 ( .A1(n20317), .A2(n20319), .ZN(n25309) );
  NAND2_X1 U4234 ( .A1(n19258), .A2(n5027), .ZN(n20427) );
  OR2_X1 U4243 ( .A1(n20507), .A2(n20216), .ZN(n25348) );
  OAI21_X1 U4248 ( .B1(n17896), .B2(n17895), .A(n17894), .ZN(n20102) );
  AOI21_X1 U4251 ( .B1(n19116), .B2(n19115), .A(n19114), .ZN(n20516) );
  OAI211_X1 U4268 ( .C1(n18773), .C2(n353), .A(n4458), .B(n4459), .ZN(n20346)
         );
  BUF_X1 U4275 ( .A(n20367), .Z(n24558) );
  AND2_X1 U4285 ( .A1(n25266), .A2(n19668), .ZN(n19673) );
  INV_X1 U4289 ( .A(n20309), .ZN(n20130) );
  OR2_X1 U4290 ( .A1(n20469), .A2(n20062), .ZN(n25302) );
  NAND2_X1 U4291 ( .A1(n4185), .A2(n20267), .ZN(n21172) );
  XNOR2_X1 U4328 ( .A(n21583), .B(n21670), .ZN(n21121) );
  XNOR2_X1 U4340 ( .A(n20903), .B(n2569), .ZN(n5503) );
  INV_X1 U4359 ( .A(n21815), .ZN(n25297) );
  XNOR2_X1 U4396 ( .A(n21244), .B(n21243), .ZN(n22792) );
  OR2_X1 U4400 ( .A1(n333), .A2(n22564), .ZN(n22406) );
  AND2_X1 U4417 ( .A1(n22131), .A2(n22968), .ZN(n25308) );
  BUF_X1 U4454 ( .A(n22139), .Z(n22337) );
  NOR2_X1 U4523 ( .A1(n22185), .A2(n22184), .ZN(n23671) );
  AND2_X1 U4713 ( .A1(n23492), .A2(n23494), .ZN(n25517) );
  OR2_X1 U4744 ( .A1(n23204), .A2(n23203), .ZN(n23208) );
  AOI21_X1 U4745 ( .B1(n22841), .B2(n22840), .A(n22839), .ZN(n24426) );
  AOI21_X1 U4746 ( .B1(n23455), .B2(n23456), .A(n25517), .ZN(n25516) );
  CLKBUF_X1 U4752 ( .A(Key[176]), .Z(n1854) );
  CLKBUF_X1 U4760 ( .A(Key[20]), .Z(n16574) );
  CLKBUF_X1 U4886 ( .A(Key[68]), .Z(n1864) );
  CLKBUF_X1 U4888 ( .A(Key[131]), .Z(n2782) );
  AND2_X1 U4950 ( .A1(n16023), .A2(n15773), .ZN(n25254) );
  OR2_X1 U4983 ( .A1(n19465), .A2(n19464), .ZN(n25255) );
  AND2_X1 U4988 ( .A1(n17242), .A2(n17241), .ZN(n25256) );
  INV_X1 U4992 ( .A(n6034), .ZN(n25325) );
  INV_X1 U4998 ( .A(n20217), .ZN(n25345) );
  XOR2_X1 U4999 ( .A(n12102), .B(n16), .Z(n25257) );
  XNOR2_X1 U5023 ( .A(n11436), .B(n11437), .ZN(n13053) );
  INV_X1 U5034 ( .A(n13053), .ZN(n25337) );
  INV_X1 U5073 ( .A(n13221), .ZN(n25292) );
  INV_X1 U5090 ( .A(n13788), .ZN(n25560) );
  XOR2_X1 U5097 ( .A(n15253), .B(n20690), .Z(n25258) );
  AND2_X1 U5104 ( .A1(n16051), .A2(n4897), .ZN(n25259) );
  INV_X1 U5131 ( .A(n25389), .ZN(n25284) );
  XNOR2_X1 U5163 ( .A(n10882), .B(n10883), .ZN(n13102) );
  INV_X1 U5168 ( .A(n17119), .ZN(n25357) );
  XOR2_X1 U5211 ( .A(n18617), .B(n18618), .Z(n25260) );
  OR2_X1 U5290 ( .A1(n25260), .A2(n19441), .ZN(n25261) );
  AND3_X1 U5310 ( .A1(n17675), .A2(n5456), .A3(n5455), .ZN(n25262) );
  AND2_X1 U5336 ( .A1(n20316), .A2(n19889), .ZN(n25263) );
  AND2_X1 U5355 ( .A1(n24982), .A2(n19578), .ZN(n25264) );
  NAND2_X1 U5375 ( .A1(n19181), .A2(n4792), .ZN(n20215) );
  INV_X1 U5387 ( .A(n20215), .ZN(n25347) );
  AND3_X1 U5400 ( .A1(n25303), .A2(n19642), .A3(n25302), .ZN(n25265) );
  OR2_X1 U5401 ( .A1(n20522), .A2(n20523), .ZN(n25266) );
  NAND2_X1 U5438 ( .A1(n13713), .A2(n13394), .ZN(n1486) );
  XNOR2_X1 U5513 ( .A(n25267), .B(n23729), .ZN(Ciphertext[137]) );
  NAND3_X1 U5588 ( .A1(n23726), .A2(n23725), .A3(n786), .ZN(n25267) );
  NAND2_X1 U5697 ( .A1(n13234), .A2(n13298), .ZN(n2842) );
  XNOR2_X2 U5716 ( .A(n11831), .B(n11830), .ZN(n13298) );
  NAND2_X1 U5721 ( .A1(n25163), .A2(n25164), .ZN(n9309) );
  XNOR2_X1 U5728 ( .A(n25268), .B(n768), .ZN(Ciphertext[120]) );
  NAND2_X1 U5732 ( .A1(n22153), .A2(n22152), .ZN(n25268) );
  OR2_X2 U5749 ( .A1(n25269), .A2(n6821), .ZN(n7985) );
  AOI21_X1 U5759 ( .B1(n6816), .B2(n6817), .A(n6894), .ZN(n25269) );
  NAND2_X1 U5762 ( .A1(n7585), .A2(n7581), .ZN(n7314) );
  OAI21_X2 U5767 ( .B1(n13654), .B2(n1899), .A(n25270), .ZN(n14644) );
  NAND3_X1 U5772 ( .A1(n13657), .A2(n13658), .A3(n13922), .ZN(n25270) );
  NAND2_X1 U5774 ( .A1(n25412), .A2(n16971), .ZN(n16915) );
  NAND3_X1 U5844 ( .A1(n535), .A2(n21294), .A3(n534), .ZN(n22539) );
  NAND2_X1 U5876 ( .A1(n6425), .A2(n5966), .ZN(n6314) );
  OAI211_X2 U5886 ( .C1(n4884), .C2(n4167), .A(n18867), .B(n25271), .ZN(n21008) );
  NAND2_X1 U5936 ( .A1(n18866), .A2(n19113), .ZN(n25271) );
  NAND2_X1 U5950 ( .A1(n4139), .A2(n19112), .ZN(n18865) );
  NOR2_X2 U6035 ( .A1(n17333), .A2(n16602), .ZN(n16917) );
  NAND2_X1 U6082 ( .A1(n24185), .A2(n965), .ZN(n17333) );
  NAND2_X1 U6168 ( .A1(n25272), .A2(n25254), .ZN(n965) );
  NAND2_X1 U6195 ( .A1(n25273), .A2(n16107), .ZN(n969) );
  NAND2_X1 U6207 ( .A1(n15854), .A2(n2478), .ZN(n25273) );
  AND3_X2 U6216 ( .A1(n3481), .A2(n3483), .A3(n3477), .ZN(n21559) );
  NAND2_X1 U6222 ( .A1(n3479), .A2(n3478), .ZN(n3477) );
  NAND2_X1 U6237 ( .A1(n5756), .A2(n16068), .ZN(n15795) );
  NAND2_X1 U6242 ( .A1(n365), .A2(n17633), .ZN(n17475) );
  NAND2_X1 U6261 ( .A1(n15606), .A2(n25274), .ZN(n879) );
  NOR2_X1 U6263 ( .A1(n294), .A2(n16051), .ZN(n25274) );
  NAND2_X1 U6274 ( .A1(n16838), .A2(n25219), .ZN(n16839) );
  NAND4_X1 U6295 ( .A1(n21821), .A2(n21818), .A3(n21820), .A4(n21819), .ZN(
        n21828) );
  NAND2_X1 U6308 ( .A1(n25395), .A2(n25275), .ZN(n21819) );
  OAI21_X1 U6309 ( .B1(n25264), .B2(n25276), .A(n280), .ZN(n1131) );
  NOR2_X1 U6311 ( .A1(n19056), .A2(n19057), .ZN(n25276) );
  NAND3_X1 U6320 ( .A1(n4894), .A2(n13437), .A3(n25445), .ZN(n2003) );
  INV_X1 U6343 ( .A(n1514), .ZN(n22475) );
  NAND2_X1 U6350 ( .A1(n22798), .A2(n22805), .ZN(n1514) );
  NAND2_X1 U6365 ( .A1(n20269), .A2(n20498), .ZN(n61) );
  NAND2_X1 U6413 ( .A1(n19074), .A2(n24700), .ZN(n20269) );
  AOI22_X1 U6425 ( .A1(n14099), .A2(n14211), .B1(n24376), .B2(n14101), .ZN(
        n14217) );
  OAI211_X2 U6444 ( .C1(n13120), .C2(n13119), .A(n2097), .B(n2980), .ZN(n14101) );
  NAND3_X1 U6455 ( .A1(n4927), .A2(n15061), .A3(n15679), .ZN(n564) );
  OR2_X1 U6496 ( .A1(n11109), .A2(n13144), .ZN(n13141) );
  NAND2_X1 U6503 ( .A1(n2555), .A2(n25277), .ZN(n2554) );
  NAND3_X1 U6507 ( .A1(n25278), .A2(n14101), .A3(n13552), .ZN(n4891) );
  INV_X1 U6513 ( .A(n24375), .ZN(n25278) );
  NAND2_X1 U6514 ( .A1(n15585), .A2(n5100), .ZN(n25279) );
  NAND2_X1 U6546 ( .A1(n25587), .A2(n3410), .ZN(n25280) );
  NAND2_X1 U6554 ( .A1(n7760), .A2(n7761), .ZN(n7392) );
  OR2_X2 U6594 ( .A1(n6172), .A2(n5068), .ZN(n7760) );
  NAND2_X1 U6603 ( .A1(n3743), .A2(n15767), .ZN(n16639) );
  NAND2_X1 U6613 ( .A1(n10533), .A2(n11146), .ZN(n714) );
  NAND2_X1 U6667 ( .A1(n24116), .A2(n21010), .ZN(n19972) );
  NAND2_X1 U6668 ( .A1(n21008), .A2(n20290), .ZN(n21010) );
  NAND2_X1 U6708 ( .A1(n23070), .A2(n23071), .ZN(n23073) );
  NAND2_X1 U6786 ( .A1(n20089), .A2(n3480), .ZN(n3479) );
  NAND3_X1 U6809 ( .A1(n20459), .A2(n20461), .A3(n24461), .ZN(n25139) );
  NAND2_X2 U6819 ( .A1(n25281), .A2(n2885), .ZN(n23748) );
  NAND3_X1 U6882 ( .A1(n22248), .A2(n22247), .A3(n22246), .ZN(n25281) );
  NAND2_X1 U6883 ( .A1(n486), .A2(n25282), .ZN(n17832) );
  NAND2_X1 U6884 ( .A1(n25562), .A2(n4683), .ZN(n25282) );
  NAND2_X1 U6928 ( .A1(n23927), .A2(n24948), .ZN(n23928) );
  NAND2_X1 U6951 ( .A1(n2604), .A2(n2093), .ZN(n14786) );
  NAND2_X1 U6960 ( .A1(n15765), .A2(n25283), .ZN(n17081) );
  OAI211_X1 U7022 ( .C1(n16246), .C2(n16247), .A(n25285), .B(n25284), .ZN(
        n25283) );
  NAND2_X1 U7109 ( .A1(n16246), .A2(n25484), .ZN(n25285) );
  XNOR2_X2 U7114 ( .A(n18672), .B(n25286), .ZN(n19173) );
  XNOR2_X1 U7115 ( .A(n18668), .B(n18667), .ZN(n25286) );
  NAND3_X1 U7137 ( .A1(n23205), .A2(n23206), .A3(n2903), .ZN(n23210) );
  NAND2_X1 U7151 ( .A1(n10119), .A2(n10118), .ZN(n11212) );
  AND3_X2 U7152 ( .A1(n1035), .A2(n1036), .A3(n25287), .ZN(n5120) );
  NAND3_X1 U7171 ( .A1(n1032), .A2(n17475), .A3(n1033), .ZN(n25287) );
  NAND2_X2 U7177 ( .A1(n20431), .A2(n5043), .ZN(n21525) );
  AOI21_X1 U7195 ( .B1(n25289), .B2(n25288), .A(n20428), .ZN(n20430) );
  INV_X1 U7261 ( .A(n3047), .ZN(n25288) );
  NAND2_X1 U7265 ( .A1(n19253), .A2(n24943), .ZN(n25289) );
  AND2_X1 U7320 ( .A1(n18959), .A2(n19466), .ZN(n18840) );
  OAI22_X1 U7325 ( .A1(n3646), .A2(n3645), .B1(n17049), .B2(n17052), .ZN(
        n17532) );
  NAND2_X1 U7353 ( .A1(n25378), .A2(n20017), .ZN(n25362) );
  NOR2_X1 U7386 ( .A1(n20137), .A2(n19991), .ZN(n20017) );
  AND2_X2 U7399 ( .A1(n21917), .A2(n22324), .ZN(n22752) );
  OAI21_X1 U7409 ( .B1(n18986), .B2(n3296), .A(n3297), .ZN(n25290) );
  XNOR2_X1 U7416 ( .A(n17839), .B(n17874), .ZN(n24192) );
  NOR2_X2 U7418 ( .A1(n16825), .A2(n807), .ZN(n17839) );
  NAND2_X1 U7446 ( .A1(n25291), .A2(n3098), .ZN(n10653) );
  NAND2_X1 U7447 ( .A1(n10804), .A2(n3100), .ZN(n25291) );
  NAND2_X1 U7448 ( .A1(n4340), .A2(n1544), .ZN(n1539) );
  NAND3_X1 U7459 ( .A1(n20433), .A2(n24940), .A3(n20434), .ZN(n20435) );
  NAND2_X1 U7472 ( .A1(n5208), .A2(n20576), .ZN(n20433) );
  OR3_X1 U7492 ( .A1(n23696), .A2(n22148), .A3(n22082), .ZN(n3441) );
  NAND3_X1 U7501 ( .A1(n25293), .A2(n13222), .A3(n25292), .ZN(n4486) );
  INV_X1 U7504 ( .A(n12919), .ZN(n25293) );
  NAND2_X1 U7518 ( .A1(n656), .A2(n658), .ZN(n6441) );
  NAND2_X1 U7526 ( .A1(n7702), .A2(n7701), .ZN(n8203) );
  NAND2_X1 U7558 ( .A1(n4353), .A2(n25294), .ZN(n15313) );
  XNOR2_X2 U7578 ( .A(n25295), .B(n14994), .ZN(n16225) );
  XNOR2_X1 U7579 ( .A(n14995), .B(n15000), .ZN(n25295) );
  NAND2_X1 U7599 ( .A1(n17338), .A2(n17337), .ZN(n645) );
  NAND2_X1 U7602 ( .A1(n19395), .A2(n19163), .ZN(n19016) );
  NAND3_X1 U7662 ( .A1(n18), .A2(n2258), .A3(n19), .ZN(n17321) );
  OAI21_X1 U7668 ( .B1(n23311), .B2(n23327), .A(n5660), .ZN(n2143) );
  OAI21_X2 U7682 ( .B1(n21788), .B2(n22063), .A(n25296), .ZN(n23769) );
  NAND2_X1 U7689 ( .A1(n21786), .A2(n25297), .ZN(n25296) );
  NAND2_X1 U7691 ( .A1(n22180), .A2(n22239), .ZN(n25298) );
  INV_X1 U7695 ( .A(n22241), .ZN(n25299) );
  NAND2_X1 U7698 ( .A1(n12973), .A2(n25300), .ZN(n14124) );
  OR2_X1 U7715 ( .A1(n12971), .A2(n5412), .ZN(n25300) );
  NAND2_X1 U7745 ( .A1(n17207), .A2(n17216), .ZN(n17210) );
  NAND2_X1 U7804 ( .A1(n12583), .A2(n12980), .ZN(n25301) );
  OAI21_X1 U7817 ( .B1(n19640), .B2(n20471), .A(n20470), .ZN(n25303) );
  XNOR2_X1 U7819 ( .A(n25304), .B(n23448), .ZN(Ciphertext[94]) );
  NAND4_X1 U7820 ( .A1(n23447), .A2(n23446), .A3(n23445), .A4(n23444), .ZN(
        n25304) );
  NAND2_X1 U7884 ( .A1(n16639), .A2(n15557), .ZN(n3744) );
  NAND3_X1 U7916 ( .A1(n1214), .A2(n15912), .A3(n3544), .ZN(n24792) );
  NAND2_X1 U7968 ( .A1(n6550), .A2(n25305), .ZN(n8484) );
  NAND2_X1 U7977 ( .A1(n10628), .A2(n44), .ZN(n25306) );
  NAND2_X1 U8057 ( .A1(n7474), .A2(n7421), .ZN(n7953) );
  AOI21_X1 U8069 ( .B1(n9557), .B2(n9556), .A(n9555), .ZN(n25307) );
  NAND2_X1 U8092 ( .A1(n5529), .A2(n5530), .ZN(n22144) );
  NOR2_X2 U8114 ( .A1(n25308), .A2(n22130), .ZN(n24349) );
  OAI21_X1 U8171 ( .B1(n25263), .B2(n25309), .A(n24917), .ZN(n19892) );
  NAND2_X1 U8183 ( .A1(n25311), .A2(n25310), .ZN(n15976) );
  NAND2_X1 U8207 ( .A1(n15973), .A2(n15970), .ZN(n25310) );
  NAND2_X1 U8226 ( .A1(n746), .A2(n25312), .ZN(n25311) );
  INV_X1 U8238 ( .A(n15973), .ZN(n25312) );
  NAND2_X1 U8242 ( .A1(n22187), .A2(n25313), .ZN(n22192) );
  OR2_X1 U8244 ( .A1(n25070), .A2(n22922), .ZN(n25313) );
  NAND2_X1 U8252 ( .A1(n22712), .A2(n22928), .ZN(n22187) );
  OAI211_X2 U8255 ( .C1(n20248), .C2(n24077), .A(n25314), .B(n20247), .ZN(
        n21087) );
  NAND2_X1 U8265 ( .A1(n24818), .A2(n24077), .ZN(n25314) );
  NAND2_X1 U8269 ( .A1(n9236), .A2(n9757), .ZN(n2268) );
  NAND2_X1 U8273 ( .A1(n2269), .A2(n1814), .ZN(n9236) );
  NAND2_X1 U8305 ( .A1(n22959), .A2(n22958), .ZN(n22034) );
  NOR2_X1 U8322 ( .A1(n7562), .A2(n7725), .ZN(n1596) );
  NAND2_X1 U8348 ( .A1(n7246), .A2(n7563), .ZN(n7562) );
  NOR2_X2 U8351 ( .A1(n23667), .A2(n5508), .ZN(n23670) );
  NAND2_X1 U8366 ( .A1(n22161), .A2(n24768), .ZN(n23667) );
  NAND2_X1 U8380 ( .A1(n19463), .A2(n25255), .ZN(n19494) );
  NAND2_X1 U8391 ( .A1(n24414), .A2(n20343), .ZN(n25315) );
  NAND2_X1 U8411 ( .A1(n3671), .A2(n20344), .ZN(n25316) );
  OAI21_X2 U8419 ( .B1(n15703), .B2(n4552), .A(n25317), .ZN(n18539) );
  NAND3_X1 U8447 ( .A1(n2338), .A2(n15701), .A3(n15700), .ZN(n25317) );
  AOI22_X1 U8460 ( .A1(n19740), .A2(n1667), .B1(n20430), .B2(n5044), .ZN(
        n25318) );
  NAND2_X1 U8462 ( .A1(n25324), .A2(n25327), .ZN(n25319) );
  NAND3_X1 U8509 ( .A1(n16127), .A2(n129), .A3(n24528), .ZN(n17173) );
  OAI21_X1 U8510 ( .B1(n7382), .B2(n7622), .A(n7616), .ZN(n6223) );
  NAND2_X1 U8512 ( .A1(n7618), .A2(n7382), .ZN(n7616) );
  NAND3_X1 U8515 ( .A1(n17287), .A2(n17284), .A3(n16951), .ZN(n24635) );
  INV_X1 U8516 ( .A(n24249), .ZN(n25508) );
  NAND2_X1 U8519 ( .A1(n25320), .A2(n849), .ZN(n16256) );
  NAND3_X1 U8528 ( .A1(n15938), .A2(n25389), .A3(n24162), .ZN(n25320) );
  OAI21_X1 U8529 ( .B1(n3031), .B2(n3030), .A(n13394), .ZN(n25321) );
  NAND2_X1 U8540 ( .A1(n7111), .A2(n7112), .ZN(n8891) );
  NAND2_X1 U8543 ( .A1(n22348), .A2(n25395), .ZN(n21821) );
  NAND2_X1 U8570 ( .A1(n16257), .A2(n17216), .ZN(n25524) );
  NOR2_X2 U8607 ( .A1(n25322), .A2(n13872), .ZN(n15120) );
  AOI21_X1 U8609 ( .B1(n3403), .B2(n3400), .A(n5440), .ZN(n25322) );
  NAND2_X1 U8627 ( .A1(n23288), .A2(n23289), .ZN(n23291) );
  NAND2_X1 U8678 ( .A1(n1030), .A2(n25261), .ZN(n19082) );
  NAND2_X1 U8732 ( .A1(n305), .A2(n10850), .ZN(n10272) );
  NAND3_X1 U8749 ( .A1(n24669), .A2(n3826), .A3(n3829), .ZN(n24633) );
  NAND3_X1 U8780 ( .A1(n7945), .A2(n7946), .A3(n7657), .ZN(n7950) );
  INV_X1 U8795 ( .A(n16191), .ZN(n25323) );
  NAND2_X1 U8799 ( .A1(n25326), .A2(n25325), .ZN(n25324) );
  NAND2_X1 U8801 ( .A1(n6499), .A2(n6434), .ZN(n25326) );
  NAND2_X1 U8821 ( .A1(n6353), .A2(n6034), .ZN(n25327) );
  NAND2_X1 U8831 ( .A1(n25328), .A2(n3410), .ZN(n2076) );
  NAND2_X1 U8846 ( .A1(n15579), .A2(n15582), .ZN(n25328) );
  NAND2_X1 U8851 ( .A1(n556), .A2(n9587), .ZN(n10612) );
  OAI21_X2 U8856 ( .B1(n138), .B2(n16242), .A(n25329), .ZN(n16578) );
  NAND2_X1 U8878 ( .A1(n24294), .A2(n24292), .ZN(n25329) );
  OAI22_X1 U8885 ( .A1(n5020), .A2(n25330), .B1(n14192), .B2(n14191), .ZN(
        n14197) );
  NAND2_X1 U8886 ( .A1(n24186), .A2(n14191), .ZN(n25330) );
  NAND2_X1 U8887 ( .A1(n1694), .A2(n4446), .ZN(n17) );
  NAND2_X1 U8892 ( .A1(n25331), .A2(n4823), .ZN(n12962) );
  NAND2_X1 U8922 ( .A1(n4822), .A2(n399), .ZN(n25331) );
  XNOR2_X1 U8950 ( .A(n15252), .B(n25258), .ZN(n15256) );
  NAND3_X1 U8996 ( .A1(n1275), .A2(n1272), .A3(n1273), .ZN(n25147) );
  XNOR2_X1 U8998 ( .A(n25332), .B(n22301), .ZN(Ciphertext[45]) );
  NAND3_X1 U9003 ( .A1(n188), .A2(n2083), .A3(n22299), .ZN(n25332) );
  OAI22_X1 U9025 ( .A1(n14270), .A2(n14271), .B1(n14273), .B2(n24368), .ZN(
        n14277) );
  NAND2_X1 U9027 ( .A1(n14344), .A2(n3059), .ZN(n24701) );
  XNOR2_X1 U9036 ( .A(n25333), .B(n17868), .ZN(n17871) );
  XNOR2_X1 U9038 ( .A(n17866), .B(n18601), .ZN(n25333) );
  NAND2_X1 U9102 ( .A1(n5404), .A2(n19678), .ZN(n21336) );
  NAND3_X2 U9135 ( .A1(n3801), .A2(n3802), .A3(n13967), .ZN(n15153) );
  NAND3_X1 U9187 ( .A1(n715), .A2(n973), .A3(n25335), .ZN(n14324) );
  NAND3_X1 U9236 ( .A1(n25337), .A2(n13057), .A3(n25336), .ZN(n25335) );
  NAND2_X1 U9238 ( .A1(n22941), .A2(n22940), .ZN(n21654) );
  NAND2_X1 U9256 ( .A1(n17559), .A2(n19264), .ZN(n3470) );
  XNOR2_X2 U9259 ( .A(n3852), .B(n3853), .ZN(n19413) );
  INV_X1 U9262 ( .A(n22483), .ZN(n25569) );
  NAND3_X1 U9263 ( .A1(n10481), .A2(n10482), .A3(n10262), .ZN(n10267) );
  NAND2_X1 U9296 ( .A1(n13744), .A2(n14168), .ZN(n14171) );
  NAND2_X2 U9323 ( .A1(n1783), .A2(n12446), .ZN(n13744) );
  NAND2_X1 U9343 ( .A1(n25338), .A2(n17374), .ZN(n17874) );
  NAND2_X1 U9344 ( .A1(n3693), .A2(n5522), .ZN(n25338) );
  NAND2_X1 U9345 ( .A1(n17574), .A2(n373), .ZN(n17370) );
  OAI21_X1 U9380 ( .B1(n7615), .B2(n7382), .A(n25339), .ZN(n7383) );
  NAND2_X1 U9382 ( .A1(n7382), .A2(n7380), .ZN(n25339) );
  NAND3_X1 U9398 ( .A1(n1217), .A2(n410), .A3(n1219), .ZN(n1215) );
  NAND3_X1 U9406 ( .A1(n25340), .A2(n1478), .A3(n22188), .ZN(n2456) );
  NAND2_X1 U9410 ( .A1(n22107), .A2(n25070), .ZN(n25340) );
  NAND2_X1 U9411 ( .A1(n25342), .A2(n24267), .ZN(n16724) );
  NAND2_X1 U9526 ( .A1(n16720), .A2(n17059), .ZN(n25342) );
  AND2_X2 U9556 ( .A1(n25343), .A2(n24272), .ZN(n19939) );
  NAND2_X1 U9559 ( .A1(n19308), .A2(n19307), .ZN(n25343) );
  NAND2_X1 U9596 ( .A1(n4328), .A2(n25344), .ZN(n20804) );
  NAND3_X1 U9643 ( .A1(n25348), .A2(n25346), .A3(n25345), .ZN(n25344) );
  NAND2_X1 U9645 ( .A1(n25347), .A2(n20507), .ZN(n25346) );
  NAND2_X1 U9689 ( .A1(n24910), .A2(n23967), .ZN(n22693) );
  NAND3_X1 U9712 ( .A1(n2600), .A2(n6686), .A3(n24579), .ZN(n5876) );
  NAND3_X1 U9812 ( .A1(n6721), .A2(n1609), .A3(n6720), .ZN(n6726) );
  NAND2_X1 U9813 ( .A1(n16367), .A2(n16206), .ZN(n16365) );
  NAND2_X1 U9849 ( .A1(n19469), .A2(n19470), .ZN(n458) );
  NAND2_X1 U9854 ( .A1(n19466), .A2(n19321), .ZN(n19469) );
  NAND2_X1 U9859 ( .A1(n11085), .A2(n10438), .ZN(n10221) );
  OR3_X1 U9873 ( .A1(n9459), .A2(n9918), .A3(n9463), .ZN(n9135) );
  NAND3_X1 U9874 ( .A1(n1968), .A2(n13994), .A3(n13993), .ZN(n1966) );
  NAND3_X1 U9889 ( .A1(n16998), .A2(n24471), .A3(n374), .ZN(n15994) );
  NAND3_X1 U9951 ( .A1(n19374), .A2(n19373), .A3(n25349), .ZN(n19774) );
  NAND2_X1 U9979 ( .A1(n19363), .A2(n25243), .ZN(n25349) );
  NAND4_X2 U10008 ( .A1(n2425), .A2(n19776), .A3(n2427), .A4(n2426), .ZN(
        n21267) );
  NOR2_X2 U10023 ( .A1(n20044), .A2(n20045), .ZN(n4294) );
  BUF_X1 U10027 ( .A(n12439), .Z(n13064) );
  AND2_X1 U10057 ( .A1(n22715), .A2(n22927), .ZN(n25557) );
  NAND3_X1 U10069 ( .A1(n10694), .A2(n11057), .A3(n11053), .ZN(n3209) );
  NAND2_X2 U10146 ( .A1(n25350), .A2(n12432), .ZN(n14165) );
  NAND3_X1 U10147 ( .A1(n2192), .A2(n12429), .A3(n12430), .ZN(n25350) );
  NAND3_X1 U10161 ( .A1(n1895), .A2(n7384), .A3(n7380), .ZN(n7201) );
  NAND2_X1 U10196 ( .A1(n4181), .A2(n25351), .ZN(n1268) );
  NAND2_X1 U10220 ( .A1(n13114), .A2(n12660), .ZN(n25351) );
  NAND2_X1 U10239 ( .A1(n17172), .A2(n17522), .ZN(n17176) );
  NAND2_X1 U10247 ( .A1(n17170), .A2(n17171), .ZN(n17172) );
  NAND3_X1 U10267 ( .A1(n3283), .A2(n23716), .A3(n23723), .ZN(n3280) );
  NAND2_X1 U10280 ( .A1(n3888), .A2(n2684), .ZN(n2683) );
  NAND3_X1 U10348 ( .A1(n17353), .A2(n4840), .A3(n4004), .ZN(n16673) );
  NAND2_X1 U10361 ( .A1(n25354), .A2(n25352), .ZN(n12599) );
  NAND2_X1 U10395 ( .A1(n25353), .A2(n13292), .ZN(n25352) );
  MUX2_X1 U10397 ( .A(n12911), .B(n13288), .S(n12593), .Z(n25353) );
  NAND2_X1 U10420 ( .A1(n25355), .A2(n12596), .ZN(n25354) );
  INV_X1 U10455 ( .A(n13292), .ZN(n25355) );
  NAND3_X2 U10458 ( .A1(n24628), .A2(n10624), .A3(n10625), .ZN(n12370) );
  OAI211_X1 U10478 ( .C1(n16472), .C2(n16473), .A(n16469), .B(n24550), .ZN(
        n25356) );
  AND3_X2 U10483 ( .A1(n21279), .A2(n5765), .A3(n4079), .ZN(n23066) );
  NAND3_X1 U10563 ( .A1(n25358), .A2(n2580), .A3(n25357), .ZN(n17105) );
  INV_X1 U10581 ( .A(n17100), .ZN(n25358) );
  NAND3_X2 U10596 ( .A1(n687), .A2(n16536), .A3(n686), .ZN(n18451) );
  XNOR2_X1 U10664 ( .A(n25359), .B(n451), .ZN(Ciphertext[83]) );
  NAND3_X1 U10673 ( .A1(n25142), .A2(n25141), .A3(n22884), .ZN(n25359) );
  XNOR2_X2 U10692 ( .A(n18236), .B(n18235), .ZN(n19186) );
  NAND2_X1 U10697 ( .A1(n10162), .A2(n10161), .ZN(n8417) );
  INV_X1 U10712 ( .A(n14189), .ZN(n25360) );
  NAND2_X1 U10721 ( .A1(n13785), .A2(n14143), .ZN(n14194) );
  OAI21_X1 U10723 ( .B1(n997), .B2(n24063), .A(n25361), .ZN(n22309) );
  NAND2_X1 U10768 ( .A1(n22308), .A2(n24063), .ZN(n25361) );
  OAI211_X2 U10789 ( .C1(n19758), .C2(n19759), .A(n19756), .B(n25362), .ZN(
        n21245) );
  NAND2_X1 U10793 ( .A1(n18768), .A2(n25363), .ZN(n18769) );
  NAND2_X1 U10794 ( .A1(n25364), .A2(n18767), .ZN(n25363) );
  INV_X1 U10806 ( .A(n19307), .ZN(n25364) );
  NAND3_X1 U10808 ( .A1(n12477), .A2(n13041), .A3(n12797), .ZN(n12480) );
  NAND2_X1 U10809 ( .A1(n13039), .A2(n13038), .ZN(n12797) );
  NAND2_X1 U10838 ( .A1(n24118), .A2(n4520), .ZN(n25548) );
  NAND2_X1 U10840 ( .A1(n19183), .A2(n18597), .ZN(n19426) );
  NAND2_X1 U10895 ( .A1(n4795), .A2(n4793), .ZN(n654) );
  NAND3_X1 U10911 ( .A1(n24344), .A2(n18166), .A3(n4647), .ZN(n18167) );
  NAND2_X1 U10949 ( .A1(n19199), .A2(n18809), .ZN(n4647) );
  OAI21_X2 U10966 ( .B1(n17950), .B2(n17949), .A(n17948), .ZN(n21532) );
  OAI21_X2 U10997 ( .B1(n17393), .B2(n3602), .A(n17392), .ZN(n18531) );
  BUF_X1 U11074 ( .A(n23904), .Z(n23896) );
  BUF_X1 U11106 ( .A(n22593), .Z(n24042) );
  OAI21_X1 U11127 ( .B1(n19699), .B2(n24378), .A(n19698), .ZN(n21300) );
  INV_X1 U11137 ( .A(n11159), .ZN(n4737) );
  CLKBUF_X1 U11159 ( .A(n22975), .Z(n25365) );
  XNOR2_X1 U11167 ( .A(n4101), .B(n4100), .ZN(n22975) );
  MUX2_X2 U11169 ( .A(n19848), .B(n19847), .S(n276), .Z(n21660) );
  INV_X1 U11218 ( .A(n12636), .ZN(n25366) );
  OAI21_X1 U11281 ( .B1(n5121), .B2(n20821), .A(n20820), .ZN(n25367) );
  OAI21_X1 U11333 ( .B1(n5121), .B2(n20821), .A(n20820), .ZN(n23228) );
  OR2_X1 U11372 ( .A1(n348), .A2(n20479), .ZN(n1008) );
  OR2_X1 U11375 ( .A1(n21885), .A2(n25368), .ZN(n25175) );
  NAND2_X1 U11407 ( .A1(n22401), .A2(n22400), .ZN(n25368) );
  XNOR2_X2 U11433 ( .A(n19769), .B(n19768), .ZN(n21816) );
  NAND2_X1 U11510 ( .A1(n13028), .A2(n13023), .ZN(n25369) );
  XOR2_X1 U11527 ( .A(n11401), .B(n12381), .Z(n12385) );
  MUX2_X1 U11528 ( .A(n25214), .B(n25058), .S(n17039), .Z(n25370) );
  AND2_X1 U11565 ( .A1(n12934), .A2(n13267), .ZN(n2632) );
  AOI21_X1 U11569 ( .B1(n5711), .B2(n20473), .A(n24704), .ZN(n21173) );
  AOI22_X1 U11571 ( .A1(n10316), .A2(n10661), .B1(n10315), .B2(n10556), .ZN(
        n12368) );
  BUF_X1 U11575 ( .A(n20778), .Z(n25372) );
  AOI21_X1 U11581 ( .B1(n19908), .B2(n19912), .A(n1755), .ZN(n20778) );
  INV_X1 U11599 ( .A(n2869), .ZN(n25373) );
  OR2_X1 U11600 ( .A1(n24908), .A2(n24451), .ZN(n19629) );
  BUF_X1 U11604 ( .A(n18902), .Z(n19275) );
  OR2_X1 U11631 ( .A1(n20491), .A2(n24078), .ZN(n20076) );
  XOR2_X1 U11641 ( .A(n18268), .B(n17110), .Z(n17112) );
  MUX2_X1 U11692 ( .A(n14944), .B(n14945), .S(n2684), .Z(n14948) );
  CLKBUF_X1 U11693 ( .A(n14943), .Z(n25458) );
  AND2_X1 U11784 ( .A1(n5290), .A2(n18765), .ZN(n25374) );
  XNOR2_X1 U11792 ( .A(n20880), .B(n20879), .ZN(n25375) );
  XNOR2_X1 U11793 ( .A(n20880), .B(n20879), .ZN(n22888) );
  OAI21_X1 U11811 ( .B1(n3686), .B2(n13062), .A(n24165), .ZN(n14360) );
  BUF_X1 U11814 ( .A(n2375), .Z(n25376) );
  OAI211_X1 U11815 ( .C1(n20456), .C2(n24357), .A(n24189), .B(n24188), .ZN(
        n25377) );
  XNOR2_X1 U11842 ( .A(n15279), .B(n15278), .ZN(n2375) );
  OAI211_X1 U11846 ( .C1(n20456), .C2(n24357), .A(n24189), .B(n24188), .ZN(
        n21402) );
  INV_X1 U11888 ( .A(n25242), .ZN(n25378) );
  OAI211_X1 U11957 ( .C1(n18974), .C2(n18975), .A(n18973), .B(n18972), .ZN(
        n1629) );
  XNOR2_X1 U11975 ( .A(n20994), .B(n20993), .ZN(n22927) );
  XNOR2_X1 U11977 ( .A(n20863), .B(n20862), .ZN(n22093) );
  OAI211_X1 U12050 ( .C1(n17169), .C2(n2430), .A(n17168), .B(n514), .ZN(n25379) );
  BUF_X1 U12060 ( .A(n23697), .Z(n23715) );
  XNOR2_X1 U12069 ( .A(n20773), .B(n20772), .ZN(n25381) );
  XNOR2_X1 U12096 ( .A(n20773), .B(n20772), .ZN(n22398) );
  AND2_X1 U12105 ( .A1(n23251), .A2(n23242), .ZN(n23235) );
  OR2_X1 U12127 ( .A1(n7045), .A2(n5264), .ZN(n24260) );
  OR2_X1 U12265 ( .A1(n17300), .A2(n16708), .ZN(n3775) );
  XOR2_X1 U12281 ( .A(n21698), .B(n21697), .Z(n25382) );
  XNOR2_X2 U12312 ( .A(n20818), .B(n25222), .ZN(n21697) );
  INV_X1 U12369 ( .A(n22655), .ZN(n22606) );
  AND3_X2 U12482 ( .A1(n3087), .A2(n4102), .A3(n4099), .ZN(n1340) );
  CLKBUF_X1 U12542 ( .A(n20373), .Z(n25383) );
  INV_X1 U12656 ( .A(n20373), .ZN(n20369) );
  INV_X1 U12675 ( .A(n16360), .ZN(n25546) );
  INV_X1 U12725 ( .A(n16105), .ZN(n25587) );
  BUF_X1 U12756 ( .A(n22059), .Z(n22241) );
  NAND3_X1 U12769 ( .A1(n1747), .A2(n1748), .A3(n14224), .ZN(n25384) );
  XOR2_X1 U12822 ( .A(n18109), .B(n18218), .Z(n16760) );
  NAND3_X1 U12864 ( .A1(n1747), .A2(n1748), .A3(n14224), .ZN(n15522) );
  NAND2_X1 U12914 ( .A1(n3076), .A2(n3075), .ZN(n25385) );
  NAND2_X1 U13127 ( .A1(n3076), .A2(n3075), .ZN(n21567) );
  NAND3_X1 U13146 ( .A1(n2724), .A2(n20177), .A3(n2725), .ZN(n25386) );
  NAND3_X1 U13158 ( .A1(n2724), .A2(n20177), .A3(n2725), .ZN(n25387) );
  NAND3_X1 U13193 ( .A1(n2724), .A2(n20177), .A3(n2725), .ZN(n21439) );
  NAND3_X2 U13234 ( .A1(n17675), .A2(n5456), .A3(n5455), .ZN(n25388) );
  OAI211_X1 U13268 ( .C1(n20423), .C2(n20422), .A(n20421), .B(n20420), .ZN(
        n21310) );
  OAI211_X1 U13346 ( .C1(n22847), .C2(n22901), .A(n25568), .B(n22904), .ZN(
        n4648) );
  OR2_X1 U13347 ( .A1(n23147), .A2(n23146), .ZN(n4627) );
  NAND2_X1 U13547 ( .A1(n21190), .A2(n2781), .ZN(n23077) );
  CLKBUF_X1 U13597 ( .A(n9237), .Z(n10031) );
  XNOR2_X1 U13651 ( .A(n14766), .B(n14767), .ZN(n25389) );
  AND3_X1 U13983 ( .A1(n638), .A2(n16632), .A3(n16631), .ZN(n17873) );
  NOR2_X1 U13993 ( .A1(n21291), .A2(n24625), .ZN(n25391) );
  NOR2_X1 U14016 ( .A1(n21291), .A2(n24625), .ZN(n23030) );
  XNOR2_X1 U14021 ( .A(n18008), .B(n18007), .ZN(n25392) );
  XNOR2_X1 U14147 ( .A(n18008), .B(n18007), .ZN(n19360) );
  XNOR2_X1 U14386 ( .A(n8656), .B(n8655), .ZN(n25393) );
  XOR2_X1 U14537 ( .A(n11561), .B(n11646), .Z(n12246) );
  XNOR2_X1 U14560 ( .A(n8656), .B(n8655), .ZN(n10108) );
  OR2_X1 U14577 ( .A1(n19257), .A2(n18831), .ZN(n18055) );
  OAI211_X1 U14588 ( .C1(n12846), .C2(n4241), .A(n2769), .B(n2770), .ZN(n14336) );
  OR2_X1 U14691 ( .A1(n21140), .A2(n22667), .ZN(n22668) );
  AOI21_X1 U14710 ( .B1(n14103), .B2(n4877), .A(n4876), .ZN(n3462) );
  OR2_X1 U14764 ( .A1(n20216), .A2(n20510), .ZN(n20200) );
  XOR2_X1 U14808 ( .A(n19832), .B(n19833), .Z(n25395) );
  AND2_X1 U14842 ( .A1(n24856), .A2(n5516), .ZN(n12003) );
  BUF_X1 U14921 ( .A(n20428), .Z(n25397) );
  AOI22_X1 U15030 ( .A1(n19236), .A2(n19237), .B1(n24310), .B2(n19234), .ZN(
        n20428) );
  XNOR2_X1 U15121 ( .A(Key[14]), .B(Plaintext[14]), .ZN(n25398) );
  XNOR2_X1 U15162 ( .A(Key[14]), .B(Plaintext[14]), .ZN(n6521) );
  OAI211_X1 U15215 ( .C1(n19010), .C2(n19171), .A(n3821), .B(n3820), .ZN(
        n20145) );
  OAI21_X1 U15269 ( .B1(n20608), .B2(n22369), .A(n20607), .ZN(n25399) );
  OAI21_X1 U15301 ( .B1(n20608), .B2(n22369), .A(n20607), .ZN(n23859) );
  OR2_X1 U15308 ( .A1(n22187), .A2(n25557), .ZN(n24782) );
  OAI21_X1 U15462 ( .B1(n20004), .B2(n2864), .A(n1420), .ZN(n21444) );
  XNOR2_X1 U15498 ( .A(n5951), .B(Key[171]), .ZN(n25401) );
  OR2_X2 U15511 ( .A1(n25402), .A2(n25403), .ZN(n7537) );
  AND3_X1 U15586 ( .A1(n6305), .A2(n6303), .A3(n6493), .ZN(n25402) );
  NOR2_X1 U15638 ( .A1(n1561), .A2(n4727), .ZN(n25403) );
  XNOR2_X1 U15656 ( .A(n5951), .B(Key[171]), .ZN(n6427) );
  OR2_X1 U15983 ( .A1(n20248), .A2(n174), .ZN(n679) );
  OAI21_X1 U16070 ( .B1(n22393), .B2(n22858), .A(n22035), .ZN(n23394) );
  AOI22_X2 U16071 ( .A1(n10204), .A2(n4507), .B1(n3443), .B2(n10203), .ZN(
        n12314) );
  XOR2_X1 U16126 ( .A(n5968), .B(Key[175]), .Z(n25404) );
  OR2_X1 U16186 ( .A1(n23672), .A2(n23671), .ZN(n25405) );
  AND2_X1 U16195 ( .A1(n19875), .A2(n20022), .ZN(n20093) );
  AOI21_X1 U16251 ( .B1(n16013), .B2(n16012), .A(n16011), .ZN(n25406) );
  OAI21_X1 U16469 ( .B1(n7199), .B2(n7198), .A(n7197), .ZN(n25407) );
  OAI21_X1 U16586 ( .B1(n7199), .B2(n7198), .A(n7197), .ZN(n8633) );
  XNOR2_X1 U16621 ( .A(n11631), .B(n11630), .ZN(n25408) );
  XNOR2_X1 U16628 ( .A(n14728), .B(n14727), .ZN(n25409) );
  XNOR2_X1 U16641 ( .A(n11631), .B(n11630), .ZN(n13050) );
  BUF_X1 U16692 ( .A(n15657), .Z(n16383) );
  NAND2_X1 U16701 ( .A1(n892), .A2(n539), .ZN(n25411) );
  NAND2_X1 U16705 ( .A1(n892), .A2(n539), .ZN(n18283) );
  BUF_X1 U16754 ( .A(n20475), .Z(n21259) );
  NAND2_X1 U16774 ( .A1(n17662), .A2(n17661), .ZN(n18559) );
  OAI211_X1 U16777 ( .C1(n24370), .C2(n20101), .A(n20100), .B(n20099), .ZN(
        n2010) );
  BUF_X1 U16786 ( .A(n17334), .Z(n25412) );
  OAI211_X1 U16792 ( .C1(n22353), .C2(n22352), .A(n22351), .B(n22350), .ZN(
        n23933) );
  OAI211_X1 U16796 ( .C1(n13591), .C2(n13864), .A(n2417), .B(n5150), .ZN(
        n25413) );
  XNOR2_X1 U16798 ( .A(n21111), .B(n21110), .ZN(n25414) );
  XNOR2_X1 U16812 ( .A(n21110), .B(n21111), .ZN(n23995) );
  XNOR2_X1 U16838 ( .A(n12394), .B(n12395), .ZN(n25415) );
  NOR3_X1 U16896 ( .A1(n12883), .A2(n12882), .A3(n13600), .ZN(n25416) );
  NOR3_X1 U16918 ( .A1(n12883), .A2(n12882), .A3(n13600), .ZN(n25417) );
  XNOR2_X1 U16927 ( .A(n12394), .B(n12395), .ZN(n13344) );
  NOR3_X1 U16947 ( .A1(n12883), .A2(n12882), .A3(n13600), .ZN(n14992) );
  XOR2_X1 U16978 ( .A(n12413), .B(n12207), .Z(n25418) );
  AND2_X1 U16992 ( .A1(n13844), .A2(n13843), .ZN(n1579) );
  XNOR2_X1 U17047 ( .A(n17788), .B(n25419), .ZN(n17794) );
  XOR2_X1 U17059 ( .A(n24488), .B(n2318), .Z(n25419) );
  NAND2_X1 U17075 ( .A1(n4430), .A2(n4429), .ZN(n25420) );
  NAND2_X1 U17178 ( .A1(n4430), .A2(n4429), .ZN(n25421) );
  NAND2_X1 U17227 ( .A1(n4430), .A2(n4429), .ZN(n20413) );
  XNOR2_X1 U17236 ( .A(n18617), .B(n18618), .ZN(n25422) );
  XNOR2_X1 U17257 ( .A(n18617), .B(n18618), .ZN(n25423) );
  XOR2_X1 U17301 ( .A(Key[98]), .B(Plaintext[98]), .Z(n25424) );
  INV_X1 U17334 ( .A(n301), .ZN(n25425) );
  NAND2_X1 U17564 ( .A1(n24734), .A2(n14305), .ZN(n25426) );
  XNOR2_X1 U17617 ( .A(n5936), .B(Key[3]), .ZN(n25427) );
  XNOR2_X1 U17659 ( .A(n5936), .B(Key[3]), .ZN(n25428) );
  INV_X1 U17691 ( .A(n16895), .ZN(n25429) );
  XNOR2_X1 U17730 ( .A(n5936), .B(Key[3]), .ZN(n6513) );
  XNOR2_X1 U17807 ( .A(n12310), .B(n12309), .ZN(n25430) );
  OAI21_X1 U17957 ( .B1(n13604), .B2(n14319), .A(n13603), .ZN(n25431) );
  XNOR2_X1 U18144 ( .A(n12310), .B(n12309), .ZN(n13352) );
  OAI21_X1 U18261 ( .B1(n13604), .B2(n14319), .A(n13603), .ZN(n15521) );
  XOR2_X1 U18333 ( .A(n12783), .B(n12782), .Z(n25432) );
  AOI22_X1 U18334 ( .A1(n14352), .A2(n16381), .B1(n15659), .B2(n14351), .ZN(
        n16955) );
  BUF_X1 U18406 ( .A(n13998), .Z(n25434) );
  BUF_X1 U18464 ( .A(n13998), .Z(n25435) );
  AOI21_X1 U18465 ( .B1(n13342), .B2(n13341), .A(n3126), .ZN(n13998) );
  OAI211_X1 U18467 ( .C1(n13780), .C2(n13779), .A(n4354), .B(n13778), .ZN(
        n25436) );
  OAI211_X1 U18492 ( .C1(n13780), .C2(n13779), .A(n4354), .B(n13778), .ZN(
        n14384) );
  XNOR2_X1 U18495 ( .A(n21984), .B(n21983), .ZN(n25438) );
  XNOR2_X1 U18648 ( .A(Key[35]), .B(Plaintext[35]), .ZN(n5904) );
  XNOR2_X1 U18676 ( .A(n21984), .B(n21983), .ZN(n22838) );
  XNOR2_X1 U18677 ( .A(n21104), .B(n21105), .ZN(n25439) );
  XNOR2_X1 U18678 ( .A(n21104), .B(n21105), .ZN(n23994) );
  OR2_X1 U18695 ( .A1(n10104), .A2(n9773), .ZN(n8643) );
  CLKBUF_X1 U18706 ( .A(n20386), .Z(n25440) );
  XNOR2_X1 U18716 ( .A(n17668), .B(n17667), .ZN(n20386) );
  XNOR2_X1 U18763 ( .A(n15060), .B(n15059), .ZN(n25441) );
  XNOR2_X1 U18788 ( .A(n21573), .B(n21721), .ZN(n25442) );
  XNOR2_X1 U18789 ( .A(n15060), .B(n15059), .ZN(n15746) );
  XNOR2_X2 U18790 ( .A(n15182), .B(n15181), .ZN(n16311) );
  OAI21_X1 U18818 ( .B1(n13885), .B2(n4293), .A(n790), .ZN(n25443) );
  OAI21_X1 U18819 ( .B1(n13885), .B2(n4293), .A(n790), .ZN(n15316) );
  CLKBUF_X1 U18910 ( .A(n9423), .Z(n25444) );
  OR2_X1 U18923 ( .A1(n21008), .A2(n20290), .ZN(n25558) );
  NOR2_X1 U18955 ( .A1(n13099), .A2(n13100), .ZN(n25445) );
  XNOR2_X1 U18966 ( .A(n15414), .B(n15413), .ZN(n25446) );
  NOR2_X1 U18983 ( .A1(n13099), .A2(n13100), .ZN(n24503) );
  AOI22_X2 U19042 ( .A1(n20357), .A2(n20356), .B1(n20355), .B2(n2168), .ZN(
        n21511) );
  XNOR2_X1 U19071 ( .A(n15256), .B(n15257), .ZN(n25447) );
  OAI21_X1 U19072 ( .B1(n18873), .B2(n18874), .A(n18872), .ZN(n20291) );
  INV_X1 U19108 ( .A(n19554), .ZN(n25448) );
  XNOR2_X1 U19109 ( .A(n16698), .B(n16697), .ZN(n19290) );
  XNOR2_X2 U19122 ( .A(n14855), .B(n14856), .ZN(n16465) );
  XNOR2_X1 U19191 ( .A(n14380), .B(n14379), .ZN(n25449) );
  XOR2_X1 U19300 ( .A(n20791), .B(n20790), .Z(n25450) );
  INV_X1 U19329 ( .A(n2624), .ZN(n25451) );
  NOR2_X1 U19330 ( .A1(n21148), .A2(n21149), .ZN(n25452) );
  NOR2_X1 U19383 ( .A1(n21148), .A2(n21149), .ZN(n23065) );
  XNOR2_X1 U19541 ( .A(n8474), .B(n8473), .ZN(n25453) );
  AND3_X2 U19542 ( .A1(n4005), .A2(n5599), .A3(n4003), .ZN(n17817) );
  INV_X1 U19546 ( .A(n20428), .ZN(n276) );
  XOR2_X1 U19549 ( .A(n2797), .B(n8570), .Z(n25454) );
  XNOR2_X1 U19578 ( .A(n2812), .B(n13544), .ZN(n25455) );
  XNOR2_X1 U19593 ( .A(n2812), .B(n13544), .ZN(n16331) );
  NOR2_X1 U19601 ( .A1(n20319), .A2(n25456), .ZN(n17568) );
  NAND2_X1 U19629 ( .A1(n19889), .A2(n19714), .ZN(n25456) );
  OR2_X1 U19635 ( .A1(n6866), .A2(n2404), .ZN(n2965) );
  XNOR2_X1 U19677 ( .A(n8723), .B(n8724), .ZN(n25457) );
  AOI22_X1 U19714 ( .A1(n12644), .A2(n12643), .B1(n12641), .B2(n12642), .ZN(
        n14943) );
  XNOR2_X1 U19729 ( .A(n17937), .B(n17936), .ZN(n25459) );
  INV_X1 U19730 ( .A(n997), .ZN(n25460) );
  BUF_X1 U19868 ( .A(n22220), .Z(n25461) );
  XNOR2_X1 U19876 ( .A(n21305), .B(n21304), .ZN(n22220) );
  INV_X1 U19976 ( .A(n14721), .ZN(n25518) );
  XNOR2_X1 U19985 ( .A(n2577), .B(n5503), .ZN(n25462) );
  XNOR2_X1 U20052 ( .A(n5503), .B(n2577), .ZN(n22782) );
  XNOR2_X1 U20053 ( .A(n9173), .B(n9172), .ZN(n25463) );
  XNOR2_X1 U20070 ( .A(n9173), .B(n9172), .ZN(n10137) );
  CLKBUF_X1 U20317 ( .A(n9554), .Z(n25464) );
  OAI211_X1 U20402 ( .C1(n16199), .C2(n3143), .A(n16201), .B(n3542), .ZN(
        n25465) );
  XOR2_X1 U20446 ( .A(n11786), .B(n11785), .Z(n25466) );
  AND2_X1 U20566 ( .A1(n24863), .A2(n25162), .ZN(n25467) );
  OR2_X1 U20581 ( .A1(n16771), .A2(n17039), .ZN(n25468) );
  XOR2_X1 U20594 ( .A(n18699), .B(n18698), .Z(n25469) );
  CLKBUF_X1 U20609 ( .A(n22449), .Z(n25471) );
  XNOR2_X1 U20628 ( .A(n17658), .B(n17659), .ZN(n25473) );
  XNOR2_X1 U20630 ( .A(n17658), .B(n17659), .ZN(n25474) );
  NOR2_X1 U20707 ( .A1(n15832), .A2(n151), .ZN(n17728) );
  XNOR2_X1 U20727 ( .A(n17658), .B(n17659), .ZN(n19487) );
  INV_X1 U20729 ( .A(n19326), .ZN(n25566) );
  XNOR2_X1 U20788 ( .A(n8838), .B(n8837), .ZN(n25475) );
  AOI21_X1 U20793 ( .B1(n19253), .B2(n24943), .A(n3047), .ZN(n25476) );
  AOI21_X1 U20800 ( .B1(n19253), .B2(n24943), .A(n3047), .ZN(n25477) );
  XNOR2_X1 U20829 ( .A(n8838), .B(n8837), .ZN(n9491) );
  OAI211_X1 U20834 ( .C1(n18726), .C2(n19376), .A(n18725), .B(n4317), .ZN(
        n25478) );
  XOR2_X1 U20857 ( .A(n20988), .B(n20987), .Z(n25479) );
  NAND3_X2 U20858 ( .A1(n2468), .A2(n2467), .A3(n2466), .ZN(n21699) );
  XOR2_X1 U20873 ( .A(Key[165]), .B(Plaintext[165]), .Z(n25480) );
  NOR2_X1 U20904 ( .A1(n4969), .A2(n4528), .ZN(n25481) );
  NOR2_X1 U20929 ( .A1(n4969), .A2(n4528), .ZN(n25482) );
  NOR2_X1 U20942 ( .A1(n4969), .A2(n4528), .ZN(n18628) );
  BUF_X1 U20972 ( .A(n21477), .Z(n25483) );
  OAI211_X1 U20980 ( .C1(n20070), .C2(n20071), .A(n1469), .B(n24722), .ZN(
        n21477) );
  XOR2_X1 U21001 ( .A(n14779), .B(n14778), .Z(n25484) );
  XNOR2_X1 U21031 ( .A(n20908), .B(n5503), .ZN(n25485) );
  XNOR2_X1 U21047 ( .A(n8190), .B(n8189), .ZN(n25486) );
  CLKBUF_X1 U21097 ( .A(n22453), .Z(n25487) );
  OAI21_X1 U21107 ( .B1(n22327), .B2(n22326), .A(n3682), .ZN(n25488) );
  XOR2_X1 U21109 ( .A(n18427), .B(n18426), .Z(n25489) );
  NOR2_X1 U21110 ( .A1(n18791), .A2(n18792), .ZN(n25490) );
  NOR2_X1 U21132 ( .A1(n18791), .A2(n18792), .ZN(n20054) );
  XNOR2_X2 U21133 ( .A(n14717), .B(n14718), .ZN(n16101) );
  AOI21_X2 U21161 ( .B1(n10380), .B2(n4928), .A(n1418), .ZN(n12207) );
  XNOR2_X2 U21175 ( .A(n861), .B(n11926), .ZN(n13318) );
  OAI21_X2 U21191 ( .B1(n3964), .B2(n13729), .A(n3298), .ZN(n15071) );
  OAI211_X1 U21208 ( .C1(n15870), .C2(n16802), .A(n25129), .B(n24685), .ZN(
        n25493) );
  OAI211_X1 U21216 ( .C1(n15870), .C2(n16802), .A(n25129), .B(n24685), .ZN(
        n18636) );
  XOR2_X1 U21253 ( .A(n11605), .B(n11606), .Z(n25494) );
  XNOR2_X1 U21310 ( .A(n21429), .B(n21633), .ZN(n25495) );
  OR3_X1 U21319 ( .A1(n25253), .A2(n7449), .A3(n7917), .ZN(n3346) );
  CLKBUF_X1 U21320 ( .A(n21368), .Z(n25496) );
  INV_X1 U21321 ( .A(n13151), .ZN(n13148) );
  OAI21_X1 U21422 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n25497) );
  NOR2_X1 U21465 ( .A1(n19509), .A2(n19508), .ZN(n25498) );
  NOR2_X1 U21469 ( .A1(n19509), .A2(n19508), .ZN(n21659) );
  XNOR2_X1 U21470 ( .A(n11919), .B(n11918), .ZN(n25499) );
  XNOR2_X1 U21482 ( .A(n13576), .B(n13577), .ZN(n25500) );
  BUF_X1 U21524 ( .A(n15515), .Z(n25501) );
  XOR2_X1 U21525 ( .A(n13939), .B(n13938), .Z(n25502) );
  NAND2_X1 U21561 ( .A1(n1054), .A2(n10895), .ZN(n10898) );
  NAND2_X1 U21591 ( .A1(n14077), .A2(n14075), .ZN(n769) );
  NAND3_X1 U21593 ( .A1(n25505), .A2(n25504), .A3(n25503), .ZN(n15274) );
  NAND2_X1 U21597 ( .A1(n2122), .A2(n14079), .ZN(n25503) );
  NAND2_X1 U21601 ( .A1(n14080), .A2(n12704), .ZN(n25505) );
  OAI21_X1 U21630 ( .B1(n10585), .B2(n25507), .A(n25506), .ZN(n9444) );
  NAND2_X1 U21665 ( .A1(n10585), .A2(n10375), .ZN(n25506) );
  NAND2_X1 U21677 ( .A1(n25509), .A2(n25508), .ZN(n1674) );
  INV_X1 U21701 ( .A(n15625), .ZN(n25510) );
  NAND4_X2 U21717 ( .A1(n5076), .A2(n5075), .A3(n1163), .A4(n1164), .ZN(n23779) );
  NAND3_X1 U21916 ( .A1(n13282), .A2(n24988), .A3(n25191), .ZN(n12610) );
  NAND2_X1 U21933 ( .A1(n23814), .A2(n23815), .ZN(n24630) );
  NAND2_X1 U21954 ( .A1(n18134), .A2(n18135), .ZN(n20328) );
  NAND2_X1 U21983 ( .A1(n25512), .A2(n25511), .ZN(n24879) );
  NAND2_X1 U22002 ( .A1(n5421), .A2(n22038), .ZN(n25511) );
  NAND2_X1 U22016 ( .A1(n22037), .A2(n603), .ZN(n25512) );
  NAND4_X2 U22070 ( .A1(n15313), .A2(n4440), .A3(n15311), .A4(n15312), .ZN(
        n15314) );
  OR2_X1 U22115 ( .A1(n9851), .A2(n9853), .ZN(n8419) );
  NOR2_X1 U22128 ( .A1(n9592), .A2(n10158), .ZN(n9853) );
  OAI21_X1 U22177 ( .B1(n19883), .B2(n25514), .A(n25513), .ZN(n19120) );
  NAND2_X1 U22178 ( .A1(n19883), .A2(n20111), .ZN(n25513) );
  INV_X1 U22230 ( .A(n20109), .ZN(n25514) );
  NAND2_X1 U22339 ( .A1(n5409), .A2(n17425), .ZN(n16644) );
  NOR2_X2 U22361 ( .A1(n1887), .A2(n25515), .ZN(n12241) );
  NAND2_X1 U22497 ( .A1(n4999), .A2(n5000), .ZN(n25515) );
  NAND2_X1 U22541 ( .A1(n22711), .A2(n21020), .ZN(n24781) );
  XNOR2_X1 U22552 ( .A(n25516), .B(n452), .ZN(Ciphertext[96]) );
  OAI21_X2 U22591 ( .B1(n20275), .B2(n20276), .A(n25519), .ZN(n21658) );
  NAND2_X1 U22597 ( .A1(n3520), .A2(n3521), .ZN(n25519) );
  NAND2_X1 U22608 ( .A1(n16138), .A2(n24747), .ZN(n25077) );
  NAND2_X1 U22616 ( .A1(n1836), .A2(n4015), .ZN(n24976) );
  NAND2_X1 U22684 ( .A1(n25523), .A2(n25520), .ZN(n8383) );
  NAND2_X1 U22685 ( .A1(n25522), .A2(n25521), .ZN(n25520) );
  INV_X1 U22687 ( .A(n9837), .ZN(n25521) );
  NAND2_X1 U22688 ( .A1(n421), .A2(n10099), .ZN(n25522) );
  NAND2_X1 U22735 ( .A1(n8381), .A2(n9837), .ZN(n25523) );
  OR2_X1 U22740 ( .A1(n20290), .A2(n20291), .ZN(n24116) );
  XNOR2_X2 U22764 ( .A(n21026), .B(n21243), .ZN(n22243) );
  AOI22_X1 U22801 ( .A1(n23805), .A2(n23003), .B1(n25525), .B2(n23005), .ZN(
        n23006) );
  NOR2_X1 U22844 ( .A1(n2411), .A2(n23790), .ZN(n25525) );
  NAND3_X1 U22897 ( .A1(n10286), .A2(n11112), .A3(n11113), .ZN(n2752) );
  NAND3_X1 U22904 ( .A1(n23681), .A2(n23678), .A3(n23679), .ZN(n23680) );
  NAND2_X1 U22906 ( .A1(n25526), .A2(n15957), .ZN(n18557) );
  NAND3_X1 U22907 ( .A1(n1909), .A2(n284), .A3(n1908), .ZN(n25526) );
  NAND2_X1 U22915 ( .A1(n6364), .A2(n25527), .ZN(n7713) );
  NAND2_X1 U22944 ( .A1(n16461), .A2(n16466), .ZN(n3271) );
  NAND2_X1 U22972 ( .A1(n25529), .A2(n25528), .ZN(n12948) );
  NAND2_X1 U22989 ( .A1(n13317), .A2(n12945), .ZN(n25528) );
  NAND2_X1 U22992 ( .A1(n12946), .A2(n25530), .ZN(n25529) );
  INV_X1 U22994 ( .A(n13317), .ZN(n25530) );
  NAND3_X1 U22998 ( .A1(n13619), .A2(n4771), .A3(n14852), .ZN(n4768) );
  NAND3_X1 U23051 ( .A1(n13054), .A2(n408), .A3(n13055), .ZN(n715) );
  AND3_X2 U23087 ( .A1(n25532), .A2(n22172), .A3(n25531), .ZN(n23689) );
  NAND2_X1 U23115 ( .A1(n4064), .A2(n22918), .ZN(n25531) );
  NAND2_X1 U23116 ( .A1(n4063), .A2(n22170), .ZN(n25532) );
  NAND2_X1 U23147 ( .A1(n20103), .A2(n20102), .ZN(n20099) );
  NAND2_X1 U23312 ( .A1(n746), .A2(n25533), .ZN(n2419) );
  NOR2_X1 U23324 ( .A1(n25502), .A2(n16397), .ZN(n25533) );
  NAND3_X1 U23325 ( .A1(n22454), .A2(n24496), .A3(n22453), .ZN(n2188) );
  NAND3_X1 U23389 ( .A1(n25534), .A2(n3404), .A3(n5256), .ZN(n3369) );
  NAND2_X1 U23396 ( .A1(n14458), .A2(n14317), .ZN(n25534) );
  NAND3_X1 U23532 ( .A1(n4537), .A2(n4534), .A3(n25535), .ZN(n24648) );
  NAND3_X1 U23615 ( .A1(n1238), .A2(n22222), .A3(n1728), .ZN(n24832) );
  NAND2_X1 U23617 ( .A1(n2918), .A2(n12580), .ZN(n12581) );
  NAND3_X1 U23662 ( .A1(n23452), .A2(n23425), .A3(n3242), .ZN(n23447) );
  NAND2_X1 U23756 ( .A1(n5703), .A2(n6984), .ZN(n8499) );
  NAND3_X2 U23757 ( .A1(n25537), .A2(n2955), .A3(n25536), .ZN(n15486) );
  NAND2_X1 U23889 ( .A1(n3533), .A2(n13426), .ZN(n25536) );
  NAND2_X1 U24006 ( .A1(n1744), .A2(n1742), .ZN(n25538) );
  NAND2_X1 U24023 ( .A1(n24144), .A2(n9208), .ZN(n135) );
  NAND2_X1 U24026 ( .A1(n2068), .A2(n19106), .ZN(n2463) );
  OAI21_X1 U24083 ( .B1(n19760), .B2(n18385), .A(n25195), .ZN(n25539) );
  OAI21_X1 U24140 ( .B1(n10453), .B2(n10756), .A(n10452), .ZN(n10454) );
  NAND2_X1 U24141 ( .A1(n10756), .A2(n3324), .ZN(n10452) );
  NAND2_X1 U24142 ( .A1(n24639), .A2(n24642), .ZN(n13538) );
  NAND3_X2 U24150 ( .A1(n4388), .A2(n4387), .A3(n13276), .ZN(n14251) );
  NAND2_X1 U24151 ( .A1(n5047), .A2(n25542), .ZN(n24325) );
  NAND2_X1 U24152 ( .A1(n21379), .A2(n25543), .ZN(n25542) );
  INV_X1 U24169 ( .A(n274), .ZN(n25543) );
  NAND2_X1 U24180 ( .A1(n2394), .A2(n2395), .ZN(n21379) );
  OAI211_X2 U24188 ( .C1(n3642), .C2(n22678), .A(n3640), .B(n25544), .ZN(
        n23967) );
  NAND2_X1 U24189 ( .A1(n22676), .A2(n23997), .ZN(n25544) );
  NAND3_X2 U24203 ( .A1(n3029), .A2(n5492), .A3(n3028), .ZN(n11302) );
  NAND2_X1 U24208 ( .A1(n5049), .A2(n22444), .ZN(n24627) );
  NAND2_X1 U24215 ( .A1(n20093), .A2(n25545), .ZN(n24845) );
  INV_X1 U24216 ( .A(n25220), .ZN(n25545) );
  NAND2_X1 U24224 ( .A1(n23319), .A2(n23317), .ZN(n2668) );
  NAND3_X1 U24228 ( .A1(n1682), .A2(n1684), .A3(n23311), .ZN(n23319) );
  AND3_X2 U24240 ( .A1(n5178), .A2(n5176), .A3(n5177), .ZN(n17171) );
  NAND3_X1 U24244 ( .A1(n3625), .A2(n3624), .A3(n2861), .ZN(n25561) );
  NAND2_X1 U24248 ( .A1(n6730), .A2(n6733), .ZN(n5001) );
  AND2_X2 U24249 ( .A1(n24518), .A2(n24517), .ZN(n23969) );
  NAND2_X1 U24262 ( .A1(n20417), .A2(n20419), .ZN(n20418) );
  NAND3_X1 U24282 ( .A1(n24919), .A2(n24456), .A3(n25546), .ZN(n19) );
  NAND2_X1 U24298 ( .A1(n19006), .A2(n19007), .ZN(n19008) );
  NAND3_X1 U24302 ( .A1(n24664), .A2(n24572), .A3(n14060), .ZN(n4222) );
  NAND2_X1 U24305 ( .A1(n14059), .A2(n14850), .ZN(n14060) );
  NAND3_X2 U24310 ( .A1(n25547), .A2(n10843), .A3(n10842), .ZN(n12381) );
  NAND3_X1 U24316 ( .A1(n2967), .A2(n11135), .A3(n10839), .ZN(n25547) );
  NAND3_X1 U24330 ( .A1(n13307), .A2(n13304), .A3(n12613), .ZN(n4791) );
  NAND3_X2 U24335 ( .A1(n5248), .A2(n5247), .A3(n5825), .ZN(n7882) );
  NAND2_X1 U24336 ( .A1(n6351), .A2(n24466), .ZN(n6504) );
  NOR2_X1 U24337 ( .A1(n25548), .A2(n10925), .ZN(n8180) );
  NAND2_X1 U24345 ( .A1(n14265), .A2(n13426), .ZN(n25549) );
  NAND2_X1 U24346 ( .A1(n22127), .A2(n22126), .ZN(n23277) );
  INV_X1 U24348 ( .A(n23263), .ZN(n25550) );
  AND2_X2 U24349 ( .A1(n3567), .A2(n3618), .ZN(n4400) );
  NAND3_X1 U24350 ( .A1(n6765), .A2(n6766), .A3(n6764), .ZN(n3567) );
  NAND2_X1 U24351 ( .A1(n23069), .A2(n21239), .ZN(n1304) );
  OAI21_X1 U24352 ( .B1(n25552), .B2(n25551), .A(n3065), .ZN(n3064) );
  INV_X1 U24353 ( .A(n12752), .ZN(n25552) );
  NAND2_X1 U24354 ( .A1(n10919), .A2(n10918), .ZN(n10921) );
  OAI21_X1 U24355 ( .B1(n17040), .B2(n25058), .A(n3949), .ZN(n3955) );
  OAI211_X2 U24356 ( .C1(n15893), .C2(n24587), .A(n15892), .B(n15891), .ZN(
        n25058) );
  NAND2_X1 U24357 ( .A1(n20185), .A2(n20191), .ZN(n19662) );
  OR2_X1 U24358 ( .A1(n25485), .A2(n21766), .ZN(n22155) );
  AOI21_X1 U24359 ( .B1(n25554), .B2(n25553), .A(n22231), .ZN(n4397) );
  NAND2_X1 U24360 ( .A1(n22056), .A2(n22226), .ZN(n25554) );
  NAND2_X1 U24361 ( .A1(n20296), .A2(n20142), .ZN(n25555) );
  NAND2_X1 U24362 ( .A1(n20011), .A2(n20301), .ZN(n25556) );
  NAND3_X1 U24363 ( .A1(n20528), .A2(n20525), .A3(n55), .ZN(n20526) );
  OAI21_X1 U24364 ( .B1(n55), .B2(n20528), .A(n25558), .ZN(n3833) );
  NAND2_X1 U24365 ( .A1(n7556), .A2(n25559), .ZN(n9016) );
  NAND2_X1 U24366 ( .A1(n3572), .A2(n3569), .ZN(n25559) );
  NAND3_X1 U24367 ( .A1(n14194), .A2(n13785), .A3(n25560), .ZN(n4202) );
  XNOR2_X1 U24368 ( .A(n17782), .B(n17781), .ZN(n19097) );
  OR2_X2 U24369 ( .A1(n3449), .A2(n15749), .ZN(n2562) );
  NAND3_X1 U24370 ( .A1(n3268), .A2(n7757), .A3(n432), .ZN(n7544) );
  NAND2_X1 U24371 ( .A1(n19522), .A2(n19523), .ZN(n18796) );
  NAND2_X1 U24372 ( .A1(n17028), .A2(n25003), .ZN(n17398) );
  NAND2_X1 U24373 ( .A1(n1069), .A2(n5324), .ZN(n4332) );
  NAND2_X1 U24374 ( .A1(n11112), .A2(n11117), .ZN(n9581) );
  NAND2_X1 U24375 ( .A1(n244), .A2(n16426), .ZN(n15649) );
  AOI22_X1 U24376 ( .A1(n1550), .A2(n20486), .B1(n20485), .B2(n20913), .ZN(
        n20490) );
  AND3_X2 U24377 ( .A1(n3311), .A2(n6778), .A3(n6779), .ZN(n7972) );
  NAND2_X1 U24378 ( .A1(n25561), .A2(n3622), .ZN(n24794) );
  NAND2_X1 U24379 ( .A1(n4686), .A2(n17109), .ZN(n25562) );
  NAND2_X1 U24380 ( .A1(n19332), .A2(n25563), .ZN(n19937) );
  NAND2_X1 U24381 ( .A1(n25565), .A2(n25564), .ZN(n25563) );
  AOI21_X1 U24382 ( .B1(n24516), .B2(n19326), .A(n4291), .ZN(n25564) );
  NAND2_X1 U24383 ( .A1(n19327), .A2(n25566), .ZN(n25565) );
  NAND2_X1 U24384 ( .A1(n25249), .A2(n10714), .ZN(n10293) );
  NAND3_X2 U24385 ( .A1(n9311), .A2(n25567), .A3(n9312), .ZN(n10714) );
  OR2_X1 U24386 ( .A1(n9313), .A2(n9314), .ZN(n25567) );
  NAND2_X1 U24387 ( .A1(n16100), .A2(n16101), .ZN(n5458) );
  XNOR2_X2 U24388 ( .A(n14713), .B(n14712), .ZN(n16100) );
  NAND3_X1 U24389 ( .A1(n23881), .A2(n107), .A3(n23882), .ZN(n24692) );
  NAND3_X1 U24390 ( .A1(n23897), .A2(n23899), .A3(n23898), .ZN(n23901) );
  NAND2_X1 U24391 ( .A1(n24825), .A2(n16072), .ZN(n16133) );
  NAND3_X1 U24392 ( .A1(n4487), .A2(n17255), .A3(n16942), .ZN(n3189) );
  NAND2_X1 U24393 ( .A1(n22901), .A2(n25569), .ZN(n25568) );
  NAND2_X1 U24394 ( .A1(n11837), .A2(n4499), .ZN(n25570) );
  XNOR2_X1 U24395 ( .A(n25571), .B(n21391), .ZN(Ciphertext[21]) );
  NAND3_X1 U24396 ( .A1(n4627), .A2(n4628), .A3(n4626), .ZN(n25571) );
  MUX2_X1 U24397 ( .A(n20567), .B(n20560), .S(n20561), .Z(n20098) );
  NAND3_X1 U24398 ( .A1(n25573), .A2(n2062), .A3(n25572), .ZN(n3993) );
  NAND2_X1 U24399 ( .A1(n2064), .A2(n287), .ZN(n25573) );
  OAI21_X1 U24400 ( .B1(n22426), .B2(n22125), .A(n25574), .ZN(n21876) );
  NAND2_X1 U24401 ( .A1(n24322), .A2(n22422), .ZN(n25574) );
  OR2_X1 U24402 ( .A1(n16365), .A2(n17183), .ZN(n15817) );
  AND2_X2 U24403 ( .A1(n25576), .A2(n25575), .ZN(n16796) );
  NAND2_X2 U24404 ( .A1(n25577), .A2(n2802), .ZN(n19986) );
  NAND3_X1 U24405 ( .A1(n19149), .A2(n19150), .A3(n19266), .ZN(n25577) );
  NAND3_X1 U24406 ( .A1(n5285), .A2(n5287), .A3(n22090), .ZN(Ciphertext[132])
         );
  NAND2_X1 U24407 ( .A1(n25578), .A2(n21067), .ZN(n21071) );
  OAI21_X1 U24408 ( .B1(n21066), .B2(n21065), .A(n25579), .ZN(n25578) );
  NAND3_X1 U24409 ( .A1(n22581), .A2(n4989), .A3(n4990), .ZN(n24789) );
  NAND2_X1 U24410 ( .A1(n21825), .A2(n21822), .ZN(n3856) );
  XNOR2_X2 U24411 ( .A(n18861), .B(n18860), .ZN(n21822) );
  NAND3_X2 U24412 ( .A1(n14238), .A2(n1342), .A3(n1343), .ZN(n15369) );
  NAND2_X1 U24413 ( .A1(n25580), .A2(n24198), .ZN(n8853) );
  NAND2_X1 U24414 ( .A1(n7470), .A2(n25154), .ZN(n25580) );
  NAND2_X1 U24415 ( .A1(n2718), .A2(n15811), .ZN(n42) );
  NAND2_X1 U24416 ( .A1(n24061), .A2(n16403), .ZN(n2718) );
  NAND2_X1 U24417 ( .A1(n10960), .A2(n4998), .ZN(n10963) );
  NAND2_X1 U24418 ( .A1(n25583), .A2(n25581), .ZN(n12628) );
  NAND2_X1 U24419 ( .A1(n13364), .A2(n25582), .ZN(n25581) );
  NOR2_X1 U24420 ( .A1(n12977), .A2(n12980), .ZN(n25582) );
  NAND2_X1 U24421 ( .A1(n25584), .A2(n12624), .ZN(n25583) );
  INV_X1 U24422 ( .A(n13364), .ZN(n25584) );
  NAND2_X1 U24423 ( .A1(n25587), .A2(n25585), .ZN(n16088) );
  INV_X1 U24424 ( .A(n16080), .ZN(n25586) );
  NOR2_X1 U24425 ( .A1(n1737), .A2(n7721), .ZN(n1736) );
  NAND3_X1 U24426 ( .A1(n269), .A2(n8531), .A3(n7087), .ZN(n7089) );
  OAI211_X1 U24427 ( .C1(n16340), .C2(n16339), .A(n25589), .B(n25588), .ZN(
        n16527) );
  NAND2_X1 U24428 ( .A1(n16337), .A2(n16336), .ZN(n25588) );
  NAND2_X1 U24429 ( .A1(n16335), .A2(n16334), .ZN(n25589) );
  NAND2_X1 U24430 ( .A1(n25590), .A2(n6525), .ZN(n7662) );
  NAND3_X1 U24431 ( .A1(n1321), .A2(n1320), .A3(n6520), .ZN(n25590) );
  OAI211_X1 U24432 ( .C1(n15961), .C2(n1329), .A(n16424), .B(n25591), .ZN(
        n17436) );
  NAND3_X1 U24433 ( .A1(n3847), .A2(n3848), .A3(n24487), .ZN(n25592) );
  NAND2_X1 U24434 ( .A1(n4973), .A2(n4755), .ZN(n4751) );
  XNOR2_X1 U24435 ( .A(n25593), .B(n15319), .ZN(n5494) );
  XNOR2_X1 U24436 ( .A(n15317), .B(n15318), .ZN(n25593) );
  NAND3_X1 U24437 ( .A1(n22548), .A2(n25595), .A3(n25594), .ZN(n22550) );
  NAND2_X1 U24438 ( .A1(n22547), .A2(n23906), .ZN(n25594) );
  NAND2_X1 U24439 ( .A1(n22546), .A2(n23879), .ZN(n25595) );
  NOR2_X1 U24440 ( .A1(n19012), .A2(n19689), .ZN(n19020) );
  NAND3_X1 U24441 ( .A1(n16458), .A2(n16459), .A3(n25596), .ZN(n4724) );
  NOR2_X1 U24442 ( .A1(n22224), .A2(n25597), .ZN(n23742) );
  NAND2_X1 U24443 ( .A1(n24832), .A2(n1237), .ZN(n25597) );
  AND2_X2 U24444 ( .A1(n16055), .A2(n16054), .ZN(n16375) );
  NAND2_X1 U24445 ( .A1(n2322), .A2(n20533), .ZN(n3076) );
  NAND2_X1 U24446 ( .A1(n19687), .A2(n19688), .ZN(n2322) );
  OAI211_X2 U24447 ( .C1(n5360), .C2(n12830), .A(n2631), .B(n12608), .ZN(
        n14850) );
  NAND3_X2 U24448 ( .A1(n14396), .A2(n14395), .A3(n14394), .ZN(n17283) );
  AOI22_X2 U24449 ( .A1(n5244), .A2(n20477), .B1(n999), .B2(n18839), .ZN(
        n25073) );
  XNOR2_X2 U24450 ( .A(n22018), .B(n22017), .ZN(n25041) );
  AND2_X2 U24451 ( .A1(n5583), .A2(n5582), .ZN(n24498) );
endmodule


module SPEEDY_Top ( clk, Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFF_X1 \reg_in_reg[191]  ( .D(Plaintext[191]), .CK(clk), .Q(reg_in[191]) );
  DFF_X1 \reg_in_reg[190]  ( .D(Plaintext[190]), .CK(clk), .Q(reg_in[190]) );
  DFF_X1 \reg_in_reg[189]  ( .D(Plaintext[189]), .CK(clk), .Q(reg_in[189]) );
  DFF_X1 \reg_in_reg[188]  ( .D(Plaintext[188]), .CK(clk), .Q(reg_in[188]) );
  DFF_X1 \reg_in_reg[187]  ( .D(Plaintext[187]), .CK(clk), .Q(reg_in[187]) );
  DFF_X1 \reg_in_reg[186]  ( .D(Plaintext[186]), .CK(clk), .Q(reg_in[186]) );
  DFF_X1 \reg_in_reg[185]  ( .D(Plaintext[185]), .CK(clk), .Q(reg_in[185]) );
  DFF_X1 \reg_in_reg[184]  ( .D(Plaintext[184]), .CK(clk), .Q(reg_in[184]) );
  DFF_X1 \reg_in_reg[183]  ( .D(Plaintext[183]), .CK(clk), .Q(reg_in[183]) );
  DFF_X1 \reg_in_reg[182]  ( .D(Plaintext[182]), .CK(clk), .Q(reg_in[182]) );
  DFF_X1 \reg_in_reg[181]  ( .D(Plaintext[181]), .CK(clk), .Q(reg_in[181]) );
  DFF_X1 \reg_in_reg[180]  ( .D(Plaintext[180]), .CK(clk), .Q(reg_in[180]) );
  DFF_X1 \reg_in_reg[179]  ( .D(Plaintext[179]), .CK(clk), .Q(reg_in[179]) );
  DFF_X1 \reg_in_reg[178]  ( .D(Plaintext[178]), .CK(clk), .Q(reg_in[178]) );
  DFF_X1 \reg_in_reg[177]  ( .D(Plaintext[177]), .CK(clk), .Q(reg_in[177]) );
  DFF_X1 \reg_in_reg[176]  ( .D(Plaintext[176]), .CK(clk), .Q(reg_in[176]) );
  DFF_X1 \reg_in_reg[175]  ( .D(Plaintext[175]), .CK(clk), .Q(reg_in[175]) );
  DFF_X1 \reg_in_reg[174]  ( .D(Plaintext[174]), .CK(clk), .Q(reg_in[174]) );
  DFF_X1 \reg_in_reg[173]  ( .D(Plaintext[173]), .CK(clk), .Q(reg_in[173]) );
  DFF_X1 \reg_in_reg[172]  ( .D(Plaintext[172]), .CK(clk), .Q(reg_in[172]) );
  DFF_X1 \reg_in_reg[171]  ( .D(Plaintext[171]), .CK(clk), .Q(reg_in[171]) );
  DFF_X1 \reg_in_reg[170]  ( .D(Plaintext[170]), .CK(clk), .Q(reg_in[170]) );
  DFF_X1 \reg_in_reg[169]  ( .D(Plaintext[169]), .CK(clk), .Q(reg_in[169]) );
  DFF_X1 \reg_in_reg[168]  ( .D(Plaintext[168]), .CK(clk), .Q(reg_in[168]) );
  DFF_X1 \reg_in_reg[167]  ( .D(Plaintext[167]), .CK(clk), .Q(reg_in[167]) );
  DFF_X1 \reg_in_reg[166]  ( .D(Plaintext[166]), .CK(clk), .Q(reg_in[166]) );
  DFF_X1 \reg_in_reg[165]  ( .D(Plaintext[165]), .CK(clk), .Q(reg_in[165]) );
  DFF_X1 \reg_in_reg[164]  ( .D(Plaintext[164]), .CK(clk), .Q(reg_in[164]) );
  DFF_X1 \reg_in_reg[163]  ( .D(Plaintext[163]), .CK(clk), .Q(reg_in[163]) );
  DFF_X1 \reg_in_reg[162]  ( .D(Plaintext[162]), .CK(clk), .Q(reg_in[162]) );
  DFF_X1 \reg_in_reg[161]  ( .D(Plaintext[161]), .CK(clk), .Q(reg_in[161]) );
  DFF_X1 \reg_in_reg[160]  ( .D(Plaintext[160]), .CK(clk), .Q(reg_in[160]) );
  DFF_X1 \reg_in_reg[159]  ( .D(Plaintext[159]), .CK(clk), .Q(reg_in[159]) );
  DFF_X1 \reg_in_reg[158]  ( .D(Plaintext[158]), .CK(clk), .Q(reg_in[158]) );
  DFF_X1 \reg_in_reg[157]  ( .D(Plaintext[157]), .CK(clk), .Q(reg_in[157]) );
  DFF_X1 \reg_in_reg[156]  ( .D(Plaintext[156]), .CK(clk), .Q(reg_in[156]) );
  DFF_X1 \reg_in_reg[155]  ( .D(Plaintext[155]), .CK(clk), .Q(reg_in[155]) );
  DFF_X1 \reg_in_reg[154]  ( .D(Plaintext[154]), .CK(clk), .Q(reg_in[154]) );
  DFF_X1 \reg_in_reg[153]  ( .D(Plaintext[153]), .CK(clk), .Q(reg_in[153]) );
  DFF_X1 \reg_in_reg[152]  ( .D(Plaintext[152]), .CK(clk), .Q(reg_in[152]) );
  DFF_X1 \reg_in_reg[151]  ( .D(Plaintext[151]), .CK(clk), .Q(reg_in[151]) );
  DFF_X1 \reg_in_reg[150]  ( .D(Plaintext[150]), .CK(clk), .Q(reg_in[150]) );
  DFF_X1 \reg_in_reg[149]  ( .D(Plaintext[149]), .CK(clk), .Q(reg_in[149]) );
  DFF_X1 \reg_in_reg[148]  ( .D(Plaintext[148]), .CK(clk), .Q(reg_in[148]) );
  DFF_X1 \reg_in_reg[147]  ( .D(Plaintext[147]), .CK(clk), .Q(reg_in[147]) );
  DFF_X1 \reg_in_reg[146]  ( .D(Plaintext[146]), .CK(clk), .Q(reg_in[146]) );
  DFF_X1 \reg_in_reg[145]  ( .D(Plaintext[145]), .CK(clk), .Q(reg_in[145]) );
  DFF_X1 \reg_in_reg[144]  ( .D(Plaintext[144]), .CK(clk), .Q(reg_in[144]) );
  DFF_X1 \reg_in_reg[143]  ( .D(Plaintext[143]), .CK(clk), .Q(reg_in[143]) );
  DFF_X1 \reg_in_reg[142]  ( .D(Plaintext[142]), .CK(clk), .Q(reg_in[142]) );
  DFF_X1 \reg_in_reg[141]  ( .D(Plaintext[141]), .CK(clk), .Q(reg_in[141]) );
  DFF_X1 \reg_in_reg[140]  ( .D(Plaintext[140]), .CK(clk), .Q(reg_in[140]) );
  DFF_X1 \reg_in_reg[139]  ( .D(Plaintext[139]), .CK(clk), .Q(reg_in[139]) );
  DFF_X1 \reg_in_reg[138]  ( .D(Plaintext[138]), .CK(clk), .Q(reg_in[138]) );
  DFF_X1 \reg_in_reg[137]  ( .D(Plaintext[137]), .CK(clk), .Q(reg_in[137]) );
  DFF_X1 \reg_in_reg[136]  ( .D(Plaintext[136]), .CK(clk), .Q(reg_in[136]) );
  DFF_X1 \reg_in_reg[135]  ( .D(Plaintext[135]), .CK(clk), .Q(reg_in[135]) );
  DFF_X1 \reg_in_reg[134]  ( .D(Plaintext[134]), .CK(clk), .Q(reg_in[134]) );
  DFF_X1 \reg_in_reg[133]  ( .D(Plaintext[133]), .CK(clk), .Q(reg_in[133]) );
  DFF_X1 \reg_in_reg[132]  ( .D(Plaintext[132]), .CK(clk), .Q(reg_in[132]) );
  DFF_X1 \reg_in_reg[131]  ( .D(Plaintext[131]), .CK(clk), .Q(reg_in[131]) );
  DFF_X1 \reg_in_reg[130]  ( .D(Plaintext[130]), .CK(clk), .Q(reg_in[130]) );
  DFF_X1 \reg_in_reg[129]  ( .D(Plaintext[129]), .CK(clk), .Q(reg_in[129]) );
  DFF_X1 \reg_in_reg[128]  ( .D(Plaintext[128]), .CK(clk), .Q(reg_in[128]) );
  DFF_X1 \reg_in_reg[127]  ( .D(Plaintext[127]), .CK(clk), .Q(reg_in[127]) );
  DFF_X1 \reg_in_reg[126]  ( .D(Plaintext[126]), .CK(clk), .Q(reg_in[126]) );
  DFF_X1 \reg_in_reg[125]  ( .D(Plaintext[125]), .CK(clk), .Q(reg_in[125]) );
  DFF_X1 \reg_in_reg[124]  ( .D(Plaintext[124]), .CK(clk), .Q(reg_in[124]) );
  DFF_X1 \reg_in_reg[123]  ( .D(Plaintext[123]), .CK(clk), .Q(reg_in[123]) );
  DFF_X1 \reg_in_reg[122]  ( .D(Plaintext[122]), .CK(clk), .Q(reg_in[122]) );
  DFF_X1 \reg_in_reg[121]  ( .D(Plaintext[121]), .CK(clk), .Q(reg_in[121]) );
  DFF_X1 \reg_in_reg[120]  ( .D(Plaintext[120]), .CK(clk), .Q(reg_in[120]) );
  DFF_X1 \reg_in_reg[119]  ( .D(Plaintext[119]), .CK(clk), .Q(reg_in[119]) );
  DFF_X1 \reg_in_reg[118]  ( .D(Plaintext[118]), .CK(clk), .Q(reg_in[118]) );
  DFF_X1 \reg_in_reg[117]  ( .D(Plaintext[117]), .CK(clk), .Q(reg_in[117]) );
  DFF_X1 \reg_in_reg[116]  ( .D(Plaintext[116]), .CK(clk), .Q(reg_in[116]) );
  DFF_X1 \reg_in_reg[115]  ( .D(Plaintext[115]), .CK(clk), .Q(reg_in[115]) );
  DFF_X1 \reg_in_reg[114]  ( .D(Plaintext[114]), .CK(clk), .Q(reg_in[114]) );
  DFF_X1 \reg_in_reg[113]  ( .D(Plaintext[113]), .CK(clk), .Q(reg_in[113]) );
  DFF_X1 \reg_in_reg[112]  ( .D(Plaintext[112]), .CK(clk), .Q(reg_in[112]) );
  DFF_X1 \reg_in_reg[111]  ( .D(Plaintext[111]), .CK(clk), .Q(reg_in[111]) );
  DFF_X1 \reg_in_reg[110]  ( .D(Plaintext[110]), .CK(clk), .Q(reg_in[110]) );
  DFF_X1 \reg_in_reg[109]  ( .D(Plaintext[109]), .CK(clk), .Q(reg_in[109]) );
  DFF_X1 \reg_in_reg[108]  ( .D(Plaintext[108]), .CK(clk), .Q(reg_in[108]) );
  DFF_X1 \reg_in_reg[107]  ( .D(Plaintext[107]), .CK(clk), .Q(reg_in[107]) );
  DFF_X1 \reg_in_reg[106]  ( .D(Plaintext[106]), .CK(clk), .Q(reg_in[106]) );
  DFF_X1 \reg_in_reg[105]  ( .D(Plaintext[105]), .CK(clk), .Q(reg_in[105]) );
  DFF_X1 \reg_in_reg[104]  ( .D(Plaintext[104]), .CK(clk), .Q(reg_in[104]) );
  DFF_X1 \reg_in_reg[103]  ( .D(Plaintext[103]), .CK(clk), .Q(reg_in[103]) );
  DFF_X1 \reg_in_reg[102]  ( .D(Plaintext[102]), .CK(clk), .Q(reg_in[102]) );
  DFF_X1 \reg_in_reg[101]  ( .D(Plaintext[101]), .CK(clk), .Q(reg_in[101]) );
  DFF_X1 \reg_in_reg[100]  ( .D(Plaintext[100]), .CK(clk), .Q(reg_in[100]) );
  DFF_X1 \reg_in_reg[99]  ( .D(Plaintext[99]), .CK(clk), .Q(reg_in[99]) );
  DFF_X1 \reg_in_reg[98]  ( .D(Plaintext[98]), .CK(clk), .Q(reg_in[98]) );
  DFF_X1 \reg_in_reg[97]  ( .D(Plaintext[97]), .CK(clk), .Q(reg_in[97]) );
  DFF_X1 \reg_in_reg[96]  ( .D(Plaintext[96]), .CK(clk), .Q(reg_in[96]) );
  DFF_X1 \reg_in_reg[95]  ( .D(Plaintext[95]), .CK(clk), .Q(reg_in[95]) );
  DFF_X1 \reg_in_reg[94]  ( .D(Plaintext[94]), .CK(clk), .Q(reg_in[94]) );
  DFF_X1 \reg_in_reg[93]  ( .D(Plaintext[93]), .CK(clk), .Q(reg_in[93]) );
  DFF_X1 \reg_in_reg[92]  ( .D(Plaintext[92]), .CK(clk), .Q(reg_in[92]) );
  DFF_X1 \reg_in_reg[91]  ( .D(Plaintext[91]), .CK(clk), .Q(reg_in[91]) );
  DFF_X1 \reg_in_reg[90]  ( .D(Plaintext[90]), .CK(clk), .Q(reg_in[90]) );
  DFF_X1 \reg_in_reg[89]  ( .D(Plaintext[89]), .CK(clk), .Q(reg_in[89]) );
  DFF_X1 \reg_in_reg[88]  ( .D(Plaintext[88]), .CK(clk), .Q(reg_in[88]) );
  DFF_X1 \reg_in_reg[87]  ( .D(Plaintext[87]), .CK(clk), .Q(reg_in[87]) );
  DFF_X1 \reg_in_reg[86]  ( .D(Plaintext[86]), .CK(clk), .Q(reg_in[86]) );
  DFF_X1 \reg_in_reg[85]  ( .D(Plaintext[85]), .CK(clk), .Q(reg_in[85]) );
  DFF_X1 \reg_in_reg[84]  ( .D(Plaintext[84]), .CK(clk), .Q(reg_in[84]) );
  DFF_X1 \reg_in_reg[83]  ( .D(Plaintext[83]), .CK(clk), .Q(reg_in[83]) );
  DFF_X1 \reg_in_reg[82]  ( .D(Plaintext[82]), .CK(clk), .Q(reg_in[82]) );
  DFF_X1 \reg_in_reg[81]  ( .D(Plaintext[81]), .CK(clk), .Q(reg_in[81]) );
  DFF_X1 \reg_in_reg[80]  ( .D(Plaintext[80]), .CK(clk), .Q(reg_in[80]) );
  DFF_X1 \reg_in_reg[79]  ( .D(Plaintext[79]), .CK(clk), .Q(reg_in[79]) );
  DFF_X1 \reg_in_reg[78]  ( .D(Plaintext[78]), .CK(clk), .Q(reg_in[78]) );
  DFF_X1 \reg_in_reg[77]  ( .D(Plaintext[77]), .CK(clk), .Q(reg_in[77]) );
  DFF_X1 \reg_in_reg[76]  ( .D(Plaintext[76]), .CK(clk), .Q(reg_in[76]) );
  DFF_X1 \reg_in_reg[75]  ( .D(Plaintext[75]), .CK(clk), .Q(reg_in[75]) );
  DFF_X1 \reg_in_reg[74]  ( .D(Plaintext[74]), .CK(clk), .Q(reg_in[74]) );
  DFF_X1 \reg_in_reg[73]  ( .D(Plaintext[73]), .CK(clk), .Q(reg_in[73]) );
  DFF_X1 \reg_in_reg[72]  ( .D(Plaintext[72]), .CK(clk), .Q(reg_in[72]) );
  DFF_X1 \reg_in_reg[71]  ( .D(Plaintext[71]), .CK(clk), .Q(reg_in[71]) );
  DFF_X1 \reg_in_reg[70]  ( .D(Plaintext[70]), .CK(clk), .Q(reg_in[70]) );
  DFF_X1 \reg_in_reg[69]  ( .D(Plaintext[69]), .CK(clk), .Q(reg_in[69]) );
  DFF_X1 \reg_in_reg[68]  ( .D(Plaintext[68]), .CK(clk), .Q(reg_in[68]) );
  DFF_X1 \reg_in_reg[67]  ( .D(Plaintext[67]), .CK(clk), .Q(reg_in[67]) );
  DFF_X1 \reg_in_reg[66]  ( .D(Plaintext[66]), .CK(clk), .Q(reg_in[66]) );
  DFF_X1 \reg_in_reg[65]  ( .D(Plaintext[65]), .CK(clk), .Q(reg_in[65]) );
  DFF_X1 \reg_in_reg[64]  ( .D(Plaintext[64]), .CK(clk), .Q(reg_in[64]) );
  DFF_X1 \reg_in_reg[63]  ( .D(Plaintext[63]), .CK(clk), .Q(reg_in[63]) );
  DFF_X1 \reg_in_reg[62]  ( .D(Plaintext[62]), .CK(clk), .Q(reg_in[62]) );
  DFF_X1 \reg_in_reg[61]  ( .D(Plaintext[61]), .CK(clk), .Q(reg_in[61]) );
  DFF_X1 \reg_in_reg[60]  ( .D(Plaintext[60]), .CK(clk), .Q(reg_in[60]) );
  DFF_X1 \reg_in_reg[59]  ( .D(Plaintext[59]), .CK(clk), .Q(reg_in[59]) );
  DFF_X1 \reg_in_reg[58]  ( .D(Plaintext[58]), .CK(clk), .Q(reg_in[58]) );
  DFF_X1 \reg_in_reg[57]  ( .D(Plaintext[57]), .CK(clk), .Q(reg_in[57]) );
  DFF_X1 \reg_in_reg[56]  ( .D(Plaintext[56]), .CK(clk), .Q(reg_in[56]) );
  DFF_X1 \reg_in_reg[55]  ( .D(Plaintext[55]), .CK(clk), .Q(reg_in[55]) );
  DFF_X1 \reg_in_reg[54]  ( .D(Plaintext[54]), .CK(clk), .Q(reg_in[54]) );
  DFF_X1 \reg_in_reg[53]  ( .D(Plaintext[53]), .CK(clk), .Q(reg_in[53]) );
  DFF_X1 \reg_in_reg[52]  ( .D(Plaintext[52]), .CK(clk), .Q(reg_in[52]) );
  DFF_X1 \reg_in_reg[51]  ( .D(Plaintext[51]), .CK(clk), .Q(reg_in[51]) );
  DFF_X1 \reg_in_reg[50]  ( .D(Plaintext[50]), .CK(clk), .Q(reg_in[50]) );
  DFF_X1 \reg_in_reg[49]  ( .D(Plaintext[49]), .CK(clk), .Q(reg_in[49]) );
  DFF_X1 \reg_in_reg[48]  ( .D(Plaintext[48]), .CK(clk), .Q(reg_in[48]) );
  DFF_X1 \reg_in_reg[47]  ( .D(Plaintext[47]), .CK(clk), .Q(reg_in[47]) );
  DFF_X1 \reg_in_reg[46]  ( .D(Plaintext[46]), .CK(clk), .Q(reg_in[46]) );
  DFF_X1 \reg_in_reg[45]  ( .D(Plaintext[45]), .CK(clk), .Q(reg_in[45]) );
  DFF_X1 \reg_in_reg[44]  ( .D(Plaintext[44]), .CK(clk), .Q(reg_in[44]) );
  DFF_X1 \reg_in_reg[43]  ( .D(Plaintext[43]), .CK(clk), .Q(reg_in[43]) );
  DFF_X1 \reg_in_reg[42]  ( .D(Plaintext[42]), .CK(clk), .Q(reg_in[42]) );
  DFF_X1 \reg_in_reg[41]  ( .D(Plaintext[41]), .CK(clk), .Q(reg_in[41]) );
  DFF_X1 \reg_in_reg[40]  ( .D(Plaintext[40]), .CK(clk), .Q(reg_in[40]) );
  DFF_X1 \reg_in_reg[39]  ( .D(Plaintext[39]), .CK(clk), .Q(reg_in[39]) );
  DFF_X1 \reg_in_reg[38]  ( .D(Plaintext[38]), .CK(clk), .Q(reg_in[38]) );
  DFF_X1 \reg_in_reg[37]  ( .D(Plaintext[37]), .CK(clk), .Q(reg_in[37]) );
  DFF_X1 \reg_in_reg[36]  ( .D(Plaintext[36]), .CK(clk), .Q(reg_in[36]) );
  DFF_X1 \reg_in_reg[35]  ( .D(Plaintext[35]), .CK(clk), .Q(reg_in[35]) );
  DFF_X1 \reg_in_reg[34]  ( .D(Plaintext[34]), .CK(clk), .Q(reg_in[34]) );
  DFF_X1 \reg_in_reg[33]  ( .D(Plaintext[33]), .CK(clk), .Q(reg_in[33]) );
  DFF_X1 \reg_in_reg[32]  ( .D(Plaintext[32]), .CK(clk), .Q(reg_in[32]) );
  DFF_X1 \reg_in_reg[31]  ( .D(Plaintext[31]), .CK(clk), .Q(reg_in[31]) );
  DFF_X1 \reg_in_reg[30]  ( .D(Plaintext[30]), .CK(clk), .Q(reg_in[30]) );
  DFF_X1 \reg_in_reg[29]  ( .D(Plaintext[29]), .CK(clk), .Q(reg_in[29]) );
  DFF_X1 \reg_in_reg[28]  ( .D(Plaintext[28]), .CK(clk), .Q(reg_in[28]) );
  DFF_X1 \reg_in_reg[27]  ( .D(Plaintext[27]), .CK(clk), .Q(reg_in[27]) );
  DFF_X1 \reg_in_reg[26]  ( .D(Plaintext[26]), .CK(clk), .Q(reg_in[26]) );
  DFF_X1 \reg_in_reg[25]  ( .D(Plaintext[25]), .CK(clk), .Q(reg_in[25]) );
  DFF_X1 \reg_in_reg[24]  ( .D(Plaintext[24]), .CK(clk), .Q(reg_in[24]) );
  DFF_X1 \reg_in_reg[23]  ( .D(Plaintext[23]), .CK(clk), .Q(reg_in[23]) );
  DFF_X1 \reg_in_reg[22]  ( .D(Plaintext[22]), .CK(clk), .Q(reg_in[22]) );
  DFF_X1 \reg_in_reg[21]  ( .D(Plaintext[21]), .CK(clk), .Q(reg_in[21]) );
  DFF_X1 \reg_in_reg[20]  ( .D(Plaintext[20]), .CK(clk), .Q(reg_in[20]) );
  DFF_X1 \reg_in_reg[19]  ( .D(Plaintext[19]), .CK(clk), .Q(reg_in[19]) );
  DFF_X1 \reg_in_reg[18]  ( .D(Plaintext[18]), .CK(clk), .Q(reg_in[18]) );
  DFF_X1 \reg_in_reg[17]  ( .D(Plaintext[17]), .CK(clk), .Q(reg_in[17]) );
  DFF_X1 \reg_in_reg[16]  ( .D(Plaintext[16]), .CK(clk), .Q(reg_in[16]) );
  DFF_X1 \reg_in_reg[15]  ( .D(Plaintext[15]), .CK(clk), .Q(reg_in[15]) );
  DFF_X1 \reg_in_reg[14]  ( .D(Plaintext[14]), .CK(clk), .Q(reg_in[14]) );
  DFF_X1 \reg_in_reg[13]  ( .D(Plaintext[13]), .CK(clk), .Q(reg_in[13]) );
  DFF_X1 \reg_in_reg[12]  ( .D(Plaintext[12]), .CK(clk), .Q(reg_in[12]) );
  DFF_X1 \reg_in_reg[11]  ( .D(Plaintext[11]), .CK(clk), .Q(reg_in[11]) );
  DFF_X1 \reg_in_reg[10]  ( .D(Plaintext[10]), .CK(clk), .Q(reg_in[10]) );
  DFF_X1 \reg_in_reg[9]  ( .D(Plaintext[9]), .CK(clk), .Q(reg_in[9]) );
  DFF_X1 \reg_in_reg[8]  ( .D(Plaintext[8]), .CK(clk), .Q(reg_in[8]) );
  DFF_X1 \reg_in_reg[7]  ( .D(Plaintext[7]), .CK(clk), .Q(reg_in[7]) );
  DFF_X1 \reg_in_reg[6]  ( .D(Plaintext[6]), .CK(clk), .Q(reg_in[6]) );
  DFF_X1 \reg_in_reg[5]  ( .D(Plaintext[5]), .CK(clk), .Q(reg_in[5]) );
  DFF_X1 \reg_in_reg[4]  ( .D(Plaintext[4]), .CK(clk), .Q(reg_in[4]) );
  DFF_X1 \reg_in_reg[3]  ( .D(Plaintext[3]), .CK(clk), .Q(reg_in[3]) );
  DFF_X1 \reg_in_reg[2]  ( .D(Plaintext[2]), .CK(clk), .Q(reg_in[2]) );
  DFF_X1 \reg_in_reg[1]  ( .D(Plaintext[1]), .CK(clk), .Q(reg_in[1]) );
  DFF_X1 \reg_in_reg[0]  ( .D(Plaintext[0]), .CK(clk), .Q(reg_in[0]) );
  DFF_X1 \reg_key_reg[191]  ( .D(Key[191]), .CK(clk), .Q(reg_key[191]) );
  DFF_X1 \reg_key_reg[190]  ( .D(Key[190]), .CK(clk), .Q(reg_key[190]) );
  DFF_X1 \reg_key_reg[189]  ( .D(Key[189]), .CK(clk), .Q(reg_key[189]) );
  DFF_X1 \reg_key_reg[188]  ( .D(Key[188]), .CK(clk), .Q(reg_key[188]) );
  DFF_X1 \reg_key_reg[187]  ( .D(Key[187]), .CK(clk), .Q(reg_key[187]) );
  DFF_X1 \reg_key_reg[184]  ( .D(Key[184]), .CK(clk), .Q(reg_key[184]) );
  DFF_X1 \reg_key_reg[179]  ( .D(Key[179]), .CK(clk), .Q(reg_key[179]) );
  DFF_X1 \reg_key_reg[178]  ( .D(Key[178]), .CK(clk), .Q(reg_key[178]) );
  DFF_X1 \reg_key_reg[177]  ( .D(Key[177]), .CK(clk), .Q(reg_key[177]) );
  DFF_X1 \reg_key_reg[173]  ( .D(Key[173]), .CK(clk), .Q(reg_key[173]) );
  DFF_X1 \reg_key_reg[171]  ( .D(Key[171]), .CK(clk), .Q(reg_key[171]) );
  DFF_X1 \reg_key_reg[169]  ( .D(Key[169]), .CK(clk), .Q(reg_key[169]) );
  DFF_X1 \reg_key_reg[165]  ( .D(Key[165]), .CK(clk), .Q(reg_key[165]) );
  DFF_X1 \reg_key_reg[160]  ( .D(Key[160]), .CK(clk), .Q(reg_key[160]) );
  DFF_X1 \reg_key_reg[156]  ( .D(Key[156]), .CK(clk), .Q(reg_key[156]) );
  DFF_X1 \reg_key_reg[151]  ( .D(Key[151]), .CK(clk), .Q(reg_key[151]) );
  DFF_X1 \reg_key_reg[149]  ( .D(Key[149]), .CK(clk), .Q(reg_key[149]) );
  DFF_X1 \reg_key_reg[143]  ( .D(Key[143]), .CK(clk), .Q(reg_key[143]) );
  DFF_X1 \reg_key_reg[140]  ( .D(Key[140]), .CK(clk), .Q(reg_key[140]) );
  DFF_X1 \reg_key_reg[137]  ( .D(Key[137]), .CK(clk), .Q(reg_key[137]) );
  DFF_X1 \reg_key_reg[135]  ( .D(Key[135]), .CK(clk), .Q(reg_key[135]) );
  DFF_X1 \reg_key_reg[132]  ( .D(Key[132]), .CK(clk), .Q(reg_key[132]) );
  DFF_X1 \reg_key_reg[125]  ( .D(Key[125]), .CK(clk), .Q(reg_key[125]) );
  DFF_X1 \reg_key_reg[123]  ( .D(Key[123]), .CK(clk), .Q(reg_key[123]) );
  DFF_X1 \reg_key_reg[120]  ( .D(Key[120]), .CK(clk), .Q(reg_key[120]) );
  DFF_X1 \reg_key_reg[119]  ( .D(Key[119]), .CK(clk), .Q(reg_key[119]) );
  DFF_X1 \reg_key_reg[118]  ( .D(Key[118]), .CK(clk), .Q(reg_key[118]) );
  DFF_X1 \reg_key_reg[109]  ( .D(Key[109]), .CK(clk), .Q(reg_key[109]) );
  DFF_X1 \reg_key_reg[108]  ( .D(Key[108]), .CK(clk), .Q(reg_key[108]) );
  DFF_X1 \reg_key_reg[105]  ( .D(Key[105]), .CK(clk), .Q(reg_key[105]) );
  DFF_X1 \reg_key_reg[104]  ( .D(Key[104]), .CK(clk), .Q(reg_key[104]) );
  DFF_X1 \reg_key_reg[103]  ( .D(Key[103]), .CK(clk), .Q(reg_key[103]) );
  DFF_X1 \reg_key_reg[101]  ( .D(Key[101]), .CK(clk), .Q(reg_key[101]) );
  DFF_X1 \reg_key_reg[100]  ( .D(Key[100]), .CK(clk), .Q(reg_key[100]) );
  DFF_X1 \reg_key_reg[96]  ( .D(Key[96]), .CK(clk), .Q(reg_key[96]) );
  DFF_X1 \reg_key_reg[95]  ( .D(Key[95]), .CK(clk), .Q(reg_key[95]) );
  DFF_X1 \reg_key_reg[82]  ( .D(Key[82]), .CK(clk), .Q(reg_key[82]) );
  DFF_X1 \reg_key_reg[81]  ( .D(Key[81]), .CK(clk), .Q(reg_key[81]) );
  DFF_X1 \reg_key_reg[80]  ( .D(Key[80]), .CK(clk), .Q(reg_key[80]) );
  DFF_X1 \reg_key_reg[76]  ( .D(Key[76]), .CK(clk), .Q(reg_key[76]) );
  DFF_X1 \reg_key_reg[71]  ( .D(Key[71]), .CK(clk), .Q(reg_key[71]) );
  DFF_X1 \reg_key_reg[66]  ( .D(Key[66]), .CK(clk), .Q(reg_key[66]) );
  DFF_X1 \reg_key_reg[65]  ( .D(Key[65]), .CK(clk), .Q(reg_key[65]) );
  DFF_X1 \reg_key_reg[60]  ( .D(Key[60]), .CK(clk), .Q(reg_key[60]) );
  DFF_X1 \reg_key_reg[59]  ( .D(Key[59]), .CK(clk), .Q(reg_key[59]) );
  DFF_X1 \reg_key_reg[58]  ( .D(Key[58]), .CK(clk), .Q(reg_key[58]) );
  DFF_X1 \reg_key_reg[51]  ( .D(Key[51]), .CK(clk), .Q(reg_key[51]) );
  DFF_X1 \reg_key_reg[48]  ( .D(Key[48]), .CK(clk), .Q(reg_key[48]) );
  DFF_X1 \reg_key_reg[45]  ( .D(Key[45]), .CK(clk), .Q(reg_key[45]) );
  DFF_X1 \reg_key_reg[44]  ( .D(Key[44]), .CK(clk), .Q(reg_key[44]) );
  DFF_X1 \reg_key_reg[38]  ( .D(Key[38]), .CK(clk), .Q(reg_key[38]) );
  DFF_X1 \reg_key_reg[36]  ( .D(Key[36]), .CK(clk), .Q(reg_key[36]) );
  DFF_X1 \reg_key_reg[30]  ( .D(Key[30]), .CK(clk), .Q(reg_key[30]) );
  DFF_X1 \reg_key_reg[28]  ( .D(Key[28]), .CK(clk), .Q(reg_key[28]) );
  DFF_X1 \reg_key_reg[25]  ( .D(Key[25]), .CK(clk), .Q(reg_key[25]) );
  DFF_X1 \reg_key_reg[24]  ( .D(Key[24]), .CK(clk), .Q(reg_key[24]) );
  DFF_X1 \reg_key_reg[21]  ( .D(Key[21]), .CK(clk), .Q(reg_key[21]) );
  DFF_X1 \reg_key_reg[20]  ( .D(Key[20]), .CK(clk), .Q(reg_key[20]) );
  DFF_X1 \reg_key_reg[18]  ( .D(Key[18]), .CK(clk), .Q(reg_key[18]) );
  DFF_X1 \reg_key_reg[10]  ( .D(Key[10]), .CK(clk), .Q(reg_key[10]) );
  DFF_X1 \reg_key_reg[9]  ( .D(Key[9]), .CK(clk), .Q(reg_key[9]) );
  DFF_X1 \reg_key_reg[6]  ( .D(Key[6]), .CK(clk), .Q(reg_key[6]) );
  DFF_X1 \reg_key_reg[5]  ( .D(Key[5]), .CK(clk), .Q(reg_key[5]) );
  DFF_X1 \reg_key_reg[4]  ( .D(Key[4]), .CK(clk), .Q(reg_key[4]) );
  DFF_X1 \reg_key_reg[3]  ( .D(Key[3]), .CK(clk), .Q(reg_key[3]) );
  DFF_X1 \Ciphertext_reg[190]  ( .D(reg_out[190]), .CK(clk), .Q(
        Ciphertext[190]) );
  DFF_X1 \Ciphertext_reg[188]  ( .D(reg_out[188]), .CK(clk), .Q(
        Ciphertext[188]) );
  DFF_X1 \Ciphertext_reg[187]  ( .D(reg_out[187]), .CK(clk), .Q(
        Ciphertext[187]) );
  DFF_X1 \Ciphertext_reg[185]  ( .D(reg_out[185]), .CK(clk), .Q(
        Ciphertext[185]) );
  DFF_X1 \Ciphertext_reg[183]  ( .D(reg_out[183]), .CK(clk), .Q(
        Ciphertext[183]) );
  DFF_X1 \Ciphertext_reg[177]  ( .D(reg_out[177]), .CK(clk), .Q(
        Ciphertext[177]) );
  DFF_X1 \Ciphertext_reg[171]  ( .D(reg_out[171]), .CK(clk), .Q(
        Ciphertext[171]) );
  DFF_X1 \Ciphertext_reg[170]  ( .D(reg_out[170]), .CK(clk), .Q(
        Ciphertext[170]) );
  DFF_X1 \Ciphertext_reg[169]  ( .D(reg_out[169]), .CK(clk), .Q(
        Ciphertext[169]) );
  DFF_X1 \Ciphertext_reg[168]  ( .D(reg_out[168]), .CK(clk), .Q(
        Ciphertext[168]) );
  DFF_X1 \Ciphertext_reg[167]  ( .D(reg_out[167]), .CK(clk), .Q(
        Ciphertext[167]) );
  DFF_X1 \Ciphertext_reg[165]  ( .D(reg_out[165]), .CK(clk), .Q(
        Ciphertext[165]) );
  DFF_X1 \Ciphertext_reg[164]  ( .D(reg_out[164]), .CK(clk), .Q(
        Ciphertext[164]) );
  DFF_X1 \Ciphertext_reg[163]  ( .D(reg_out[163]), .CK(clk), .Q(
        Ciphertext[163]) );
  DFF_X1 \Ciphertext_reg[160]  ( .D(reg_out[160]), .CK(clk), .Q(
        Ciphertext[160]) );
  DFF_X1 \Ciphertext_reg[159]  ( .D(reg_out[159]), .CK(clk), .Q(
        Ciphertext[159]) );
  DFF_X1 \Ciphertext_reg[158]  ( .D(reg_out[158]), .CK(clk), .Q(
        Ciphertext[158]) );
  DFF_X1 \Ciphertext_reg[155]  ( .D(reg_out[155]), .CK(clk), .Q(
        Ciphertext[155]) );
  DFF_X1 \Ciphertext_reg[152]  ( .D(reg_out[152]), .CK(clk), .Q(
        Ciphertext[152]) );
  DFF_X1 \Ciphertext_reg[149]  ( .D(reg_out[149]), .CK(clk), .Q(
        Ciphertext[149]) );
  DFF_X1 \Ciphertext_reg[148]  ( .D(reg_out[148]), .CK(clk), .Q(
        Ciphertext[148]) );
  DFF_X1 \Ciphertext_reg[147]  ( .D(reg_out[147]), .CK(clk), .Q(
        Ciphertext[147]) );
  DFF_X1 \Ciphertext_reg[145]  ( .D(reg_out[145]), .CK(clk), .Q(
        Ciphertext[145]) );
  DFF_X1 \Ciphertext_reg[143]  ( .D(reg_out[143]), .CK(clk), .Q(
        Ciphertext[143]) );
  DFF_X1 \Ciphertext_reg[142]  ( .D(reg_out[142]), .CK(clk), .Q(
        Ciphertext[142]) );
  DFF_X1 \Ciphertext_reg[141]  ( .D(reg_out[141]), .CK(clk), .Q(
        Ciphertext[141]) );
  DFF_X1 \Ciphertext_reg[140]  ( .D(reg_out[140]), .CK(clk), .Q(
        Ciphertext[140]) );
  DFF_X1 \Ciphertext_reg[139]  ( .D(reg_out[139]), .CK(clk), .Q(
        Ciphertext[139]) );
  DFF_X1 \Ciphertext_reg[138]  ( .D(reg_out[138]), .CK(clk), .Q(
        Ciphertext[138]) );
  DFF_X1 \Ciphertext_reg[137]  ( .D(reg_out[137]), .CK(clk), .Q(
        Ciphertext[137]) );
  DFF_X1 \Ciphertext_reg[136]  ( .D(reg_out[136]), .CK(clk), .Q(
        Ciphertext[136]) );
  DFF_X1 \Ciphertext_reg[135]  ( .D(reg_out[135]), .CK(clk), .Q(
        Ciphertext[135]) );
  DFF_X1 \Ciphertext_reg[131]  ( .D(reg_out[131]), .CK(clk), .Q(
        Ciphertext[131]) );
  DFF_X1 \Ciphertext_reg[130]  ( .D(reg_out[130]), .CK(clk), .Q(
        Ciphertext[130]) );
  DFF_X1 \Ciphertext_reg[129]  ( .D(reg_out[129]), .CK(clk), .Q(
        Ciphertext[129]) );
  DFF_X1 \Ciphertext_reg[128]  ( .D(reg_out[128]), .CK(clk), .Q(
        Ciphertext[128]) );
  DFF_X1 \Ciphertext_reg[126]  ( .D(reg_out[126]), .CK(clk), .Q(
        Ciphertext[126]) );
  DFF_X1 \Ciphertext_reg[125]  ( .D(reg_out[125]), .CK(clk), .Q(
        Ciphertext[125]) );
  DFF_X1 \Ciphertext_reg[122]  ( .D(reg_out[122]), .CK(clk), .Q(
        Ciphertext[122]) );
  DFF_X1 \Ciphertext_reg[120]  ( .D(reg_out[120]), .CK(clk), .Q(
        Ciphertext[120]) );
  DFF_X1 \Ciphertext_reg[118]  ( .D(reg_out[118]), .CK(clk), .Q(
        Ciphertext[118]) );
  DFF_X1 \Ciphertext_reg[116]  ( .D(reg_out[116]), .CK(clk), .Q(
        Ciphertext[116]) );
  DFF_X1 \Ciphertext_reg[112]  ( .D(reg_out[112]), .CK(clk), .Q(
        Ciphertext[112]) );
  DFF_X1 \Ciphertext_reg[108]  ( .D(reg_out[108]), .CK(clk), .Q(
        Ciphertext[108]) );
  DFF_X1 \Ciphertext_reg[106]  ( .D(reg_out[106]), .CK(clk), .Q(
        Ciphertext[106]) );
  DFF_X1 \Ciphertext_reg[101]  ( .D(reg_out[101]), .CK(clk), .Q(
        Ciphertext[101]) );
  DFF_X1 \Ciphertext_reg[98]  ( .D(reg_out[98]), .CK(clk), .Q(Ciphertext[98])
         );
  DFF_X1 \Ciphertext_reg[92]  ( .D(reg_out[92]), .CK(clk), .Q(Ciphertext[92])
         );
  DFF_X1 \Ciphertext_reg[91]  ( .D(reg_out[91]), .CK(clk), .Q(Ciphertext[91])
         );
  DFF_X1 \Ciphertext_reg[89]  ( .D(reg_out[89]), .CK(clk), .Q(Ciphertext[89])
         );
  DFF_X1 \Ciphertext_reg[88]  ( .D(reg_out[88]), .CK(clk), .Q(Ciphertext[88])
         );
  DFF_X1 \Ciphertext_reg[87]  ( .D(reg_out[87]), .CK(clk), .Q(Ciphertext[87])
         );
  DFF_X1 \Ciphertext_reg[86]  ( .D(reg_out[86]), .CK(clk), .Q(Ciphertext[86])
         );
  DFF_X1 \Ciphertext_reg[84]  ( .D(reg_out[84]), .CK(clk), .Q(Ciphertext[84])
         );
  DFF_X1 \Ciphertext_reg[83]  ( .D(reg_out[83]), .CK(clk), .Q(Ciphertext[83])
         );
  DFF_X1 \Ciphertext_reg[82]  ( .D(reg_out[82]), .CK(clk), .Q(Ciphertext[82])
         );
  DFF_X1 \Ciphertext_reg[77]  ( .D(reg_out[77]), .CK(clk), .Q(Ciphertext[77])
         );
  DFF_X1 \Ciphertext_reg[74]  ( .D(reg_out[74]), .CK(clk), .Q(Ciphertext[74])
         );
  DFF_X1 \Ciphertext_reg[72]  ( .D(reg_out[72]), .CK(clk), .Q(Ciphertext[72])
         );
  DFF_X1 \Ciphertext_reg[64]  ( .D(reg_out[64]), .CK(clk), .Q(Ciphertext[64])
         );
  DFF_X1 \Ciphertext_reg[62]  ( .D(reg_out[62]), .CK(clk), .Q(Ciphertext[62])
         );
  DFF_X1 \Ciphertext_reg[57]  ( .D(reg_out[57]), .CK(clk), .Q(Ciphertext[57])
         );
  DFF_X1 \Ciphertext_reg[56]  ( .D(reg_out[56]), .CK(clk), .Q(Ciphertext[56])
         );
  DFF_X1 \Ciphertext_reg[54]  ( .D(reg_out[54]), .CK(clk), .Q(Ciphertext[54])
         );
  DFF_X1 \Ciphertext_reg[49]  ( .D(reg_out[49]), .CK(clk), .Q(Ciphertext[49])
         );
  DFF_X1 \Ciphertext_reg[46]  ( .D(reg_out[46]), .CK(clk), .Q(Ciphertext[46])
         );
  DFF_X1 \Ciphertext_reg[41]  ( .D(reg_out[41]), .CK(clk), .Q(Ciphertext[41])
         );
  DFF_X1 \Ciphertext_reg[37]  ( .D(reg_out[37]), .CK(clk), .Q(Ciphertext[37])
         );
  DFF_X1 \Ciphertext_reg[35]  ( .D(reg_out[35]), .CK(clk), .Q(Ciphertext[35])
         );
  DFF_X1 \Ciphertext_reg[34]  ( .D(reg_out[34]), .CK(clk), .Q(Ciphertext[34])
         );
  DFF_X1 \Ciphertext_reg[33]  ( .D(reg_out[33]), .CK(clk), .Q(Ciphertext[33])
         );
  DFF_X1 \Ciphertext_reg[32]  ( .D(reg_out[32]), .CK(clk), .Q(Ciphertext[32])
         );
  DFF_X1 \Ciphertext_reg[31]  ( .D(reg_out[31]), .CK(clk), .Q(Ciphertext[31])
         );
  DFF_X1 \Ciphertext_reg[30]  ( .D(reg_out[30]), .CK(clk), .Q(Ciphertext[30])
         );
  DFF_X1 \Ciphertext_reg[29]  ( .D(reg_out[29]), .CK(clk), .Q(Ciphertext[29])
         );
  DFF_X1 \Ciphertext_reg[28]  ( .D(reg_out[28]), .CK(clk), .Q(Ciphertext[28])
         );
  DFF_X1 \Ciphertext_reg[26]  ( .D(reg_out[26]), .CK(clk), .Q(Ciphertext[26])
         );
  DFF_X1 \Ciphertext_reg[23]  ( .D(reg_out[23]), .CK(clk), .Q(Ciphertext[23])
         );
  DFF_X1 \Ciphertext_reg[18]  ( .D(reg_out[18]), .CK(clk), .Q(Ciphertext[18])
         );
  DFF_X1 \Ciphertext_reg[17]  ( .D(reg_out[17]), .CK(clk), .Q(Ciphertext[17])
         );
  DFF_X1 \Ciphertext_reg[15]  ( .D(reg_out[15]), .CK(clk), .Q(Ciphertext[15])
         );
  DFF_X1 \Ciphertext_reg[14]  ( .D(reg_out[14]), .CK(clk), .Q(Ciphertext[14])
         );
  DFF_X1 \Ciphertext_reg[13]  ( .D(reg_out[13]), .CK(clk), .Q(Ciphertext[13])
         );
  DFF_X1 \Ciphertext_reg[11]  ( .D(reg_out[11]), .CK(clk), .Q(Ciphertext[11])
         );
  DFF_X1 \Ciphertext_reg[10]  ( .D(reg_out[10]), .CK(clk), .Q(Ciphertext[10])
         );
  DFF_X1 \Ciphertext_reg[8]  ( .D(reg_out[8]), .CK(clk), .Q(Ciphertext[8]) );
  DFF_X1 \Ciphertext_reg[6]  ( .D(reg_out[6]), .CK(clk), .Q(Ciphertext[6]) );
  DFF_X1 \Ciphertext_reg[5]  ( .D(reg_out[5]), .CK(clk), .Q(Ciphertext[5]) );
  DFF_X1 \Ciphertext_reg[4]  ( .D(reg_out[4]), .CK(clk), .Q(Ciphertext[4]) );
  DFF_X1 \Ciphertext_reg[2]  ( .D(reg_out[2]), .CK(clk), .Q(Ciphertext[2]) );
  DFF_X1 \Ciphertext_reg[0]  ( .D(reg_out[0]), .CK(clk), .Q(Ciphertext[0]) );
  DFF_X1 \reg_key_reg[14]  ( .D(Key[14]), .CK(clk), .Q(reg_key[14]) );
  DFF_X1 \reg_key_reg[122]  ( .D(Key[122]), .CK(clk), .Q(reg_key[122]) );
  DFF_X1 \reg_key_reg[86]  ( .D(Key[86]), .CK(clk), .Q(reg_key[86]) );
  DFF_X1 \Ciphertext_reg[100]  ( .D(reg_out[100]), .CK(clk), .Q(
        Ciphertext[100]) );
  DFF_X1 \reg_key_reg[111]  ( .D(Key[111]), .CK(clk), .Q(reg_key[111]) );
  DFF_X1 \reg_key_reg[54]  ( .D(Key[54]), .CK(clk), .Q(reg_key[54]) );
  DFF_X1 \reg_key_reg[61]  ( .D(Key[61]), .CK(clk), .Q(reg_key[61]) );
  DFF_X1 \reg_key_reg[116]  ( .D(Key[116]), .CK(clk), .Q(reg_key[116]) );
  DFF_X1 \reg_key_reg[158]  ( .D(Key[158]), .CK(clk), .Q(reg_key[158]) );
  DFF_X1 \reg_key_reg[15]  ( .D(Key[15]), .CK(clk), .Q(reg_key[15]) );
  DFF_X1 \reg_key_reg[185]  ( .D(Key[185]), .CK(clk), .Q(reg_key[185]) );
  DFF_X1 \reg_key_reg[13]  ( .D(Key[13]), .CK(clk), .Q(reg_key[13]) );
  DFF_X1 \reg_key_reg[8]  ( .D(Key[8]), .CK(clk), .Q(reg_key[8]) );
  DFF_X1 \reg_key_reg[2]  ( .D(Key[2]), .CK(clk), .Q(reg_key[2]) );
  DFF_X1 \reg_key_reg[29]  ( .D(Key[29]), .CK(clk), .Q(reg_key[29]) );
  DFF_X1 \reg_key_reg[74]  ( .D(Key[74]), .CK(clk), .Q(reg_key[74]) );
  DFF_X1 \reg_key_reg[98]  ( .D(Key[98]), .CK(clk), .Q(reg_key[98]) );
  DFF_X1 \reg_key_reg[83]  ( .D(Key[83]), .CK(clk), .Q(reg_key[83]) );
  DFF_X1 \reg_key_reg[183]  ( .D(Key[183]), .CK(clk), .Q(reg_key[183]) );
  DFF_X1 \reg_key_reg[107]  ( .D(Key[107]), .CK(clk), .Q(reg_key[107]) );
  DFF_X1 \reg_key_reg[146]  ( .D(Key[146]), .CK(clk), .Q(reg_key[146]) );
  DFF_X1 \reg_key_reg[56]  ( .D(Key[56]), .CK(clk), .Q(reg_key[56]) );
  DFF_X1 \reg_key_reg[152]  ( .D(Key[152]), .CK(clk), .Q(reg_key[152]) );
  DFF_X1 \reg_key_reg[63]  ( .D(Key[63]), .CK(clk), .Q(reg_key[63]) );
  DFF_X1 \reg_key_reg[134]  ( .D(Key[134]), .CK(clk), .Q(reg_key[134]) );
  DFF_X1 \reg_key_reg[106]  ( .D(Key[106]), .CK(clk), .Q(reg_key[106]) );
  DFF_X1 \reg_key_reg[41]  ( .D(Key[41]), .CK(clk), .Q(reg_key[41]) );
  DFF_X1 \reg_key_reg[16]  ( .D(Key[16]), .CK(clk), .Q(reg_key[16]) );
  DFF_X1 \reg_key_reg[35]  ( .D(Key[35]), .CK(clk), .Q(reg_key[35]) );
  DFF_X1 \reg_key_reg[102]  ( .D(Key[102]), .CK(clk), .Q(reg_key[102]) );
  DFF_X1 \reg_key_reg[27]  ( .D(Key[27]), .CK(clk), .Q(reg_key[27]) );
  DFF_X1 \Ciphertext_reg[124]  ( .D(reg_out[124]), .CK(clk), .Q(
        Ciphertext[124]) );
  DFF_X1 \reg_key_reg[22]  ( .D(Key[22]), .CK(clk), .Q(reg_key[22]) );
  DFF_X1 \reg_key_reg[163]  ( .D(Key[163]), .CK(clk), .Q(reg_key[163]) );
  DFF_X1 \reg_key_reg[159]  ( .D(Key[159]), .CK(clk), .Q(reg_key[159]) );
  DFF_X1 \reg_key_reg[155]  ( .D(Key[155]), .CK(clk), .Q(reg_key[155]) );
  DFF_X1 \reg_key_reg[147]  ( .D(Key[147]), .CK(clk), .Q(reg_key[147]) );
  DFF_X1 \reg_key_reg[49]  ( .D(Key[49]), .CK(clk), .Q(reg_key[49]) );
  DFF_X1 \reg_key_reg[92]  ( .D(Key[92]), .CK(clk), .Q(reg_key[92]) );
  DFF_X1 \reg_key_reg[186]  ( .D(Key[186]), .CK(clk), .Q(reg_key[186]) );
  DFF_X1 \reg_key_reg[182]  ( .D(Key[182]), .CK(clk), .Q(reg_key[182]) );
  DFF_X1 \reg_key_reg[84]  ( .D(Key[84]), .CK(clk), .Q(reg_key[84]) );
  DFF_X1 \reg_key_reg[131]  ( .D(Key[131]), .CK(clk), .Q(reg_key[131]) );
  DFF_X1 \reg_key_reg[170]  ( .D(Key[170]), .CK(clk), .Q(reg_key[170]) );
  DFF_X1 \reg_key_reg[72]  ( .D(Key[72]), .CK(clk), .Q(reg_key[72]) );
  DFF_X1 \reg_key_reg[68]  ( .D(Key[68]), .CK(clk), .Q(reg_key[68]) );
  DFF_X1 \reg_key_reg[17]  ( .D(Key[17]), .CK(clk), .Q(reg_key[17]) );
  DFF_X1 \reg_key_reg[154]  ( .D(Key[154]), .CK(clk), .Q(reg_key[154]) );
  DFF_X1 \reg_key_reg[150]  ( .D(Key[150]), .CK(clk), .Q(reg_key[150]) );
  DFF_X1 \reg_key_reg[99]  ( .D(Key[99]), .CK(clk), .Q(reg_key[99]) );
  DFF_X1 \reg_key_reg[1]  ( .D(Key[1]), .CK(clk), .Q(reg_key[1]) );
  DFF_X1 \reg_key_reg[138]  ( .D(Key[138]), .CK(clk), .Q(reg_key[138]) );
  DFF_X1 \reg_key_reg[40]  ( .D(Key[40]), .CK(clk), .Q(reg_key[40]) );
  DFF_X1 \reg_key_reg[87]  ( .D(Key[87]), .CK(clk), .Q(reg_key[87]) );
  DFF_X1 \reg_key_reg[181]  ( .D(Key[181]), .CK(clk), .Q(reg_key[181]) );
  DFF_X1 \reg_key_reg[130]  ( .D(Key[130]), .CK(clk), .Q(reg_key[130]) );
  DFF_X1 \reg_key_reg[32]  ( .D(Key[32]), .CK(clk), .Q(reg_key[32]) );
  DFF_X1 \reg_key_reg[79]  ( .D(Key[79]), .CK(clk), .Q(reg_key[79]) );
  DFF_X1 \reg_key_reg[75]  ( .D(Key[75]), .CK(clk), .Q(reg_key[75]) );
  DFF_X1 \reg_key_reg[114]  ( .D(Key[114]), .CK(clk), .Q(reg_key[114]) );
  DFF_X1 \reg_key_reg[161]  ( .D(Key[161]), .CK(clk), .Q(reg_key[161]) );
  DFF_X1 \reg_key_reg[157]  ( .D(Key[157]), .CK(clk), .Q(reg_key[157]) );
  DFF_X1 \reg_key_reg[12]  ( .D(Key[12]), .CK(clk), .Q(reg_key[12]) );
  DFF_X1 \reg_key_reg[153]  ( .D(Key[153]), .CK(clk), .Q(reg_key[153]) );
  DFF_X1 \reg_key_reg[55]  ( .D(Key[55]), .CK(clk), .Q(reg_key[55]) );
  DFF_X1 \reg_key_reg[145]  ( .D(Key[145]), .CK(clk), .Q(reg_key[145]) );
  DFF_X1 \reg_key_reg[94]  ( .D(Key[94]), .CK(clk), .Q(reg_key[94]) );
  DFF_X1 \reg_key_reg[141]  ( .D(Key[141]), .CK(clk), .Q(reg_key[141]) );
  DFF_X1 \reg_key_reg[43]  ( .D(Key[43]), .CK(clk), .Q(reg_key[43]) );
  DFF_X1 \reg_key_reg[39]  ( .D(Key[39]), .CK(clk), .Q(reg_key[39]) );
  DFF_X1 \reg_key_reg[133]  ( .D(Key[133]), .CK(clk), .Q(reg_key[133]) );
  DFF_X1 \reg_key_reg[176]  ( .D(Key[176]), .CK(clk), .Q(reg_key[176]) );
  DFF_X1 \reg_key_reg[31]  ( .D(Key[31]), .CK(clk), .Q(reg_key[31]) );
  DFF_X1 \reg_key_reg[78]  ( .D(Key[78]), .CK(clk), .Q(reg_key[78]) );
  DFF_X1 \reg_key_reg[121]  ( .D(Key[121]), .CK(clk), .Q(reg_key[121]) );
  DFF_X1 \reg_key_reg[23]  ( .D(Key[23]), .CK(clk), .Q(reg_key[23]) );
  DFF_X1 \reg_key_reg[117]  ( .D(Key[117]), .CK(clk), .Q(reg_key[117]) );
  DFF_X1 \reg_key_reg[19]  ( .D(Key[19]), .CK(clk), .Q(reg_key[19]) );
  DFF_X1 \reg_key_reg[113]  ( .D(Key[113]), .CK(clk), .Q(reg_key[113]) );
  DFF_X1 \reg_key_reg[11]  ( .D(Key[11]), .CK(clk), .Q(reg_key[11]) );
  DFF_X1 \reg_key_reg[7]  ( .D(Key[7]), .CK(clk), .Q(reg_key[7]) );
  DFF_X1 \reg_key_reg[50]  ( .D(Key[50]), .CK(clk), .Q(reg_key[50]) );
  DFF_X1 \reg_key_reg[144]  ( .D(Key[144]), .CK(clk), .Q(reg_key[144]) );
  DFF_X1 \reg_key_reg[42]  ( .D(Key[42]), .CK(clk), .Q(reg_key[42]) );
  DFF_X1 \reg_key_reg[89]  ( .D(Key[89]), .CK(clk), .Q(reg_key[89]) );
  DFF_X1 \reg_key_reg[85]  ( .D(Key[85]), .CK(clk), .Q(reg_key[85]) );
  DFF_X1 \reg_key_reg[34]  ( .D(Key[34]), .CK(clk), .Q(reg_key[34]) );
  DFF_X1 \reg_key_reg[128]  ( .D(Key[128]), .CK(clk), .Q(reg_key[128]) );
  DFF_X1 \reg_key_reg[26]  ( .D(Key[26]), .CK(clk), .Q(reg_key[26]) );
  DFF_X1 \reg_key_reg[90]  ( .D(Key[90]), .CK(clk), .Q(reg_key[90]) );
  DFF_X1 \reg_key_reg[93]  ( .D(Key[93]), .CK(clk), .Q(reg_key[93]) );
  DFF_X1 \reg_key_reg[52]  ( .D(Key[52]), .CK(clk), .Q(reg_key[52]) );
  DFF_X1 \reg_key_reg[167]  ( .D(Key[167]), .CK(clk), .Q(reg_key[167]) );
  DFF_X1 \reg_key_reg[53]  ( .D(Key[53]), .CK(clk), .Q(reg_key[53]) );
  DFF_X1 \reg_key_reg[64]  ( .D(Key[64]), .CK(clk), .Q(reg_key[64]) );
  DFF_X1 \reg_key_reg[91]  ( .D(Key[91]), .CK(clk), .Q(reg_key[91]) );
  DFF_X1 \reg_key_reg[126]  ( .D(Key[126]), .CK(clk), .Q(reg_key[126]) );
  DFF_X1 \reg_key_reg[175]  ( .D(Key[175]), .CK(clk), .Q(reg_key[175]) );
  DFF_X1 \reg_key_reg[33]  ( .D(Key[33]), .CK(clk), .Q(reg_key[33]) );
  DFF_X1 \reg_key_reg[112]  ( .D(Key[112]), .CK(clk), .Q(reg_key[112]) );
  DFF_X1 \reg_key_reg[139]  ( .D(Key[139]), .CK(clk), .Q(reg_key[139]) );
  DFF_X1 \reg_key_reg[127]  ( .D(Key[127]), .CK(clk), .Q(reg_key[127]) );
  DFF_X1 \reg_key_reg[142]  ( .D(Key[142]), .CK(clk), .Q(reg_key[142]) );
  DFF_X1 \reg_key_reg[110]  ( .D(Key[110]), .CK(clk), .Q(reg_key[110]) );
  DFF_X1 \reg_key_reg[62]  ( .D(Key[62]), .CK(clk), .Q(reg_key[62]) );
  DFF_X1 \reg_key_reg[164]  ( .D(Key[164]), .CK(clk), .Q(reg_key[164]) );
  DFF_X1 \reg_key_reg[97]  ( .D(Key[97]), .CK(clk), .Q(reg_key[97]) );
  DFF_X1 \reg_key_reg[168]  ( .D(Key[168]), .CK(clk), .Q(reg_key[168]) );
  DFF_X1 \reg_key_reg[115]  ( .D(Key[115]), .CK(clk), .Q(reg_key[115]) );
  DFF_X1 \reg_key_reg[162]  ( .D(Key[162]), .CK(clk), .Q(reg_key[162]) );
  DFF_X1 \reg_key_reg[37]  ( .D(Key[37]), .CK(clk), .Q(reg_key[37]) );
  DFF_X1 \reg_key_reg[129]  ( .D(Key[129]), .CK(clk), .Q(reg_key[129]) );
  DFF_X1 \reg_key_reg[124]  ( .D(Key[124]), .CK(clk), .Q(reg_key[124]) );
  DFF_X1 \reg_key_reg[69]  ( .D(Key[69]), .CK(clk), .Q(reg_key[69]) );
  DFF_X1 \reg_key_reg[73]  ( .D(Key[73]), .CK(clk), .Q(reg_key[73]) );
  DFF_X1 \reg_key_reg[46]  ( .D(Key[46]), .CK(clk), .Q(reg_key[46]) );
  DFF_X1 \reg_key_reg[57]  ( .D(Key[57]), .CK(clk), .Q(reg_key[57]) );
  DFF_X1 \reg_key_reg[180]  ( .D(Key[180]), .CK(clk), .Q(reg_key[180]) );
  DFF_X1 \reg_key_reg[77]  ( .D(Key[77]), .CK(clk), .Q(reg_key[77]) );
  DFF_X1 \reg_key_reg[47]  ( .D(Key[47]), .CK(clk), .Q(reg_key[47]) );
  DFF_X1 \reg_key_reg[0]  ( .D(Key[0]), .CK(clk), .Q(reg_key[0]) );
  DFF_X1 \reg_key_reg[67]  ( .D(Key[67]), .CK(clk), .Q(reg_key[67]) );
  DFF_X1 \reg_key_reg[166]  ( .D(Key[166]), .CK(clk), .Q(reg_key[166]) );
  DFF_X1 \reg_key_reg[136]  ( .D(Key[136]), .CK(clk), .Q(reg_key[136]) );
  DFF_X1 \reg_key_reg[70]  ( .D(Key[70]), .CK(clk), .Q(reg_key[70]) );
  DFF_X1 \reg_key_reg[148]  ( .D(Key[148]), .CK(clk), .Q(reg_key[148]) );
  DFF_X1 \reg_key_reg[88]  ( .D(Key[88]), .CK(clk), .Q(reg_key[88]) );
  DFF_X1 \reg_key_reg[174]  ( .D(Key[174]), .CK(clk), .Q(reg_key[174]) );
  DFFRS_X1 \Ciphertext_reg[42]  ( .D(reg_out[42]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Ciphertext[42]) );
  DFF_X1 \Ciphertext_reg[21]  ( .D(reg_out[21]), .CK(clk), .Q(Ciphertext[21])
         );
  DFF_X1 \Ciphertext_reg[65]  ( .D(reg_out[65]), .CK(clk), .Q(Ciphertext[65])
         );
  DFF_X1 \Ciphertext_reg[105]  ( .D(reg_out[105]), .CK(clk), .Q(
        Ciphertext[105]) );
  DFF_X1 \Ciphertext_reg[27]  ( .D(reg_out[27]), .CK(clk), .Q(Ciphertext[27])
         );
  DFF_X1 \Ciphertext_reg[133]  ( .D(reg_out[133]), .CK(clk), .Q(
        Ciphertext[133]) );
  DFF_X1 \Ciphertext_reg[154]  ( .D(reg_out[154]), .CK(clk), .Q(
        Ciphertext[154]) );
  DFF_X1 \Ciphertext_reg[103]  ( .D(reg_out[103]), .CK(clk), .Q(
        Ciphertext[103]) );
  DFF_X1 \Ciphertext_reg[73]  ( .D(reg_out[73]), .CK(clk), .Q(Ciphertext[73])
         );
  DFF_X1 \Ciphertext_reg[90]  ( .D(reg_out[90]), .CK(clk), .Q(Ciphertext[90])
         );
  DFF_X1 \Ciphertext_reg[39]  ( .D(reg_out[39]), .CK(clk), .Q(Ciphertext[39])
         );
  DFF_X1 \Ciphertext_reg[132]  ( .D(reg_out[132]), .CK(clk), .Q(
        Ciphertext[132]) );
  DFF_X1 \Ciphertext_reg[79]  ( .D(reg_out[79]), .CK(clk), .Q(Ciphertext[79])
         );
  DFF_X1 \Ciphertext_reg[3]  ( .D(reg_out[3]), .CK(clk), .Q(Ciphertext[3]) );
  DFF_X1 \Ciphertext_reg[50]  ( .D(reg_out[50]), .CK(clk), .Q(Ciphertext[50])
         );
  DFF_X1 \Ciphertext_reg[24]  ( .D(reg_out[24]), .CK(clk), .Q(Ciphertext[24])
         );
  DFF_X1 \Ciphertext_reg[80]  ( .D(reg_out[80]), .CK(clk), .Q(Ciphertext[80])
         );
  DFF_X1 \Ciphertext_reg[157]  ( .D(reg_out[157]), .CK(clk), .Q(
        Ciphertext[157]) );
  DFF_X1 \Ciphertext_reg[114]  ( .D(reg_out[114]), .CK(clk), .Q(
        Ciphertext[114]) );
  DFF_X1 \Ciphertext_reg[94]  ( .D(reg_out[94]), .CK(clk), .Q(Ciphertext[94])
         );
  DFF_X1 \Ciphertext_reg[38]  ( .D(reg_out[38]), .CK(clk), .Q(Ciphertext[38])
         );
  DFF_X1 \Ciphertext_reg[68]  ( .D(reg_out[68]), .CK(clk), .Q(Ciphertext[68])
         );
  DFF_X1 \Ciphertext_reg[70]  ( .D(reg_out[70]), .CK(clk), .Q(Ciphertext[70])
         );
  DFF_X1 \Ciphertext_reg[45]  ( .D(reg_out[45]), .CK(clk), .Q(Ciphertext[45])
         );
  DFF_X1 \Ciphertext_reg[7]  ( .D(reg_out[7]), .CK(clk), .Q(Ciphertext[7]) );
  DFF_X1 \Ciphertext_reg[191]  ( .D(reg_out[191]), .CK(clk), .Q(
        Ciphertext[191]) );
  DFF_X1 \Ciphertext_reg[180]  ( .D(reg_out[180]), .CK(clk), .Q(
        Ciphertext[180]) );
  DFF_X2 \reg_key_reg[172]  ( .D(Key[172]), .CK(clk), .Q(reg_key[172]) );
  DFF_X2 \Ciphertext_reg[176]  ( .D(reg_out[176]), .CK(clk), .Q(
        Ciphertext[176]) );
  DFF_X1 \Ciphertext_reg[172]  ( .D(reg_out[172]), .CK(clk), .Q(
        Ciphertext[172]) );
  SPEEDY_Rounds6_0 SPEEDY_instance ( .Plaintext(reg_in), .Key(reg_key), 
        .Ciphertext(reg_out) );
  DFFRS_X1 \Ciphertext_reg[53]  ( .D(reg_out[53]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Ciphertext[53]) );
  DFFS_X1 \Ciphertext_reg[96]  ( .D(reg_out[96]), .CK(clk), .SN(1'b1), .Q(
        Ciphertext[96]) );
  DFF_X1 \Ciphertext_reg[1]  ( .D(reg_out[1]), .CK(clk), .Q(Ciphertext[1]) );
  DFF_X1 \Ciphertext_reg[69]  ( .D(reg_out[69]), .CK(clk), .Q(Ciphertext[69])
         );
  DFF_X1 \Ciphertext_reg[63]  ( .D(reg_out[63]), .CK(clk), .Q(Ciphertext[63])
         );
  DFF_X1 \Ciphertext_reg[19]  ( .D(reg_out[19]), .CK(clk), .Q(Ciphertext[19])
         );
  DFF_X1 \Ciphertext_reg[175]  ( .D(reg_out[175]), .CK(clk), .Q(
        Ciphertext[175]) );
  DFF_X1 \Ciphertext_reg[104]  ( .D(reg_out[104]), .CK(clk), .Q(
        Ciphertext[104]) );
  DFF_X1 \Ciphertext_reg[117]  ( .D(reg_out[117]), .CK(clk), .Q(
        Ciphertext[117]) );
  DFF_X1 \Ciphertext_reg[67]  ( .D(reg_out[67]), .CK(clk), .Q(Ciphertext[67])
         );
  DFF_X1 \Ciphertext_reg[115]  ( .D(reg_out[115]), .CK(clk), .Q(
        Ciphertext[115]) );
  DFF_X1 \Ciphertext_reg[151]  ( .D(reg_out[151]), .CK(clk), .Q(
        Ciphertext[151]) );
  DFF_X1 \Ciphertext_reg[44]  ( .D(reg_out[44]), .CK(clk), .Q(Ciphertext[44])
         );
  DFF_X1 \Ciphertext_reg[109]  ( .D(reg_out[109]), .CK(clk), .Q(
        Ciphertext[109]) );
  DFF_X1 \Ciphertext_reg[43]  ( .D(reg_out[43]), .CK(clk), .Q(Ciphertext[43])
         );
  DFF_X1 \Ciphertext_reg[20]  ( .D(reg_out[20]), .CK(clk), .Q(Ciphertext[20])
         );
  DFF_X1 \Ciphertext_reg[178]  ( .D(reg_out[178]), .CK(clk), .Q(
        Ciphertext[178]) );
  DFF_X1 \Ciphertext_reg[81]  ( .D(reg_out[81]), .CK(clk), .Q(Ciphertext[81])
         );
  DFF_X1 \Ciphertext_reg[127]  ( .D(reg_out[127]), .CK(clk), .Q(
        Ciphertext[127]) );
  DFF_X1 \Ciphertext_reg[99]  ( .D(reg_out[99]), .CK(clk), .Q(Ciphertext[99])
         );
  DFF_X1 \Ciphertext_reg[85]  ( .D(reg_out[85]), .CK(clk), .Q(Ciphertext[85])
         );
  DFF_X1 \Ciphertext_reg[97]  ( .D(reg_out[97]), .CK(clk), .Q(Ciphertext[97])
         );
  DFF_X1 \Ciphertext_reg[36]  ( .D(reg_out[36]), .CK(clk), .Q(Ciphertext[36])
         );
  DFF_X1 \Ciphertext_reg[166]  ( .D(reg_out[166]), .CK(clk), .Q(
        Ciphertext[166]) );
  DFF_X1 \Ciphertext_reg[60]  ( .D(reg_out[60]), .CK(clk), .Q(Ciphertext[60])
         );
  DFF_X1 \Ciphertext_reg[119]  ( .D(reg_out[119]), .CK(clk), .Q(
        Ciphertext[119]) );
  DFF_X1 \Ciphertext_reg[150]  ( .D(reg_out[150]), .CK(clk), .Q(
        Ciphertext[150]) );
  DFF_X1 \Ciphertext_reg[111]  ( .D(reg_out[111]), .CK(clk), .Q(
        Ciphertext[111]) );
  DFF_X1 \Ciphertext_reg[102]  ( .D(reg_out[102]), .CK(clk), .Q(
        Ciphertext[102]) );
  DFF_X1 \Ciphertext_reg[134]  ( .D(reg_out[134]), .CK(clk), .Q(
        Ciphertext[134]) );
  DFF_X1 \Ciphertext_reg[144]  ( .D(reg_out[144]), .CK(clk), .Q(
        Ciphertext[144]) );
  DFF_X1 \Ciphertext_reg[182]  ( .D(reg_out[182]), .CK(clk), .Q(
        Ciphertext[182]) );
  DFF_X1 \Ciphertext_reg[52]  ( .D(reg_out[52]), .CK(clk), .Q(Ciphertext[52])
         );
  DFF_X1 \Ciphertext_reg[16]  ( .D(reg_out[16]), .CK(clk), .Q(Ciphertext[16])
         );
  DFF_X1 \Ciphertext_reg[161]  ( .D(reg_out[161]), .CK(clk), .Q(
        Ciphertext[161]) );
  DFF_X1 \Ciphertext_reg[186]  ( .D(reg_out[186]), .CK(clk), .Q(
        Ciphertext[186]) );
  DFF_X1 \Ciphertext_reg[179]  ( .D(reg_out[179]), .CK(clk), .Q(
        Ciphertext[179]) );
  DFF_X1 \Ciphertext_reg[61]  ( .D(reg_out[61]), .CK(clk), .Q(Ciphertext[61])
         );
  DFF_X1 \Ciphertext_reg[95]  ( .D(reg_out[95]), .CK(clk), .Q(Ciphertext[95])
         );
  DFF_X1 \Ciphertext_reg[107]  ( .D(reg_out[107]), .CK(clk), .Q(
        Ciphertext[107]) );
  DFF_X1 \Ciphertext_reg[75]  ( .D(reg_out[75]), .CK(clk), .Q(Ciphertext[75])
         );
  DFF_X1 \Ciphertext_reg[110]  ( .D(reg_out[110]), .CK(clk), .Q(
        Ciphertext[110]) );
  DFF_X1 \Ciphertext_reg[51]  ( .D(reg_out[51]), .CK(clk), .Q(Ciphertext[51])
         );
  DFF_X1 \Ciphertext_reg[184]  ( .D(reg_out[184]), .CK(clk), .Q(
        Ciphertext[184]) );
  DFF_X1 \Ciphertext_reg[71]  ( .D(reg_out[71]), .CK(clk), .Q(Ciphertext[71])
         );
  DFF_X1 \Ciphertext_reg[123]  ( .D(reg_out[123]), .CK(clk), .Q(
        Ciphertext[123]) );
  DFF_X1 \Ciphertext_reg[58]  ( .D(reg_out[58]), .CK(clk), .Q(Ciphertext[58])
         );
  DFF_X1 \Ciphertext_reg[93]  ( .D(reg_out[93]), .CK(clk), .Q(Ciphertext[93])
         );
  DFF_X1 \Ciphertext_reg[66]  ( .D(reg_out[66]), .CK(clk), .Q(Ciphertext[66])
         );
  DFF_X1 \Ciphertext_reg[76]  ( .D(reg_out[76]), .CK(clk), .Q(Ciphertext[76])
         );
  DFF_X1 \Ciphertext_reg[25]  ( .D(reg_out[25]), .CK(clk), .Q(Ciphertext[25])
         );
  DFF_X1 \Ciphertext_reg[113]  ( .D(reg_out[113]), .CK(clk), .Q(
        Ciphertext[113]) );
  DFF_X1 \Ciphertext_reg[59]  ( .D(reg_out[59]), .CK(clk), .Q(Ciphertext[59])
         );
  DFF_X1 \Ciphertext_reg[48]  ( .D(reg_out[48]), .CK(clk), .Q(Ciphertext[48])
         );
  DFF_X1 \Ciphertext_reg[156]  ( .D(reg_out[156]), .CK(clk), .Q(
        Ciphertext[156]) );
  DFF_X1 \Ciphertext_reg[174]  ( .D(reg_out[174]), .CK(clk), .Q(
        Ciphertext[174]) );
  DFF_X1 \Ciphertext_reg[9]  ( .D(reg_out[9]), .CK(clk), .Q(Ciphertext[9]) );
  DFF_X1 \Ciphertext_reg[153]  ( .D(reg_out[153]), .CK(clk), .Q(
        Ciphertext[153]) );
  DFF_X1 \Ciphertext_reg[47]  ( .D(reg_out[47]), .CK(clk), .Q(Ciphertext[47])
         );
  DFF_X1 \Ciphertext_reg[173]  ( .D(reg_out[173]), .CK(clk), .Q(
        Ciphertext[173]) );
  DFF_X1 \Ciphertext_reg[146]  ( .D(reg_out[146]), .CK(clk), .Q(
        Ciphertext[146]) );
  DFF_X1 \Ciphertext_reg[55]  ( .D(reg_out[55]), .CK(clk), .Q(Ciphertext[55])
         );
  DFF_X1 \Ciphertext_reg[162]  ( .D(reg_out[162]), .CK(clk), .Q(
        Ciphertext[162]) );
  DFF_X1 \Ciphertext_reg[78]  ( .D(reg_out[78]), .CK(clk), .Q(Ciphertext[78])
         );
  DFF_X1 \Ciphertext_reg[121]  ( .D(reg_out[121]), .CK(clk), .Q(
        Ciphertext[121]) );
  DFF_X1 \Ciphertext_reg[181]  ( .D(reg_out[181]), .CK(clk), .Q(
        Ciphertext[181]) );
  DFF_X1 \Ciphertext_reg[22]  ( .D(reg_out[22]), .CK(clk), .Q(Ciphertext[22])
         );
  DFF_X1 \Ciphertext_reg[40]  ( .D(reg_out[40]), .CK(clk), .Q(Ciphertext[40])
         );
  DFF_X1 \Ciphertext_reg[189]  ( .D(reg_out[189]), .CK(clk), .Q(
        Ciphertext[189]) );
  DFF_X1 \Ciphertext_reg[12]  ( .D(reg_out[12]), .CK(clk), .Q(Ciphertext[12])
         );
endmodule

