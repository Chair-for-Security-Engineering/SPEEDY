module SPEEDY_Rounds7_0 ( Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  wire   n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19,
         n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37,
         n39, n40, n41, n42, n43, n44, n46, n48, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n63, n64, n66, n69, n71, n72, n73, n75, n76,
         n77, n79, n80, n81, n82, n84, n85, n87, n88, n89, n91, n92, n96, n97,
         n100, n101, n104, n105, n106, n107, n109, n111, n112, n113, n114,
         n117, n118, n119, n120, n121, n122, n123, n125, n127, n128, n130,
         n132, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n153, n155, n156, n157, n159,
         n161, n162, n163, n165, n167, n168, n169, n170, n171, n172, n174,
         n175, n178, n179, n180, n181, n182, n183, n184, n186, n187, n188,
         n189, n190, n191, n192, n193, n195, n196, n197, n198, n199, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n215, n216, n217, n219, n220, n221, n223, n224, n225, n226,
         n227, n229, n231, n232, n233, n235, n237, n238, n240, n241, n242,
         n243, n244, n245, n248, n249, n250, n251, n252, n253, n255, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n283, n284, n285, n287, n292, n293, n294, n295, n296, n297,
         n300, n301, n303, n306, n307, n308, n320, n321, n323, n324, n325,
         n326, n329, n333, n336, n337, n339, n341, n342, n349, n351, n355,
         n359, n363, n365, n370, n371, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n393, n394, n395, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n412, n413, n414, n415,
         n416, n417, n418, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n449, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n468, n469, n470, n471, n473, n474, n475, n476, n477, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n538, n539, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n577, n578, n579, n580, n581, n582, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n612, n613, n614, n615, n616, n617, n618, n619, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n678, n679,
         n680, n681, n683, n686, n688, n689, n690, n691, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n717, n719, n720,
         n721, n722, n724, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n753, n754, n755, n756, n757,
         n758, n760, n761, n762, n763, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n790, n792, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n834, n835, n836, n837, n839, n840, n841, n842,
         n843, n844, n846, n847, n848, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n903, n905, n906, n907, n908, n909, n910, n912, n913,
         n914, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n951, n952, n953, n954, n956, n957, n958, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n977, n980, n981, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1028, n1029, n1030, n1032,
         n1033, n1034, n1035, n1037, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1073, n1075, n1076, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1094, n1095, n1096, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1137, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1148, n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1169,
         n1170, n1171, n1172, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1196, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1223, n1224,
         n1225, n1226, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1326, n1327, n1328, n1329, n1330,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1342,
         n1344, n1345, n1346, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1361, n1362, n1363, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1410,
         n1411, n1412, n1413, n1415, n1416, n1417, n1418, n1419, n1420, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1433, n1434,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1487, n1489, n1490, n1491,
         n1493, n1494, n1495, n1496, n1497, n1498, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1558, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1574, n1575, n1576, n1577, n1580,
         n1581, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1634, n1635, n1637,
         n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1673, n1674, n1675, n1676, n1679, n1681, n1683,
         n1684, n1685, n1686, n1687, n1688, n1690, n1691, n1692, n1693, n1694,
         n1695, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1720, n1721, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1828, n1829, n1830, n1831, n1832, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1861, n1862, n1863, n1864, n1865, n1868,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1883, n1884, n1885, n1886, n1887, n1888, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1933, n1934,
         n1938, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2096, n2097, n2098, n2099, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2157, n2158, n2159, n2160, n2161, n2162, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2196, n2199, n2200,
         n2201, n2202, n2203, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2234, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2246, n2247, n2248, n2250, n2251, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2278, n2281, n2282,
         n2283, n2285, n2286, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2323, n2324, n2325, n2326, n2327,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2355, n2357, n2358, n2359, n2360,
         n2361, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2437, n2438, n2439, n2440, n2441, n2442, n2444, n2445,
         n2446, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2480, n2481, n2482, n2483, n2484, n2485, n2487, n2488, n2489, n2490,
         n2491, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2514, n2516, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2538,
         n2539, n2541, n2542, n2544, n2545, n2546, n2547, n2549, n2551, n2552,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2589, n2590, n2591, n2592, n2593, n2594,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2655, n2656, n2657, n2658, n2659,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2675, n2676, n2677, n2678, n2680, n2681, n2682, n2683, n2684,
         n2685, n2687, n2688, n2689, n2690, n2691, n2692, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2704, n2705, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2882,
         n2883, n2884, n2885, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2911, n2912, n2913, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2934, n2935, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2954, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2999, n3001, n3002, n3003, n3004, n3005, n3006,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3097, n3099, n3100, n3101,
         n3103, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3121, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3210, n3211,
         n3212, n3213, n3214, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3254, n3255,
         n3256, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3266, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3325, n3326, n3328, n3329, n3330, n3331, n3332, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3356, n3357, n3359, n3360, n3361, n3362, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3382, n3383, n3384, n3385, n3386, n3387, n3390, n3391, n3392,
         n3393, n3395, n3396, n3397, n3400, n3401, n3402, n3403, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3413, n3414, n3415, n3416, n3417,
         n3418, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3466, n3467, n3468, n3469,
         n3470, n3471, n3473, n3474, n3475, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3745,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3768, n3770, n3771, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3917, n3918, n3919, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3983, n3984, n3985, n3986, n3987,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4132, n4133,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4184, n4185, n4186, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4206, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4258,
         n4259, n4260, n4261, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4290,
         n4291, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4438, n4439, n4440, n4441, n4442, n4443, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4472, n4473, n4474, n4476, n4477, n4478, n4479, n4480, n4482, n4483,
         n4484, n4485, n4486, n4487, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4705, n4706, n4707, n4708, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4741, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4772, n4773, n4774, n4776, n4777, n4778, n4779, n4780,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4900,
         n4901, n4902, n4903, n4904, n4905, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4950, n4951, n4953, n4954,
         n4955, n4956, n4957, n4959, n4960, n4961, n4962, n4963, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5066, n5067, n5068, n5069, n5070,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5086, n5087, n5088, n5089, n5090, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5109, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5146, n5147, n5148, n5149,
         n5150, n5151, n5154, n5155, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5184, n5185, n5186, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5221, n5222, n5223, n5224, n5225, n5226,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5248,
         n5250, n5251, n5252, n5253, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5272, n5273,
         n5274, n5275, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5287, n5288, n5289, n5291, n5292, n5293, n5294, n5295, n5297,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5341,
         n5342, n5343, n5344, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5381, n5382, n5383,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5439, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5504, n5505, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5581, n5582, n5584, n5585, n5586,
         n5587, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5709, n5710, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5763, n5764, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5801, n5802, n5803, n5804, n5805, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5830, n5831, n5832, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5862, n5863, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6097, n6098, n6099,
         n6100, n6101, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6128, n6130, n6132, n6133,
         n6134, n6135, n6136, n6137, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6252, n6253, n6254, n6255, n6256, n6257, n6259, n6260,
         n6261, n6262, n6264, n6265, n6266, n6267, n6268, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6304, n6305, n6306, n6307, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6332, n6333, n6335, n6336,
         n6337, n6338, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6396, n6397, n6398, n6399, n6400, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6461, n6462, n6464, n6465, n6466,
         n6467, n6468, n6469, n6472, n6474, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6487, n6488, n6489, n6490, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6524,
         n6526, n6527, n6528, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6584, n6585, n6586, n6587, n6588, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6631, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6642, n6643, n6644, n6645,
         n6646, n6647, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6677,
         n6678, n6679, n6680, n6681, n6683, n6685, n6686, n6687, n6688, n6689,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6727, n6728, n6729, n6730, n6731, n6733,
         n6734, n6735, n6736, n6737, n6738, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6777, n6778, n6779, n6780, n6782, n6783, n6785, n6786, n6787,
         n6788, n6789, n6790, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7013, n7014, n7015, n7016,
         n7017, n7018, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7451, n7452, n7454, n7456,
         n7457, n7458, n7459, n7460, n7461, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8094, n8097,
         n8098, n8099, n8100, n8101, n8102, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8326, n8327, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8359, n8360, n8361, n8362, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8426, n8427, n8428, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8540, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8715, n8716, n8717, n8718, n8719, n8720,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8779, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9368, n9369, n9370, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10406, n10407, n10408, n10409, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10482, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10492, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10511, n10512, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10589, n10590, n10591, n10592,
         n10593, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10611, n10612, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10867, n10868, n10869, n10870, n10871, n10872, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10976, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11174, n11175, n11176, n11178, n11179, n11180, n11181,
         n11183, n11184, n11185, n11186, n11187, n11188, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11264, n11265, n11266, n11267,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11650, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11841, n11843, n11844, n11845,
         n11846, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11907, n11908, n11909, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12037,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12083, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12106,
         n12107, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12255,
         n12256, n12257, n12258, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12938, n12939, n12940,
         n12941, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13620, n13621, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13732, n13733, n13734, n13735, n13736, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13778, n13779, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13898,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13938, n13939, n13940, n13941,
         n13943, n13944, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14197, n14198, n14199, n14200, n14202, n14203, n14204,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14511, n14512, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14960, n14961, n14962, n14963, n14964, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15040,
         n15041, n15042, n15043, n15044, n15046, n15047, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15920, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16848, n16849, n16850, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16964, n16965, n16966, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16985, n16986, n16987, n16988,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17029, n17030, n17031,
         n17033, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17049, n17051,
         n17052, n17053, n17054, n17055, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17087, n17088, n17089, n17090, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17128, n17129, n17130,
         n17131, n17132, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17164, n17165,
         n17166, n17167, n17169, n17170, n17171, n17172, n17173, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17368, n17369, n17370, n17371, n17372, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17610, n17611, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17785, n17788, n17789, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17801, n17802, n17803, n17804, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17895, n17896, n17897, n17898, n17899,
         n17900, n17902, n17903, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17915, n17916, n17917, n17918,
         n17919, n17920, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18015, n18016, n18017, n18018,
         n18019, n18020, n18022, n18023, n18024, n18025, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18576, n18577, n18578, n18579, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18833, n18834, n18835,
         n18836, n18837, n18838, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19187,
         n19188, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19254, n19256,
         n19257, n19258, n19259, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19832, n19833, n19834,
         n19836, n19837, n19838, n19839, n19841, n19842, n19843, n19844,
         n19846, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19906, n19907, n19908, n19909, n19911, n19912, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19923,
         n19924, n19925, n19926, n19927, n19928, n19930, n19931, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20077,
         n20078, n20079, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20268, n20269,
         n20270, n20271, n20272, n20273, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20400, n20401,
         n20402, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20520, n20521, n20522, n20523, n20524, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20537, n20539, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20570,
         n20571, n20572, n20573, n20574, n20575, n20577, n20578, n20579,
         n20580, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21047, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21101,
         n21102, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21161, n21162, n21163, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21467, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21499, n21500,
         n21501, n21503, n21504, n21505, n21506, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21864, n21865, n21866, n21867, n21868, n21870,
         n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
         n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
         n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
         n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
         n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
         n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918,
         n21919, n21920, n21921, n21922, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
         n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
         n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077,
         n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
         n22086, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
         n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102,
         n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110,
         n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
         n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
         n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
         n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
         n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
         n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
         n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
         n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
         n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
         n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
         n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206,
         n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
         n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230,
         n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
         n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
         n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278,
         n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
         n22287, n22288, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22633, n22634, n22635, n22636,
         n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
         n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
         n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
         n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
         n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
         n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
         n22685, n22686, n22688, n22689, n22690, n22691, n22692, n22693,
         n22694, n22695, n22696, n22697, n22698, n22699, n22701, n22702,
         n22703, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,
         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22841,
         n22842, n22843, n22844, n22845, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
         n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890,
         n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
         n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
         n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
         n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
         n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
         n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
         n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
         n22955, n22956, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22967, n22968, n22969, n22970, n22971, n22972,
         n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980,
         n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
         n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
         n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
         n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23014,
         n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022,
         n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030,
         n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038,
         n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046,
         n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054,
         n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062,
         n23063, n23065, n23066, n23067, n23068, n23069, n23070, n23072,
         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23096, n23097, n23098,
         n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106,
         n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
         n23115, n23116, n23117, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23159, n23161, n23162, n23163, n23164, n23165,
         n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173,
         n23174, n23175, n23176, n23177, n23179, n23180, n23181, n23182,
         n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190,
         n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23200,
         n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
         n23209, n23210, n23211, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23224, n23225, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23235, n23236,
         n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244,
         n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252,
         n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260,
         n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268,
         n23269, n23270, n23271, n23272, n23273, n23274, n23276, n23277,
         n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285,
         n23286, n23287, n23289, n23290, n23291, n23292, n23293, n23294,
         n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302,
         n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23311,
         n23313, n23314, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23326, n23327, n23328, n23329, n23330,
         n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
         n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346,
         n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23422, n23423, n23424, n23426, n23427, n23428, n23429,
         n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
         n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445,
         n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23454,
         n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462,
         n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470,
         n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478,
         n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486,
         n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
         n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502,
         n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510,
         n23511, n23512, n23513, n23514, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23531, n23532, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23593, n23594, n23595, n23596,
         n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604,
         n23605, n23606, n23607, n23608, n23610, n23611, n23612, n23613,
         n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622,
         n23623, n23624, n23625, n23626, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23662, n23663, n23664,
         n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,
         n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
         n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688,
         n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,
         n23697, n23698, n23699, n23700, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23751, n23752, n23753, n23754,
         n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
         n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
         n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778,
         n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
         n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
         n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
         n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
         n23811, n23812, n23813, n23814, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23825, n23827, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23837, n23838, n23839, n23840,
         n23841, n23842, n23843, n23845, n23846, n23848, n23849, n23850,
         n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860,
         n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868,
         n23869, n23870, n23871, n23874, n23875, n23876, n23877, n23878,
         n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886,
         n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894,
         n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23926, n23927, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23944, n23945, n23946,
         n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954,
         n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
         n23963, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23984, n23985, n23986, n23987, n23988,
         n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23997,
         n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24006,
         n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
         n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24024,
         n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
         n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
         n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048,
         n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
         n24057, n24058, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24104, n24105, n24106,
         n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114,
         n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122,
         n24123, n24124, n24125, n24126, n24128, n24129, n24130, n24131,
         n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140,
         n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148,
         n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156,
         n24157, n24158, n24159, n24160, n24162, n24163, n24164, n24165,
         n24166, n24167, n24168, n24169, n24170, n24171, n24173, n24174,
         n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182,
         n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
         n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198,
         n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206,
         n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
         n24215, n24216, n24218, n24219, n24220, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
         n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255,
         n24256, n24257, n24258, n24259, n24261, n24262, n24263, n24264,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24282,
         n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
         n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
         n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306,
         n24307, n24308, n24310, n24311, n24312, n24314, n24315, n24316,
         n24317, n24318, n24319, n24322, n24323, n24324, n24325, n24326,
         n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334,
         n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342,
         n24343, n24345, n24347, n24348, n24349, n24350, n24351, n24352,
         n24353, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24376, n24377, n24378,
         n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
         n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
         n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402,
         n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410,
         n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418,
         n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426,
         n24427, n24428, n24429, n24430, n24433, n24434, n24435, n24436,
         n24437, n24439, n24440, n24441, n24442, n24443, n24444, n24445,
         n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453,
         n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
         n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
         n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477,
         n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24486,
         n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494,
         n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
         n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510,
         n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518,
         n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
         n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534,
         n24535, n24537, n24538, n24539, n24540, n24541, n24542, n24543,
         n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
         n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
         n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567,
         n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
         n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
         n24592, n24593, n24595, n24596, n24597, n24598, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24623, n24624, n24625, n24626,
         n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
         n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642,
         n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
         n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24690, n24691, n24692,
         n24693, n24694, n24695, n24696, n24697, n24699, n24700, n24701,
         n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710,
         n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
         n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726,
         n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734,
         n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742,
         n24743, n24744, n24745, n24746, n24747, n24748, n24750, n24751,
         n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24760,
         n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,
         n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
         n24777, n24778, n24779, n24780, n24781, n24782, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24816, n24817, n24821, n24822,
         n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830,
         n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
         n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846,
         n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
         n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862,
         n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870,
         n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878,
         n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886,
         n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894,
         n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902,
         n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910,
         n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918,
         n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926,
         n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934,
         n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942,
         n24943, n24944, n24945, n24948, n24949, n24950, n24951, n24952,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24998, n24999, n25001, n25002, n25003, n25004,
         n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
         n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
         n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
         n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
         n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044,
         n25045, n25046, n25047, n25048, n25049, n25050, n25052, n25053,
         n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061,
         n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069,
         n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077,
         n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085,
         n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
         n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
         n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
         n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117,
         n25119, n25120, n25122, n25123, n25124, n25126, n25127, n25128,
         n25129, n25130, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25404, n25405,
         n25406, n25408, n25409, n25410, n25411, n25412, n25413, n25414,
         n25415, n25416, n25417, n25418, n25419, n25421, n25422, n25423,
         n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431,
         n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439,
         n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
         n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455,
         n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463,
         n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
         n25472, n25473, n25474, n25475, n25476, n25478, n25479, n25480,
         n25481, n25482, n25483, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
         n25629, n25631, n25632, n25633, n25634, n25635, n25636, n25637,
         n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
         n25646, n25647, n25649, n25650, n25651, n25652, n25653, n25654,
         n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662,
         n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670,
         n25671, n25672, n25674, n25675, n25676, n25677, n25678, n25679,
         n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
         n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695,
         n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
         n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711,
         n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719,
         n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
         n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
         n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
         n25744, n25745, n25746, n25747, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25844,
         n25845, n25846, n25847, n25848, n25849, n25851, n25852, n25853,
         n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861,
         n25862, n25864, n25865, n25866, n25867, n25868, n25869, n25870,
         n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878,
         n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
         n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894,
         n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902,
         n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
         n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918,
         n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926,
         n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934,
         n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
         n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950,
         n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
         n25959, n25960, n25961, n25963, n25964, n25965, n25966, n25968,
         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26066, n26067, n26068,
         n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076,
         n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084,
         n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092,
         n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100,
         n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
         n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116,
         n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124,
         n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132,
         n26133, n26135, n26136, n26137, n26138, n26139, n26140, n26141,
         n26142, n26144, n26145, n26146, n26147, n26148, n26151, n26153,
         n26154, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26166, n26168, n26169, n26170, n26171, n26172, n26173,
         n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181,
         n26182, n26183, n26184, n26185, n26186, n26187, n26189, n26190,
         n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
         n26199, n26200, n26201, n26203, n26204, n26205, n26206, n26207,
         n26208, n26209, n26210, n26212, n26213, n26214, n26215, n26216,
         n26217, n26218, n26219, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26332, n26333,
         n26334, n26335, n26336, n26337, n26338, n26339, n26341, n26342,
         n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350,
         n26351, n26352, n26354, n26355, n26356, n26357, n26358, n26359,
         n26360, n26361, n26362, n26363, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26389, n26390, n26392, n26394, n26395, n26396,
         n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404,
         n26406, n26408, n26409, n26410, n26412, n26413, n26414, n26415,
         n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
         n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
         n26432, n26433, n26434, n26435, n26436, n26437, n26439, n26440,
         n26441, n26442, n26443, n26444, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508,
         n26509, n26510, n26511, n26512, n26513, n26515, n26516, n26517,
         n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525,
         n26528, n26529, n26530, n26531, n26532, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26592, n26593, n26594, n26595, n26596,
         n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
         n26605, n26606, n26608, n26609, n26610, n26611, n26612, n26613,
         n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
         n26622, n26623, n26624, n26625, n26626, n26628, n26630, n26631,
         n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
         n26640, n26641, n26643, n26644, n26645, n26646, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26708,
         n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
         n26717, n26718, n26719, n26720, n26721, n26723, n26724, n26725,
         n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
         n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741,
         n26742, n26743, n26744, n26746, n26747, n26748, n26749, n26751,
         n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759,
         n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
         n26768, n26769, n26771, n26772, n26773, n26774, n26775, n26776,
         n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784,
         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
         n26793, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26846, n26848, n26849, n26850, n26851, n26852,
         n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
         n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868,
         n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876,
         n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
         n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
         n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
         n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908,
         n26909, n26910, n26911, n26912, n26914, n26915, n26916, n26917,
         n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925,
         n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
         n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
         n26942, n26943, n26944, n26946, n26948, n26949, n26950, n26951,
         n26952, n26953, n26954, n26956, n26957, n26958, n26959, n26960,
         n26961, n26962, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27041, n27043, n27044,
         n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052,
         n27053, n27054, n27055, n27056, n27057, n27058, n27060, n27061,
         n27062, n27063, n27064, n27065, n27066, n27067, n27069, n27070,
         n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078,
         n27079, n27080, n27081, n27083, n27084, n27085, n27086, n27087,
         n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
         n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
         n27104, n27105, n27106, n27107, n27109, n27110, n27111, n27112,
         n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120,
         n27121, n27122, n27123, n27124, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27175, n27177, n27178, n27179, n27180,
         n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
         n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
         n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205,
         n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213,
         n27214, n27215, n27216, n27217, n27219, n27220, n27221, n27222,
         n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
         n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238,
         n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246,
         n27247, n27248, n27249, n27250, n27252, n27253, n27254, n27255,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27374, n27375, n27376, n27377, n27378, n27379, n27380,
         n27381, n27382, n27384, n27385, n27386, n27387, n27388, n27389,
         n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397,
         n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405,
         n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413,
         n27414, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
         n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431,
         n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439,
         n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447,
         n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27456,
         n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
         n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,
         n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,
         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,
         n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
         n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,
         n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,
         n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,
         n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528,
         n27529, n27530, n27531, n27532, n27533, n27534, n27537, n27538,
         n27539, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27588,
         n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596,
         n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
         n27605, n27606, n27607, n27608, n27609, n27610, n27612, n27613,
         n27614, n27615, n27616, n27617, n27619, n27620, n27621, n27622,
         n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630,
         n27631, n27632, n27633, n27634, n27636, n27637, n27638, n27639,
         n27640, n27641, n27642, n27643, n27645, n27646, n27647, n27648,
         n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656,
         n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664,
         n27666, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
         n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
         n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
         n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
         n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
         n27707, n27708, n27709, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27736, n27737, n27738, n27739, n27740,
         n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
         n27749, n27750, n27751, n27752, n27755, n27757, n27758, n27759,
         n27760, n27761, n27762, n27764, n27765, n27766, n27767, n27768,
         n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776,
         n27777, n27778, n27779, n27780, n27782, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27811, n27812,
         n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
         n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
         n27829, n27830, n27831, n27832, n27833, n27834, n27836, n27837,
         n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
         n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853,
         n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861,
         n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
         n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877,
         n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885,
         n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893,
         n27894, n27898, n27899, n27900, n27901, n27902, n27903, n27904,
         n27905, n27906, n27907, n27908, n27909, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27940, n27941, n27942, n27943, n27944, n27947, n27948,
         n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
         n27957, n27958, n27960, n27961, n27962, n27963, n27964, n27965,
         n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27974,
         n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982,
         n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990,
         n27991, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28078, n28079, n28080, n28081, n28083,
         n28084, n28086, n28087, n28088, n28089, n28090, n28091, n28092,
         n28093, n28094, n28095, n28096, n28097, n28099, n28100, n28101,
         n28102, n28103, n28104, n28105, n28107, n28108, n28109, n28110,
         n28111, n28112, n28114, n28115, n28116, n28121, n28122, n28126,
         n28130, n28133, n28140, n28142, n28143, n28144, n28147, n28149,
         n28155, n28157, n28161, n28162, n28164, n28171, n28172, n28173,
         n28174, n28175, n28176, n28177, n28179, n28180, n28181, n28182,
         n28183, n28184, n28185, n28186, n28187, n28188, n28191, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28210,
         n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218,
         n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226,
         n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28235,
         n28236, n28237, n28238, n28240, n28241, n28242, n28243, n28244,
         n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
         n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
         n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
         n28269, n28270, n28271, n28273, n28274, n28275, n28276, n28277,
         n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
         n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28294,
         n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302,
         n28303, n28305, n28306, n28307, n28308, n28309, n28310, n28311,
         n28312, n28313, n28314, n28315, n28316, n28317, n28319, n28320,
         n28321, n28322, n28323, n28324, n28326, n28327, n28329, n28330,
         n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28339,
         n28340, n28341, n28343, n28344, n28345, n28347, n28348, n28349,
         n28351, n28352, n28353, n28354, n28355, n28357, n28358, n28359,
         n28360, n28361, n28362, n28363, n28364, n28365, n28367, n28368,
         n28369, n28370, n28371, n28372, n28373, n28376, n28377, n28378,
         n28379, n28380, n28381, n28383, n28384, n28385, n28386, n28387,
         n28388, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
         n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404,
         n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412,
         n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
         n28421, n28422, n28423, n28424, n28425, n28426, n28428, n28429,
         n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437,
         n28438, n28439, n28440, n28441, n28442, n28444, n28445, n28446,
         n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454,
         n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462,
         n28465, n28466, n28467, n28468, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28499,
         n28500, n28501, n28503, n28504, n28505, n28506, n28507, n28508,
         n28509, n28510, n28512, n28513, n28514, n28515, n28516, n28517,
         n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525,
         n28526, n28527, n28528, n28530, n28531, n28532, n28534, n28535,
         n28536, n28538, n28540, n28541, n28542, n28543, n28544, n28545,
         n28547, n28548, n28549, n28550, n28551, n28552, n28554, n28555,
         n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
         n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572,
         n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580,
         n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588,
         n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596,
         n28597, n28598, n28600, n28601, n28602, n28603, n28604, n28605,
         n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613,
         n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621,
         n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28630,
         n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638,
         n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
         n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654,
         n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662,
         n28663, n28665, n28666, n28667, n28668, n28669, n28670, n28671,
         n28672, n28674, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28698,
         n28699, n28701, n28702, n28703, n28704, n28706, n28707, n28708,
         n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716,
         n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28725,
         n28726, n28727, n28728, n28729, n28730, n28732, n28733, n28734,
         n28736, n28737, n28738, n28739, n28741, n28742, n28743, n28744,
         n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752,
         n28753, n28754, n28756, n28757, n28759, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28771, n28775,
         n28776, n28779, n28783, n28785, n28789, n28790, n28791, n28792,
         n28793, n28794, n28796, n28797, n28798, n28800, n28801, n28802,
         n28803, n28804, n28805, n28806, n28807, n28808, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28836,
         n28837, n28838, n28839, n28840, n28841, n28842, n28844, n28845,
         n28847, n28848, n28849, n28851, n28852, n28853, n28854, n28855,
         n28856, n28857, n28858, n28860, n28861, n28862, n28863, n28864,
         n28866, n28867, n28869, n28871, n28872, n28874, n28875, n28876,
         n28877, n28878, n28879, n28882, n28883, n28885, n28886, n28887,
         n28888, n28889, n28890, n28891, n28892, n28894, n28895, n28896,
         n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904,
         n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912,
         n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920,
         n28921, n28922, n28923, n28924, n28928, n28929, n28930, n28931,
         n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940,
         n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
         n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956,
         n28958, n28960, n28961, n28962, n28963, n28964, n28965, n28966,
         n28967, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
         n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
         n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992,
         n28993, n28994, n28995, n28996, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29069, n29070, n29071, n29072, n29073, n29074,
         n29075, n29076, n29077, n29078, n29079, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29114, n29115, n29116,
         n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124,
         n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132,
         n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140,
         n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149,
         n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157,
         n29158, n29159, n29160, n29161, n29163, n29164, n29165, n29166,
         n29168, n29169, n29171, n29172, n29173, n29174, n29175, n29176,
         n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184,
         n29185, n29186, n29187, n29188, n29189, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29201, n29202,
         n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
         n29211, n29212, n29214, n29215, n29217, n29218, n29219, n29220,
         n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228,
         n29229, n29230, n29231, n29232, n29233, n29235, n29236, n29237,
         n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245,
         n29246, n29247, n29248, n29249, n29251, n29253, n29255, n29256,
         n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264,
         n29265, n29268, n29269, n29270, n29271, n29272, n29273, n29274,
         n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
         n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290,
         n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298,
         n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306,
         n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
         n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322,
         n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
         n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338,
         n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346,
         n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354,
         n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362,
         n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370,
         n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378,
         n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
         n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
         n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
         n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
         n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
         n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434,
         n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442,
         n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450,
         n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
         n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466,
         n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
         n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482,
         n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490,
         n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514,
         n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538,
         n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546,
         n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554,
         n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562,
         n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570,
         n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578,
         n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
         n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594,
         n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
         n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610,
         n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
         n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
         n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
         n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642,
         n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
         n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
         n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666,
         n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
         n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682,
         n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690,
         n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
         n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706,
         n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
         n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722,
         n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730,
         n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738,
         n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
         n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754,
         n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
         n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
         n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778,
         n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786,
         n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794,
         n29795, n29796, n29797, n29798, n29799, n29800, n29801;

  NAND2_X1 U1 ( .A1(n26973), .A2(n28213), .ZN(n114) );
  AOI22_X1 U2 ( .A1(n27917), .A2(n27918), .B1(n27907), .B2(n27906), .ZN(n27914) );
  INV_X1 U3 ( .A(n27671), .ZN(n85) );
  BUF_X1 U6 ( .A(n26652), .Z(n27539) );
  AND3_X1 U7 ( .A1(n278), .A2(n923), .A3(n921), .ZN(n27877) );
  INV_X1 U8 ( .A(n3722), .ZN(n27978) );
  AND3_X1 U9 ( .A1(n4064), .A2(n2013), .A3(n4063), .ZN(n25914) );
  OR2_X1 U14 ( .A1(n23051), .A2(n24341), .ZN(n1223) );
  INV_X1 U16 ( .A(n24758), .ZN(n171) );
  OAI21_X2 U18 ( .B1(n23019), .B2(n23018), .A(n23017), .ZN(n24688) );
  OR2_X1 U22 ( .A1(n28460), .A2(n23078), .ZN(n23838) );
  OR2_X1 U25 ( .A1(n3940), .A2(n23825), .ZN(n4483) );
  OR2_X1 U29 ( .A1(n20858), .A2(n21159), .ZN(n14) );
  OR2_X1 U30 ( .A1(n20933), .A2(n20533), .ZN(n1342) );
  INV_X1 U32 ( .A(n21495), .ZN(n44) );
  AND2_X1 U33 ( .A1(n21481), .A2(n21483), .ZN(n20368) );
  NOR2_X1 U34 ( .A1(n21481), .A2(n21574), .ZN(n20849) );
  INV_X1 U35 ( .A(n21497), .ZN(n7) );
  BUF_X1 U39 ( .A(n20225), .Z(n20503) );
  OR2_X1 U41 ( .A1(n17849), .A2(n18137), .ZN(n18142) );
  OAI211_X1 U42 ( .C1(n18506), .C2(n18216), .A(n28763), .B(n18217), .ZN(n2045)
         );
  OR2_X1 U43 ( .A1(n18252), .A2(n17771), .ZN(n3086) );
  AND2_X1 U44 ( .A1(n18101), .A2(n18449), .ZN(n106) );
  OR2_X1 U48 ( .A1(n5200), .A2(n18173), .ZN(n1137) );
  OR2_X1 U49 ( .A1(n18324), .A2(n18263), .ZN(n18323) );
  AND2_X1 U50 ( .A1(n18306), .A2(n17679), .ZN(n17680) );
  INV_X1 U52 ( .A(n18465), .ZN(n145) );
  INV_X1 U53 ( .A(n18270), .ZN(n48) );
  AND3_X1 U54 ( .A1(n17187), .A2(n17186), .A3(n17185), .ZN(n18122) );
  OR2_X1 U57 ( .A1(n18507), .A2(n29496), .ZN(n18074) );
  INV_X1 U58 ( .A(n18213), .ZN(n511) );
  OR2_X1 U62 ( .A1(n16917), .A2(n16916), .ZN(n186) );
  OAI22_X1 U64 ( .A1(n17315), .A2(n17316), .B1(n4220), .B2(n17562), .ZN(n792)
         );
  NOR2_X1 U65 ( .A1(n17528), .A2(n17524), .ZN(n17182) );
  OR2_X1 U66 ( .A1(n16811), .A2(n16812), .ZN(n3302) );
  XNOR2_X1 U68 ( .A(n15068), .B(n15067), .ZN(n17435) );
  XNOR2_X1 U69 ( .A(n16256), .B(n15977), .ZN(n16627) );
  OR2_X1 U70 ( .A1(n15399), .A2(n13638), .ZN(n6856) );
  OR2_X1 U73 ( .A1(n15370), .A2(n15009), .ZN(n3783) );
  OR2_X1 U74 ( .A1(n5049), .A2(n15274), .ZN(n217) );
  AND2_X1 U75 ( .A1(n15046), .A2(n15342), .ZN(n15229) );
  OR2_X1 U81 ( .A1(n13766), .A2(n14481), .ZN(n140) );
  OR2_X1 U83 ( .A1(n14037), .A2(n60), .ZN(n13722) );
  AND2_X1 U84 ( .A1(n29565), .A2(n29306), .ZN(n12121) );
  OR2_X1 U85 ( .A1(n14365), .A2(n14091), .ZN(n731) );
  NOR2_X1 U87 ( .A1(n12887), .A2(n1841), .ZN(n245) );
  INV_X1 U88 ( .A(n14452), .ZN(n190) );
  INV_X1 U89 ( .A(n13589), .ZN(n58) );
  INV_X1 U90 ( .A(n29089), .ZN(n60) );
  OAI21_X1 U92 ( .B1(n30), .B2(n14400), .A(n29), .ZN(n2112) );
  INV_X1 U93 ( .A(n14398), .ZN(n30) );
  XNOR2_X1 U94 ( .A(n12606), .B(n12605), .ZN(n14292) );
  AND2_X1 U95 ( .A1(n11985), .A2(n11986), .ZN(n163) );
  NAND3_X1 U96 ( .A1(n11697), .A2(n11696), .A3(n11695), .ZN(n13484) );
  OR2_X1 U97 ( .A1(n10900), .A2(n919), .ZN(n172) );
  OAI211_X1 U98 ( .C1(n12297), .C2(n12296), .A(n12295), .B(n12294), .ZN(n13121) );
  OR2_X1 U99 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  AND3_X1 U103 ( .A1(n4902), .A2(n11172), .A3(n11171), .ZN(n11194) );
  OR2_X1 U105 ( .A1(n4789), .A2(n4790), .ZN(n11417) );
  AND2_X1 U106 ( .A1(n10963), .A2(n10956), .ZN(n9859) );
  OAI21_X1 U108 ( .B1(n11289), .B2(n11290), .A(n11077), .ZN(n5717) );
  INV_X1 U111 ( .A(n11113), .ZN(n242) );
  AND3_X1 U119 ( .A1(n1417), .A2(n1418), .A3(n7574), .ZN(n15) );
  OR2_X1 U120 ( .A1(n8360), .A2(n9037), .ZN(n6189) );
  INV_X1 U121 ( .A(n9374), .ZN(n11) );
  BUF_X1 U122 ( .A(n7679), .Z(n9210) );
  INV_X1 U123 ( .A(n9122), .ZN(n81) );
  AND3_X1 U127 ( .A1(n5493), .A2(n7780), .A3(n7779), .ZN(n8427) );
  OAI211_X1 U128 ( .C1(n7425), .C2(n7426), .A(n3929), .B(n1358), .ZN(n8740) );
  INV_X1 U129 ( .A(n8215), .ZN(n8212) );
  BUF_X1 U130 ( .A(n8221), .Z(n7827) );
  AND2_X1 U137 ( .A1(n29621), .A2(n26125), .ZN(n26860) );
  OR2_X1 U140 ( .A1(n1807), .A2(n29043), .ZN(n24418) );
  AOI22_X1 U142 ( .A1(n21426), .A2(n5827), .B1(n20129), .B2(n6937), .ZN(n5622)
         );
  AND2_X1 U146 ( .A1(n26917), .A2(n26172), .ZN(n26553) );
  BUF_X1 U147 ( .A(n14630), .Z(n15394) );
  OR2_X1 U149 ( .A1(n11282), .A2(n10518), .ZN(n10519) );
  AND2_X1 U150 ( .A1(n20299), .A2(n20443), .ZN(n128) );
  AND2_X1 U153 ( .A1(n17336), .A2(n17155), .ZN(n15581) );
  OR2_X1 U154 ( .A1(n17336), .A2(n17155), .ZN(n241) );
  AND2_X1 U158 ( .A1(n27711), .A2(n27724), .ZN(n27694) );
  AND2_X1 U160 ( .A1(n20547), .A2(n20546), .ZN(n19960) );
  OR2_X1 U165 ( .A1(n24347), .A2(n24436), .ZN(n24442) );
  OAI21_X1 U166 ( .B1(n29090), .B2(n85), .A(n84), .ZN(n27658) );
  OR2_X1 U167 ( .A1(n11195), .A2(n11194), .ZN(n179) );
  XNOR2_X1 U171 ( .A(n18568), .B(n18567), .ZN(n20077) );
  INV_X1 U172 ( .A(n3315), .ZN(n184) );
  OR2_X1 U173 ( .A1(n15098), .A2(n3315), .ZN(n183) );
  OR3_X1 U175 ( .A1(n395), .A2(n26880), .A3(n27300), .ZN(n26882) );
  OR2_X1 U176 ( .A1(n26166), .A2(n29054), .ZN(n4399) );
  OR2_X1 U177 ( .A1(n26410), .A2(n26797), .ZN(n56) );
  AND2_X1 U179 ( .A1(n23403), .A2(n23214), .ZN(n23749) );
  OR2_X1 U181 ( .A1(n15402), .A2(n13639), .ZN(n14896) );
  AOI21_X1 U185 ( .B1(n9202), .B2(n9199), .A(n231), .ZN(n2196) );
  OR2_X1 U188 ( .A1(n2794), .A2(n27739), .ZN(n1216) );
  OR2_X1 U190 ( .A1(n26965), .A2(n27497), .ZN(n225) );
  OAI21_X1 U191 ( .B1(n17997), .B2(n17883), .A(n3283), .ZN(n2468) );
  OR2_X1 U193 ( .A1(n1533), .A2(n25628), .ZN(n1532) );
  OR3_X1 U195 ( .A1(n28567), .A2(n2823), .A3(n24020), .ZN(n275) );
  BUF_X1 U196 ( .A(n27407), .Z(n342) );
  OAI21_X1 U199 ( .B1(n22970), .B2(n22969), .A(n22968), .ZN(n26023) );
  BUF_X1 U204 ( .A(n14358), .Z(n14272) );
  OAI211_X1 U205 ( .C1(n487), .C2(n28418), .A(n23838), .B(n23837), .ZN(n1162)
         );
  OR2_X1 U206 ( .A1(n29057), .A2(n29647), .ZN(n17693) );
  NAND3_X1 U209 ( .A1(n24447), .A2(n24756), .A3(n24218), .ZN(n24219) );
  AND2_X2 U210 ( .A1(n23561), .A2(n23560), .ZN(n24447) );
  NOR2_X1 U211 ( .A1(n14392), .A2(n1), .ZN(n2207) );
  INV_X1 U212 ( .A(n14391), .ZN(n1) );
  NAND2_X1 U213 ( .A1(n6048), .A2(n15284), .ZN(n14391) );
  NAND2_X1 U215 ( .A1(n28762), .A2(n3784), .ZN(n2) );
  NAND2_X1 U220 ( .A1(n9), .A2(n6), .ZN(n19832) );
  NAND2_X1 U221 ( .A1(n8), .A2(n7), .ZN(n6) );
  NAND2_X1 U222 ( .A1(n28789), .A2(n20865), .ZN(n8) );
  NAND2_X1 U223 ( .A1(n19830), .A2(n21497), .ZN(n9) );
  NAND3_X2 U237 ( .A1(n6218), .A2(n19900), .A3(n6219), .ZN(n3838) );
  OR2_X1 U239 ( .A1(n11921), .A2(n11853), .ZN(n3521) );
  NAND2_X1 U242 ( .A1(n12), .A2(n10), .ZN(n8571) );
  NAND2_X1 U243 ( .A1(n9370), .A2(n11), .ZN(n10) );
  NAND2_X1 U244 ( .A1(n8569), .A2(n8929), .ZN(n9370) );
  NAND2_X1 U245 ( .A1(n9373), .A2(n9374), .ZN(n12) );
  NAND3_X1 U246 ( .A1(n24123), .A2(n24125), .A3(n24124), .ZN(n153) );
  NAND3_X1 U250 ( .A1(n3119), .A2(n21161), .A3(n13), .ZN(n22656) );
  NAND2_X1 U253 ( .A1(n8208), .A2(n7700), .ZN(n7423) );
  NAND2_X1 U254 ( .A1(n3579), .A2(n3581), .ZN(n888) );
  BUF_X1 U257 ( .A(n22829), .Z(n355) );
  XNOR2_X1 U258 ( .A(n9673), .B(n4601), .ZN(n11163) );
  NAND3_X1 U267 ( .A1(n16), .A2(n17848), .A3(n3264), .ZN(n6443) );
  NAND2_X1 U268 ( .A1(n2811), .A2(n17847), .ZN(n16) );
  NAND2_X1 U275 ( .A1(n6829), .A2(n16974), .ZN(n17717) );
  NAND2_X1 U276 ( .A1(n18270), .A2(n18511), .ZN(n1124) );
  NAND2_X1 U277 ( .A1(n29647), .A2(n18508), .ZN(n18270) );
  NAND3_X1 U278 ( .A1(n7871), .A2(n7053), .A3(n7960), .ZN(n7055) );
  NAND2_X1 U280 ( .A1(n6679), .A2(n12050), .ZN(n6678) );
  NAND3_X1 U284 ( .A1(n19), .A2(n12240), .A3(n4617), .ZN(n4616) );
  NAND2_X1 U285 ( .A1(n12159), .A2(n11969), .ZN(n19) );
  AND4_X2 U291 ( .A1(n5502), .A2(n5504), .A3(n24627), .A4(n24626), .ZN(n27025)
         );
  NAND2_X1 U295 ( .A1(n22), .A2(n11185), .ZN(n11327) );
  NAND3_X1 U299 ( .A1(n18933), .A2(n21286), .A3(n21291), .ZN(n24) );
  NAND2_X1 U300 ( .A1(n21704), .A2(n21277), .ZN(n21374) );
  OR2_X1 U301 ( .A1(n8258), .A2(n28615), .ZN(n7468) );
  NAND2_X1 U305 ( .A1(n8608), .A2(n8320), .ZN(n8747) );
  OR2_X1 U306 ( .A1(n702), .A2(n20160), .ZN(n273) );
  NOR2_X2 U308 ( .A1(n6824), .A2(n25422), .ZN(n27442) );
  NAND2_X1 U310 ( .A1(n25), .A2(n11470), .ZN(n12955) );
  NAND3_X1 U314 ( .A1(n14466), .A2(n4840), .A3(n13678), .ZN(n13680) );
  AND3_X2 U315 ( .A1(n1946), .A2(n5437), .A3(n5435), .ZN(n21497) );
  OR2_X1 U316 ( .A1(n10726), .A2(n10929), .ZN(n10933) );
  AOI21_X1 U317 ( .B1(n23519), .B2(n21058), .A(n23516), .ZN(n21059) );
  NAND2_X1 U318 ( .A1(n23682), .A2(n29544), .ZN(n23519) );
  NAND2_X1 U319 ( .A1(n17201), .A2(n17203), .ZN(n2741) );
  AND2_X1 U320 ( .A1(n19054), .A2(n20178), .ZN(n20055) );
  NAND2_X1 U324 ( .A1(n14400), .A2(n14399), .ZN(n29) );
  NAND3_X1 U325 ( .A1(n2890), .A2(n8849), .A3(n8850), .ZN(n8854) );
  AND2_X2 U326 ( .A1(n7538), .A2(n7539), .ZN(n9060) );
  NAND2_X1 U327 ( .A1(n17430), .A2(n31), .ZN(n18398) );
  NAND3_X1 U329 ( .A1(n5025), .A2(n14897), .A3(n14896), .ZN(n14898) );
  NAND2_X1 U331 ( .A1(n5658), .A2(n21495), .ZN(n5657) );
  XNOR2_X2 U332 ( .A(n7117), .B(Key[8]), .ZN(n7164) );
  NAND2_X1 U333 ( .A1(n35), .A2(n32), .ZN(n4259) );
  NAND2_X1 U334 ( .A1(n34), .A2(n28171), .ZN(n32) );
  NAND2_X1 U336 ( .A1(n5847), .A2(n13583), .ZN(n34) );
  NAND2_X1 U337 ( .A1(n4260), .A2(n13730), .ZN(n35) );
  NAND3_X1 U338 ( .A1(n3167), .A2(n7771), .A3(n7770), .ZN(n7772) );
  NAND3_X1 U339 ( .A1(n24125), .A2(n24705), .A3(n24338), .ZN(n5836) );
  AND2_X2 U341 ( .A1(n5898), .A2(n5897), .ZN(n21982) );
  INV_X1 U343 ( .A(n14738), .ZN(n36) );
  NAND2_X1 U344 ( .A1(n7716), .A2(n7717), .ZN(n7720) );
  NAND3_X1 U346 ( .A1(n11321), .A2(n11322), .A3(n11181), .ZN(n37) );
  NAND2_X1 U347 ( .A1(n11324), .A2(n29316), .ZN(n39) );
  NAND2_X1 U352 ( .A1(n3753), .A2(n18286), .ZN(n40) );
  NAND3_X1 U354 ( .A1(n8998), .A2(n9435), .A3(n8996), .ZN(n41) );
  NAND2_X1 U355 ( .A1(n42), .A2(n16942), .ZN(n6643) );
  NAND3_X1 U359 ( .A1(n11063), .A2(n1851), .A3(n10641), .ZN(n2084) );
  NAND2_X1 U361 ( .A1(n28789), .A2(n44), .ZN(n43) );
  INV_X1 U364 ( .A(n7266), .ZN(n7709) );
  XNOR2_X1 U365 ( .A(n16051), .B(n16620), .ZN(n16196) );
  NOR2_X1 U366 ( .A1(n20293), .A2(n19815), .ZN(n20122) );
  NAND3_X1 U368 ( .A1(n3175), .A2(n6352), .A3(n3488), .ZN(n14696) );
  OR2_X1 U369 ( .A1(n18449), .A2(n18451), .ZN(n1026) );
  NAND3_X1 U373 ( .A1(n4130), .A2(n27031), .A3(n4132), .ZN(n3611) );
  NAND2_X1 U374 ( .A1(n19060), .A2(n20221), .ZN(n19062) );
  NAND2_X1 U375 ( .A1(n29587), .A2(n20222), .ZN(n19060) );
  NAND2_X1 U377 ( .A1(n48), .A2(n18271), .ZN(n46) );
  MUX2_X1 U380 ( .A(n11708), .B(n11648), .S(n11417), .Z(n11408) );
  AND2_X1 U381 ( .A1(n23968), .A2(n24209), .ZN(n23116) );
  AND2_X1 U388 ( .A1(n12321), .A2(n12050), .ZN(n77) );
  NAND2_X1 U393 ( .A1(n50), .A2(n1048), .ZN(n12504) );
  NAND2_X1 U394 ( .A1(n11647), .A2(n743), .ZN(n50) );
  NOR2_X2 U395 ( .A1(n162), .A2(n51), .ZN(n24949) );
  NAND2_X1 U397 ( .A1(n24475), .A2(n53), .ZN(n52) );
  INV_X1 U398 ( .A(n6348), .ZN(n53) );
  NAND2_X1 U399 ( .A1(n23841), .A2(n6348), .ZN(n54) );
  OR2_X2 U400 ( .A1(n10831), .A2(n10832), .ZN(n11648) );
  OAI21_X1 U402 ( .B1(n14662), .B2(n14663), .A(n55), .ZN(n14665) );
  INV_X1 U403 ( .A(n14660), .ZN(n55) );
  NAND2_X1 U405 ( .A1(n10808), .A2(n10544), .ZN(n10805) );
  NAND3_X1 U406 ( .A1(n461), .A2(n28415), .A3(n25008), .ZN(n4141) );
  MUX2_X2 U411 ( .A(n9477), .B(n13082), .S(n13081), .Z(n13051) );
  NAND2_X1 U414 ( .A1(n1717), .A2(n3833), .ZN(n1716) );
  OR2_X2 U418 ( .A1(n2832), .A2(n7589), .ZN(n7875) );
  OAI211_X1 U421 ( .C1(n13720), .C2(n60), .A(n59), .B(n58), .ZN(n57) );
  OAI21_X1 U425 ( .B1(n6904), .B2(n21471), .A(n21232), .ZN(n21233) );
  INV_X1 U428 ( .A(n8187), .ZN(n8936) );
  NAND2_X1 U433 ( .A1(n28894), .A2(n20616), .ZN(n20256) );
  NAND3_X1 U439 ( .A1(n9188), .A2(n9185), .A3(n9184), .ZN(n887) );
  NAND2_X1 U440 ( .A1(n9012), .A2(n8910), .ZN(n8482) );
  NAND3_X2 U443 ( .A1(n2676), .A2(n7412), .A3(n7414), .ZN(n2677) );
  NAND2_X1 U446 ( .A1(n18171), .A2(n17780), .ZN(n1563) );
  BUF_X1 U448 ( .A(n27271), .Z(n27923) );
  INV_X1 U449 ( .A(n21467), .ZN(n19793) );
  NAND2_X1 U450 ( .A1(n5953), .A2(n21113), .ZN(n21467) );
  NAND2_X1 U452 ( .A1(n1436), .A2(n17447), .ZN(n1468) );
  OR2_X1 U455 ( .A1(n28796), .A2(n23408), .ZN(n23748) );
  NAND2_X1 U459 ( .A1(n14122), .A2(n14366), .ZN(n14093) );
  OAI21_X1 U460 ( .B1(n28800), .B2(n17464), .A(n63), .ZN(n5251) );
  NAND2_X1 U461 ( .A1(n17466), .A2(n4246), .ZN(n63) );
  NAND3_X2 U463 ( .A1(n64), .A2(n13765), .A3(n13766), .ZN(n15207) );
  NAND2_X1 U464 ( .A1(n6744), .A2(n13947), .ZN(n64) );
  NAND3_X1 U467 ( .A1(n66), .A2(n16152), .A3(n519), .ZN(n2457) );
  OAI21_X1 U470 ( .B1(n23192), .B2(n23193), .A(n28764), .ZN(n3158) );
  XNOR2_X2 U475 ( .A(n15969), .B(n15970), .ZN(n17277) );
  OAI211_X2 U476 ( .C1(n14060), .C2(n4185), .A(n4184), .B(n4181), .ZN(n16232)
         );
  AND2_X1 U477 ( .A1(n11033), .A2(n11248), .ZN(n10525) );
  NAND2_X1 U478 ( .A1(n69), .A2(n18180), .ZN(n17792) );
  NAND2_X1 U479 ( .A1(n17788), .A2(n17789), .ZN(n69) );
  NAND2_X1 U480 ( .A1(n4477), .A2(n4476), .ZN(n17789) );
  NAND2_X1 U482 ( .A1(n6399), .A2(n6400), .ZN(n20876) );
  NAND2_X1 U484 ( .A1(n4446), .A2(n12208), .ZN(n71) );
  NAND2_X1 U486 ( .A1(n6117), .A2(n20914), .ZN(n73) );
  AND2_X2 U490 ( .A1(n76), .A2(n75), .ZN(n21291) );
  NAND2_X1 U491 ( .A1(n18891), .A2(n18892), .ZN(n75) );
  NAND2_X1 U492 ( .A1(n5424), .A2(n3911), .ZN(n76) );
  NAND2_X1 U493 ( .A1(n566), .A2(n77), .ZN(n11771) );
  NOR2_X2 U497 ( .A1(n17682), .A2(n17681), .ZN(n19637) );
  MUX2_X2 U503 ( .A(n25986), .B(n25985), .S(n27013), .Z(n28019) );
  NAND2_X1 U504 ( .A1(n80), .A2(n79), .ZN(n6172) );
  NAND2_X1 U505 ( .A1(n9125), .A2(n9122), .ZN(n79) );
  NAND2_X1 U506 ( .A1(n1651), .A2(n1793), .ZN(n80) );
  NAND2_X1 U510 ( .A1(n15393), .A2(n15392), .ZN(n82) );
  INV_X1 U513 ( .A(n18603), .ZN(n18604) );
  NAND3_X1 U514 ( .A1(n28142), .A2(n18600), .A3(n17989), .ZN(n18603) );
  NOR2_X1 U515 ( .A1(n28522), .A2(n24804), .ZN(n24805) );
  NAND2_X1 U518 ( .A1(n400), .A2(n27701), .ZN(n27163) );
  NAND2_X1 U520 ( .A1(n29091), .A2(n27672), .ZN(n84) );
  BUF_X1 U521 ( .A(n27728), .Z(n1826) );
  NOR2_X1 U522 ( .A1(n17347), .A2(n29632), .ZN(n16949) );
  MUX2_X1 U532 ( .A(n9229), .B(n9232), .S(n9233), .Z(n7000) );
  NAND2_X1 U535 ( .A1(n6961), .A2(n6960), .ZN(n87) );
  OAI21_X1 U538 ( .B1(n6061), .B2(n14792), .A(n14970), .ZN(n88) );
  INV_X1 U539 ( .A(n12517), .ZN(n12077) );
  MUX2_X1 U540 ( .A(n12271), .B(n12578), .S(n12517), .Z(n11567) );
  NOR2_X2 U541 ( .A1(n11098), .A2(n11097), .ZN(n12517) );
  NAND2_X1 U544 ( .A1(n432), .A2(n89), .ZN(n6165) );
  NOR2_X1 U545 ( .A1(n5258), .A2(n10431), .ZN(n89) );
  INV_X1 U547 ( .A(n28105), .ZN(n91) );
  NAND3_X1 U548 ( .A1(n13944), .A2(n13941), .A3(n15025), .ZN(n13950) );
  OAI21_X1 U549 ( .B1(n26236), .B2(n26753), .A(n92), .ZN(n26756) );
  NAND2_X1 U550 ( .A1(n26753), .A2(n28575), .ZN(n92) );
  BUF_X1 U552 ( .A(n15165), .Z(n1850) );
  NAND3_X1 U555 ( .A1(n13651), .A2(n14303), .A3(n13817), .ZN(n13650) );
  NAND2_X1 U557 ( .A1(n27124), .A2(n27190), .ZN(n26336) );
  OR2_X1 U559 ( .A1(n26338), .A2(n26339), .ZN(n96) );
  NAND3_X1 U561 ( .A1(n19899), .A2(n20645), .A3(n19927), .ZN(n6218) );
  NAND3_X1 U568 ( .A1(n7493), .A2(n7491), .A3(n28219), .ZN(n9313) );
  AND3_X2 U572 ( .A1(n983), .A2(n3736), .A3(n7459), .ZN(n8320) );
  XNOR2_X2 U575 ( .A(n100), .B(n2113), .ZN(n14400) );
  XNOR2_X1 U576 ( .A(n12448), .B(n12449), .ZN(n100) );
  NAND3_X2 U582 ( .A1(n101), .A2(n1602), .A3(n1601), .ZN(n19452) );
  NAND2_X1 U583 ( .A1(n18088), .A2(n527), .ZN(n101) );
  INV_X1 U584 ( .A(n20560), .ZN(n20561) );
  NAND2_X1 U585 ( .A1(n19849), .A2(n20208), .ZN(n20560) );
  NAND3_X1 U586 ( .A1(n23182), .A2(n23181), .A3(n28765), .ZN(n24241) );
  NAND2_X1 U589 ( .A1(n948), .A2(n4913), .ZN(n951) );
  NAND3_X1 U591 ( .A1(n24016), .A2(n4639), .A3(n5799), .ZN(n6215) );
  AND4_X2 U594 ( .A1(n11286), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n12176) );
  NAND2_X1 U598 ( .A1(n15271), .A2(n5948), .ZN(n15956) );
  AND2_X1 U599 ( .A1(n17564), .A2(n17772), .ZN(n17577) );
  NAND3_X1 U602 ( .A1(n104), .A2(n5623), .A3(n4732), .ZN(n17329) );
  NAND2_X1 U603 ( .A1(n18138), .A2(n18137), .ZN(n104) );
  NAND3_X1 U605 ( .A1(n1798), .A2(n1799), .A3(n6500), .ZN(n18193) );
  OAI21_X2 U606 ( .B1(n18751), .B2(n20087), .A(n18750), .ZN(n21000) );
  NAND3_X1 U607 ( .A1(n8701), .A2(n8703), .A3(n105), .ZN(n10231) );
  OAI21_X1 U610 ( .B1(n20793), .B2(n107), .A(n21198), .ZN(n20796) );
  NOR2_X1 U611 ( .A1(n21512), .A2(n21199), .ZN(n107) );
  NAND2_X1 U613 ( .A1(n17861), .A2(n18511), .ZN(n5228) );
  NAND2_X1 U614 ( .A1(n10838), .A2(n10835), .ZN(n10836) );
  XNOR2_X1 U625 ( .A(n109), .B(n2509), .ZN(Ciphertext[140]) );
  NAND3_X1 U626 ( .A1(n26524), .A2(n26525), .A3(n26523), .ZN(n109) );
  XNOR2_X2 U632 ( .A(n16562), .B(n16561), .ZN(n17106) );
  XNOR2_X2 U645 ( .A(n9486), .B(n9485), .ZN(n11318) );
  NOR2_X1 U648 ( .A1(n29595), .A2(n18423), .ZN(n111) );
  INV_X1 U649 ( .A(n4805), .ZN(n112) );
  NAND2_X1 U650 ( .A1(n17822), .A2(n29594), .ZN(n113) );
  NOR3_X1 U651 ( .A1(n21692), .A2(n21348), .A3(n6314), .ZN(n20963) );
  XNOR2_X1 U653 ( .A(n22338), .B(n22717), .ZN(n22519) );
  NAND2_X2 U656 ( .A1(n1207), .A2(n8901), .ZN(n10328) );
  NAND3_X1 U658 ( .A1(n1651), .A2(n8897), .A3(n29304), .ZN(n1714) );
  OAI22_X1 U660 ( .A1(n7716), .A2(n8134), .B1(n7718), .B2(n29646), .ZN(n2506)
         );
  MUX2_X2 U662 ( .A(n11448), .B(n11447), .S(n12361), .Z(n13166) );
  NAND2_X1 U663 ( .A1(n12115), .A2(n6281), .ZN(n12113) );
  NAND2_X1 U667 ( .A1(n8861), .A2(n4585), .ZN(n4584) );
  NOR2_X1 U668 ( .A1(n8378), .A2(n9075), .ZN(n8861) );
  NAND3_X1 U671 ( .A1(n10718), .A2(n11137), .A3(n11142), .ZN(n10107) );
  NOR2_X1 U672 ( .A1(n27615), .A2(n114), .ZN(n27623) );
  NAND2_X1 U674 ( .A1(n479), .A2(n23419), .ZN(n22806) );
  NAND2_X1 U679 ( .A1(n13642), .A2(n13641), .ZN(n16322) );
  NAND2_X1 U681 ( .A1(n8536), .A2(n8734), .ZN(n8542) );
  NAND2_X1 U682 ( .A1(n3558), .A2(n12058), .ZN(n11295) );
  NAND3_X1 U689 ( .A1(n5552), .A2(n23222), .A3(n5553), .ZN(n24538) );
  OAI211_X1 U698 ( .C1(n27746), .C2(n27736), .A(n119), .B(n118), .ZN(n27738)
         );
  NAND2_X1 U699 ( .A1(n27733), .A2(n27749), .ZN(n118) );
  NAND2_X1 U700 ( .A1(n27734), .A2(n27757), .ZN(n119) );
  NAND3_X1 U701 ( .A1(n8006), .A2(n120), .A3(n9099), .ZN(n8005) );
  NAND2_X1 U702 ( .A1(n9100), .A2(n8664), .ZN(n120) );
  NAND3_X1 U704 ( .A1(n8168), .A2(n8159), .A3(n8158), .ZN(n8164) );
  NAND2_X1 U705 ( .A1(n121), .A2(n14802), .ZN(n3287) );
  NAND2_X1 U706 ( .A1(n3506), .A2(n3507), .ZN(n121) );
  NAND3_X1 U709 ( .A1(n1181), .A2(n4681), .A3(n17275), .ZN(n4613) );
  BUF_X1 U710 ( .A(n7198), .Z(n7406) );
  NAND2_X1 U720 ( .A1(n10549), .A2(n10492), .ZN(n11112) );
  INV_X1 U722 ( .A(n18190), .ZN(n122) );
  INV_X1 U723 ( .A(n18188), .ZN(n123) );
  NAND2_X1 U726 ( .A1(n11609), .A2(n4404), .ZN(n125) );
  NAND2_X1 U732 ( .A1(n29321), .A2(n8024), .ZN(n8022) );
  NAND2_X1 U734 ( .A1(n21007), .A2(n4266), .ZN(n2343) );
  OAI22_X1 U736 ( .A1(n8708), .A2(n8876), .B1(n8710), .B2(n8709), .ZN(n127) );
  NAND2_X1 U737 ( .A1(n415), .A2(n128), .ZN(n6840) );
  NAND2_X1 U738 ( .A1(n7843), .A2(n8024), .ZN(n7010) );
  NAND3_X1 U739 ( .A1(n10453), .A2(n130), .A3(n287), .ZN(n6330) );
  INV_X1 U741 ( .A(n11881), .ZN(n130) );
  NAND3_X2 U743 ( .A1(n16552), .A2(n16551), .A3(n16553), .ZN(n18354) );
  NAND2_X1 U749 ( .A1(n24893), .A2(n24532), .ZN(n132) );
  NAND3_X1 U752 ( .A1(n9362), .A2(n10959), .A3(n10686), .ZN(n897) );
  NOR2_X1 U763 ( .A1(n6424), .A2(n23772), .ZN(n136) );
  NAND3_X1 U765 ( .A1(n6709), .A2(n26907), .A3(n6710), .ZN(n6708) );
  AND3_X2 U767 ( .A1(n3720), .A2(n6887), .A3(n6888), .ZN(n27457) );
  XNOR2_X1 U769 ( .A(n19331), .B(n19408), .ZN(n19119) );
  NOR2_X1 U771 ( .A1(n22967), .A2(n137), .ZN(n22968) );
  NOR2_X1 U772 ( .A1(n6686), .A2(n23127), .ZN(n137) );
  NAND2_X2 U776 ( .A1(n2620), .A2(n138), .ZN(n24347) );
  NAND2_X1 U780 ( .A1(n8574), .A2(n8579), .ZN(n8767) );
  NOR2_X2 U782 ( .A1(n13820), .A2(n13819), .ZN(n16366) );
  NAND2_X1 U784 ( .A1(n3089), .A2(n10916), .ZN(n139) );
  NAND3_X1 U786 ( .A1(n141), .A2(n12140), .A3(n140), .ZN(n15407) );
  NAND2_X1 U793 ( .A1(n21425), .A2(n5827), .ZN(n21086) );
  NAND2_X1 U798 ( .A1(n626), .A2(n8217), .ZN(n8215) );
  NAND2_X1 U799 ( .A1(n144), .A2(n143), .ZN(n5492) );
  AOI21_X1 U800 ( .B1(n18465), .B2(n6079), .A(n18471), .ZN(n143) );
  NAND2_X1 U801 ( .A1(n145), .A2(n17916), .ZN(n144) );
  OR2_X2 U802 ( .A1(n14588), .A2(n14587), .ZN(n16257) );
  NAND2_X1 U803 ( .A1(n148), .A2(n147), .ZN(n146) );
  NAND2_X1 U804 ( .A1(n24683), .A2(n23902), .ZN(n147) );
  INV_X1 U806 ( .A(n24683), .ZN(n149) );
  NAND2_X1 U807 ( .A1(n21564), .A2(n21563), .ZN(n21115) );
  NAND2_X1 U808 ( .A1(n20756), .A2(n21565), .ZN(n21563) );
  AOI21_X1 U810 ( .B1(n17002), .B2(n17276), .A(n17272), .ZN(n15981) );
  XNOR2_X1 U812 ( .A(n9577), .B(n9878), .ZN(n10123) );
  NAND2_X1 U814 ( .A1(n3230), .A2(n3231), .ZN(n27958) );
  AND2_X1 U822 ( .A1(n15060), .A2(n15360), .ZN(n15357) );
  NAND2_X1 U833 ( .A1(n6761), .A2(n1315), .ZN(n1314) );
  OR2_X2 U837 ( .A1(n8487), .A2(n8486), .ZN(n9125) );
  OR2_X1 U839 ( .A1(n14106), .A2(n14107), .ZN(n14235) );
  NAND2_X1 U843 ( .A1(n1003), .A2(n1004), .ZN(n1002) );
  AOI21_X1 U845 ( .B1(n208), .B2(n7943), .A(n29317), .ZN(n155) );
  AOI22_X2 U847 ( .A1(n17372), .A2(n17371), .B1(n17370), .B2(n17369), .ZN(
        n18404) );
  OR2_X1 U848 ( .A1(n14842), .A2(n14600), .ZN(n14071) );
  XNOR2_X1 U850 ( .A(n156), .B(n26590), .ZN(Ciphertext[48]) );
  NAND4_X1 U851 ( .A1(n5367), .A2(n5369), .A3(n26589), .A4(n26588), .ZN(n156)
         );
  NOR2_X1 U855 ( .A1(n23179), .A2(n157), .ZN(n23182) );
  NOR3_X1 U856 ( .A1(n1838), .A2(n23645), .A3(n23640), .ZN(n157) );
  NAND3_X1 U858 ( .A1(n5035), .A2(n25453), .A3(n29100), .ZN(n25470) );
  NAND2_X1 U859 ( .A1(n2418), .A2(n2420), .ZN(n9190) );
  OAI21_X1 U863 ( .B1(n21420), .B2(n20806), .A(n20805), .ZN(n20807) );
  NOR2_X1 U864 ( .A1(n5000), .A2(n20899), .ZN(n21420) );
  NAND2_X1 U865 ( .A1(n15464), .A2(n15160), .ZN(n785) );
  NAND2_X1 U867 ( .A1(n18478), .A2(n18304), .ZN(n18309) );
  BUF_X1 U871 ( .A(n10534), .Z(n10659) );
  NAND3_X1 U873 ( .A1(n14385), .A2(n14382), .A3(n14381), .ZN(n14383) );
  XNOR2_X1 U875 ( .A(n29580), .B(n19637), .ZN(n19430) );
  XNOR2_X1 U877 ( .A(n21789), .B(n22094), .ZN(n22689) );
  AND2_X2 U878 ( .A1(n20927), .A2(n4566), .ZN(n21789) );
  OAI21_X1 U887 ( .B1(n21163), .B2(n4148), .A(n21609), .ZN(n159) );
  NAND3_X1 U890 ( .A1(n24412), .A2(n24711), .A3(n24714), .ZN(n24413) );
  NAND2_X1 U893 ( .A1(n161), .A2(n20858), .ZN(n20530) );
  NAND2_X1 U894 ( .A1(n21157), .A2(n21159), .ZN(n161) );
  NAND2_X2 U898 ( .A1(n23015), .A2(n3743), .ZN(n24682) );
  AOI21_X2 U899 ( .B1(n20489), .B2(n20488), .A(n20487), .ZN(n21611) );
  NAND4_X2 U900 ( .A1(n2653), .A2(n5477), .A3(n2651), .A4(n2650), .ZN(n22633)
         );
  OR2_X2 U903 ( .A1(n6537), .A2(n23056), .ZN(n24713) );
  BUF_X1 U909 ( .A(n23010), .Z(n23011) );
  NAND2_X1 U913 ( .A1(n8930), .A2(n9147), .ZN(n8935) );
  XNOR2_X2 U914 ( .A(Key[1]), .B(Plaintext[1]), .ZN(n7890) );
  OR2_X1 U915 ( .A1(n8658), .A2(n8116), .ZN(n8497) );
  AND3_X2 U916 ( .A1(n23076), .A2(n1206), .A3(n3337), .ZN(n24374) );
  AOI22_X1 U918 ( .A1(n27001), .A2(n27045), .B1(n27003), .B2(n27002), .ZN(
        n27009) );
  NAND3_X1 U920 ( .A1(n5291), .A2(n23283), .A3(n6279), .ZN(n5293) );
  NAND2_X1 U921 ( .A1(n25423), .A2(n25424), .ZN(n25425) );
  OAI22_X1 U922 ( .A1(n23850), .A2(n24100), .B1(n23875), .B2(n24489), .ZN(n162) );
  NAND2_X1 U923 ( .A1(n377), .A2(n26560), .ZN(n948) );
  NAND3_X1 U924 ( .A1(n14065), .A2(n14064), .A3(n14325), .ZN(n3125) );
  NAND2_X1 U925 ( .A1(n694), .A2(n15335), .ZN(n693) );
  NAND2_X1 U926 ( .A1(n3415), .A2(n3416), .ZN(n17782) );
  XNOR2_X1 U936 ( .A(n165), .B(n8573), .ZN(n11199) );
  XNOR2_X1 U937 ( .A(n9668), .B(n9940), .ZN(n165) );
  NOR2_X1 U941 ( .A1(n6941), .A2(n167), .ZN(n23065) );
  NOR2_X1 U942 ( .A1(n23147), .A2(n1837), .ZN(n167) );
  NAND2_X1 U947 ( .A1(n14780), .A2(n15432), .ZN(n168) );
  NAND2_X1 U948 ( .A1(n14779), .A2(n15030), .ZN(n169) );
  AOI21_X1 U953 ( .B1(n170), .B2(n20618), .A(n20616), .ZN(n19923) );
  NAND2_X1 U954 ( .A1(n20617), .A2(n500), .ZN(n170) );
  NAND3_X1 U955 ( .A1(n171), .A2(n24760), .A3(n378), .ZN(n24763) );
  OAI211_X2 U958 ( .C1(n13908), .C2(n14051), .A(n5730), .B(n5386), .ZN(n13922)
         );
  XNOR2_X2 U959 ( .A(n16584), .B(n16583), .ZN(n17470) );
  BUF_X2 U960 ( .A(n10939), .Z(n11952) );
  OAI211_X2 U961 ( .C1(n19778), .C2(n19777), .A(n5075), .B(n5074), .ZN(n21140)
         );
  OAI22_X1 U969 ( .A1(n17823), .A2(n512), .B1(n4802), .B2(n17824), .ZN(n174)
         );
  AND3_X2 U978 ( .A1(n3535), .A2(n941), .A3(n939), .ZN(n18195) );
  AND2_X2 U979 ( .A1(n6120), .A2(n6121), .ZN(n25396) );
  NAND2_X1 U983 ( .A1(n1178), .A2(n2390), .ZN(n20298) );
  NAND3_X1 U986 ( .A1(n3291), .A2(n23601), .A3(n3292), .ZN(n24870) );
  NAND4_X2 U987 ( .A1(n175), .A2(n11015), .A3(n11016), .A4(n11018), .ZN(n12253) );
  NAND2_X1 U988 ( .A1(n1999), .A2(n6108), .ZN(n175) );
  MUX2_X1 U989 ( .A(n18215), .B(n18506), .S(n18213), .Z(n17728) );
  XNOR2_X2 U991 ( .A(n12910), .B(n12909), .ZN(n14287) );
  NAND2_X1 U992 ( .A1(n12402), .A2(n12407), .ZN(n11800) );
  OR2_X2 U993 ( .A1(n4462), .A2(n4461), .ZN(n12402) );
  INV_X1 U998 ( .A(n10250), .ZN(n9674) );
  OAI21_X2 U1003 ( .B1(n22448), .B2(n1740), .A(n178), .ZN(n24734) );
  NAND2_X1 U1004 ( .A1(n639), .A2(n23192), .ZN(n178) );
  NAND2_X1 U1005 ( .A1(n1040), .A2(n1082), .ZN(n19887) );
  NAND3_X1 U1006 ( .A1(n15448), .A2(n15322), .A3(n15446), .ZN(n15016) );
  INV_X1 U1007 ( .A(n8925), .ZN(n7403) );
  NAND2_X1 U1008 ( .A1(n9340), .A2(n6718), .ZN(n8925) );
  XNOR2_X1 U1009 ( .A(n18756), .B(n27225), .ZN(n18704) );
  BUF_X1 U1010 ( .A(n25120), .Z(n27182) );
  AOI21_X2 U1011 ( .B1(n26402), .B2(n26401), .A(n26400), .ZN(n27561) );
  XNOR2_X2 U1012 ( .A(n12643), .B(n12642), .ZN(n14451) );
  OAI21_X2 U1013 ( .B1(n15688), .B2(n2133), .A(n15687), .ZN(n18490) );
  OAI22_X1 U1014 ( .A1(n24118), .A2(n24435), .B1(n23886), .B2(n24119), .ZN(
        n24122) );
  NAND2_X1 U1015 ( .A1(n5837), .A2(n179), .ZN(n6850) );
  NAND2_X1 U1016 ( .A1(n4341), .A2(n11195), .ZN(n5837) );
  XNOR2_X1 U1020 ( .A(n16594), .B(n16595), .ZN(n180) );
  XNOR2_X1 U1021 ( .A(n181), .B(n9254), .ZN(n9608) );
  XNOR2_X1 U1022 ( .A(n9241), .B(n9242), .ZN(n181) );
  NAND2_X1 U1026 ( .A1(n24551), .A2(n24555), .ZN(n24550) );
  AND3_X2 U1028 ( .A1(n182), .A2(n3754), .A3(n26399), .ZN(n27203) );
  OAI21_X1 U1029 ( .B1(n25122), .B2(n25123), .A(n25034), .ZN(n182) );
  OAI21_X1 U1030 ( .B1(n15099), .B2(n14677), .A(n183), .ZN(n14682) );
  OAI211_X2 U1031 ( .C1(n24553), .C2(n24174), .A(n5510), .B(n5508), .ZN(n26083) );
  OAI21_X1 U1032 ( .B1(n14170), .B2(n14169), .A(n14167), .ZN(n4073) );
  NAND3_X1 U1038 ( .A1(n8492), .A2(n8630), .A3(n9100), .ZN(n8493) );
  NOR2_X2 U1039 ( .A1(n16929), .A2(n16930), .ZN(n19272) );
  OAI211_X1 U1040 ( .C1(n12159), .C2(n12241), .A(n187), .B(n12037), .ZN(n4615)
         );
  NAND2_X1 U1041 ( .A1(n188), .A2(n12241), .ZN(n187) );
  INV_X1 U1042 ( .A(n12244), .ZN(n188) );
  NAND2_X1 U1048 ( .A1(n191), .A2(n190), .ZN(n189) );
  NAND2_X1 U1049 ( .A1(n14176), .A2(n14177), .ZN(n191) );
  NAND2_X1 U1050 ( .A1(n14179), .A2(n14452), .ZN(n192) );
  NAND2_X1 U1052 ( .A1(n193), .A2(n18138), .ZN(n914) );
  NAND3_X1 U1055 ( .A1(n29086), .A2(n29559), .A3(n17101), .ZN(n17103) );
  NAND3_X1 U1056 ( .A1(n11114), .A2(n29627), .A3(n28205), .ZN(n2867) );
  NAND2_X2 U1057 ( .A1(n5739), .A2(n5740), .ZN(n5234) );
  NAND3_X2 U1059 ( .A1(n2405), .A2(n8306), .A3(n8307), .ZN(n8955) );
  NAND2_X1 U1062 ( .A1(n21230), .A2(n21408), .ZN(n195) );
  OAI22_X1 U1064 ( .A1(n17693), .A2(n18516), .B1(n18270), .B2(n418), .ZN(
        n17694) );
  NAND3_X2 U1066 ( .A1(n6915), .A2(n2915), .A3(n9038), .ZN(n10350) );
  AND3_X2 U1068 ( .A1(n866), .A2(n275), .A3(n865), .ZN(n25381) );
  NAND3_X1 U1071 ( .A1(n9027), .A2(n9031), .A3(n9028), .ZN(n9033) );
  NAND3_X1 U1074 ( .A1(n22084), .A2(n6099), .A3(n28428), .ZN(n6585) );
  NAND3_X1 U1075 ( .A1(n197), .A2(n4924), .A3(n4919), .ZN(n4918) );
  NAND2_X1 U1076 ( .A1(n27243), .A2(n27402), .ZN(n197) );
  NOR2_X1 U1078 ( .A1(n5697), .A2(n198), .ZN(n5696) );
  NOR2_X1 U1079 ( .A1(n199), .A2(n5530), .ZN(n198) );
  NAND2_X1 U1080 ( .A1(n201), .A2(n23301), .ZN(n199) );
  INV_X1 U1082 ( .A(n22686), .ZN(n201) );
  NOR2_X2 U1085 ( .A1(n202), .A2(n24355), .ZN(n25149) );
  OAI21_X1 U1086 ( .B1(n24353), .B2(n28416), .A(n24352), .ZN(n202) );
  NAND3_X1 U1089 ( .A1(n7010), .A2(n6299), .A3(n29106), .ZN(n7014) );
  NAND2_X1 U1092 ( .A1(n204), .A2(n7163), .ZN(n2692) );
  NOR2_X1 U1093 ( .A1(n614), .A2(n7770), .ZN(n204) );
  NAND2_X1 U1094 ( .A1(n7585), .A2(n7580), .ZN(n7074) );
  NAND3_X1 U1097 ( .A1(n17905), .A2(n3866), .A3(n17903), .ZN(n3864) );
  XNOR2_X2 U1099 ( .A(n6986), .B(Key[90]), .ZN(n7424) );
  NAND3_X1 U1102 ( .A1(n1338), .A2(n3817), .A3(n11033), .ZN(n1336) );
  AND3_X2 U1103 ( .A1(n19009), .A2(n19008), .A3(n19007), .ZN(n21287) );
  NAND2_X1 U1107 ( .A1(n29547), .A2(n18410), .ZN(n18027) );
  MUX2_X1 U1113 ( .A(n11990), .B(n10863), .S(n12512), .Z(n10117) );
  NAND2_X2 U1117 ( .A1(n23374), .A2(n205), .ZN(n25931) );
  OR2_X2 U1119 ( .A1(n7461), .A2(n7460), .ZN(n8605) );
  NAND2_X1 U1120 ( .A1(n207), .A2(n206), .ZN(n20596) );
  NAND2_X1 U1121 ( .A1(n21591), .A2(n21322), .ZN(n206) );
  NAND2_X1 U1122 ( .A1(n20575), .A2(n20889), .ZN(n207) );
  NAND2_X1 U1123 ( .A1(n8301), .A2(n7942), .ZN(n208) );
  NAND3_X1 U1127 ( .A1(n5233), .A2(n18393), .A3(n17766), .ZN(n5232) );
  NAND2_X1 U1129 ( .A1(n4266), .A2(n20698), .ZN(n19733) );
  OAI211_X1 U1133 ( .C1(n27858), .C2(n447), .A(n209), .B(n4533), .ZN(n4535) );
  INV_X1 U1134 ( .A(n210), .ZN(n209) );
  OAI22_X1 U1135 ( .A1(n26646), .A2(n29095), .B1(n27859), .B2(n27851), .ZN(
        n210) );
  OAI211_X1 U1136 ( .C1(n17463), .C2(n28800), .A(n528), .B(n17280), .ZN(n4286)
         );
  AOI22_X2 U1137 ( .A1(n18338), .A2(n18339), .B1(n18336), .B2(n18337), .ZN(
        n19384) );
  OAI22_X1 U1139 ( .A1(n212), .A2(n211), .B1(n17057), .B2(n17542), .ZN(n17059)
         );
  INV_X1 U1140 ( .A(n17055), .ZN(n211) );
  NAND2_X1 U1141 ( .A1(n17213), .A2(n15787), .ZN(n212) );
  NAND3_X1 U1144 ( .A1(n20628), .A2(n28186), .A3(n20623), .ZN(n6883) );
  NAND2_X1 U1145 ( .A1(n213), .A2(n3279), .ZN(n7646) );
  NAND2_X1 U1146 ( .A1(n251), .A2(n7985), .ZN(n213) );
  NAND2_X1 U1148 ( .A1(n4856), .A2(n7100), .ZN(n7761) );
  AND3_X2 U1151 ( .A1(n216), .A2(n1363), .A3(n215), .ZN(n18087) );
  NAND2_X1 U1152 ( .A1(n16823), .A2(n17710), .ZN(n215) );
  NAND2_X1 U1153 ( .A1(n1366), .A2(n1365), .ZN(n216) );
  OR2_X2 U1154 ( .A1(n5465), .A2(n11615), .ZN(n13450) );
  NAND2_X1 U1157 ( .A1(n1909), .A2(n8058), .ZN(n8352) );
  NAND3_X1 U1158 ( .A1(n7765), .A2(n4855), .A3(n7764), .ZN(n1909) );
  NAND4_X2 U1161 ( .A1(n11745), .A2(n12360), .A3(n11744), .A4(n11743), .ZN(
        n13039) );
  OR2_X1 U1166 ( .A1(n7909), .A2(n8290), .ZN(n2898) );
  NAND2_X1 U1171 ( .A1(n15400), .A2(n28518), .ZN(n13636) );
  OAI21_X1 U1172 ( .B1(n1285), .B2(n10681), .A(n10680), .ZN(n10682) );
  NAND2_X1 U1173 ( .A1(n1285), .A2(n28608), .ZN(n10680) );
  NAND2_X1 U1174 ( .A1(n16550), .A2(n16547), .ZN(n699) );
  XNOR2_X2 U1176 ( .A(n1756), .B(n1755), .ZN(n20511) );
  NAND2_X1 U1179 ( .A1(n1255), .A2(n14498), .ZN(n2488) );
  AND2_X2 U1182 ( .A1(n6527), .A2(n6531), .ZN(n22271) );
  NAND2_X1 U1184 ( .A1(n221), .A2(n220), .ZN(n219) );
  NAND2_X1 U1185 ( .A1(n4685), .A2(n5004), .ZN(n221) );
  AOI21_X1 U1186 ( .B1(n223), .B2(n15409), .A(n15108), .ZN(n3918) );
  INV_X1 U1187 ( .A(n3922), .ZN(n223) );
  BUF_X2 U1188 ( .A(n17687), .Z(n20941) );
  AND3_X2 U1195 ( .A1(n874), .A2(n1518), .A3(n1613), .ZN(n15668) );
  NAND3_X1 U1196 ( .A1(n1643), .A2(n29138), .A3(n6306), .ZN(n1306) );
  NAND2_X1 U1197 ( .A1(n26428), .A2(n26381), .ZN(n26429) );
  XNOR2_X2 U1198 ( .A(n7122), .B(Key[38]), .ZN(n8141) );
  NAND3_X1 U1206 ( .A1(n7827), .A2(n7825), .A3(n7824), .ZN(n7826) );
  NAND3_X1 U1208 ( .A1(n5604), .A2(n5605), .A3(n225), .ZN(n2380) );
  NAND2_X1 U1215 ( .A1(n226), .A2(n5956), .ZN(n1020) );
  NAND2_X1 U1216 ( .A1(n794), .A2(n13647), .ZN(n226) );
  OAI21_X1 U1218 ( .B1(n17210), .B2(n17824), .A(n227), .ZN(n5551) );
  NAND3_X2 U1223 ( .A1(n5960), .A2(n8528), .A3(n5959), .ZN(n9755) );
  NOR2_X1 U1227 ( .A1(n23083), .A2(n23082), .ZN(n1777) );
  NAND2_X1 U1232 ( .A1(n4484), .A2(n229), .ZN(n5080) );
  OAI21_X1 U1233 ( .B1(n23845), .B2(n23722), .A(n23721), .ZN(n229) );
  NAND3_X1 U1240 ( .A1(n7685), .A2(n7843), .A3(n7515), .ZN(n7519) );
  AND2_X1 U1241 ( .A1(n28451), .A2(n27244), .ZN(n27948) );
  INV_X1 U1244 ( .A(n4880), .ZN(n19283) );
  NAND2_X1 U1245 ( .A1(n1231), .A2(n1232), .ZN(n4880) );
  BUF_X1 U1246 ( .A(n8592), .Z(n8978) );
  NAND2_X1 U1247 ( .A1(n5389), .A2(n29481), .ZN(n5388) );
  INV_X1 U1249 ( .A(n15071), .ZN(n14639) );
  NAND4_X2 U1250 ( .A1(n12940), .A2(n12939), .A3(n12941), .A4(n6562), .ZN(
        n15071) );
  NAND3_X1 U1251 ( .A1(n6479), .A2(n11486), .A3(n4744), .ZN(n11306) );
  NAND3_X1 U1257 ( .A1(n12190), .A2(n2483), .A3(n11724), .ZN(n11723) );
  NAND2_X1 U1258 ( .A1(n232), .A2(n5148), .ZN(n5147) );
  NAND3_X1 U1259 ( .A1(n7868), .A2(n7173), .A3(n7867), .ZN(n232) );
  BUF_X1 U1260 ( .A(n7233), .Z(n7592) );
  NAND2_X1 U1261 ( .A1(n17939), .A2(n17601), .ZN(n17943) );
  OAI211_X2 U1262 ( .C1(n16151), .C2(n16853), .A(n16150), .B(n3587), .ZN(
        n17939) );
  NAND3_X1 U1266 ( .A1(n705), .A2(n706), .A3(n12167), .ZN(n233) );
  NAND2_X2 U1270 ( .A1(n4268), .A2(n4267), .ZN(n21253) );
  XNOR2_X2 U1272 ( .A(n6979), .B(Key[99]), .ZN(n7635) );
  AND2_X2 U1277 ( .A1(n1469), .A2(n1471), .ZN(n27340) );
  NAND3_X1 U1280 ( .A1(n8856), .A2(n8857), .A3(n28212), .ZN(n881) );
  OAI21_X1 U1282 ( .B1(n2549), .B2(n13877), .A(n235), .ZN(n2607) );
  NAND2_X1 U1283 ( .A1(n13877), .A2(n14402), .ZN(n235) );
  NAND2_X1 U1285 ( .A1(n237), .A2(n17435), .ZN(n4427) );
  OAI21_X1 U1287 ( .B1(n8428), .B2(n1909), .A(n238), .ZN(n8432) );
  AND2_X1 U1293 ( .A1(n21000), .A2(n20972), .ZN(n20968) );
  NAND2_X1 U1295 ( .A1(n16774), .A2(n17016), .ZN(n16865) );
  OAI211_X2 U1296 ( .C1(n7927), .C2(n8216), .A(n2556), .B(n7627), .ZN(n9200)
         );
  NAND4_X2 U1297 ( .A1(n16793), .A2(n16796), .A3(n16794), .A4(n16795), .ZN(
        n19549) );
  AOI22_X1 U1300 ( .A1(n28437), .A2(n27120), .B1(n26512), .B2(n402), .ZN(
        n27122) );
  OAI22_X1 U1302 ( .A1(n18749), .A2(n19755), .B1(n29114), .B2(n20040), .ZN(
        n18750) );
  NAND2_X1 U1303 ( .A1(n29104), .A2(n20090), .ZN(n19755) );
  NAND2_X1 U1304 ( .A1(n15125), .A2(n14998), .ZN(n13985) );
  NAND3_X2 U1311 ( .A1(n4619), .A2(n4620), .A3(n4622), .ZN(n16377) );
  NAND2_X1 U1318 ( .A1(n8926), .A2(n9131), .ZN(n240) );
  BUF_X2 U1319 ( .A(n26374), .Z(n26950) );
  NAND3_X1 U1327 ( .A1(n11291), .A2(n11077), .A3(n11076), .ZN(n4352) );
  NAND2_X1 U1332 ( .A1(n11115), .A2(n11114), .ZN(n243) );
  NAND4_X2 U1335 ( .A1(n8697), .A2(n8694), .A3(n8695), .A4(n8696), .ZN(n10232)
         );
  MUX2_X2 U1350 ( .A(n15524), .B(n15523), .S(n18478), .Z(n19495) );
  NAND3_X1 U1351 ( .A1(n29475), .A2(n6419), .A3(n5188), .ZN(n26317) );
  XNOR2_X2 U1352 ( .A(n4961), .B(n12918), .ZN(n14285) );
  NAND2_X1 U1355 ( .A1(n14761), .A2(n14762), .ZN(n14765) );
  OAI211_X2 U1356 ( .C1(n21129), .C2(n21497), .A(n21128), .B(n244), .ZN(n22409) );
  NAND3_X1 U1357 ( .A1(n21126), .A2(n21127), .A3(n21497), .ZN(n244) );
  NAND3_X1 U1360 ( .A1(n530), .A2(n29636), .A3(n17379), .ZN(n16876) );
  AOI21_X1 U1363 ( .B1(n28761), .B2(n28200), .A(n245), .ZN(n2295) );
  NAND3_X2 U1365 ( .A1(n248), .A2(n8423), .A3(n8424), .ZN(n12202) );
  OAI21_X1 U1368 ( .B1(n250), .B2(n8223), .A(n249), .ZN(n8226) );
  NAND2_X1 U1369 ( .A1(n8223), .A2(n8224), .ZN(n249) );
  INV_X1 U1370 ( .A(n8225), .ZN(n250) );
  OAI21_X1 U1371 ( .B1(n15102), .B2(n15105), .A(n14936), .ZN(n6022) );
  NAND2_X1 U1373 ( .A1(n5838), .A2(n11622), .ZN(n6705) );
  NAND3_X1 U1374 ( .A1(n4926), .A2(n4925), .A3(n26820), .ZN(n3263) );
  NAND2_X1 U1376 ( .A1(n7191), .A2(n7641), .ZN(n251) );
  OAI21_X1 U1379 ( .B1(n4100), .B2(n16911), .A(n252), .ZN(n15848) );
  NAND2_X1 U1380 ( .A1(n4099), .A2(n16911), .ZN(n252) );
  OR2_X1 U1382 ( .A1(n11330), .A2(n10821), .ZN(n5366) );
  OR2_X2 U1385 ( .A1(n6485), .A2(n5732), .ZN(n18353) );
  OR2_X2 U1386 ( .A1(n10845), .A2(n10846), .ZN(n4617) );
  XNOR2_X1 U1387 ( .A(n253), .B(n11575), .ZN(n11577) );
  OAI211_X1 U1395 ( .C1(n26603), .C2(n6859), .A(n2053), .B(n255), .ZN(n6858)
         );
  NAND2_X1 U1396 ( .A1(n28026), .A2(n28030), .ZN(n255) );
  NAND2_X1 U1401 ( .A1(n1599), .A2(n14471), .ZN(n1598) );
  NAND2_X1 U1403 ( .A1(n3914), .A2(n17197), .ZN(n18414) );
  AND2_X2 U1404 ( .A1(n2705), .A2(n2704), .ZN(n19511) );
  NAND2_X1 U1406 ( .A1(n19981), .A2(n29066), .ZN(n702) );
  MUX2_X2 U1408 ( .A(n25596), .B(n25595), .S(n29482), .Z(n28035) );
  XNOR2_X1 U1412 ( .A(n9754), .B(n9992), .ZN(n10376) );
  BUF_X1 U1414 ( .A(n26322), .Z(n26992) );
  NAND2_X1 U1417 ( .A1(n257), .A2(n24750), .ZN(n2880) );
  OAI21_X1 U1418 ( .B1(n24746), .B2(n28550), .A(n4980), .ZN(n257) );
  NAND2_X1 U1421 ( .A1(n1527), .A2(n8760), .ZN(n8759) );
  NAND3_X1 U1425 ( .A1(n15315), .A2(n15319), .A3(n15308), .ZN(n14855) );
  NAND2_X2 U1428 ( .A1(n649), .A2(n19979), .ZN(n4937) );
  NAND3_X2 U1429 ( .A1(n14857), .A2(n1067), .A3(n14858), .ZN(n16165) );
  NAND2_X1 U1430 ( .A1(n398), .A2(n27041), .ZN(n4487) );
  AOI22_X1 U1433 ( .A1(n27886), .A2(n27885), .B1(n27884), .B2(n27923), .ZN(
        n27888) );
  NOR2_X2 U1436 ( .A1(n15590), .A2(n15589), .ZN(n18292) );
  BUF_X1 U1439 ( .A(n15239), .Z(n15234) );
  NAND3_X1 U1440 ( .A1(n24531), .A2(n24894), .A3(n24530), .ZN(n24537) );
  OR2_X1 U1441 ( .A1(n7231), .A2(n441), .ZN(n7871) );
  OAI21_X1 U1443 ( .B1(n8899), .B2(n1793), .A(n610), .ZN(n1792) );
  OAI211_X1 U1444 ( .C1(n8908), .C2(n1770), .A(n9016), .B(n1769), .ZN(n1771)
         );
  OR2_X1 U1445 ( .A1(n8752), .A2(n9529), .ZN(n749) );
  NOR2_X1 U1446 ( .A1(n8908), .A2(n9014), .ZN(n8662) );
  AOI22_X1 U1447 ( .A1(n8092), .A2(n9047), .B1(n5945), .B2(n8091), .ZN(n9577)
         );
  XNOR2_X1 U1449 ( .A(n9749), .B(n748), .ZN(n9946) );
  AND2_X1 U1450 ( .A1(n6779), .A2(n11004), .ZN(n1380) );
  XNOR2_X1 U1451 ( .A(n1396), .B(n1397), .ZN(n11227) );
  XNOR2_X1 U1458 ( .A(n16131), .B(n15854), .ZN(n16267) );
  OR2_X1 U1459 ( .A1(n28775), .A2(n17374), .ZN(n4652) );
  AND2_X1 U1460 ( .A1(n18493), .A2(n28633), .ZN(n18495) );
  INV_X1 U1461 ( .A(n21047), .ZN(n21412) );
  AND2_X1 U1464 ( .A1(n23338), .A2(n29108), .ZN(n1263) );
  XNOR2_X1 U1465 ( .A(n271), .B(n22432), .ZN(n23469) );
  OR2_X1 U1467 ( .A1(n24765), .A2(n24767), .ZN(n3054) );
  OR2_X1 U1469 ( .A1(n6198), .A2(n630), .ZN(n1301) );
  XNOR2_X1 U1471 ( .A(n277), .B(n25212), .ZN(n26480) );
  OR2_X1 U1472 ( .A1(n26476), .A2(n26186), .ZN(n24204) );
  INV_X1 U1474 ( .A(n29538), .ZN(n27372) );
  AND3_X1 U1475 ( .A1(n631), .A2(n8270), .A3(n7485), .ZN(n258) );
  XOR2_X1 U1476 ( .A(n16603), .B(n16476), .Z(n259) );
  XOR2_X1 U1477 ( .A(n9505), .B(n653), .Z(n260) );
  AND3_X1 U1478 ( .A1(n7765), .A2(n4855), .A3(n7764), .ZN(n261) );
  BUF_X1 U1479 ( .A(n10793), .Z(n12155) );
  BUF_X1 U1481 ( .A(n17206), .Z(n18129) );
  XNOR2_X1 U1482 ( .A(n25223), .B(n25222), .ZN(n26727) );
  AND3_X1 U1484 ( .A1(n11069), .A2(n1851), .A3(n11243), .ZN(n262) );
  NAND2_X2 U1485 ( .A1(n5089), .A2(n10115), .ZN(n12507) );
  AND2_X2 U1486 ( .A1(n3941), .A2(n3942), .ZN(n3946) );
  OR2_X1 U1489 ( .A1(n13310), .A2(n13309), .ZN(n263) );
  AND2_X1 U1494 ( .A1(n14144), .A2(n2974), .ZN(n265) );
  XOR2_X1 U1495 ( .A(n16313), .B(n634), .Z(n266) );
  NOR2_X2 U1496 ( .A1(n13792), .A2(n13791), .ZN(n15070) );
  AND2_X2 U1501 ( .A1(n17036), .A2(n17035), .ZN(n18332) );
  XOR2_X1 U1502 ( .A(n19622), .B(n3728), .Z(n267) );
  OR2_X1 U1504 ( .A1(n20121), .A2(n20302), .ZN(n268) );
  OR3_X1 U1506 ( .A1(n21587), .A2(n21586), .A3(n21585), .ZN(n269) );
  OR3_X1 U1507 ( .A1(n22142), .A2(n21624), .A3(n22141), .ZN(n270) );
  XOR2_X1 U1509 ( .A(n22430), .B(n22429), .Z(n271) );
  XOR2_X1 U1511 ( .A(n28450), .B(n3622), .Z(n272) );
  XOR2_X1 U1512 ( .A(n21947), .B(n1538), .Z(n274) );
  OR3_X1 U1514 ( .A1(n23897), .A2(n25006), .A3(n25005), .ZN(n276) );
  XOR2_X1 U1515 ( .A(n25211), .B(n25467), .Z(n277) );
  OR2_X1 U1517 ( .A1(n28228), .A2(n925), .ZN(n278) );
  XNOR2_X1 U1521 ( .A(n9546), .B(n9545), .ZN(n11037) );
  XNOR2_X1 U1523 ( .A(n24360), .B(n24359), .ZN(n26466) );
  XNOR2_X1 U1528 ( .A(n25292), .B(n25291), .ZN(n26717) );
  NAND4_X2 U1539 ( .A1(n8567), .A2(n8568), .A3(n8566), .A4(n8565), .ZN(n10436)
         );
  AOI22_X2 U1542 ( .A1(n16921), .A2(n17414), .B1(n15811), .B2(n15522), .ZN(
        n17679) );
  NOR2_X2 U1551 ( .A1(n5967), .A2(n16769), .ZN(n18109) );
  BUF_X1 U1552 ( .A(n23448), .Z(n292) );
  XNOR2_X1 U1553 ( .A(n22739), .B(n22738), .ZN(n23448) );
  AND2_X1 U1557 ( .A1(n11782), .A2(n11778), .ZN(n11784) );
  OR2_X1 U1561 ( .A1(n16807), .A2(n29574), .ZN(n16672) );
  BUF_X1 U1564 ( .A(n27378), .Z(n294) );
  OAI21_X1 U1566 ( .B1(n5582), .B2(n26485), .A(n26199), .ZN(n27378) );
  XNOR2_X1 U1570 ( .A(n18965), .B(n18964), .ZN(n20224) );
  BUF_X2 U1575 ( .A(n26090), .Z(n300) );
  INV_X1 U1576 ( .A(n26865), .ZN(n401) );
  OAI211_X1 U1578 ( .C1(n8795), .C2(n9034), .A(n8794), .B(n8793), .ZN(n10222)
         );
  XNOR2_X2 U1580 ( .A(n4531), .B(n16007), .ZN(n16977) );
  NAND2_X2 U1582 ( .A1(n24563), .A2(n24562), .ZN(n25947) );
  BUF_X1 U1584 ( .A(n12226), .Z(n303) );
  BUF_X1 U1593 ( .A(n27028), .Z(n307) );
  OAI22_X1 U1594 ( .A1(n26925), .A2(n28711), .B1(n23864), .B2(n29552), .ZN(
        n27028) );
  BUF_X2 U1595 ( .A(n14122), .Z(n308) );
  XNOR2_X1 U1596 ( .A(n12959), .B(n12958), .ZN(n14122) );
  NAND3_X2 U1598 ( .A1(n14503), .A2(n264), .A3(n14502), .ZN(n16558) );
  XNOR2_X2 U1599 ( .A(n7086), .B(Key[3]), .ZN(n7315) );
  AND3_X2 U1602 ( .A1(n2709), .A2(n2710), .A3(n3553), .ZN(n13445) );
  OR2_X1 U1606 ( .A1(n29541), .A2(n27364), .ZN(n799) );
  OR2_X1 U1607 ( .A1(n27074), .A2(n29622), .ZN(n3771) );
  OAI211_X1 U1617 ( .C1(n14284), .C2(n14081), .A(n13823), .B(n13822), .ZN(
        n14981) );
  XNOR2_X1 U1621 ( .A(n3582), .B(n16169), .ZN(n17466) );
  XNOR2_X2 U1623 ( .A(n21828), .B(n21827), .ZN(n23768) );
  AND2_X2 U1624 ( .A1(n21725), .A2(n21724), .ZN(n24747) );
  BUF_X1 U1626 ( .A(n16289), .Z(n320) );
  OAI211_X1 U1627 ( .C1(n4514), .C2(n4515), .A(n5016), .B(n4512), .ZN(n16289)
         );
  AND2_X1 U1628 ( .A1(n26731), .A2(n26480), .ZN(n26485) );
  NOR2_X2 U1629 ( .A1(n6601), .A2(n5441), .ZN(n22896) );
  BUF_X1 U1636 ( .A(n27718), .Z(n326) );
  AOI21_X1 U1637 ( .B1(n27690), .B2(n27688), .A(n27687), .ZN(n27718) );
  XNOR2_X2 U1640 ( .A(n1609), .B(Key[25]), .ZN(n7792) );
  OAI22_X1 U1641 ( .A1(n15032), .A2(n14825), .B1(n1644), .B2(n14826), .ZN(
        n14780) );
  OAI21_X2 U1646 ( .B1(n24136), .B2(n24135), .A(n24134), .ZN(n5275) );
  XNOR2_X1 U1649 ( .A(n24402), .B(n24401), .ZN(n26458) );
  XNOR2_X2 U1651 ( .A(n15672), .B(n15671), .ZN(n4218) );
  NAND2_X2 U1652 ( .A1(n10909), .A2(n10910), .ZN(n13414) );
  XNOR2_X2 U1654 ( .A(n4600), .B(n9933), .ZN(n11113) );
  AOI21_X2 U1661 ( .B1(n15378), .B2(n15377), .A(n15376), .ZN(n16081) );
  AND3_X2 U1665 ( .A1(n1477), .A2(n1479), .A3(n1476), .ZN(n26029) );
  AOI21_X2 U1666 ( .B1(n20775), .B2(n20774), .A(n20773), .ZN(n22219) );
  MUX2_X2 U1671 ( .A(n23237), .B(n23236), .S(n23716), .Z(n24653) );
  BUF_X1 U1674 ( .A(n337), .Z(n336) );
  OAI21_X2 U1675 ( .B1(n24083), .B2(n23506), .A(n23505), .ZN(n25751) );
  BUF_X2 U1681 ( .A(n23777), .Z(n339) );
  NOR2_X2 U1682 ( .A1(n18084), .A2(n6228), .ZN(n19717) );
  BUF_X1 U1685 ( .A(n8269), .Z(n341) );
  XNOR2_X1 U1686 ( .A(Key[147]), .B(Plaintext[147]), .ZN(n8269) );
  NAND3_X2 U1687 ( .A1(n1392), .A2(n5614), .A3(n1393), .ZN(n16563) );
  AOI22_X2 U1689 ( .A1(n23495), .A2(n23323), .B1(n23321), .B2(n23322), .ZN(
        n24672) );
  NOR3_X1 U1691 ( .A1(n25612), .A2(n25611), .A3(n25610), .ZN(n27407) );
  NOR2_X2 U1695 ( .A1(n19759), .A2(n19758), .ZN(n22143) );
  NOR2_X1 U1700 ( .A1(n470), .A2(n23946), .ZN(n1483) );
  AND2_X1 U1701 ( .A1(n20609), .A2(n29508), .ZN(n899) );
  OAI211_X2 U1703 ( .C1(n4374), .C2(n4373), .A(n4372), .B(n4371), .ZN(n19669)
         );
  OAI211_X2 U1705 ( .C1(n14100), .C2(n14099), .A(n3750), .B(n3749), .ZN(n15217) );
  OR2_X1 U1709 ( .A1(n4088), .A2(n13060), .ZN(n14350) );
  NOR2_X2 U1711 ( .A1(n17755), .A2(n5688), .ZN(n19045) );
  XNOR2_X2 U1725 ( .A(Key[35]), .B(Plaintext[35]), .ZN(n8161) );
  XNOR2_X2 U1727 ( .A(n7115), .B(Key[6]), .ZN(n7116) );
  NOR2_X2 U1731 ( .A1(n17946), .A2(n17945), .ZN(n19267) );
  NOR2_X2 U1733 ( .A1(n17126), .A2(n17125), .ZN(n18136) );
  BUF_X1 U1739 ( .A(n7369), .Z(n370) );
  XNOR2_X1 U1740 ( .A(Key[89]), .B(Plaintext[89]), .ZN(n7369) );
  NOR2_X2 U1751 ( .A1(n4648), .A2(n4602), .ZN(n24668) );
  XNOR2_X2 U1758 ( .A(n26009), .B(n26010), .ZN(n27155) );
  OAI22_X1 U1759 ( .A1(n27795), .A2(n27821), .B1(n29469), .B2(n27819), .ZN(
        n27823) );
  INV_X1 U1761 ( .A(n28025), .ZN(n376) );
  INV_X1 U1766 ( .A(n26459), .ZN(n377) );
  INV_X1 U1768 ( .A(n24215), .ZN(n378) );
  CLKBUF_X1 U1769 ( .A(n22935), .Z(n23449) );
  INV_X1 U1770 ( .A(n23266), .ZN(n379) );
  INV_X1 U1771 ( .A(n23587), .ZN(n380) );
  OAI21_X1 U1774 ( .B1(n3953), .B2(n3952), .A(n3951), .ZN(n21530) );
  INV_X1 U1775 ( .A(n21000), .ZN(n381) );
  INV_X1 U1776 ( .A(n20477), .ZN(n382) );
  INV_X1 U1779 ( .A(n20488), .ZN(n384) );
  INV_X1 U1780 ( .A(n20166), .ZN(n385) );
  INV_X1 U1781 ( .A(n20601), .ZN(n386) );
  INV_X1 U1784 ( .A(n16879), .ZN(n17382) );
  XNOR2_X1 U1785 ( .A(n16089), .B(n16088), .ZN(n17456) );
  INV_X1 U1786 ( .A(n17463), .ZN(n387) );
  NAND4_X1 U1788 ( .A1(n14859), .A2(n14862), .A3(n14860), .A4(n14861), .ZN(
        n16313) );
  BUF_X1 U1789 ( .A(n15323), .Z(n546) );
  INV_X1 U1790 ( .A(n13789), .ZN(n388) );
  XNOR2_X1 U1792 ( .A(n11670), .B(n5805), .ZN(n14479) );
  INV_X1 U1793 ( .A(n14016), .ZN(n389) );
  NAND2_X1 U1795 ( .A1(n12188), .A2(n12187), .ZN(n12128) );
  INV_X1 U1798 ( .A(n11004), .ZN(n10997) );
  INV_X1 U1799 ( .A(n10963), .ZN(n10780) );
  INV_X1 U1802 ( .A(n10948), .ZN(n391) );
  CLKBUF_X1 U1805 ( .A(n7101), .Z(n8179) );
  CLKBUF_X1 U1811 ( .A(Key[25]), .Z(n1175) );
  CLKBUF_X1 U1812 ( .A(Key[35]), .Z(n3116) );
  CLKBUF_X1 U1813 ( .A(Key[46]), .Z(n2325) );
  CLKBUF_X1 U1815 ( .A(Key[56]), .Z(n3029) );
  CLKBUF_X1 U1816 ( .A(Key[123]), .Z(n3380) );
  CLKBUF_X1 U1818 ( .A(Key[147]), .Z(n21537) );
  CLKBUF_X1 U1819 ( .A(Key[188]), .Z(n3751) );
  CLKBUF_X1 U1820 ( .A(Key[52]), .Z(n3635) );
  CLKBUF_X1 U1821 ( .A(Key[38]), .Z(n2984) );
  CLKBUF_X1 U1822 ( .A(Key[17]), .Z(n3317) );
  CLKBUF_X1 U1823 ( .A(Key[57]), .Z(n3686) );
  CLKBUF_X1 U1824 ( .A(Key[132]), .Z(n2522) );
  CLKBUF_X1 U1825 ( .A(Key[145]), .Z(n3154) );
  CLKBUF_X1 U1827 ( .A(Key[41]), .Z(n3528) );
  CLKBUF_X1 U1828 ( .A(Key[54]), .Z(n1179) );
  CLKBUF_X1 U1830 ( .A(Key[65]), .Z(n1246) );
  CLKBUF_X1 U1831 ( .A(Key[191]), .Z(n3607) );
  CLKBUF_X1 U1834 ( .A(Key[2]), .Z(n3586) );
  CLKBUF_X1 U1835 ( .A(Key[64]), .Z(n1887) );
  CLKBUF_X1 U1836 ( .A(Key[107]), .Z(n3662) );
  AOI21_X1 U1837 ( .B1(n802), .B2(n27366), .A(n29387), .ZN(n801) );
  INV_X1 U1838 ( .A(n6568), .ZN(n393) );
  INV_X1 U1841 ( .A(n27549), .ZN(n394) );
  INV_X1 U1843 ( .A(n27308), .ZN(n395) );
  OR2_X1 U1845 ( .A1(n1427), .A2(n1622), .ZN(n5582) );
  OAI21_X1 U1850 ( .B1(n26482), .B2(n1622), .A(n29501), .ZN(n1470) );
  INV_X1 U1851 ( .A(n29054), .ZN(n1279) );
  OR2_X1 U1852 ( .A1(n4678), .A2(n26426), .ZN(n2033) );
  NOR3_X1 U1853 ( .A1(n26927), .A2(n26926), .A3(n26581), .ZN(n24823) );
  AND2_X1 U1854 ( .A1(n26995), .A2(n29481), .ZN(n26735) );
  OR3_X1 U1855 ( .A1(n28532), .A2(n26632), .A3(n29481), .ZN(n25971) );
  INV_X1 U1856 ( .A(n28783), .ZN(n398) );
  CLKBUF_X1 U1857 ( .A(n25666), .Z(n26475) );
  CLKBUF_X1 U1858 ( .A(n25119), .Z(n26357) );
  INV_X1 U1860 ( .A(n27052), .ZN(n399) );
  INV_X1 U1861 ( .A(n27700), .ZN(n400) );
  INV_X1 U1862 ( .A(n26835), .ZN(n402) );
  XNOR2_X1 U1863 ( .A(n25261), .B(n25366), .ZN(n1254) );
  OAI21_X1 U1865 ( .B1(n24506), .B2(n24263), .A(n24262), .ZN(n26090) );
  OAI22_X1 U1867 ( .A1(n24506), .A2(n28523), .B1(n24505), .B2(n24806), .ZN(
        n25844) );
  OR2_X1 U1868 ( .A1(n24258), .A2(n23467), .ZN(n1250) );
  NAND2_X1 U1870 ( .A1(n28415), .A2(n25008), .ZN(n1522) );
  OR2_X1 U1872 ( .A1(n24484), .A2(n24046), .ZN(n966) );
  AND3_X1 U1873 ( .A1(n3723), .A2(n4254), .A3(n6822), .ZN(n1955) );
  CLKBUF_X1 U1874 ( .A(n23962), .Z(n24468) );
  OR2_X1 U1875 ( .A1(n23045), .A2(n477), .ZN(n1805) );
  INV_X1 U1876 ( .A(n24435), .ZN(n403) );
  OAI211_X1 U1877 ( .C1(n23061), .C2(n23344), .A(n4137), .B(n4138), .ZN(n23867) );
  INV_X1 U1878 ( .A(n24672), .ZN(n404) );
  OR2_X1 U1881 ( .A1(n481), .A2(n22531), .ZN(n1531) );
  MUX2_X1 U1882 ( .A(n480), .B(n23062), .S(n23417), .Z(n23063) );
  INV_X1 U1884 ( .A(n960), .ZN(n23622) );
  INV_X1 U1885 ( .A(n4231), .ZN(n405) );
  INV_X1 U1886 ( .A(n23612), .ZN(n406) );
  CLKBUF_X1 U1887 ( .A(n23825), .Z(n23829) );
  INV_X1 U1891 ( .A(n23820), .ZN(n407) );
  INV_X1 U1896 ( .A(n23432), .ZN(n408) );
  INV_X1 U1897 ( .A(n23250), .ZN(n409) );
  XNOR2_X1 U1898 ( .A(n22684), .B(n1818), .ZN(n23773) );
  XNOR2_X1 U1899 ( .A(n22459), .B(n621), .ZN(n22382) );
  AND2_X1 U1900 ( .A1(n5014), .A2(n5013), .ZN(n22320) );
  AOI22_X1 U1902 ( .A1(n21556), .A2(n21555), .B1(n21554), .B2(n21553), .ZN(
        n22829) );
  OR2_X1 U1905 ( .A1(n20886), .A2(n21322), .ZN(n21590) );
  INV_X1 U1909 ( .A(n1925), .ZN(n1924) );
  INV_X1 U1911 ( .A(n21679), .ZN(n412) );
  OAI22_X1 U1912 ( .A1(n821), .A2(n20474), .B1(n2062), .B2(n382), .ZN(n21328)
         );
  NAND2_X1 U1914 ( .A1(n20134), .A2(n507), .ZN(n6770) );
  AOI21_X1 U1915 ( .B1(n19920), .B2(n20619), .A(n500), .ZN(n1565) );
  NAND2_X1 U1917 ( .A1(n20586), .A2(n20587), .ZN(n1429) );
  INV_X1 U1918 ( .A(n19949), .ZN(n20587) );
  OAI21_X1 U1919 ( .B1(n502), .B2(n20109), .A(n703), .ZN(n20111) );
  INV_X1 U1920 ( .A(n20049), .ZN(n413) );
  INV_X1 U1921 ( .A(n20282), .ZN(n19808) );
  OR2_X1 U1923 ( .A1(n505), .A2(n20549), .ZN(n5982) );
  XNOR2_X1 U1924 ( .A(n19037), .B(n19038), .ZN(n20477) );
  XNOR2_X1 U1925 ( .A(n18953), .B(n18952), .ZN(n20166) );
  INV_X1 U1927 ( .A(n20088), .ZN(n414) );
  XNOR2_X1 U1929 ( .A(n16982), .B(n16983), .ZN(n20549) );
  INV_X1 U1930 ( .A(n19947), .ZN(n416) );
  XNOR2_X1 U1931 ( .A(n19504), .B(n19503), .ZN(n6843) );
  XNOR2_X1 U1932 ( .A(n19191), .B(n19452), .ZN(n19540) );
  OR2_X1 U1936 ( .A1(n18466), .A2(n1384), .ZN(n1383) );
  OR2_X1 U1937 ( .A1(n17875), .A2(n525), .ZN(n1034) );
  OR2_X1 U1938 ( .A1(n18449), .A2(n18198), .ZN(n18452) );
  AND2_X1 U1940 ( .A1(n510), .A2(n18507), .ZN(n1125) );
  AND2_X1 U1941 ( .A1(n17618), .A2(n17617), .ZN(n17825) );
  AND2_X1 U1942 ( .A1(n29044), .A2(n527), .ZN(n18189) );
  INV_X1 U1944 ( .A(n18411), .ZN(n417) );
  OR2_X1 U1945 ( .A1(n18242), .A2(n522), .ZN(n2786) );
  INV_X1 U1946 ( .A(n18507), .ZN(n418) );
  INV_X1 U1948 ( .A(n18148), .ZN(n420) );
  OAI21_X1 U1949 ( .B1(n926), .B2(n533), .A(n17394), .ZN(n1367) );
  AOI21_X1 U1950 ( .B1(n17281), .B2(n528), .A(n784), .ZN(n783) );
  NAND2_X1 U1952 ( .A1(n16067), .A2(n1464), .ZN(n17941) );
  OAI211_X1 U1953 ( .C1(n29373), .C2(n17492), .A(n4314), .B(n1153), .ZN(n4313)
         );
  INV_X1 U1954 ( .A(n6371), .ZN(n1090) );
  INV_X1 U1955 ( .A(n16812), .ZN(n421) );
  INV_X1 U1958 ( .A(n17259), .ZN(n422) );
  INV_X1 U1959 ( .A(n17571), .ZN(n423) );
  XNOR2_X1 U1961 ( .A(n16624), .B(n16623), .ZN(n16803) );
  OAI21_X1 U1964 ( .B1(n14788), .B2(n552), .A(n14787), .ZN(n16077) );
  AND3_X1 U1966 ( .A1(n1571), .A2(n552), .A3(n1570), .ZN(n13820) );
  NAND3_X1 U1968 ( .A1(n5197), .A2(n15153), .A3(n5196), .ZN(n16434) );
  OAI211_X1 U1969 ( .C1(n15518), .C2(n15519), .A(n15517), .B(n15516), .ZN(
        n15928) );
  INV_X1 U1971 ( .A(n15323), .ZN(n1926) );
  INV_X1 U1973 ( .A(n15343), .ZN(n425) );
  NAND2_X1 U1975 ( .A1(n13810), .A2(n13809), .ZN(n15182) );
  INV_X1 U1977 ( .A(n15370), .ZN(n426) );
  OAI21_X1 U1978 ( .B1(n14150), .B2(n557), .A(n713), .ZN(n14151) );
  OAI211_X1 U1979 ( .C1(n13934), .C2(n14158), .A(n646), .B(n558), .ZN(n645) );
  INV_X1 U1981 ( .A(n14358), .ZN(n13829) );
  OR2_X1 U1986 ( .A1(n14061), .A2(n13652), .ZN(n14322) );
  INV_X1 U1988 ( .A(n14293), .ZN(n428) );
  INV_X1 U1992 ( .A(n13069), .ZN(n429) );
  OR2_X1 U1994 ( .A1(n11930), .A2(n568), .ZN(n1489) );
  INV_X1 U1995 ( .A(n11951), .ZN(n11862) );
  NAND2_X1 U1997 ( .A1(n29137), .A2(n11778), .ZN(n11552) );
  NAND3_X1 U1998 ( .A1(n11051), .A2(n11050), .A3(n11049), .ZN(n12266) );
  INV_X1 U2000 ( .A(n12150), .ZN(n430) );
  INV_X1 U2001 ( .A(n10939), .ZN(n11945) );
  NAND2_X1 U2002 ( .A1(n9292), .A2(n9291), .ZN(n13086) );
  NOR2_X1 U2003 ( .A1(n1375), .A2(n9654), .ZN(n9692) );
  AOI21_X1 U2004 ( .B1(n10923), .B2(n10922), .A(n10921), .ZN(n10939) );
  OAI21_X1 U2009 ( .B1(n1359), .B2(n391), .A(n6366), .ZN(n11984) );
  NOR2_X1 U2010 ( .A1(n391), .A2(n10972), .ZN(n10969) );
  OR2_X1 U2011 ( .A1(n595), .A2(n11210), .ZN(n11082) );
  AND2_X1 U2012 ( .A1(n11210), .A2(n595), .ZN(n6604) );
  INV_X1 U2016 ( .A(n11207), .ZN(n432) );
  XNOR2_X1 U2017 ( .A(n9571), .B(n9926), .ZN(n1338) );
  INV_X1 U2019 ( .A(n11337), .ZN(n434) );
  XNOR2_X1 U2020 ( .A(n10349), .B(n1855), .ZN(n1854) );
  INV_X1 U2022 ( .A(n11218), .ZN(n435) );
  OAI21_X1 U2023 ( .B1(n606), .B2(n7328), .A(n7327), .ZN(n10007) );
  OAI211_X1 U2025 ( .C1(n8379), .C2(n882), .A(n881), .B(n880), .ZN(n10207) );
  OR2_X1 U2026 ( .A1(n937), .A2(n7714), .ZN(n2915) );
  INV_X1 U2027 ( .A(n8617), .ZN(n882) );
  OR2_X1 U2028 ( .A1(n8617), .A2(n28212), .ZN(n880) );
  INV_X1 U2033 ( .A(n8983), .ZN(n436) );
  OAI211_X1 U2034 ( .C1(n7659), .C2(n29317), .A(n7402), .B(n7401), .ZN(n9134)
         );
  OR2_X1 U2037 ( .A1(n7690), .A2(n7817), .ZN(n7501) );
  NOR2_X1 U2039 ( .A1(n7089), .A2(n29112), .ZN(n3188) );
  INV_X1 U2040 ( .A(n7997), .ZN(n437) );
  INV_X1 U2041 ( .A(n7775), .ZN(n438) );
  XNOR2_X1 U2042 ( .A(n7136), .B(Key[51]), .ZN(n7742) );
  CLKBUF_X1 U2044 ( .A(Key[174]), .Z(n3462) );
  CLKBUF_X1 U2046 ( .A(Key[93]), .Z(n1172) );
  CLKBUF_X1 U2047 ( .A(Key[49]), .Z(n1928) );
  CLKBUF_X1 U2048 ( .A(Key[159]), .Z(n1927) );
  CLKBUF_X1 U2049 ( .A(Key[20]), .Z(n3770) );
  CLKBUF_X1 U2050 ( .A(Key[10]), .Z(n2402) );
  CLKBUF_X1 U2051 ( .A(Key[86]), .Z(n2511) );
  CLKBUF_X1 U2054 ( .A(Key[149]), .Z(n3180) );
  CLKBUF_X1 U2055 ( .A(Key[142]), .Z(n3386) );
  CLKBUF_X1 U2056 ( .A(Key[110]), .Z(n1193) );
  CLKBUF_X1 U2057 ( .A(Key[50]), .Z(n3697) );
  CLKBUF_X1 U2058 ( .A(Key[27]), .Z(n3493) );
  CLKBUF_X1 U2059 ( .A(Key[23]), .Z(n3622) );
  CLKBUF_X1 U2060 ( .A(Key[72]), .Z(n3212) );
  CLKBUF_X1 U2061 ( .A(Key[103]), .Z(n2505) );
  CLKBUF_X1 U2062 ( .A(Key[96]), .Z(n3374) );
  CLKBUF_X1 U2064 ( .A(Key[13]), .Z(n5059) );
  CLKBUF_X1 U2065 ( .A(Key[94]), .Z(n1119) );
  CLKBUF_X1 U2066 ( .A(Key[81]), .Z(n2476) );
  CLKBUF_X1 U2067 ( .A(Key[179]), .Z(n1247) );
  CLKBUF_X1 U2068 ( .A(Key[104]), .Z(n3625) );
  CLKBUF_X1 U2069 ( .A(Key[146]), .Z(n2577) );
  CLKBUF_X1 U2070 ( .A(Key[16]), .Z(n730) );
  CLKBUF_X1 U2071 ( .A(Key[3]), .Z(n1187) );
  CLKBUF_X1 U2072 ( .A(Key[37]), .Z(n1248) );
  CLKBUF_X1 U2073 ( .A(Key[67]), .Z(n2441) );
  CLKBUF_X1 U2074 ( .A(Key[88]), .Z(n3114) );
  CLKBUF_X1 U2075 ( .A(Key[74]), .Z(n22489) );
  CLKBUF_X1 U2076 ( .A(Key[128]), .Z(n3211) );
  CLKBUF_X1 U2077 ( .A(Key[8]), .Z(n2973) );
  CLKBUF_X1 U2078 ( .A(Key[97]), .Z(n2509) );
  CLKBUF_X1 U2079 ( .A(Key[160]), .Z(n1046) );
  CLKBUF_X1 U2080 ( .A(Key[121]), .Z(n1184) );
  CLKBUF_X1 U2082 ( .A(Key[181]), .Z(n2385) );
  CLKBUF_X1 U2083 ( .A(Key[60]), .Z(n2541) );
  CLKBUF_X1 U2084 ( .A(Key[85]), .Z(n3067) );
  CLKBUF_X1 U2085 ( .A(Key[18]), .Z(n2381) );
  CLKBUF_X1 U2086 ( .A(Key[11]), .Z(n21865) );
  INV_X1 U2087 ( .A(n7369), .ZN(n439) );
  CLKBUF_X1 U2088 ( .A(Key[90]), .Z(n3035) );
  CLKBUF_X1 U2089 ( .A(Key[135]), .Z(n3457) );
  CLKBUF_X1 U2090 ( .A(Key[173]), .Z(n24897) );
  CLKBUF_X1 U2092 ( .A(Key[106]), .Z(n3244) );
  CLKBUF_X1 U2093 ( .A(Key[51]), .Z(n22072) );
  CLKBUF_X1 U2094 ( .A(Key[140]), .Z(n3109) );
  CLKBUF_X1 U2095 ( .A(Key[24]), .Z(n1196) );
  CLKBUF_X1 U2098 ( .A(Key[9]), .Z(n3606) );
  CLKBUF_X1 U2100 ( .A(Key[168]), .Z(n3508) );
  CLKBUF_X1 U2101 ( .A(Key[78]), .Z(n857) );
  CLKBUF_X1 U2103 ( .A(Key[118]), .Z(n3232) );
  CLKBUF_X1 U2105 ( .A(Key[114]), .Z(n3336) );
  CLKBUF_X1 U2106 ( .A(Key[34]), .Z(n2602) );
  CLKBUF_X1 U2107 ( .A(Key[69]), .Z(n3321) );
  CLKBUF_X1 U2109 ( .A(Key[22]), .Z(n2446) );
  INV_X1 U2110 ( .A(n3029), .ZN(n440) );
  CLKBUF_X1 U2111 ( .A(Key[21]), .Z(n1133) );
  CLKBUF_X1 U2112 ( .A(Key[156]), .Z(n2353) );
  CLKBUF_X1 U2114 ( .A(Key[58]), .Z(n2544) );
  CLKBUF_X1 U2115 ( .A(Key[42]), .Z(n2306) );
  CLKBUF_X1 U2116 ( .A(Key[43]), .Z(n3378) );
  CLKBUF_X1 U2117 ( .A(Key[163]), .Z(n3191) );
  CLKBUF_X1 U2118 ( .A(Key[115]), .Z(n2912) );
  CLKBUF_X1 U2119 ( .A(Key[75]), .Z(n3372) );
  CLKBUF_X1 U2120 ( .A(Key[61]), .Z(n1062) );
  CLKBUF_X1 U2121 ( .A(Key[155]), .Z(n27956) );
  CLKBUF_X1 U2122 ( .A(Key[178]), .Z(n3463) );
  CLKBUF_X1 U2123 ( .A(Key[87]), .Z(n3482) );
  CLKBUF_X1 U2124 ( .A(Key[184]), .Z(n3323) );
  CLKBUF_X1 U2126 ( .A(Key[136]), .Z(n2996) );
  CLKBUF_X1 U2128 ( .A(Key[177]), .Z(n2889) );
  CLKBUF_X1 U2129 ( .A(Key[80]), .Z(n3660) );
  CLKBUF_X1 U2130 ( .A(Key[190]), .Z(n1923) );
  CLKBUF_X1 U2131 ( .A(Key[82]), .Z(n3516) );
  CLKBUF_X1 U2132 ( .A(Key[157]), .Z(n900) );
  CLKBUF_X1 U2133 ( .A(Key[164]), .Z(n3728) );
  CLKBUF_X1 U2134 ( .A(Key[176]), .Z(n27231) );
  CLKBUF_X1 U2135 ( .A(Key[170]), .Z(n1123) );
  CLKBUF_X1 U2136 ( .A(Key[108]), .Z(n26531) );
  CLKBUF_X1 U2137 ( .A(Key[12]), .Z(n2411) );
  CLKBUF_X1 U2139 ( .A(Key[55]), .Z(n2982) );
  CLKBUF_X1 U2141 ( .A(Key[113]), .Z(n3451) );
  CLKBUF_X1 U2142 ( .A(Key[109]), .Z(n2404) );
  CLKBUF_X1 U2145 ( .A(Key[169]), .Z(n3369) );
  CLKBUF_X1 U2146 ( .A(Key[63]), .Z(n3334) );
  CLKBUF_X1 U2147 ( .A(Key[40]), .Z(n891) );
  CLKBUF_X1 U2149 ( .A(Key[120]), .Z(n2274) );
  CLKBUF_X1 U2150 ( .A(Key[14]), .Z(n2894) );
  CLKBUF_X1 U2151 ( .A(Key[33]), .Z(n3633) );
  CLKBUF_X1 U2153 ( .A(Key[127]), .Z(n2981) );
  CLKBUF_X1 U2154 ( .A(Key[141]), .Z(n3752) );
  CLKBUF_X1 U2155 ( .A(Key[28]), .Z(n2995) );
  CLKBUF_X1 U2156 ( .A(Key[76]), .Z(n2598) );
  CLKBUF_X1 U2158 ( .A(Key[148]), .Z(n1161) );
  CLKBUF_X1 U2159 ( .A(Key[137]), .Z(n3742) );
  OR2_X1 U2161 ( .A1(n26145), .A2(n27727), .ZN(n26147) );
  OR2_X1 U2162 ( .A1(n28005), .A2(n28006), .ZN(n1546) );
  AOI22_X1 U2164 ( .A1(n28027), .A2(n376), .B1(n25601), .B2(n28035), .ZN(
        n26664) );
  NOR2_X1 U2165 ( .A1(n27586), .A2(n27585), .ZN(n931) );
  INV_X1 U2166 ( .A(n1548), .ZN(n28000) );
  INV_X1 U2167 ( .A(n27862), .ZN(n27873) );
  AOI211_X1 U2168 ( .C1(n27431), .C2(n27430), .A(n1821), .B(n1820), .ZN(n1819)
         );
  OAI21_X1 U2169 ( .B1(n27387), .B2(n27408), .A(n26960), .ZN(n27403) );
  AND2_X1 U2170 ( .A1(n27387), .A2(n25629), .ZN(n27409) );
  INV_X1 U2171 ( .A(n25629), .ZN(n27400) );
  OR2_X1 U2172 ( .A1(n397), .A2(n27759), .ZN(n2794) );
  INV_X1 U2173 ( .A(n6095), .ZN(n27526) );
  NOR3_X1 U2175 ( .A1(n27429), .A2(n27426), .A3(n27425), .ZN(n1821) );
  INV_X1 U2176 ( .A(n27573), .ZN(n27553) );
  NOR2_X1 U2177 ( .A1(n29056), .A2(n28111), .ZN(n1691) );
  NOR2_X1 U2178 ( .A1(n28089), .A2(n28111), .ZN(n28109) );
  NOR2_X1 U2179 ( .A1(n27830), .A2(n27829), .ZN(n27100) );
  OR2_X1 U2180 ( .A1(n27938), .A2(n27244), .ZN(n1011) );
  OR2_X1 U2181 ( .A1(n28016), .A2(n28017), .ZN(n1548) );
  NOR2_X1 U2182 ( .A1(n27855), .A2(n26641), .ZN(n26696) );
  INV_X1 U2184 ( .A(n27362), .ZN(n27370) );
  INV_X1 U2185 ( .A(n28179), .ZN(n930) );
  INV_X1 U2187 ( .A(n27588), .ZN(n933) );
  NOR2_X1 U2188 ( .A1(n27582), .A2(n27590), .ZN(n27589) );
  INV_X1 U2189 ( .A(n27439), .ZN(n26829) );
  NOR2_X1 U2190 ( .A1(n26069), .A2(n26068), .ZN(n27728) );
  AND3_X1 U2191 ( .A1(n27429), .A2(n27428), .A3(n27427), .ZN(n1820) );
  AND3_X1 U2192 ( .A1(n5735), .A2(n24825), .A3(n24824), .ZN(n6568) );
  NOR2_X1 U2194 ( .A1(n25201), .A2(n25200), .ZN(n27549) );
  NOR2_X1 U2195 ( .A1(n27547), .A2(n26652), .ZN(n27200) );
  INV_X1 U2196 ( .A(n27630), .ZN(n442) );
  OAI211_X1 U2197 ( .C1(n26361), .C2(n1076), .A(n2033), .B(n1075), .ZN(n27614)
         );
  INV_X1 U2198 ( .A(n28019), .ZN(n443) );
  INV_X1 U2199 ( .A(n27301), .ZN(n444) );
  INV_X1 U2200 ( .A(n28016), .ZN(n445) );
  AND2_X1 U2203 ( .A1(n3703), .A2(n3702), .ZN(n27286) );
  NOR2_X1 U2204 ( .A1(n1968), .A2(n26262), .ZN(n27597) );
  INV_X1 U2205 ( .A(n27213), .ZN(n446) );
  INV_X1 U2208 ( .A(n27863), .ZN(n27871) );
  NAND3_X1 U2209 ( .A1(n798), .A2(n29055), .A3(n4173), .ZN(n27362) );
  INV_X1 U2210 ( .A(n27859), .ZN(n447) );
  NOR2_X1 U2213 ( .A1(n26743), .A2(n26744), .ZN(n28090) );
  INV_X1 U2215 ( .A(n27465), .ZN(n449) );
  MUX2_X1 U2218 ( .A(n26509), .B(n26508), .S(n27084), .Z(n26639) );
  OAI21_X1 U2220 ( .B1(n27122), .B2(n26516), .A(n26515), .ZN(n27854) );
  NOR2_X1 U2221 ( .A1(n26635), .A2(n26634), .ZN(n27972) );
  OAI21_X1 U2222 ( .B1(n26301), .B2(n27904), .A(n25953), .ZN(n27863) );
  AOI21_X1 U2223 ( .B1(n27151), .B2(n401), .A(n27152), .ZN(n3590) );
  NOR2_X1 U2224 ( .A1(n26356), .A2(n28650), .ZN(n27186) );
  AND2_X1 U2225 ( .A1(n28575), .A2(n26761), .ZN(n1169) );
  NAND2_X1 U2226 ( .A1(n27012), .A2(n399), .ZN(n1535) );
  INV_X1 U2228 ( .A(n1622), .ZN(n1472) );
  AND2_X1 U2229 ( .A1(n26727), .A2(n26480), .ZN(n1533) );
  NOR2_X1 U2231 ( .A1(n26241), .A2(n26753), .ZN(n25650) );
  BUF_X1 U2232 ( .A(n26729), .Z(n26482) );
  NOR2_X1 U2233 ( .A1(n26200), .A2(n26235), .ZN(n26741) );
  OAI21_X1 U2234 ( .B1(n26461), .B2(n26457), .A(n28578), .ZN(n949) );
  AOI21_X1 U2235 ( .B1(n28504), .B2(n27161), .A(n27701), .ZN(n5994) );
  OR2_X1 U2236 ( .A1(n27124), .A2(n28513), .ZN(n5486) );
  OR3_X1 U2237 ( .A1(n26426), .A2(n26382), .A3(n26381), .ZN(n26383) );
  INV_X1 U2238 ( .A(n26736), .ZN(n826) );
  INV_X1 U2240 ( .A(n25406), .ZN(n26469) );
  INV_X1 U2241 ( .A(n27067), .ZN(n922) );
  XNOR2_X1 U2244 ( .A(n6436), .B(n25064), .ZN(n4820) );
  OR2_X1 U2245 ( .A1(n26997), .A2(n26733), .ZN(n26736) );
  XNOR2_X1 U2247 ( .A(n23941), .B(n23940), .ZN(n26448) );
  BUF_X1 U2250 ( .A(n25676), .Z(n27041) );
  XNOR2_X1 U2253 ( .A(n24988), .B(n24989), .ZN(n27169) );
  INV_X1 U2254 ( .A(n26727), .ZN(n1622) );
  INV_X1 U2256 ( .A(n25365), .ZN(n26928) );
  XNOR2_X1 U2261 ( .A(n25742), .B(n25741), .ZN(n5263) );
  XNOR2_X1 U2264 ( .A(n25804), .B(n25805), .ZN(n26841) );
  INV_X1 U2267 ( .A(n26919), .ZN(n454) );
  XNOR2_X1 U2269 ( .A(n24695), .B(n24696), .ZN(n25365) );
  XNOR2_X1 U2270 ( .A(n4084), .B(n4082), .ZN(n26740) );
  INV_X1 U2271 ( .A(n27704), .ZN(n455) );
  INV_X1 U2272 ( .A(n26941), .ZN(n456) );
  XNOR2_X1 U2273 ( .A(n25587), .B(n25586), .ZN(n26995) );
  INV_X1 U2274 ( .A(n26917), .ZN(n457) );
  XNOR2_X1 U2276 ( .A(n23893), .B(n23892), .ZN(n26179) );
  NOR2_X1 U2278 ( .A1(n24981), .A2(n24980), .ZN(n25411) );
  XNOR2_X1 U2279 ( .A(n1303), .B(n25891), .ZN(n1302) );
  XNOR2_X1 U2280 ( .A(n25262), .B(n26070), .ZN(n25081) );
  INV_X1 U2282 ( .A(n24870), .ZN(n25944) );
  XNOR2_X1 U2283 ( .A(n25703), .B(n5146), .ZN(n26101) );
  AND3_X1 U2284 ( .A1(n4691), .A2(n4694), .A3(n4690), .ZN(n25369) );
  NOR2_X1 U2285 ( .A1(n24615), .A2(n5136), .ZN(n25876) );
  NOR2_X1 U2287 ( .A1(n3567), .A2(n24122), .ZN(n25268) );
  NOR2_X1 U2288 ( .A1(n22871), .A2(n22872), .ZN(n25293) );
  OR2_X1 U2289 ( .A1(n820), .A2(n3654), .ZN(n1458) );
  AND4_X1 U2295 ( .A1(n276), .A2(n1517), .A3(n25007), .A4(n1515), .ZN(n1514)
         );
  OAI211_X1 U2296 ( .C1(n24442), .C2(n24441), .A(n24440), .B(n24439), .ZN(
        n25564) );
  OR2_X1 U2297 ( .A1(n1283), .A2(n24589), .ZN(n1282) );
  OR2_X1 U2300 ( .A1(n24649), .A2(n672), .ZN(n24660) );
  INV_X1 U2302 ( .A(n966), .ZN(n24482) );
  OAI22_X1 U2303 ( .A1(n24083), .A2(n24408), .B1(n6266), .B2(n24405), .ZN(
        n24407) );
  AND2_X1 U2304 ( .A1(n23971), .A2(n24479), .ZN(n1655) );
  NOR2_X1 U2305 ( .A1(n24806), .A2(n803), .ZN(n24263) );
  INV_X1 U2308 ( .A(n24454), .ZN(n458) );
  INV_X1 U2309 ( .A(n29555), .ZN(n1274) );
  NOR2_X1 U2311 ( .A1(n24467), .A2(n24582), .ZN(n1203) );
  INV_X1 U2312 ( .A(n24278), .ZN(n24590) );
  INV_X1 U2313 ( .A(n1808), .ZN(n24338) );
  NOR2_X1 U2314 ( .A1(n25793), .A2(n25794), .ZN(n25800) );
  AND2_X1 U2315 ( .A1(n24745), .A2(n24751), .ZN(n24616) );
  INV_X1 U2316 ( .A(n24612), .ZN(n459) );
  INV_X1 U2317 ( .A(n23389), .ZN(n811) );
  OR2_X1 U2318 ( .A1(n831), .A2(n24592), .ZN(n2586) );
  AND2_X1 U2319 ( .A1(n24739), .A2(n24735), .ZN(n24604) );
  NOR2_X1 U2320 ( .A1(n22867), .A2(n22866), .ZN(n24173) );
  INV_X1 U2321 ( .A(n24706), .ZN(n24417) );
  NAND2_X1 U2322 ( .A1(n24339), .A2(n24340), .ZN(n3731) );
  OR2_X1 U2323 ( .A1(n24388), .A2(n24077), .ZN(n24135) );
  AND2_X1 U2324 ( .A1(n4849), .A2(n2557), .ZN(n1856) );
  INV_X1 U2325 ( .A(n831), .ZN(n4693) );
  AND2_X1 U2326 ( .A1(n25008), .A2(n24138), .ZN(n1516) );
  INV_X1 U2327 ( .A(n24804), .ZN(n24162) );
  OR2_X1 U2328 ( .A1(n24241), .A2(n24559), .ZN(n1726) );
  OR2_X1 U2330 ( .A1(n24133), .A2(n24081), .ZN(n1617) );
  INV_X1 U2332 ( .A(n3061), .ZN(n673) );
  INV_X1 U2334 ( .A(n29695), .ZN(n460) );
  OR2_X1 U2335 ( .A1(n24629), .A2(n4364), .ZN(n24531) );
  OR2_X1 U2336 ( .A1(n23897), .A2(n25008), .ZN(n1515) );
  INV_X1 U2337 ( .A(n24747), .ZN(n1631) );
  INV_X1 U2338 ( .A(n24457), .ZN(n1426) );
  INV_X1 U2339 ( .A(n29309), .ZN(n24775) );
  INV_X1 U2340 ( .A(n24369), .ZN(n461) );
  INV_X1 U2341 ( .A(n24745), .ZN(n462) );
  AND2_X1 U2342 ( .A1(n24891), .A2(n24631), .ZN(n23982) );
  OR2_X1 U2347 ( .A1(n25008), .A2(n24138), .ZN(n1448) );
  INV_X1 U2348 ( .A(n23945), .ZN(n463) );
  INV_X1 U2349 ( .A(n1955), .ZN(n464) );
  AND2_X1 U2350 ( .A1(n5696), .A2(n5698), .ZN(n24555) );
  INV_X1 U2354 ( .A(n24635), .ZN(n465) );
  OAI211_X1 U2355 ( .C1(n23741), .C2(n23383), .A(n1638), .B(n1637), .ZN(n24133) );
  OAI21_X1 U2356 ( .B1(n23444), .B2(n4794), .A(n2169), .ZN(n1498) );
  NOR2_X1 U2358 ( .A1(n21929), .A2(n6310), .ZN(n6309) );
  OAI21_X1 U2359 ( .B1(n23424), .B2(n23426), .A(n23115), .ZN(n24483) );
  INV_X1 U2360 ( .A(n24310), .ZN(n466) );
  OR2_X1 U2362 ( .A1(n24367), .A2(n24138), .ZN(n1551) );
  INV_X1 U2364 ( .A(n24972), .ZN(n468) );
  NAND2_X1 U2366 ( .A1(n5080), .A2(n24093), .ZN(n24489) );
  AND2_X1 U2367 ( .A1(n23805), .A2(n22742), .ZN(n1240) );
  AND3_X1 U2368 ( .A1(n6609), .A2(n6608), .A3(n6607), .ZN(n24337) );
  INV_X1 U2369 ( .A(n24211), .ZN(n469) );
  AOI21_X1 U2370 ( .B1(n1531), .B2(n22863), .A(n23835), .ZN(n22867) );
  AOI22_X1 U2371 ( .A1(n23690), .A2(n23802), .B1(n23689), .B2(n23688), .ZN(
        n24205) );
  INV_X1 U2372 ( .A(n24779), .ZN(n470) );
  OR2_X1 U2376 ( .A1(n23440), .A2(n23441), .ZN(n1228) );
  INV_X1 U2378 ( .A(n24509), .ZN(n471) );
  AND2_X1 U2380 ( .A1(n23189), .A2(n1286), .ZN(n23757) );
  OR2_X1 U2381 ( .A1(n23253), .A2(n23252), .ZN(n867) );
  OAI22_X1 U2382 ( .A1(n6054), .A2(n2141), .B1(n943), .B2(n23735), .ZN(n22009)
         );
  OR2_X1 U2383 ( .A1(n2066), .A2(n23558), .ZN(n1556) );
  OR3_X1 U2384 ( .A1(n23180), .A2(n23645), .A3(n23643), .ZN(n23181) );
  OAI21_X1 U2385 ( .B1(n808), .B2(n23787), .A(n23036), .ZN(n1642) );
  OR2_X1 U2386 ( .A1(n23395), .A2(n23396), .ZN(n907) );
  AND2_X1 U2387 ( .A1(n754), .A2(n755), .ZN(n23402) );
  OR2_X1 U2388 ( .A1(n23384), .A2(n23385), .ZN(n1637) );
  AND2_X1 U2389 ( .A1(n23442), .A2(n23370), .ZN(n23444) );
  NOR2_X1 U2390 ( .A1(n23626), .A2(n23566), .ZN(n23274) );
  NOR2_X1 U2391 ( .A1(n23074), .A2(n28653), .ZN(n23811) );
  OR2_X1 U2392 ( .A1(n23538), .A2(n1913), .ZN(n712) );
  AND3_X1 U2393 ( .A1(n28594), .A2(n23807), .A3(n29102), .ZN(n23814) );
  AND2_X1 U2394 ( .A1(n22451), .A2(n22452), .ZN(n23704) );
  NAND2_X1 U2395 ( .A1(n23787), .A2(n23786), .ZN(n1641) );
  AND2_X1 U2396 ( .A1(n23305), .A2(n22686), .ZN(n23303) );
  OR2_X1 U2397 ( .A1(n23808), .A2(n29102), .ZN(n1284) );
  OR2_X1 U2398 ( .A1(n23073), .A2(n23099), .ZN(n2400) );
  INV_X1 U2399 ( .A(n23615), .ZN(n760) );
  OR2_X1 U2401 ( .A1(n23829), .A2(n23382), .ZN(n23383) );
  OR2_X1 U2405 ( .A1(n23735), .A2(n23736), .ZN(n755) );
  XNOR2_X1 U2406 ( .A(n21782), .B(n21781), .ZN(n23767) );
  XNOR2_X1 U2407 ( .A(n4228), .B(n22924), .ZN(n23461) );
  INV_X1 U2409 ( .A(n23784), .ZN(n473) );
  XNOR2_X1 U2410 ( .A(n22203), .B(n22202), .ZN(n23612) );
  INV_X1 U2411 ( .A(n23679), .ZN(n474) );
  INV_X1 U2412 ( .A(n23825), .ZN(n885) );
  XNOR2_X1 U2415 ( .A(n22276), .B(n2393), .ZN(n23633) );
  INV_X1 U2416 ( .A(n23787), .ZN(n475) );
  XNOR2_X1 U2417 ( .A(n22324), .B(n22323), .ZN(n23762) );
  INV_X1 U2418 ( .A(n379), .ZN(n476) );
  INV_X1 U2419 ( .A(n23557), .ZN(n477) );
  XNOR2_X1 U2421 ( .A(n22816), .B(n22817), .ZN(n23820) );
  INV_X1 U2423 ( .A(n23647), .ZN(n641) );
  CLKBUF_X1 U2425 ( .A(n23258), .Z(n23398) );
  INV_X1 U2426 ( .A(n22979), .ZN(n23405) );
  INV_X1 U2429 ( .A(n22946), .ZN(n23385) );
  INV_X1 U2430 ( .A(n23416), .ZN(n479) );
  OR2_X1 U2431 ( .A1(n23733), .A2(n23258), .ZN(n754) );
  INV_X1 U2432 ( .A(n23099), .ZN(n480) );
  INV_X1 U2433 ( .A(n23077), .ZN(n481) );
  INV_X1 U2434 ( .A(n23382), .ZN(n482) );
  INV_X1 U2436 ( .A(n23419), .ZN(n483) );
  INV_X1 U2437 ( .A(n28164), .ZN(n484) );
  INV_X1 U2439 ( .A(n23418), .ZN(n485) );
  INV_X1 U2440 ( .A(n23360), .ZN(n486) );
  XNOR2_X1 U2441 ( .A(n22425), .B(n22424), .ZN(n23647) );
  INV_X1 U2443 ( .A(n28460), .ZN(n487) );
  XNOR2_X1 U2447 ( .A(n21835), .B(n21834), .ZN(n23777) );
  XNOR2_X1 U2448 ( .A(n22390), .B(n1451), .ZN(n23618) );
  XNOR2_X1 U2449 ( .A(n1500), .B(n22711), .ZN(n1055) );
  XNOR2_X1 U2450 ( .A(n22610), .B(n22007), .ZN(n4968) );
  XNOR2_X1 U2451 ( .A(n22156), .B(n22155), .ZN(n23587) );
  XNOR2_X1 U2454 ( .A(n22522), .B(n3372), .ZN(n1538) );
  XNOR2_X1 U2455 ( .A(n22912), .B(n21990), .ZN(n22533) );
  XNOR2_X1 U2456 ( .A(n22923), .B(n1501), .ZN(n1500) );
  INV_X1 U2457 ( .A(n22710), .ZN(n1501) );
  XNOR2_X1 U2460 ( .A(n21982), .B(n22110), .ZN(n22395) );
  XNOR2_X1 U2461 ( .A(n22245), .B(n3635), .ZN(n6389) );
  XNOR2_X1 U2462 ( .A(n22830), .B(n22525), .ZN(n21847) );
  INV_X1 U2464 ( .A(n22690), .ZN(n22169) );
  AND2_X1 U2468 ( .A1(n20991), .A2(n20990), .ZN(n22006) );
  INV_X1 U2470 ( .A(n22099), .ZN(n22098) );
  AND2_X1 U2471 ( .A1(n20185), .A2(n5018), .ZN(n22132) );
  NAND3_X1 U2472 ( .A1(n270), .A2(n3889), .A3(n3891), .ZN(n1271) );
  OAI211_X1 U2476 ( .C1(n21619), .C2(n21618), .A(n21617), .B(n21616), .ZN(
        n22813) );
  AND3_X1 U2478 ( .A1(n1289), .A2(n269), .A3(n1288), .ZN(n3486) );
  OR2_X1 U2479 ( .A1(n19859), .A2(n4467), .ZN(n4466) );
  OAI211_X1 U2480 ( .C1(n21619), .C2(n20906), .A(n20524), .B(n20523), .ZN(
        n22609) );
  AND3_X1 U2482 ( .A1(n650), .A2(n648), .A3(n647), .ZN(n3578) );
  OR2_X1 U2486 ( .A1(n21748), .A2(n20658), .ZN(n1327) );
  AOI22_X1 U2487 ( .A1(n1621), .A2(n21550), .B1(n21553), .B2(n21547), .ZN(
        n21181) );
  AND2_X1 U2488 ( .A1(n21178), .A2(n21179), .ZN(n879) );
  OAI21_X1 U2489 ( .B1(n21015), .B2(n21016), .A(n22404), .ZN(n1720) );
  AOI21_X1 U2490 ( .B1(n21236), .B2(n21237), .A(n21748), .ZN(n952) );
  OAI21_X1 U2491 ( .B1(n20844), .B2(n1814), .A(n21125), .ZN(n1083) );
  AND2_X1 U2493 ( .A1(n20848), .A2(n21481), .ZN(n854) );
  OR2_X1 U2494 ( .A1(n28791), .A2(n21334), .ZN(n4776) );
  OR2_X1 U2495 ( .A1(n4960), .A2(n20744), .ZN(n3119) );
  AND2_X1 U2497 ( .A1(n21306), .A2(n21311), .ZN(n906) );
  INV_X1 U2498 ( .A(n21171), .ZN(n21409) );
  NOR2_X1 U2499 ( .A1(n20688), .A2(n20689), .ZN(n21716) );
  INV_X1 U2500 ( .A(n21090), .ZN(n701) );
  INV_X1 U2501 ( .A(n21530), .ZN(n1543) );
  INV_X1 U2502 ( .A(n21532), .ZN(n1540) );
  OR2_X1 U2504 ( .A1(n20886), .A2(n21587), .ZN(n1288) );
  INV_X1 U2505 ( .A(n20786), .ZN(n21930) );
  NOR2_X1 U2507 ( .A1(n22286), .A2(n22290), .ZN(n1693) );
  INV_X1 U2508 ( .A(n21221), .ZN(n20703) );
  OR2_X1 U2509 ( .A1(n21113), .A2(n21464), .ZN(n4224) );
  INV_X1 U2511 ( .A(n20988), .ZN(n20914) );
  OR2_X1 U2516 ( .A1(n20854), .A2(n21145), .ZN(n2427) );
  INV_X1 U2517 ( .A(n21213), .ZN(n489) );
  INV_X1 U2518 ( .A(n21574), .ZN(n21485) );
  INV_X1 U2519 ( .A(n20783), .ZN(n21550) );
  AND2_X1 U2520 ( .A1(n21014), .A2(n21429), .ZN(n21016) );
  INV_X1 U2521 ( .A(n21736), .ZN(n21471) );
  NOR2_X1 U2524 ( .A1(n20878), .A2(n20877), .ZN(n20879) );
  INV_X1 U2525 ( .A(n21119), .ZN(n21117) );
  INV_X1 U2527 ( .A(n21408), .ZN(n490) );
  INV_X1 U2529 ( .A(n20393), .ZN(n21541) );
  AND2_X1 U2530 ( .A1(n21599), .A2(n21600), .ZN(n20905) );
  AND2_X1 U2531 ( .A1(n6771), .A2(n6770), .ZN(n20899) );
  AND2_X1 U2532 ( .A1(n21679), .A2(n21674), .ZN(n21449) );
  OR2_X1 U2534 ( .A1(n19980), .A2(n6114), .ZN(n649) );
  OR2_X1 U2535 ( .A1(n21118), .A2(n21145), .ZN(n21141) );
  INV_X1 U2537 ( .A(n21078), .ZN(n491) );
  OR2_X1 U2545 ( .A1(n6577), .A2(n19994), .ZN(n1462) );
  INV_X1 U2546 ( .A(n21143), .ZN(n492) );
  INV_X1 U2548 ( .A(n21473), .ZN(n493) );
  OR2_X1 U2549 ( .A1(n20045), .A2(n19985), .ZN(n18884) );
  NOR2_X1 U2550 ( .A1(n20328), .A2(n28491), .ZN(n1335) );
  INV_X1 U2551 ( .A(n20744), .ZN(n494) );
  AND2_X1 U2552 ( .A1(n681), .A2(n680), .ZN(n20139) );
  INV_X1 U2555 ( .A(n20533), .ZN(n495) );
  OAI211_X1 U2556 ( .C1(n20198), .C2(n20588), .A(n1428), .B(n1429), .ZN(n21679) );
  OR2_X1 U2560 ( .A1(n18848), .A2(n836), .ZN(n835) );
  INV_X1 U2561 ( .A(n21704), .ZN(n496) );
  INV_X1 U2562 ( .A(n21400), .ZN(n497) );
  AOI21_X1 U2563 ( .B1(n19808), .B2(n20284), .A(n20283), .ZN(n680) );
  INV_X1 U2568 ( .A(n21362), .ZN(n19458) );
  INV_X1 U2569 ( .A(n6840), .ZN(n21248) );
  INV_X1 U2572 ( .A(n20248), .ZN(n20636) );
  NOR2_X1 U2573 ( .A1(n20354), .A2(n20478), .ZN(n20474) );
  AND2_X1 U2574 ( .A1(n20162), .A2(n29066), .ZN(n19872) );
  AND2_X1 U2575 ( .A1(n384), .A2(n20486), .ZN(n869) );
  AND2_X1 U2576 ( .A1(n19765), .A2(n20049), .ZN(n18848) );
  INV_X1 U2577 ( .A(n21353), .ZN(n20517) );
  OR2_X1 U2579 ( .A1(n4657), .A2(n19973), .ZN(n4656) );
  OR2_X1 U2581 ( .A1(n20607), .A2(n20441), .ZN(n20612) );
  INV_X1 U2582 ( .A(n19993), .ZN(n20222) );
  INV_X1 U2583 ( .A(n20549), .ZN(n1781) );
  XNOR2_X1 U2584 ( .A(n19674), .B(n19673), .ZN(n20137) );
  INV_X1 U2586 ( .A(n20504), .ZN(n1626) );
  BUF_X1 U2587 ( .A(n18699), .Z(n20379) );
  INV_X1 U2589 ( .A(n20637), .ZN(n498) );
  OR2_X1 U2591 ( .A1(n20299), .A2(n20130), .ZN(n1178) );
  XNOR2_X1 U2592 ( .A(n19545), .B(n19544), .ZN(n19554) );
  XNOR2_X1 U2593 ( .A(n19319), .B(n19318), .ZN(n1881) );
  AND2_X1 U2594 ( .A1(n20209), .A2(n19851), .ZN(n20397) );
  OR2_X1 U2595 ( .A1(n19993), .A2(n20166), .ZN(n20221) );
  INV_X1 U2596 ( .A(n20209), .ZN(n20394) );
  XNOR2_X1 U2597 ( .A(n19352), .B(n19353), .ZN(n19920) );
  OR2_X1 U2598 ( .A1(n20458), .A2(n4569), .ZN(n20275) );
  INV_X1 U2599 ( .A(n20182), .ZN(n499) );
  INV_X1 U2600 ( .A(n20431), .ZN(n500) );
  XNOR2_X1 U2601 ( .A(n18623), .B(n19690), .ZN(n20567) );
  XNOR2_X1 U2602 ( .A(n18911), .B(n18910), .ZN(n20144) );
  XNOR2_X1 U2604 ( .A(n1757), .B(n19617), .ZN(n1755) );
  INV_X1 U2607 ( .A(n21355), .ZN(n501) );
  BUF_X1 U2609 ( .A(n19093), .Z(n20239) );
  XNOR2_X1 U2610 ( .A(n774), .B(n773), .ZN(n20618) );
  INV_X1 U2611 ( .A(n28140), .ZN(n503) );
  XNOR2_X1 U2612 ( .A(n17655), .B(n17656), .ZN(n20580) );
  XNOR2_X1 U2613 ( .A(n17606), .B(n17605), .ZN(n20414) );
  XNOR2_X1 U2615 ( .A(n18678), .B(n18679), .ZN(n20375) );
  INV_X1 U2616 ( .A(n20178), .ZN(n504) );
  XNOR2_X1 U2619 ( .A(n5211), .B(n18721), .ZN(n20088) );
  XNOR2_X1 U2621 ( .A(n5161), .B(n19484), .ZN(n19315) );
  XNOR2_X1 U2622 ( .A(n18116), .B(n18115), .ZN(n19947) );
  XNOR2_X1 U2623 ( .A(n19591), .B(n775), .ZN(n774) );
  INV_X1 U2624 ( .A(n19855), .ZN(n505) );
  INV_X1 U2625 ( .A(n20284), .ZN(n506) );
  XNOR2_X1 U2626 ( .A(n19225), .B(n3087), .ZN(n1757) );
  XNOR2_X1 U2627 ( .A(n1823), .B(n1822), .ZN(n20130) );
  INV_X1 U2628 ( .A(n19270), .ZN(n1054) );
  XNOR2_X1 U2631 ( .A(n18804), .B(n18805), .ZN(n20098) );
  XNOR2_X1 U2632 ( .A(n18985), .B(n18986), .ZN(n20173) );
  INV_X1 U2633 ( .A(n6843), .ZN(n507) );
  XNOR2_X1 U2634 ( .A(n1504), .B(n19349), .ZN(n19445) );
  XNOR2_X1 U2635 ( .A(n1825), .B(n1824), .ZN(n1822) );
  XNOR2_X1 U2636 ( .A(n19330), .B(n267), .ZN(n773) );
  XNOR2_X1 U2637 ( .A(n18782), .B(n19332), .ZN(n19175) );
  NOR2_X1 U2638 ( .A1(n18594), .A2(n2341), .ZN(n19300) );
  INV_X1 U2640 ( .A(n1733), .ZN(n1783) );
  XNOR2_X1 U2642 ( .A(n19481), .B(n19483), .ZN(n1825) );
  XNOR2_X1 U2644 ( .A(n1733), .B(n19207), .ZN(n19528) );
  XNOR2_X1 U2645 ( .A(n19192), .B(n1741), .ZN(n19356) );
  INV_X1 U2646 ( .A(n19086), .ZN(n18906) );
  XNOR2_X1 U2647 ( .A(n19206), .B(n18695), .ZN(n19330) );
  INV_X1 U2648 ( .A(n19490), .ZN(n18085) );
  NAND2_X1 U2649 ( .A1(n2150), .A2(n2147), .ZN(n19475) );
  INV_X1 U2650 ( .A(n19246), .ZN(n19616) );
  INV_X1 U2651 ( .A(n19349), .ZN(n1505) );
  INV_X1 U2653 ( .A(n19228), .ZN(n1503) );
  XNOR2_X1 U2655 ( .A(n19482), .B(n22072), .ZN(n1824) );
  OR2_X1 U2661 ( .A1(n1455), .A2(n17602), .ZN(n19490) );
  AND3_X1 U2663 ( .A1(n1506), .A2(n18066), .A3(n18065), .ZN(n19349) );
  NAND2_X1 U2664 ( .A1(n16981), .A2(n3544), .ZN(n19483) );
  NOR2_X1 U2666 ( .A1(n5178), .A2(n17936), .ZN(n19323) );
  NOR2_X1 U2672 ( .A1(n17591), .A2(n17590), .ZN(n18725) );
  AND3_X1 U2673 ( .A1(n2045), .A2(n5857), .A3(n5985), .ZN(n19122) );
  AND3_X1 U2676 ( .A1(n2770), .A2(n2771), .A3(n17757), .ZN(n19273) );
  AND2_X1 U2678 ( .A1(n17638), .A2(n6930), .ZN(n19305) );
  AND2_X1 U2682 ( .A1(n18181), .A2(n18444), .ZN(n18448) );
  INV_X1 U2683 ( .A(n18100), .ZN(n18199) );
  MUX2_X1 U2686 ( .A(n18219), .B(n18218), .S(n18217), .Z(n18877) );
  OAI21_X1 U2687 ( .B1(n17652), .B2(n17653), .A(n17651), .ZN(n18773) );
  INV_X1 U2688 ( .A(n3439), .ZN(n1731) );
  OR2_X1 U2689 ( .A1(n18098), .A2(n18444), .ZN(n1304) );
  INV_X1 U2691 ( .A(n18173), .ZN(n1708) );
  AND2_X1 U2692 ( .A1(n17942), .A2(n17941), .ZN(n1433) );
  AND2_X1 U2694 ( .A1(n18304), .A2(n18306), .ZN(n17933) );
  INV_X1 U2695 ( .A(n17793), .ZN(n671) );
  OR2_X1 U2696 ( .A1(n18333), .A2(n817), .ZN(n17652) );
  OR2_X1 U2697 ( .A1(n18195), .A2(n18449), .ZN(n18100) );
  AND2_X1 U2698 ( .A1(n15734), .A2(n18490), .ZN(n18016) );
  AND2_X1 U2699 ( .A1(n17858), .A2(n18285), .ZN(n18521) );
  INV_X1 U2700 ( .A(n420), .ZN(n1758) );
  AND2_X1 U2701 ( .A1(n18261), .A2(n18263), .ZN(n697) );
  AND2_X1 U2702 ( .A1(n17842), .A2(n18242), .ZN(n2787) );
  AND2_X1 U2704 ( .A1(n17564), .A2(n17771), .ZN(n1378) );
  INV_X1 U2705 ( .A(n18706), .ZN(n876) );
  NOR2_X1 U2706 ( .A1(n18333), .A2(n18334), .ZN(n1180) );
  OR2_X1 U2707 ( .A1(n18402), .A2(n18232), .ZN(n1524) );
  AND2_X1 U2708 ( .A1(n18268), .A2(n18326), .ZN(n1717) );
  INV_X1 U2709 ( .A(n18422), .ZN(n1530) );
  OR2_X1 U2711 ( .A1(n17132), .A2(n17131), .ZN(n18137) );
  NAND2_X1 U2712 ( .A1(n6643), .A2(n6642), .ZN(n18537) );
  INV_X1 U2713 ( .A(n18342), .ZN(n17906) );
  AND2_X1 U2714 ( .A1(n15892), .A2(n18299), .ZN(n18061) );
  OAI21_X1 U2715 ( .B1(n17717), .B2(n17431), .A(n5329), .ZN(n18522) );
  INV_X1 U2716 ( .A(n817), .ZN(n4412) );
  OR2_X1 U2720 ( .A1(n17939), .A2(n17872), .ZN(n1436) );
  INV_X1 U2722 ( .A(n18040), .ZN(n17824) );
  AND2_X1 U2723 ( .A1(n18421), .A2(n17802), .ZN(n1577) );
  AND2_X1 U2724 ( .A1(n18040), .A2(n18421), .ZN(n1576) );
  INV_X1 U2725 ( .A(n17864), .ZN(n509) );
  NAND4_X1 U2726 ( .A1(n679), .A2(n16893), .A3(n16892), .A4(n16894), .ZN(
        n18511) );
  OAI211_X1 U2727 ( .C1(n16825), .C2(n4571), .A(n4113), .B(n4112), .ZN(n18476)
         );
  OAI21_X1 U2728 ( .B1(n1509), .B2(n17037), .A(n1508), .ZN(n18299) );
  INV_X1 U2729 ( .A(n1384), .ZN(n17916) );
  INV_X1 U2730 ( .A(n18508), .ZN(n510) );
  INV_X1 U2733 ( .A(n18441), .ZN(n513) );
  OAI21_X1 U2736 ( .B1(n17513), .B2(n4273), .A(n4705), .ZN(n17696) );
  INV_X1 U2737 ( .A(n18506), .ZN(n515) );
  AND2_X1 U2738 ( .A1(n18251), .A2(n18017), .ZN(n17961) );
  AND2_X1 U2739 ( .A1(n18020), .A2(n18017), .ZN(n17959) );
  NOR2_X1 U2741 ( .A1(n17021), .A2(n17020), .ZN(n17854) );
  INV_X1 U2742 ( .A(n18172), .ZN(n516) );
  AND2_X1 U2743 ( .A1(n1665), .A2(n1667), .ZN(n17781) );
  INV_X1 U2745 ( .A(n17601), .ZN(n517) );
  INV_X1 U2746 ( .A(n19560), .ZN(n18188) );
  OR2_X1 U2748 ( .A1(n17059), .A2(n17058), .ZN(n817) );
  OAI211_X1 U2751 ( .C1(n387), .C2(n1666), .A(n4286), .B(n4285), .ZN(n17872)
         );
  INV_X1 U2752 ( .A(n17939), .ZN(n519) );
  AND2_X1 U2753 ( .A1(n17008), .A2(n2827), .ZN(n17715) );
  INV_X1 U2754 ( .A(n17667), .ZN(n824) );
  OR2_X1 U2755 ( .A1(n2819), .A2(n17710), .ZN(n1363) );
  INV_X1 U2758 ( .A(n18402), .ZN(n521) );
  INV_X1 U2759 ( .A(n18236), .ZN(n522) );
  OAI21_X1 U2760 ( .B1(n17467), .B2(n4246), .A(n1481), .ZN(n16674) );
  INV_X1 U2761 ( .A(n18178), .ZN(n523) );
  AND3_X1 U2762 ( .A1(n4900), .A2(n4901), .A3(n16700), .ZN(n5814) );
  OAI21_X1 U2763 ( .B1(n422), .B2(n16782), .A(n16781), .ZN(n17902) );
  INV_X1 U2764 ( .A(n17941), .ZN(n525) );
  NAND3_X1 U2767 ( .A1(n1387), .A2(n17436), .A3(n16828), .ZN(n19560) );
  AND2_X1 U2768 ( .A1(n1253), .A2(n1252), .ZN(n17292) );
  OR2_X1 U2770 ( .A1(n16906), .A2(n17566), .ZN(n15892) );
  OR2_X1 U2771 ( .A1(n16787), .A2(n2826), .ZN(n1226) );
  AND2_X1 U2772 ( .A1(n29513), .A2(n17570), .ZN(n17318) );
  OR2_X1 U2773 ( .A1(n17361), .A2(n17365), .ZN(n15717) );
  NOR3_X1 U2774 ( .A1(n17512), .A2(n4273), .A3(n17830), .ZN(n4272) );
  INV_X1 U2776 ( .A(n6465), .ZN(n1181) );
  INV_X1 U2777 ( .A(n16883), .ZN(n17526) );
  AND2_X1 U2779 ( .A1(n17467), .A2(n4246), .ZN(n784) );
  OR2_X1 U2780 ( .A1(n16543), .A2(n17120), .ZN(n17462) );
  OR2_X1 U2781 ( .A1(n2768), .A2(n17229), .ZN(n1307) );
  NOR2_X1 U2782 ( .A1(n17279), .A2(n17278), .ZN(n779) );
  AND2_X1 U2784 ( .A1(n2122), .A2(n17552), .ZN(n17051) );
  XNOR2_X1 U2785 ( .A(n16402), .B(n16403), .ZN(n16883) );
  OR2_X1 U2786 ( .A1(n17396), .A2(n14871), .ZN(n16825) );
  INV_X1 U2787 ( .A(n17262), .ZN(n1657) );
  NOR2_X1 U2789 ( .A1(n424), .A2(n16879), .ZN(n17384) );
  INV_X1 U2790 ( .A(n4246), .ZN(n528) );
  OR2_X1 U2791 ( .A1(n17293), .A2(n17393), .ZN(n1253) );
  OR2_X1 U2793 ( .A1(n17830), .A2(n17829), .ZN(n16547) );
  AOI21_X1 U2795 ( .B1(n29559), .B2(n1466), .A(n16860), .ZN(n1465) );
  AND2_X1 U2796 ( .A1(n17569), .A2(n29138), .ZN(n4317) );
  NOR2_X1 U2797 ( .A1(n17229), .A2(n17569), .ZN(n1507) );
  INV_X1 U2798 ( .A(n17106), .ZN(n796) );
  INV_X1 U2801 ( .A(n6002), .ZN(n16790) );
  AND3_X1 U2802 ( .A1(n17275), .A2(n17277), .A3(n17276), .ZN(n780) );
  AOI21_X1 U2803 ( .B1(n29737), .B2(n1482), .A(n17464), .ZN(n17094) );
  OR2_X1 U2804 ( .A1(n17258), .A2(n1438), .ZN(n1437) );
  OR2_X1 U2805 ( .A1(n16541), .A2(n16810), .ZN(n16543) );
  OR2_X1 U2807 ( .A1(n4316), .A2(n17566), .ZN(n6417) );
  INV_X1 U2808 ( .A(n17437), .ZN(n529) );
  INV_X1 U2809 ( .A(n17396), .ZN(n17294) );
  INV_X1 U2811 ( .A(n17528), .ZN(n17158) );
  INV_X1 U2812 ( .A(n17375), .ZN(n530) );
  XNOR2_X1 U2813 ( .A(n6650), .B(n6649), .ZN(n17542) );
  INV_X1 U2818 ( .A(n16706), .ZN(n531) );
  BUF_X1 U2820 ( .A(n16736), .Z(n17488) );
  INV_X1 U2821 ( .A(n17315), .ZN(n532) );
  XNOR2_X1 U2826 ( .A(n16507), .B(n16508), .ZN(n17452) );
  INV_X1 U2827 ( .A(n17277), .ZN(n17001) );
  INV_X1 U2828 ( .A(n17124), .ZN(n1816) );
  INV_X1 U2829 ( .A(n17467), .ZN(n1482) );
  CLKBUF_X1 U2832 ( .A(n16668), .Z(n17258) );
  XNOR2_X1 U2833 ( .A(n16142), .B(n1575), .ZN(n1438) );
  XNOR2_X1 U2834 ( .A(n14914), .B(n14913), .ZN(n17397) );
  XNOR2_X1 U2835 ( .A(n15653), .B(n15652), .ZN(n17552) );
  XNOR2_X1 U2837 ( .A(n16420), .B(n16419), .ZN(n17528) );
  INV_X1 U2838 ( .A(n17393), .ZN(n533) );
  INV_X1 U2840 ( .A(n16803), .ZN(n534) );
  INV_X1 U2841 ( .A(n15731), .ZN(n535) );
  XNOR2_X1 U2843 ( .A(n16064), .B(n16063), .ZN(n17097) );
  INV_X1 U2844 ( .A(n17062), .ZN(n536) );
  XNOR2_X1 U2846 ( .A(n15564), .B(n6929), .ZN(n16937) );
  XNOR2_X1 U2847 ( .A(n1778), .B(n1348), .ZN(n17356) );
  XNOR2_X1 U2849 ( .A(n15794), .B(n15793), .ZN(n17545) );
  XNOR2_X1 U2851 ( .A(n6160), .B(n6158), .ZN(n17137) );
  XNOR2_X1 U2852 ( .A(n15778), .B(n15777), .ZN(n6649) );
  XNOR2_X1 U2854 ( .A(n16163), .B(n16164), .ZN(n17463) );
  INV_X1 U2857 ( .A(n29632), .ZN(n542) );
  XNOR2_X1 U2858 ( .A(n16434), .B(n4323), .ZN(n16050) );
  XNOR2_X1 U2859 ( .A(n15982), .B(n15940), .ZN(n16201) );
  XNOR2_X1 U2860 ( .A(n16233), .B(n1259), .ZN(n1258) );
  XNOR2_X1 U2861 ( .A(n14719), .B(n16422), .ZN(n16145) );
  INV_X1 U2862 ( .A(n16278), .ZN(n16281) );
  XNOR2_X1 U2863 ( .A(n1310), .B(n15668), .ZN(n16278) );
  NAND2_X1 U2864 ( .A1(n14866), .A2(n4324), .ZN(n4323) );
  INV_X1 U2865 ( .A(n16232), .ZN(n769) );
  XNOR2_X1 U2867 ( .A(n15900), .B(n16023), .ZN(n16302) );
  AND2_X1 U2868 ( .A1(n14800), .A2(n2190), .ZN(n15760) );
  INV_X1 U2869 ( .A(n16304), .ZN(n16131) );
  XNOR2_X1 U2870 ( .A(n16230), .B(n16090), .ZN(n1259) );
  XNOR2_X1 U2873 ( .A(n16084), .B(n2116), .ZN(n16205) );
  AND2_X1 U2874 ( .A1(n6760), .A2(n6758), .ZN(n16585) );
  NAND2_X1 U2876 ( .A1(n14911), .A2(n14910), .ZN(n16070) );
  AND3_X1 U2880 ( .A1(n6090), .A2(n6089), .A3(n6088), .ZN(n15992) );
  NOR2_X1 U2882 ( .A1(n14528), .A2(n14527), .ZN(n16024) );
  NOR2_X1 U2883 ( .A1(n2208), .A2(n2207), .ZN(n15565) );
  NAND3_X1 U2884 ( .A1(n14673), .A2(n14674), .A3(n2699), .ZN(n2700) );
  OAI21_X1 U2887 ( .B1(n4955), .B2(n4957), .A(n14110), .ZN(n16332) );
  OAI211_X1 U2889 ( .C1(n14532), .C2(n14533), .A(n14531), .B(n14530), .ZN(
        n16052) );
  OR2_X1 U2890 ( .A1(n15131), .A2(n15132), .ZN(n1597) );
  OAI211_X1 U2892 ( .C1(n14940), .C2(n15406), .A(n14939), .B(n14938), .ZN(
        n16241) );
  OAI21_X1 U2893 ( .B1(n15227), .B2(n1149), .A(n1148), .ZN(n3923) );
  OR2_X1 U2894 ( .A1(n756), .A2(n15288), .ZN(n4184) );
  INV_X1 U2895 ( .A(n16172), .ZN(n543) );
  AND2_X1 U2896 ( .A1(n14855), .A2(n14856), .ZN(n1067) );
  AND2_X1 U2897 ( .A1(n15373), .A2(n15374), .ZN(n1662) );
  OAI22_X1 U2899 ( .A1(n15353), .A2(n5238), .B1(n14191), .B2(n15228), .ZN(
        n16176) );
  INV_X1 U2901 ( .A(n15458), .ZN(n1701) );
  BUF_X1 U2902 ( .A(n14882), .Z(n14884) );
  INV_X1 U2903 ( .A(n15185), .ZN(n972) );
  MUX2_X1 U2904 ( .A(n15187), .B(n13818), .S(n15190), .Z(n13819) );
  AND2_X1 U2905 ( .A1(n15310), .A2(n15272), .ZN(n1095) );
  NAND3_X1 U2906 ( .A1(n4259), .A2(n13732), .A3(n14070), .ZN(n15373) );
  OAI21_X1 U2907 ( .B1(n14737), .B2(n15009), .A(n837), .ZN(n14738) );
  OAI211_X1 U2909 ( .C1(n15275), .C2(n15274), .A(n15514), .B(n1328), .ZN(n1518) );
  OR2_X1 U2910 ( .A1(n14220), .A2(n15047), .ZN(n3615) );
  OR2_X1 U2912 ( .A1(n15371), .A2(n15370), .ZN(n683) );
  AND2_X1 U2914 ( .A1(n15290), .A2(n15292), .ZN(n15040) );
  INV_X1 U2916 ( .A(n15115), .ZN(n544) );
  OR2_X1 U2917 ( .A1(n29380), .A2(n15394), .ZN(n1326) );
  INV_X1 U2919 ( .A(n15001), .ZN(n1745) );
  AND2_X1 U2922 ( .A1(n14835), .A2(n2456), .ZN(n2455) );
  INV_X1 U2923 ( .A(n15447), .ZN(n15322) );
  INV_X1 U2924 ( .A(n15117), .ZN(n1001) );
  INV_X1 U2925 ( .A(n15190), .ZN(n14785) );
  OR2_X1 U2926 ( .A1(n15456), .A2(n28803), .ZN(n3079) );
  INV_X1 U2928 ( .A(n15160), .ZN(n545) );
  INV_X1 U2930 ( .A(n15119), .ZN(n1005) );
  INV_X1 U2931 ( .A(n15190), .ZN(n547) );
  AND2_X1 U2933 ( .A1(n5666), .A2(n2304), .ZN(n15155) );
  INV_X1 U2936 ( .A(n15444), .ZN(n548) );
  AND2_X1 U2939 ( .A1(n14550), .A2(n14549), .ZN(n1809) );
  NAND3_X1 U2941 ( .A1(n14441), .A2(n14442), .A3(n14443), .ZN(n14923) );
  INV_X1 U2942 ( .A(n15127), .ZN(n1744) );
  INV_X1 U2945 ( .A(n15102), .ZN(n549) );
  BUF_X1 U2946 ( .A(n14153), .Z(n15360) );
  AND3_X1 U2947 ( .A1(n14904), .A2(n14905), .A3(n14906), .ZN(n14908) );
  INV_X1 U2948 ( .A(n15152), .ZN(n5198) );
  INV_X1 U2949 ( .A(n15222), .ZN(n550) );
  INV_X1 U2950 ( .A(n15123), .ZN(n551) );
  NAND4_X1 U2952 ( .A1(n4435), .A2(n4432), .A3(n13688), .A4(n4431), .ZN(n14992) );
  AOI21_X1 U2953 ( .B1(n13773), .B2(n13774), .A(n13772), .ZN(n14963) );
  AND2_X1 U2956 ( .A1(n1628), .A2(n1629), .ZN(n1627) );
  OAI21_X1 U2957 ( .B1(n13793), .B2(n13217), .A(n13216), .ZN(n15085) );
  INV_X1 U2958 ( .A(n15182), .ZN(n552) );
  OR2_X1 U2960 ( .A1(n13797), .A2(n13796), .ZN(n1569) );
  AND2_X1 U2962 ( .A1(n13709), .A2(n13708), .ZN(n15246) );
  BUF_X1 U2963 ( .A(n14115), .Z(n15248) );
  NAND2_X1 U2964 ( .A1(n14139), .A2(n14140), .ZN(n4992) );
  OAI21_X1 U2966 ( .B1(n14770), .B2(n14771), .A(n14769), .ZN(n14713) );
  INV_X1 U2967 ( .A(n15456), .ZN(n553) );
  AOI21_X1 U2970 ( .B1(n830), .B2(n14273), .A(n4666), .ZN(n15513) );
  OAI21_X1 U2971 ( .B1(n815), .B2(n13903), .A(n814), .ZN(n13904) );
  NOR2_X1 U2972 ( .A1(n13751), .A2(n13750), .ZN(n15151) );
  OR2_X1 U2976 ( .A1(n4074), .A2(n14168), .ZN(n998) );
  OR2_X1 U2977 ( .A1(n5409), .A2(n14437), .ZN(n727) );
  OR2_X1 U2979 ( .A1(n4837), .A2(n28986), .ZN(n5015) );
  INV_X1 U2982 ( .A(n4666), .ZN(n829) );
  AND2_X1 U2984 ( .A1(n11372), .A2(n1580), .ZN(n1776) );
  NAND3_X1 U2988 ( .A1(n14429), .A2(n14428), .A3(n28199), .ZN(n14430) );
  INV_X1 U2989 ( .A(n4893), .ZN(n14355) );
  CLKBUF_X1 U2990 ( .A(n13257), .Z(n14320) );
  AND2_X1 U2991 ( .A1(n14244), .A2(n28172), .ZN(n956) );
  AOI21_X1 U2992 ( .B1(n13903), .B2(n389), .A(n1661), .ZN(n1660) );
  OR2_X1 U2993 ( .A1(n1320), .A2(n14452), .ZN(n1322) );
  BUF_X1 U2994 ( .A(n13775), .Z(n14250) );
  INV_X1 U2995 ( .A(n1742), .ZN(n13614) );
  INV_X1 U2996 ( .A(n28804), .ZN(n4012) );
  AND2_X1 U2997 ( .A1(n29589), .A2(n4425), .ZN(n815) );
  OR2_X1 U2998 ( .A1(n13999), .A2(n14038), .ZN(n1016) );
  AND2_X1 U2999 ( .A1(n14480), .A2(n13936), .ZN(n644) );
  XNOR2_X1 U3002 ( .A(n13225), .B(n4041), .ZN(n14043) );
  INV_X1 U3003 ( .A(n13595), .ZN(n14146) );
  INV_X1 U3004 ( .A(n13716), .ZN(n13903) );
  INV_X1 U3005 ( .A(n14158), .ZN(n14474) );
  AND2_X1 U3006 ( .A1(n29589), .A2(n13902), .ZN(n1661) );
  OR3_X1 U3007 ( .A1(n14285), .A2(n14083), .A3(n14084), .ZN(n14283) );
  INV_X1 U3008 ( .A(n14217), .ZN(n555) );
  INV_X1 U3011 ( .A(n14322), .ZN(n1346) );
  INV_X1 U3013 ( .A(n14327), .ZN(n14323) );
  INV_X1 U3014 ( .A(n5531), .ZN(n6351) );
  AND2_X1 U3015 ( .A1(n14593), .A2(n14101), .ZN(n12938) );
  XNOR2_X1 U3016 ( .A(n13276), .B(n13275), .ZN(n14053) );
  INV_X1 U3017 ( .A(n13837), .ZN(n556) );
  INV_X1 U3018 ( .A(n14381), .ZN(n557) );
  INV_X1 U3019 ( .A(n14479), .ZN(n558) );
  XNOR2_X1 U3020 ( .A(n12526), .B(n12525), .ZN(n13874) );
  XNOR2_X1 U3021 ( .A(n13041), .B(n1956), .ZN(n14126) );
  INV_X1 U3022 ( .A(n14122), .ZN(n559) );
  XNOR2_X1 U3023 ( .A(n12710), .B(n12709), .ZN(n14200) );
  INV_X1 U3024 ( .A(n14309), .ZN(n560) );
  XNOR2_X1 U3025 ( .A(n3624), .B(n13011), .ZN(n4166) );
  INV_X1 U3026 ( .A(n1368), .ZN(n13901) );
  INV_X1 U3027 ( .A(n14083), .ZN(n561) );
  XNOR2_X1 U3029 ( .A(n13498), .B(n13499), .ZN(n13589) );
  XNOR2_X1 U3030 ( .A(n11370), .B(n11369), .ZN(n14101) );
  INV_X1 U3032 ( .A(n14435), .ZN(n562) );
  XNOR2_X1 U3033 ( .A(n12439), .B(n12438), .ZN(n14399) );
  XNOR2_X1 U3035 ( .A(n13367), .B(n13368), .ZN(n13716) );
  XNOR2_X1 U3038 ( .A(n12821), .B(n12820), .ZN(n13953) );
  XNOR2_X1 U3039 ( .A(n12694), .B(n12695), .ZN(n14455) );
  INV_X1 U3040 ( .A(n14238), .ZN(n563) );
  XNOR2_X1 U3041 ( .A(n13268), .B(n13267), .ZN(n13816) );
  XNOR2_X1 U3042 ( .A(n11410), .B(n3687), .ZN(n13943) );
  XNOR2_X1 U3043 ( .A(n12873), .B(n12874), .ZN(n12878) );
  XNOR2_X1 U3045 ( .A(n12832), .B(n12829), .ZN(n1085) );
  XNOR2_X1 U3046 ( .A(n12901), .B(n1780), .ZN(n12902) );
  INV_X1 U3047 ( .A(n14123), .ZN(n564) );
  XNOR2_X1 U3049 ( .A(n12884), .B(n12885), .ZN(n4041) );
  XNOR2_X1 U3051 ( .A(n13101), .B(n13348), .ZN(n13246) );
  INV_X1 U3052 ( .A(n12461), .ZN(n13298) );
  XNOR2_X1 U3053 ( .A(n12504), .B(n12813), .ZN(n13521) );
  AND2_X1 U3054 ( .A1(n5468), .A2(n5467), .ZN(n13227) );
  XNOR2_X1 U3055 ( .A(n13297), .B(n1664), .ZN(n13501) );
  OR2_X1 U3057 ( .A1(n6645), .A2(n15576), .ZN(n961) );
  INV_X1 U3058 ( .A(n6645), .ZN(n962) );
  XNOR2_X1 U3059 ( .A(n12799), .B(n1293), .ZN(n13346) );
  NOR2_X1 U3060 ( .A1(n11407), .A2(n5076), .ZN(n12747) );
  NAND2_X1 U3061 ( .A1(n11931), .A2(n1491), .ZN(n1293) );
  BUF_X1 U3065 ( .A(n12608), .Z(n13359) );
  AND2_X1 U3066 ( .A1(n4017), .A2(n11956), .ZN(n860) );
  NAND3_X1 U3067 ( .A1(n2604), .A2(n12002), .A3(n2603), .ZN(n12879) );
  AND2_X1 U3068 ( .A1(n4102), .A2(n12130), .ZN(n13538) );
  INV_X1 U3071 ( .A(n12529), .ZN(n565) );
  OAI211_X1 U3077 ( .C1(n12256), .C2(n11598), .A(n11597), .B(n11596), .ZN(
        n13504) );
  NAND2_X1 U3078 ( .A1(n11691), .A2(n11690), .ZN(n13043) );
  AND4_X1 U3079 ( .A1(n10955), .A2(n10954), .A3(n10953), .A4(n10952), .ZN(
        n13069) );
  OR2_X1 U3082 ( .A1(n12280), .A2(n4105), .ZN(n12284) );
  OR2_X1 U3090 ( .A1(n12103), .A2(n12164), .ZN(n705) );
  OR2_X1 U3091 ( .A1(n375), .A2(n776), .ZN(n11541) );
  OR2_X1 U3092 ( .A1(n12027), .A2(n1291), .ZN(n1107) );
  AOI22_X1 U3093 ( .A1(n11862), .A2(n11861), .B1(n11860), .B2(n11947), .ZN(
        n1526) );
  INV_X1 U3094 ( .A(n12288), .ZN(n1103) );
  INV_X1 U3095 ( .A(n11844), .ZN(n706) );
  OAI21_X1 U3096 ( .B1(n12177), .B2(n11413), .A(n11412), .ZN(n12788) );
  AND2_X1 U3097 ( .A1(n1484), .A2(n11715), .ZN(n11650) );
  OR2_X1 U3099 ( .A1(n11703), .A2(n12205), .ZN(n11439) );
  AND2_X1 U3101 ( .A1(n13086), .A2(n13081), .ZN(n11812) );
  INV_X1 U3103 ( .A(n9692), .ZN(n12210) );
  INV_X1 U3104 ( .A(n11648), .ZN(n1706) );
  OR2_X1 U3105 ( .A1(n11417), .A2(n11648), .ZN(n11714) );
  AND2_X1 U3106 ( .A1(n12354), .A2(n12352), .ZN(n1371) );
  CLKBUF_X1 U3107 ( .A(n12293), .Z(n12061) );
  OR2_X1 U3108 ( .A1(n1890), .A2(n12177), .ZN(n1318) );
  INV_X1 U3109 ( .A(n12508), .ZN(n1746) );
  INV_X1 U3110 ( .A(n11505), .ZN(n12280) );
  INV_X1 U3111 ( .A(n12315), .ZN(n566) );
  INV_X1 U3113 ( .A(n11551), .ZN(n1453) );
  INV_X1 U3115 ( .A(n11867), .ZN(n11360) );
  OR2_X1 U3117 ( .A1(n5905), .A2(n10935), .ZN(n11947) );
  OAI21_X1 U3118 ( .B1(n10911), .B2(n10452), .A(n10451), .ZN(n11876) );
  INV_X1 U3119 ( .A(n11852), .ZN(n11547) );
  INV_X1 U3122 ( .A(n11715), .ZN(n1485) );
  NOR2_X1 U3123 ( .A1(n12337), .A2(n11473), .ZN(n1292) );
  INV_X1 U3128 ( .A(n12266), .ZN(n568) );
  AND2_X1 U3129 ( .A1(n12508), .A2(n12507), .ZN(n11616) );
  OR2_X1 U3130 ( .A1(n11980), .A2(n12226), .ZN(n11981) );
  AND4_X2 U3132 ( .A1(n10107), .A2(n10104), .A3(n10106), .A4(n10105), .ZN(
        n12508) );
  AOI22_X1 U3133 ( .A1(n11107), .A2(n11106), .B1(n11217), .B2(n11105), .ZN(
        n12577) );
  OAI21_X1 U3135 ( .B1(n11143), .B2(n11142), .A(n1452), .ZN(n11780) );
  NAND2_X1 U3137 ( .A1(n6720), .A2(n3570), .ZN(n11969) );
  INV_X1 U3139 ( .A(n12181), .ZN(n570) );
  INV_X1 U3142 ( .A(n12132), .ZN(n12265) );
  INV_X1 U3144 ( .A(n11536), .ZN(n572) );
  INV_X1 U3145 ( .A(n12146), .ZN(n573) );
  INV_X1 U3146 ( .A(n11855), .ZN(n574) );
  INV_X1 U3148 ( .A(n11574), .ZN(n575) );
  INV_X1 U3150 ( .A(n10863), .ZN(n577) );
  INV_X1 U3152 ( .A(n12050), .ZN(n12316) );
  OAI211_X1 U3153 ( .C1(n10844), .C2(n10523), .A(n11039), .B(n4145), .ZN(
        n12328) );
  OR2_X1 U3155 ( .A1(n10542), .A2(n10541), .ZN(n989) );
  OAI211_X1 U3156 ( .C1(n1975), .C2(n2143), .A(n1399), .B(n1400), .ZN(n12163)
         );
  AND2_X1 U3157 ( .A1(n10755), .A2(n10756), .ZN(n11672) );
  INV_X1 U3159 ( .A(n11463), .ZN(n578) );
  INV_X1 U3160 ( .A(n11856), .ZN(n579) );
  AND4_X1 U3161 ( .A1(n2086), .A2(n10642), .A3(n2085), .A4(n2084), .ZN(n11962)
         );
  OR2_X1 U3162 ( .A1(n10996), .A2(n10995), .ZN(n1786) );
  NAND2_X1 U3165 ( .A1(n10652), .A2(n10884), .ZN(n1261) );
  INV_X1 U3166 ( .A(n11901), .ZN(n580) );
  OR2_X1 U3167 ( .A1(n3801), .A2(n10694), .ZN(n12194) );
  OR2_X1 U3168 ( .A1(n10963), .A2(n10956), .ZN(n3413) );
  INV_X1 U3169 ( .A(n10726), .ZN(n10928) );
  AND2_X1 U3171 ( .A1(n10893), .A2(n11290), .ZN(n1736) );
  OR2_X1 U3172 ( .A1(n11082), .A2(n11083), .ZN(n1399) );
  CLKBUF_X1 U3173 ( .A(n11323), .Z(n11328) );
  OR2_X1 U3174 ( .A1(n1703), .A2(n1338), .ZN(n10526) );
  OR2_X1 U3176 ( .A1(n10520), .A2(n10884), .ZN(n1260) );
  OR2_X1 U3177 ( .A1(n11241), .A2(n11244), .ZN(n787) );
  INV_X1 U3178 ( .A(n28624), .ZN(n1357) );
  AND2_X1 U3179 ( .A1(n11121), .A2(n11119), .ZN(n10506) );
  NOR2_X1 U3180 ( .A1(n969), .A2(n10806), .ZN(n10741) );
  INV_X1 U3181 ( .A(n11209), .ZN(n11213) );
  INV_X1 U3182 ( .A(n1338), .ZN(n1704) );
  NOR2_X1 U3183 ( .A1(n433), .A2(n11210), .ZN(n1975) );
  INV_X1 U3190 ( .A(n28407), .ZN(n10998) );
  OR2_X1 U3193 ( .A1(n11064), .A2(n11067), .ZN(n11068) );
  INV_X1 U3194 ( .A(n11199), .ZN(n581) );
  XNOR2_X1 U3195 ( .A(n10416), .B(n10415), .ZN(n11207) );
  INV_X1 U3196 ( .A(n11196), .ZN(n3585) );
  CLKBUF_X1 U3197 ( .A(n10882), .Z(n11211) );
  INV_X1 U3198 ( .A(n11064), .ZN(n11244) );
  XNOR2_X1 U3199 ( .A(n9809), .B(n9808), .ZN(n10786) );
  XNOR2_X1 U3203 ( .A(n8376), .B(n8377), .ZN(n11166) );
  INV_X1 U3204 ( .A(n10970), .ZN(n1285) );
  INV_X1 U3206 ( .A(n2690), .ZN(n11255) );
  OR2_X1 U3207 ( .A1(n11243), .A2(n11240), .ZN(n1760) );
  OR2_X1 U3208 ( .A1(n11315), .A2(n2690), .ZN(n1537) );
  CLKBUF_X1 U3209 ( .A(n10524), .Z(n11248) );
  XNOR2_X1 U3210 ( .A(n10301), .B(n10300), .ZN(n11294) );
  XNOR2_X1 U3212 ( .A(n8775), .B(n8774), .ZN(n11337) );
  INV_X1 U3213 ( .A(n11149), .ZN(n582) );
  XNOR2_X1 U3218 ( .A(n9302), .B(n9915), .ZN(n10300) );
  INV_X1 U3219 ( .A(n11282), .ZN(n584) );
  INV_X1 U3221 ( .A(n11084), .ZN(n10883) );
  INV_X1 U3222 ( .A(n1854), .ZN(n585) );
  XNOR2_X1 U3223 ( .A(n9968), .B(n9967), .ZN(n10502) );
  XNOR2_X1 U3224 ( .A(n8620), .B(n8621), .ZN(n11196) );
  INV_X1 U3225 ( .A(n11033), .ZN(n586) );
  INV_X1 U3227 ( .A(n11093), .ZN(n587) );
  XNOR2_X1 U3229 ( .A(n9720), .B(n9719), .ZN(n11226) );
  INV_X1 U3231 ( .A(n10930), .ZN(n588) );
  INV_X1 U3232 ( .A(n10984), .ZN(n589) );
  XNOR2_X1 U3234 ( .A(n10389), .B(n10390), .ZN(n11094) );
  INV_X1 U3235 ( .A(n10932), .ZN(n590) );
  XNOR2_X1 U3236 ( .A(n10213), .B(n10214), .ZN(n11066) );
  INV_X1 U3237 ( .A(n10976), .ZN(n591) );
  XNOR2_X1 U3238 ( .A(n1761), .B(n10187), .ZN(n11243) );
  XNOR2_X1 U3241 ( .A(n9629), .B(n9379), .ZN(n9721) );
  INV_X1 U3243 ( .A(n10752), .ZN(n593) );
  INV_X1 U3244 ( .A(n11253), .ZN(n594) );
  INV_X1 U3246 ( .A(n11084), .ZN(n595) );
  XNOR2_X1 U3249 ( .A(n654), .B(n10207), .ZN(n9590) );
  XNOR2_X1 U3250 ( .A(n10322), .B(n9295), .ZN(n9977) );
  XNOR2_X1 U3251 ( .A(n655), .B(n10310), .ZN(n9956) );
  AND2_X1 U3253 ( .A1(n2596), .A2(n2597), .ZN(n10228) );
  XNOR2_X1 U3256 ( .A(n4479), .B(n10353), .ZN(n10433) );
  OR2_X1 U3257 ( .A1(n8606), .A2(n963), .ZN(n10246) );
  INV_X1 U3259 ( .A(n9648), .ZN(n9900) );
  XNOR2_X1 U3262 ( .A(n9696), .B(n10171), .ZN(n9596) );
  AND2_X1 U3269 ( .A1(n2290), .A2(n5330), .ZN(n10359) );
  XNOR2_X1 U3271 ( .A(n9426), .B(n10357), .ZN(n9722) );
  INV_X1 U3273 ( .A(n9505), .ZN(n654) );
  AND2_X1 U3275 ( .A1(n10233), .A2(n8724), .ZN(n8606) );
  AND2_X1 U3277 ( .A1(n843), .A2(n842), .ZN(n10064) );
  NAND4_X1 U3281 ( .A1(n4728), .A2(n8689), .A3(n8690), .A4(n9024), .ZN(n9899)
         );
  OR2_X1 U3285 ( .A1(n7575), .A2(n8537), .ZN(n1355) );
  OAI21_X1 U3288 ( .B1(n970), .B2(n8355), .A(n8354), .ZN(n971) );
  NAND4_X1 U3290 ( .A1(n9049), .A2(n4730), .A3(n4731), .A4(n8691), .ZN(n10227)
         );
  NAND3_X1 U3292 ( .A1(n8417), .A2(n8416), .A3(n8415), .ZN(n10073) );
  OR2_X1 U3293 ( .A1(n7575), .A2(n8537), .ZN(n1416) );
  MUX2_X1 U3294 ( .A(n8960), .B(n8959), .S(n8958), .Z(n9613) );
  OAI21_X1 U3295 ( .B1(n744), .B2(n8120), .A(n5449), .ZN(n9992) );
  OAI22_X1 U3296 ( .A1(n9340), .A2(n8755), .B1(n1934), .B2(n8754), .ZN(n8756)
         );
  MUX2_X1 U3297 ( .A(n7001), .B(n7000), .S(n9045), .Z(n9732) );
  INV_X1 U3298 ( .A(n8993), .ZN(n1047) );
  AND3_X1 U3299 ( .A1(n2861), .A2(n2860), .A3(n2863), .ZN(n10302) );
  OR2_X1 U3300 ( .A1(n8483), .A2(n440), .ZN(n1710) );
  OR2_X1 U3301 ( .A1(n1788), .A2(n8760), .ZN(n1790) );
  OAI21_X1 U3302 ( .B1(n8426), .B2(n8427), .A(n8078), .ZN(n8120) );
  OR2_X1 U3305 ( .A1(n9049), .A2(n9235), .ZN(n1117) );
  NOR2_X1 U3306 ( .A1(n844), .A2(n9137), .ZN(n843) );
  AOI21_X1 U3307 ( .B1(n8920), .B2(n8919), .A(n8918), .ZN(n9647) );
  OR2_X1 U3308 ( .A1(n8610), .A2(n9530), .ZN(n714) );
  AND2_X1 U3310 ( .A1(n9135), .A2(n9134), .ZN(n844) );
  AND2_X1 U3311 ( .A1(n6747), .A2(n9374), .ZN(n8570) );
  NOR2_X1 U3312 ( .A1(n9140), .A2(n638), .ZN(n637) );
  OR2_X1 U3313 ( .A1(n5568), .A2(n5945), .ZN(n9238) );
  NOR2_X1 U3314 ( .A1(n8819), .A2(n8594), .ZN(n8823) );
  INV_X1 U3315 ( .A(n8058), .ZN(n8426) );
  NOR2_X1 U3316 ( .A1(n9438), .A2(n8777), .ZN(n8993) );
  OR2_X1 U3317 ( .A1(n8931), .A2(n9148), .ZN(n8761) );
  MUX2_X1 U3318 ( .A(n8661), .B(n8482), .S(n9016), .Z(n8483) );
  AND2_X1 U3319 ( .A1(n8961), .A2(n9171), .ZN(n9173) );
  OR2_X1 U3320 ( .A1(n8827), .A2(n8586), .ZN(n8465) );
  INV_X1 U3321 ( .A(n8699), .ZN(n8403) );
  OAI211_X1 U3322 ( .C1(n9140), .C2(n8562), .A(n8561), .B(n1803), .ZN(n2336)
         );
  OR2_X1 U3323 ( .A1(n1934), .A2(n9133), .ZN(n1670) );
  OR2_X1 U3324 ( .A1(n8764), .A2(n8763), .ZN(n9564) );
  OR2_X1 U3326 ( .A1(n9013), .A2(n9014), .ZN(n1615) );
  AND2_X1 U3327 ( .A1(n4938), .A2(n7091), .ZN(n1839) );
  OAI21_X1 U3328 ( .B1(n8924), .B2(n6718), .A(n1934), .ZN(n8552) );
  INV_X1 U3329 ( .A(n9037), .ZN(n1634) );
  OR2_X1 U3330 ( .A1(n8782), .A2(n9186), .ZN(n8784) );
  OR2_X1 U3331 ( .A1(n9148), .A2(n8929), .ZN(n1528) );
  OR2_X1 U3332 ( .A1(n8983), .A2(n8981), .ZN(n8408) );
  AND2_X1 U3335 ( .A1(n9125), .A2(n8899), .ZN(n1794) );
  AND2_X1 U3336 ( .A1(n8500), .A2(n8652), .ZN(n7906) );
  INV_X1 U3337 ( .A(n1910), .ZN(n8430) );
  INV_X1 U3338 ( .A(n9122), .ZN(n1793) );
  CLKBUF_X1 U3339 ( .A(n8777), .Z(n9208) );
  OAI21_X1 U3340 ( .B1(n8353), .B2(n8077), .A(n8427), .ZN(n745) );
  INV_X1 U3341 ( .A(n8963), .ZN(n9170) );
  OR2_X1 U3344 ( .A1(n8183), .A2(n8182), .ZN(n8980) );
  INV_X1 U3345 ( .A(n9144), .ZN(n638) );
  INV_X1 U3347 ( .A(n8981), .ZN(n596) );
  INV_X1 U3350 ( .A(n9228), .ZN(n597) );
  OR2_X1 U3351 ( .A1(n7476), .A2(n7475), .ZN(n8848) );
  INV_X1 U3352 ( .A(n9139), .ZN(n598) );
  INV_X1 U3353 ( .A(n8562), .ZN(n599) );
  AOI21_X1 U3355 ( .B1(n1586), .B2(n1587), .A(n1589), .ZN(n8326) );
  INV_X1 U3356 ( .A(n8792), .ZN(n9035) );
  INV_X1 U3357 ( .A(n9132), .ZN(n600) );
  INV_X1 U3358 ( .A(n9134), .ZN(n601) );
  INV_X1 U3360 ( .A(n8977), .ZN(n602) );
  OAI211_X1 U3362 ( .C1(n7725), .C2(n8043), .A(n7724), .B(n7723), .ZN(n9007)
         );
  INV_X1 U3363 ( .A(n8579), .ZN(n603) );
  INV_X1 U3365 ( .A(n9171), .ZN(n605) );
  OR2_X1 U3368 ( .A1(n7217), .A2(n742), .ZN(n3301) );
  OAI21_X1 U3369 ( .B1(n5911), .B2(n8247), .A(n5910), .ZN(n8966) );
  NAND3_X1 U3370 ( .A1(n1352), .A2(n1351), .A3(n1349), .ZN(n8384) );
  INV_X1 U3371 ( .A(n9421), .ZN(n606) );
  INV_X1 U3373 ( .A(n1589), .ZN(n1585) );
  OR2_X1 U3374 ( .A1(n7317), .A2(n7775), .ZN(n1586) );
  INV_X1 U3375 ( .A(n8819), .ZN(n607) );
  AOI21_X1 U3376 ( .B1(n1568), .B2(n5256), .A(n5255), .ZN(n7973) );
  INV_X1 U3377 ( .A(n9016), .ZN(n608) );
  NAND4_X1 U3378 ( .A1(n7182), .A2(n7183), .A3(n7181), .A4(n7180), .ZN(n8733)
         );
  OAI211_X1 U3380 ( .C1(n7704), .C2(n7840), .A(n7702), .B(n7703), .ZN(n8792)
         );
  AOI22_X1 U3382 ( .A1(n7209), .A2(n7208), .B1(n7207), .B2(n7206), .ZN(n8525)
         );
  OR2_X1 U3383 ( .A1(n7766), .A2(n4856), .ZN(n4855) );
  AOI22_X1 U3385 ( .A1(n8052), .A2(n8132), .B1(n8051), .B2(n8050), .ZN(n9363)
         );
  INV_X1 U3386 ( .A(n9396), .ZN(n609) );
  OR2_X1 U3390 ( .A1(n7385), .A2(n6748), .ZN(n9374) );
  NOR2_X1 U3391 ( .A1(n7316), .A2(n1700), .ZN(n1589) );
  INV_X1 U3392 ( .A(n3654), .ZN(n771) );
  AND3_X1 U3393 ( .A1(n7381), .A2(n7380), .A3(n7379), .ZN(n8929) );
  OAI21_X1 U3394 ( .B1(n7864), .B2(n7172), .A(n5149), .ZN(n5148) );
  AND2_X1 U3395 ( .A1(n7290), .A2(n7759), .ZN(n2630) );
  OR2_X1 U3396 ( .A1(n8260), .A2(n28614), .ZN(n1198) );
  AND2_X1 U3398 ( .A1(n8044), .A2(n7722), .ZN(n889) );
  INV_X1 U3399 ( .A(n1354), .ZN(n1350) );
  BUF_X1 U3400 ( .A(n7399), .Z(n8304) );
  BUF_X1 U3401 ( .A(n7400), .Z(n8305) );
  AND2_X1 U3404 ( .A1(n7368), .A2(n439), .ZN(n1295) );
  OR2_X1 U3405 ( .A1(n7456), .A2(n7040), .ZN(n7645) );
  OR2_X1 U3406 ( .A1(n7793), .A2(n7150), .ZN(n2545) );
  INV_X1 U3407 ( .A(n7283), .ZN(n8150) );
  INV_X1 U3409 ( .A(n7742), .ZN(n7744) );
  BUF_X1 U3410 ( .A(n7283), .Z(n7542) );
  INV_X1 U3411 ( .A(n7793), .ZN(n3810) );
  CLKBUF_X1 U3413 ( .A(n7405), .Z(n8276) );
  INV_X1 U3415 ( .A(n2804), .ZN(n1911) );
  INV_X1 U3416 ( .A(n7456), .ZN(n612) );
  XNOR2_X1 U3417 ( .A(n7038), .B(Key[154]), .ZN(n7641) );
  INV_X1 U3418 ( .A(n7349), .ZN(n8168) );
  INV_X1 U3419 ( .A(n27742), .ZN(n5633) );
  BUF_X1 U3421 ( .A(n7488), .Z(n8264) );
  INV_X1 U3422 ( .A(n8173), .ZN(n613) );
  INV_X1 U3423 ( .A(n3083), .ZN(n653) );
  BUF_X1 U3424 ( .A(n7082), .Z(n7303) );
  XNOR2_X1 U3425 ( .A(n7109), .B(Key[190]), .ZN(n7897) );
  INV_X1 U3428 ( .A(n2511), .ZN(n1782) );
  INV_X1 U3429 ( .A(n7164), .ZN(n614) );
  INV_X1 U3430 ( .A(n7089), .ZN(n1354) );
  CLKBUF_X1 U3431 ( .A(n7466), .Z(n7946) );
  CLKBUF_X1 U3432 ( .A(n7589), .Z(n7960) );
  INV_X1 U3433 ( .A(n8131), .ZN(n615) );
  INV_X1 U3434 ( .A(n3482), .ZN(n1412) );
  INV_X1 U3436 ( .A(n7839), .ZN(n7367) );
  INV_X1 U3437 ( .A(n7817), .ZN(n616) );
  XNOR2_X1 U3438 ( .A(n7154), .B(Key[30]), .ZN(n7348) );
  INV_X1 U3439 ( .A(n3752), .ZN(n1229) );
  INV_X1 U3441 ( .A(n2350), .ZN(n927) );
  CLKBUF_X1 U3442 ( .A(n7150), .Z(n7541) );
  INV_X1 U3443 ( .A(n7250), .ZN(n617) );
  XNOR2_X1 U3444 ( .A(n6996), .B(Key[121]), .ZN(n7912) );
  INV_X1 U3445 ( .A(n7268), .ZN(n618) );
  CLKBUF_X1 U3447 ( .A(Key[73]), .Z(n2523) );
  CLKBUF_X1 U3448 ( .A(Key[83]), .Z(n27452) );
  XNOR2_X1 U3452 ( .A(Key[77]), .B(Plaintext[77]), .ZN(n7851) );
  CLKBUF_X1 U3453 ( .A(Key[180]), .Z(n2987) );
  CLKBUF_X1 U3454 ( .A(Key[187]), .Z(n26825) );
  INV_X1 U3455 ( .A(n7836), .ZN(n619) );
  INV_X1 U3457 ( .A(Plaintext[25]), .ZN(n1609) );
  INV_X1 U3458 ( .A(n3219), .ZN(n621) );
  INV_X1 U3459 ( .A(n1179), .ZN(n622) );
  CLKBUF_X1 U3460 ( .A(Key[68]), .Z(n26680) );
  CLKBUF_X1 U3461 ( .A(Key[129]), .Z(n3276) );
  INV_X1 U3464 ( .A(n3751), .ZN(n623) );
  CLKBUF_X1 U3468 ( .A(Key[139]), .Z(n3501) );
  CLKBUF_X1 U3469 ( .A(Key[48]), .Z(n3650) );
  INV_X1 U3470 ( .A(n3528), .ZN(n625) );
  INV_X1 U3471 ( .A(n7924), .ZN(n626) );
  INV_X1 U3472 ( .A(n7626), .ZN(n627) );
  INV_X1 U3473 ( .A(n3686), .ZN(n628) );
  CLKBUF_X1 U3474 ( .A(Key[32]), .Z(n3003) );
  INV_X1 U3475 ( .A(n3697), .ZN(n629) );
  CLKBUF_X1 U3479 ( .A(Key[98]), .Z(n3666) );
  INV_X1 U3480 ( .A(n26665), .ZN(n630) );
  INV_X1 U3481 ( .A(n8269), .ZN(n631) );
  CLKBUF_X1 U3482 ( .A(Key[182]), .Z(n3710) );
  CLKBUF_X1 U3487 ( .A(Key[130]), .Z(n26032) );
  CLKBUF_X1 U3489 ( .A(Key[119]), .Z(n27298) );
  INV_X1 U3490 ( .A(n3423), .ZN(n632) );
  CLKBUF_X1 U3491 ( .A(Key[91]), .Z(n3134) );
  INV_X1 U3492 ( .A(n3742), .ZN(n633) );
  INV_X1 U3494 ( .A(n1175), .ZN(n634) );
  INV_X1 U3495 ( .A(n2325), .ZN(n635) );
  NAND2_X1 U3498 ( .A1(n9140), .A2(n638), .ZN(n2928) );
  NAND2_X1 U3499 ( .A1(n8561), .A2(n636), .ZN(n8567) );
  NOR2_X1 U3500 ( .A1(n9140), .A2(n599), .ZN(n636) );
  NAND2_X1 U3501 ( .A1(n599), .A2(n637), .ZN(n8189) );
  NAND2_X1 U3503 ( .A1(n641), .A2(n28391), .ZN(n23048) );
  OAI21_X1 U3504 ( .B1(n641), .B2(n23470), .A(n23469), .ZN(n23471) );
  INV_X1 U3505 ( .A(n640), .ZN(n639) );
  OAI211_X1 U3506 ( .C1(n661), .C2(n641), .A(n23193), .B(n640), .ZN(n660) );
  NAND2_X1 U3508 ( .A1(n14474), .A2(n644), .ZN(n643) );
  XNOR2_X2 U3509 ( .A(n11735), .B(n11734), .ZN(n14158) );
  NAND2_X1 U3510 ( .A1(n13934), .A2(n14480), .ZN(n646) );
  NAND3_X1 U3511 ( .A1(n21410), .A2(n21408), .A3(n21412), .ZN(n647) );
  NAND3_X1 U3513 ( .A1(n20663), .A2(n21047), .A3(n4937), .ZN(n648) );
  NAND2_X1 U3514 ( .A1(n490), .A2(n651), .ZN(n650) );
  NOR2_X1 U3515 ( .A1(n21171), .A2(n21047), .ZN(n651) );
  NAND2_X1 U3517 ( .A1(n652), .A2(n10523), .ZN(n11041) );
  XNOR2_X1 U3520 ( .A(n654), .B(n9941), .ZN(n8835) );
  XNOR2_X1 U3521 ( .A(n654), .B(n10271), .ZN(n10274) );
  OAI21_X2 U3522 ( .B1(n8983), .B2(n8411), .A(n8410), .ZN(n655) );
  XNOR2_X1 U3523 ( .A(n655), .B(n1187), .ZN(n9484) );
  XNOR2_X1 U3524 ( .A(n655), .B(n10073), .ZN(n8418) );
  XNOR2_X1 U3525 ( .A(n10272), .B(n655), .ZN(n8844) );
  XNOR2_X1 U3526 ( .A(n655), .B(n10353), .ZN(n10354) );
  NAND2_X1 U3527 ( .A1(n21143), .A2(n21117), .ZN(n21146) );
  AOI21_X1 U3528 ( .B1(n21145), .B2(n492), .A(n21119), .ZN(n657) );
  NAND2_X1 U3529 ( .A1(n657), .A2(n21141), .ZN(n656) );
  OAI21_X2 U3530 ( .B1(n19781), .B2(n20081), .A(n19780), .ZN(n21143) );
  NAND2_X1 U3531 ( .A1(n492), .A2(n20852), .ZN(n658) );
  NAND2_X1 U3533 ( .A1(n659), .A2(n21314), .ZN(n3531) );
  NAND2_X1 U3534 ( .A1(n659), .A2(n21138), .ZN(n21139) );
  NAND2_X1 U3535 ( .A1(n20723), .A2(n20724), .ZN(n659) );
  NAND2_X1 U3536 ( .A1(n24324), .A2(n24677), .ZN(n3480) );
  NAND2_X1 U3537 ( .A1(n24397), .A2(n24678), .ZN(n24324) );
  NAND3_X2 U3538 ( .A1(n660), .A2(n2046), .A3(n662), .ZN(n24678) );
  INV_X1 U3539 ( .A(n23318), .ZN(n661) );
  NAND2_X1 U3540 ( .A1(n1740), .A2(n23654), .ZN(n662) );
  NAND2_X1 U3542 ( .A1(n26734), .A2(n26995), .ZN(n663) );
  NAND2_X1 U3543 ( .A1(n29486), .A2(n25972), .ZN(n664) );
  OAI21_X1 U3544 ( .B1(n11782), .B2(n11550), .A(n11785), .ZN(n666) );
  NAND2_X1 U3546 ( .A1(n11786), .A2(n11502), .ZN(n667) );
  NAND2_X1 U3547 ( .A1(n17793), .A2(n513), .ZN(n668) );
  NAND2_X1 U3549 ( .A1(n17739), .A2(n17740), .ZN(n669) );
  NAND2_X1 U3550 ( .A1(n17738), .A2(n671), .ZN(n670) );
  NAND2_X1 U3551 ( .A1(n510), .A2(n18072), .ZN(n18076) );
  AOI21_X1 U3553 ( .B1(n24029), .B2(n24651), .A(n673), .ZN(n6664) );
  NAND2_X1 U3554 ( .A1(n3061), .A2(n629), .ZN(n672) );
  NAND3_X1 U3556 ( .A1(n24657), .A2(n24656), .A3(n673), .ZN(n24658) );
  NAND2_X1 U3557 ( .A1(n17658), .A2(n17657), .ZN(n993) );
  OR2_X1 U3559 ( .A1(n17436), .A2(n17437), .ZN(n4988) );
  NAND2_X1 U3560 ( .A1(n15489), .A2(n15485), .ZN(n5644) );
  NAND3_X1 U3561 ( .A1(n1541), .A2(n1540), .A3(n21535), .ZN(n1539) );
  NAND3_X1 U3563 ( .A1(n23271), .A2(n23272), .A3(n23273), .ZN(n674) );
  XNOR2_X1 U3564 ( .A(n675), .B(n26003), .ZN(Ciphertext[6]) );
  NAND3_X1 U3565 ( .A1(n26002), .A2(n26000), .A3(n26001), .ZN(n675) );
  NOR2_X1 U3567 ( .A1(n26180), .A2(n24204), .ZN(n25611) );
  NAND2_X1 U3568 ( .A1(n1480), .A2(n18340), .ZN(n18347) );
  NAND3_X1 U3574 ( .A1(n7765), .A2(n4855), .A3(n7764), .ZN(n1910) );
  OAI21_X1 U3575 ( .B1(n23486), .B2(n23154), .A(n23155), .ZN(n1390) );
  NAND3_X1 U3576 ( .A1(n678), .A2(n11529), .A3(n13087), .ZN(n11530) );
  NAND2_X1 U3577 ( .A1(n13084), .A2(n11980), .ZN(n678) );
  NAND2_X1 U3579 ( .A1(n16890), .A2(n17078), .ZN(n679) );
  NAND3_X1 U3580 ( .A1(n2216), .A2(n18600), .A3(n2215), .ZN(n2214) );
  NAND2_X1 U3582 ( .A1(n26817), .A2(n27025), .ZN(n26816) );
  INV_X1 U3583 ( .A(n17838), .ZN(n17839) );
  NAND2_X1 U3586 ( .A1(n17715), .A2(n17431), .ZN(n5329) );
  NAND3_X1 U3587 ( .A1(n6686), .A2(n24547), .A3(n23126), .ZN(n865) );
  NAND2_X1 U3588 ( .A1(n19938), .A2(n506), .ZN(n681) );
  NAND2_X1 U3591 ( .A1(n17663), .A2(n17947), .ZN(n757) );
  NAND3_X1 U3592 ( .A1(n17596), .A2(n686), .A3(n29024), .ZN(n17594) );
  NAND2_X1 U3595 ( .A1(n13872), .A2(n13703), .ZN(n4837) );
  OAI211_X2 U3597 ( .C1(n14884), .C2(n14585), .A(n14584), .B(n688), .ZN(n16256) );
  NAND2_X1 U3598 ( .A1(n14884), .A2(n14582), .ZN(n688) );
  INV_X1 U3599 ( .A(n690), .ZN(n689) );
  NAND2_X1 U3602 ( .A1(n691), .A2(n14275), .ZN(n14834) );
  NAND2_X1 U3603 ( .A1(n14361), .A2(n28507), .ZN(n691) );
  OAI21_X2 U3604 ( .B1(n4656), .B2(n19517), .A(n19516), .ZN(n21806) );
  NAND3_X1 U3605 ( .A1(n17416), .A2(n3234), .A3(n15811), .ZN(n17417) );
  INV_X1 U3606 ( .A(n8790), .ZN(n7606) );
  NAND2_X1 U3607 ( .A1(n8414), .A2(n8788), .ZN(n8790) );
  INV_X1 U3610 ( .A(n15047), .ZN(n694) );
  NAND2_X1 U3611 ( .A1(n15336), .A2(n15047), .ZN(n695) );
  OAI21_X1 U3612 ( .B1(n18441), .B2(n523), .A(n696), .ZN(n18098) );
  NAND2_X1 U3613 ( .A1(n18441), .A2(n18179), .ZN(n696) );
  NOR2_X2 U3614 ( .A1(n19012), .A2(n19011), .ZN(n21292) );
  NAND2_X1 U3618 ( .A1(n21090), .A2(n5817), .ZN(n20801) );
  AND2_X1 U3620 ( .A1(n20790), .A2(n20791), .ZN(n698) );
  OAI21_X1 U3621 ( .B1(n28203), .B2(n12206), .A(n1221), .ZN(n11833) );
  NAND2_X1 U3622 ( .A1(n699), .A2(n4270), .ZN(n5791) );
  NAND2_X1 U3623 ( .A1(n2296), .A2(n700), .ZN(n20789) );
  NAND2_X1 U3624 ( .A1(n20802), .A2(n701), .ZN(n700) );
  NAND2_X1 U3625 ( .A1(n20109), .A2(n20322), .ZN(n703) );
  NAND2_X1 U3626 ( .A1(n15253), .A2(n707), .ZN(n15254) );
  NAND3_X1 U3627 ( .A1(n15251), .A2(n15250), .A3(n15252), .ZN(n707) );
  NAND3_X2 U3628 ( .A1(n3765), .A2(n708), .A3(n2288), .ZN(n12760) );
  NAND3_X1 U3629 ( .A1(n1061), .A2(n12400), .A3(n11800), .ZN(n708) );
  XNOR2_X1 U3630 ( .A(n18608), .B(n19299), .ZN(n19683) );
  NOR2_X1 U3632 ( .A1(n26505), .A2(n26506), .ZN(n26638) );
  NOR2_X1 U3633 ( .A1(n24846), .A2(n709), .ZN(n24857) );
  NOR2_X1 U3634 ( .A1(n26361), .A2(n26425), .ZN(n709) );
  XNOR2_X1 U3635 ( .A(n710), .B(n21573), .ZN(n21584) );
  XNOR2_X1 U3636 ( .A(n21566), .B(n22271), .ZN(n710) );
  NAND2_X1 U3640 ( .A1(n14150), .A2(n14382), .ZN(n713) );
  XNOR2_X1 U3643 ( .A(n22315), .B(n22077), .ZN(n21341) );
  XNOR2_X1 U3644 ( .A(n22596), .B(n21325), .ZN(n22315) );
  NAND2_X1 U3645 ( .A1(n26648), .A2(n29532), .ZN(n26979) );
  NAND2_X1 U3647 ( .A1(n2708), .A2(n22084), .ZN(n1635) );
  OR2_X1 U3648 ( .A1(n7640), .A2(n612), .ZN(n983) );
  OR3_X1 U3650 ( .A1(n14380), .A2(n13837), .A3(n14381), .ZN(n6105) );
  INV_X1 U3651 ( .A(n24616), .ZN(n1262) );
  NAND2_X1 U3653 ( .A1(n16895), .A2(n16896), .ZN(n715) );
  NAND2_X1 U3656 ( .A1(n6072), .A2(n8760), .ZN(n8930) );
  INV_X1 U3657 ( .A(n15010), .ZN(n14865) );
  NAND2_X1 U3658 ( .A1(n14863), .A2(n15370), .ZN(n15010) );
  AND2_X1 U3659 ( .A1(n11308), .A2(n11053), .ZN(n10852) );
  OAI21_X1 U3660 ( .B1(n2132), .B2(n24322), .A(n24324), .ZN(n2131) );
  OAI21_X1 U3661 ( .B1(n20639), .B2(n717), .A(n20638), .ZN(n20640) );
  OAI21_X1 U3662 ( .B1(n20633), .B2(n28538), .A(n20632), .ZN(n717) );
  NAND3_X1 U3663 ( .A1(n20202), .A2(n20302), .A3(n20304), .ZN(n19948) );
  NAND2_X1 U3664 ( .A1(n719), .A2(n3717), .ZN(n3716) );
  NAND2_X1 U3665 ( .A1(n810), .A2(n3954), .ZN(n719) );
  MUX2_X2 U3666 ( .A(n24393), .B(n24394), .S(n24683), .Z(n25689) );
  NAND2_X1 U3667 ( .A1(n1744), .A2(n15004), .ZN(n14746) );
  NAND2_X1 U3668 ( .A1(n23369), .A2(n23368), .ZN(n24316) );
  NAND2_X1 U3669 ( .A1(n2508), .A2(n720), .ZN(n18667) );
  NAND3_X1 U3670 ( .A1(n1523), .A2(n18234), .A3(n1524), .ZN(n720) );
  OR2_X1 U3671 ( .A1(n5817), .A2(n21089), .ZN(n20186) );
  NAND3_X1 U3672 ( .A1(n4355), .A2(n2064), .A3(n4354), .ZN(n4353) );
  OR3_X1 U3674 ( .A1(n24140), .A2(n25009), .A3(n24139), .ZN(n2153) );
  NAND2_X1 U3675 ( .A1(n3207), .A2(n721), .ZN(n19192) );
  OAI21_X1 U3676 ( .B1(n18377), .B2(n18378), .A(n3283), .ZN(n721) );
  OAI21_X1 U3677 ( .B1(n11460), .B2(n11459), .A(n390), .ZN(n722) );
  NAND2_X1 U3678 ( .A1(n6403), .A2(n18327), .ZN(n3757) );
  NAND3_X1 U3679 ( .A1(n836), .A2(n19762), .A3(n20063), .ZN(n1699) );
  NAND2_X1 U3680 ( .A1(n18765), .A2(n19761), .ZN(n836) );
  NAND2_X1 U3683 ( .A1(n15072), .A2(n15071), .ZN(n14641) );
  NAND2_X1 U3684 ( .A1(n20553), .A2(n20406), .ZN(n20407) );
  NAND2_X1 U3686 ( .A1(n22391), .A2(n23567), .ZN(n724) );
  INV_X1 U3688 ( .A(n23567), .ZN(n726) );
  NAND3_X2 U3689 ( .A1(n728), .A2(n727), .A3(n4300), .ZN(n15389) );
  NAND2_X1 U3690 ( .A1(n3851), .A2(n14432), .ZN(n728) );
  INV_X1 U3691 ( .A(n7906), .ZN(n944) );
  XNOR2_X1 U3692 ( .A(n729), .B(n25361), .ZN(Ciphertext[10]) );
  OAI211_X1 U3693 ( .C1(n6806), .C2(n29387), .A(n3623), .B(n5359), .ZN(n729)
         );
  INV_X1 U3694 ( .A(n17844), .ZN(n17607) );
  NAND2_X1 U3695 ( .A1(n18242), .A2(n17969), .ZN(n17844) );
  NAND3_X1 U3696 ( .A1(n19837), .A2(n19750), .A3(n29143), .ZN(n5100) );
  NOR2_X1 U3697 ( .A1(n14000), .A2(n14036), .ZN(n1019) );
  INV_X1 U3698 ( .A(n22977), .ZN(n23252) );
  AOI21_X1 U3700 ( .B1(n26990), .B2(n28521), .A(n29622), .ZN(n26994) );
  NOR2_X1 U3702 ( .A1(n780), .A2(n779), .ZN(n778) );
  NOR2_X1 U3703 ( .A1(n19345), .A2(n19890), .ZN(n19369) );
  NAND2_X1 U3704 ( .A1(n14370), .A2(n731), .ZN(n5796) );
  AOI21_X1 U3705 ( .B1(n7735), .B2(n7736), .A(n7734), .ZN(n732) );
  INV_X1 U3706 ( .A(n893), .ZN(n14832) );
  NAND2_X1 U3707 ( .A1(n733), .A2(n564), .ZN(n893) );
  NAND2_X1 U3708 ( .A1(n14092), .A2(n14093), .ZN(n733) );
  NAND2_X1 U3710 ( .A1(n12928), .A2(n561), .ZN(n734) );
  NAND2_X1 U3711 ( .A1(n12927), .A2(n14083), .ZN(n735) );
  AND2_X2 U3712 ( .A1(n737), .A2(n736), .ZN(n22671) );
  NAND2_X1 U3713 ( .A1(n19460), .A2(n21717), .ZN(n736) );
  NAND2_X1 U3714 ( .A1(n738), .A2(n19461), .ZN(n737) );
  NAND2_X1 U3715 ( .A1(n19419), .A2(n19418), .ZN(n738) );
  AOI21_X1 U3717 ( .B1(n29547), .B2(n17818), .A(n18122), .ZN(n739) );
  XNOR2_X2 U3718 ( .A(n19031), .B(n19030), .ZN(n20480) );
  NAND2_X1 U3719 ( .A1(n740), .A2(n1779), .ZN(n17360) );
  NAND2_X1 U3720 ( .A1(n28793), .A2(n17356), .ZN(n740) );
  NAND2_X1 U3721 ( .A1(n28175), .A2(n28559), .ZN(n10754) );
  XNOR2_X1 U3722 ( .A(n10078), .B(n10077), .ZN(n10556) );
  NAND2_X1 U3724 ( .A1(n742), .A2(n8284), .ZN(n7673) );
  NAND2_X1 U3725 ( .A1(n742), .A2(n8280), .ZN(n7669) );
  NAND2_X1 U3726 ( .A1(n742), .A2(n8276), .ZN(n8277) );
  NAND3_X1 U3727 ( .A1(n8282), .A2(n8281), .A3(n742), .ZN(n8283) );
  NAND2_X1 U3728 ( .A1(n7215), .A2(n742), .ZN(n7216) );
  OAI21_X1 U3730 ( .B1(n743), .B2(n1485), .A(n12143), .ZN(n12148) );
  NAND2_X1 U3731 ( .A1(n573), .A2(n11712), .ZN(n743) );
  NOR2_X1 U3732 ( .A1(n1910), .A2(n745), .ZN(n744) );
  INV_X1 U3733 ( .A(n7312), .ZN(n7804) );
  NAND2_X1 U3735 ( .A1(n7804), .A2(n7898), .ZN(n746) );
  NAND2_X1 U3736 ( .A1(n7805), .A2(n7804), .ZN(n747) );
  XNOR2_X1 U3737 ( .A(n748), .B(n10228), .ZN(n9724) );
  XNOR2_X1 U3738 ( .A(n748), .B(n1895), .ZN(n9988) );
  NAND2_X1 U3740 ( .A1(n4858), .A2(n4860), .ZN(n750) );
  NAND3_X1 U3741 ( .A1(n750), .A2(n820), .A3(n3654), .ZN(n772) );
  NAND2_X1 U3742 ( .A1(n750), .A2(n820), .ZN(n1459) );
  AND2_X2 U3743 ( .A1(n751), .A2(n753), .ZN(n24369) );
  NAND2_X1 U3746 ( .A1(n23259), .A2(n23735), .ZN(n753) );
  NAND2_X1 U3747 ( .A1(n14600), .A2(n15284), .ZN(n756) );
  NAND2_X1 U3748 ( .A1(n17665), .A2(n757), .ZN(n4191) );
  INV_X1 U3749 ( .A(n7231), .ZN(n758) );
  NAND2_X1 U3750 ( .A1(n758), .A2(n7589), .ZN(n3740) );
  NAND2_X1 U3751 ( .A1(n758), .A2(n441), .ZN(n5120) );
  NAND3_X1 U3752 ( .A1(n7592), .A2(n7591), .A3(n758), .ZN(n7593) );
  NAND3_X1 U3753 ( .A1(n7873), .A2(n7957), .A3(n758), .ZN(n7054) );
  NAND3_X1 U3755 ( .A1(n10929), .A2(n762), .A3(n761), .ZN(n763) );
  NAND2_X1 U3756 ( .A1(n590), .A2(n10726), .ZN(n761) );
  NAND2_X1 U3757 ( .A1(n588), .A2(n10932), .ZN(n762) );
  XNOR2_X2 U3758 ( .A(n9474), .B(n9473), .ZN(n10726) );
  NAND2_X1 U3759 ( .A1(n765), .A2(n763), .ZN(n11878) );
  NAND2_X1 U3761 ( .A1(n10460), .A2(n10927), .ZN(n765) );
  NAND3_X1 U3762 ( .A1(n17392), .A2(n766), .A3(n5021), .ZN(n17391) );
  NAND2_X1 U3763 ( .A1(n18248), .A2(n18709), .ZN(n766) );
  NAND2_X1 U3764 ( .A1(n5023), .A2(n18706), .ZN(n17392) );
  NAND2_X1 U3765 ( .A1(n26735), .A2(n26736), .ZN(n767) );
  NAND2_X1 U3766 ( .A1(n26734), .A2(n28532), .ZN(n28100) );
  NAND3_X1 U3767 ( .A1(n2094), .A2(n26736), .A3(n29486), .ZN(n768) );
  XNOR2_X1 U3768 ( .A(n16232), .B(n622), .ZN(n14602) );
  XNOR2_X1 U3769 ( .A(n543), .B(n16232), .ZN(n15991) );
  XNOR2_X1 U3770 ( .A(n769), .B(n16400), .ZN(n15619) );
  NAND3_X1 U3771 ( .A1(n4858), .A2(n4860), .A3(n771), .ZN(n770) );
  XNOR2_X1 U3773 ( .A(n1733), .B(n19332), .ZN(n775) );
  INV_X1 U3774 ( .A(n375), .ZN(n777) );
  NAND3_X1 U3776 ( .A1(n4349), .A2(n12235), .A3(n777), .ZN(n11681) );
  NAND2_X1 U3777 ( .A1(n17274), .A2(n6465), .ZN(n781) );
  NAND2_X1 U3778 ( .A1(n17273), .A2(n1181), .ZN(n782) );
  AOI21_X1 U3779 ( .B1(n4734), .B2(n785), .A(n15462), .ZN(n15468) );
  NAND2_X1 U3781 ( .A1(n18503), .A2(n515), .ZN(n17866) );
  NAND2_X1 U3782 ( .A1(n18502), .A2(n515), .ZN(n5985) );
  OAI211_X2 U3783 ( .C1(n788), .C2(n1851), .A(n787), .B(n786), .ZN(n12050) );
  NAND2_X1 U3784 ( .A1(n11245), .A2(n11244), .ZN(n786) );
  MUX2_X1 U3785 ( .A(n1900), .B(n11240), .S(n11244), .Z(n788) );
  INV_X1 U3787 ( .A(n4220), .ZN(n790) );
  XNOR2_X2 U3788 ( .A(n15759), .B(n15758), .ZN(n4220) );
  OR2_X1 U3789 ( .A1(n14301), .A2(n13816), .ZN(n794) );
  NAND2_X1 U3790 ( .A1(n13816), .A2(n14053), .ZN(n13647) );
  NAND2_X1 U3791 ( .A1(n17520), .A2(n795), .ZN(n16743) );
  NOR2_X1 U3792 ( .A1(n17106), .A2(n29406), .ZN(n795) );
  NAND2_X1 U3793 ( .A1(n17473), .A2(n796), .ZN(n3812) );
  OAI21_X1 U3794 ( .B1(n29364), .B2(n22286), .A(n21187), .ZN(n797) );
  NAND2_X1 U3795 ( .A1(n22023), .A2(n22290), .ZN(n21187) );
  NAND2_X1 U3797 ( .A1(n797), .A2(n22288), .ZN(n3857) );
  NAND2_X1 U3798 ( .A1(n800), .A2(n799), .ZN(n26809) );
  NAND2_X1 U3799 ( .A1(n27362), .A2(n27366), .ZN(n800) );
  AOI21_X1 U3800 ( .B1(n26809), .B2(n28562), .A(n801), .ZN(n26810) );
  NAND2_X1 U3801 ( .A1(n27362), .A2(n29538), .ZN(n802) );
  INV_X1 U3803 ( .A(n24804), .ZN(n803) );
  OAI21_X2 U3804 ( .B1(n23788), .B2(n807), .A(n804), .ZN(n24806) );
  NAND2_X1 U3805 ( .A1(n24027), .A2(n24263), .ZN(n2807) );
  NAND2_X1 U3806 ( .A1(n805), .A2(n23788), .ZN(n804) );
  OAI21_X1 U3807 ( .B1(n23785), .B2(n475), .A(n806), .ZN(n805) );
  NAND2_X1 U3808 ( .A1(n23785), .A2(n23786), .ZN(n806) );
  MUX2_X1 U3809 ( .A(n808), .B(n473), .S(n23036), .Z(n807) );
  INV_X1 U3810 ( .A(n23783), .ZN(n808) );
  OAI21_X2 U3811 ( .B1(n23757), .B2(n23034), .A(n3192), .ZN(n24804) );
  NAND2_X1 U3812 ( .A1(n20946), .A2(n28185), .ZN(n2724) );
  AND2_X1 U3813 ( .A1(n21501), .A2(n20944), .ZN(n20946) );
  INV_X1 U3814 ( .A(n24341), .ZN(n5571) );
  NAND2_X1 U3815 ( .A1(n24708), .A2(n24341), .ZN(n24125) );
  OR2_X1 U3818 ( .A1(n1908), .A2(n810), .ZN(n825) );
  NAND2_X1 U3819 ( .A1(n20456), .A2(n810), .ZN(n3953) );
  NAND2_X1 U3820 ( .A1(n20636), .A2(n20635), .ZN(n810) );
  NAND2_X1 U3821 ( .A1(n29470), .A2(n24386), .ZN(n813) );
  NAND3_X1 U3822 ( .A1(n24133), .A2(n24386), .A3(n29470), .ZN(n812) );
  NAND2_X1 U3823 ( .A1(n5307), .A2(n813), .ZN(n24134) );
  INV_X1 U3824 ( .A(n2874), .ZN(n814) );
  NAND2_X1 U3825 ( .A1(n18334), .A2(n817), .ZN(n18331) );
  NAND2_X1 U3827 ( .A1(n18370), .A2(n817), .ZN(n4213) );
  NAND2_X1 U3828 ( .A1(n17652), .A2(n816), .ZN(n18002) );
  NAND2_X1 U3829 ( .A1(n817), .A2(n18332), .ZN(n816) );
  OAI211_X1 U3831 ( .C1(n5728), .C2(n29470), .A(n24081), .B(n24135), .ZN(n818)
         );
  NAND3_X1 U3832 ( .A1(n616), .A2(n7017), .A3(n7692), .ZN(n3637) );
  XNOR2_X2 U3833 ( .A(Plaintext[83]), .B(Key[83]), .ZN(n7692) );
  XNOR2_X2 U3834 ( .A(n819), .B(Key[78]), .ZN(n7817) );
  INV_X1 U3835 ( .A(Plaintext[78]), .ZN(n819) );
  NAND2_X1 U3836 ( .A1(n4857), .A2(n23911), .ZN(n820) );
  NAND2_X1 U3837 ( .A1(n822), .A2(n382), .ZN(n821) );
  NAND2_X1 U3838 ( .A1(n383), .A2(n20476), .ZN(n822) );
  NAND3_X1 U3839 ( .A1(n5310), .A2(n28527), .A3(n823), .ZN(n23407) );
  NAND2_X1 U3840 ( .A1(n23405), .A2(n2239), .ZN(n823) );
  NAND3_X1 U3842 ( .A1(n2746), .A2(n20456), .A3(n825), .ZN(n21532) );
  OAI211_X1 U3843 ( .C1(n28102), .C2(n826), .A(n28101), .B(n28100), .ZN(n28104) );
  NAND2_X1 U3845 ( .A1(n14272), .A2(n14359), .ZN(n827) );
  NAND2_X1 U3846 ( .A1(n14271), .A2(n4166), .ZN(n14361) );
  NAND2_X1 U3849 ( .A1(n831), .A2(n24141), .ZN(n3541) );
  NAND2_X1 U3851 ( .A1(n24277), .A2(n831), .ZN(n5094) );
  NOR2_X1 U3852 ( .A1(n24590), .A2(n831), .ZN(n23855) );
  OAI21_X1 U3853 ( .B1(n24277), .B2(n831), .A(n24592), .ZN(n23856) );
  NAND2_X1 U3854 ( .A1(n24279), .A2(n831), .ZN(n5118) );
  OAI22_X1 U3855 ( .A1(n24593), .A2(n4692), .B1(n4966), .B2(n831), .ZN(n4152)
         );
  NAND2_X1 U3857 ( .A1(n23854), .A2(n831), .ZN(n840) );
  NAND2_X1 U3858 ( .A1(n3251), .A2(n831), .ZN(n5117) );
  NAND2_X1 U3859 ( .A1(n832), .A2(n20522), .ZN(n21334) );
  NAND2_X1 U3860 ( .A1(n1200), .A2(n1199), .ZN(n832) );
  OAI21_X1 U3861 ( .B1(n8786), .B2(n8717), .A(n8716), .ZN(n8791) );
  NAND2_X1 U3862 ( .A1(n834), .A2(n8788), .ZN(n8716) );
  INV_X1 U3863 ( .A(n8414), .ZN(n834) );
  INV_X1 U3864 ( .A(n8414), .ZN(n8720) );
  NAND2_X1 U3865 ( .A1(n8791), .A2(n8790), .ZN(n1294) );
  NAND3_X1 U3867 ( .A1(n15009), .A2(n15372), .A3(n14863), .ZN(n837) );
  OAI211_X2 U3868 ( .C1(n14374), .C2(n13594), .A(n4330), .B(n13727), .ZN(
        n14863) );
  NAND2_X1 U3869 ( .A1(n15370), .A2(n15371), .ZN(n14737) );
  OAI21_X1 U3870 ( .B1(n24474), .B2(n24471), .A(n53), .ZN(n6123) );
  MUX2_X1 U3872 ( .A(n23876), .B(n23875), .S(n6348), .Z(n23877) );
  NAND2_X1 U3873 ( .A1(n20483), .A2(n20485), .ZN(n20241) );
  XNOR2_X2 U3874 ( .A(n22708), .B(n22709), .ZN(n23442) );
  INV_X1 U3875 ( .A(n17565), .ZN(n1166) );
  OAI22_X1 U3876 ( .A1(n8343), .A2(n9133), .B1(n1670), .B2(n600), .ZN(n839) );
  INV_X1 U3877 ( .A(n20598), .ZN(n20273) );
  NAND2_X1 U3880 ( .A1(n23855), .A2(n24593), .ZN(n841) );
  NAND2_X1 U3881 ( .A1(n9136), .A2(n601), .ZN(n842) );
  NAND2_X1 U3882 ( .A1(n846), .A2(n28567), .ZN(n866) );
  NAND2_X1 U3884 ( .A1(n24019), .A2(n24541), .ZN(n846) );
  XNOR2_X1 U3885 ( .A(n847), .B(n26601), .ZN(Ciphertext[144]) );
  NAND4_X1 U3886 ( .A1(n26600), .A2(n26598), .A3(n26597), .A4(n26599), .ZN(
        n847) );
  NAND2_X1 U3887 ( .A1(n5514), .A2(n15419), .ZN(n3705) );
  AOI21_X2 U3889 ( .B1(n11418), .B2(n12146), .A(n848), .ZN(n12595) );
  AOI21_X1 U3890 ( .B1(n11416), .B2(n11417), .A(n11645), .ZN(n848) );
  INV_X1 U3891 ( .A(n1287), .ZN(n23060) );
  NAND2_X1 U3892 ( .A1(n23343), .A2(n23338), .ZN(n1287) );
  NAND3_X1 U3894 ( .A1(n14204), .A2(n2959), .A3(n14459), .ZN(n12704) );
  NAND3_X1 U3899 ( .A1(n4547), .A2(n4548), .A3(n14575), .ZN(n2731) );
  OAI21_X1 U3901 ( .B1(n16779), .B2(n17262), .A(n17258), .ZN(n16151) );
  OAI22_X1 U3902 ( .A1(n18430), .A2(n850), .B1(n17814), .B2(n18148), .ZN(
        n17817) );
  NAND2_X1 U3903 ( .A1(n18431), .A2(n18433), .ZN(n850) );
  NAND2_X1 U3904 ( .A1(n17517), .A2(n17518), .ZN(n17472) );
  NAND2_X1 U3905 ( .A1(n23336), .A2(n851), .ZN(n25761) );
  OAI21_X2 U3907 ( .B1(n24190), .B2(n24191), .A(n24189), .ZN(n25440) );
  OAI22_X1 U3908 ( .A1(n25669), .A2(n25670), .B1(n26474), .B2(n26181), .ZN(
        n852) );
  NAND2_X1 U3911 ( .A1(n3830), .A2(n13582), .ZN(n13645) );
  AND2_X1 U3914 ( .A1(n20351), .A2(n20783), .ZN(n20931) );
  NAND2_X1 U3915 ( .A1(n20847), .A2(n854), .ZN(n5942) );
  NAND2_X1 U3916 ( .A1(n21485), .A2(n20749), .ZN(n20847) );
  OAI21_X1 U3917 ( .B1(n28225), .B2(n406), .A(n855), .ZN(n23001) );
  NAND2_X1 U3918 ( .A1(n28225), .A2(n379), .ZN(n855) );
  NOR3_X1 U3919 ( .A1(n24617), .A2(n28550), .A3(n1631), .ZN(n24620) );
  XNOR2_X1 U3922 ( .A(n10029), .B(n9934), .ZN(n10287) );
  OR2_X1 U3923 ( .A1(n11594), .A2(n11932), .ZN(n11597) );
  AOI22_X1 U3924 ( .A1(n18508), .A2(n18271), .B1(n18273), .B2(n29057), .ZN(
        n856) );
  NAND2_X1 U3926 ( .A1(n8963), .A2(n605), .ZN(n2289) );
  XNOR2_X1 U3927 ( .A(n858), .B(n10391), .ZN(n9357) );
  INV_X1 U3928 ( .A(n9447), .ZN(n858) );
  NAND2_X1 U3929 ( .A1(n18297), .A2(n28745), .ZN(n2459) );
  AND2_X2 U3930 ( .A1(n7360), .A2(n7361), .ZN(n9148) );
  XNOR2_X1 U3931 ( .A(n859), .B(n8940), .ZN(n10472) );
  XNOR2_X1 U3932 ( .A(n8952), .B(n9523), .ZN(n859) );
  OR2_X1 U3934 ( .A1(n20972), .A2(n20966), .ZN(n21215) );
  NAND2_X1 U3935 ( .A1(n10853), .A2(n10851), .ZN(n11162) );
  NAND2_X1 U3936 ( .A1(n861), .A2(n18248), .ZN(n1784) );
  NAND2_X1 U3937 ( .A1(n863), .A2(n862), .ZN(n861) );
  NAND2_X1 U3938 ( .A1(n18707), .A2(n17353), .ZN(n862) );
  OR2_X1 U3940 ( .A1(n13888), .A2(n14317), .ZN(n12585) );
  INV_X1 U3941 ( .A(n15223), .ZN(n15227) );
  XNOR2_X1 U3942 ( .A(n16871), .B(n16870), .ZN(n20405) );
  OAI22_X1 U3944 ( .A1(n20548), .A2(n19857), .B1(n5982), .B2(n6315), .ZN(
        n21696) );
  XNOR2_X1 U3945 ( .A(n864), .B(n10285), .ZN(n5562) );
  XNOR2_X1 U3946 ( .A(n10284), .B(n10283), .ZN(n864) );
  OAI21_X1 U3947 ( .B1(n1736), .B2(n1735), .A(n11077), .ZN(n1734) );
  OR2_X1 U3949 ( .A1(n9140), .A2(n598), .ZN(n1127) );
  NAND2_X1 U3950 ( .A1(n27191), .A2(n27190), .ZN(n26290) );
  NOR2_X1 U3951 ( .A1(n23254), .A2(n867), .ZN(n23255) );
  NAND2_X1 U3952 ( .A1(n27645), .A2(n868), .ZN(n26672) );
  NAND2_X1 U3953 ( .A1(n27641), .A2(n27639), .ZN(n868) );
  NAND2_X1 U3954 ( .A1(n20001), .A2(n869), .ZN(n6137) );
  XNOR2_X1 U3955 ( .A(n16377), .B(n3856), .ZN(n16121) );
  OR2_X1 U3956 ( .A1(n29585), .A2(n27191), .ZN(n26138) );
  NAND2_X1 U3957 ( .A1(n18231), .A2(n18398), .ZN(n18397) );
  OAI21_X1 U3958 ( .B1(n12363), .B2(n12361), .A(n870), .ZN(n10899) );
  NOR2_X1 U3961 ( .A1(n15036), .A2(n15290), .ZN(n4955) );
  OAI211_X1 U3962 ( .C1(n21692), .C2(n21242), .A(n6311), .B(n21348), .ZN(n6312) );
  NAND2_X1 U3963 ( .A1(n1165), .A2(n1167), .ZN(n871) );
  INV_X1 U3964 ( .A(n21645), .ZN(n21042) );
  NAND2_X1 U3965 ( .A1(n10110), .A2(n10704), .ZN(n10708) );
  NAND2_X1 U3967 ( .A1(n1673), .A2(n1674), .ZN(n872) );
  NAND2_X2 U3969 ( .A1(n5970), .A2(n5969), .ZN(n15900) );
  XNOR2_X1 U3970 ( .A(n22357), .B(n22600), .ZN(n22361) );
  NAND2_X1 U3971 ( .A1(n5349), .A2(n24435), .ZN(n873) );
  NAND2_X1 U3972 ( .A1(n6293), .A2(n14605), .ZN(n874) );
  OAI21_X1 U3973 ( .B1(n18707), .B2(n876), .A(n875), .ZN(n18250) );
  NAND2_X1 U3974 ( .A1(n18707), .A2(n18404), .ZN(n875) );
  NAND2_X1 U3975 ( .A1(n2690), .A2(n11022), .ZN(n11316) );
  INV_X1 U3976 ( .A(n21511), .ZN(n20463) );
  NAND2_X1 U3977 ( .A1(n21532), .A2(n21534), .ZN(n21511) );
  XOR2_X1 U3978 ( .A(n16482), .B(n16478), .Z(n1094) );
  NAND3_X1 U3979 ( .A1(n877), .A2(n3342), .A3(n3343), .ZN(n18305) );
  NAND2_X1 U3980 ( .A1(n14694), .A2(n29600), .ZN(n877) );
  OAI21_X1 U3982 ( .B1(n23556), .B2(n23636), .A(n5143), .ZN(n878) );
  MUX2_X1 U3983 ( .A(n24068), .B(n24067), .S(n24677), .Z(n24069) );
  AOI22_X1 U3984 ( .A1(n26483), .A2(n1623), .B1(n29501), .B2(n26484), .ZN(
        n26487) );
  INV_X1 U3985 ( .A(n22514), .ZN(n21182) );
  INV_X1 U3986 ( .A(n21549), .ZN(n1621) );
  INV_X1 U3987 ( .A(n18333), .ZN(n1650) );
  NAND2_X1 U3988 ( .A1(n883), .A2(n8569), .ZN(n7387) );
  OAI21_X1 U3989 ( .B1(n9150), .B2(n8929), .A(n9374), .ZN(n883) );
  OAI211_X1 U3991 ( .C1(n28181), .C2(n23741), .A(n886), .B(n885), .ZN(n884) );
  NAND2_X1 U3992 ( .A1(n23741), .A2(n482), .ZN(n886) );
  NAND2_X1 U3995 ( .A1(n6832), .A2(n12513), .ZN(n3382) );
  NOR2_X2 U3996 ( .A1(n12715), .A2(n888), .ZN(n15420) );
  NAND2_X1 U3997 ( .A1(n25617), .A2(n27395), .ZN(n25621) );
  NAND2_X1 U3998 ( .A1(n17164), .A2(n28775), .ZN(n4293) );
  NAND2_X1 U3999 ( .A1(n890), .A2(n889), .ZN(n7724) );
  NAND2_X1 U4000 ( .A1(n7721), .A2(n7336), .ZN(n890) );
  NAND2_X1 U4003 ( .A1(n18382), .A2(n17881), .ZN(n18350) );
  NAND2_X1 U4004 ( .A1(n903), .A2(n905), .ZN(n23754) );
  NAND2_X1 U4005 ( .A1(n12510), .A2(n11990), .ZN(n6833) );
  NAND2_X1 U4006 ( .A1(n8740), .A2(n9073), .ZN(n9072) );
  AOI21_X1 U4008 ( .B1(n23796), .B2(n23321), .A(n23039), .ZN(n24336) );
  XNOR2_X1 U4009 ( .A(n892), .B(n19356), .ZN(n19358) );
  XNOR2_X1 U4010 ( .A(n19355), .B(n19354), .ZN(n892) );
  AND2_X1 U4011 ( .A1(n4478), .A2(n17361), .ZN(n17047) );
  NAND2_X1 U4012 ( .A1(n12206), .A2(n4037), .ZN(n4446) );
  AOI22_X1 U4013 ( .A1(n11851), .A2(n11853), .B1(n11852), .B2(n11921), .ZN(
        n11854) );
  OR2_X1 U4014 ( .A1(n14665), .A2(n14666), .ZN(n1053) );
  NAND3_X1 U4015 ( .A1(n5529), .A2(n20230), .A3(n4557), .ZN(n5528) );
  NAND2_X1 U4018 ( .A1(n1354), .A2(n29112), .ZN(n7088) );
  NAND3_X1 U4019 ( .A1(n24996), .A2(n24995), .A3(n894), .ZN(n24998) );
  NAND2_X1 U4021 ( .A1(n897), .A2(n895), .ZN(n10968) );
  NAND2_X1 U4022 ( .A1(n10687), .A2(n10961), .ZN(n895) );
  INV_X1 U4023 ( .A(n10959), .ZN(n896) );
  NOR2_X1 U4025 ( .A1(n11070), .A2(n262), .ZN(n898) );
  NAND2_X1 U4026 ( .A1(n20614), .A2(n899), .ZN(n1082) );
  AOI22_X1 U4027 ( .A1(n28036), .A2(n28037), .B1(n28034), .B2(n28035), .ZN(
        n28042) );
  NAND2_X1 U4028 ( .A1(n26661), .A2(n26662), .ZN(n28036) );
  AND3_X2 U4029 ( .A1(n23092), .A2(n23091), .A3(n3990), .ZN(n24380) );
  NAND3_X1 U4030 ( .A1(n9436), .A2(n9210), .A3(n8996), .ZN(n7680) );
  NAND2_X1 U4031 ( .A1(n7662), .A2(n8271), .ZN(n901) );
  NAND2_X1 U4034 ( .A1(n23744), .A2(n24514), .ZN(n905) );
  OR2_X1 U4035 ( .A1(n20479), .A2(n20480), .ZN(n4556) );
  NAND2_X1 U4036 ( .A1(n20298), .A2(n5933), .ZN(n20301) );
  NAND2_X1 U4038 ( .A1(n23848), .A2(n23845), .ZN(n908) );
  OAI21_X1 U4039 ( .B1(n909), .B2(n29227), .A(n21706), .ZN(n21711) );
  AOI21_X1 U4040 ( .B1(n21702), .B2(n21705), .A(n496), .ZN(n909) );
  NAND3_X1 U4041 ( .A1(n23911), .A2(n23389), .A3(n24077), .ZN(n23410) );
  OR2_X1 U4042 ( .A1(n21443), .A2(n21656), .ZN(n1109) );
  NAND2_X1 U4043 ( .A1(n14284), .A2(n14283), .ZN(n14290) );
  NAND2_X1 U4044 ( .A1(n7909), .A2(n8287), .ZN(n7474) );
  OAI211_X1 U4046 ( .C1(n23415), .C2(n23417), .A(n2435), .B(n23419), .ZN(n910)
         );
  OAI22_X1 U4048 ( .A1(n23807), .A2(n29102), .B1(n28594), .B2(n28653), .ZN(
        n22745) );
  NAND2_X1 U4050 ( .A1(n14079), .A2(n13744), .ZN(n912) );
  NAND2_X1 U4052 ( .A1(n914), .A2(n17846), .ZN(n913) );
  NAND2_X1 U4053 ( .A1(n917), .A2(n18144), .ZN(n916) );
  NAND2_X1 U4054 ( .A1(n918), .A2(n18143), .ZN(n917) );
  NAND2_X1 U4055 ( .A1(n2811), .A2(n18137), .ZN(n918) );
  OAI211_X1 U4057 ( .C1(n17526), .C2(n17157), .A(n920), .B(n17181), .ZN(n5919)
         );
  NAND2_X1 U4058 ( .A1(n17157), .A2(n17528), .ZN(n920) );
  NAND2_X1 U4059 ( .A1(n27865), .A2(n27877), .ZN(n27866) );
  NAND2_X1 U4060 ( .A1(n25720), .A2(n922), .ZN(n921) );
  NAND3_X1 U4061 ( .A1(n924), .A2(n3332), .A3(n27069), .ZN(n923) );
  NAND2_X1 U4062 ( .A1(n29076), .A2(n29520), .ZN(n924) );
  NAND2_X1 U4063 ( .A1(n28545), .A2(n29520), .ZN(n925) );
  INV_X1 U4064 ( .A(n14871), .ZN(n17400) );
  INV_X1 U4065 ( .A(n16825), .ZN(n926) );
  XNOR2_X1 U4066 ( .A(n928), .B(n927), .ZN(Ciphertext[87]) );
  NAND3_X1 U4067 ( .A1(n936), .A2(n932), .A3(n929), .ZN(n928) );
  NAND2_X1 U4068 ( .A1(n931), .A2(n930), .ZN(n929) );
  INV_X1 U4069 ( .A(n27591), .ZN(n27585) );
  NAND2_X1 U4070 ( .A1(n934), .A2(n933), .ZN(n932) );
  NOR2_X1 U4071 ( .A1(n27589), .A2(n935), .ZN(n934) );
  AND2_X1 U4072 ( .A1(n27591), .A2(n27590), .ZN(n935) );
  NAND2_X1 U4073 ( .A1(n27592), .A2(n1901), .ZN(n936) );
  AND2_X1 U4074 ( .A1(n2502), .A2(n937), .ZN(n938) );
  NAND2_X1 U4075 ( .A1(n8433), .A2(n9029), .ZN(n937) );
  INV_X1 U4076 ( .A(n17159), .ZN(n940) );
  NAND2_X1 U4077 ( .A1(n940), .A2(n424), .ZN(n939) );
  NAND2_X1 U4078 ( .A1(n17384), .A2(n18069), .ZN(n941) );
  XNOR2_X1 U4079 ( .A(n942), .B(n18145), .ZN(n18167) );
  XNOR2_X1 U4080 ( .A(n19469), .B(n942), .ZN(n19470) );
  XNOR2_X1 U4081 ( .A(n942), .B(n19017), .ZN(n19018) );
  XNOR2_X1 U4082 ( .A(n19370), .B(n18134), .ZN(n942) );
  NAND2_X1 U4083 ( .A1(n2141), .A2(n23258), .ZN(n943) );
  NAND4_X2 U4084 ( .A1(n8636), .A2(n8638), .A3(n8637), .A4(n944), .ZN(n10160)
         );
  NAND2_X1 U4085 ( .A1(n945), .A2(n2325), .ZN(n947) );
  NAND3_X1 U4087 ( .A1(n24587), .A2(n6055), .A3(n635), .ZN(n946) );
  XNOR2_X1 U4088 ( .A(n945), .B(n3232), .ZN(n24925) );
  XNOR2_X1 U4089 ( .A(n945), .B(n3516), .ZN(n25168) );
  XNOR2_X1 U4090 ( .A(n945), .B(n3114), .ZN(n25576) );
  XNOR2_X1 U4091 ( .A(n945), .B(n3635), .ZN(n25938) );
  XNOR2_X1 U4092 ( .A(n25785), .B(n945), .ZN(n25467) );
  NAND2_X1 U4093 ( .A1(n951), .A2(n949), .ZN(n25362) );
  XNOR2_X2 U4095 ( .A(n24574), .B(n24573), .ZN(n26560) );
  NAND2_X1 U4096 ( .A1(n954), .A2(n953), .ZN(n15301) );
  NAND2_X1 U4097 ( .A1(n14172), .A2(n957), .ZN(n953) );
  NAND3_X1 U4098 ( .A1(n14244), .A2(n957), .A3(n28172), .ZN(n954) );
  OAI21_X2 U4099 ( .B1(n956), .B2(n14172), .A(n957), .ZN(n15436) );
  NAND2_X1 U4100 ( .A1(n6573), .A2(n958), .ZN(n957) );
  OR2_X1 U4101 ( .A1(n13943), .A2(n15194), .ZN(n958) );
  AND2_X1 U4102 ( .A1(n14239), .A2(n14240), .ZN(n6573) );
  NAND2_X1 U4103 ( .A1(n23618), .A2(n960), .ZN(n23626) );
  NOR2_X1 U4104 ( .A1(n23566), .A2(n960), .ZN(n22986) );
  NAND3_X1 U4105 ( .A1(n23566), .A2(n23621), .A3(n960), .ZN(n23272) );
  OAI21_X1 U4106 ( .B1(n23570), .B2(n23571), .A(n960), .ZN(n23572) );
  OAI211_X1 U4107 ( .C1(n6646), .C2(n962), .A(n1947), .B(n961), .ZN(n13222) );
  NAND3_X1 U4108 ( .A1(n581), .A2(n3585), .A3(n10563), .ZN(n10511) );
  NAND2_X1 U4109 ( .A1(n20299), .A2(n20443), .ZN(n19924) );
  NAND2_X1 U4111 ( .A1(n10237), .A2(n3116), .ZN(n963) );
  XNOR2_X1 U4112 ( .A(n25933), .B(n26100), .ZN(n25112) );
  NAND3_X1 U4113 ( .A1(n965), .A2(n966), .A3(n24486), .ZN(n964) );
  OR2_X1 U4114 ( .A1(n24481), .A2(n24480), .ZN(n965) );
  NAND2_X1 U4115 ( .A1(n968), .A2(n6539), .ZN(n6538) );
  NOR2_X1 U4116 ( .A1(n17015), .A2(n968), .ZN(n17021) );
  NAND2_X1 U4117 ( .A1(n10808), .A2(n28627), .ZN(n969) );
  NAND2_X1 U4119 ( .A1(n261), .A2(n8427), .ZN(n8354) );
  INV_X1 U4120 ( .A(n8352), .ZN(n970) );
  NAND2_X1 U4122 ( .A1(n547), .A2(n15185), .ZN(n1570) );
  OAI21_X1 U4123 ( .B1(n14784), .B2(n972), .A(n15182), .ZN(n14532) );
  NAND2_X1 U4124 ( .A1(n15186), .A2(n972), .ZN(n1571) );
  OAI211_X1 U4125 ( .C1(n15190), .C2(n15183), .A(n15186), .B(n972), .ZN(n14800) );
  NAND2_X1 U4126 ( .A1(n13801), .A2(n13802), .ZN(n973) );
  NAND2_X1 U4127 ( .A1(n13800), .A2(n14312), .ZN(n974) );
  NAND2_X1 U4128 ( .A1(n18071), .A2(n18070), .ZN(n975) );
  NOR2_X1 U4129 ( .A1(n29496), .A2(n2032), .ZN(n18075) );
  NOR2_X2 U4130 ( .A1(n975), .A2(n5814), .ZN(n18510) );
  NAND2_X1 U4132 ( .A1(n626), .A2(n977), .ZN(n7436) );
  INV_X1 U4133 ( .A(n8217), .ZN(n977) );
  NAND2_X1 U4134 ( .A1(n14934), .A2(n14935), .ZN(n6286) );
  NAND2_X1 U4138 ( .A1(n24071), .A2(n24316), .ZN(n980) );
  MUX2_X1 U4141 ( .A(n11549), .B(n11922), .S(n11852), .Z(n10095) );
  AND2_X2 U4142 ( .A1(n6151), .A2(n10004), .ZN(n11852) );
  NAND2_X1 U4143 ( .A1(n3580), .A2(n427), .ZN(n981) );
  NAND2_X1 U4148 ( .A1(n23885), .A2(n24437), .ZN(n5349) );
  NAND2_X1 U4149 ( .A1(n24436), .A2(n24347), .ZN(n23885) );
  NOR2_X1 U4150 ( .A1(n23154), .A2(n23482), .ZN(n984) );
  NAND2_X1 U4153 ( .A1(n987), .A2(n15115), .ZN(n986) );
  NAND2_X1 U4154 ( .A1(n14740), .A2(n15117), .ZN(n987) );
  NAND2_X1 U4155 ( .A1(n1003), .A2(n544), .ZN(n988) );
  NAND2_X1 U4156 ( .A1(n990), .A2(n989), .ZN(n11536) );
  NAND2_X1 U4157 ( .A1(n10540), .A2(n10760), .ZN(n990) );
  NAND2_X1 U4158 ( .A1(n13586), .A2(n13602), .ZN(n13592) );
  NAND2_X1 U4159 ( .A1(n2248), .A2(n8350), .ZN(n2247) );
  AOI21_X1 U4161 ( .B1(n19880), .B2(n19881), .A(n20028), .ZN(n19885) );
  NAND3_X2 U4164 ( .A1(n3070), .A2(n3069), .A3(n3068), .ZN(n19440) );
  NAND2_X1 U4165 ( .A1(n14076), .A2(n14253), .ZN(n14096) );
  NAND2_X1 U4166 ( .A1(n991), .A2(n2824), .ZN(n2821) );
  NAND2_X1 U4167 ( .A1(n2822), .A2(n28567), .ZN(n991) );
  INV_X1 U4168 ( .A(n1650), .ZN(n1087) );
  OAI211_X2 U4169 ( .C1(n493), .C2(n21391), .A(n21390), .B(n992), .ZN(n22326)
         );
  NAND2_X1 U4170 ( .A1(n21388), .A2(n21387), .ZN(n992) );
  NOR2_X2 U4172 ( .A1(n994), .A2(n993), .ZN(n19123) );
  XNOR2_X1 U4175 ( .A(n22922), .B(n272), .ZN(n21996) );
  NAND2_X1 U4177 ( .A1(n997), .A2(n996), .ZN(n8058) );
  NAND2_X1 U4178 ( .A1(n7806), .A2(n7805), .ZN(n996) );
  INV_X1 U4179 ( .A(n20441), .ZN(n1081) );
  NAND2_X1 U4180 ( .A1(n11183), .A2(n11323), .ZN(n11186) );
  NAND2_X1 U4181 ( .A1(n8605), .A2(n9081), .ZN(n8850) );
  NAND2_X1 U4182 ( .A1(n4072), .A2(n998), .ZN(n15342) );
  INV_X1 U4184 ( .A(n24240), .ZN(n25794) );
  NAND2_X1 U4185 ( .A1(n999), .A2(n23186), .ZN(n24240) );
  NAND2_X1 U4186 ( .A1(n23184), .A2(n23566), .ZN(n999) );
  NAND2_X1 U4187 ( .A1(n17221), .A2(n29142), .ZN(n15847) );
  NAND2_X1 U4188 ( .A1(n5179), .A2(n5561), .ZN(n5178) );
  NOR2_X1 U4189 ( .A1(n12260), .A2(n11622), .ZN(n11581) );
  NAND2_X1 U4191 ( .A1(n1002), .A2(n1001), .ZN(n1000) );
  NAND2_X1 U4192 ( .A1(n15113), .A2(n15119), .ZN(n1003) );
  NAND2_X1 U4193 ( .A1(n15114), .A2(n1005), .ZN(n1004) );
  NAND2_X1 U4194 ( .A1(n15118), .A2(n15117), .ZN(n1006) );
  XNOR2_X1 U4195 ( .A(n9352), .B(n10335), .ZN(n9242) );
  NOR2_X1 U4196 ( .A1(n3155), .A2(n258), .ZN(n1007) );
  NAND3_X1 U4197 ( .A1(n17173), .A2(n29635), .A3(n16874), .ZN(n1799) );
  NAND2_X1 U4199 ( .A1(n1009), .A2(n17858), .ZN(n3540) );
  NAND3_X1 U4200 ( .A1(n17718), .A2(n5329), .A3(n17719), .ZN(n1009) );
  AOI22_X2 U4203 ( .A1(n7249), .A2(n8135), .B1(n1010), .B2(n615), .ZN(n8553)
         );
  OAI211_X1 U4205 ( .C1(n4998), .C2(n27926), .A(n27950), .B(n1011), .ZN(n4999)
         );
  INV_X1 U4206 ( .A(n29082), .ZN(n6615) );
  NAND2_X1 U4209 ( .A1(n3833), .A2(n3834), .ZN(n3832) );
  AND2_X1 U4210 ( .A1(n20483), .A2(n20484), .ZN(n19791) );
  NAND2_X1 U4211 ( .A1(n4058), .A2(n4059), .ZN(n18265) );
  INV_X1 U4212 ( .A(n18263), .ZN(n18262) );
  AND2_X1 U4215 ( .A1(n1166), .A2(n29098), .ZN(n1723) );
  INV_X1 U4216 ( .A(n17439), .ZN(n16962) );
  INV_X1 U4217 ( .A(n11780), .ZN(n11421) );
  INV_X1 U4218 ( .A(n18042), .ZN(n16862) );
  XNOR2_X1 U4219 ( .A(n10196), .B(n10197), .ZN(n11064) );
  INV_X1 U4220 ( .A(n21705), .ZN(n21373) );
  XNOR2_X1 U4222 ( .A(n15742), .B(n15743), .ZN(n16837) );
  AOI21_X1 U4224 ( .B1(n1013), .B2(n1012), .A(n24405), .ZN(n23910) );
  NAND2_X1 U4225 ( .A1(n3797), .A2(n24085), .ZN(n1012) );
  NAND2_X1 U4226 ( .A1(n6265), .A2(n24404), .ZN(n1013) );
  XNOR2_X2 U4227 ( .A(n1015), .B(n19281), .ZN(n19985) );
  XNOR2_X1 U4228 ( .A(n3659), .B(n18876), .ZN(n1015) );
  NAND2_X1 U4230 ( .A1(n20020), .A2(n19795), .ZN(n20518) );
  NAND2_X1 U4231 ( .A1(n6465), .A2(n17275), .ZN(n1017) );
  NAND2_X1 U4232 ( .A1(n16844), .A2(n539), .ZN(n1018) );
  OAI21_X1 U4234 ( .B1(n8579), .B2(n606), .A(n604), .ZN(n8771) );
  NAND3_X1 U4235 ( .A1(n7585), .A2(n7584), .A3(n7884), .ZN(n7304) );
  NAND2_X1 U4236 ( .A1(n1930), .A2(n21471), .ZN(n21475) );
  NAND2_X1 U4237 ( .A1(n1021), .A2(n5625), .ZN(n5624) );
  OR2_X1 U4239 ( .A1(n28478), .A2(n13646), .ZN(n5341) );
  OAI211_X1 U4240 ( .C1(n18153), .C2(n18154), .A(n18158), .B(n1022), .ZN(n1232) );
  NAND2_X1 U4241 ( .A1(n17825), .A2(n18154), .ZN(n1022) );
  NAND2_X1 U4242 ( .A1(n1309), .A2(n1023), .ZN(n15011) );
  INV_X1 U4243 ( .A(n1024), .ZN(n1023) );
  AOI21_X1 U4244 ( .B1(n14614), .B2(n14615), .A(n632), .ZN(n1024) );
  NAND2_X1 U4245 ( .A1(n15302), .A2(n15436), .ZN(n13944) );
  NAND2_X1 U4246 ( .A1(n1026), .A2(n1025), .ZN(n17810) );
  XNOR2_X2 U4248 ( .A(n7030), .B(Key[63]), .ZN(n7266) );
  NAND2_X1 U4249 ( .A1(n1028), .A2(n7915), .ZN(n1797) );
  OAI21_X1 U4250 ( .B1(n29568), .B2(n7909), .A(n7474), .ZN(n1028) );
  NAND3_X1 U4251 ( .A1(n15131), .A2(n14999), .A3(n15132), .ZN(n5866) );
  NAND2_X1 U4252 ( .A1(n14998), .A2(n15123), .ZN(n15131) );
  NAND2_X1 U4253 ( .A1(n26380), .A2(n1076), .ZN(n1029) );
  INV_X1 U4254 ( .A(n26425), .ZN(n1030) );
  NAND2_X1 U4256 ( .A1(n29321), .A2(n7846), .ZN(n6299) );
  NAND2_X1 U4258 ( .A1(n7522), .A2(n7268), .ZN(n1033) );
  OAI211_X1 U4261 ( .C1(n3440), .C2(n623), .A(n1730), .B(n1729), .ZN(n19433)
         );
  NAND3_X1 U4262 ( .A1(n2318), .A2(n2838), .A3(n2317), .ZN(n18867) );
  NAND2_X1 U4263 ( .A1(n1035), .A2(n20136), .ZN(n20138) );
  NAND2_X1 U4264 ( .A1(n19896), .A2(n2152), .ZN(n1035) );
  AND2_X2 U4267 ( .A1(n12624), .A2(n12625), .ZN(n3315) );
  NAND2_X1 U4269 ( .A1(n3737), .A2(n3739), .ZN(n18466) );
  OAI21_X1 U4270 ( .B1(n28015), .B2(n445), .A(n1037), .ZN(n28012) );
  NAND2_X1 U4271 ( .A1(n28015), .A2(n28017), .ZN(n1037) );
  NOR2_X1 U4273 ( .A1(n28104), .A2(n28103), .ZN(n1690) );
  INV_X1 U4275 ( .A(n4617), .ZN(n12037) );
  XNOR2_X1 U4276 ( .A(n10045), .B(n10411), .ZN(n1572) );
  AOI21_X2 U4277 ( .B1(n15354), .B2(n15353), .A(n15352), .ZN(n16279) );
  XNOR2_X1 U4278 ( .A(n9930), .B(n3073), .ZN(n9743) );
  NAND3_X1 U4280 ( .A1(n15434), .A2(n15431), .A3(n15432), .ZN(n14022) );
  NAND2_X1 U4284 ( .A1(n18136), .A2(n17846), .ZN(n17849) );
  OR2_X1 U4287 ( .A1(n18311), .A2(n17920), .ZN(n4629) );
  NAND3_X1 U4288 ( .A1(n24412), .A2(n24714), .A3(n28524), .ZN(n24411) );
  NOR2_X1 U4290 ( .A1(n21653), .A2(n6275), .ZN(n20244) );
  NAND2_X1 U4291 ( .A1(n17972), .A2(n17973), .ZN(n19409) );
  NAND3_X1 U4292 ( .A1(n20607), .A2(n1081), .A3(n20611), .ZN(n1040) );
  AOI21_X1 U4294 ( .B1(n5303), .B2(n20494), .A(n6834), .ZN(n1041) );
  NAND2_X1 U4295 ( .A1(n2514), .A2(n2516), .ZN(n1042) );
  INV_X1 U4296 ( .A(n20938), .ZN(n21309) );
  NAND2_X1 U4297 ( .A1(n1043), .A2(n20938), .ZN(n1315) );
  NAND3_X1 U4298 ( .A1(n20308), .A2(n20307), .A3(n20309), .ZN(n20938) );
  INV_X1 U4299 ( .A(n21306), .ZN(n1043) );
  OAI21_X1 U4301 ( .B1(n20055), .B2(n1044), .A(n2555), .ZN(n20058) );
  AOI21_X1 U4302 ( .B1(n20054), .B2(n20172), .A(n6114), .ZN(n1044) );
  NAND2_X1 U4303 ( .A1(n20917), .A2(n21287), .ZN(n20918) );
  NOR2_X1 U4304 ( .A1(n20986), .A2(n21288), .ZN(n20917) );
  AND2_X1 U4306 ( .A1(n1938), .A2(n7675), .ZN(n7678) );
  INV_X1 U4309 ( .A(n18421), .ZN(n4805) );
  OAI22_X1 U4310 ( .A1(n1456), .A2(n525), .B1(n17762), .B2(n17943), .ZN(n1455)
         );
  NAND2_X1 U4313 ( .A1(n13803), .A2(n14292), .ZN(n13804) );
  NAND3_X1 U4316 ( .A1(n5129), .A2(n5594), .A3(n8579), .ZN(n1045) );
  NAND2_X1 U4318 ( .A1(n11714), .A2(n11650), .ZN(n1048) );
  INV_X1 U4319 ( .A(n16815), .ZN(n1091) );
  OAI22_X1 U4320 ( .A1(n21893), .A2(n28444), .B1(n23689), .B2(n23537), .ZN(
        n23690) );
  NOR2_X2 U4321 ( .A1(n23528), .A2(n1049), .ZN(n24765) );
  NOR3_X1 U4322 ( .A1(n23527), .A2(n23662), .A3(n23526), .ZN(n1049) );
  NAND2_X1 U4324 ( .A1(n3936), .A2(n21562), .ZN(n1050) );
  NAND2_X1 U4325 ( .A1(n15434), .A2(n15030), .ZN(n5407) );
  NAND2_X1 U4326 ( .A1(n27340), .A2(n29052), .ZN(n27348) );
  NAND2_X1 U4327 ( .A1(n1052), .A2(n1051), .ZN(n1256) );
  NAND2_X1 U4328 ( .A1(n1622), .A2(n29579), .ZN(n1051) );
  NAND2_X1 U4329 ( .A1(n26726), .A2(n26727), .ZN(n1052) );
  NAND2_X1 U4331 ( .A1(n23600), .A2(n23467), .ZN(n23601) );
  NAND2_X1 U4332 ( .A1(n2656), .A2(n6526), .ZN(n17990) );
  NAND2_X1 U4333 ( .A1(n14664), .A2(n1053), .ZN(n15304) );
  XNOR2_X1 U4334 ( .A(n19271), .B(n1054), .ZN(n20272) );
  OR2_X1 U4336 ( .A1(n8265), .A2(n341), .ZN(n2472) );
  OAI21_X1 U4338 ( .B1(n22878), .B2(n4385), .A(n22743), .ZN(n22744) );
  AOI21_X1 U4339 ( .B1(n8459), .B2(n8524), .A(n8680), .ZN(n1056) );
  XNOR2_X1 U4340 ( .A(n19315), .B(n1057), .ZN(n18694) );
  XNOR2_X1 U4341 ( .A(n18689), .B(n18880), .ZN(n1057) );
  NAND2_X1 U4342 ( .A1(n1059), .A2(n1058), .ZN(n8577) );
  NAND2_X1 U4343 ( .A1(n8576), .A2(n29395), .ZN(n1058) );
  NAND2_X1 U4344 ( .A1(n1060), .A2(n8749), .ZN(n1059) );
  NAND2_X1 U4345 ( .A1(n9532), .A2(n9530), .ZN(n1060) );
  NAND2_X1 U4346 ( .A1(n1256), .A2(n1532), .ZN(n25629) );
  NAND2_X1 U4348 ( .A1(n2167), .A2(n12281), .ZN(n1061) );
  NAND2_X1 U4352 ( .A1(n1063), .A2(n12231), .ZN(n11987) );
  NAND2_X1 U4353 ( .A1(n9433), .A2(n11981), .ZN(n1063) );
  NAND2_X1 U4354 ( .A1(n13083), .A2(n303), .ZN(n9433) );
  XOR2_X1 U4356 ( .A(n13543), .B(n440), .Z(n6270) );
  OR2_X1 U4358 ( .A1(n2228), .A2(n10871), .ZN(n1163) );
  NAND2_X1 U4361 ( .A1(n18144), .A2(n526), .ZN(n17845) );
  OAI211_X1 U4362 ( .C1(n28206), .C2(n10742), .A(n28876), .B(n1064), .ZN(
        n10744) );
  NAND2_X1 U4364 ( .A1(n1066), .A2(n1065), .ZN(n14524) );
  NAND2_X1 U4365 ( .A1(n425), .A2(n15046), .ZN(n1065) );
  NAND2_X1 U4366 ( .A1(n15227), .A2(n15343), .ZN(n1066) );
  OAI21_X1 U4369 ( .B1(n27954), .B2(n27965), .A(n28636), .ZN(n1068) );
  NAND2_X1 U4370 ( .A1(n1069), .A2(n20322), .ZN(n3341) );
  OAI22_X1 U4371 ( .A1(n19956), .A2(n20319), .B1(n20324), .B2(n20323), .ZN(
        n1069) );
  NAND2_X1 U4372 ( .A1(n11782), .A2(n11502), .ZN(n11420) );
  OAI211_X1 U4373 ( .C1(n1292), .C2(n12343), .A(n1070), .B(n11474), .ZN(n11475) );
  NAND2_X1 U4374 ( .A1(n1290), .A2(n431), .ZN(n1070) );
  NAND2_X1 U4375 ( .A1(n1071), .A2(n11253), .ZN(n4649) );
  NAND2_X1 U4376 ( .A1(n11258), .A2(n11318), .ZN(n1071) );
  NAND3_X1 U4377 ( .A1(n15434), .A2(n15030), .A3(n14821), .ZN(n14023) );
  OR2_X1 U4379 ( .A1(n17277), .A2(n17276), .ZN(n17004) );
  INV_X1 U4380 ( .A(n1073), .ZN(n22875) );
  NAND2_X1 U4383 ( .A1(n26432), .A2(n26361), .ZN(n1075) );
  INV_X1 U4384 ( .A(n26425), .ZN(n1076) );
  XNOR2_X1 U4385 ( .A(n19267), .B(n6319), .ZN(n17974) );
  INV_X1 U4386 ( .A(n12677), .ZN(n1511) );
  NAND2_X1 U4388 ( .A1(n12239), .A2(n11514), .ZN(n4140) );
  NAND2_X1 U4389 ( .A1(n1450), .A2(n4141), .ZN(n1449) );
  AOI21_X1 U4392 ( .B1(n2246), .B2(n24461), .A(n24809), .ZN(n23951) );
  NAND3_X1 U4395 ( .A1(n1220), .A2(n1219), .A3(n10989), .ZN(n1080) );
  NAND2_X1 U4396 ( .A1(n11551), .A2(n11784), .ZN(n1140) );
  NAND2_X1 U4398 ( .A1(n1198), .A2(n7388), .ZN(n7392) );
  NAND2_X1 U4399 ( .A1(n21570), .A2(n21567), .ZN(n1084) );
  XNOR2_X2 U4400 ( .A(n1085), .B(n2293), .ZN(n14393) );
  OAI211_X1 U4401 ( .C1(n27326), .C2(n28641), .A(n27325), .B(n1086), .ZN(
        Ciphertext[148]) );
  NAND4_X1 U4402 ( .A1(n27323), .A2(n27320), .A3(n27322), .A4(n27321), .ZN(
        n1086) );
  XOR2_X1 U4407 ( .A(n22589), .B(n2522), .Z(n1773) );
  OAI21_X1 U4408 ( .B1(n18001), .B2(n18334), .A(n1087), .ZN(n1649) );
  NAND3_X1 U4409 ( .A1(n4586), .A2(n13724), .A3(n4331), .ZN(n4330) );
  OAI211_X1 U4410 ( .C1(n29086), .C2(n1091), .A(n1090), .B(n1089), .ZN(n1088)
         );
  NAND2_X1 U4411 ( .A1(n29086), .A2(n1466), .ZN(n1089) );
  NAND3_X1 U4412 ( .A1(n15434), .A2(n15432), .A3(n15030), .ZN(n15034) );
  NOR2_X2 U4413 ( .A1(n18030), .A2(n1092), .ZN(n18981) );
  OAI22_X1 U4414 ( .A1(n18027), .A2(n417), .B1(n29547), .B2(n18029), .ZN(n1092) );
  NAND2_X1 U4416 ( .A1(n7706), .A2(n7853), .ZN(n2590) );
  NAND2_X1 U4417 ( .A1(n7496), .A2(n7494), .ZN(n7706) );
  INV_X1 U4420 ( .A(n4270), .ZN(n17512) );
  XNOR2_X2 U4422 ( .A(n1094), .B(n5784), .ZN(n4270) );
  NAND2_X1 U4424 ( .A1(n15271), .A2(n1095), .ZN(n14615) );
  XOR2_X1 U4425 ( .A(n16246), .B(n15639), .Z(n1348) );
  NAND2_X1 U4430 ( .A1(n8874), .A2(n8699), .ZN(n8710) );
  OAI21_X1 U4431 ( .B1(n1334), .B2(n20517), .A(n20329), .ZN(n1099) );
  NAND3_X1 U4432 ( .A1(n14190), .A2(n14189), .A3(n14188), .ZN(n15223) );
  INV_X1 U4433 ( .A(n17954), .ZN(n20314) );
  OAI211_X1 U4434 ( .C1(n11280), .C2(n584), .A(n1100), .B(n585), .ZN(n3018) );
  NAND2_X1 U4435 ( .A1(n11280), .A2(n11281), .ZN(n1100) );
  NAND2_X1 U4437 ( .A1(n12079), .A2(n12296), .ZN(n1101) );
  NAND3_X1 U4438 ( .A1(n1104), .A2(n11482), .A3(n1103), .ZN(n1102) );
  INV_X1 U4439 ( .A(n11796), .ZN(n1104) );
  NAND2_X1 U4440 ( .A1(n618), .A2(n7266), .ZN(n8027) );
  XNOR2_X2 U4441 ( .A(n7027), .B(Key[65]), .ZN(n7268) );
  XNOR2_X1 U4442 ( .A(n28566), .B(n22641), .ZN(n22565) );
  NAND2_X1 U4443 ( .A1(n2619), .A2(n24437), .ZN(n24120) );
  INV_X1 U4444 ( .A(n19923), .ZN(n1105) );
  NAND2_X1 U4445 ( .A1(n1106), .A2(n13976), .ZN(n13977) );
  NAND2_X1 U4447 ( .A1(n1108), .A2(n2256), .ZN(n9292) );
  NAND2_X1 U4448 ( .A1(n2255), .A2(n10946), .ZN(n1108) );
  NAND2_X1 U4449 ( .A1(n18415), .A2(n18416), .ZN(n18417) );
  NAND2_X1 U4452 ( .A1(n21660), .A2(n21656), .ZN(n1110) );
  NAND2_X1 U4453 ( .A1(n8304), .A2(n7942), .ZN(n7659) );
  NAND3_X1 U4454 ( .A1(n13857), .A2(n13858), .A3(n29036), .ZN(n13860) );
  NAND2_X1 U4456 ( .A1(n15557), .A2(n542), .ZN(n1591) );
  NAND2_X1 U4458 ( .A1(n13585), .A2(n13645), .ZN(n1111) );
  NOR2_X2 U4459 ( .A1(n11667), .A2(n11668), .ZN(n13048) );
  MUX2_X1 U4460 ( .A(n1883), .B(n24372), .S(n24373), .Z(n24381) );
  NAND2_X1 U4462 ( .A1(n15395), .A2(n1112), .ZN(n1164) );
  NAND2_X1 U4463 ( .A1(n14723), .A2(n15144), .ZN(n1112) );
  NAND2_X1 U4465 ( .A1(n1594), .A2(n17348), .ZN(n1593) );
  NAND2_X1 U4468 ( .A1(n7920), .A2(n7619), .ZN(n7921) );
  OAI21_X1 U4469 ( .B1(n8228), .B2(n8227), .A(n8226), .ZN(n8230) );
  NAND2_X1 U4470 ( .A1(n18124), .A2(n18589), .ZN(n5475) );
  NAND2_X1 U4471 ( .A1(n1115), .A2(n2944), .ZN(n7537) );
  NAND2_X1 U4472 ( .A1(n8162), .A2(n7349), .ZN(n1115) );
  OAI21_X1 U4473 ( .B1(n11318), .B2(n594), .A(n1116), .ZN(n11259) );
  NAND2_X1 U4474 ( .A1(n11318), .A2(n2690), .ZN(n1116) );
  NAND2_X1 U4477 ( .A1(n9046), .A2(n5945), .ZN(n1118) );
  NAND4_X2 U4479 ( .A1(n2635), .A2(n18142), .A3(n2633), .A4(n18139), .ZN(
        n18852) );
  OR2_X1 U4480 ( .A1(n4188), .A2(n17259), .ZN(n1374) );
  INV_X1 U4482 ( .A(n17025), .ZN(n1121) );
  NAND2_X1 U4483 ( .A1(n17026), .A2(n17025), .ZN(n1122) );
  NAND3_X2 U4484 ( .A1(n5525), .A2(n5524), .A3(n11808), .ZN(n12776) );
  NAND2_X1 U4485 ( .A1(n4799), .A2(n14429), .ZN(n14199) );
  OAI21_X1 U4486 ( .B1(n1125), .B2(n18511), .A(n1124), .ZN(n18274) );
  NAND3_X1 U4487 ( .A1(n5931), .A2(n15284), .A3(n2893), .ZN(n5930) );
  NAND2_X1 U4489 ( .A1(n1127), .A2(n1126), .ZN(n9145) );
  NAND2_X1 U4490 ( .A1(n599), .A2(n9140), .ZN(n1126) );
  NAND2_X1 U4491 ( .A1(n13308), .A2(n263), .ZN(n15083) );
  OR2_X1 U4493 ( .A1(n24082), .A2(n24081), .ZN(n1128) );
  NAND2_X1 U4495 ( .A1(n1131), .A2(n1130), .ZN(n1129) );
  AOI21_X1 U4496 ( .B1(n17157), .B2(n16706), .A(n17181), .ZN(n1130) );
  NAND2_X1 U4497 ( .A1(n17526), .A2(n531), .ZN(n1131) );
  NAND2_X1 U4499 ( .A1(n1625), .A2(n6605), .ZN(n1132) );
  NAND2_X1 U4500 ( .A1(n24998), .A2(n24999), .ZN(n25052) );
  NAND2_X1 U4501 ( .A1(n1135), .A2(n1134), .ZN(n15332) );
  NAND2_X1 U4502 ( .A1(n16968), .A2(n17421), .ZN(n1134) );
  NAND2_X1 U4503 ( .A1(n17305), .A2(n17012), .ZN(n1135) );
  AND2_X1 U4506 ( .A1(n13803), .A2(n13699), .ZN(n12614) );
  NAND2_X1 U4507 ( .A1(n1561), .A2(n1137), .ZN(n6342) );
  XNOR2_X1 U4508 ( .A(n22710), .B(n22923), .ZN(n5841) );
  INV_X1 U4509 ( .A(n15184), .ZN(n15186) );
  INV_X1 U4510 ( .A(n10287), .ZN(n9311) );
  NOR2_X1 U4512 ( .A1(n11000), .A2(n10997), .ZN(n10683) );
  NAND2_X1 U4513 ( .A1(n11233), .A2(n11234), .ZN(n3442) );
  AOI21_X1 U4514 ( .B1(n23221), .B2(n23222), .A(n23220), .ZN(n23225) );
  NAND2_X1 U4515 ( .A1(n2708), .A2(n23700), .ZN(n23221) );
  NAND2_X1 U4516 ( .A1(n28810), .A2(n7935), .ZN(n7609) );
  NAND2_X1 U4519 ( .A1(n23740), .A2(n23741), .ZN(n23742) );
  NAND2_X1 U4520 ( .A1(n2911), .A2(n21624), .ZN(n3227) );
  NAND2_X1 U4521 ( .A1(n20381), .A2(n20567), .ZN(n18624) );
  XNOR2_X2 U4522 ( .A(n12397), .B(n12398), .ZN(n5584) );
  NAND2_X1 U4524 ( .A1(n1620), .A2(n7837), .ZN(n1139) );
  XNOR2_X1 U4526 ( .A(n9627), .B(n10079), .ZN(n1141) );
  OAI21_X1 U4527 ( .B1(n27603), .B2(n27604), .A(n1142), .ZN(n27606) );
  OAI21_X1 U4528 ( .B1(n27602), .B2(n27607), .A(n27617), .ZN(n1142) );
  XOR2_X1 U4529 ( .A(n16616), .B(n16141), .Z(n1575) );
  XOR2_X1 U4530 ( .A(n22000), .B(n22204), .Z(n1640) );
  NAND2_X1 U4531 ( .A1(n6663), .A2(n18197), .ZN(n1143) );
  OAI21_X1 U4532 ( .B1(n24243), .B2(n24242), .A(n1144), .ZN(n24244) );
  NAND2_X1 U4533 ( .A1(n1217), .A2(n1145), .ZN(n1144) );
  AND2_X1 U4534 ( .A1(n24240), .A2(n24241), .ZN(n1145) );
  INV_X1 U4535 ( .A(n4295), .ZN(n1801) );
  NAND2_X1 U4536 ( .A1(n9232), .A2(n9229), .ZN(n8544) );
  OAI21_X2 U4537 ( .B1(n6994), .B2(n6993), .A(n6992), .ZN(n9232) );
  NAND2_X1 U4539 ( .A1(n11065), .A2(n11242), .ZN(n1146) );
  NAND2_X1 U4541 ( .A1(n3924), .A2(n15343), .ZN(n1148) );
  NAND2_X1 U4542 ( .A1(n550), .A2(n425), .ZN(n1149) );
  NAND2_X1 U4544 ( .A1(n1808), .A2(n24341), .ZN(n5795) );
  NAND2_X1 U4547 ( .A1(n8663), .A2(n284), .ZN(n1789) );
  NAND2_X1 U4549 ( .A1(n24590), .A2(n24141), .ZN(n24144) );
  NAND2_X1 U4552 ( .A1(n23075), .A2(n23285), .ZN(n1150) );
  NAND2_X1 U4553 ( .A1(n23808), .A2(n23810), .ZN(n1151) );
  NAND2_X1 U4554 ( .A1(n2416), .A2(n15484), .ZN(n16921) );
  NAND2_X1 U4557 ( .A1(n17492), .A2(n536), .ZN(n1153) );
  NAND2_X1 U4558 ( .A1(n10778), .A2(n10958), .ZN(n10779) );
  NAND3_X1 U4559 ( .A1(n15733), .A2(n15732), .A3(n17236), .ZN(n18488) );
  NAND2_X1 U4560 ( .A1(n1154), .A2(n21547), .ZN(n20932) );
  NAND2_X1 U4561 ( .A1(n21553), .A2(n21519), .ZN(n1154) );
  OAI21_X1 U4562 ( .B1(n27715), .B2(n26126), .A(n1155), .ZN(n27696) );
  INV_X1 U4563 ( .A(n26889), .ZN(n1155) );
  NAND2_X1 U4564 ( .A1(n4980), .A2(n1156), .ZN(n21727) );
  NAND2_X1 U4565 ( .A1(n28223), .A2(n462), .ZN(n1156) );
  NAND2_X1 U4570 ( .A1(n1158), .A2(n442), .ZN(n2414) );
  NAND2_X1 U4571 ( .A1(n27627), .A2(n27632), .ZN(n1158) );
  NAND2_X1 U4573 ( .A1(n1159), .A2(n760), .ZN(n23218) );
  NAND2_X1 U4574 ( .A1(n23217), .A2(n476), .ZN(n1159) );
  NAND2_X2 U4575 ( .A1(n1160), .A2(n6146), .ZN(n13226) );
  NAND2_X1 U4576 ( .A1(n6145), .A2(n6658), .ZN(n1160) );
  NAND2_X1 U4577 ( .A1(n18034), .A2(n18033), .ZN(n17621) );
  OR2_X1 U4579 ( .A1(n8221), .A2(n7371), .ZN(n1358) );
  AOI22_X1 U4580 ( .A1(n26793), .A2(n28710), .B1(n26575), .B2(n26576), .ZN(
        n26925) );
  NAND2_X1 U4582 ( .A1(n1245), .A2(n5926), .ZN(n22298) );
  NOR3_X1 U4584 ( .A1(n25231), .A2(n25230), .A3(n26485), .ZN(n25238) );
  NAND2_X1 U4586 ( .A1(n19871), .A2(n3400), .ZN(n19879) );
  XOR2_X1 U4587 ( .A(n16495), .B(n15855), .Z(n1234) );
  OAI21_X1 U4588 ( .B1(n4557), .B2(n20474), .A(n5528), .ZN(n20739) );
  XNOR2_X1 U4589 ( .A(n22712), .B(n20923), .ZN(n1502) );
  AOI21_X1 U4590 ( .B1(n5761), .B2(n26748), .A(n5035), .ZN(n26634) );
  NAND2_X1 U4591 ( .A1(n27169), .A2(n28573), .ZN(n24990) );
  XNOR2_X1 U4592 ( .A(n25412), .B(n1302), .ZN(n24982) );
  NAND2_X1 U4594 ( .A1(n1166), .A2(n17227), .ZN(n1165) );
  NAND2_X1 U4595 ( .A1(n4717), .A2(n29138), .ZN(n1167) );
  XNOR2_X2 U4596 ( .A(n12591), .B(n12592), .ZN(n13803) );
  NAND2_X1 U4599 ( .A1(n17219), .A2(n17220), .ZN(n17223) );
  OR2_X1 U4600 ( .A1(n10517), .A2(n1854), .ZN(n10520) );
  OR2_X1 U4601 ( .A1(n7715), .A2(n6860), .ZN(n8793) );
  AND2_X1 U4602 ( .A1(n11113), .A2(n10461), .ZN(n1494) );
  NOR2_X1 U4604 ( .A1(n25650), .A2(n1169), .ZN(n25276) );
  NAND3_X1 U4605 ( .A1(n28494), .A2(n6621), .A3(n27372), .ZN(n6620) );
  NAND2_X1 U4606 ( .A1(n17205), .A2(n17818), .ZN(n1170) );
  NAND4_X2 U4607 ( .A1(n6192), .A2(n6189), .A3(n6190), .A4(n6191), .ZN(n10384)
         );
  NAND2_X1 U4608 ( .A1(n8362), .A2(n8361), .ZN(n1171) );
  NAND2_X1 U4609 ( .A1(n9012), .A2(n9016), .ZN(n5676) );
  NAND2_X1 U4611 ( .A1(n17232), .A2(n17361), .ZN(n17236) );
  INV_X1 U4612 ( .A(n17263), .ZN(n16991) );
  NAND2_X1 U4613 ( .A1(n18136), .A2(n526), .ZN(n2719) );
  NAND2_X1 U4614 ( .A1(n24303), .A2(n24369), .ZN(n1450) );
  NAND2_X1 U4615 ( .A1(n16725), .A2(n17481), .ZN(n4368) );
  NAND3_X1 U4617 ( .A1(n598), .A2(n9140), .A3(n8185), .ZN(n9141) );
  OAI21_X1 U4619 ( .B1(n4815), .B2(n11319), .A(n11318), .ZN(n1174) );
  NAND2_X1 U4620 ( .A1(n8147), .A2(n7792), .ZN(n7794) );
  NAND2_X1 U4622 ( .A1(n18174), .A2(n18171), .ZN(n1395) );
  AND3_X1 U4623 ( .A1(n23678), .A2(n23676), .A3(n23131), .ZN(n23365) );
  INV_X1 U4624 ( .A(n23469), .ZN(n23649) );
  NAND2_X1 U4625 ( .A1(n23469), .A2(n23647), .ZN(n22433) );
  NAND2_X1 U4626 ( .A1(n1441), .A2(n1443), .ZN(n17946) );
  NAND2_X1 U4627 ( .A1(n8360), .A2(n8433), .ZN(n8362) );
  NAND2_X1 U4629 ( .A1(n23684), .A2(n29544), .ZN(n1176) );
  NAND2_X1 U4630 ( .A1(n23685), .A2(n28457), .ZN(n1177) );
  NAND2_X1 U4631 ( .A1(n18087), .A2(n16985), .ZN(n16843) );
  NAND3_X1 U4632 ( .A1(n1546), .A2(n1547), .A3(n28004), .ZN(n1545) );
  NAND2_X1 U4633 ( .A1(n18332), .A2(n1180), .ZN(n1973) );
  INV_X1 U4634 ( .A(n7840), .ZN(n7420) );
  NAND2_X1 U4635 ( .A1(n7835), .A2(n7840), .ZN(n3112) );
  XNOR2_X2 U4636 ( .A(Key[87]), .B(Plaintext[87]), .ZN(n7840) );
  XOR2_X1 U4637 ( .A(n21855), .B(n6364), .Z(n1818) );
  AOI21_X1 U4638 ( .B1(n17710), .B2(n17572), .A(n423), .ZN(n1366) );
  XNOR2_X1 U4639 ( .A(n10252), .B(n1713), .ZN(n10254) );
  NOR2_X2 U4640 ( .A1(n21648), .A2(n1182), .ZN(n22067) );
  OAI21_X1 U4641 ( .B1(n21647), .B2(n21749), .A(n21646), .ZN(n1182) );
  XNOR2_X1 U4643 ( .A(n19650), .B(n1183), .ZN(n19282) );
  XNOR2_X1 U4644 ( .A(n19279), .B(n19280), .ZN(n1183) );
  NAND2_X1 U4645 ( .A1(n21458), .A2(n21457), .ZN(n20846) );
  XNOR2_X1 U4647 ( .A(n1185), .B(n26106), .ZN(n2902) );
  INV_X1 U4648 ( .A(n26107), .ZN(n1185) );
  NAND2_X1 U4649 ( .A1(n7912), .A2(n7628), .ZN(n8291) );
  AOI21_X1 U4650 ( .B1(n27630), .B2(n27616), .A(n1186), .ZN(n27622) );
  NAND3_X1 U4652 ( .A1(n29600), .A2(n29299), .A3(n17263), .ZN(n3878) );
  NAND2_X1 U4653 ( .A1(n14516), .A2(n1904), .ZN(n13668) );
  NAND2_X1 U4654 ( .A1(n13979), .A2(n14743), .ZN(n14516) );
  NAND3_X1 U4655 ( .A1(n1353), .A2(n1700), .A3(n7888), .ZN(n1352) );
  NAND2_X1 U4656 ( .A1(n1413), .A2(n20165), .ZN(n1188) );
  NAND2_X1 U4657 ( .A1(n1415), .A2(n19993), .ZN(n1189) );
  NAND2_X1 U4658 ( .A1(n8371), .A2(n8372), .ZN(n8373) );
  OR2_X1 U4659 ( .A1(n11168), .A2(n11166), .ZN(n10823) );
  OAI211_X1 U4660 ( .C1(n11336), .C2(n11338), .A(n1190), .B(n10558), .ZN(n2521) );
  NOR2_X1 U4662 ( .A1(n18468), .A2(n1191), .ZN(n6077) );
  NAND2_X1 U4663 ( .A1(n18472), .A2(n18469), .ZN(n1191) );
  NAND2_X1 U4665 ( .A1(n9231), .A2(n6590), .ZN(n5158) );
  NAND2_X1 U4666 ( .A1(n21213), .A2(n21211), .ZN(n21020) );
  NAND2_X1 U4667 ( .A1(n4217), .A2(n17421), .ZN(n16791) );
  NAND2_X1 U4668 ( .A1(n1737), .A2(n16789), .ZN(n4217) );
  NAND2_X1 U4671 ( .A1(n504), .A2(n29584), .ZN(n2555) );
  OAI21_X1 U4672 ( .B1(n24677), .B2(n24678), .A(n1194), .ZN(n24399) );
  NAND2_X1 U4673 ( .A1(n24677), .A2(n24395), .ZN(n1194) );
  INV_X1 U4674 ( .A(n5714), .ZN(n1738) );
  NAND2_X1 U4675 ( .A1(n5645), .A2(n5644), .ZN(n1244) );
  NOR2_X2 U4676 ( .A1(n1356), .A2(n14606), .ZN(n15309) );
  NAND2_X1 U4679 ( .A1(n21680), .A2(n21675), .ZN(n21672) );
  NAND2_X1 U4680 ( .A1(n10586), .A2(n11468), .ZN(n2589) );
  NAND2_X1 U4681 ( .A1(n3700), .A2(n3699), .ZN(n3698) );
  NAND3_X1 U4682 ( .A1(n21401), .A2(n21749), .A3(n20658), .ZN(n4647) );
  NAND2_X1 U4685 ( .A1(n20518), .A2(n501), .ZN(n1199) );
  NAND2_X1 U4686 ( .A1(n1201), .A2(n28126), .ZN(n1200) );
  NAND2_X1 U4687 ( .A1(n20520), .A2(n20517), .ZN(n1201) );
  NAND2_X1 U4689 ( .A1(n1204), .A2(n1203), .ZN(n1202) );
  NAND2_X1 U4692 ( .A1(n6451), .A2(n6452), .ZN(n21283) );
  OR2_X1 U4693 ( .A1(n14468), .A2(n4840), .ZN(n1628) );
  OR2_X1 U4694 ( .A1(n18068), .A2(n18067), .ZN(n1506) );
  NAND2_X1 U4695 ( .A1(n7802), .A2(n7803), .ZN(n7806) );
  NAND2_X1 U4696 ( .A1(n23805), .A2(n28594), .ZN(n1206) );
  INV_X1 U4697 ( .A(n15491), .ZN(n14703) );
  XNOR2_X1 U4698 ( .A(n1505), .B(n19243), .ZN(n19020) );
  XNOR2_X2 U4699 ( .A(Key[41]), .B(Plaintext[41]), .ZN(n7336) );
  AOI21_X1 U4702 ( .B1(n27097), .B2(n27531), .A(n1208), .ZN(n27098) );
  OAI22_X1 U4703 ( .A1(n27509), .A2(n27527), .B1(n27531), .B2(n27221), .ZN(
        n1208) );
  XNOR2_X1 U4704 ( .A(n1209), .B(n9917), .ZN(n9920) );
  XNOR2_X1 U4705 ( .A(n9918), .B(n1920), .ZN(n1209) );
  NAND3_X1 U4706 ( .A1(n8905), .A2(n6147), .A3(n9013), .ZN(n8907) );
  NAND2_X1 U4707 ( .A1(n1596), .A2(n29632), .ZN(n1592) );
  NAND2_X1 U4708 ( .A1(n1593), .A2(n1595), .ZN(n1596) );
  NAND2_X1 U4709 ( .A1(n16687), .A2(n6380), .ZN(n6379) );
  AOI21_X1 U4711 ( .B1(n6469), .B2(n28822), .A(n26949), .ZN(n1210) );
  NAND2_X1 U4712 ( .A1(n5903), .A2(n5904), .ZN(n3089) );
  NAND2_X1 U4713 ( .A1(n3147), .A2(n23771), .ZN(n6543) );
  NAND2_X1 U4714 ( .A1(n1211), .A2(n7835), .ZN(n7842) );
  NAND2_X1 U4715 ( .A1(n619), .A2(n7369), .ZN(n1211) );
  AND2_X2 U4716 ( .A1(n1213), .A2(n1212), .ZN(n16586) );
  NAND2_X1 U4717 ( .A1(n14809), .A2(n14810), .ZN(n1212) );
  NAND2_X1 U4718 ( .A1(n14811), .A2(n14812), .ZN(n1213) );
  NAND2_X1 U4719 ( .A1(n14715), .A2(n13922), .ZN(n14811) );
  MUX2_X1 U4721 ( .A(n11286), .B(n11285), .S(n11284), .Z(n1214) );
  OAI22_X1 U4722 ( .A1(n4423), .A2(n2974), .B1(n13903), .B2(n13902), .ZN(
        n14020) );
  NAND2_X1 U4724 ( .A1(n17481), .A2(n17476), .ZN(n3171) );
  INV_X1 U4726 ( .A(n24559), .ZN(n1217) );
  NAND3_X1 U4727 ( .A1(n17663), .A2(n18343), .A3(n17906), .ZN(n4075) );
  NAND2_X1 U4728 ( .A1(n2769), .A2(n17569), .ZN(n2768) );
  XNOR2_X1 U4729 ( .A(n1218), .B(n22413), .ZN(n22417) );
  XNOR2_X1 U4730 ( .A(n22412), .B(n22411), .ZN(n1218) );
  NAND2_X1 U4731 ( .A1(n6636), .A2(n21465), .ZN(n3936) );
  NAND2_X1 U4734 ( .A1(n10985), .A2(n589), .ZN(n1219) );
  NAND2_X1 U4735 ( .A1(n3804), .A2(n10984), .ZN(n1220) );
  OAI21_X1 U4736 ( .B1(n14045), .B2(n13906), .A(n14049), .ZN(n14052) );
  NAND2_X1 U4737 ( .A1(n12206), .A2(n12111), .ZN(n1221) );
  XNOR2_X2 U4738 ( .A(n3663), .B(n10300), .ZN(n10972) );
  OAI21_X1 U4739 ( .B1(n17815), .B2(n18045), .A(n1224), .ZN(n17816) );
  NAND3_X1 U4740 ( .A1(n1894), .A2(n18148), .A3(n18430), .ZN(n1224) );
  MUX2_X1 U4743 ( .A(n27551), .B(n27571), .S(n27573), .Z(n27219) );
  XNOR2_X1 U4746 ( .A(n1230), .B(n1229), .ZN(Ciphertext[64]) );
  NAND3_X1 U4747 ( .A1(n27284), .A2(n5331), .A3(n27283), .ZN(n1230) );
  OR2_X1 U4748 ( .A1(n1914), .A2(n28444), .ZN(n23024) );
  INV_X1 U4749 ( .A(n17827), .ZN(n1231) );
  NAND2_X1 U4750 ( .A1(n27088), .A2(n27084), .ZN(n27020) );
  XNOR2_X1 U4751 ( .A(n1234), .B(n16627), .ZN(n1233) );
  INV_X1 U4752 ( .A(n7967), .ZN(n1568) );
  NAND3_X1 U4755 ( .A1(n4348), .A2(n4347), .A3(n17673), .ZN(n18520) );
  XNOR2_X1 U4756 ( .A(n10251), .B(n1709), .ZN(n1713) );
  AOI21_X1 U4758 ( .B1(n7281), .B2(n7282), .A(n8150), .ZN(n1237) );
  NAND2_X1 U4760 ( .A1(n1238), .A2(n12300), .ZN(n2219) );
  NAND2_X1 U4762 ( .A1(n23813), .A2(n1239), .ZN(n24472) );
  NOR2_X1 U4763 ( .A1(n1240), .A2(n23814), .ZN(n1239) );
  OAI22_X1 U4765 ( .A1(n15847), .A2(n17553), .B1(n17224), .B2(n17556), .ZN(
        n1241) );
  OR2_X2 U4768 ( .A1(n1242), .A2(n7588), .ZN(n8718) );
  NAND2_X1 U4769 ( .A1(n2236), .A2(n2237), .ZN(n1242) );
  NAND2_X1 U4771 ( .A1(n1244), .A2(n15268), .ZN(n1243) );
  NAND2_X1 U4773 ( .A1(n24100), .A2(n29051), .ZN(n23875) );
  OAI211_X1 U4775 ( .C1(n24973), .C2(n24258), .A(n471), .B(n468), .ZN(n24259)
         );
  NAND2_X1 U4777 ( .A1(n468), .A2(n23467), .ZN(n1249) );
  MUX2_X1 U4780 ( .A(n468), .B(n23467), .S(n24976), .Z(n24014) );
  OAI21_X2 U4781 ( .B1(n17292), .B2(n28729), .A(n6524), .ZN(n6526) );
  NAND2_X1 U4782 ( .A1(n17400), .A2(n17397), .ZN(n1252) );
  XNOR2_X1 U4783 ( .A(n1254), .B(n25728), .ZN(n25733) );
  XNOR2_X1 U4784 ( .A(n1254), .B(n25015), .ZN(n24170) );
  XNOR2_X1 U4785 ( .A(n1254), .B(n25432), .ZN(n25433) );
  INV_X1 U4787 ( .A(n29037), .ZN(n1255) );
  XNOR2_X1 U4790 ( .A(n16093), .B(n16091), .ZN(n1257) );
  NAND2_X1 U4791 ( .A1(n1261), .A2(n1260), .ZN(n10654) );
  NAND2_X1 U4794 ( .A1(n1265), .A2(n1817), .ZN(n1264) );
  NAND2_X1 U4795 ( .A1(n1419), .A2(n16803), .ZN(n1265) );
  NAND2_X1 U4796 ( .A1(n17477), .A2(n3883), .ZN(n1419) );
  XNOR2_X1 U4797 ( .A(n1266), .B(n1271), .ZN(n1270) );
  OR2_X1 U4799 ( .A1(n3237), .A2(n628), .ZN(n1268) );
  NAND2_X1 U4800 ( .A1(n3237), .A2(n21088), .ZN(n22394) );
  OR2_X1 U4801 ( .A1(n21088), .A2(n628), .ZN(n1269) );
  INV_X1 U4802 ( .A(n1271), .ZN(n22773) );
  XNOR2_X1 U4803 ( .A(n1270), .B(n22395), .ZN(n3338) );
  NAND2_X1 U4804 ( .A1(n5505), .A2(n26489), .ZN(n1280) );
  NOR2_X1 U4805 ( .A1(n24678), .A2(n29555), .ZN(n24673) );
  NAND3_X1 U4806 ( .A1(n6406), .A2(n24674), .A3(n1272), .ZN(n24680) );
  NAND2_X1 U4807 ( .A1(n1274), .A2(n1273), .ZN(n1272) );
  NOR2_X1 U4808 ( .A1(n24678), .A2(n404), .ZN(n1273) );
  AOI21_X1 U4809 ( .B1(n29054), .B2(n26928), .A(n26927), .ZN(n1281) );
  NAND2_X1 U4810 ( .A1(n1276), .A2(n1275), .ZN(n26712) );
  NAND2_X1 U4811 ( .A1(n27433), .A2(n27439), .ZN(n1275) );
  NAND2_X1 U4812 ( .A1(n26829), .A2(n27434), .ZN(n1276) );
  OAI211_X2 U4813 ( .C1(n1279), .C2(n26166), .A(n1278), .B(n1277), .ZN(n27439)
         );
  NAND2_X1 U4814 ( .A1(n1280), .A2(n1281), .ZN(n1278) );
  NAND2_X1 U4817 ( .A1(n23074), .A2(n23285), .ZN(n22878) );
  NAND2_X1 U4818 ( .A1(n5265), .A2(n1285), .ZN(n4171) );
  NAND2_X1 U4819 ( .A1(n10723), .A2(n1285), .ZN(n10725) );
  NAND2_X1 U4820 ( .A1(n5743), .A2(n1286), .ZN(n5742) );
  NAND2_X1 U4821 ( .A1(n23474), .A2(n29620), .ZN(n1286) );
  NAND2_X1 U4822 ( .A1(n4546), .A2(n17977), .ZN(n17976) );
  NAND2_X1 U4823 ( .A1(n1287), .A2(n23428), .ZN(n23424) );
  NAND3_X1 U4824 ( .A1(n21591), .A2(n5983), .A3(n1921), .ZN(n4962) );
  NAND2_X1 U4825 ( .A1(n21588), .A2(n29569), .ZN(n1289) );
  AOI21_X1 U4826 ( .B1(n21323), .B2(n21588), .A(n1921), .ZN(n21324) );
  NOR2_X1 U4827 ( .A1(n1291), .A2(n12337), .ZN(n1290) );
  INV_X1 U4828 ( .A(n12026), .ZN(n1291) );
  INV_X1 U4829 ( .A(n20354), .ZN(n19032) );
  XNOR2_X1 U4831 ( .A(n1293), .B(n13556), .ZN(n13152) );
  XNOR2_X1 U4832 ( .A(n1293), .B(n12854), .ZN(n11939) );
  XNOR2_X1 U4833 ( .A(n13263), .B(n1293), .ZN(n12435) );
  XNOR2_X1 U4834 ( .A(n13244), .B(n1293), .ZN(n12538) );
  NAND2_X1 U4835 ( .A1(n1296), .A2(n1295), .ZN(n1297) );
  NAND2_X1 U4836 ( .A1(n7367), .A2(n7840), .ZN(n1296) );
  NAND2_X1 U4837 ( .A1(n7370), .A2(n370), .ZN(n1298) );
  NAND3_X1 U4838 ( .A1(n23075), .A2(n23074), .A3(n29102), .ZN(n22743) );
  OAI21_X1 U4839 ( .B1(n23074), .B2(n23806), .A(n23810), .ZN(n22638) );
  NAND2_X1 U4840 ( .A1(n24263), .A2(n28522), .ZN(n1299) );
  OAI21_X1 U4842 ( .B1(n24298), .B2(n1301), .A(n1300), .ZN(n1303) );
  OAI21_X1 U4843 ( .B1(n24298), .B2(n6198), .A(n630), .ZN(n1300) );
  NOR2_X2 U4844 ( .A1(n18096), .A2(n18091), .ZN(n17793) );
  NAND2_X1 U4845 ( .A1(n1308), .A2(n10937), .ZN(n9417) );
  AND2_X1 U4846 ( .A1(n1308), .A2(n10936), .ZN(n11005) );
  NAND2_X1 U4847 ( .A1(n11002), .A2(n28407), .ZN(n3640) );
  NOR2_X1 U4848 ( .A1(n11002), .A2(n28407), .ZN(n10684) );
  OAI21_X1 U4849 ( .B1(n10999), .B2(n10936), .A(n1308), .ZN(n9693) );
  NAND3_X1 U4850 ( .A1(n11002), .A2(n5573), .A3(n28407), .ZN(n11007) );
  NAND3_X1 U4851 ( .A1(n14614), .A2(n14615), .A3(n632), .ZN(n1309) );
  XNOR2_X1 U4852 ( .A(n1310), .B(n857), .ZN(n16046) );
  XNOR2_X1 U4853 ( .A(n15070), .B(n1310), .ZN(n15796) );
  XNOR2_X1 U4854 ( .A(n9645), .B(n9746), .ZN(n9687) );
  NAND3_X1 U4856 ( .A1(n8961), .A2(n8963), .A3(n9171), .ZN(n1311) );
  OAI21_X1 U4858 ( .B1(n21269), .B2(n20818), .A(n20711), .ZN(n1312) );
  NAND2_X1 U4859 ( .A1(n21266), .A2(n20816), .ZN(n20818) );
  NOR2_X2 U4860 ( .A1(n20876), .A2(n20877), .ZN(n21269) );
  NAND2_X1 U4862 ( .A1(n6362), .A2(n1314), .ZN(n6363) );
  NAND2_X1 U4863 ( .A1(n1314), .A2(n21150), .ZN(n21151) );
  NAND3_X1 U4864 ( .A1(n1318), .A2(n12181), .A3(n1319), .ZN(n1317) );
  NAND2_X1 U4866 ( .A1(n10441), .A2(n570), .ZN(n1316) );
  NAND2_X1 U4867 ( .A1(n1890), .A2(n12124), .ZN(n1319) );
  INV_X1 U4868 ( .A(n14177), .ZN(n1320) );
  NAND2_X1 U4870 ( .A1(n13850), .A2(n1322), .ZN(n1321) );
  NAND2_X1 U4871 ( .A1(n1324), .A2(n1323), .ZN(n4299) );
  NAND2_X1 U4872 ( .A1(n14991), .A2(n15389), .ZN(n1323) );
  NAND2_X1 U4873 ( .A1(n1326), .A2(n15145), .ZN(n1324) );
  AOI21_X1 U4875 ( .B1(n21644), .B2(n1327), .A(n21643), .ZN(n21648) );
  NAND2_X1 U4876 ( .A1(n15275), .A2(n15513), .ZN(n1328) );
  NAND3_X2 U4877 ( .A1(n1748), .A2(n1749), .A3(n6511), .ZN(n15274) );
  AOI21_X1 U4879 ( .B1(n2930), .B2(n2931), .A(n20567), .ZN(n1329) );
  OAI21_X1 U4880 ( .B1(n6237), .B2(n97), .A(n6236), .ZN(n1330) );
  NAND2_X1 U4883 ( .A1(n17458), .A2(n421), .ZN(n1332) );
  NAND3_X1 U4884 ( .A1(n17116), .A2(n16812), .A3(n17118), .ZN(n1333) );
  NAND2_X1 U4885 ( .A1(n29083), .A2(n29539), .ZN(n17458) );
  AND2_X1 U4887 ( .A1(n415), .A2(n6843), .ZN(n5934) );
  NAND2_X1 U4888 ( .A1(n6840), .A2(n507), .ZN(n6839) );
  NAND2_X1 U4889 ( .A1(n19505), .A2(n507), .ZN(n6838) );
  NAND2_X1 U4890 ( .A1(n19796), .A2(n28126), .ZN(n1334) );
  OAI211_X2 U4891 ( .C1(n2843), .C2(n1337), .A(n1521), .B(n1336), .ZN(n12132)
         );
  INV_X1 U4892 ( .A(n1704), .ZN(n1337) );
  NAND2_X1 U4893 ( .A1(n3820), .A2(n1338), .ZN(n10838) );
  NAND2_X1 U4894 ( .A1(n3817), .A2(n1338), .ZN(n1440) );
  OAI22_X1 U4897 ( .A1(n1340), .A2(n22011), .B1(n20762), .B2(n4828), .ZN(n1339) );
  NAND2_X1 U4899 ( .A1(n21823), .A2(n4828), .ZN(n1340) );
  AOI21_X1 U4900 ( .B1(n21077), .B2(n1342), .A(n21823), .ZN(n22014) );
  XNOR2_X2 U4901 ( .A(n13149), .B(n13148), .ZN(n14327) );
  OAI211_X1 U4903 ( .C1(n14324), .C2(n13653), .A(n14322), .B(n14323), .ZN(
        n1344) );
  NAND2_X1 U4904 ( .A1(n1346), .A2(n14328), .ZN(n1345) );
  NAND3_X1 U4906 ( .A1(n3731), .A2(n6506), .A3(n1808), .ZN(n2460) );
  NAND3_X1 U4907 ( .A1(n7774), .A2(n1350), .A3(n438), .ZN(n1349) );
  NAND2_X1 U4908 ( .A1(n3188), .A2(n438), .ZN(n1351) );
  NAND2_X1 U4909 ( .A1(n7774), .A2(n7777), .ZN(n1353) );
  XNOR2_X1 U4910 ( .A(n10019), .B(n1884), .ZN(n8883) );
  NAND2_X1 U4911 ( .A1(n8739), .A2(n8369), .ZN(n1417) );
  NAND3_X1 U4912 ( .A1(n11213), .A2(n11212), .A3(n1357), .ZN(n11214) );
  AOI21_X1 U4913 ( .B1(n1358), .B2(n7696), .A(n7695), .ZN(n7699) );
  OR2_X1 U4914 ( .A1(n10680), .A2(n29577), .ZN(n11983) );
  NAND2_X1 U4915 ( .A1(n11984), .A2(n11983), .ZN(n12231) );
  AND2_X1 U4916 ( .A1(n5265), .A2(n10970), .ZN(n1359) );
  OAI21_X1 U4919 ( .B1(n17562), .B2(n532), .A(n4220), .ZN(n1361) );
  NAND2_X1 U4920 ( .A1(n4873), .A2(n17561), .ZN(n1362) );
  NAND2_X1 U4921 ( .A1(n4220), .A2(n17315), .ZN(n17561) );
  OR2_X1 U4922 ( .A1(n17313), .A2(n17312), .ZN(n4873) );
  NAND2_X1 U4923 ( .A1(n423), .A2(n17570), .ZN(n2819) );
  NAND2_X1 U4924 ( .A1(n17320), .A2(n17707), .ZN(n1365) );
  NAND3_X1 U4926 ( .A1(n389), .A2(n1368), .A3(n4425), .ZN(n3741) );
  OR2_X1 U4927 ( .A1(n14144), .A2(n1368), .ZN(n6924) );
  NAND2_X1 U4928 ( .A1(n4423), .A2(n1368), .ZN(n14018) );
  NAND2_X1 U4929 ( .A1(n265), .A2(n13901), .ZN(n4421) );
  OAI21_X1 U4930 ( .B1(n389), .B2(n1368), .A(n14141), .ZN(n14145) );
  NAND2_X1 U4931 ( .A1(n1368), .A2(n2974), .ZN(n14141) );
  NAND3_X1 U4932 ( .A1(n12355), .A2(n1370), .A3(n1369), .ZN(n12461) );
  NAND2_X1 U4933 ( .A1(n10586), .A2(n1371), .ZN(n1370) );
  NAND3_X1 U4935 ( .A1(n4085), .A2(n1374), .A3(n17262), .ZN(n1373) );
  NOR2_X1 U4936 ( .A1(n12207), .A2(n12210), .ZN(n12209) );
  NAND2_X1 U4937 ( .A1(n9653), .A2(n11043), .ZN(n1375) );
  OAI21_X1 U4938 ( .B1(n28370), .B2(n17582), .A(n1377), .ZN(n1376) );
  NAND2_X1 U4939 ( .A1(n524), .A2(n17771), .ZN(n6912) );
  NAND2_X1 U4940 ( .A1(n524), .A2(n1378), .ZN(n1377) );
  NAND2_X1 U4941 ( .A1(n7373), .A2(n1379), .ZN(n7374) );
  NAND3_X1 U4942 ( .A1(n8227), .A2(n28721), .A3(n8221), .ZN(n1379) );
  INV_X1 U4943 ( .A(n6988), .ZN(n8227) );
  NAND2_X1 U4944 ( .A1(n592), .A2(n1380), .ZN(n2554) );
  XNOR2_X1 U4946 ( .A(n9745), .B(n9744), .ZN(n11010) );
  INV_X1 U4947 ( .A(n11010), .ZN(n1381) );
  OAI21_X1 U4948 ( .B1(n10628), .B2(n11235), .A(n11012), .ZN(n10579) );
  NAND2_X1 U4949 ( .A1(n1381), .A2(n11235), .ZN(n11012) );
  INV_X1 U4950 ( .A(n11010), .ZN(n6108) );
  NOR2_X1 U4951 ( .A1(n16338), .A2(n1382), .ZN(n16493) );
  AND2_X1 U4952 ( .A1(n6079), .A2(n1384), .ZN(n1382) );
  NAND2_X1 U4953 ( .A1(n1384), .A2(n18466), .ZN(n18472) );
  AND2_X1 U4954 ( .A1(n18467), .A2(n1384), .ZN(n18314) );
  AOI21_X1 U4955 ( .B1(n17915), .B2(n1384), .A(n18006), .ZN(n18010) );
  NAND2_X1 U4956 ( .A1(n16442), .A2(n1383), .ZN(n16492) );
  NAND2_X1 U4958 ( .A1(n603), .A2(n1386), .ZN(n9580) );
  NAND2_X1 U4959 ( .A1(n7912), .A2(n8290), .ZN(n7913) );
  NAND2_X1 U4960 ( .A1(n1388), .A2(n1961), .ZN(n14969) );
  NAND2_X1 U4961 ( .A1(n13470), .A2(n13469), .ZN(n1388) );
  OAI211_X1 U4962 ( .C1(n8914), .C2(n9107), .A(n8071), .B(n8669), .ZN(n8072)
         );
  NAND2_X1 U4963 ( .A1(n8071), .A2(n8669), .ZN(n8916) );
  NAND2_X1 U4965 ( .A1(n23155), .A2(n1641), .ZN(n1391) );
  MUX2_X1 U4966 ( .A(n17535), .B(n17536), .S(n18242), .Z(n17538) );
  NAND3_X1 U4967 ( .A1(n14696), .A2(n14845), .A3(n14695), .ZN(n1393) );
  NAND2_X1 U4968 ( .A1(n28198), .A2(n14842), .ZN(n1394) );
  NAND2_X1 U4969 ( .A1(n1395), .A2(n18170), .ZN(n2591) );
  NAND2_X1 U4970 ( .A1(n18169), .A2(n1395), .ZN(n18177) );
  NOR2_X1 U4971 ( .A1(n10622), .A2(n11227), .ZN(n10624) );
  XNOR2_X1 U4972 ( .A(n9956), .B(n260), .ZN(n1396) );
  XNOR2_X1 U4973 ( .A(n9722), .B(n9721), .ZN(n1397) );
  NAND2_X1 U4974 ( .A1(n436), .A2(n1398), .ZN(n8988) );
  NOR2_X1 U4975 ( .A1(n609), .A2(n8981), .ZN(n1398) );
  NAND3_X1 U4976 ( .A1(n10883), .A2(n11209), .A3(n11085), .ZN(n1400) );
  OAI21_X1 U4978 ( .B1(n12429), .B2(n12428), .A(n5134), .ZN(n1401) );
  OR2_X1 U4979 ( .A1(n12354), .A2(n580), .ZN(n5134) );
  OR2_X1 U4980 ( .A1(n7088), .A2(n438), .ZN(n1404) );
  NAND2_X1 U4981 ( .A1(n1403), .A2(n1402), .ZN(n4938) );
  NAND2_X1 U4982 ( .A1(n7088), .A2(n1700), .ZN(n1402) );
  NAND2_X1 U4983 ( .A1(n4939), .A2(n438), .ZN(n1403) );
  OAI21_X1 U4985 ( .B1(n17316), .B2(n790), .A(n1406), .ZN(n1405) );
  OR2_X1 U4986 ( .A1(n4220), .A2(n17315), .ZN(n1406) );
  NAND3_X1 U4988 ( .A1(n27301), .A2(n6150), .A3(n395), .ZN(n1407) );
  XNOR2_X1 U4989 ( .A(n1410), .B(n1412), .ZN(Ciphertext[70]) );
  NAND3_X1 U4990 ( .A1(n5425), .A2(n29493), .A3(n444), .ZN(n1411) );
  NAND2_X1 U4992 ( .A1(n20223), .A2(n297), .ZN(n1415) );
  NAND2_X1 U4993 ( .A1(n6578), .A2(n20219), .ZN(n20223) );
  NAND2_X1 U4994 ( .A1(n6901), .A2(n8734), .ZN(n1418) );
  NOR2_X1 U4995 ( .A1(n1419), .A2(n16723), .ZN(n17667) );
  INV_X1 U4997 ( .A(n29307), .ZN(n1420) );
  NAND2_X1 U5000 ( .A1(n1425), .A2(n1423), .ZN(n1422) );
  NAND2_X1 U5001 ( .A1(n29309), .A2(n23945), .ZN(n1423) );
  NAND3_X1 U5002 ( .A1(n470), .A2(n463), .A3(n29309), .ZN(n1424) );
  OR2_X1 U5003 ( .A1(n1427), .A2(n1470), .ZN(n1469) );
  NOR2_X1 U5004 ( .A1(n26484), .A2(n26731), .ZN(n1427) );
  NAND2_X1 U5005 ( .A1(n20197), .A2(n20589), .ZN(n1428) );
  INV_X1 U5007 ( .A(n13802), .ZN(n1430) );
  NAND2_X1 U5008 ( .A1(n14319), .A2(n14317), .ZN(n13802) );
  OR2_X1 U5009 ( .A1(n13802), .A2(n560), .ZN(n13712) );
  OAI21_X1 U5010 ( .B1(n13258), .B2(n1430), .A(n560), .ZN(n2331) );
  NAND2_X1 U5012 ( .A1(n28191), .A2(n17941), .ZN(n17763) );
  NAND2_X1 U5013 ( .A1(n28191), .A2(n1433), .ZN(n17944) );
  NOR2_X1 U5014 ( .A1(n1434), .A2(n17942), .ZN(n17602) );
  NAND2_X1 U5015 ( .A1(n525), .A2(n17762), .ZN(n1434) );
  NAND3_X1 U5016 ( .A1(n17937), .A2(n17939), .A3(n28191), .ZN(n16189) );
  INV_X1 U5017 ( .A(n1438), .ZN(n1574) );
  NAND2_X1 U5018 ( .A1(n1657), .A2(n1438), .ZN(n16852) );
  NAND3_X1 U5019 ( .A1(n1658), .A2(n1657), .A3(n1437), .ZN(n1656) );
  OAI21_X1 U5020 ( .B1(n16780), .B2(n16850), .A(n1438), .ZN(n16781) );
  NAND2_X1 U5021 ( .A1(n501), .A2(n20261), .ZN(n19794) );
  NAND3_X1 U5022 ( .A1(n501), .A2(n20261), .A3(n28133), .ZN(n21362) );
  NAND2_X1 U5023 ( .A1(n1439), .A2(n5716), .ZN(n12080) );
  OAI22_X1 U5024 ( .A1(n11251), .A2(n11250), .B1(n29149), .B2(n586), .ZN(n1439) );
  NAND2_X1 U5025 ( .A1(n1440), .A2(n3818), .ZN(n11251) );
  XNOR2_X2 U5026 ( .A(n9578), .B(n9933), .ZN(n11033) );
  NAND2_X1 U5027 ( .A1(n1442), .A2(n17941), .ZN(n1463) );
  NAND2_X1 U5028 ( .A1(n1442), .A2(n17939), .ZN(n1441) );
  NAND2_X1 U5029 ( .A1(n17940), .A2(n519), .ZN(n1443) );
  XNOR2_X1 U5030 ( .A(n22334), .B(n21955), .ZN(n22809) );
  NAND2_X1 U5032 ( .A1(n21450), .A2(n21675), .ZN(n1445) );
  INV_X1 U5033 ( .A(n1617), .ZN(n6111) );
  OAI211_X1 U5034 ( .C1(n28431), .C2(n22084), .A(n1635), .B(n6099), .ZN(n1446)
         );
  XNOR2_X1 U5035 ( .A(n25508), .B(n2602), .ZN(n24306) );
  NOR2_X2 U5036 ( .A1(n1449), .A2(n1447), .ZN(n25508) );
  AOI21_X1 U5037 ( .B1(n1448), .B2(n24305), .A(n23897), .ZN(n1447) );
  XNOR2_X1 U5038 ( .A(n2532), .B(n22389), .ZN(n1451) );
  NAND2_X1 U5039 ( .A1(n1453), .A2(n29137), .ZN(n1668) );
  NOR2_X1 U5041 ( .A1(n15132), .A2(n15127), .ZN(n1454) );
  NAND2_X1 U5043 ( .A1(n1454), .A2(n13632), .ZN(n13635) );
  NAND2_X1 U5044 ( .A1(n17943), .A2(n1457), .ZN(n1456) );
  NAND2_X1 U5045 ( .A1(n517), .A2(n28656), .ZN(n1457) );
  XNOR2_X1 U5046 ( .A(n1459), .B(n27894), .ZN(n25837) );
  XNOR2_X1 U5047 ( .A(n1459), .B(n25351), .ZN(n25082) );
  NAND2_X1 U5048 ( .A1(n21230), .A2(n21409), .ZN(n4632) );
  NAND2_X1 U5050 ( .A1(n1467), .A2(n1465), .ZN(n1464) );
  INV_X1 U5051 ( .A(n16679), .ZN(n1466) );
  NAND2_X1 U5052 ( .A1(n16814), .A2(n17282), .ZN(n1467) );
  AOI22_X1 U5053 ( .A1(n25641), .A2(n29579), .B1(n1473), .B2(n1472), .ZN(n1471) );
  NOR2_X1 U5054 ( .A1(n26480), .A2(n29579), .ZN(n1473) );
  XNOR2_X1 U5056 ( .A(n26029), .B(n4263), .ZN(n25507) );
  NAND2_X1 U5057 ( .A1(n23502), .A2(n23945), .ZN(n1476) );
  NAND2_X1 U5058 ( .A1(n1478), .A2(n458), .ZN(n1477) );
  AOI21_X1 U5059 ( .B1(n24780), .B2(n23946), .A(n23945), .ZN(n1478) );
  NAND2_X1 U5060 ( .A1(n24454), .A2(n24775), .ZN(n1479) );
  NAND2_X1 U5062 ( .A1(n17280), .A2(n4246), .ZN(n1481) );
  NAND2_X1 U5064 ( .A1(n1485), .A2(n11708), .ZN(n11709) );
  NAND2_X1 U5065 ( .A1(n11648), .A2(n12145), .ZN(n1484) );
  NAND2_X1 U5066 ( .A1(n15286), .A2(n14696), .ZN(n15287) );
  AND2_X1 U5068 ( .A1(n14842), .A2(n28996), .ZN(n15286) );
  NAND2_X1 U5071 ( .A1(n11645), .A2(n1487), .ZN(n3143) );
  NOR2_X1 U5072 ( .A1(n573), .A2(n11715), .ZN(n1487) );
  NAND2_X1 U5075 ( .A1(n11437), .A2(n12265), .ZN(n1490) );
  NAND2_X1 U5077 ( .A1(n1493), .A2(n11552), .ZN(n11554) );
  NAND2_X1 U5078 ( .A1(n1669), .A2(n1493), .ZN(n11504) );
  NAND2_X1 U5079 ( .A1(n11115), .A2(n11113), .ZN(n4128) );
  NAND2_X1 U5080 ( .A1(n11115), .A2(n1494), .ZN(n4630) );
  NAND3_X1 U5082 ( .A1(n24484), .A2(n1496), .A3(n1497), .ZN(n1495) );
  NAND2_X1 U5083 ( .A1(n29597), .A2(n24209), .ZN(n1496) );
  NAND2_X1 U5084 ( .A1(n24480), .A2(n24479), .ZN(n1497) );
  INV_X1 U5086 ( .A(n19229), .ZN(n1504) );
  XNOR2_X1 U5087 ( .A(n19349), .B(n1503), .ZN(n19518) );
  NOR2_X1 U5088 ( .A1(n4317), .A2(n1507), .ZN(n1509) );
  NAND2_X1 U5089 ( .A1(n15884), .A2(n17037), .ZN(n1508) );
  XNOR2_X1 U5090 ( .A(n12677), .B(n1510), .ZN(n13177) );
  INV_X1 U5091 ( .A(n13175), .ZN(n1510) );
  XNOR2_X1 U5092 ( .A(n1511), .B(n13380), .ZN(n13383) );
  XNOR2_X1 U5093 ( .A(n22459), .B(n633), .ZN(n21779) );
  NAND3_X1 U5094 ( .A1(n1513), .A2(n7796), .A3(n7794), .ZN(n1512) );
  NAND2_X1 U5095 ( .A1(n7541), .A2(n7793), .ZN(n1513) );
  XNOR2_X2 U5096 ( .A(n7149), .B(Key[24]), .ZN(n7793) );
  NAND2_X1 U5097 ( .A1(n1516), .A2(n28528), .ZN(n25007) );
  NAND2_X1 U5098 ( .A1(n25009), .A2(n28528), .ZN(n1517) );
  INV_X1 U5099 ( .A(n15514), .ZN(n15510) );
  AND2_X1 U5100 ( .A1(n1519), .A2(n14438), .ZN(n3851) );
  INV_X1 U5101 ( .A(n1876), .ZN(n1519) );
  OR2_X1 U5102 ( .A1(n14438), .A2(n1841), .ZN(n13959) );
  OAI21_X1 U5103 ( .B1(n13957), .B2(n13671), .A(n28200), .ZN(n4300) );
  OAI21_X2 U5104 ( .B1(n28200), .B2(n13849), .A(n13848), .ZN(n15168) );
  NAND3_X1 U5105 ( .A1(n586), .A2(n11248), .A3(n29148), .ZN(n1521) );
  INV_X1 U5107 ( .A(n18232), .ZN(n18401) );
  NAND2_X1 U5108 ( .A1(n18399), .A2(n18232), .ZN(n1523) );
  NAND2_X1 U5109 ( .A1(n390), .A2(n11867), .ZN(n6304) );
  NAND2_X1 U5110 ( .A1(n4126), .A2(n11116), .ZN(n1525) );
  XNOR2_X2 U5112 ( .A(n25266), .B(n25265), .ZN(n26753) );
  XNOR2_X1 U5115 ( .A(n22592), .B(n6938), .ZN(n23825) );
  OAI21_X2 U5116 ( .B1(n21297), .B2(n21296), .A(n21295), .ZN(n22644) );
  NAND2_X1 U5119 ( .A1(n9146), .A2(n8929), .ZN(n1529) );
  OR2_X2 U5120 ( .A1(n7374), .A2(n7375), .ZN(n9146) );
  AOI21_X1 U5121 ( .B1(n1530), .B2(n18042), .A(n29595), .ZN(n18044) );
  AND2_X2 U5122 ( .A1(n16855), .A2(n16854), .ZN(n18042) );
  INV_X1 U5123 ( .A(n22531), .ZN(n23833) );
  INV_X1 U5124 ( .A(n1534), .ZN(n27941) );
  OAI211_X1 U5125 ( .C1(n27016), .C2(n27017), .A(n1536), .B(n1535), .ZN(n1534)
         );
  NAND2_X1 U5126 ( .A1(n28441), .A2(n28451), .ZN(n1775) );
  NAND2_X1 U5127 ( .A1(n27011), .A2(n28446), .ZN(n1536) );
  INV_X1 U5128 ( .A(n11315), .ZN(n2689) );
  NAND2_X1 U5129 ( .A1(n4327), .A2(n1537), .ZN(n4329) );
  AOI21_X1 U5130 ( .B1(n2094), .B2(n29486), .A(n26735), .ZN(n28102) );
  NAND2_X1 U5132 ( .A1(n21533), .A2(n21534), .ZN(n1541) );
  NAND3_X1 U5133 ( .A1(n1544), .A2(n21536), .A3(n1543), .ZN(n1542) );
  INV_X1 U5134 ( .A(n21531), .ZN(n1544) );
  XNOR2_X1 U5135 ( .A(n1545), .B(n28007), .ZN(Ciphertext[171]) );
  NAND3_X1 U5136 ( .A1(n1548), .A2(n28002), .A3(n443), .ZN(n1547) );
  NAND3_X1 U5137 ( .A1(n23897), .A2(n25006), .A3(n28415), .ZN(n1549) );
  NAND2_X1 U5138 ( .A1(n1550), .A2(n1549), .ZN(n4558) );
  NAND2_X1 U5139 ( .A1(n4559), .A2(n1551), .ZN(n1550) );
  NAND2_X1 U5140 ( .A1(n12321), .A2(n12050), .ZN(n1552) );
  NAND3_X1 U5141 ( .A1(n12318), .A2(n12319), .A3(n1552), .ZN(n2979) );
  NAND2_X1 U5142 ( .A1(n428), .A2(n14295), .ZN(n13805) );
  NAND2_X1 U5143 ( .A1(n13806), .A2(n428), .ZN(n13702) );
  NAND2_X1 U5144 ( .A1(n17712), .A2(n18263), .ZN(n3834) );
  NAND2_X1 U5146 ( .A1(n16919), .A2(n790), .ZN(n1553) );
  NAND2_X1 U5147 ( .A1(n16920), .A2(n17317), .ZN(n1554) );
  NAND2_X1 U5150 ( .A1(n23555), .A2(n477), .ZN(n1555) );
  MUX2_X1 U5151 ( .A(n24635), .B(n24634), .S(n24633), .Z(n25793) );
  NAND2_X1 U5152 ( .A1(n23187), .A2(n23557), .ZN(n1558) );
  NAND2_X1 U5155 ( .A1(n1562), .A2(n1563), .ZN(n1561) );
  NAND2_X1 U5156 ( .A1(n18173), .A2(n18170), .ZN(n1562) );
  NAND2_X1 U5157 ( .A1(n20432), .A2(n1565), .ZN(n1564) );
  INV_X1 U5159 ( .A(n19920), .ZN(n20255) );
  OAI21_X1 U5164 ( .B1(n7678), .B2(n4697), .A(n1567), .ZN(n6540) );
  NAND2_X1 U5165 ( .A1(n7676), .A2(n4697), .ZN(n1567) );
  NAND3_X2 U5166 ( .A1(n1569), .A2(n4251), .A3(n4252), .ZN(n15190) );
  XNOR2_X1 U5167 ( .A(n1572), .B(n10188), .ZN(n1761) );
  XNOR2_X1 U5168 ( .A(n1572), .B(n9518), .ZN(n9522) );
  XNOR2_X1 U5169 ( .A(n9805), .B(n1572), .ZN(n9809) );
  AOI21_X1 U5170 ( .B1(n17262), .B2(n1574), .A(n17260), .ZN(n16782) );
  NAND2_X1 U5173 ( .A1(n16850), .A2(n1574), .ZN(n16150) );
  INV_X1 U5179 ( .A(n12938), .ZN(n1580) );
  MUX2_X1 U5181 ( .A(n16995), .B(n16992), .S(n17263), .Z(n1581) );
  NAND2_X1 U5182 ( .A1(n28176), .A2(n1865), .ZN(n6542) );
  NAND2_X1 U5186 ( .A1(n1584), .A2(n1585), .ZN(n8574) );
  NAND2_X1 U5187 ( .A1(n1586), .A2(n1587), .ZN(n1584) );
  OAI21_X1 U5188 ( .B1(n7777), .B2(n7890), .A(n1354), .ZN(n1588) );
  NAND2_X1 U5189 ( .A1(n7317), .A2(n1588), .ZN(n1587) );
  NAND2_X1 U5190 ( .A1(n1590), .A2(n14264), .ZN(n13615) );
  NAND2_X1 U5191 ( .A1(n14267), .A2(n1742), .ZN(n1590) );
  NAND2_X1 U5192 ( .A1(n1743), .A2(n14260), .ZN(n1742) );
  NAND2_X1 U5194 ( .A1(n14099), .A2(n14259), .ZN(n14267) );
  INV_X1 U5197 ( .A(n17025), .ZN(n1594) );
  NAND2_X1 U5198 ( .A1(n5420), .A2(n17025), .ZN(n1595) );
  NAND2_X1 U5200 ( .A1(n14659), .A2(n14658), .ZN(n15018) );
  NAND2_X1 U5201 ( .A1(n1598), .A2(n14467), .ZN(n14659) );
  NAND2_X1 U5202 ( .A1(n14185), .A2(n13933), .ZN(n1599) );
  NAND2_X1 U5203 ( .A1(n14466), .A2(n1600), .ZN(n14658) );
  NAND2_X1 U5204 ( .A1(n13933), .A2(n3843), .ZN(n1600) );
  OR2_X1 U5205 ( .A1(n14469), .A2(n14464), .ZN(n3843) );
  NAND3_X1 U5206 ( .A1(n527), .A2(n29044), .A3(n18087), .ZN(n1601) );
  NAND3_X1 U5207 ( .A1(n16843), .A2(n29125), .A3(n1603), .ZN(n1602) );
  OR2_X1 U5208 ( .A1(n18087), .A2(n18188), .ZN(n1603) );
  NOR2_X1 U5209 ( .A1(n19561), .A2(n18190), .ZN(n18088) );
  NAND3_X1 U5212 ( .A1(n7792), .A2(n1607), .A3(n7796), .ZN(n1606) );
  INV_X1 U5213 ( .A(n7542), .ZN(n1607) );
  OAI21_X1 U5214 ( .B1(n7792), .B2(n7541), .A(n8150), .ZN(n1608) );
  OAI211_X1 U5215 ( .C1(n12063), .C2(n12289), .A(n12062), .B(n1610), .ZN(
        n12697) );
  NAND3_X1 U5216 ( .A1(n12060), .A2(n29498), .A3(n1611), .ZN(n1610) );
  NAND3_X1 U5217 ( .A1(n12058), .A2(n12061), .A3(n12290), .ZN(n1611) );
  NAND3_X1 U5219 ( .A1(n7839), .A2(n370), .A3(n7840), .ZN(n1612) );
  NAND2_X1 U5220 ( .A1(n14604), .A2(n15515), .ZN(n1613) );
  AOI21_X1 U5221 ( .B1(n1616), .B2(n1615), .A(n608), .ZN(n1614) );
  NAND2_X1 U5222 ( .A1(n6147), .A2(n9014), .ZN(n1616) );
  NAND2_X1 U5223 ( .A1(n1617), .A2(n28401), .ZN(n4860) );
  NAND2_X1 U5225 ( .A1(n15731), .A2(n17232), .ZN(n17045) );
  INV_X1 U5226 ( .A(n17362), .ZN(n17232) );
  XNOR2_X1 U5228 ( .A(n19540), .B(n18639), .ZN(n1619) );
  NAND2_X1 U5229 ( .A1(n8210), .A2(n8211), .ZN(n1620) );
  OR2_X1 U5230 ( .A1(n7836), .A2(n7839), .ZN(n8211) );
  NAND3_X1 U5231 ( .A1(n21551), .A2(n1621), .A3(n21177), .ZN(n20930) );
  NAND2_X1 U5232 ( .A1(n21552), .A2(n1621), .ZN(n21522) );
  MUX2_X1 U5233 ( .A(n20351), .B(n21551), .S(n21549), .Z(n20784) );
  INV_X1 U5236 ( .A(n26480), .ZN(n1623) );
  NOR2_X1 U5237 ( .A1(n1624), .A2(n20504), .ZN(n1625) );
  INV_X1 U5238 ( .A(n20506), .ZN(n1624) );
  OAI21_X1 U5240 ( .B1(n6605), .B2(n29601), .A(n1626), .ZN(n19150) );
  NAND3_X1 U5241 ( .A1(n11963), .A2(n12219), .A3(n2846), .ZN(n11535) );
  NAND2_X1 U5242 ( .A1(n11963), .A2(n12219), .ZN(n11697) );
  NAND3_X1 U5243 ( .A1(n14466), .A2(n4840), .A3(n14467), .ZN(n1629) );
  NOR2_X1 U5245 ( .A1(n19791), .A2(n20486), .ZN(n1804) );
  NAND2_X1 U5248 ( .A1(n24746), .A2(n1632), .ZN(n24266) );
  NAND2_X1 U5249 ( .A1(n24617), .A2(n24747), .ZN(n1632) );
  MUX2_X2 U5250 ( .A(n21726), .B(n21727), .S(n24747), .Z(n25901) );
  NAND3_X1 U5251 ( .A1(n9034), .A2(n9035), .A3(n1634), .ZN(n2502) );
  NAND3_X1 U5253 ( .A1(n6472), .A2(n23739), .A3(n6474), .ZN(n1638) );
  XNOR2_X1 U5255 ( .A(n22777), .B(n1640), .ZN(n21742) );
  OR2_X1 U5256 ( .A1(n6081), .A2(n1642), .ZN(n24687) );
  NAND2_X1 U5257 ( .A1(n4118), .A2(n17569), .ZN(n1643) );
  XNOR2_X2 U5258 ( .A(n15868), .B(n16237), .ZN(n17569) );
  AND2_X2 U5259 ( .A1(n1646), .A2(n1645), .ZN(n1644) );
  INV_X2 U5260 ( .A(n1644), .ZN(n15434) );
  NAND2_X1 U5261 ( .A1(n15027), .A2(n1644), .ZN(n15028) );
  NAND2_X1 U5262 ( .A1(n1644), .A2(n14821), .ZN(n14683) );
  NAND3_X1 U5263 ( .A1(n15032), .A2(n1644), .A3(n15031), .ZN(n15033) );
  MUX2_X1 U5264 ( .A(n14823), .B(n14822), .S(n1644), .Z(n14829) );
  INV_X1 U5265 ( .A(n14014), .ZN(n1645) );
  NAND2_X1 U5266 ( .A1(n14015), .A2(n14351), .ZN(n1646) );
  NAND2_X1 U5267 ( .A1(n1648), .A2(n1647), .ZN(n18373) );
  NAND2_X1 U5268 ( .A1(n4412), .A2(n18333), .ZN(n1647) );
  NAND2_X1 U5269 ( .A1(n18371), .A2(n1650), .ZN(n1648) );
  MUX2_X1 U5270 ( .A(n1650), .B(n18370), .S(n18337), .Z(n18374) );
  NAND2_X1 U5271 ( .A1(n1649), .A2(n17061), .ZN(n19096) );
  MUX2_X1 U5272 ( .A(n1651), .B(n8485), .S(n81), .Z(n8489) );
  NAND3_X1 U5273 ( .A1(n24457), .A2(n24777), .A3(n24775), .ZN(n1654) );
  NAND2_X1 U5274 ( .A1(n24212), .A2(n29597), .ZN(n1652) );
  NAND2_X1 U5275 ( .A1(n1655), .A2(n24480), .ZN(n1653) );
  INV_X1 U5276 ( .A(n24211), .ZN(n24480) );
  NAND2_X1 U5277 ( .A1(n17258), .A2(n17259), .ZN(n1658) );
  NAND2_X1 U5278 ( .A1(n13717), .A2(n13900), .ZN(n1659) );
  XNOR2_X1 U5279 ( .A(n6647), .B(n1664), .ZN(n12707) );
  AND3_X1 U5281 ( .A1(n11971), .A2(n11972), .A3(n11973), .ZN(n1663) );
  XNOR2_X1 U5282 ( .A(n12644), .B(n1664), .ZN(n12588) );
  XNOR2_X1 U5283 ( .A(n11975), .B(n1664), .ZN(n11988) );
  NAND2_X1 U5284 ( .A1(n20368), .A2(n21581), .ZN(n6694) );
  AOI21_X1 U5285 ( .B1(n29737), .B2(n387), .A(n1666), .ZN(n1665) );
  INV_X1 U5286 ( .A(n17464), .ZN(n1666) );
  NAND2_X1 U5287 ( .A1(n528), .A2(n17280), .ZN(n1667) );
  NAND2_X1 U5288 ( .A1(n11420), .A2(n1668), .ZN(n1669) );
  NAND2_X1 U5289 ( .A1(n1669), .A2(n3900), .ZN(n11425) );
  NAND2_X1 U5290 ( .A1(n8342), .A2(n9132), .ZN(n8755) );
  INV_X1 U5291 ( .A(n1934), .ZN(n8342) );
  OAI22_X1 U5293 ( .A1(n14400), .A2(n28804), .B1(n13963), .B2(n29628), .ZN(
        n1671) );
  NAND2_X1 U5295 ( .A1(n21212), .A2(n28790), .ZN(n1673) );
  NAND2_X1 U5296 ( .A1(n5855), .A2(n22023), .ZN(n1674) );
  XNOR2_X1 U5297 ( .A(n22783), .B(n3317), .ZN(n22785) );
  NAND3_X1 U5298 ( .A1(n479), .A2(n28626), .A3(n483), .ZN(n1675) );
  AND2_X1 U5302 ( .A1(n24204), .A2(n1679), .ZN(n25321) );
  NAND2_X1 U5303 ( .A1(n28561), .A2(n28547), .ZN(n1679) );
  OAI21_X1 U5306 ( .B1(n1683), .B2(n26498), .A(n27372), .ZN(n1681) );
  NOR2_X1 U5308 ( .A1(n26497), .A2(n27364), .ZN(n1683) );
  INV_X1 U5309 ( .A(n25995), .ZN(n1684) );
  XNOR2_X1 U5310 ( .A(n16596), .B(n16393), .ZN(n16116) );
  OAI211_X2 U5311 ( .C1(n14739), .C2(n5198), .A(n5815), .B(n1685), .ZN(n16596)
         );
  NAND3_X1 U5312 ( .A1(n15379), .A2(n15384), .A3(n2203), .ZN(n1685) );
  INV_X1 U5313 ( .A(n12420), .ZN(n12980) );
  XNOR2_X1 U5314 ( .A(n11432), .B(n1686), .ZN(n11445) );
  XNOR2_X1 U5315 ( .A(n1687), .B(n12420), .ZN(n1686) );
  INV_X1 U5316 ( .A(n13179), .ZN(n1687) );
  XNOR2_X1 U5317 ( .A(n1688), .B(n28108), .ZN(Ciphertext[190]) );
  NAND2_X1 U5321 ( .A1(n1693), .A2(n489), .ZN(n1692) );
  NAND2_X1 U5322 ( .A1(n1695), .A2(n28790), .ZN(n1694) );
  MUX2_X1 U5323 ( .A(n22286), .B(n22290), .S(n21211), .Z(n1695) );
  NAND2_X1 U5325 ( .A1(n29294), .A2(n17179), .ZN(n1697) );
  AOI21_X1 U5328 ( .B1(n1698), .B2(n7628), .A(n7914), .ZN(n6999) );
  NAND2_X1 U5329 ( .A1(n7396), .A2(n1698), .ZN(n1796) );
  NAND2_X1 U5330 ( .A1(n7912), .A2(n7911), .ZN(n1698) );
  INV_X1 U5331 ( .A(n28692), .ZN(n1700) );
  OR2_X1 U5332 ( .A1(n28608), .A2(n591), .ZN(n10678) );
  NAND3_X1 U5333 ( .A1(n5267), .A2(n5265), .A3(n391), .ZN(n10950) );
  NAND3_X1 U5334 ( .A1(n6368), .A2(n6367), .A3(n391), .ZN(n6366) );
  NAND3_X1 U5336 ( .A1(n553), .A2(n15180), .A3(n15459), .ZN(n1702) );
  INV_X1 U5337 ( .A(n15180), .ZN(n15457) );
  NAND2_X1 U5338 ( .A1(n1934), .A2(n9134), .ZN(n8343) );
  NAND2_X1 U5339 ( .A1(n1934), .A2(n9133), .ZN(n9131) );
  NAND2_X1 U5340 ( .A1(n8753), .A2(n1934), .ZN(n7411) );
  NAND2_X1 U5341 ( .A1(n7397), .A2(n1934), .ZN(n7414) );
  NAND2_X1 U5342 ( .A1(n11248), .A2(n29666), .ZN(n1703) );
  NAND2_X1 U5343 ( .A1(n3819), .A2(n1704), .ZN(n3814) );
  NAND2_X1 U5344 ( .A1(n1706), .A2(n12145), .ZN(n11711) );
  AOI21_X1 U5345 ( .B1(n1706), .B2(n11645), .A(n11715), .ZN(n11647) );
  OAI21_X1 U5346 ( .B1(n12144), .B2(n1706), .A(n1705), .ZN(n5636) );
  NAND2_X1 U5347 ( .A1(n12147), .A2(n1706), .ZN(n1705) );
  NAND2_X1 U5348 ( .A1(n1707), .A2(n11322), .ZN(n6510) );
  NAND2_X1 U5349 ( .A1(n11184), .A2(n1707), .ZN(n8992) );
  NAND3_X1 U5350 ( .A1(n11181), .A2(n10473), .A3(n1707), .ZN(n3906) );
  INV_X1 U5351 ( .A(n10810), .ZN(n1707) );
  AND2_X1 U5352 ( .A1(n516), .A2(n18173), .ZN(n5223) );
  OAI21_X1 U5354 ( .B1(n17689), .B2(n4884), .A(n1708), .ZN(n16821) );
  OR2_X1 U5356 ( .A1(n8484), .A2(n440), .ZN(n1711) );
  NAND3_X1 U5357 ( .A1(n1710), .A2(n1711), .A3(n1712), .ZN(n1709) );
  NAND3_X1 U5358 ( .A1(n8483), .A2(n8484), .A3(n440), .ZN(n1712) );
  NAND2_X1 U5359 ( .A1(n4060), .A2(n610), .ZN(n1715) );
  XNOR2_X1 U5360 ( .A(n10328), .B(n625), .ZN(n8902) );
  NAND2_X1 U5361 ( .A1(n17896), .A2(n18322), .ZN(n1718) );
  NAND2_X2 U5362 ( .A1(n1721), .A2(n5999), .ZN(n18261) );
  NAND2_X1 U5364 ( .A1(n6417), .A2(n29138), .ZN(n16906) );
  OAI22_X1 U5366 ( .A1(n27758), .A2(n1724), .B1(n27740), .B2(n27741), .ZN(
        n27743) );
  INV_X1 U5367 ( .A(n27229), .ZN(n1724) );
  OR2_X1 U5368 ( .A1(n27732), .A2(n27759), .ZN(n27229) );
  NAND2_X1 U5370 ( .A1(n1725), .A2(n14667), .ZN(n14668) );
  INV_X1 U5371 ( .A(n15020), .ZN(n1725) );
  AND2_X1 U5372 ( .A1(n465), .A2(n24559), .ZN(n23989) );
  OAI21_X1 U5373 ( .B1(n24242), .B2(n1727), .A(n1726), .ZN(n24194) );
  INV_X1 U5374 ( .A(n24633), .ZN(n1727) );
  NAND2_X1 U5375 ( .A1(n402), .A2(n26837), .ZN(n1728) );
  OAI211_X1 U5377 ( .C1(n28631), .C2(n402), .A(n27120), .B(n1728), .ZN(n2270)
         );
  NAND2_X1 U5378 ( .A1(n3440), .A2(n3439), .ZN(n1733) );
  NAND2_X1 U5380 ( .A1(n1731), .A2(n3751), .ZN(n1730) );
  XNOR2_X1 U5381 ( .A(n1783), .B(n1732), .ZN(n19036) );
  INV_X1 U5382 ( .A(n19320), .ZN(n1732) );
  NAND2_X1 U5383 ( .A1(n5563), .A2(n1734), .ZN(n10533) );
  NOR2_X1 U5384 ( .A1(n11290), .A2(n29116), .ZN(n1735) );
  INV_X1 U5385 ( .A(n14240), .ZN(n2714) );
  NAND2_X1 U5386 ( .A1(n17615), .A2(n4217), .ZN(n3250) );
  NAND2_X1 U5387 ( .A1(n1738), .A2(n6002), .ZN(n1737) );
  NAND2_X1 U5389 ( .A1(n1739), .A2(n26228), .ZN(n26233) );
  NAND2_X1 U5390 ( .A1(n1740), .A2(n23648), .ZN(n5555) );
  XNOR2_X1 U5391 ( .A(n1741), .B(n3516), .ZN(n18666) );
  XNOR2_X1 U5392 ( .A(n18912), .B(n1741), .ZN(n16696) );
  XNOR2_X1 U5393 ( .A(n18913), .B(n1741), .ZN(n19133) );
  INV_X1 U5394 ( .A(n14260), .ZN(n13611) );
  INV_X1 U5395 ( .A(n14267), .ZN(n13613) );
  INV_X1 U5396 ( .A(n14268), .ZN(n1743) );
  NOR2_X1 U5397 ( .A1(n1744), .A2(n14998), .ZN(n15126) );
  NOR2_X1 U5398 ( .A1(n1745), .A2(n15127), .ZN(n13986) );
  NAND2_X1 U5399 ( .A1(n1745), .A2(n15004), .ZN(n14685) );
  NAND2_X1 U5400 ( .A1(n14686), .A2(n1745), .ZN(n14687) );
  NAND2_X1 U5401 ( .A1(n1746), .A2(n12507), .ZN(n10864) );
  NOR2_X1 U5402 ( .A1(n577), .A2(n12508), .ZN(n11989) );
  NAND3_X1 U5404 ( .A1(n12512), .A2(n577), .A3(n1746), .ZN(n11992) );
  NAND3_X1 U5405 ( .A1(n1747), .A2(n10165), .A3(n10166), .ZN(n10168) );
  NAND2_X1 U5406 ( .A1(n10572), .A2(n10883), .ZN(n1747) );
  NAND2_X1 U5407 ( .A1(n15511), .A2(n15274), .ZN(n15509) );
  MUX2_X1 U5408 ( .A(n14356), .B(n14357), .S(n4893), .Z(n1749) );
  MUX2_X1 U5410 ( .A(n9243), .B(n9041), .S(n9247), .Z(n1750) );
  XNOR2_X1 U5411 ( .A(n1751), .B(n21847), .ZN(n21852) );
  XNOR2_X1 U5412 ( .A(n21849), .B(n21848), .ZN(n1751) );
  NAND2_X1 U5414 ( .A1(n1753), .A2(n1752), .ZN(n5023) );
  NAND2_X1 U5416 ( .A1(n17360), .A2(n17359), .ZN(n1753) );
  XNOR2_X1 U5417 ( .A(n19231), .B(n19227), .ZN(n1756) );
  MUX2_X1 U5419 ( .A(n2853), .B(n18430), .S(n18431), .Z(n1759) );
  AND2_X1 U5420 ( .A1(n11068), .A2(n1760), .ZN(n5063) );
  INV_X1 U5421 ( .A(n11067), .ZN(n10880) );
  NAND2_X1 U5422 ( .A1(n3189), .A2(n1762), .ZN(n6049) );
  AOI21_X1 U5423 ( .B1(n23680), .B2(n474), .A(n28457), .ZN(n1762) );
  INV_X1 U5424 ( .A(n12166), .ZN(n12102) );
  NAND2_X1 U5426 ( .A1(n21033), .A2(n21473), .ZN(n1763) );
  NAND2_X1 U5427 ( .A1(n1765), .A2(n493), .ZN(n1764) );
  NAND2_X1 U5428 ( .A1(n1766), .A2(n21472), .ZN(n1765) );
  NAND2_X1 U5429 ( .A1(n29314), .A2(n21736), .ZN(n1766) );
  AND3_X2 U5430 ( .A1(n3341), .A2(n2956), .A3(n19957), .ZN(n21736) );
  NOR2_X1 U5431 ( .A1(n9247), .A2(n28211), .ZN(n6344) );
  NAND3_X1 U5432 ( .A1(n9248), .A2(n28211), .A3(n1768), .ZN(n9249) );
  INV_X1 U5433 ( .A(n9247), .ZN(n1768) );
  INV_X1 U5434 ( .A(n9014), .ZN(n1770) );
  NAND2_X1 U5435 ( .A1(n9015), .A2(n9014), .ZN(n1769) );
  OAI211_X2 U5436 ( .C1(n9019), .C2(n5674), .A(n9017), .B(n1771), .ZN(n10362)
         );
  XNOR2_X1 U5437 ( .A(n22651), .B(n1773), .ZN(n1772) );
  OAI21_X1 U5438 ( .B1(n1775), .B2(n27925), .A(n1774), .ZN(n27022) );
  NAND3_X1 U5439 ( .A1(n27925), .A2(n27944), .A3(n27938), .ZN(n1774) );
  AOI21_X2 U5440 ( .B1(n1776), .B2(n11371), .A(n1969), .ZN(n14893) );
  XNOR2_X1 U5442 ( .A(n15975), .B(n266), .ZN(n1778) );
  NAND2_X1 U5443 ( .A1(n17354), .A2(n17355), .ZN(n1779) );
  XNOR2_X1 U5444 ( .A(n12420), .B(n565), .ZN(n1780) );
  NOR2_X1 U5445 ( .A1(n505), .A2(n1781), .ZN(n19963) );
  XNOR2_X1 U5446 ( .A(n18959), .B(n1782), .ZN(n18577) );
  XNOR2_X1 U5447 ( .A(n18959), .B(n624), .ZN(n18977) );
  XNOR2_X1 U5448 ( .A(n1783), .B(n18959), .ZN(n17982) );
  OAI21_X1 U5449 ( .B1(n23604), .B2(n23606), .A(n1785), .ZN(n23249) );
  NAND2_X1 U5450 ( .A1(n23607), .A2(n23606), .ZN(n1785) );
  NAND2_X1 U5452 ( .A1(n3455), .A2(n3453), .ZN(n1787) );
  NAND2_X1 U5453 ( .A1(n12251), .A2(n12252), .ZN(n11934) );
  INV_X1 U5454 ( .A(n11934), .ZN(n11020) );
  INV_X1 U5455 ( .A(n8760), .ZN(n8569) );
  NAND3_X1 U5456 ( .A1(n6747), .A2(n9374), .A3(n6072), .ZN(n1791) );
  NAND2_X1 U5457 ( .A1(n9148), .A2(n9149), .ZN(n1788) );
  XNOR2_X2 U5459 ( .A(n13071), .B(n13072), .ZN(n4893) );
  AND2_X2 U5462 ( .A1(n1797), .A2(n1796), .ZN(n1934) );
  INV_X1 U5463 ( .A(n18101), .ZN(n16717) );
  NAND2_X1 U5464 ( .A1(n18193), .A2(n16718), .ZN(n18101) );
  NAND2_X1 U5466 ( .A1(n530), .A2(n29635), .ZN(n1800) );
  NAND2_X1 U5467 ( .A1(n16874), .A2(n17375), .ZN(n1802) );
  NAND2_X1 U5468 ( .A1(n8562), .A2(n9139), .ZN(n1803) );
  NAND2_X1 U5469 ( .A1(n29526), .A2(n21705), .ZN(n19187) );
  OAI22_X2 U5470 ( .A1(n1804), .A2(n20482), .B1(n20238), .B2(n19092), .ZN(
        n21705) );
  NAND2_X1 U5471 ( .A1(n5571), .A2(n1808), .ZN(n24415) );
  OAI21_X1 U5472 ( .B1(n24709), .B2(n1808), .A(n24417), .ZN(n1807) );
  NAND2_X1 U5473 ( .A1(n24710), .A2(n1808), .ZN(n5749) );
  AND2_X1 U5474 ( .A1(n1809), .A2(n15171), .ZN(n6925) );
  NAND2_X1 U5475 ( .A1(n1810), .A2(n20276), .ZN(n22657) );
  NAND2_X1 U5476 ( .A1(n2666), .A2(n1810), .ZN(n2665) );
  NAND2_X1 U5478 ( .A1(n8242), .A2(n616), .ZN(n3655) );
  OR2_X1 U5479 ( .A1(n11038), .A2(n28612), .ZN(n10671) );
  MUX2_X1 U5480 ( .A(n11273), .B(n28147), .S(n11038), .Z(n10673) );
  NOR2_X1 U5481 ( .A1(n11039), .A2(n1811), .ZN(n10846) );
  INV_X1 U5482 ( .A(n11038), .ZN(n1811) );
  NAND3_X1 U5484 ( .A1(n607), .A2(n602), .A3(n8594), .ZN(n1813) );
  INV_X1 U5485 ( .A(n21124), .ZN(n1814) );
  AND2_X1 U5486 ( .A1(n20842), .A2(n3838), .ZN(n20844) );
  NAND2_X1 U5487 ( .A1(n439), .A2(n7835), .ZN(n8210) );
  MUX2_X1 U5488 ( .A(n15896), .B(n15897), .S(n15434), .Z(n15898) );
  NAND2_X1 U5491 ( .A1(n16690), .A2(n534), .ZN(n1817) );
  INV_X1 U5492 ( .A(n11085), .ZN(n11212) );
  XNOR2_X1 U5493 ( .A(n1819), .B(n2476), .ZN(Ciphertext[28]) );
  NAND2_X1 U5494 ( .A1(n1622), .A2(n26485), .ZN(n26486) );
  XNOR2_X1 U5496 ( .A(n19308), .B(n4976), .ZN(n1823) );
  XNOR2_X1 U5497 ( .A(n7068), .B(Key[175]), .ZN(n7584) );
  XNOR2_X1 U5499 ( .A(n22647), .B(n22648), .ZN(n1829) );
  XNOR2_X1 U5500 ( .A(n22647), .B(n22648), .ZN(n23430) );
  INV_X1 U5501 ( .A(n14331), .ZN(n1830) );
  OR2_X1 U5502 ( .A1(n10546), .A2(n10545), .ZN(n1831) );
  XNOR2_X1 U5504 ( .A(n9982), .B(n9983), .ZN(n1834) );
  INV_X1 U5505 ( .A(n20109), .ZN(n1835) );
  INV_X1 U5506 ( .A(n578), .ZN(n1836) );
  XNOR2_X1 U5507 ( .A(n5862), .B(n22885), .ZN(n1837) );
  NAND2_X1 U5508 ( .A1(n19826), .A2(n19825), .ZN(n20865) );
  AOI21_X1 U5509 ( .B1(n10503), .B2(n10502), .A(n3458), .ZN(n11463) );
  XNOR2_X1 U5510 ( .A(n5862), .B(n22885), .ZN(n23145) );
  XNOR2_X1 U5512 ( .A(n22244), .B(n22243), .ZN(n1838) );
  XNOR2_X1 U5513 ( .A(n22244), .B(n22243), .ZN(n22992) );
  OAI211_X1 U5514 ( .C1(n8761), .C2(n8760), .A(n8759), .B(n8758), .ZN(n10151)
         );
  INV_X1 U5515 ( .A(n21016), .ZN(n1840) );
  INV_X1 U5516 ( .A(n14435), .ZN(n1841) );
  NAND2_X1 U5517 ( .A1(n7821), .A2(n7424), .ZN(n1842) );
  AND2_X1 U5518 ( .A1(n14834), .A2(n14833), .ZN(n2456) );
  NAND2_X1 U5519 ( .A1(n20016), .A2(n1844), .ZN(n1845) );
  NAND2_X1 U5520 ( .A1(n20015), .A2(n20014), .ZN(n1846) );
  NAND2_X1 U5521 ( .A1(n1845), .A2(n1846), .ZN(n20669) );
  INV_X1 U5522 ( .A(n20014), .ZN(n1844) );
  XNOR2_X1 U5525 ( .A(n2805), .B(n21825), .ZN(n22582) );
  INV_X1 U5527 ( .A(n15165), .ZN(n1848) );
  AND2_X1 U5528 ( .A1(n3844), .A2(n3846), .ZN(n1849) );
  OAI211_X1 U5531 ( .C1(n8882), .C2(n8881), .A(n8880), .B(n8879), .ZN(n1853)
         );
  XOR2_X1 U5533 ( .A(n10347), .B(n10348), .Z(n1855) );
  NAND2_X1 U5537 ( .A1(n11713), .A2(n3174), .ZN(n1857) );
  NAND2_X1 U5538 ( .A1(n3407), .A2(n20692), .ZN(n1858) );
  NAND2_X1 U5539 ( .A1(n3407), .A2(n20692), .ZN(n1859) );
  NAND2_X1 U5541 ( .A1(n11713), .A2(n3174), .ZN(n13269) );
  XOR2_X1 U5544 ( .A(n13005), .B(n13260), .Z(n12389) );
  OR2_X1 U5547 ( .A1(n18061), .A2(n17931), .ZN(n1863) );
  NAND4_X1 U5549 ( .A1(n15933), .A2(n15932), .A3(n15934), .A4(n17404), .ZN(
        n18057) );
  XNOR2_X1 U5550 ( .A(n4967), .B(n4968), .ZN(n23733) );
  OR2_X1 U5551 ( .A1(n26419), .A2(n26914), .ZN(n1864) );
  XNOR2_X1 U5552 ( .A(n3141), .B(n5195), .ZN(n1865) );
  OAI211_X1 U5553 ( .C1(n8939), .C2(n9144), .A(n8938), .B(n8937), .ZN(n1868)
         );
  AOI21_X1 U5556 ( .B1(n24004), .B2(n24547), .A(n24003), .ZN(n1871) );
  XNOR2_X1 U5557 ( .A(n6071), .B(n25390), .ZN(n1872) );
  XNOR2_X2 U5558 ( .A(n25400), .B(n25401), .ZN(n26914) );
  XNOR2_X1 U5559 ( .A(n3141), .B(n5195), .ZN(n10940) );
  OAI211_X1 U5560 ( .C1(n8939), .C2(n9144), .A(n8938), .B(n8937), .ZN(n9894)
         );
  XNOR2_X1 U5562 ( .A(n6071), .B(n25390), .ZN(n26565) );
  INV_X1 U5563 ( .A(n23138), .ZN(n1873) );
  AND2_X1 U5564 ( .A1(n25597), .A2(n25654), .ZN(n26742) );
  XNOR2_X1 U5565 ( .A(n25338), .B(n25339), .ZN(n1874) );
  OR2_X1 U5566 ( .A1(n20337), .A2(n3144), .ZN(n1875) );
  XNOR2_X1 U5567 ( .A(n12878), .B(n12877), .ZN(n1876) );
  AOI21_X1 U5568 ( .B1(n8582), .B2(n8583), .A(n8581), .ZN(n1877) );
  AOI21_X1 U5569 ( .B1(n8582), .B2(n8583), .A(n8581), .ZN(n1878) );
  XNOR2_X1 U5570 ( .A(n9445), .B(n9444), .ZN(n1879) );
  XNOR2_X1 U5571 ( .A(n12878), .B(n12877), .ZN(n14434) );
  AOI21_X1 U5572 ( .B1(n8582), .B2(n8583), .A(n8581), .ZN(n9517) );
  XNOR2_X1 U5573 ( .A(n19319), .B(n19318), .ZN(n20630) );
  NAND2_X1 U5575 ( .A1(n6579), .A2(n5940), .ZN(n1883) );
  OAI21_X1 U5576 ( .B1(n9868), .B2(n12186), .A(n9867), .ZN(n1885) );
  NAND2_X1 U5577 ( .A1(n6579), .A2(n5940), .ZN(n23995) );
  AND2_X1 U5578 ( .A1(n15691), .A2(n323), .ZN(n1886) );
  BUF_X1 U5579 ( .A(n11247), .Z(n12321) );
  XOR2_X1 U5581 ( .A(n18520), .B(n19427), .Z(n19234) );
  NAND3_X1 U5582 ( .A1(n4623), .A2(n17550), .A3(n17551), .ZN(n1888) );
  OAI211_X1 U5585 ( .C1(n9065), .C2(n9064), .A(n5537), .B(n5536), .ZN(n1891)
         );
  OAI211_X1 U5586 ( .C1(n9065), .C2(n9064), .A(n5537), .B(n5536), .ZN(n1892)
         );
  OAI211_X1 U5587 ( .C1(n9065), .C2(n9064), .A(n5537), .B(n5536), .ZN(n9661)
         );
  AOI22_X1 U5588 ( .A1(n6610), .A2(n23390), .B1(n6279), .B2(n23837), .ZN(n1893) );
  INV_X1 U5589 ( .A(n18433), .ZN(n1894) );
  XNOR2_X1 U5591 ( .A(n13253), .B(n13252), .ZN(n1896) );
  OR2_X1 U5592 ( .A1(n6635), .A2(n19801), .ZN(n1897) );
  XNOR2_X1 U5593 ( .A(n8706), .B(n8707), .ZN(n1898) );
  XNOR2_X1 U5594 ( .A(Key[21]), .B(Plaintext[21]), .ZN(n1899) );
  AOI22_X1 U5595 ( .A1(n6610), .A2(n23390), .B1(n6279), .B2(n23837), .ZN(
        n23393) );
  XNOR2_X1 U5596 ( .A(n8706), .B(n8707), .ZN(n10828) );
  XNOR2_X1 U5599 ( .A(n10175), .B(n10174), .ZN(n1900) );
  OR2_X1 U5600 ( .A1(n1968), .A2(n26262), .ZN(n1901) );
  NAND4_X1 U5601 ( .A1(n7187), .A2(n7186), .A3(n7185), .A4(n7184), .ZN(n1902)
         );
  NAND4_X1 U5603 ( .A1(n13658), .A2(n13659), .A3(n13702), .A4(n13657), .ZN(
        n1904) );
  NOR2_X1 U5604 ( .A1(n11110), .A2(n11109), .ZN(n1905) );
  NOR2_X1 U5605 ( .A1(n11110), .A2(n11109), .ZN(n1906) );
  INV_X1 U5607 ( .A(n498), .ZN(n1908) );
  NAND4_X1 U5608 ( .A1(n7187), .A2(n7186), .A3(n7185), .A4(n7184), .ZN(n9542)
         );
  NAND4_X1 U5609 ( .A1(n13658), .A2(n13659), .A3(n13702), .A4(n13657), .ZN(
        n15119) );
  XNOR2_X1 U5610 ( .A(n24971), .B(n24970), .ZN(n26386) );
  XNOR2_X1 U5611 ( .A(n19401), .B(n19400), .ZN(n20637) );
  INV_X1 U5613 ( .A(n1914), .ZN(n1913) );
  XNOR2_X1 U5615 ( .A(n19271), .B(n19270), .ZN(n1915) );
  XNOR2_X1 U5616 ( .A(n19271), .B(n19270), .ZN(n1916) );
  OAI21_X1 U5617 ( .B1(n9155), .B2(n9154), .A(n9153), .ZN(n1917) );
  OAI21_X1 U5618 ( .B1(n9155), .B2(n9154), .A(n9153), .ZN(n1918) );
  INV_X1 U5619 ( .A(n4861), .ZN(n1919) );
  NOR2_X1 U5620 ( .A1(n26355), .A2(n26354), .ZN(n27629) );
  XNOR2_X1 U5621 ( .A(n21874), .B(n21873), .ZN(n4726) );
  OAI21_X1 U5622 ( .B1(n9155), .B2(n9154), .A(n9153), .ZN(n10412) );
  INV_X1 U5624 ( .A(n20886), .ZN(n1921) );
  OAI21_X1 U5625 ( .B1(n23879), .B2(n23878), .A(n23877), .ZN(n1922) );
  OAI21_X1 U5627 ( .B1(n23879), .B2(n23878), .A(n23877), .ZN(n25107) );
  XNOR2_X1 U5629 ( .A(n6717), .B(n19018), .ZN(n20354) );
  XNOR2_X1 U5631 ( .A(n9982), .B(n9983), .ZN(n10498) );
  XNOR2_X1 U5635 ( .A(n9667), .B(n9666), .ZN(n10853) );
  XNOR2_X1 U5637 ( .A(n13253), .B(n13252), .ZN(n14047) );
  XNOR2_X1 U5638 ( .A(n24088), .B(n24089), .ZN(n26186) );
  OR2_X1 U5639 ( .A1(n8033), .A2(n8032), .ZN(n4061) );
  AOI21_X1 U5640 ( .B1(n7424), .B2(n7697), .A(n7824), .ZN(n7698) );
  OR2_X1 U5641 ( .A1(n4552), .A2(n7827), .ZN(n4550) );
  OR2_X1 U5642 ( .A1(n7856), .A2(n617), .ZN(n7857) );
  INV_X1 U5643 ( .A(n8910), .ZN(n5674) );
  XNOR2_X1 U5644 ( .A(n10137), .B(n10294), .ZN(n9736) );
  XNOR2_X1 U5646 ( .A(n10382), .B(n5896), .ZN(n5895) );
  AND2_X1 U5647 ( .A1(n10860), .A2(n10859), .ZN(n3570) );
  AOI22_X1 U5648 ( .A1(n5753), .A2(n2680), .B1(n4591), .B2(n11165), .ZN(n2678)
         );
  AND2_X1 U5649 ( .A1(n5526), .A2(n11806), .ZN(n5525) );
  XNOR2_X1 U5651 ( .A(n13291), .B(n12776), .ZN(n13513) );
  XNOR2_X1 U5652 ( .A(n13218), .B(n6821), .ZN(n6819) );
  XNOR2_X1 U5653 ( .A(n13219), .B(n1196), .ZN(n6821) );
  INV_X1 U5654 ( .A(n13674), .ZN(n14492) );
  INV_X1 U5655 ( .A(n14434), .ZN(n14437) );
  XNOR2_X1 U5656 ( .A(n13194), .B(n13193), .ZN(n13793) );
  INV_X1 U5657 ( .A(n13943), .ZN(n15199) );
  OR2_X1 U5658 ( .A1(n14070), .A2(n3798), .ZN(n3175) );
  INV_X1 U5659 ( .A(n14616), .ZN(n6797) );
  OR2_X1 U5660 ( .A1(n5678), .A2(n14916), .ZN(n14502) );
  NOR2_X1 U5661 ( .A1(n17259), .A2(n29574), .ZN(n16853) );
  INV_X1 U5662 ( .A(n17659), .ZN(n18317) );
  NOR2_X1 U5663 ( .A1(n18313), .A2(n18314), .ZN(n18318) );
  OR2_X1 U5664 ( .A1(n524), .A2(n2558), .ZN(n17777) );
  OAI211_X1 U5665 ( .C1(n18490), .C2(n18491), .A(n18487), .B(n3826), .ZN(n3825) );
  XNOR2_X1 U5666 ( .A(n3222), .B(n22697), .ZN(n21826) );
  OAI211_X1 U5667 ( .C1(n7165), .C2(n7279), .A(n5282), .B(n2692), .ZN(n7175)
         );
  OR2_X1 U5669 ( .A1(n7533), .A2(n8014), .ZN(n8018) );
  XNOR2_X1 U5670 ( .A(n6977), .B(Key[101]), .ZN(n7830) );
  NOR2_X1 U5671 ( .A1(n7657), .A2(n8304), .ZN(n7207) );
  INV_X1 U5672 ( .A(n29317), .ZN(n8297) );
  INV_X1 U5673 ( .A(n7692), .ZN(n8243) );
  OR2_X1 U5674 ( .A1(n7690), .A2(n7376), .ZN(n3511) );
  OR2_X1 U5676 ( .A1(n8927), .A2(n9132), .ZN(n3101) );
  XNOR2_X1 U5678 ( .A(n4508), .B(n4507), .ZN(n4505) );
  XNOR2_X1 U5679 ( .A(n9714), .B(n6916), .ZN(n10620) );
  OR2_X1 U5680 ( .A1(n6272), .A2(n11198), .ZN(n4710) );
  AND3_X1 U5682 ( .A1(n3046), .A2(n3047), .A3(n11282), .ZN(n10653) );
  OR2_X1 U5683 ( .A1(n11583), .A2(n10869), .ZN(n6328) );
  NAND2_X1 U5684 ( .A1(n11813), .A2(n11814), .ZN(n12985) );
  NOR2_X1 U5685 ( .A1(n11809), .A2(n11982), .ZN(n4021) );
  OR2_X1 U5686 ( .A1(n14426), .A2(n12534), .ZN(n13871) );
  NOR2_X1 U5687 ( .A1(n4046), .A2(n6482), .ZN(n6481) );
  OR2_X1 U5688 ( .A1(n11714), .A2(n11715), .ZN(n3174) );
  XNOR2_X1 U5689 ( .A(n5122), .B(n4041), .ZN(n14440) );
  XNOR2_X1 U5690 ( .A(n12778), .B(n12779), .ZN(n14494) );
  XNOR2_X1 U5691 ( .A(n6895), .B(n12584), .ZN(n14309) );
  INV_X1 U5692 ( .A(n13257), .ZN(n14312) );
  INV_X1 U5693 ( .A(n14106), .ZN(n14231) );
  INV_X1 U5694 ( .A(n14440), .ZN(n14432) );
  OR2_X1 U5695 ( .A1(n14379), .A2(n4258), .ZN(n14384) );
  INV_X1 U5696 ( .A(n15402), .ZN(n14943) );
  OR2_X1 U5697 ( .A1(n6699), .A2(n15503), .ZN(n15267) );
  OR2_X1 U5698 ( .A1(n15077), .A2(n15073), .ZN(n14569) );
  AND2_X1 U5699 ( .A1(n15511), .A2(n15275), .ZN(n15279) );
  NAND2_X1 U5701 ( .A1(n13601), .A2(n5024), .ZN(n16477) );
  AND2_X1 U5702 ( .A1(n4288), .A2(n4287), .ZN(n6080) );
  AOI22_X1 U5703 ( .A1(n3841), .A2(n3784), .B1(n426), .B2(n3840), .ZN(n4324)
         );
  INV_X1 U5704 ( .A(n4493), .ZN(n15862) );
  XNOR2_X1 U5705 ( .A(n15212), .B(n3792), .ZN(n15745) );
  INV_X1 U5706 ( .A(n17710), .ZN(n4156) );
  OR2_X1 U5707 ( .A1(n15154), .A2(n15155), .ZN(n5196) );
  OR2_X1 U5708 ( .A1(n17190), .A2(n424), .ZN(n4241) );
  INV_X1 U5709 ( .A(n4687), .ZN(n17124) );
  AND2_X1 U5712 ( .A1(n6337), .A2(n6336), .ZN(n3529) );
  INV_X1 U5713 ( .A(n18106), .ZN(n17903) );
  OAI21_X1 U5715 ( .B1(n2707), .B2(n18537), .A(n17699), .ZN(n2704) );
  XNOR2_X1 U5717 ( .A(n19701), .B(n18638), .ZN(n2993) );
  INV_X1 U5719 ( .A(n20205), .ZN(n4340) );
  XNOR2_X1 U5720 ( .A(n19465), .B(n18653), .ZN(n18815) );
  OR2_X1 U5721 ( .A1(n17761), .A2(n525), .ZN(n5417) );
  INV_X1 U5722 ( .A(n19480), .ZN(n4976) );
  XNOR2_X1 U5723 ( .A(n19273), .B(n19535), .ZN(n19084) );
  AND2_X1 U5724 ( .A1(n19938), .A2(n506), .ZN(n2487) );
  XNOR2_X1 U5725 ( .A(n19483), .B(n19085), .ZN(n19634) );
  OAI21_X1 U5727 ( .B1(n18406), .B2(n5021), .A(n18706), .ZN(n17778) );
  OR2_X1 U5728 ( .A1(n17862), .A2(n18516), .ZN(n17863) );
  INV_X1 U5730 ( .A(n4569), .ZN(n4306) );
  AOI21_X1 U5731 ( .B1(n20404), .B2(n20549), .A(n3747), .ZN(n19857) );
  AND2_X1 U5732 ( .A1(n20551), .A2(n20405), .ZN(n3747) );
  OR2_X1 U5733 ( .A1(n20401), .A2(n5680), .ZN(n20566) );
  XNOR2_X1 U5734 ( .A(n19479), .B(n19478), .ZN(n20133) );
  XNOR2_X1 U5735 ( .A(n4030), .B(n19492), .ZN(n19493) );
  INV_X1 U5737 ( .A(n23642), .ZN(n2138) );
  XNOR2_X1 U5738 ( .A(n22231), .B(n22230), .ZN(n23177) );
  INV_X1 U5739 ( .A(n23102), .ZN(n22686) );
  INV_X1 U5744 ( .A(n23227), .ZN(n23399) );
  INV_X1 U5745 ( .A(n23289), .ZN(n4950) );
  XNOR2_X1 U5746 ( .A(n6017), .B(n21988), .ZN(n21989) );
  INV_X1 U5748 ( .A(n23702), .ZN(n6099) );
  XNOR2_X1 U5749 ( .A(n22588), .B(n22587), .ZN(n22592) );
  OR2_X1 U5750 ( .A1(n23770), .A2(n23769), .ZN(n6355) );
  OR2_X1 U5751 ( .A1(n4561), .A2(n23611), .ZN(n4560) );
  AOI21_X1 U5752 ( .B1(n4336), .B2(n23803), .A(n2004), .ZN(n2835) );
  XNOR2_X1 U5753 ( .A(n25738), .B(n25921), .ZN(n25563) );
  INV_X1 U5754 ( .A(n7584), .ZN(n7885) );
  OR2_X1 U5755 ( .A1(n8141), .A2(n7560), .ZN(n7565) );
  OR2_X1 U5756 ( .A1(n7840), .A2(n7836), .ZN(n7368) );
  OR2_X1 U5757 ( .A1(n6209), .A2(n7506), .ZN(n7133) );
  OR2_X1 U5758 ( .A1(n7912), .A2(n7911), .ZN(n8286) );
  OR2_X1 U5759 ( .A1(n8018), .A2(n28161), .ZN(n6807) );
  OR2_X1 U5762 ( .A1(n8716), .A2(n8786), .ZN(n7607) );
  INV_X1 U5765 ( .A(n8073), .ZN(n9100) );
  OR2_X1 U5766 ( .A1(n9026), .A2(n9228), .ZN(n3675) );
  INV_X1 U5767 ( .A(n10087), .ZN(n10009) );
  AND2_X1 U5768 ( .A1(n8974), .A2(n8819), .ZN(n6689) );
  OR2_X1 U5770 ( .A1(n9398), .A2(n8983), .ZN(n3139) );
  INV_X1 U5771 ( .A(n10251), .ZN(n5995) );
  XNOR2_X1 U5772 ( .A(n9626), .B(n9754), .ZN(n9683) );
  INV_X1 U5773 ( .A(n11123), .ZN(n11118) );
  INV_X1 U5774 ( .A(n9590), .ZN(n4807) );
  NOR2_X1 U5775 ( .A1(n9034), .A2(n8792), .ZN(n6860) );
  AND2_X1 U5776 ( .A1(n8330), .A2(n9144), .ZN(n2335) );
  XNOR2_X1 U5777 ( .A(n10228), .B(n10184), .ZN(n10046) );
  INV_X1 U5778 ( .A(n8742), .ZN(n2908) );
  INV_X1 U5779 ( .A(n11144), .ZN(n10806) );
  XNOR2_X1 U5780 ( .A(n8063), .B(n8062), .ZN(n11149) );
  XNOR2_X1 U5781 ( .A(n10206), .B(n10205), .ZN(n11240) );
  OAI21_X1 U5782 ( .B1(n12132), .B2(n12266), .A(n12267), .ZN(n5964) );
  INV_X1 U5783 ( .A(n12504), .ZN(n12867) );
  OR2_X1 U5784 ( .A1(n6282), .A2(n6281), .ZN(n6280) );
  OR2_X1 U5785 ( .A1(n12151), .A2(n11856), .ZN(n3796) );
  OR2_X1 U5786 ( .A1(n10771), .A2(n567), .ZN(n2538) );
  OAI21_X1 U5787 ( .B1(n11879), .B2(n11876), .A(n11582), .ZN(n6561) );
  NOR2_X1 U5789 ( .A1(n11297), .A2(n3558), .ZN(n3557) );
  OR2_X1 U5790 ( .A1(n11837), .A2(n3653), .ZN(n3646) );
  XNOR2_X1 U5791 ( .A(n12738), .B(n12632), .ZN(n13220) );
  OR2_X1 U5792 ( .A1(n569), .A2(n10701), .ZN(n2217) );
  INV_X1 U5793 ( .A(n14126), .ZN(n4897) );
  OR2_X1 U5794 ( .A1(n29089), .A2(n13589), .ZN(n2144) );
  XNOR2_X1 U5795 ( .A(n6052), .B(n13439), .ZN(n14373) );
  XNOR2_X1 U5796 ( .A(n13438), .B(n13437), .ZN(n6052) );
  XNOR2_X1 U5799 ( .A(n12419), .B(n12418), .ZN(n14398) );
  XNOR2_X1 U5800 ( .A(n12757), .B(n12756), .ZN(n14464) );
  INV_X1 U5801 ( .A(n16090), .ZN(n16282) );
  XNOR2_X1 U5802 ( .A(n11203), .B(n11202), .ZN(n14106) );
  OR2_X1 U5804 ( .A1(n13871), .A2(n13706), .ZN(n3435) );
  XNOR2_X1 U5805 ( .A(n12375), .B(n12376), .ZN(n14408) );
  INV_X1 U5806 ( .A(n13877), .ZN(n4509) );
  XNOR2_X1 U5807 ( .A(n2172), .B(n13462), .ZN(n2171) );
  XNOR2_X1 U5808 ( .A(n6297), .B(n6298), .ZN(n2173) );
  XNOR2_X1 U5811 ( .A(n13273), .B(n4501), .ZN(n11543) );
  OR2_X1 U5812 ( .A1(n5531), .A2(n13730), .ZN(n3799) );
  OR2_X1 U5813 ( .A1(n14321), .A2(n14320), .ZN(n6794) );
  OR3_X1 U5814 ( .A1(n29306), .A2(n14165), .A3(n14481), .ZN(n3408) );
  INV_X1 U5815 ( .A(n16567), .ZN(n15723) );
  INV_X1 U5816 ( .A(n15135), .ZN(n15252) );
  OR2_X1 U5817 ( .A1(n15025), .A2(n15444), .ZN(n4491) );
  AND2_X1 U5818 ( .A1(n14111), .A2(n2727), .ZN(n2726) );
  AND2_X1 U5819 ( .A1(n14484), .A2(n14166), .ZN(n4074) );
  OR2_X1 U5820 ( .A1(n14896), .A2(n5025), .ZN(n6851) );
  XNOR2_X1 U5821 ( .A(n4765), .B(n4766), .ZN(n17315) );
  INV_X1 U5822 ( .A(n17492), .ZN(n17496) );
  INV_X1 U5823 ( .A(n14846), .ZN(n5614) );
  OR2_X1 U5824 ( .A1(n15091), .A2(n15090), .ZN(n3022) );
  INV_X1 U5825 ( .A(n16937), .ZN(n17340) );
  XNOR2_X1 U5827 ( .A(n15817), .B(n15790), .ZN(n5621) );
  XNOR2_X1 U5829 ( .A(n16012), .B(n15977), .ZN(n16224) );
  XNOR2_X1 U5830 ( .A(n14561), .B(n14562), .ZN(n17269) );
  NOR2_X1 U5832 ( .A1(n28768), .A2(n17012), .ZN(n17423) );
  XNOR2_X1 U5833 ( .A(n15575), .B(n6319), .ZN(n15577) );
  OR2_X1 U5834 ( .A1(n17469), .A2(n17516), .ZN(n2610) );
  XNOR2_X1 U5835 ( .A(n16050), .B(n259), .ZN(n4588) );
  INV_X1 U5836 ( .A(n16918), .ZN(n17314) );
  XNOR2_X1 U5837 ( .A(n15883), .B(n15882), .ZN(n17567) );
  INV_X1 U5838 ( .A(n17484), .ZN(n4271) );
  XNOR2_X1 U5840 ( .A(n2671), .B(n16610), .ZN(n17110) );
  XNOR2_X1 U5841 ( .A(n1977), .B(n16140), .ZN(n2671) );
  XNOR2_X1 U5842 ( .A(n16090), .B(n5892), .ZN(n13926) );
  AND2_X1 U5843 ( .A1(n29406), .A2(n17110), .ZN(n17473) );
  OR2_X1 U5844 ( .A1(n17570), .A2(n423), .ZN(n4157) );
  XNOR2_X1 U5845 ( .A(n6870), .B(n6869), .ZN(n17143) );
  AND2_X1 U5846 ( .A1(n17528), .A2(n16706), .ZN(n6161) );
  XNOR2_X1 U5847 ( .A(n15860), .B(n15861), .ZN(n4316) );
  INV_X1 U5848 ( .A(n17355), .ZN(n4283) );
  INV_X1 U5850 ( .A(n17553), .ZN(n16913) );
  INV_X1 U5851 ( .A(n17524), .ZN(n4979) );
  INV_X1 U5853 ( .A(n17361), .ZN(n17046) );
  OR2_X1 U5854 ( .A1(n17546), .A2(n211), .ZN(n2375) );
  INV_X1 U5855 ( .A(n18035), .ZN(n2500) );
  XNOR2_X1 U5856 ( .A(n19445), .B(n3255), .ZN(n4339) );
  XNOR2_X1 U5857 ( .A(n18691), .B(n4029), .ZN(n3255) );
  INV_X1 U5858 ( .A(n20221), .ZN(n20168) );
  XNOR2_X1 U5859 ( .A(n17334), .B(n17333), .ZN(n20406) );
  INV_X1 U5860 ( .A(n20547), .ZN(n6261) );
  INV_X1 U5861 ( .A(n21092), .ZN(n20145) );
  XNOR2_X1 U5862 ( .A(n19648), .B(n19649), .ZN(n20282) );
  INV_X1 U5863 ( .A(n20475), .ZN(n5408) );
  INV_X1 U5864 ( .A(n415), .ZN(n5935) );
  XNOR2_X1 U5865 ( .A(n19633), .B(n6535), .ZN(n6534) );
  BUF_X1 U5866 ( .A(n20176), .Z(n20171) );
  AND2_X1 U5868 ( .A1(n28658), .A2(n29145), .ZN(n20084) );
  NOR2_X1 U5869 ( .A1(n20176), .A2(n6114), .ZN(n19052) );
  OR2_X1 U5870 ( .A1(n20099), .A2(n18887), .ZN(n20042) );
  AND2_X1 U5871 ( .A1(n5056), .A2(n20099), .ZN(n2715) );
  INV_X1 U5872 ( .A(n29146), .ZN(n18837) );
  INV_X1 U5873 ( .A(n20334), .ZN(n20005) );
  INV_X1 U5874 ( .A(n20406), .ZN(n20556) );
  XNOR2_X1 U5875 ( .A(n16869), .B(n5062), .ZN(n16870) );
  XNOR2_X1 U5876 ( .A(n5539), .B(n5538), .ZN(n20319) );
  AND2_X1 U5877 ( .A1(n20388), .A2(n20539), .ZN(n19958) );
  OR2_X1 U5878 ( .A1(n19820), .A2(n20539), .ZN(n19959) );
  AND2_X1 U5879 ( .A1(n20293), .A2(n20125), .ZN(n19973) );
  INV_X1 U5880 ( .A(n20039), .ZN(n20087) );
  XNOR2_X1 U5881 ( .A(n18734), .B(n18733), .ZN(n2735) );
  XNOR2_X1 U5882 ( .A(n4838), .B(n4030), .ZN(n6701) );
  OAI21_X1 U5884 ( .B1(n20444), .B2(n3247), .A(n3246), .ZN(n20448) );
  INV_X1 U5885 ( .A(n4567), .ZN(n4570) );
  OR2_X1 U5886 ( .A1(n20153), .A2(n28188), .ZN(n5034) );
  INV_X1 U5887 ( .A(n22386), .ZN(n21325) );
  INV_X1 U5889 ( .A(n3838), .ZN(n20841) );
  XNOR2_X1 U5891 ( .A(n6837), .B(n6836), .ZN(n23637) );
  XNOR2_X1 U5892 ( .A(n22572), .B(n22573), .ZN(n23827) );
  XNOR2_X1 U5893 ( .A(n21386), .B(n21385), .ZN(n23338) );
  XNOR2_X1 U5894 ( .A(n21911), .B(n21910), .ZN(n23492) );
  OR2_X1 U5895 ( .A1(n23149), .A2(n23461), .ZN(n4892) );
  INV_X1 U5896 ( .A(n23493), .ZN(n6608) );
  OR2_X1 U5898 ( .A1(n23741), .A2(n22944), .ZN(n3149) );
  INV_X1 U5899 ( .A(n23564), .ZN(n22995) );
  INV_X1 U5900 ( .A(n4003), .ZN(n23761) );
  INV_X1 U5903 ( .A(n23637), .ZN(n23557) );
  INV_X1 U5904 ( .A(n2141), .ZN(n23397) );
  OAI21_X1 U5905 ( .B1(n4256), .B2(n4255), .A(n22996), .ZN(n4254) );
  OR2_X1 U5906 ( .A1(n23646), .A2(n23645), .ZN(n3723) );
  NOR2_X1 U5907 ( .A1(n23529), .A2(n23531), .ZN(n5482) );
  NAND2_X1 U5908 ( .A1(n23677), .A2(n3901), .ZN(n24808) );
  OR2_X1 U5909 ( .A1(n23360), .A2(n23673), .ZN(n2575) );
  AOI21_X1 U5910 ( .B1(n6267), .B2(n24404), .A(n24405), .ZN(n23306) );
  INV_X1 U5911 ( .A(n3797), .ZN(n6267) );
  INV_X1 U5912 ( .A(n6110), .ZN(n25179) );
  XNOR2_X1 U5913 ( .A(n25398), .B(n25249), .ZN(n25069) );
  XNOR2_X1 U5915 ( .A(n25907), .B(n25906), .ZN(n26510) );
  XNOR2_X1 U5916 ( .A(n3837), .B(n25191), .ZN(n25915) );
  NAND2_X1 U5917 ( .A1(n24150), .A2(n5922), .ZN(n25546) );
  OAI22_X1 U5918 ( .A1(n5137), .A2(n5138), .B1(n24612), .B2(n24611), .ZN(n5136) );
  NAND2_X1 U5919 ( .A1(n24614), .A2(n29109), .ZN(n5138) );
  XNOR2_X1 U5920 ( .A(n23244), .B(n23243), .ZN(n23862) );
  INV_X1 U5921 ( .A(n25418), .ZN(n26792) );
  INV_X1 U5922 ( .A(n26278), .ZN(n26798) );
  XNOR2_X1 U5923 ( .A(n24923), .B(n24925), .ZN(n5754) );
  OR2_X1 U5924 ( .A1(n26868), .A2(n27110), .ZN(n26310) );
  AND2_X1 U5926 ( .A1(n7162), .A2(n7320), .ZN(n7279) );
  OR2_X1 U5927 ( .A1(n7865), .A2(n7308), .ZN(n3664) );
  OR2_X1 U5928 ( .A1(n7787), .A2(n7330), .ZN(n7293) );
  INV_X1 U5929 ( .A(n7591), .ZN(n7957) );
  OAI21_X1 U5931 ( .B1(n7303), .B2(n7305), .A(n7237), .ZN(n5173) );
  OR2_X1 U5932 ( .A1(n8525), .A2(n8687), .ZN(n9223) );
  NAND2_X1 U5933 ( .A1(n6316), .A2(n8898), .ZN(n6318) );
  OAI21_X1 U5934 ( .B1(n8840), .B2(n8839), .A(n8961), .ZN(n3182) );
  OR2_X1 U5935 ( .A1(n8842), .A2(n605), .ZN(n3181) );
  INV_X1 U5936 ( .A(n10372), .ZN(n10201) );
  OR2_X1 U5937 ( .A1(n8762), .A2(n9566), .ZN(n7273) );
  INV_X1 U5938 ( .A(n8472), .ZN(n6662) );
  OAI21_X1 U5940 ( .B1(n6344), .B2(n9042), .A(n8110), .ZN(n7159) );
  XNOR2_X1 U5943 ( .A(n9786), .B(n9785), .ZN(n5984) );
  XNOR2_X1 U5944 ( .A(n8649), .B(n10334), .ZN(n11144) );
  XNOR2_X1 U5945 ( .A(n9639), .B(n10426), .ZN(n10189) );
  XNOR2_X1 U5946 ( .A(n10265), .B(n10302), .ZN(n9961) );
  AND2_X1 U5947 ( .A1(n7413), .A2(n7411), .ZN(n2676) );
  OR2_X1 U5948 ( .A1(n8407), .A2(n3297), .ZN(n3296) );
  XNOR2_X1 U5949 ( .A(n10007), .B(n4714), .ZN(n10424) );
  OR2_X1 U5950 ( .A1(n9224), .A2(n8685), .ZN(n5959) );
  OR2_X1 U5951 ( .A1(n8802), .A2(n8801), .ZN(n8803) );
  INV_X1 U5952 ( .A(n11335), .ZN(n11341) );
  NOR2_X1 U5954 ( .A1(n3804), .A2(n10989), .ZN(n3803) );
  AND2_X1 U5955 ( .A1(n10775), .A2(n6108), .ZN(n5706) );
  XNOR2_X1 U5956 ( .A(n9683), .B(n10027), .ZN(n4589) );
  INV_X1 U5957 ( .A(n11056), .ZN(n10851) );
  INV_X1 U5958 ( .A(n11350), .ZN(n3161) );
  INV_X1 U5959 ( .A(n333), .ZN(n6816) );
  OR2_X1 U5960 ( .A1(n10911), .A2(n10913), .ZN(n5904) );
  XNOR2_X1 U5961 ( .A(n9811), .B(n9887), .ZN(n2662) );
  INV_X1 U5962 ( .A(n11090), .ZN(n5277) );
  XNOR2_X1 U5963 ( .A(n6133), .B(n6135), .ZN(n11022) );
  XNOR2_X1 U5964 ( .A(n5414), .B(n5413), .ZN(n10937) );
  XNOR2_X1 U5965 ( .A(n9683), .B(n9416), .ZN(n5413) );
  XNOR2_X1 U5966 ( .A(n5411), .B(n5410), .ZN(n5414) );
  INV_X1 U5967 ( .A(n10936), .ZN(n11002) );
  INV_X1 U5968 ( .A(n10620), .ZN(n11099) );
  OR2_X1 U5969 ( .A1(n11056), .A2(n10855), .ZN(n10856) );
  OR2_X1 U5970 ( .A1(n591), .A2(n2211), .ZN(n2210) );
  XNOR2_X1 U5972 ( .A(n9350), .B(n10046), .ZN(n5860) );
  INV_X1 U5973 ( .A(n6108), .ZN(n5710) );
  AND2_X1 U5974 ( .A1(n11933), .A2(n12070), .ZN(n11595) );
  INV_X1 U5975 ( .A(n12559), .ZN(n13034) );
  XNOR2_X1 U5976 ( .A(n12377), .B(n4277), .ZN(n12379) );
  INV_X1 U5977 ( .A(n12788), .ZN(n4277) );
  OR2_X1 U5978 ( .A1(n12080), .A2(n29499), .ZN(n5715) );
  INV_X1 U5979 ( .A(n285), .ZN(n12322) );
  INV_X1 U5981 ( .A(n12472), .ZN(n13231) );
  INV_X1 U5982 ( .A(n12236), .ZN(n11979) );
  AND2_X1 U5985 ( .A1(n12330), .A2(n6431), .ZN(n3281) );
  OR2_X1 U5986 ( .A1(n12003), .A2(n12004), .ZN(n2603) );
  INV_X1 U5987 ( .A(n13538), .ZN(n12885) );
  XNOR2_X1 U5988 ( .A(n12542), .B(n13493), .ZN(n13315) );
  XNOR2_X1 U5989 ( .A(n13406), .B(n13538), .ZN(n13027) );
  INV_X1 U5990 ( .A(n13872), .ZN(n14428) );
  INV_X1 U5992 ( .A(n11676), .ZN(n11674) );
  XNOR2_X1 U5994 ( .A(n12658), .B(n12723), .ZN(n13243) );
  OR2_X1 U5998 ( .A1(n6581), .A2(n28201), .ZN(n6519) );
  INV_X1 U5999 ( .A(n12978), .ZN(n4375) );
  INV_X1 U6000 ( .A(n28805), .ZN(n4433) );
  NOR2_X1 U6001 ( .A1(n14475), .A2(n13936), .ZN(n14473) );
  OR2_X1 U6002 ( .A1(n14480), .A2(n14157), .ZN(n13847) );
  XNOR2_X1 U6003 ( .A(n4199), .B(n4198), .ZN(n14487) );
  XNOR2_X1 U6004 ( .A(n4200), .B(n12065), .ZN(n4199) );
  XNOR2_X1 U6005 ( .A(n12064), .B(n2916), .ZN(n4200) );
  INV_X1 U6006 ( .A(n14450), .ZN(n2972) );
  XNOR2_X1 U6007 ( .A(n11669), .B(n3870), .ZN(n5805) );
  AOI21_X1 U6008 ( .B1(n14232), .B2(n14102), .A(n4054), .ZN(n14104) );
  AND2_X1 U6009 ( .A1(n4056), .A2(n14106), .ZN(n2608) );
  INV_X1 U6010 ( .A(n15431), .ZN(n15031) );
  XNOR2_X1 U6012 ( .A(n13338), .B(n2570), .ZN(n11838) );
  XNOR2_X1 U6013 ( .A(n4474), .B(n13035), .ZN(n2570) );
  OR2_X1 U6014 ( .A1(n15494), .A2(n14702), .ZN(n6246) );
  XNOR2_X1 U6015 ( .A(n12635), .B(n12636), .ZN(n14177) );
  OR2_X1 U6016 ( .A1(n14498), .A2(n29036), .ZN(n13973) );
  XNOR2_X1 U6017 ( .A(n12963), .B(n12964), .ZN(n14123) );
  AND2_X1 U6019 ( .A1(n15053), .A2(n15261), .ZN(n2161) );
  INV_X1 U6020 ( .A(n15310), .ZN(n15315) );
  NOR2_X1 U6021 ( .A1(n4088), .A2(n4897), .ZN(n4896) );
  AND2_X1 U6022 ( .A1(n14262), .A2(n14259), .ZN(n13747) );
  INV_X1 U6025 ( .A(n15515), .ZN(n6293) );
  OAI211_X1 U6026 ( .C1(n15249), .C2(n15247), .A(n13715), .B(n13714), .ZN(
        n16126) );
  OR2_X1 U6027 ( .A1(n15053), .A2(n14761), .ZN(n6391) );
  INV_X1 U6028 ( .A(n4811), .ZN(n16384) );
  INV_X1 U6029 ( .A(n15073), .ZN(n14571) );
  INV_X1 U6031 ( .A(n4992), .ZN(n6674) );
  OR2_X1 U6032 ( .A1(n15266), .A2(n14922), .ZN(n5722) );
  INV_X1 U6033 ( .A(n3673), .ZN(n4492) );
  OR2_X1 U6034 ( .A1(n14598), .A2(n14762), .ZN(n3550) );
  XNOR2_X1 U6035 ( .A(n3856), .B(n16373), .ZN(n16640) );
  XNOR2_X1 U6036 ( .A(n16084), .B(n2117), .ZN(n16643) );
  OR2_X1 U6039 ( .A1(n14728), .A2(n15395), .ZN(n3605) );
  OR2_X1 U6040 ( .A1(n13519), .A2(n14884), .ZN(n3487) );
  INV_X1 U6041 ( .A(n17298), .ZN(n5430) );
  NOR2_X1 U6042 ( .A1(n5471), .A2(n17143), .ZN(n17087) );
  XNOR2_X1 U6043 ( .A(n15106), .B(n16229), .ZN(n16191) );
  BUF_X1 U6044 ( .A(n14871), .Z(n17395) );
  BUF_X1 U6045 ( .A(n16679), .Z(n17282) );
  AND2_X1 U6047 ( .A1(n4414), .A2(n4413), .ZN(n17828) );
  AOI21_X1 U6048 ( .B1(n17074), .B2(n17505), .A(n17829), .ZN(n4414) );
  INV_X1 U6049 ( .A(n17556), .ZN(n16916) );
  INV_X1 U6050 ( .A(n538), .ZN(n4314) );
  OR2_X1 U6051 ( .A1(n29547), .A2(n18028), .ZN(n3932) );
  OR2_X1 U6052 ( .A1(n18410), .A2(n18121), .ZN(n18416) );
  XNOR2_X1 U6054 ( .A(n5859), .B(n16658), .ZN(n17438) );
  NAND2_X1 U6055 ( .A1(n17081), .A2(n6067), .ZN(n18589) );
  INV_X1 U6056 ( .A(n17151), .ZN(n6067) );
  NOR2_X1 U6057 ( .A1(n28194), .A2(n5891), .ZN(n16973) );
  OR2_X1 U6059 ( .A1(n2825), .A2(n5891), .ZN(n2827) );
  AND2_X1 U6060 ( .A1(n18305), .A2(n18306), .ZN(n6576) );
  NAND2_X1 U6062 ( .A1(n4830), .A2(n4829), .ZN(n17834) );
  OAI211_X1 U6064 ( .C1(n17518), .C2(n17470), .A(n6889), .B(n17516), .ZN(
        n17084) );
  AND2_X1 U6065 ( .A1(n17017), .A2(n17016), .ZN(n4866) );
  AND3_X1 U6066 ( .A1(n17844), .A2(n18241), .A3(n3848), .ZN(n3847) );
  AND3_X1 U6067 ( .A1(n524), .A2(n18018), .A3(n1888), .ZN(n6429) );
  OR2_X1 U6068 ( .A1(n18251), .A2(n1888), .ZN(n18254) );
  AND2_X1 U6069 ( .A1(n18216), .A2(n18215), .ZN(n4824) );
  OR2_X1 U6070 ( .A1(n17596), .A2(n18227), .ZN(n5747) );
  OR2_X1 U6071 ( .A1(n18261), .A2(n18324), .ZN(n17986) );
  OR2_X1 U6072 ( .A1(n17815), .A2(n4762), .ZN(n4761) );
  OR2_X1 U6073 ( .A1(n17266), .A2(n29298), .ZN(n16971) );
  OAI21_X1 U6074 ( .B1(n18445), .B2(n4928), .A(n4927), .ZN(n19252) );
  AOI21_X1 U6075 ( .B1(n18178), .B2(n4930), .A(n4929), .ZN(n4928) );
  XNOR2_X1 U6076 ( .A(n19389), .B(n3385), .ZN(n19048) );
  XNOR2_X1 U6077 ( .A(n6445), .B(n4883), .ZN(n19026) );
  INV_X1 U6078 ( .A(n19103), .ZN(n6445) );
  OR2_X1 U6080 ( .A1(n17693), .A2(n18078), .ZN(n18079) );
  OAI22_X1 U6081 ( .A1(n18311), .A2(n17918), .B1(n6225), .B2(n18355), .ZN(
        n17922) );
  NOR2_X1 U6082 ( .A1(n2776), .A2(n18123), .ZN(n2775) );
  AND2_X1 U6083 ( .A1(n2778), .A2(n17818), .ZN(n2776) );
  AND2_X1 U6084 ( .A1(n4210), .A2(n4212), .ZN(n3402) );
  XNOR2_X1 U6085 ( .A(n19152), .B(n4746), .ZN(n4745) );
  AND2_X1 U6086 ( .A1(n18376), .A2(n18380), .ZN(n17166) );
  XNOR2_X1 U6087 ( .A(n19496), .B(n28516), .ZN(n19402) );
  XNOR2_X1 U6088 ( .A(n19553), .B(n19552), .ZN(n20451) );
  INV_X1 U6090 ( .A(n18691), .ZN(n4030) );
  OR2_X1 U6092 ( .A1(n17756), .A2(n18243), .ZN(n2771) );
  INV_X1 U6093 ( .A(n18653), .ZN(n19568) );
  AND2_X1 U6094 ( .A1(n5000), .A2(n21425), .ZN(n20896) );
  AND2_X1 U6095 ( .A1(n21087), .A2(n5827), .ZN(n20895) );
  XNOR2_X1 U6096 ( .A(n19543), .B(n2993), .ZN(n19544) );
  OAI22_X1 U6097 ( .A1(n19174), .A2(n5491), .B1(n19692), .B2(n5490), .ZN(
        n19176) );
  INV_X1 U6098 ( .A(n5225), .ZN(n5303) );
  NOR2_X1 U6099 ( .A1(n499), .A2(n6834), .ZN(n2797) );
  AND2_X1 U6100 ( .A1(n19752), .A2(n5937), .ZN(n19781) );
  INV_X1 U6101 ( .A(n19761), .ZN(n20069) );
  OR2_X1 U6102 ( .A1(n20089), .A2(n29114), .ZN(n6399) );
  OR2_X1 U6103 ( .A1(n5684), .A2(n20713), .ZN(n20714) );
  OR2_X1 U6104 ( .A1(n20715), .A2(n5684), .ZN(n5683) );
  AND2_X1 U6106 ( .A1(n20451), .A2(n19554), .ZN(n21063) );
  OR2_X1 U6107 ( .A1(n28491), .A2(n21359), .ZN(n4167) );
  OR2_X1 U6108 ( .A1(n19935), .A2(n20607), .ZN(n19936) );
  INV_X1 U6109 ( .A(n20647), .ZN(n5783) );
  INV_X1 U6110 ( .A(n2081), .ZN(n4096) );
  NAND2_X1 U6111 ( .A1(n20229), .A2(n29426), .ZN(n3852) );
  INV_X1 U6112 ( .A(n21642), .ZN(n21402) );
  AND2_X1 U6113 ( .A1(n5778), .A2(n20088), .ZN(n18749) );
  INV_X1 U6114 ( .A(n3238), .ZN(n5928) );
  AND2_X1 U6115 ( .A1(n4242), .A2(n19974), .ZN(n3243) );
  INV_X1 U6116 ( .A(n21253), .ZN(n2125) );
  OR2_X1 U6117 ( .A1(n21078), .A2(n495), .ZN(n21076) );
  AND2_X1 U6118 ( .A1(n21075), .A2(n21071), .ZN(n2992) );
  INV_X1 U6119 ( .A(n21075), .ZN(n2989) );
  OR2_X1 U6120 ( .A1(n21052), .A2(n21051), .ZN(n3039) );
  OR2_X1 U6122 ( .A1(n19921), .A2(n28894), .ZN(n20257) );
  OAI211_X1 U6123 ( .C1(n21818), .C2(n20108), .A(n5124), .B(n5123), .ZN(n22099) );
  OR2_X1 U6124 ( .A1(n20043), .A2(n20151), .ZN(n4409) );
  NOR2_X1 U6126 ( .A1(n20152), .A2(n18887), .ZN(n18831) );
  INV_X1 U6127 ( .A(n21875), .ZN(n22093) );
  OR2_X1 U6128 ( .A1(n20557), .A2(n20556), .ZN(n3193) );
  INV_X1 U6129 ( .A(n19743), .ZN(n4362) );
  AND2_X1 U6130 ( .A1(n5443), .A2(n5442), .ZN(n5441) );
  OR2_X1 U6131 ( .A1(n29530), .A2(n21309), .ZN(n5442) );
  INV_X1 U6132 ( .A(n21567), .ZN(n6247) );
  XNOR2_X1 U6134 ( .A(n22337), .B(n6504), .ZN(n22852) );
  OR2_X1 U6135 ( .A1(n21542), .A2(n20393), .ZN(n2725) );
  XNOR2_X1 U6136 ( .A(n22811), .B(n22363), .ZN(n21454) );
  AND2_X1 U6137 ( .A1(n23768), .A2(n23765), .ZN(n5355) );
  XNOR2_X1 U6138 ( .A(n22710), .B(n22320), .ZN(n22545) );
  OAI21_X1 U6139 ( .B1(n481), .B2(n29602), .A(n22962), .ZN(n2367) );
  INV_X1 U6140 ( .A(n22923), .ZN(n4229) );
  XNOR2_X1 U6141 ( .A(n22882), .B(n3321), .ZN(n3091) );
  OAI21_X1 U6142 ( .B1(n20955), .B2(n20802), .A(n2296), .ZN(n21102) );
  OAI21_X1 U6143 ( .B1(n21449), .B2(n21673), .A(n3132), .ZN(n3131) );
  OAI21_X1 U6144 ( .B1(n20830), .B2(n20831), .A(n412), .ZN(n20832) );
  INV_X1 U6145 ( .A(n21675), .ZN(n3132) );
  OR2_X1 U6147 ( .A1(n21572), .A2(n21571), .ZN(n3562) );
  OR2_X1 U6148 ( .A1(n20950), .A2(n21538), .ZN(n5878) );
  XNOR2_X1 U6149 ( .A(n22896), .B(n22692), .ZN(n22502) );
  OR2_X1 U6150 ( .A1(n21202), .A2(n21509), .ZN(n3288) );
  NAND2_X1 U6152 ( .A1(n21393), .A2(n21392), .ZN(n2395) );
  AOI22_X1 U6153 ( .A1(n4143), .A2(n20031), .B1(n3588), .B2(n21638), .ZN(
        n20035) );
  NOR2_X1 U6154 ( .A1(n21392), .A2(n21632), .ZN(n3588) );
  XNOR2_X1 U6155 ( .A(n28449), .B(n3451), .ZN(n5840) );
  OR2_X1 U6156 ( .A1(n21261), .A2(n21718), .ZN(n3407) );
  OR2_X1 U6157 ( .A1(n28789), .A2(n21497), .ZN(n6750) );
  OR2_X1 U6158 ( .A1(n20928), .A2(n21198), .ZN(n4566) );
  INV_X1 U6160 ( .A(n5080), .ZN(n24092) );
  INV_X1 U6161 ( .A(n23492), .ZN(n23791) );
  XNOR2_X1 U6162 ( .A(n22466), .B(n22465), .ZN(n23392) );
  OR2_X1 U6163 ( .A1(n23127), .A2(n23126), .ZN(n23128) );
  NOR2_X1 U6165 ( .A1(n24120), .A2(n29726), .ZN(n23888) );
  INV_X1 U6166 ( .A(n24305), .ZN(n24365) );
  OAI21_X1 U6167 ( .B1(n24673), .B2(n23334), .A(n2130), .ZN(n25444) );
  AND2_X1 U6168 ( .A1(n24323), .A2(n404), .ZN(n4025) );
  AND2_X1 U6169 ( .A1(n24547), .A2(n24160), .ZN(n2820) );
  XNOR2_X1 U6170 ( .A(n24254), .B(n24255), .ZN(n25406) );
  XNOR2_X1 U6171 ( .A(n25191), .B(n4861), .ZN(n24784) );
  AND3_X1 U6172 ( .A1(n5479), .A2(n5478), .A3(n220), .ZN(n23698) );
  OR2_X1 U6173 ( .A1(n24817), .A2(n24809), .ZN(n5479) );
  OR2_X1 U6174 ( .A1(n24237), .A2(n24195), .ZN(n24571) );
  OR2_X1 U6175 ( .A1(n24551), .A2(n24552), .ZN(n5509) );
  OR2_X1 U6176 ( .A1(n5094), .A2(n24593), .ZN(n4690) );
  INV_X1 U6177 ( .A(n24257), .ZN(n2175) );
  XNOR2_X1 U6178 ( .A(n28465), .B(n3493), .ZN(n5431) );
  XNOR2_X1 U6179 ( .A(n5146), .B(n26899), .ZN(n25140) );
  OR2_X1 U6182 ( .A1(n24972), .A2(n24256), .ZN(n3121) );
  OAI21_X1 U6183 ( .B1(n24716), .B2(n4136), .A(n4135), .ZN(n23869) );
  XNOR2_X1 U6184 ( .A(n25546), .B(n26093), .ZN(n26007) );
  NOR2_X1 U6185 ( .A1(n5105), .A2(n24227), .ZN(n5104) );
  NAND2_X1 U6186 ( .A1(n2880), .A2(n2878), .ZN(n4161) );
  INV_X1 U6187 ( .A(n24237), .ZN(n6239) );
  AND2_X1 U6189 ( .A1(n24711), .A2(n24713), .ZN(n23070) );
  XNOR2_X1 U6190 ( .A(n26083), .B(n26053), .ZN(n25533) );
  XNOR2_X1 U6193 ( .A(n26101), .B(n25411), .ZN(n2812) );
  INV_X1 U6194 ( .A(n24797), .ZN(n25786) );
  XNOR2_X1 U6195 ( .A(n25577), .B(n25282), .ZN(n25875) );
  XNOR2_X1 U6196 ( .A(n25430), .B(n25369), .ZN(n25898) );
  OR2_X1 U6197 ( .A1(n26466), .A2(n26191), .ZN(n26192) );
  AND2_X1 U6198 ( .A1(n29028), .A2(n25406), .ZN(n6685) );
  XNOR2_X1 U6199 ( .A(n1958), .B(n25311), .ZN(n4643) );
  AND2_X1 U6200 ( .A1(n26581), .A2(n26927), .ZN(n4401) );
  INV_X1 U6201 ( .A(n26927), .ZN(n4402) );
  XNOR2_X1 U6202 ( .A(n24982), .B(n24983), .ZN(n26385) );
  OR2_X1 U6203 ( .A1(n27055), .A2(n27902), .ZN(n26851) );
  XNOR2_X1 U6205 ( .A(n3168), .B(n25712), .ZN(n27063) );
  AND2_X1 U6207 ( .A1(n29524), .A2(n29058), .ZN(n27001) );
  OR2_X1 U6208 ( .A1(n26623), .A2(n27050), .ZN(n26246) );
  NOR2_X1 U6209 ( .A1(n28468), .A2(n27548), .ZN(n2617) );
  INV_X1 U6210 ( .A(n27287), .ZN(n27281) );
  OAI21_X1 U6211 ( .B1(n29022), .B2(n27772), .A(n6419), .ZN(n6418) );
  AND2_X1 U6212 ( .A1(n7584), .A2(n7303), .ZN(n3004) );
  INV_X1 U6213 ( .A(n7257), .ZN(n6209) );
  AND2_X1 U6214 ( .A1(n29639), .A2(n7488), .ZN(n7664) );
  INV_X1 U6215 ( .A(n7585), .ZN(n2224) );
  NOR2_X1 U6216 ( .A1(n7580), .A2(n7071), .ZN(n2223) );
  INV_X1 U6217 ( .A(n8724), .ZN(n10241) );
  OR2_X1 U6218 ( .A1(n8720), .A2(n8787), .ZN(n4322) );
  AND2_X1 U6219 ( .A1(n8810), .A2(n8523), .ZN(n3225) );
  NAND3_X1 U6220 ( .A1(n3094), .A2(n8283), .A3(n3093), .ZN(n8956) );
  OR2_X1 U6221 ( .A1(n8285), .A2(n8284), .ZN(n3093) );
  INV_X1 U6222 ( .A(n8658), .ZN(n8501) );
  AND2_X1 U6223 ( .A1(n2740), .A2(n2739), .ZN(n7302) );
  OR2_X1 U6224 ( .A1(n9004), .A2(n9184), .ZN(n3755) );
  OR3_X1 U6226 ( .A1(n9184), .A2(n8782), .A3(n9009), .ZN(n7755) );
  OR2_X1 U6227 ( .A1(n8642), .A2(n8984), .ZN(n9176) );
  OR2_X1 U6229 ( .A1(n8752), .A2(n8751), .ZN(n3050) );
  OR2_X1 U6232 ( .A1(n6590), .A2(n5944), .ZN(n4730) );
  NAND4_X1 U6233 ( .A1(n8076), .A2(n2698), .A3(n8075), .A4(n8074), .ZN(n10028)
         );
  INV_X1 U6234 ( .A(n9097), .ZN(n2698) );
  AND2_X1 U6235 ( .A1(n8666), .A2(n8490), .ZN(n9097) );
  OAI211_X1 U6237 ( .C1(n610), .C2(n8897), .A(n3274), .B(n2980), .ZN(n3273) );
  OR2_X1 U6239 ( .A1(n8888), .A2(n8886), .ZN(n8010) );
  XNOR2_X1 U6240 ( .A(n9794), .B(n2677), .ZN(n9658) );
  OR2_X1 U6241 ( .A1(n9026), .A2(n597), .ZN(n3780) );
  XNOR2_X1 U6242 ( .A(n10144), .B(n1225), .ZN(n4507) );
  OR2_X1 U6243 ( .A1(n11166), .A2(n10820), .ZN(n2103) );
  OR2_X1 U6244 ( .A1(n8327), .A2(n606), .ZN(n3609) );
  AND2_X1 U6245 ( .A1(n9120), .A2(n9119), .ZN(n4969) );
  MUX2_X1 U6246 ( .A(n9149), .B(n11), .S(n9146), .Z(n9155) );
  AND2_X1 U6247 ( .A1(n8338), .A2(n8337), .ZN(n2712) );
  XNOR2_X1 U6248 ( .A(n9296), .B(n9977), .ZN(n5268) );
  XNOR2_X1 U6249 ( .A(n9931), .B(n4713), .ZN(n10303) );
  OR2_X1 U6250 ( .A1(n8753), .A2(n9132), .ZN(n8341) );
  OR2_X1 U6251 ( .A1(n8631), .A2(n8490), .ZN(n8494) );
  XNOR2_X1 U6252 ( .A(n10227), .B(n9899), .ZN(n9825) );
  OR2_X1 U6253 ( .A1(n8852), .A2(n9079), .ZN(n7493) );
  OR2_X1 U6254 ( .A1(n8851), .A2(n8724), .ZN(n7491) );
  OR2_X1 U6255 ( .A1(n11351), .A2(n11350), .ZN(n11190) );
  INV_X1 U6256 ( .A(n11165), .ZN(n9686) );
  NOR2_X1 U6257 ( .A1(n8422), .A2(n10821), .ZN(n2127) );
  OR2_X1 U6258 ( .A1(n10522), .A2(n279), .ZN(n11276) );
  INV_X1 U6259 ( .A(n10051), .ZN(n10730) );
  OR2_X1 U6260 ( .A1(n5366), .A2(n28208), .ZN(n4902) );
  AND2_X1 U6262 ( .A1(n11435), .A2(n12266), .ZN(n2466) );
  XNOR2_X1 U6264 ( .A(n1990), .B(n8845), .ZN(n11335) );
  INV_X1 U6265 ( .A(n12206), .ZN(n4038) );
  OR2_X1 U6266 ( .A1(n4037), .A2(n12109), .ZN(n2683) );
  INV_X1 U6267 ( .A(n11671), .ZN(n5079) );
  OR2_X1 U6268 ( .A1(n11165), .A2(n11053), .ZN(n11309) );
  AND2_X1 U6269 ( .A1(n10833), .A2(n11033), .ZN(n4801) );
  NOR2_X1 U6270 ( .A1(n11047), .A2(n11261), .ZN(n6515) );
  AND2_X1 U6272 ( .A1(n11185), .A2(n11186), .ZN(n3907) );
  OR2_X1 U6273 ( .A1(n10431), .A2(n5279), .ZN(n10577) );
  AND2_X1 U6274 ( .A1(n10620), .A2(n11226), .ZN(n10623) );
  NOR2_X1 U6275 ( .A1(n11990), .A2(n10863), .ZN(n11617) );
  INV_X1 U6276 ( .A(n12566), .ZN(n13557) );
  AOI21_X1 U6277 ( .B1(n12512), .B2(n10863), .A(n6374), .ZN(n5090) );
  NOR2_X1 U6278 ( .A1(n12211), .A2(n12111), .ZN(n4449) );
  INV_X1 U6279 ( .A(n10648), .ZN(n12343) );
  INV_X1 U6280 ( .A(n12200), .ZN(n11807) );
  AND2_X1 U6281 ( .A1(n11007), .A2(n11006), .ZN(n3013) );
  INV_X1 U6282 ( .A(n11990), .ZN(n5637) );
  INV_X1 U6283 ( .A(n3653), .ZN(n3108) );
  OR2_X1 U6284 ( .A1(n10923), .A2(n10920), .ZN(n3776) );
  AND2_X1 U6285 ( .A1(n11195), .A2(n11194), .ZN(n12261) );
  INV_X1 U6286 ( .A(n4341), .ZN(n11954) );
  INV_X1 U6288 ( .A(n10905), .ZN(n11927) );
  INV_X1 U6289 ( .A(n11921), .ZN(n11549) );
  NOR2_X1 U6291 ( .A1(n11022), .A2(n11315), .ZN(n3882) );
  AND2_X1 U6292 ( .A1(n3817), .A2(n11248), .ZN(n3275) );
  OR2_X1 U6293 ( .A1(n11540), .A2(n572), .ZN(n6659) );
  INV_X1 U6294 ( .A(n4474), .ZN(n12808) );
  OR2_X1 U6295 ( .A1(n10685), .A2(n28405), .ZN(n6780) );
  OR2_X1 U6296 ( .A1(n10691), .A2(n4538), .ZN(n4537) );
  AND2_X1 U6297 ( .A1(n10957), .A2(n10962), .ZN(n6775) );
  OR2_X1 U6299 ( .A1(n11116), .A2(n11115), .ZN(n3807) );
  AND2_X1 U6300 ( .A1(n12042), .A2(n11962), .ZN(n12043) );
  OR2_X1 U6301 ( .A1(n11963), .A2(n11968), .ZN(n2976) );
  OR2_X1 U6302 ( .A1(n11514), .A2(n12244), .ZN(n3021) );
  AOI21_X1 U6303 ( .B1(n12155), .B2(n12991), .A(n430), .ZN(n11387) );
  OR2_X1 U6304 ( .A1(n5964), .A2(n2008), .ZN(n4997) );
  INV_X1 U6305 ( .A(n13457), .ZN(n6298) );
  XNOR2_X1 U6306 ( .A(n13460), .B(n13459), .ZN(n2172) );
  OR2_X1 U6307 ( .A1(n14593), .A2(n14101), .ZN(n4150) );
  AND2_X1 U6308 ( .A1(n2440), .A2(n11946), .ZN(n11950) );
  AND2_X1 U6310 ( .A1(n15503), .A2(n15506), .ZN(n5575) );
  NOR2_X1 U6311 ( .A1(n12146), .A2(n11715), .ZN(n5169) );
  OR2_X1 U6312 ( .A1(n11415), .A2(n11715), .ZN(n3688) );
  INV_X1 U6314 ( .A(n12377), .ZN(n13562) );
  XNOR2_X1 U6315 ( .A(n2975), .B(n13209), .ZN(n13402) );
  INV_X1 U6316 ( .A(n13025), .ZN(n2975) );
  OR3_X1 U6317 ( .A1(n15180), .A2(n28803), .A3(n15174), .ZN(n13841) );
  OR2_X1 U6318 ( .A1(n14407), .A2(n5584), .ZN(n4974) );
  AND2_X1 U6319 ( .A1(n14398), .A2(n13877), .ZN(n4009) );
  INV_X1 U6320 ( .A(n28806), .ZN(n2959) );
  INV_X1 U6321 ( .A(n14166), .ZN(n13947) );
  AND2_X1 U6322 ( .A1(n14241), .A2(n15194), .ZN(n6571) );
  AND2_X1 U6323 ( .A1(n14078), .A2(n14250), .ZN(n5789) );
  AND2_X1 U6324 ( .A1(n14165), .A2(n14487), .ZN(n13948) );
  OAI211_X1 U6325 ( .C1(n5693), .C2(n14181), .A(n5451), .B(n1320), .ZN(n15345)
         );
  INV_X1 U6326 ( .A(n14480), .ZN(n14161) );
  OR2_X1 U6328 ( .A1(n14084), .A2(n14287), .ZN(n14080) );
  NAND2_X1 U6329 ( .A1(n1848), .A2(n15171), .ZN(n13865) );
  OR2_X1 U6330 ( .A1(n14262), .A2(n14259), .ZN(n13761) );
  OR2_X1 U6331 ( .A1(n15491), .A2(n15485), .ZN(n14618) );
  OAI211_X1 U6332 ( .C1(n14575), .C2(n2733), .A(n2732), .B(n2731), .ZN(n16304)
         );
  OAI21_X1 U6333 ( .B1(n14172), .B2(n14173), .A(n15199), .ZN(n3012) );
  INV_X1 U6334 ( .A(n16283), .ZN(n16486) );
  INV_X1 U6335 ( .A(n14645), .ZN(n2191) );
  OR2_X1 U6336 ( .A1(n13847), .A2(n293), .ZN(n6725) );
  NOR2_X1 U6337 ( .A1(n4992), .A2(n15060), .ZN(n15062) );
  AOI21_X1 U6339 ( .B1(n14496), .B2(n14154), .A(n6798), .ZN(n14501) );
  AND2_X1 U6340 ( .A1(n14495), .A2(n14494), .ZN(n6798) );
  OR2_X1 U6341 ( .A1(n14453), .A2(n1320), .ZN(n5641) );
  OR2_X1 U6342 ( .A1(n15164), .A2(n15464), .ZN(n4677) );
  OR2_X1 U6343 ( .A1(n15010), .A2(n15374), .ZN(n6877) );
  OAI211_X1 U6344 ( .C1(n15008), .C2(n426), .A(n15369), .B(n3783), .ZN(n6880)
         );
  AOI22_X1 U6345 ( .A1(n2608), .A2(n14230), .B1(n14108), .B2(n14107), .ZN(
        n14109) );
  OAI22_X1 U6346 ( .A1(n14390), .A2(n14601), .B1(n15288), .B2(n14391), .ZN(
        n2208) );
  OR2_X1 U6347 ( .A1(n15691), .A2(n13989), .ZN(n4407) );
  AND2_X1 U6348 ( .A1(n13932), .A2(n2493), .ZN(n13930) );
  AND2_X1 U6349 ( .A1(n14784), .A2(n15184), .ZN(n14533) );
  AND2_X1 U6350 ( .A1(n14677), .A2(n15098), .ZN(n4660) );
  AND2_X1 U6351 ( .A1(n15183), .A2(n15182), .ZN(n13818) );
  AND2_X1 U6353 ( .A1(n15015), .A2(n15014), .ZN(n15320) );
  OR2_X1 U6354 ( .A1(n14516), .A2(n15115), .ZN(n5444) );
  INV_X1 U6355 ( .A(n14928), .ZN(n14960) );
  INV_X1 U6356 ( .A(n14697), .ZN(n15512) );
  INV_X1 U6357 ( .A(n13587), .ZN(n14038) );
  OAI21_X1 U6358 ( .B1(n15335), .B2(n15338), .A(n28802), .ZN(n15240) );
  OR2_X1 U6359 ( .A1(n15104), .A2(n15420), .ZN(n5379) );
  XNOR2_X1 U6360 ( .A(n15397), .B(n1957), .ZN(n17296) );
  OR2_X1 U6361 ( .A1(n14187), .A2(n12743), .ZN(n14189) );
  OR2_X1 U6362 ( .A1(n14261), .A2(n3395), .ZN(n3750) );
  OR2_X1 U6363 ( .A1(n14098), .A2(n3396), .ZN(n3749) );
  OAI21_X1 U6364 ( .B1(n13758), .B2(n15152), .A(n2448), .ZN(n16318) );
  OAI21_X1 U6365 ( .B1(n28222), .B2(n2028), .A(n15056), .ZN(n2162) );
  AND3_X1 U6366 ( .A1(n15264), .A2(n4097), .A3(n2738), .ZN(n14711) );
  OR2_X1 U6367 ( .A1(n15260), .A2(n15054), .ZN(n2738) );
  XNOR2_X1 U6368 ( .A(n6454), .B(n16625), .ZN(n6453) );
  AND2_X1 U6369 ( .A1(n14021), .A2(n14024), .ZN(n3782) );
  INV_X1 U6370 ( .A(n16878), .ZN(n17388) );
  XNOR2_X1 U6371 ( .A(n16051), .B(n1967), .ZN(n16525) );
  OR2_X1 U6372 ( .A1(n14706), .A2(n15506), .ZN(n6216) );
  OR2_X1 U6373 ( .A1(n14641), .A2(n15082), .ZN(n2592) );
  AND2_X1 U6374 ( .A1(n2744), .A2(n14982), .ZN(n2743) );
  OR2_X1 U6375 ( .A1(n14797), .A2(n14534), .ZN(n2742) );
  XNOR2_X1 U6376 ( .A(n15545), .B(n6295), .ZN(n15874) );
  INV_X1 U6377 ( .A(n3856), .ZN(n6295) );
  AND2_X1 U6378 ( .A1(n17348), .A2(n29632), .ZN(n16948) );
  XNOR2_X1 U6379 ( .A(n28406), .B(n4852), .ZN(n16203) );
  AND2_X1 U6380 ( .A1(n16724), .A2(n4687), .ZN(n6559) );
  XNOR2_X1 U6381 ( .A(n15909), .B(n5406), .ZN(n15682) );
  INV_X1 U6382 ( .A(n16377), .ZN(n5406) );
  XNOR2_X1 U6383 ( .A(n15660), .B(n15659), .ZN(n16944) );
  INV_X1 U6384 ( .A(n15174), .ZN(n3080) );
  OR2_X1 U6385 ( .A1(n15326), .A2(n15014), .ZN(n2699) );
  INV_X1 U6386 ( .A(n3565), .ZN(n4978) );
  INV_X1 U6388 ( .A(n16467), .ZN(n6296) );
  NOR2_X1 U6389 ( .A1(n4218), .A2(n17548), .ZN(n16946) );
  INV_X1 U6390 ( .A(n17338), .ZN(n17201) );
  OR2_X1 U6392 ( .A1(n17459), .A2(n16812), .ZN(n16813) );
  AND2_X1 U6396 ( .A1(n16860), .A2(n16814), .ZN(n16687) );
  INV_X1 U6397 ( .A(n17137), .ZN(n17502) );
  OR2_X1 U6398 ( .A1(n17304), .A2(n6002), .ZN(n6001) );
  AND2_X1 U6399 ( .A1(n17304), .A2(n17421), .ZN(n17616) );
  OR2_X1 U6400 ( .A1(n4269), .A2(n17830), .ZN(n2856) );
  INV_X1 U6401 ( .A(n4218), .ZN(n2133) );
  NOR2_X1 U6402 ( .A1(n5398), .A2(n17552), .ZN(n2632) );
  AND2_X1 U6404 ( .A1(n18197), .A2(n16718), .ZN(n4174) );
  AOI21_X1 U6405 ( .B1(n511), .B2(n18500), .A(n18506), .ZN(n5392) );
  AND2_X1 U6407 ( .A1(n18325), .A2(n18262), .ZN(n4058) );
  OR2_X1 U6408 ( .A1(n337), .A2(n17437), .ZN(n17308) );
  AND3_X1 U6409 ( .A1(n18441), .A2(n4929), .A3(n18444), .ZN(n4786) );
  OR2_X1 U6410 ( .A1(n18012), .A2(n18480), .ZN(n5179) );
  INV_X1 U6412 ( .A(n17336), .ZN(n2664) );
  INV_X1 U6413 ( .A(n387), .ZN(n6830) );
  OR2_X1 U6414 ( .A1(n17441), .A2(n336), .ZN(n5458) );
  NAND2_X1 U6415 ( .A1(n3250), .A2(n17422), .ZN(n18231) );
  AND2_X1 U6416 ( .A1(n17695), .A2(n18276), .ZN(n17804) );
  AND2_X1 U6417 ( .A1(n18124), .A2(n17834), .ZN(n17840) );
  AND2_X1 U6418 ( .A1(n18596), .A2(n18595), .ZN(n2341) );
  INV_X1 U6419 ( .A(n18332), .ZN(n18372) );
  AND2_X1 U6420 ( .A1(n18232), .A2(n18402), .ZN(n3285) );
  OAI21_X1 U6421 ( .B1(n17715), .B2(n17720), .A(n6588), .ZN(n18526) );
  OR2_X1 U6422 ( .A1(n17990), .A2(n6927), .ZN(n6713) );
  OR2_X1 U6423 ( .A1(n15647), .A2(n28793), .ZN(n5610) );
  OR2_X1 U6424 ( .A1(n16714), .A2(n4283), .ZN(n5609) );
  OR2_X1 U6425 ( .A1(n518), .A2(n18356), .ZN(n2317) );
  OR2_X1 U6426 ( .A1(n6030), .A2(n16611), .ZN(n2838) );
  OR2_X1 U6427 ( .A1(n4059), .A2(n18268), .ZN(n4119) );
  AND2_X1 U6429 ( .A1(n6230), .A2(n6229), .ZN(n6228) );
  AND2_X1 U6430 ( .A1(n18285), .A2(n18081), .ZN(n18083) );
  INV_X1 U6431 ( .A(n19706), .ZN(n3284) );
  AOI22_X1 U6432 ( .A1(n16980), .A2(n18523), .B1(n18524), .B2(n373), .ZN(
        n16981) );
  INV_X1 U6433 ( .A(n19111), .ZN(n18980) );
  INV_X1 U6435 ( .A(n5492), .ZN(n5491) );
  AND2_X1 U6436 ( .A1(n20193), .A2(n20414), .ZN(n20578) );
  OR2_X1 U6437 ( .A1(n17918), .A2(n18354), .ZN(n5842) );
  INV_X1 U6438 ( .A(n20200), .ZN(n20304) );
  XNOR2_X1 U6439 ( .A(n18857), .B(n18856), .ZN(n19269) );
  INV_X1 U6440 ( .A(n18877), .ZN(n3403) );
  OR2_X1 U6441 ( .A1(n17639), .A2(n29125), .ZN(n17640) );
  OR2_X1 U6445 ( .A1(n18458), .A2(n18459), .ZN(n6670) );
  AND2_X1 U6446 ( .A1(n18455), .A2(n18456), .ZN(n6671) );
  INV_X1 U6447 ( .A(n20302), .ZN(n5436) );
  INV_X1 U6448 ( .A(n18690), .ZN(n18927) );
  XNOR2_X1 U6449 ( .A(n19139), .B(n1179), .ZN(n5746) );
  XNOR2_X1 U6450 ( .A(n18867), .B(n19108), .ZN(n19599) );
  XNOR2_X1 U6451 ( .A(n19247), .B(n4030), .ZN(n19248) );
  OR2_X1 U6452 ( .A1(n18042), .A2(n18423), .ZN(n4802) );
  OAI21_X1 U6453 ( .B1(n18202), .B2(n18201), .A(n18200), .ZN(n6488) );
  XNOR2_X1 U6454 ( .A(n19252), .B(n18948), .ZN(n6276) );
  AND2_X1 U6455 ( .A1(n20533), .A2(n20933), .ZN(n5125) );
  OR2_X1 U6456 ( .A1(n20144), .A2(n21091), .ZN(n5854) );
  INV_X1 U6457 ( .A(n21087), .ZN(n21426) );
  AND2_X1 U6458 ( .A1(n20283), .A2(n20282), .ZN(n19896) );
  NOR2_X1 U6459 ( .A1(n20443), .A2(n20299), .ZN(n20446) );
  OR2_X1 U6460 ( .A1(n22145), .A2(n22139), .ZN(n21030) );
  NOR2_X1 U6461 ( .A1(n20406), .A2(n28501), .ZN(n6315) );
  XNOR2_X1 U6462 ( .A(n5522), .B(n5521), .ZN(n5520) );
  AND2_X1 U6464 ( .A1(n20474), .A2(n5408), .ZN(n21275) );
  OR2_X1 U6465 ( .A1(n20477), .A2(n20475), .ZN(n20352) );
  OR2_X1 U6466 ( .A1(n21143), .A2(n4395), .ZN(n4394) );
  AND2_X1 U6467 ( .A1(n20351), .A2(n21547), .ZN(n20362) );
  OAI21_X1 U6468 ( .B1(n18846), .B2(n18776), .A(n19765), .ZN(n5469) );
  OR2_X1 U6470 ( .A1(n20450), .A2(n5375), .ZN(n2747) );
  OR2_X1 U6471 ( .A1(n20183), .A2(n499), .ZN(n19185) );
  OR2_X1 U6472 ( .A1(n20721), .A2(n21599), .ZN(n5720) );
  INV_X1 U6473 ( .A(n22320), .ZN(n22379) );
  OR2_X1 U6474 ( .A1(n20466), .A2(n21932), .ZN(n20184) );
  AND2_X1 U6475 ( .A1(n21119), .A2(n21144), .ZN(n21122) );
  NAND3_X1 U6476 ( .A1(n21412), .A2(n4937), .A3(n28184), .ZN(n2653) );
  INV_X1 U6478 ( .A(n5684), .ZN(n5983) );
  OAI21_X1 U6479 ( .B1(n21447), .B2(n21080), .A(n20213), .ZN(n21959) );
  NOR2_X1 U6480 ( .A1(n21674), .A2(n21679), .ZN(n21080) );
  INV_X1 U6481 ( .A(n22633), .ZN(n22691) );
  OR2_X1 U6482 ( .A1(n21625), .A2(n22145), .ZN(n21028) );
  OR2_X1 U6483 ( .A1(n22149), .A2(n22148), .ZN(n2097) );
  AND2_X1 U6485 ( .A1(n20276), .A2(n6016), .ZN(n2666) );
  AND2_X1 U6486 ( .A1(n20269), .A2(n2669), .ZN(n2668) );
  OR2_X1 U6487 ( .A1(n21645), .A2(n21642), .ZN(n4071) );
  OR2_X1 U6488 ( .A1(n22288), .A2(n21208), .ZN(n3858) );
  AOI21_X1 U6489 ( .B1(n6240), .B2(n20781), .A(n20780), .ZN(n20885) );
  INV_X1 U6490 ( .A(n5782), .ZN(n5780) );
  OR2_X1 U6491 ( .A1(n20441), .A2(n20440), .ZN(n3547) );
  XNOR2_X1 U6492 ( .A(n22822), .B(n22132), .ZN(n22571) );
  XNOR2_X1 U6493 ( .A(n22132), .B(n21959), .ZN(n22800) );
  INV_X1 U6494 ( .A(n20885), .ZN(n22787) );
  XNOR2_X1 U6495 ( .A(n5395), .B(n22903), .ZN(n6364) );
  XNOR2_X1 U6496 ( .A(n22337), .B(n634), .ZN(n5395) );
  OR2_X1 U6497 ( .A1(n20888), .A2(n20889), .ZN(n6039) );
  AND2_X1 U6498 ( .A1(n21237), .A2(n21399), .ZN(n21751) );
  XNOR2_X1 U6499 ( .A(n6141), .B(n22791), .ZN(n22164) );
  NAND2_X1 U6500 ( .A1(n4638), .A2(n4634), .ZN(n22594) );
  OR2_X1 U6502 ( .A1(n21382), .A2(n4266), .ZN(n4265) );
  OR2_X1 U6503 ( .A1(n29488), .A2(n21269), .ZN(n6427) );
  INV_X1 U6504 ( .A(n20989), .ZN(n6116) );
  XNOR2_X1 U6505 ( .A(n21903), .B(n22488), .ZN(n22727) );
  OR2_X1 U6506 ( .A1(n21257), .A2(n5772), .ZN(n3319) );
  XNOR2_X1 U6507 ( .A(n22417), .B(n22416), .ZN(n23651) );
  OR2_X1 U6508 ( .A1(n23733), .A2(n2141), .ZN(n2951) );
  OR2_X1 U6510 ( .A1(n23790), .A2(n23492), .ZN(n23319) );
  OR2_X1 U6511 ( .A1(n21445), .A2(n20833), .ZN(n6349) );
  XNOR2_X1 U6512 ( .A(n20682), .B(n20681), .ZN(n3887) );
  NOR2_X1 U6513 ( .A1(n2138), .A2(n1838), .ZN(n4255) );
  NOR2_X1 U6514 ( .A1(n28390), .A2(n29074), .ZN(n4256) );
  INV_X1 U6515 ( .A(n23177), .ZN(n23645) );
  OR2_X1 U6517 ( .A1(n23501), .A2(n28554), .ZN(n5354) );
  INV_X1 U6518 ( .A(n4726), .ZN(n23537) );
  OR2_X1 U6519 ( .A1(n23800), .A2(n28444), .ZN(n23536) );
  AND2_X1 U6520 ( .A1(n22284), .A2(n29061), .ZN(n23554) );
  AOI22_X1 U6521 ( .A1(n5541), .A2(n23835), .B1(n23833), .B2(n23834), .ZN(
        n4532) );
  AND2_X1 U6522 ( .A1(n23662), .A2(n23163), .ZN(n23524) );
  INV_X1 U6523 ( .A(n23769), .ZN(n23499) );
  OR2_X1 U6525 ( .A1(n23765), .A2(n23764), .ZN(n23501) );
  OR2_X1 U6527 ( .A1(n23586), .A2(n23262), .ZN(n4234) );
  NOR2_X1 U6528 ( .A1(n23455), .A2(n23456), .ZN(n23357) );
  XNOR2_X1 U6529 ( .A(n22922), .B(n4229), .ZN(n4228) );
  AND2_X1 U6530 ( .A1(n29120), .A2(n28523), .ZN(n6596) );
  NOR2_X1 U6531 ( .A1(n24581), .A2(n24468), .ZN(n3295) );
  OR2_X1 U6532 ( .A1(n23789), .A2(n23790), .ZN(n6609) );
  OR2_X1 U6533 ( .A1(n23809), .A2(n22742), .ZN(n2202) );
  OR2_X1 U6534 ( .A1(n24709), .A2(n24341), .ZN(n24705) );
  INV_X1 U6535 ( .A(n23606), .ZN(n5347) );
  XNOR2_X1 U6537 ( .A(n22137), .B(n22138), .ZN(n23712) );
  OR2_X1 U6538 ( .A1(n23228), .A2(n23227), .ZN(n23229) );
  AND2_X1 U6539 ( .A1(n2823), .A2(n23126), .ZN(n2822) );
  OR2_X1 U6540 ( .A1(n4664), .A2(n24376), .ZN(n3205) );
  INV_X1 U6541 ( .A(n24613), .ZN(n24057) );
  OR2_X1 U6542 ( .A1(n24593), .A2(n24141), .ZN(n3481) );
  INV_X1 U6543 ( .A(n23467), .ZN(n6787) );
  NAND4_X1 U6544 ( .A1(n6109), .A2(n23409), .A3(n23410), .A4(n23507), .ZN(
        n6110) );
  NOR2_X1 U6545 ( .A1(n24614), .A2(n29109), .ZN(n5217) );
  NAND2_X1 U6546 ( .A1(n24339), .A2(n24334), .ZN(n24709) );
  AND2_X1 U6547 ( .A1(n24706), .A2(n24708), .ZN(n5751) );
  OR2_X1 U6548 ( .A1(n23042), .A2(n23632), .ZN(n23043) );
  INV_X1 U6549 ( .A(n2153), .ZN(n2154) );
  INV_X1 U6551 ( .A(n22747), .ZN(n23979) );
  AND2_X1 U6552 ( .A1(n5210), .A2(n25007), .ZN(n24065) );
  AOI22_X1 U6553 ( .A1(n23303), .A2(n5699), .B1(n5530), .B2(n4019), .ZN(n4177)
         );
  INV_X1 U6554 ( .A(n24582), .ZN(n24054) );
  OAI211_X1 U6555 ( .C1(n22998), .C2(n23563), .A(n2623), .B(n2622), .ZN(n24437) );
  INV_X1 U6557 ( .A(n24188), .ZN(n2240) );
  BUF_X1 U6558 ( .A(n24984), .Z(n25781) );
  XNOR2_X1 U6560 ( .A(n24958), .B(n24957), .ZN(n26384) );
  INV_X1 U6562 ( .A(n5263), .ZN(n25750) );
  AND2_X1 U6563 ( .A1(n29622), .A2(n5263), .ZN(n27079) );
  INV_X1 U6564 ( .A(n25815), .ZN(n27086) );
  AND2_X1 U6565 ( .A1(n26614), .A2(n27067), .ZN(n27065) );
  AND2_X1 U6566 ( .A1(n24501), .A2(n24500), .ZN(n3206) );
  XNOR2_X1 U6567 ( .A(n26118), .B(n25849), .ZN(n25311) );
  INV_X1 U6569 ( .A(n27038), .ZN(n5314) );
  BUF_X1 U6570 ( .A(n25633), .Z(n26960) );
  NOR2_X1 U6571 ( .A1(n23862), .A2(n25418), .ZN(n23863) );
  NAND2_X1 U6572 ( .A1(n24575), .A2(n26560), .ZN(n5504) );
  NOR2_X1 U6573 ( .A1(n377), .A2(n4913), .ZN(n24575) );
  NOR2_X1 U6574 ( .A1(n26435), .A2(n26935), .ZN(n26558) );
  OR2_X1 U6575 ( .A1(n28471), .A2(n28423), .ZN(n2323) );
  OR2_X1 U6576 ( .A1(n26801), .A2(n26800), .ZN(n6322) );
  AND2_X1 U6577 ( .A1(n26132), .A2(n28642), .ZN(n26260) );
  INV_X1 U6581 ( .A(n2145), .ZN(n27123) );
  INV_X1 U6582 ( .A(n26851), .ZN(n27838) );
  INV_X1 U6583 ( .A(n26310), .ZN(n26866) );
  NOR2_X1 U6584 ( .A1(n26125), .A2(n27140), .ZN(n26519) );
  INV_X1 U6585 ( .A(n26507), .ZN(n27087) );
  OR2_X1 U6586 ( .A1(n26251), .A2(n26733), .ZN(n5390) );
  OR2_X1 U6587 ( .A1(n5388), .A2(n26995), .ZN(n5391) );
  OR2_X1 U6588 ( .A1(n27043), .A2(n29058), .ZN(n4497) );
  AND2_X1 U6589 ( .A1(n27052), .A2(n25983), .ZN(n27017) );
  XNOR2_X1 U6591 ( .A(n2153), .B(n1928), .ZN(n25257) );
  OR2_X1 U6592 ( .A1(n26222), .A2(n29159), .ZN(n28101) );
  INV_X1 U6593 ( .A(n26652), .ZN(n27537) );
  INV_X1 U6594 ( .A(n27038), .ZN(n27209) );
  NOR2_X1 U6595 ( .A1(n26197), .A2(n26196), .ZN(n5373) );
  AND2_X1 U6597 ( .A1(n342), .A2(n26960), .ZN(n4921) );
  AND2_X1 U6598 ( .A1(n27465), .A2(n29468), .ZN(n6712) );
  INV_X1 U6599 ( .A(n27525), .ZN(n4809) );
  NOR3_X1 U6600 ( .A1(n27505), .A2(n27527), .A3(n27523), .ZN(n27513) );
  OR2_X1 U6601 ( .A1(n26804), .A2(n26280), .ZN(n3075) );
  OR2_X1 U6602 ( .A1(n26785), .A2(n6070), .ZN(n3703) );
  NOR2_X1 U6603 ( .A1(n26787), .A2(n26788), .ZN(n3702) );
  AND2_X1 U6605 ( .A1(n26880), .A2(n27301), .ZN(n27259) );
  OAI21_X1 U6606 ( .B1(n26918), .B2(n26782), .A(n26920), .ZN(n6633) );
  NOR2_X1 U6607 ( .A1(n27547), .A2(n27203), .ZN(n27546) );
  AND2_X1 U6608 ( .A1(n27567), .A2(n3087), .ZN(n2268) );
  AOI21_X1 U6609 ( .B1(n28421), .B2(n6724), .A(n26935), .ZN(n6723) );
  NOR2_X1 U6610 ( .A1(n27591), .A2(n27596), .ZN(n27592) );
  INV_X1 U6612 ( .A(n27672), .ZN(n5877) );
  NOR2_X1 U6614 ( .A1(n27780), .A2(n29070), .ZN(n27769) );
  NAND2_X1 U6616 ( .A1(n6025), .A2(n6024), .ZN(n27772) );
  OR2_X1 U6617 ( .A1(n6008), .A2(n26297), .ZN(n6024) );
  INV_X1 U6618 ( .A(n27826), .ZN(n2378) );
  AND2_X1 U6619 ( .A1(n27827), .A2(n27841), .ZN(n2767) );
  OAI211_X1 U6620 ( .C1(n27056), .C2(n27902), .A(n5301), .B(n26849), .ZN(n5300) );
  AND3_X1 U6621 ( .A1(n26624), .A2(n28446), .A3(n26246), .ZN(n26626) );
  OAI22_X1 U6622 ( .A1(n4411), .A2(n27041), .B1(n28783), .B2(n28130), .ZN(
        n25555) );
  AOI21_X1 U6623 ( .B1(n25506), .B2(n25505), .A(n25504), .ZN(n6857) );
  OR2_X1 U6624 ( .A1(n7828), .A2(n7635), .ZN(n8203) );
  INV_X1 U6625 ( .A(n8207), .ZN(n3447) );
  INV_X1 U6626 ( .A(n7318), .ZN(n6384) );
  OR2_X1 U6627 ( .A1(n7349), .A2(n8158), .ZN(n2944) );
  AND2_X1 U6628 ( .A1(n7288), .A2(n4856), .ZN(n2624) );
  AND2_X1 U6629 ( .A1(n7499), .A2(n7500), .ZN(n8589) );
  AND2_X1 U6630 ( .A1(n7986), .A2(n631), .ZN(n7662) );
  NAND2_X1 U6632 ( .A1(n5160), .A2(n9045), .ZN(n5159) );
  OR2_X1 U6633 ( .A1(n9041), .A2(n9243), .ZN(n9244) );
  INV_X1 U6634 ( .A(n8941), .ZN(n9566) );
  OR2_X1 U6635 ( .A1(n8141), .A2(n7336), .ZN(n7723) );
  INV_X1 U6636 ( .A(n8465), .ZN(n8463) );
  INV_X1 U6637 ( .A(n7279), .ZN(n2115) );
  INV_X1 U6638 ( .A(n7320), .ZN(n5242) );
  INV_X1 U6639 ( .A(n8610), .ZN(n8609) );
  INV_X1 U6640 ( .A(n8762), .ZN(n9561) );
  OR2_X1 U6641 ( .A1(n7550), .A2(n7330), .ZN(n7789) );
  AND2_X1 U6642 ( .A1(n7330), .A2(n7782), .ZN(n2670) );
  INV_X1 U6645 ( .A(n7914), .ZN(n3329) );
  NOR2_X1 U6647 ( .A1(n6908), .A2(n29304), .ZN(n6316) );
  AND2_X1 U6649 ( .A1(n7585), .A2(n7303), .ZN(n5558) );
  INV_X1 U6650 ( .A(n7664), .ZN(n2099) );
  OR2_X1 U6651 ( .A1(n7485), .A2(n7665), .ZN(n7486) );
  OR2_X1 U6652 ( .A1(n8873), .A2(n8877), .ZN(n8532) );
  OR2_X1 U6653 ( .A1(n7313), .A2(n7898), .ZN(n6545) );
  AOI22_X1 U6654 ( .A1(n8245), .A2(n8246), .B1(n8243), .B2(n8244), .ZN(n5911)
         );
  OR2_X1 U6655 ( .A1(n7924), .A2(n7626), .ZN(n8218) );
  OR2_X1 U6656 ( .A1(n7520), .A2(n29321), .ZN(n5072) );
  INV_X1 U6657 ( .A(n8035), .ZN(n7510) );
  OR2_X1 U6658 ( .A1(n7376), .A2(n7692), .ZN(n8242) );
  OR2_X1 U6659 ( .A1(n8560), .A2(n8562), .ZN(n8568) );
  AND2_X1 U6660 ( .A1(n8490), .A2(n9095), .ZN(n2977) );
  AND2_X1 U6661 ( .A1(n8955), .A2(n8801), .ZN(n8472) );
  OR2_X1 U6662 ( .A1(n6908), .A2(n284), .ZN(n2980) );
  INV_X1 U6663 ( .A(n9531), .ZN(n6892) );
  AND2_X1 U6664 ( .A1(n7258), .A2(n29629), .ZN(n2170) );
  AND2_X1 U6665 ( .A1(n8685), .A2(n8687), .ZN(n4729) );
  INV_X1 U6667 ( .A(n8872), .ZN(n9061) );
  AND2_X1 U6668 ( .A1(n7216), .A2(n3301), .ZN(n3300) );
  OR2_X1 U6669 ( .A1(n8685), .A2(n8687), .ZN(n9026) );
  INV_X1 U6670 ( .A(n8717), .ZN(n4321) );
  OR2_X1 U6671 ( .A1(n7594), .A2(n7870), .ZN(n6801) );
  OR2_X1 U6672 ( .A1(n7604), .A2(n7864), .ZN(n3034) );
  OR2_X1 U6674 ( .A1(n9227), .A2(n597), .ZN(n8102) );
  OAI22_X1 U6675 ( .A1(n8234), .A2(n7619), .B1(n6973), .B2(n7919), .ZN(n6976)
         );
  INV_X1 U6677 ( .A(n7114), .ZN(n8829) );
  OR2_X1 U6678 ( .A1(n8827), .A2(n8192), .ZN(n8464) );
  INV_X1 U6679 ( .A(n8327), .ZN(n5594) );
  AND3_X1 U6680 ( .A1(n8498), .A2(n8497), .A3(n8651), .ZN(n3128) );
  INV_X1 U6681 ( .A(n9029), .ZN(n9027) );
  INV_X1 U6682 ( .A(n9034), .ZN(n7714) );
  OR2_X1 U6685 ( .A1(n7748), .A2(n7749), .ZN(n2358) );
  OAI21_X1 U6686 ( .B1(n8873), .B2(n8403), .A(n8404), .ZN(n3297) );
  OR2_X1 U6687 ( .A1(n7736), .A2(n7268), .ZN(n3115) );
  AND2_X1 U6688 ( .A1(n7792), .A2(n28149), .ZN(n2546) );
  OR3_X1 U6690 ( .A1(n8958), .A2(n8802), .A3(n8955), .ZN(n8316) );
  OR2_X1 U6691 ( .A1(n8154), .A2(n7550), .ZN(n3282) );
  INV_X1 U6692 ( .A(n8886), .ZN(n8334) );
  INV_X1 U6693 ( .A(n8605), .ZN(n2320) );
  OR2_X1 U6694 ( .A1(n8914), .A2(n8669), .ZN(n8512) );
  BUF_X1 U6695 ( .A(n8499), .Z(n8652) );
  INV_X1 U6696 ( .A(n8499), .ZN(n8656) );
  AOI21_X1 U6697 ( .B1(n7383), .B2(n617), .A(n3639), .ZN(n6748) );
  INV_X1 U6698 ( .A(n6718), .ZN(n8753) );
  INV_X1 U6699 ( .A(n8320), .ZN(n9533) );
  OAI211_X1 U6700 ( .C1(n7989), .C2(n7990), .A(n7988), .B(n7987), .ZN(n8664)
         );
  OR2_X1 U6701 ( .A1(n8211), .A2(n439), .ZN(n3117) );
  OR2_X1 U6702 ( .A1(n8811), .A2(n2238), .ZN(n8679) );
  OR2_X1 U6703 ( .A1(n8292), .A2(n8287), .ZN(n2568) );
  AND2_X1 U6705 ( .A1(n9196), .A2(n329), .ZN(n9199) );
  INV_X1 U6706 ( .A(n8726), .ZN(n8603) );
  INV_X1 U6707 ( .A(n8984), .ZN(n8982) );
  OR2_X1 U6708 ( .A1(n8157), .A2(n8156), .ZN(n6874) );
  INV_X1 U6709 ( .A(n8966), .ZN(n8837) );
  OAI21_X1 U6710 ( .B1(n3225), .B2(n29241), .A(n3224), .ZN(n8255) );
  AOI22_X1 U6711 ( .A1(n9168), .A2(n9167), .B1(n9165), .B2(n9166), .ZN(n9312)
         );
  NOR2_X1 U6712 ( .A1(n28638), .A2(n11197), .ZN(n5916) );
  INV_X1 U6713 ( .A(n9684), .ZN(n10146) );
  OR2_X1 U6714 ( .A1(n10497), .A2(n10502), .ZN(n11133) );
  XNOR2_X1 U6715 ( .A(n301), .B(n9991), .ZN(n5410) );
  AND2_X1 U6716 ( .A1(n8734), .A2(n8733), .ZN(n2983) );
  AND2_X1 U6717 ( .A1(n9221), .A2(n9220), .ZN(n2352) );
  OR2_X1 U6719 ( .A1(n8855), .A2(n9070), .ZN(n8862) );
  OAI211_X1 U6720 ( .C1(n9012), .C2(n8910), .A(n9015), .B(n6147), .ZN(n8085)
         );
  INV_X1 U6721 ( .A(n11163), .ZN(n3904) );
  XNOR2_X1 U6723 ( .A(n9312), .B(n9991), .ZN(n10373) );
  OR2_X1 U6724 ( .A1(n10740), .A2(n582), .ZN(n6703) );
  AND2_X1 U6725 ( .A1(n28876), .A2(n11149), .ZN(n10512) );
  OR2_X1 U6726 ( .A1(n10806), .A2(n28627), .ZN(n6360) );
  INV_X1 U6727 ( .A(n11778), .ZN(n11553) );
  AND2_X1 U6728 ( .A1(n10966), .A2(n10965), .ZN(n4715) );
  OR2_X1 U6729 ( .A1(n10872), .A2(n435), .ZN(n2283) );
  OR2_X1 U6730 ( .A1(n4908), .A2(n11094), .ZN(n2464) );
  OAI21_X1 U6731 ( .B1(n10505), .B2(n4383), .A(n11121), .ZN(n9914) );
  OR2_X1 U6732 ( .A1(n10504), .A2(n10507), .ZN(n3460) );
  INV_X1 U6733 ( .A(n29149), .ZN(n3816) );
  INV_X1 U6734 ( .A(n12158), .ZN(n12157) );
  AND2_X1 U6735 ( .A1(n10713), .A2(n1834), .ZN(n4553) );
  OR2_X1 U6736 ( .A1(n4844), .A2(n11599), .ZN(n4843) );
  OR2_X1 U6739 ( .A1(n12058), .A2(n11795), .ZN(n12060) );
  AND2_X1 U6740 ( .A1(n28174), .A2(n29122), .ZN(n6386) );
  AND2_X1 U6741 ( .A1(n12236), .A2(n375), .ZN(n5008) );
  INV_X1 U6742 ( .A(n11491), .ZN(n12302) );
  OR2_X1 U6743 ( .A1(n10713), .A2(n5672), .ZN(n11131) );
  AND2_X1 U6744 ( .A1(n11114), .A2(n11113), .ZN(n5109) );
  OR2_X1 U6745 ( .A1(n12109), .A2(n12110), .ZN(n6282) );
  OR2_X1 U6746 ( .A1(n10819), .A2(n10820), .ZN(n3536) );
  OR2_X1 U6747 ( .A1(n11152), .A2(n5150), .ZN(n10802) );
  XNOR2_X1 U6748 ( .A(n10086), .B(n10089), .ZN(n6183) );
  XNOR2_X1 U6749 ( .A(n10085), .B(n10090), .ZN(n6184) );
  INV_X1 U6750 ( .A(n29078), .ZN(n9348) );
  AND2_X1 U6751 ( .A1(n4296), .A2(n2690), .ZN(n2688) );
  INV_X1 U6752 ( .A(n11332), .ZN(n4463) );
  INV_X1 U6753 ( .A(n11956), .ZN(n5603) );
  OR2_X1 U6754 ( .A1(n10972), .A2(n10970), .ZN(n6368) );
  OR2_X1 U6755 ( .A1(n11551), .A2(n11778), .ZN(n5170) );
  INV_X1 U6756 ( .A(n11206), .ZN(n5258) );
  AND2_X1 U6757 ( .A1(n11754), .A2(n11536), .ZN(n11756) );
  AND2_X1 U6758 ( .A1(n10603), .A2(n10966), .ZN(n3322) );
  INV_X1 U6759 ( .A(n12156), .ZN(n12159) );
  INV_X1 U6760 ( .A(n12507), .ZN(n6374) );
  AND2_X1 U6761 ( .A1(n11955), .A2(n12257), .ZN(n4018) );
  OAI21_X1 U6762 ( .B1(n10637), .B2(n5281), .A(n11093), .ZN(n5280) );
  NOR2_X1 U6763 ( .A1(n10431), .A2(n11207), .ZN(n5281) );
  INV_X1 U6764 ( .A(n11640), .ZN(n11401) );
  AND2_X1 U6765 ( .A1(n12151), .A2(n12150), .ZN(n3603) );
  AND2_X1 U6767 ( .A1(n5533), .A2(n11193), .ZN(n4903) );
  INV_X1 U6768 ( .A(n11458), .ZN(n11874) );
  INV_X1 U6769 ( .A(n11980), .ZN(n11809) );
  AND2_X1 U6770 ( .A1(n6482), .A2(n10717), .ZN(n11489) );
  OR2_X1 U6771 ( .A1(n6411), .A2(n10851), .ZN(n3934) );
  INV_X1 U6772 ( .A(n574), .ZN(n3201) );
  INV_X1 U6774 ( .A(n13444), .ZN(n12600) );
  OR2_X1 U6775 ( .A1(n12156), .A2(n12158), .ZN(n11512) );
  OR2_X1 U6776 ( .A1(n10894), .A2(n11290), .ZN(n6430) );
  OR2_X1 U6777 ( .A1(n12177), .A2(n12181), .ZN(n3604) );
  AND2_X1 U6778 ( .A1(n12516), .A2(n12517), .ZN(n11941) );
  OR2_X1 U6779 ( .A1(n12270), .A2(n28202), .ZN(n12075) );
  OAI21_X1 U6781 ( .B1(n10883), .B2(n11086), .A(n11212), .ZN(n2143) );
  OR2_X1 U6782 ( .A1(n10918), .A2(n2968), .ZN(n10105) );
  INV_X1 U6783 ( .A(n13086), .ZN(n11810) );
  INV_X1 U6784 ( .A(n3871), .ZN(n4297) );
  OR2_X1 U6785 ( .A1(n10113), .A2(n10946), .ZN(n6373) );
  OR2_X1 U6786 ( .A1(n10927), .A2(n10930), .ZN(n2948) );
  OR2_X1 U6787 ( .A1(n11487), .A2(n11787), .ZN(n6480) );
  INV_X1 U6788 ( .A(n12077), .ZN(n5947) );
  AND2_X1 U6789 ( .A1(n12339), .A2(n12338), .ZN(n12028) );
  OR2_X1 U6790 ( .A1(n10648), .A2(n12338), .ZN(n12030) );
  OR2_X1 U6791 ( .A1(n11340), .A2(n11335), .ZN(n11342) );
  OR2_X1 U6792 ( .A1(n11344), .A2(n11345), .ZN(n2580) );
  NOR2_X1 U6793 ( .A1(n4105), .A2(n11505), .ZN(n6132) );
  AND2_X1 U6794 ( .A1(n12303), .A2(n11491), .ZN(n11608) );
  OR2_X1 U6797 ( .A1(n28568), .A2(n333), .ZN(n4101) );
  OR2_X1 U6798 ( .A1(n12155), .A2(n12150), .ZN(n12099) );
  AND3_X1 U6799 ( .A1(n7813), .A2(n28206), .A3(n10808), .ZN(n4389) );
  INV_X1 U6800 ( .A(n12145), .ZN(n11708) );
  AND2_X1 U6801 ( .A1(n11417), .A2(n11648), .ZN(n12142) );
  INV_X1 U6802 ( .A(n11599), .ZN(n12204) );
  OR2_X1 U6803 ( .A1(n10859), .A2(n11181), .ZN(n9055) );
  OR2_X1 U6804 ( .A1(n11043), .A2(n11260), .ZN(n11051) );
  INV_X1 U6805 ( .A(n12284), .ZN(n12279) );
  AND2_X1 U6806 ( .A1(n11859), .A2(n11944), .ZN(n11860) );
  INV_X1 U6807 ( .A(n12332), .ZN(n12018) );
  INV_X1 U6810 ( .A(n12273), .ZN(n4869) );
  OR2_X1 U6811 ( .A1(n12346), .A2(n12338), .ZN(n3592) );
  AND2_X1 U6812 ( .A1(n12206), .A2(n12109), .ZN(n11373) );
  AND2_X1 U6813 ( .A1(n3113), .A2(n11316), .ZN(n9502) );
  OR2_X1 U6814 ( .A1(n10993), .A2(n10992), .ZN(n2165) );
  OAI211_X1 U6815 ( .C1(n10628), .C2(n3441), .A(n2413), .B(n6108), .ZN(n2847)
         );
  INV_X1 U6816 ( .A(n11962), .ZN(n12221) );
  OR2_X1 U6817 ( .A1(n10569), .A2(n10795), .ZN(n3103) );
  OR2_X1 U6818 ( .A1(n6604), .A2(n10572), .ZN(n10574) );
  INV_X1 U6819 ( .A(n12453), .ZN(n13080) );
  XNOR2_X1 U6820 ( .A(n13445), .B(n3374), .ZN(n12262) );
  INV_X1 U6821 ( .A(n2981), .ZN(n4502) );
  INV_X1 U6822 ( .A(n4298), .ZN(n12064) );
  INV_X1 U6823 ( .A(n14600), .ZN(n6048) );
  INV_X1 U6824 ( .A(n13523), .ZN(n12816) );
  AOI21_X1 U6825 ( .B1(n12315), .B2(n5464), .A(n11615), .ZN(n5463) );
  OR2_X1 U6826 ( .A1(n14146), .A2(n3860), .ZN(n3859) );
  INV_X1 U6827 ( .A(n12799), .ZN(n12568) );
  INV_X1 U6828 ( .A(n12632), .ZN(n12603) );
  INV_X1 U6829 ( .A(n13521), .ZN(n13520) );
  INV_X1 U6831 ( .A(n14262), .ZN(n3071) );
  OR2_X1 U6832 ( .A1(n11682), .A2(n12236), .ZN(n10676) );
  OR2_X1 U6833 ( .A1(n5578), .A2(n12232), .ZN(n10674) );
  INV_X1 U6834 ( .A(n12813), .ZN(n13144) );
  AND2_X1 U6835 ( .A1(n5058), .A2(n14376), .ZN(n5057) );
  OR2_X1 U6836 ( .A1(n14434), .A2(n14433), .ZN(n12887) );
  OR2_X1 U6837 ( .A1(n14842), .A2(n15285), .ZN(n5931) );
  OR2_X1 U6838 ( .A1(n14695), .A2(n15285), .ZN(n2893) );
  INV_X1 U6839 ( .A(n14047), .ZN(n6011) );
  OAI211_X1 U6840 ( .C1(n2112), .C2(n28804), .A(n2111), .B(n2110), .ZN(n14621)
         );
  OR2_X1 U6841 ( .A1(n13868), .A2(n28805), .ZN(n3228) );
  OR2_X1 U6842 ( .A1(n14195), .A2(n14193), .ZN(n4500) );
  OR2_X1 U6843 ( .A1(n14451), .A2(n14178), .ZN(n13932) );
  NOR2_X1 U6844 ( .A1(n14294), .A2(n14295), .ZN(n13808) );
  INV_X1 U6845 ( .A(n13306), .ZN(n14291) );
  AND2_X1 U6846 ( .A1(n13893), .A2(n13892), .ZN(n4836) );
  INV_X1 U6847 ( .A(n15388), .ZN(n6517) );
  AND2_X1 U6848 ( .A1(n14142), .A2(n2000), .ZN(n13410) );
  AND2_X1 U6850 ( .A1(n14773), .A2(n14807), .ZN(n14555) );
  AND2_X1 U6851 ( .A1(n15103), .A2(n15420), .ZN(n5381) );
  INV_X1 U6853 ( .A(n13639), .ZN(n13637) );
  INV_X1 U6854 ( .A(n2974), .ZN(n2874) );
  INV_X1 U6857 ( .A(n14373), .ZN(n13726) );
  INV_X1 U6858 ( .A(n14763), .ZN(n4162) );
  OR2_X1 U6859 ( .A1(n15208), .A2(n14928), .ZN(n13785) );
  AOI21_X1 U6860 ( .B1(n28195), .B2(n6854), .A(n28196), .ZN(n6853) );
  INV_X1 U6861 ( .A(n14944), .ZN(n6854) );
  INV_X1 U6862 ( .A(n15046), .ZN(n15226) );
  OR2_X1 U6863 ( .A1(n2974), .A2(n29589), .ZN(n3379) );
  OR2_X1 U6866 ( .A1(n4436), .A2(n28805), .ZN(n4431) );
  AND2_X1 U6867 ( .A1(n29320), .A2(n293), .ZN(n3868) );
  AND3_X1 U6868 ( .A1(n3843), .A2(n13854), .A3(n4840), .ZN(n5598) );
  OR2_X1 U6869 ( .A1(n14839), .A2(n4359), .ZN(n4358) );
  INV_X1 U6870 ( .A(n14969), .ZN(n14793) );
  INV_X1 U6871 ( .A(n5378), .ZN(n14397) );
  INV_X1 U6873 ( .A(n14534), .ZN(n15460) );
  INV_X1 U6874 ( .A(n15503), .ZN(n15497) );
  INV_X1 U6875 ( .A(n14922), .ZN(n15500) );
  INV_X1 U6876 ( .A(n13785), .ZN(n14796) );
  INV_X1 U6877 ( .A(n16388), .ZN(n16471) );
  OAI21_X1 U6878 ( .B1(n2800), .B2(n15209), .A(n15201), .ZN(n2691) );
  AND3_X1 U6880 ( .A1(n14746), .A2(n14747), .A3(n14998), .ZN(n4720) );
  INV_X1 U6881 ( .A(n13796), .ZN(n6640) );
  OR2_X1 U6882 ( .A1(n15238), .A2(n15239), .ZN(n14220) );
  AND2_X1 U6883 ( .A1(n14415), .A2(n6232), .ZN(n6231) );
  INV_X1 U6884 ( .A(n14826), .ZN(n15430) );
  OR2_X1 U6885 ( .A1(n4893), .A2(n14354), .ZN(n14013) );
  OR2_X1 U6886 ( .A1(n13815), .A2(n14408), .ZN(n4284) );
  AND2_X1 U6887 ( .A1(n14969), .A2(n14972), .ZN(n14792) );
  OR2_X1 U6888 ( .A1(n15361), .A2(n4992), .ZN(n15363) );
  AND2_X1 U6889 ( .A1(n15486), .A2(n15491), .ZN(n6245) );
  INV_X1 U6890 ( .A(n15071), .ZN(n5229) );
  AND2_X1 U6891 ( .A1(n15182), .A2(n15190), .ZN(n14645) );
  AOI22_X1 U6892 ( .A1(n13799), .A2(n14063), .B1(n14064), .B2(n13798), .ZN(
        n3564) );
  OR2_X1 U6893 ( .A1(n13817), .A2(n14303), .ZN(n5283) );
  INV_X1 U6894 ( .A(n14533), .ZN(n14649) );
  AND2_X1 U6896 ( .A1(n3348), .A2(n14346), .ZN(n4121) );
  MUX2_X1 U6897 ( .A(n15108), .B(n15410), .S(n14937), .Z(n5788) );
  OR2_X1 U6898 ( .A1(n15109), .A2(n15406), .ZN(n5785) );
  OR2_X1 U6900 ( .A1(n15310), .A2(n15306), .ZN(n5189) );
  INV_X1 U6902 ( .A(n15155), .ZN(n2203) );
  NAND2_X1 U6903 ( .A1(n14733), .A2(n15248), .ZN(n4622) );
  OR2_X1 U6904 ( .A1(n14730), .A2(n15246), .ZN(n4619) );
  INV_X1 U6905 ( .A(n17232), .ZN(n4478) );
  AND2_X1 U6906 ( .A1(n3926), .A2(n15224), .ZN(n3925) );
  OR2_X1 U6907 ( .A1(n13840), .A2(n14007), .ZN(n2561) );
  OR2_X1 U6908 ( .A1(n14134), .A2(n14342), .ZN(n6235) );
  OR2_X1 U6909 ( .A1(n3799), .A2(n3798), .ZN(n13732) );
  OR2_X1 U6910 ( .A1(n15369), .A2(n14737), .ZN(n4458) );
  NOR2_X1 U6911 ( .A1(n14761), .A2(n14248), .ZN(n2729) );
  AOI21_X1 U6912 ( .B1(n14917), .B2(n15489), .A(n14916), .ZN(n5643) );
  AND2_X1 U6913 ( .A1(n6457), .A2(n15316), .ZN(n6456) );
  OR2_X1 U6914 ( .A1(n16888), .A2(n17139), .ZN(n2185) );
  XNOR2_X1 U6915 ( .A(n15281), .B(n15280), .ZN(n5714) );
  OAI211_X1 U6916 ( .C1(n15243), .C2(n15355), .A(n6675), .B(n6674), .ZN(n6673)
         );
  AOI21_X1 U6917 ( .B1(n14149), .B2(n15361), .A(n14751), .ZN(n6672) );
  XNOR2_X1 U6918 ( .A(n2700), .B(n16176), .ZN(n16591) );
  AND2_X1 U6920 ( .A1(n15420), .A2(n15101), .ZN(n14935) );
  XNOR2_X1 U6921 ( .A(n16556), .B(n27422), .ZN(n15568) );
  XNOR2_X1 U6922 ( .A(n16084), .B(n27730), .ZN(n15630) );
  INV_X1 U6923 ( .A(n15781), .ZN(n15654) );
  INV_X1 U6924 ( .A(n17555), .ZN(n17220) );
  OAI21_X1 U6925 ( .B1(n15084), .B2(n4407), .A(n13305), .ZN(n13313) );
  INV_X1 U6926 ( .A(n3374), .ZN(n3138) );
  XNOR2_X1 U6927 ( .A(n16606), .B(n5513), .ZN(n6159) );
  OR2_X1 U6928 ( .A1(n15326), .A2(n15327), .ZN(n3626) );
  OR2_X1 U6929 ( .A1(n14540), .A2(n15202), .ZN(n14541) );
  OAI21_X1 U6930 ( .B1(n14964), .B2(n14539), .A(n14963), .ZN(n14542) );
  AND2_X1 U6931 ( .A1(n17556), .A2(n17553), .ZN(n4099) );
  OR2_X1 U6932 ( .A1(n17455), .A2(n16797), .ZN(n5987) );
  OR2_X1 U6933 ( .A1(n17155), .A2(n28564), .ZN(n5226) );
  INV_X1 U6934 ( .A(n18467), .ZN(n17915) );
  INV_X1 U6935 ( .A(n17138), .ZN(n6727) );
  AND3_X1 U6936 ( .A1(n16612), .A2(n17497), .A3(n17498), .ZN(n18222) );
  OAI21_X1 U6937 ( .B1(n17530), .B2(n17531), .A(n17529), .ZN(n18224) );
  AND2_X1 U6938 ( .A1(n17830), .A2(n4270), .ZN(n5808) );
  AND2_X1 U6939 ( .A1(n17412), .A2(n16831), .ZN(n2485) );
  INV_X1 U6940 ( .A(n17745), .ZN(n2499) );
  AND2_X1 U6941 ( .A1(n17864), .A2(n18527), .ZN(n18541) );
  AOI21_X1 U6943 ( .B1(n18215), .B2(n18216), .A(n520), .ZN(n17868) );
  INV_X1 U6945 ( .A(n18526), .ZN(n5909) );
  OR2_X1 U6947 ( .A1(n18506), .A2(n18215), .ZN(n5157) );
  NOR2_X1 U6948 ( .A1(n18215), .A2(n520), .ZN(n18214) );
  AND2_X1 U6949 ( .A1(n18018), .A2(n18251), .ZN(n2316) );
  AND2_X1 U6950 ( .A1(n1888), .A2(n18020), .ZN(n2814) );
  OR2_X1 U6951 ( .A1(n18471), .A2(n18469), .ZN(n17659) );
  INV_X1 U6952 ( .A(n2819), .ZN(n17709) );
  NOR2_X1 U6953 ( .A1(n18539), .A2(n18260), .ZN(n2707) );
  OR2_X1 U6955 ( .A1(n5695), .A2(n17540), .ZN(n5694) );
  INV_X1 U6956 ( .A(n17261), .ZN(n16779) );
  OR2_X1 U6957 ( .A1(n3880), .A2(n17269), .ZN(n2985) );
  OAI211_X1 U6958 ( .C1(n16802), .C2(n534), .A(n16727), .B(n5585), .ZN(n17695)
         );
  INV_X1 U6960 ( .A(n17347), .ZN(n17345) );
  OR2_X1 U6961 ( .A1(n17439), .A2(n17437), .ZN(n5639) );
  XNOR2_X1 U6962 ( .A(n16464), .B(n4977), .ZN(n16428) );
  AND2_X1 U6963 ( .A1(n16762), .A2(n5398), .ZN(n4787) );
  INV_X1 U6964 ( .A(n17046), .ZN(n6180) );
  MUX2_X1 U6965 ( .A(n16678), .B(n16677), .S(n17456), .Z(n16932) );
  OR2_X1 U6966 ( .A1(n18595), .A2(n17834), .ZN(n3450) );
  INV_X1 U6967 ( .A(n17695), .ZN(n17803) );
  INV_X1 U6968 ( .A(n17719), .ZN(n18524) );
  INV_X1 U6969 ( .A(n18529), .ZN(n18539) );
  AND2_X1 U6970 ( .A1(n18538), .A2(n18537), .ZN(n18054) );
  AND2_X1 U6971 ( .A1(n17942), .A2(n17872), .ZN(n17940) );
  AND2_X1 U6972 ( .A1(n5383), .A2(n18379), .ZN(n17997) );
  OR2_X1 U6973 ( .A1(n2985), .A2(n16996), .ZN(n3343) );
  INV_X1 U6974 ( .A(n17402), .ZN(n4571) );
  OR2_X1 U6975 ( .A1(n14915), .A2(n17402), .ZN(n4112) );
  NOR2_X1 U6977 ( .A1(n20147), .A2(n4877), .ZN(n19010) );
  OAI21_X1 U6978 ( .B1(n17390), .B2(n424), .A(n3090), .ZN(n4040) );
  AND2_X1 U6980 ( .A1(n17562), .A2(n17314), .ZN(n4763) );
  OR2_X1 U6981 ( .A1(n17551), .A2(n17548), .ZN(n17245) );
  AND3_X1 U6982 ( .A1(n17569), .A2(n17229), .A3(n29098), .ZN(n17230) );
  AND2_X1 U6983 ( .A1(n16547), .A2(n16548), .ZN(n16552) );
  OR2_X1 U6984 ( .A1(n16550), .A2(n17508), .ZN(n16551) );
  INV_X1 U6985 ( .A(n3812), .ZN(n16661) );
  AND2_X1 U6986 ( .A1(n18380), .A2(n18379), .ZN(n17165) );
  INV_X1 U6987 ( .A(n17969), .ZN(n18238) );
  INV_X1 U6989 ( .A(n6526), .ZN(n18600) );
  OR2_X1 U6990 ( .A1(n18354), .A2(n18353), .ZN(n5084) );
  OR2_X1 U6991 ( .A1(n18355), .A2(n18353), .ZN(n5589) );
  INV_X1 U6992 ( .A(n17126), .ZN(n3471) );
  AND2_X1 U6993 ( .A1(n18449), .A2(n18195), .ZN(n18454) );
  OAI21_X1 U6994 ( .B1(n16833), .B2(n16834), .A(n16916), .ZN(n16835) );
  OR2_X1 U6995 ( .A1(n17518), .A2(n17516), .ZN(n17108) );
  INV_X1 U6996 ( .A(n18260), .ZN(n2151) );
  OR2_X1 U6997 ( .A1(n4706), .A2(n17451), .ZN(n4702) );
  INV_X1 U6998 ( .A(n5759), .ZN(n19585) );
  AND2_X1 U6999 ( .A1(n17978), .A2(n17979), .ZN(n3439) );
  AOI21_X1 U7000 ( .B1(n18500), .B2(n18213), .A(n18216), .ZN(n5692) );
  INV_X1 U7001 ( .A(n3597), .ZN(n2758) );
  OR2_X1 U7002 ( .A1(n18122), .A2(n18416), .ZN(n3933) );
  OAI211_X1 U7003 ( .C1(n2242), .C2(n17209), .A(n2243), .B(n2241), .ZN(n18690)
         );
  AND2_X1 U7004 ( .A1(n17837), .A2(n18591), .ZN(n2242) );
  INV_X1 U7005 ( .A(n2855), .ZN(n2123) );
  OR2_X1 U7006 ( .A1(n18109), .A2(n17798), .ZN(n18458) );
  OR2_X1 U7007 ( .A1(n18456), .A2(n18107), .ZN(n6038) );
  AND2_X1 U7008 ( .A1(n6912), .A2(n17584), .ZN(n17585) );
  OR2_X1 U7009 ( .A1(n16907), .A2(n17037), .ZN(n5999) );
  INV_X1 U7010 ( .A(n18180), .ZN(n18444) );
  OR2_X1 U7011 ( .A1(n17254), .A2(n17251), .ZN(n5081) );
  INV_X1 U7012 ( .A(n18589), .ZN(n18128) );
  OR2_X1 U7013 ( .A1(n17802), .A2(n18422), .ZN(n17823) );
  NOR2_X1 U7014 ( .A1(n4707), .A2(n18215), .ZN(n4450) );
  INV_X1 U7015 ( .A(n18248), .ZN(n18406) );
  INV_X1 U7016 ( .A(n17858), .ZN(n2694) );
  INV_X1 U7017 ( .A(n18081), .ZN(n18523) );
  AND2_X1 U7018 ( .A1(n18242), .A2(n18236), .ZN(n17967) );
  INV_X1 U7019 ( .A(n18268), .ZN(n18329) );
  AND2_X1 U7020 ( .A1(n18261), .A2(n18268), .ZN(n16930) );
  INV_X1 U7021 ( .A(n16718), .ZN(n18451) );
  AND2_X1 U7023 ( .A1(n18528), .A2(n17701), .ZN(n17703) );
  AND3_X1 U7024 ( .A1(n21066), .A2(n21065), .A3(n21064), .ZN(n21663) );
  OAI211_X1 U7026 ( .C1(n18239), .C2(n29034), .A(n2785), .B(n2784), .ZN(n19354) );
  OR2_X1 U7027 ( .A1(n18230), .A2(n1887), .ZN(n2723) );
  AND2_X1 U7028 ( .A1(n21091), .A2(n29134), .ZN(n20149) );
  AND3_X1 U7029 ( .A1(n4412), .A2(n18371), .A3(n18337), .ZN(n5164) );
  XNOR2_X1 U7030 ( .A(n18735), .B(n6653), .ZN(n18569) );
  INV_X1 U7031 ( .A(n20032), .ZN(n3717) );
  OR2_X1 U7032 ( .A1(n16867), .A2(n5059), .ZN(n5060) );
  INV_X1 U7033 ( .A(n20109), .ZN(n20320) );
  INV_X1 U7034 ( .A(n19669), .ZN(n18726) );
  INV_X1 U7035 ( .A(n3232), .ZN(n4881) );
  OR2_X1 U7036 ( .A1(n17212), .A2(n17211), .ZN(n3719) );
  INV_X1 U7037 ( .A(n19491), .ZN(n6489) );
  AOI21_X1 U7038 ( .B1(n18525), .B2(n18526), .A(n5325), .ZN(n5324) );
  INV_X1 U7039 ( .A(n16990), .ZN(n19525) );
  INV_X1 U7040 ( .A(n19687), .ZN(n5952) );
  OR2_X1 U7041 ( .A1(n20088), .A2(n20090), .ZN(n4006) );
  INV_X1 U7042 ( .A(n20563), .ZN(n20395) );
  AND2_X1 U7043 ( .A1(n20064), .A2(n413), .ZN(n20068) );
  OR2_X1 U7044 ( .A1(n20374), .A2(n19841), .ZN(n20070) );
  AND2_X1 U7045 ( .A1(n19814), .A2(n19815), .ZN(n4657) );
  NOR2_X1 U7046 ( .A1(n2641), .A2(n21442), .ZN(n2640) );
  INV_X1 U7047 ( .A(n2735), .ZN(n20093) );
  OR2_X1 U7048 ( .A1(n20875), .A2(n20814), .ZN(n21265) );
  INV_X1 U7049 ( .A(n20155), .ZN(n19773) );
  OAI21_X1 U7050 ( .B1(n28186), .B2(n20334), .A(n3186), .ZN(n20007) );
  AND2_X1 U7051 ( .A1(n20966), .A2(n21218), .ZN(n20999) );
  OR2_X1 U7052 ( .A1(n20200), .A2(n20205), .ZN(n4338) );
  AND2_X1 U7053 ( .A1(n20121), .A2(n20120), .ZN(n20891) );
  AND2_X1 U7054 ( .A1(n20205), .A2(n20201), .ZN(n2978) );
  OR2_X1 U7055 ( .A1(n20148), .A2(n20146), .ZN(n5794) );
  OR2_X1 U7056 ( .A1(n5334), .A2(n20580), .ZN(n5333) );
  INV_X1 U7057 ( .A(n20404), .ZN(n20554) );
  INV_X1 U7059 ( .A(n21156), .ZN(n3401) );
  AOI22_X1 U7060 ( .A1(n5935), .A2(n20446), .B1(n5934), .B2(n5933), .ZN(n6771)
         );
  AND3_X1 U7061 ( .A1(n21587), .A2(n20591), .A3(n3789), .ZN(n20594) );
  OR2_X1 U7062 ( .A1(n20404), .A2(n20549), .ZN(n20408) );
  OR2_X1 U7063 ( .A1(n20401), .A2(n20208), .ZN(n19743) );
  NOR2_X1 U7064 ( .A1(n20498), .A2(n1624), .ZN(n20008) );
  AND2_X1 U7065 ( .A1(n4148), .A2(n21334), .ZN(n2307) );
  OR2_X1 U7066 ( .A1(n20226), .A2(n1624), .ZN(n5385) );
  OR2_X1 U7067 ( .A1(n21664), .A2(n21665), .ZN(n3692) );
  INV_X1 U7068 ( .A(n5151), .ZN(n21662) );
  OR2_X1 U7069 ( .A1(n4312), .A2(n4309), .ZN(n4308) );
  OR2_X1 U7070 ( .A1(n20513), .A2(n20509), .ZN(n4909) );
  AND2_X1 U7071 ( .A1(n20623), .A2(n20626), .ZN(n6059) );
  AOI21_X1 U7072 ( .B1(n20500), .B2(n20504), .A(n3761), .ZN(n6635) );
  INV_X1 U7074 ( .A(n5106), .ZN(n19860) );
  NOR2_X1 U7075 ( .A1(n21541), .A2(n21539), .ZN(n21499) );
  OR2_X1 U7076 ( .A1(n21500), .A2(n28611), .ZN(n20779) );
  AND2_X1 U7078 ( .A1(n20645), .A2(n21063), .ZN(n5782) );
  NAND2_X1 U7079 ( .A1(n4874), .A2(n4878), .ZN(n20954) );
  AND2_X1 U7080 ( .A1(n21389), .A2(n21387), .ZN(n2572) );
  AND2_X1 U7081 ( .A1(n19993), .A2(n20165), .ZN(n19991) );
  INV_X1 U7083 ( .A(n6314), .ZN(n6311) );
  OR2_X1 U7084 ( .A1(n21265), .A2(n21269), .ZN(n6396) );
  OR2_X1 U7085 ( .A1(n21481), .A2(n21577), .ZN(n6698) );
  INV_X1 U7086 ( .A(n19505), .ZN(n6842) );
  OR2_X1 U7088 ( .A1(n20107), .A2(n20106), .ZN(n3126) );
  OR2_X1 U7089 ( .A1(n20183), .A2(n20182), .ZN(n3076) );
  NOR2_X1 U7090 ( .A1(n21615), .A2(n2339), .ZN(n2338) );
  INV_X1 U7091 ( .A(n21610), .ZN(n2339) );
  INV_X1 U7092 ( .A(n21163), .ZN(n21619) );
  OR2_X1 U7093 ( .A1(n21601), .A2(n21596), .ZN(n21597) );
  OR2_X1 U7094 ( .A1(n19417), .A2(n20688), .ZN(n19418) );
  OR2_X1 U7096 ( .A1(n20746), .A2(n20858), .ZN(n4959) );
  OR2_X1 U7097 ( .A1(n20644), .A2(n5783), .ZN(n4267) );
  INV_X1 U7098 ( .A(n20833), .ZN(n21654) );
  OR2_X1 U7099 ( .A1(n20217), .A2(n5303), .ZN(n2799) );
  INV_X1 U7101 ( .A(n21140), .ZN(n20851) );
  AOI21_X1 U7102 ( .B1(n19779), .B2(n29146), .A(n20084), .ZN(n19780) );
  OR2_X1 U7103 ( .A1(n21311), .A2(n21306), .ZN(n20768) );
  OR2_X1 U7104 ( .A1(n21265), .A2(n29553), .ZN(n6425) );
  OR2_X1 U7105 ( .A1(n19058), .A2(n20174), .ZN(n19009) );
  AND2_X1 U7107 ( .A1(n19966), .A2(n21032), .ZN(n2091) );
  INV_X1 U7108 ( .A(n5194), .ZN(n19965) );
  INV_X1 U7109 ( .A(n5827), .ZN(n21421) );
  NOR2_X1 U7111 ( .A1(n20954), .A2(n20953), .ZN(n21934) );
  AND2_X1 U7112 ( .A1(n3560), .A2(n3559), .ZN(n21936) );
  OR2_X1 U7113 ( .A1(n18787), .A2(n2804), .ZN(n2803) );
  OR2_X1 U7114 ( .A1(n22026), .A2(n22290), .ZN(n3548) );
  INV_X1 U7115 ( .A(n22618), .ZN(n6863) );
  BUF_X1 U7116 ( .A(n21625), .Z(n5339) );
  OR2_X1 U7117 ( .A1(n20600), .A2(n386), .ZN(n4933) );
  INV_X1 U7118 ( .A(n20362), .ZN(n2830) );
  AOI21_X1 U7119 ( .B1(n6533), .B2(n6532), .A(n21106), .ZN(n6531) );
  INV_X1 U7120 ( .A(n21029), .ZN(n6533) );
  OR2_X1 U7121 ( .A1(n20239), .A2(n6512), .ZN(n20003) );
  INV_X1 U7122 ( .A(n21461), .ZN(n5176) );
  INV_X1 U7123 ( .A(n21638), .ZN(n21631) );
  OR2_X1 U7125 ( .A1(n20865), .A2(n20864), .ZN(n21494) );
  OR2_X1 U7127 ( .A1(n5560), .A2(n4877), .ZN(n6894) );
  OR2_X1 U7128 ( .A1(n21113), .A2(n5953), .ZN(n5544) );
  INV_X1 U7129 ( .A(n21464), .ZN(n21560) );
  OAI21_X1 U7130 ( .B1(n5782), .B2(n20646), .A(n5781), .ZN(n20721) );
  INV_X1 U7132 ( .A(n5273), .ZN(n21439) );
  AOI22_X1 U7133 ( .A1(n20232), .A2(n383), .B1(n20231), .B2(n19032), .ZN(n5273) );
  NOR2_X1 U7134 ( .A1(n21655), .A2(n21657), .ZN(n21443) );
  INV_X1 U7135 ( .A(n3954), .ZN(n3952) );
  INV_X1 U7136 ( .A(n21534), .ZN(n21198) );
  INV_X1 U7137 ( .A(n21519), .ZN(n21180) );
  XNOR2_X1 U7138 ( .A(n21825), .B(n3380), .ZN(n3222) );
  INV_X1 U7139 ( .A(n22464), .ZN(n4862) );
  INV_X1 U7140 ( .A(n22337), .ZN(n21889) );
  INV_X1 U7141 ( .A(n22800), .ZN(n20214) );
  XNOR2_X1 U7142 ( .A(n29549), .B(n5797), .ZN(n22706) );
  INV_X1 U7143 ( .A(n3643), .ZN(n5797) );
  AND2_X1 U7144 ( .A1(n339), .A2(n23772), .ZN(n23488) );
  INV_X1 U7145 ( .A(n21872), .ZN(n2752) );
  XNOR2_X1 U7146 ( .A(n22204), .B(n4565), .ZN(n22206) );
  INV_X1 U7147 ( .A(n21789), .ZN(n4565) );
  OR2_X1 U7148 ( .A1(n23741), .A2(n29564), .ZN(n6472) );
  OR2_X1 U7149 ( .A1(n21462), .A2(n20841), .ZN(n3620) );
  OAI21_X1 U7150 ( .B1(n21568), .B2(n21460), .A(n6247), .ZN(n3621) );
  OR2_X1 U7151 ( .A1(n20276), .A2(n6016), .ZN(n6015) );
  AOI21_X1 U7152 ( .B1(n1974), .B2(n20271), .A(n2668), .ZN(n2667) );
  OR2_X1 U7153 ( .A1(n4071), .A2(n21749), .ZN(n6528) );
  AND2_X1 U7154 ( .A1(n23303), .A2(n4178), .ZN(n5697) );
  INV_X1 U7155 ( .A(n4178), .ZN(n5699) );
  INV_X1 U7156 ( .A(n2637), .ZN(n21894) );
  OR2_X1 U7157 ( .A1(n23738), .A2(n23827), .ZN(n3940) );
  AND2_X1 U7158 ( .A1(n23769), .A2(n28554), .ZN(n5237) );
  NOR2_X1 U7159 ( .A1(n23250), .A2(n23406), .ZN(n5042) );
  INV_X1 U7160 ( .A(n23777), .ZN(n23514) );
  BUF_X1 U7161 ( .A(n23167), .Z(n23169) );
  INV_X1 U7163 ( .A(n23656), .ZN(n4772) );
  INV_X1 U7164 ( .A(n24269), .ZN(n2937) );
  NOR2_X1 U7165 ( .A1(n24726), .A2(n24596), .ZN(n5767) );
  OR2_X1 U7166 ( .A1(n5741), .A2(n5448), .ZN(n23191) );
  INV_X1 U7167 ( .A(n407), .ZN(n2281) );
  INV_X1 U7168 ( .A(n4086), .ZN(n4429) );
  INV_X1 U7169 ( .A(n24503), .ZN(n6600) );
  OR2_X1 U7170 ( .A1(n23221), .A2(n6099), .ZN(n5552) );
  OR2_X1 U7171 ( .A1(n24437), .A2(n24436), .ZN(n24121) );
  AND2_X1 U7172 ( .A1(n22977), .A2(n23250), .ZN(n23746) );
  NOR2_X1 U7173 ( .A1(n24288), .A2(n24596), .ZN(n24598) );
  NOR2_X1 U7174 ( .A1(n4020), .A2(n29018), .ZN(n4019) );
  AND2_X1 U7175 ( .A1(n23768), .A2(n23767), .ZN(n6358) );
  OR2_X1 U7176 ( .A1(n2779), .A2(n23651), .ZN(n3135) );
  AOI21_X1 U7177 ( .B1(n22949), .B2(n23398), .A(n23736), .ZN(n22010) );
  NOR2_X1 U7179 ( .A1(n23005), .A2(n23787), .ZN(n6081) );
  INV_X1 U7180 ( .A(n23408), .ZN(n2239) );
  INV_X1 U7181 ( .A(n24447), .ZN(n24761) );
  INV_X1 U7182 ( .A(n23772), .ZN(n23778) );
  INV_X1 U7183 ( .A(n24735), .ZN(n3310) );
  OR2_X1 U7185 ( .A1(n23735), .A2(n2141), .ZN(n3502) );
  INV_X1 U7186 ( .A(n23790), .ZN(n23320) );
  OR2_X1 U7187 ( .A1(n24097), .A2(n24098), .ZN(n3599) );
  INV_X1 U7188 ( .A(n24676), .ZN(n6406) );
  OR2_X1 U7189 ( .A1(n23344), .A2(n23339), .ZN(n6195) );
  OAI211_X1 U7190 ( .C1(n23146), .C2(n4872), .A(n4892), .B(n4891), .ZN(n24295)
         );
  NAND2_X1 U7191 ( .A1(n24610), .A2(n24614), .ZN(n6746) );
  OR2_X1 U7192 ( .A1(n23441), .A2(n2842), .ZN(n23092) );
  NAND2_X1 U7193 ( .A1(n24655), .A2(n2810), .ZN(n24656) );
  OR2_X1 U7194 ( .A1(n23205), .A2(n24555), .ZN(n22747) );
  OAI21_X1 U7196 ( .B1(n3519), .B2(n407), .A(n3518), .ZN(n4175) );
  INV_X1 U7197 ( .A(n5591), .ZN(n3519) );
  INV_X1 U7198 ( .A(n4917), .ZN(n22869) );
  OR2_X1 U7199 ( .A1(n23457), .A2(n23460), .ZN(n23464) );
  OR2_X1 U7200 ( .A1(n23099), .A2(n23418), .ZN(n23100) );
  AND2_X1 U7202 ( .A1(n24666), .A2(n24383), .ZN(n24315) );
  NOR2_X1 U7203 ( .A1(n4851), .A2(n4232), .ZN(n4602) );
  NOR2_X1 U7204 ( .A1(n24592), .A2(n24591), .ZN(n24279) );
  AND2_X1 U7205 ( .A1(n3612), .A2(n23096), .ZN(n22929) );
  INV_X1 U7206 ( .A(n24589), .ZN(n2997) );
  AND2_X1 U7207 ( .A1(n24728), .A2(n24595), .ZN(n5768) );
  INV_X1 U7208 ( .A(n24726), .ZN(n24291) );
  INV_X1 U7209 ( .A(n24479), .ZN(n24210) );
  INV_X1 U7210 ( .A(n23867), .ZN(n24714) );
  NOR2_X1 U7211 ( .A1(n24700), .A2(n24428), .ZN(n24429) );
  INV_X1 U7212 ( .A(n23435), .ZN(n3986) );
  AND2_X1 U7213 ( .A1(n28524), .A2(n24716), .ZN(n24106) );
  INV_X1 U7214 ( .A(n24713), .ZN(n24412) );
  AND2_X1 U7215 ( .A1(n24331), .A2(n2134), .ZN(n3630) );
  NOR2_X1 U7216 ( .A1(n24631), .A2(n24532), .ZN(n24227) );
  NOR2_X1 U7217 ( .A1(n24383), .A2(n24666), .ZN(n24075) );
  INV_X1 U7218 ( .A(n24800), .ZN(n24802) );
  AND2_X1 U7219 ( .A1(n23798), .A2(n23799), .ZN(n6599) );
  AND2_X1 U7220 ( .A1(n4125), .A2(n4124), .ZN(n20656) );
  NOR2_X1 U7221 ( .A1(n24637), .A2(n24636), .ZN(n25797) );
  INV_X1 U7222 ( .A(n23599), .ZN(n23597) );
  AND2_X1 U7223 ( .A1(n24817), .A2(n24809), .ZN(n24496) );
  INV_X1 U7225 ( .A(n2649), .ZN(n24683) );
  OR2_X1 U7226 ( .A1(n405), .A2(n2697), .ZN(n3743) );
  INV_X1 U7227 ( .A(n4596), .ZN(n4595) );
  NOR2_X1 U7228 ( .A1(n24645), .A2(n24638), .ZN(n2107) );
  INV_X1 U7229 ( .A(n24665), .ZN(n4605) );
  INV_X1 U7230 ( .A(n23994), .ZN(n24376) );
  OAI21_X1 U7231 ( .B1(n6211), .B2(n23829), .A(n2188), .ZN(n22947) );
  NAND2_X1 U7232 ( .A1(n23721), .A2(n23394), .ZN(n4473) );
  OR2_X1 U7233 ( .A1(n23287), .A2(n2202), .ZN(n2612) );
  AND2_X1 U7234 ( .A1(n6741), .A2(n24584), .ZN(n22130) );
  INV_X1 U7235 ( .A(n24133), .ZN(n23389) );
  INV_X1 U7236 ( .A(n24081), .ZN(n24386) );
  INV_X1 U7237 ( .A(n24138), .ZN(n25006) );
  INV_X1 U7238 ( .A(n25008), .ZN(n24304) );
  AND2_X1 U7239 ( .A1(n24757), .A2(n24756), .ZN(n2865) );
  AND2_X1 U7240 ( .A1(n24757), .A2(n24447), .ZN(n2866) );
  AND2_X1 U7241 ( .A1(n24800), .A2(n24502), .ZN(n4335) );
  NOR2_X1 U7242 ( .A1(n24789), .A2(n4576), .ZN(n4575) );
  INV_X1 U7246 ( .A(n23004), .ZN(n5350) );
  AND2_X1 U7247 ( .A1(n3199), .A2(n23840), .ZN(n5309) );
  OR2_X1 U7248 ( .A1(n24758), .A2(n24447), .ZN(n24448) );
  INV_X1 U7249 ( .A(n5168), .ZN(n5137) );
  OR2_X1 U7250 ( .A1(n23281), .A2(n23392), .ZN(n5292) );
  NOR2_X1 U7252 ( .A1(n29467), .A2(n26447), .ZN(n26160) );
  OR2_X1 U7253 ( .A1(n6422), .A2(n5633), .ZN(n5632) );
  OR2_X1 U7255 ( .A1(n26386), .A2(n27165), .ZN(n3190) );
  OR2_X1 U7256 ( .A1(n24708), .A2(n24707), .ZN(n5750) );
  INV_X1 U7257 ( .A(n24963), .ZN(n26120) );
  AND3_X1 U7258 ( .A1(n24138), .A2(n24369), .A3(n25008), .ZN(n24139) );
  OAI21_X1 U7259 ( .B1(n26739), .B2(n25655), .A(n26737), .ZN(n5422) );
  NOR2_X1 U7260 ( .A1(n25618), .A2(n280), .ZN(n27392) );
  NOR2_X1 U7261 ( .A1(n25404), .A2(n27395), .ZN(n26463) );
  INV_X1 U7262 ( .A(n26447), .ZN(n3498) );
  OR2_X1 U7263 ( .A1(n26447), .A2(n26448), .ZN(n3497) );
  OR2_X1 U7264 ( .A1(n26920), .A2(n4820), .ZN(n3066) );
  INV_X1 U7265 ( .A(n4820), .ZN(n26173) );
  AND2_X1 U7266 ( .A1(n26172), .A2(n26919), .ZN(n26918) );
  OR2_X1 U7267 ( .A1(n26366), .A2(n29293), .ZN(n2139) );
  OR2_X1 U7268 ( .A1(n27181), .A2(n25034), .ZN(n26270) );
  XNOR2_X1 U7269 ( .A(n24918), .B(n24919), .ZN(n2145) );
  OAI211_X1 U7270 ( .C1(n26858), .C2(n28487), .A(n27138), .B(n29633), .ZN(
        n27688) );
  NOR2_X1 U7271 ( .A1(n28536), .A2(n27131), .ZN(n4080) );
  INV_X1 U7272 ( .A(n27175), .ZN(n27173) );
  OAI211_X1 U7273 ( .C1(n27073), .C2(n27072), .A(n3786), .B(n3785), .ZN(n27080) );
  AOI21_X1 U7274 ( .B1(n28101), .B2(n5036), .A(n26747), .ZN(n26635) );
  AND2_X1 U7275 ( .A1(n5144), .A2(n26251), .ZN(n26253) );
  OR2_X1 U7276 ( .A1(n29482), .A2(n26995), .ZN(n5144) );
  AND2_X1 U7277 ( .A1(n26757), .A2(n29479), .ZN(n6625) );
  NOR2_X1 U7278 ( .A1(n28107), .A2(n28794), .ZN(n28110) );
  OR2_X1 U7279 ( .A1(n25665), .A2(n26723), .ZN(n6288) );
  AND2_X1 U7281 ( .A1(n29541), .A2(n623), .ZN(n6621) );
  NOR2_X1 U7282 ( .A1(n27362), .A2(n25358), .ZN(n25360) );
  OR2_X1 U7283 ( .A1(n27377), .A2(n27213), .ZN(n4091) );
  OR2_X1 U7284 ( .A1(n27213), .A2(n28393), .ZN(n5374) );
  OR2_X1 U7285 ( .A1(n5581), .A2(n27382), .ZN(n4033) );
  OR2_X1 U7286 ( .A1(n27394), .A2(n6685), .ZN(n27396) );
  INV_X1 U7287 ( .A(n27425), .ZN(n6738) );
  AOI21_X1 U7288 ( .B1(n26171), .B2(n26782), .A(n26917), .ZN(n4816) );
  AND2_X1 U7289 ( .A1(n29468), .A2(n449), .ZN(n27446) );
  OAI211_X1 U7290 ( .C1(n26926), .C2(n4400), .A(n2050), .B(n4399), .ZN(n4823)
         );
  AOI21_X1 U7291 ( .B1(n5505), .B2(n4402), .A(n4401), .ZN(n4400) );
  OR2_X1 U7292 ( .A1(n27498), .A2(n27493), .ZN(n5605) );
  AOI21_X1 U7293 ( .B1(n6768), .B2(n26935), .A(n456), .ZN(n6766) );
  OAI21_X1 U7294 ( .B1(n26562), .B2(n26561), .A(n26457), .ZN(n2966) );
  BUF_X1 U7295 ( .A(n27526), .Z(n27505) );
  NOR2_X1 U7296 ( .A1(n27524), .A2(n3067), .ZN(n4164) );
  INV_X1 U7297 ( .A(n26151), .ZN(n26921) );
  AND2_X1 U7298 ( .A1(n6095), .A2(n27527), .ZN(n27524) );
  OR2_X1 U7299 ( .A1(n27286), .A2(n2438), .ZN(n2437) );
  NOR2_X1 U7300 ( .A1(n27304), .A2(n27306), .ZN(n6226) );
  MUX2_X1 U7301 ( .A(n26261), .B(n26260), .S(n27168), .Z(n26262) );
  OAI21_X1 U7302 ( .B1(n26381), .B2(n26426), .A(n4944), .ZN(n26277) );
  INV_X1 U7303 ( .A(n27628), .ZN(n27617) );
  INV_X1 U7304 ( .A(n27614), .ZN(n27627) );
  INV_X1 U7305 ( .A(n27650), .ZN(n27636) );
  OR2_X1 U7306 ( .A1(n28655), .A2(n27663), .ZN(n5874) );
  AND2_X1 U7307 ( .A1(n27165), .A2(n27166), .ZN(n6185) );
  INV_X1 U7308 ( .A(n27662), .ZN(n27676) );
  INV_X1 U7309 ( .A(n29117), .ZN(n4250) );
  AND2_X1 U7310 ( .A1(n26311), .A2(n26310), .ZN(n6669) );
  OR2_X1 U7311 ( .A1(n26867), .A2(n29048), .ZN(n3220) );
  OR2_X1 U7312 ( .A1(n29118), .A2(n27772), .ZN(n4248) );
  INV_X1 U7313 ( .A(n27777), .ZN(n27780) );
  NOR2_X1 U7314 ( .A1(n27795), .A2(n27807), .ZN(n27791) );
  OR3_X1 U7315 ( .A1(n29232), .A2(n27790), .A3(n27817), .ZN(n6902) );
  OR2_X1 U7316 ( .A1(n27109), .A2(n26332), .ZN(n3589) );
  AND2_X1 U7317 ( .A1(n3791), .A2(n27859), .ZN(n5294) );
  INV_X1 U7318 ( .A(n27855), .ZN(n3791) );
  NOR2_X1 U7319 ( .A1(n27855), .A2(n27859), .ZN(n4536) );
  OR2_X1 U7320 ( .A1(n27051), .A2(n28446), .ZN(n3351) );
  AND2_X1 U7321 ( .A1(n27925), .A2(n27244), .ZN(n27934) );
  OR2_X1 U7322 ( .A1(n28456), .A2(n27982), .ZN(n3271) );
  NOR2_X1 U7323 ( .A1(n4499), .A2(n398), .ZN(n4498) );
  AOI21_X1 U7324 ( .B1(n4411), .B2(n25968), .A(n27003), .ZN(n25970) );
  AND2_X1 U7325 ( .A1(n29161), .A2(n376), .ZN(n5017) );
  AND2_X1 U7326 ( .A1(n28063), .A2(n28067), .ZN(n28047) );
  OR2_X1 U7327 ( .A1(n26761), .A2(n26754), .ZN(n26238) );
  AND2_X1 U7328 ( .A1(n28065), .A2(n28066), .ZN(n28052) );
  INV_X1 U7329 ( .A(n28101), .ZN(n5037) );
  NOR2_X1 U7330 ( .A1(n28591), .A2(n28107), .ZN(n3691) );
  INV_X1 U7331 ( .A(n2541), .ZN(n3897) );
  INV_X1 U7332 ( .A(n3554), .ZN(n5649) );
  INV_X1 U7333 ( .A(n3660), .ZN(n4923) );
  INV_X1 U7334 ( .A(n3493), .ZN(n3610) );
  INV_X1 U7335 ( .A(n27286), .ZN(n27280) );
  INV_X1 U7336 ( .A(n27259), .ZN(n5426) );
  AND3_X1 U7337 ( .A1(n2267), .A2(n27570), .A3(n27569), .ZN(Ciphertext[79]) );
  OR2_X1 U7338 ( .A1(n27227), .A2(n27732), .ZN(n2792) );
  OR2_X1 U7339 ( .A1(n26872), .A2(n27101), .ZN(n2376) );
  OR2_X1 U7341 ( .A1(n26544), .A2(n3378), .ZN(n26550) );
  OAI21_X1 U7342 ( .B1(n28438), .B2(n4998), .A(n3571), .ZN(n27246) );
  OR2_X1 U7343 ( .A1(n28037), .A2(n26602), .ZN(n5850) );
  OR3_X1 U7344 ( .A1(n22140), .A2(n21627), .A3(n21624), .ZN(n1940) );
  INV_X1 U7345 ( .A(n7867), .ZN(n5149) );
  XNOR2_X1 U7347 ( .A(n13281), .B(n13282), .ZN(n14304) );
  INV_X1 U7348 ( .A(n29610), .ZN(n4751) );
  INV_X1 U7350 ( .A(n20444), .ZN(n5933) );
  INV_X1 U7351 ( .A(n26510), .ZN(n5299) );
  INV_X1 U7352 ( .A(n27854), .ZN(n5295) );
  INV_X1 U7354 ( .A(n20323), .ZN(n2181) );
  XNOR2_X1 U7355 ( .A(n9389), .B(n4716), .ZN(n10687) );
  OR2_X1 U7356 ( .A1(n21601), .A2(n21314), .ZN(n1941) );
  OR2_X1 U7357 ( .A1(n29594), .A2(n18421), .ZN(n1942) );
  INV_X1 U7359 ( .A(n14399), .ZN(n2549) );
  NAND3_X1 U7360 ( .A1(n6899), .A2(n3839), .A3(n4873), .ZN(n17772) );
  INV_X1 U7361 ( .A(n11022), .ZN(n11314) );
  OR2_X1 U7362 ( .A1(n18229), .A2(n29023), .ZN(n1943) );
  XNOR2_X1 U7363 ( .A(n13094), .B(n13093), .ZN(n14132) );
  XNOR2_X1 U7364 ( .A(n12425), .B(n12424), .ZN(n14401) );
  OR3_X1 U7365 ( .A1(n26195), .A2(n29617), .A3(n26469), .ZN(n1944) );
  OR2_X1 U7366 ( .A1(n333), .A2(n6815), .ZN(n1945) );
  OR2_X1 U7367 ( .A1(n20306), .A2(n19947), .ZN(n1946) );
  OR2_X1 U7368 ( .A1(n11361), .A2(n15576), .ZN(n1947) );
  OR2_X1 U7369 ( .A1(n21626), .A2(n22139), .ZN(n1948) );
  OR2_X1 U7370 ( .A1(n19939), .A2(n28657), .ZN(n1949) );
  AND2_X1 U7371 ( .A1(n28536), .A2(n28480), .ZN(n1950) );
  OR2_X1 U7373 ( .A1(n498), .A2(n20636), .ZN(n1951) );
  AND2_X1 U7374 ( .A1(n2735), .A2(n20088), .ZN(n1952) );
  OR2_X1 U7375 ( .A1(n17502), .A2(n17140), .ZN(n1953) );
  OR2_X1 U7376 ( .A1(n17764), .A2(n28073), .ZN(n1954) );
  INV_X1 U7377 ( .A(n1928), .ZN(n4359) );
  INV_X1 U7378 ( .A(n24141), .ZN(n24277) );
  INV_X1 U7379 ( .A(n12264), .ZN(n12134) );
  NAND2_X1 U7380 ( .A1(n9865), .A2(n12194), .ZN(n11816) );
  INV_X1 U7381 ( .A(n6114), .ZN(n20174) );
  INV_X1 U7382 ( .A(n7362), .ZN(n3431) );
  INV_X1 U7383 ( .A(n12231), .ZN(n13087) );
  XOR2_X1 U7384 ( .A(n13040), .B(n13510), .Z(n1956) );
  INV_X1 U7385 ( .A(n27701), .ZN(n6008) );
  INV_X1 U7386 ( .A(n17829), .ZN(n4273) );
  XOR2_X1 U7387 ( .A(n15396), .B(n16468), .Z(n1957) );
  XOR2_X1 U7388 ( .A(n25249), .B(n3607), .Z(n1958) );
  OAI211_X1 U7392 ( .C1(n11952), .C2(n11951), .A(n11950), .B(n11949), .ZN(
        n13008) );
  INV_X1 U7393 ( .A(n20443), .ZN(n3247) );
  INV_X1 U7394 ( .A(n23305), .ZN(n4020) );
  INV_X1 U7395 ( .A(n4037), .ZN(n12207) );
  INV_X1 U7396 ( .A(n23764), .ZN(n4759) );
  XNOR2_X1 U7397 ( .A(n26078), .B(n26079), .ZN(n27136) );
  AND2_X1 U7399 ( .A1(n14193), .A2(n14192), .ZN(n1959) );
  INV_X1 U7401 ( .A(n10453), .ZN(n11875) );
  INV_X1 U7402 ( .A(n18233), .ZN(n18399) );
  INV_X1 U7403 ( .A(n21481), .ZN(n21580) );
  INV_X1 U7404 ( .A(n17359), .ZN(n2449) );
  OR2_X1 U7406 ( .A1(n14366), .A2(n14123), .ZN(n1960) );
  OR2_X1 U7407 ( .A1(n13907), .A2(n14051), .ZN(n1961) );
  INV_X1 U7408 ( .A(n23529), .ZN(n23697) );
  INV_X1 U7410 ( .A(n18179), .ZN(n4929) );
  OR2_X1 U7411 ( .A1(n21369), .A2(n21716), .ZN(n1962) );
  AND2_X1 U7412 ( .A1(n5919), .A2(n5921), .ZN(n1963) );
  OR2_X1 U7413 ( .A1(n15395), .A2(n15394), .ZN(n1964) );
  OR2_X1 U7414 ( .A1(n28506), .A2(n5193), .ZN(n1965) );
  INV_X1 U7415 ( .A(n2846), .ZN(n12224) );
  AND2_X1 U7416 ( .A1(n6704), .A2(n6703), .ZN(n1966) );
  INV_X1 U7417 ( .A(n9312), .ZN(n5412) );
  INV_X1 U7418 ( .A(n24751), .ZN(n2879) );
  NOR2_X1 U7419 ( .A1(n26260), .A2(n6087), .ZN(n1968) );
  INV_X1 U7420 ( .A(n22143), .ZN(n6532) );
  AOI21_X1 U7421 ( .B1(n27021), .B2(n27020), .A(n27019), .ZN(n27938) );
  INV_X1 U7422 ( .A(n18595), .ZN(n5476) );
  INV_X1 U7425 ( .A(n15415), .ZN(n3922) );
  AND2_X1 U7426 ( .A1(n14101), .A2(n14231), .ZN(n1969) );
  AND3_X1 U7427 ( .A1(n20294), .A2(n19814), .A3(n19818), .ZN(n1970) );
  NAND2_X1 U7428 ( .A1(n27010), .A2(n27013), .ZN(n1971) );
  OR2_X1 U7429 ( .A1(n19829), .A2(n20588), .ZN(n1972) );
  INV_X1 U7430 ( .A(n21346), .ZN(n3260) );
  XNOR2_X1 U7431 ( .A(n25941), .B(n5186), .ZN(n26299) );
  INV_X1 U7432 ( .A(n17552), .ZN(n4624) );
  INV_X1 U7434 ( .A(n18171), .ZN(n4884) );
  AND2_X1 U7435 ( .A1(n20270), .A2(n3666), .ZN(n1974) );
  INV_X1 U7436 ( .A(n22013), .ZN(n4828) );
  INV_X1 U7437 ( .A(n18527), .ZN(n18535) );
  XNOR2_X1 U7438 ( .A(n9405), .B(n9404), .ZN(n11003) );
  INV_X1 U7439 ( .A(n23768), .ZN(n6462) );
  INV_X1 U7440 ( .A(n10786), .ZN(n4538) );
  INV_X1 U7441 ( .A(n23827), .ZN(n2187) );
  AOI22_X1 U7442 ( .A1(n22745), .A2(n23285), .B1(n22638), .B2(n28594), .ZN(
        n23922) );
  INV_X1 U7443 ( .A(n23922), .ZN(n5168) );
  OR3_X1 U7446 ( .A1(n24502), .A2(n24800), .A3(n24804), .ZN(n1976) );
  XNOR2_X1 U7447 ( .A(n6890), .B(n16537), .ZN(n17065) );
  XNOR2_X1 U7448 ( .A(n7229), .B(n7230), .ZN(n10544) );
  XNOR2_X1 U7449 ( .A(n19600), .B(n19601), .ZN(n20322) );
  INV_X1 U7450 ( .A(n20322), .ZN(n2180) );
  XNOR2_X1 U7451 ( .A(n19142), .B(n19143), .ZN(n20339) );
  INV_X1 U7452 ( .A(n20451), .ZN(n5377) );
  XNOR2_X1 U7453 ( .A(n21799), .B(n21798), .ZN(n23763) );
  XNOR2_X1 U7454 ( .A(n15587), .B(n15586), .ZN(n17335) );
  XNOR2_X1 U7455 ( .A(n25395), .B(n25394), .ZN(n26911) );
  XNOR2_X1 U7457 ( .A(Plaintext[84]), .B(Key[84]), .ZN(n7839) );
  XNOR2_X1 U7459 ( .A(n21992), .B(n21993), .ZN(n23736) );
  XOR2_X1 U7460 ( .A(n16605), .B(n16604), .Z(n1977) );
  AND3_X1 U7461 ( .A1(n26927), .A2(n26489), .A3(n26933), .ZN(n1978) );
  INV_X1 U7462 ( .A(n18203), .ZN(n3995) );
  XNOR2_X1 U7463 ( .A(n24488), .B(n25529), .ZN(n26459) );
  INV_X1 U7464 ( .A(n18033), .ZN(n18155) );
  XOR2_X1 U7465 ( .A(n16339), .B(n16405), .Z(n1979) );
  INV_X1 U7466 ( .A(n27410), .ZN(n4922) );
  XNOR2_X1 U7467 ( .A(n25258), .B(n25259), .ZN(n26761) );
  NAND2_X1 U7469 ( .A1(n25159), .A2(n25158), .ZN(n27202) );
  XNOR2_X1 U7471 ( .A(n18822), .B(n18823), .ZN(n20099) );
  XOR2_X1 U7473 ( .A(n15801), .B(n2995), .Z(n1980) );
  XOR2_X1 U7474 ( .A(n18778), .B(n19225), .Z(n1981) );
  XNOR2_X1 U7475 ( .A(n18555), .B(n18554), .ZN(n19843) );
  XNOR2_X1 U7476 ( .A(n22559), .B(n22560), .ZN(n23738) );
  XOR2_X1 U7477 ( .A(n19110), .B(n1927), .Z(n1982) );
  XOR2_X1 U7478 ( .A(n10363), .B(n3244), .Z(n1983) );
  XNOR2_X1 U7479 ( .A(n20839), .B(n20838), .ZN(n23658) );
  XOR2_X1 U7480 ( .A(n22633), .B(n28294), .Z(n1984) );
  XOR2_X1 U7481 ( .A(n9575), .B(n9512), .Z(n1985) );
  XNOR2_X1 U7482 ( .A(n8455), .B(n8454), .ZN(n10748) );
  XOR2_X1 U7483 ( .A(n13445), .B(n13446), .Z(n1987) );
  XOR2_X1 U7484 ( .A(n9466), .B(n9465), .Z(n1988) );
  XOR2_X1 U7485 ( .A(n19704), .B(n2995), .Z(n1989) );
  XNOR2_X1 U7486 ( .A(n22804), .B(n22803), .ZN(n23418) );
  XNOR2_X1 U7487 ( .A(n22335), .B(n22336), .ZN(n23760) );
  INV_X1 U7488 ( .A(n18251), .ZN(n2834) );
  INV_X1 U7489 ( .A(n6504), .ZN(n22427) );
  XOR2_X1 U7490 ( .A(n8844), .B(n8843), .Z(n1990) );
  AND2_X1 U7493 ( .A1(n8014), .A2(n7141), .ZN(n1991) );
  INV_X1 U7494 ( .A(n21145), .ZN(n21120) );
  OR2_X1 U7495 ( .A1(n18451), .A2(n18198), .ZN(n1992) );
  OR3_X1 U7496 ( .A1(n11979), .A2(n1986), .A3(n375), .ZN(n1993) );
  INV_X1 U7497 ( .A(n22991), .ZN(n22996) );
  AND2_X1 U7498 ( .A1(n27191), .A2(n28513), .ZN(n1994) );
  OR3_X1 U7499 ( .A1(n27175), .A2(n27177), .A3(n27178), .ZN(n1995) );
  OR3_X1 U7500 ( .A1(n26920), .A2(n26782), .A3(n26919), .ZN(n1996) );
  INV_X1 U7501 ( .A(n21095), .ZN(n20147) );
  INV_X1 U7502 ( .A(n20137), .ZN(n2152) );
  XOR2_X1 U7503 ( .A(n16052), .B(n16476), .Z(n1998) );
  AND2_X1 U7504 ( .A1(n11235), .A2(n3441), .ZN(n1999) );
  OR2_X1 U7505 ( .A1(n13716), .A2(n13902), .ZN(n2000) );
  XNOR2_X1 U7506 ( .A(n15579), .B(n15580), .ZN(n17204) );
  NAND2_X1 U7507 ( .A1(n4640), .A2(n20169), .ZN(n21089) );
  XNOR2_X1 U7508 ( .A(n16209), .B(n16210), .ZN(n16887) );
  AND2_X1 U7510 ( .A1(n15382), .A2(n15383), .ZN(n2001) );
  INV_X1 U7511 ( .A(n19995), .ZN(n19997) );
  INV_X1 U7512 ( .A(n18500), .ZN(n18217) );
  AND2_X1 U7513 ( .A1(n15420), .A2(n15102), .ZN(n2002) );
  XOR2_X1 U7514 ( .A(n13552), .B(n27225), .Z(n2003) );
  AND2_X1 U7515 ( .A1(n23801), .A2(n23802), .ZN(n2004) );
  INV_X1 U7516 ( .A(n20858), .ZN(n4960) );
  INV_X1 U7517 ( .A(n2108), .ZN(n4109) );
  XNOR2_X1 U7519 ( .A(Key[0]), .B(Plaintext[0]), .ZN(n7889) );
  AND2_X1 U7522 ( .A1(n9062), .A2(n8872), .ZN(n2006) );
  AND2_X1 U7523 ( .A1(n20064), .A2(n20069), .ZN(n2007) );
  INV_X1 U7524 ( .A(n18261), .ZN(n3833) );
  AND2_X1 U7525 ( .A1(n11574), .A2(n12132), .ZN(n2008) );
  OR2_X1 U7526 ( .A1(n14948), .A2(n15073), .ZN(n2009) );
  INV_X1 U7527 ( .A(n7830), .ZN(n8205) );
  AND2_X1 U7529 ( .A1(n27851), .A2(n27854), .ZN(n2010) );
  OR2_X1 U7530 ( .A1(n27704), .A2(n27161), .ZN(n2011) );
  OR3_X1 U7531 ( .A1(n12578), .A2(n12272), .A3(n12270), .ZN(n2012) );
  OR3_X1 U7532 ( .A1(n24794), .A2(n2937), .A3(n24791), .ZN(n2013) );
  OR3_X1 U7533 ( .A1(n26362), .A2(n26799), .A3(n29573), .ZN(n2014) );
  AND2_X1 U7534 ( .A1(n25239), .A2(n27395), .ZN(n2015) );
  AND2_X1 U7535 ( .A1(n23663), .A2(n23662), .ZN(n2016) );
  INV_X1 U7536 ( .A(n22141), .ZN(n21627) );
  AND2_X1 U7537 ( .A1(n14302), .A2(n29611), .ZN(n2017) );
  OR2_X1 U7538 ( .A1(n14373), .A2(n3860), .ZN(n2018) );
  OR2_X1 U7539 ( .A1(n17686), .A2(n28779), .ZN(n2019) );
  AND2_X1 U7540 ( .A1(n14131), .A2(n13842), .ZN(n2020) );
  INV_X1 U7541 ( .A(n16977), .ZN(n16774) );
  INV_X1 U7542 ( .A(n13602), .ZN(n15404) );
  AND2_X1 U7543 ( .A1(n28090), .A2(n4359), .ZN(n2021) );
  OR2_X1 U7544 ( .A1(n21634), .A2(n21638), .ZN(n2022) );
  OR2_X1 U7545 ( .A1(n20283), .A2(n28657), .ZN(n2023) );
  AND2_X1 U7547 ( .A1(n8593), .A2(n8817), .ZN(n2024) );
  XOR2_X1 U7548 ( .A(n12883), .B(n623), .Z(n2025) );
  AND2_X1 U7549 ( .A1(n21603), .A2(n28442), .ZN(n2026) );
  INV_X1 U7550 ( .A(n6741), .ZN(n24578) );
  AND2_X1 U7551 ( .A1(n12266), .A2(n12267), .ZN(n2027) );
  AND2_X1 U7552 ( .A1(n15054), .A2(n14763), .ZN(n2028) );
  AND2_X1 U7553 ( .A1(n8955), .A2(n8956), .ZN(n2029) );
  AND2_X1 U7554 ( .A1(n17004), .A2(n17003), .ZN(n2030) );
  OR2_X1 U7555 ( .A1(n18588), .A2(n17206), .ZN(n2031) );
  AND2_X1 U7556 ( .A1(n4900), .A2(n4901), .ZN(n2032) );
  XOR2_X1 U7557 ( .A(n10250), .B(n3003), .Z(n2034) );
  XOR2_X1 U7558 ( .A(n10137), .B(n2912), .Z(n2035) );
  INV_X1 U7559 ( .A(n24403), .ZN(n2762) );
  INV_X1 U7560 ( .A(n23648), .ZN(n23654) );
  OR2_X1 U7561 ( .A1(n23612), .A2(n28582), .ZN(n2036) );
  AND2_X1 U7562 ( .A1(n5435), .A2(n5437), .ZN(n2037) );
  INV_X1 U7563 ( .A(n27827), .ZN(n27825) );
  OR2_X1 U7565 ( .A1(n27134), .A2(n27129), .ZN(n2038) );
  INV_X1 U7566 ( .A(n5383), .ZN(n18380) );
  INV_X1 U7567 ( .A(n24709), .ZN(n5752) );
  AND2_X1 U7568 ( .A1(n5399), .A2(n4795), .ZN(n2039) );
  AND2_X1 U7570 ( .A1(n15382), .A2(n15151), .ZN(n2040) );
  OR2_X1 U7571 ( .A1(n22142), .A2(n19760), .ZN(n2041) );
  AND2_X1 U7572 ( .A1(n24515), .A2(n24514), .ZN(n3671) );
  AND2_X1 U7573 ( .A1(n8077), .A2(n8428), .ZN(n2042) );
  OR2_X1 U7574 ( .A1(n26455), .A2(n26454), .ZN(n2043) );
  OR2_X1 U7575 ( .A1(n18129), .A2(n17839), .ZN(n2044) );
  NOR2_X1 U7576 ( .A1(n13684), .A2(n3580), .ZN(n14989) );
  INV_X1 U7577 ( .A(n14989), .ZN(n3210) );
  OR2_X1 U7580 ( .A1(n23469), .A2(n3135), .ZN(n2046) );
  INV_X1 U7581 ( .A(n12201), .ZN(n5825) );
  OR2_X1 U7582 ( .A1(n5777), .A2(n15235), .ZN(n2047) );
  NAND2_X1 U7583 ( .A1(n17527), .A2(n6161), .ZN(n2048) );
  INV_X1 U7584 ( .A(n10558), .ZN(n11345) );
  INV_X1 U7585 ( .A(n27843), .ZN(n27828) );
  AND2_X1 U7586 ( .A1(n2259), .A2(n2258), .ZN(n2049) );
  NAND2_X1 U7587 ( .A1(n26929), .A2(n26489), .ZN(n2050) );
  OR2_X1 U7588 ( .A1(n26234), .A2(n26235), .ZN(n2051) );
  XNOR2_X1 U7589 ( .A(n9489), .B(n9490), .ZN(n11253) );
  OR2_X1 U7590 ( .A1(n17156), .A2(n17336), .ZN(n2052) );
  NAND3_X1 U7591 ( .A1(n29161), .A2(n29032), .A3(n29031), .ZN(n2053) );
  OR2_X1 U7592 ( .A1(n23724), .A2(n22455), .ZN(n2054) );
  AND2_X1 U7594 ( .A1(n3811), .A2(n5620), .ZN(n2055) );
  AND2_X1 U7595 ( .A1(n29572), .A2(n17395), .ZN(n2056) );
  INV_X1 U7596 ( .A(n15828), .ZN(n15007) );
  OR2_X1 U7597 ( .A1(n17386), .A2(n17385), .ZN(n2057) );
  NAND2_X1 U7598 ( .A1(n23141), .A2(n5773), .ZN(n2058) );
  OR2_X1 U7599 ( .A1(n7651), .A2(n29081), .ZN(n2059) );
  INV_X1 U7600 ( .A(n21586), .ZN(n3789) );
  INV_X1 U7601 ( .A(n11550), .ZN(n3900) );
  AND2_X1 U7602 ( .A1(n27938), .A2(n28439), .ZN(n2060) );
  OR2_X1 U7603 ( .A1(n17313), .A2(n17315), .ZN(n2061) );
  AND2_X1 U7606 ( .A1(n20476), .A2(n20475), .ZN(n2062) );
  INV_X1 U7607 ( .A(n11194), .ZN(n5838) );
  INV_X1 U7608 ( .A(n21575), .ZN(n21577) );
  OAI211_X1 U7609 ( .C1(n20070), .C2(n20379), .A(n20071), .B(n19842), .ZN(
        n21575) );
  INV_X1 U7610 ( .A(n24155), .ZN(n24523) );
  NAND2_X1 U7611 ( .A1(n28206), .A2(n11144), .ZN(n2063) );
  NAND2_X1 U7612 ( .A1(n25750), .A2(n27076), .ZN(n2064) );
  OR2_X1 U7613 ( .A1(n24609), .A2(n29109), .ZN(n2065) );
  OR2_X1 U7614 ( .A1(n23637), .A2(n29061), .ZN(n2066) );
  AND2_X1 U7615 ( .A1(n20783), .A2(n21177), .ZN(n2067) );
  OR2_X1 U7616 ( .A1(n3830), .A2(n13910), .ZN(n2068) );
  OR2_X1 U7617 ( .A1(n17342), .A2(n16711), .ZN(n2069) );
  AND2_X1 U7618 ( .A1(n23839), .A2(n23392), .ZN(n2070) );
  OR2_X1 U7619 ( .A1(n7534), .A2(n7749), .ZN(n2071) );
  INV_X1 U7621 ( .A(n11430), .ZN(n2748) );
  OR2_X1 U7622 ( .A1(n4097), .A2(n15261), .ZN(n2073) );
  OR2_X1 U7623 ( .A1(n11927), .A2(n11852), .ZN(n2074) );
  OR2_X1 U7624 ( .A1(n14142), .A2(n13900), .ZN(n2075) );
  INV_X1 U7625 ( .A(n28035), .ZN(n6859) );
  INV_X1 U7626 ( .A(n20580), .ZN(n20416) );
  AND2_X1 U7627 ( .A1(n28506), .A2(n5192), .ZN(n2076) );
  OAI21_X1 U7628 ( .B1(n3986), .B2(n23434), .A(n3985), .ZN(n24509) );
  INV_X1 U7629 ( .A(n12257), .ZN(n6687) );
  INV_X1 U7630 ( .A(n24794), .ZN(n4576) );
  INV_X1 U7632 ( .A(n10497), .ZN(n2646) );
  INV_X1 U7633 ( .A(n17977), .ZN(n18234) );
  BUF_X1 U7634 ( .A(n10622), .Z(n11896) );
  INV_X1 U7636 ( .A(n21656), .ZN(n21440) );
  NAND3_X1 U7638 ( .A1(n27076), .A2(n28521), .A3(n29622), .ZN(n2078) );
  INV_X1 U7639 ( .A(n18383), .ZN(n3283) );
  INV_X1 U7640 ( .A(n8929), .ZN(n5958) );
  OR2_X1 U7641 ( .A1(n23576), .A2(n23956), .ZN(n2079) );
  OR2_X1 U7642 ( .A1(n7633), .A2(n7915), .ZN(n2080) );
  AND2_X1 U7643 ( .A1(n4581), .A2(n20282), .ZN(n2081) );
  OR2_X1 U7644 ( .A1(n20321), .A2(n2180), .ZN(n2082) );
  INV_X1 U7646 ( .A(n17088), .ZN(n17504) );
  INV_X1 U7647 ( .A(n3501), .ZN(n5513) );
  INV_X1 U7648 ( .A(n900), .ZN(n4501) );
  INV_X1 U7649 ( .A(n3666), .ZN(n6016) );
  INV_X1 U7650 ( .A(n1172), .ZN(n4607) );
  INV_X1 U7651 ( .A(n72), .ZN(n4070) );
  INV_X1 U7652 ( .A(n1923), .ZN(n4222) );
  INV_X1 U7653 ( .A(n3036), .ZN(n2116) );
  INV_X1 U7654 ( .A(n3062), .ZN(n6653) );
  INV_X1 U7655 ( .A(n26032), .ZN(n2117) );
  INV_X1 U7656 ( .A(n1215), .ZN(n5892) );
  INV_X1 U7657 ( .A(n3003), .ZN(n6174) );
  INV_X1 U7658 ( .A(n3710), .ZN(n5802) );
  INV_X1 U7659 ( .A(n15576), .ZN(n6319) );
  NAND2_X1 U7660 ( .A1(n2083), .A2(n21032), .ZN(n21389) );
  NAND3_X1 U7661 ( .A1(n2091), .A2(n19965), .A3(n2083), .ZN(n21731) );
  OAI21_X1 U7662 ( .B1(n19963), .B2(n20548), .A(n20556), .ZN(n2083) );
  NAND2_X1 U7663 ( .A1(n10640), .A2(n11242), .ZN(n2085) );
  NAND2_X1 U7664 ( .A1(n10639), .A2(n1900), .ZN(n2086) );
  NAND2_X1 U7665 ( .A1(n10629), .A2(n11235), .ZN(n2087) );
  OAI22_X1 U7666 ( .A1(n2090), .A2(n7619), .B1(n2088), .B2(n5946), .ZN(n6060)
         );
  NAND2_X1 U7667 ( .A1(n8236), .A2(n2089), .ZN(n2088) );
  INV_X1 U7668 ( .A(n6973), .ZN(n2089) );
  NAND2_X1 U7669 ( .A1(n7919), .A2(n5946), .ZN(n2090) );
  INV_X1 U7670 ( .A(n8231), .ZN(n5946) );
  INV_X1 U7671 ( .A(n6973), .ZN(n8234) );
  XNOR2_X2 U7672 ( .A(n6970), .B(Key[107]), .ZN(n6973) );
  OAI21_X1 U7673 ( .B1(n28114), .B2(n29480), .A(n2092), .ZN(n2093) );
  OAI21_X1 U7674 ( .B1(n28109), .B2(n28110), .A(n28075), .ZN(n2092) );
  XNOR2_X1 U7675 ( .A(n2093), .B(n28116), .ZN(Ciphertext[191]) );
  NAND2_X1 U7676 ( .A1(n26996), .A2(n28532), .ZN(n2094) );
  NAND2_X1 U7677 ( .A1(n2096), .A2(n20222), .ZN(n6577) );
  XNOR2_X1 U7680 ( .A(n2098), .B(n22697), .ZN(n22151) );
  NAND2_X1 U7681 ( .A1(n22147), .A2(n2097), .ZN(n2098) );
  XNOR2_X1 U7682 ( .A(n2098), .B(n22525), .ZN(n22470) );
  NAND2_X1 U7685 ( .A1(n6260), .A2(n6259), .ZN(n2101) );
  NOR2_X1 U7687 ( .A1(n20829), .A2(n2101), .ZN(n20831) );
  OR2_X1 U7688 ( .A1(n2103), .A2(n10821), .ZN(n4945) );
  NOR2_X1 U7689 ( .A1(n4463), .A2(n2102), .ZN(n4462) );
  AND2_X1 U7690 ( .A1(n2103), .A2(n11331), .ZN(n2102) );
  NAND2_X1 U7691 ( .A1(n2104), .A2(n8941), .ZN(n3595) );
  INV_X1 U7692 ( .A(n8553), .ZN(n2104) );
  NAND2_X1 U7693 ( .A1(n24641), .A2(n2107), .ZN(n2105) );
  NAND2_X1 U7694 ( .A1(n23176), .A2(n24195), .ZN(n2106) );
  NAND2_X1 U7696 ( .A1(n27193), .A2(n29585), .ZN(n26140) );
  OAI211_X1 U7697 ( .C1(n4243), .C2(n29585), .A(n27123), .B(n28595), .ZN(
        n26292) );
  NAND2_X1 U7698 ( .A1(n1994), .A2(n29585), .ZN(n4110) );
  MUX2_X1 U7699 ( .A(n27193), .B(n26291), .S(n4109), .Z(n26294) );
  XNOR2_X2 U7700 ( .A(n12434), .B(n4510), .ZN(n13877) );
  NAND3_X1 U7701 ( .A1(n28804), .A2(n13877), .A3(n14402), .ZN(n2110) );
  NAND2_X1 U7703 ( .A1(n14403), .A2(n4509), .ZN(n2111) );
  XNOR2_X1 U7704 ( .A(n29140), .B(n12450), .ZN(n2113) );
  NAND2_X1 U7705 ( .A1(n2114), .A2(n17497), .ZN(n5587) );
  NOR2_X1 U7706 ( .A1(n17496), .A2(n2114), .ZN(n18223) );
  NAND2_X1 U7707 ( .A1(n538), .A2(n17062), .ZN(n2114) );
  NAND2_X1 U7708 ( .A1(n4052), .A2(n2115), .ZN(n4051) );
  NAND2_X1 U7710 ( .A1(n2119), .A2(n23446), .ZN(n2118) );
  NAND2_X1 U7712 ( .A1(n2118), .A2(n2120), .ZN(n22740) );
  NAND2_X1 U7713 ( .A1(n2119), .A2(n23449), .ZN(n4916) );
  NAND2_X1 U7714 ( .A1(n23109), .A2(n23442), .ZN(n2120) );
  NAND2_X1 U7715 ( .A1(n2121), .A2(n5397), .ZN(n4795) );
  NOR2_X1 U7716 ( .A1(n16946), .A2(n2122), .ZN(n2121) );
  INV_X1 U7717 ( .A(n17242), .ZN(n2122) );
  NAND2_X1 U7718 ( .A1(n18149), .A2(n2855), .ZN(n17814) );
  NOR2_X1 U7719 ( .A1(n18148), .A2(n2123), .ZN(n18151) );
  NOR2_X1 U7720 ( .A1(n3467), .A2(n2855), .ZN(n18049) );
  NAND3_X1 U7721 ( .A1(n420), .A2(n2123), .A3(n3467), .ZN(n18434) );
  XNOR2_X1 U7723 ( .A(n18763), .B(n18764), .ZN(n2124) );
  XNOR2_X2 U7724 ( .A(n2124), .B(n3912), .ZN(n20049) );
  AND2_X1 U7725 ( .A1(n20066), .A2(n413), .ZN(n6477) );
  NAND2_X1 U7726 ( .A1(n2125), .A2(n21811), .ZN(n21382) );
  NOR2_X1 U7727 ( .A1(n19732), .A2(n2125), .ZN(n20983) );
  NOR2_X1 U7728 ( .A1(n21809), .A2(n2125), .ZN(n20980) );
  NAND3_X1 U7729 ( .A1(n21809), .A2(n21806), .A3(n2125), .ZN(n21255) );
  NAND3_X1 U7730 ( .A1(n21809), .A2(n19732), .A3(n2125), .ZN(n19734) );
  NAND2_X1 U7731 ( .A1(n2127), .A2(n28208), .ZN(n10745) );
  NAND2_X1 U7733 ( .A1(n10467), .A2(n2127), .ZN(n8423) );
  NOR2_X1 U7734 ( .A1(n29310), .A2(n2128), .ZN(n10233) );
  INV_X1 U7735 ( .A(n8605), .ZN(n2128) );
  NAND2_X1 U7736 ( .A1(n2129), .A2(n9087), .ZN(n9088) );
  INV_X1 U7737 ( .A(n9081), .ZN(n2129) );
  INV_X1 U7738 ( .A(n2131), .ZN(n2130) );
  NAND2_X1 U7739 ( .A1(n24676), .A2(n29555), .ZN(n2132) );
  MUX2_X1 U7740 ( .A(n29483), .B(n17548), .S(n4218), .Z(n17054) );
  NAND2_X1 U7741 ( .A1(n4787), .A2(n2133), .ZN(n16763) );
  OAI22_X1 U7742 ( .A1(n2134), .A2(n24426), .B1(n28531), .B2(n24772), .ZN(
        n24430) );
  NAND2_X1 U7743 ( .A1(n5248), .A2(n24769), .ZN(n2134) );
  NAND2_X1 U7746 ( .A1(n2137), .A2(n13718), .ZN(n13723) );
  NAND2_X1 U7749 ( .A1(n27134), .A2(n29293), .ZN(n2140) );
  NAND2_X1 U7750 ( .A1(n23256), .A2(n2141), .ZN(n23732) );
  NOR2_X1 U7751 ( .A1(n23398), .A2(n2141), .ZN(n22950) );
  MUX2_X1 U7752 ( .A(n3432), .B(n22949), .S(n23397), .Z(n23232) );
  NAND2_X1 U7753 ( .A1(n11377), .A2(n12102), .ZN(n11655) );
  XNOR2_X2 U7754 ( .A(Key[11]), .B(Plaintext[11]), .ZN(n7770) );
  INV_X1 U7755 ( .A(n12104), .ZN(n11662) );
  NAND2_X1 U7757 ( .A1(n11659), .A2(n29116), .ZN(n2142) );
  AOI21_X1 U7758 ( .B1(n2144), .B2(n14037), .A(n14036), .ZN(n14042) );
  NAND2_X1 U7759 ( .A1(n28513), .A2(n27190), .ZN(n24920) );
  MUX2_X1 U7760 ( .A(n27190), .B(n28513), .S(n27191), .Z(n27192) );
  MUX2_X1 U7761 ( .A(n28595), .B(n4227), .S(n27123), .Z(n27126) );
  NAND2_X1 U7762 ( .A1(n6177), .A2(n2146), .ZN(n16957) );
  NAND2_X1 U7763 ( .A1(n18537), .A2(n18527), .ZN(n2146) );
  NAND2_X1 U7764 ( .A1(n2148), .A2(n18536), .ZN(n2147) );
  NAND2_X1 U7765 ( .A1(n18537), .A2(n2149), .ZN(n2148) );
  NAND2_X1 U7766 ( .A1(n18538), .A2(n18527), .ZN(n2149) );
  NAND2_X1 U7767 ( .A1(n16957), .A2(n2151), .ZN(n2150) );
  XNOR2_X1 U7768 ( .A(n2154), .B(n2509), .ZN(n24671) );
  XNOR2_X1 U7769 ( .A(n25773), .B(n2154), .ZN(n25099) );
  XNOR2_X1 U7770 ( .A(n25391), .B(n2154), .ZN(n25735) );
  NAND3_X1 U7773 ( .A1(n17496), .A2(n4314), .A3(n17062), .ZN(n2157) );
  NAND2_X1 U7774 ( .A1(n2159), .A2(n17492), .ZN(n2158) );
  XNOR2_X2 U7775 ( .A(n16308), .B(n16307), .ZN(n17492) );
  NAND2_X1 U7776 ( .A1(n17497), .A2(n17491), .ZN(n2159) );
  NAND2_X1 U7777 ( .A1(n2161), .A2(n6207), .ZN(n2160) );
  INV_X1 U7778 ( .A(n14761), .ZN(n15261) );
  NAND2_X1 U7780 ( .A1(n2164), .A2(n10991), .ZN(n11694) );
  NAND2_X1 U7781 ( .A1(n10635), .A2(n2165), .ZN(n2164) );
  NAND2_X1 U7783 ( .A1(n12286), .A2(n2166), .ZN(n11625) );
  INV_X1 U7784 ( .A(n12281), .ZN(n2166) );
  INV_X1 U7785 ( .A(n12407), .ZN(n2167) );
  INV_X1 U7786 ( .A(n2168), .ZN(n9567) );
  NAND2_X1 U7788 ( .A1(n23110), .A2(n4794), .ZN(n2169) );
  NAND2_X1 U7790 ( .A1(n6209), .A2(n7506), .ZN(n4129) );
  XNOR2_X2 U7791 ( .A(n7022), .B(Key[56]), .ZN(n7257) );
  NAND2_X1 U7792 ( .A1(n2174), .A2(n23468), .ZN(n25282) );
  NAND3_X1 U7793 ( .A1(n2176), .A2(n6786), .A3(n2175), .ZN(n2174) );
  NAND2_X1 U7794 ( .A1(n6788), .A2(n6787), .ZN(n2176) );
  NAND2_X1 U7795 ( .A1(n20325), .A2(n502), .ZN(n2177) );
  NAND3_X1 U7797 ( .A1(n20324), .A2(n2181), .A3(n2180), .ZN(n2179) );
  NAND2_X1 U7798 ( .A1(n2884), .A2(n20320), .ZN(n2182) );
  OAI21_X1 U7799 ( .B1(n2183), .B2(n17088), .A(n1953), .ZN(n17207) );
  NAND2_X1 U7800 ( .A1(n2186), .A2(n2184), .ZN(n2183) );
  NAND2_X1 U7801 ( .A1(n17501), .A2(n2185), .ZN(n2184) );
  NAND2_X1 U7802 ( .A1(n29127), .A2(n16888), .ZN(n17501) );
  INV_X1 U7803 ( .A(n17087), .ZN(n2186) );
  NAND2_X1 U7804 ( .A1(n23385), .A2(n23825), .ZN(n2189) );
  NAND3_X1 U7805 ( .A1(n23385), .A2(n23825), .A3(n2187), .ZN(n2188) );
  AND2_X1 U7806 ( .A1(n2189), .A2(n3940), .ZN(n23743) );
  AND2_X1 U7807 ( .A1(n4483), .A2(n2189), .ZN(n24090) );
  NAND2_X1 U7808 ( .A1(n20841), .A2(n21459), .ZN(n21571) );
  NAND2_X1 U7810 ( .A1(n2192), .A2(n2191), .ZN(n2190) );
  NAND2_X1 U7811 ( .A1(n14799), .A2(n547), .ZN(n2192) );
  NAND2_X1 U7812 ( .A1(n15185), .A2(n14784), .ZN(n14799) );
  NAND2_X1 U7813 ( .A1(n11487), .A2(n28436), .ZN(n2360) );
  OAI211_X1 U7814 ( .C1(n11430), .C2(n11487), .A(n10717), .B(n2193), .ZN(n2303) );
  INV_X1 U7816 ( .A(n11787), .ZN(n2194) );
  NAND2_X1 U7818 ( .A1(n2200), .A2(n2199), .ZN(n4954) );
  NAND2_X1 U7819 ( .A1(n523), .A2(n18441), .ZN(n2199) );
  NAND2_X1 U7820 ( .A1(n18444), .A2(n18178), .ZN(n2200) );
  NAND2_X1 U7821 ( .A1(n18090), .A2(n18093), .ZN(n18180) );
  NAND2_X1 U7822 ( .A1(n16755), .A2(n16756), .ZN(n18178) );
  AND2_X1 U7823 ( .A1(n22745), .A2(n2202), .ZN(n2201) );
  NAND2_X1 U7824 ( .A1(n2203), .A2(n15379), .ZN(n15380) );
  NAND2_X1 U7825 ( .A1(n2040), .A2(n15155), .ZN(n5815) );
  OAI21_X1 U7826 ( .B1(n15384), .B2(n2203), .A(n2001), .ZN(n15385) );
  INV_X1 U7827 ( .A(n24240), .ZN(n2205) );
  INV_X1 U7829 ( .A(n15565), .ZN(n15452) );
  XNOR2_X1 U7830 ( .A(n15565), .B(n2206), .ZN(n15852) );
  INV_X1 U7831 ( .A(n15940), .ZN(n2206) );
  OAI211_X1 U7832 ( .C1(n28555), .C2(n20614), .A(n20611), .B(n19935), .ZN(
        n4587) );
  OR2_X1 U7833 ( .A1(n29646), .A2(n8131), .ZN(n8050) );
  INV_X1 U7834 ( .A(n7129), .ZN(n8049) );
  OR2_X1 U7835 ( .A1(n6000), .A2(n14091), .ZN(n4721) );
  INV_X1 U7836 ( .A(n24520), .ZN(n3618) );
  XNOR2_X1 U7838 ( .A(n25948), .B(n1172), .ZN(n24529) );
  NOR2_X1 U7839 ( .A1(n17487), .A2(n17489), .ZN(n17151) );
  OR2_X1 U7840 ( .A1(n4884), .A2(n28649), .ZN(n3349) );
  OR2_X1 U7841 ( .A1(n10995), .A2(n10786), .ZN(n10597) );
  NOR2_X1 U7842 ( .A1(n4231), .A2(n5773), .ZN(n4769) );
  AND3_X1 U7843 ( .A1(n5774), .A2(n23011), .A3(n4231), .ZN(n4848) );
  INV_X1 U7844 ( .A(n19025), .ZN(n4883) );
  OAI21_X1 U7845 ( .B1(n8670), .B2(n9107), .A(n8914), .ZN(n8920) );
  INV_X1 U7846 ( .A(n8670), .ZN(n8511) );
  XNOR2_X1 U7847 ( .A(n22526), .B(n21980), .ZN(n22880) );
  AND2_X1 U7848 ( .A1(n7488), .A2(n341), .ZN(n3298) );
  XNOR2_X1 U7849 ( .A(n19685), .B(n3686), .ZN(n4043) );
  XNOR2_X1 U7850 ( .A(n19685), .B(n27811), .ZN(n4746) );
  XNOR2_X1 U7851 ( .A(n15971), .B(n3661), .ZN(n16140) );
  MUX2_X1 U7853 ( .A(n6608), .B(n23792), .S(n23790), .Z(n23498) );
  NOR2_X1 U7854 ( .A1(n5764), .A2(n2640), .ZN(n2639) );
  OR2_X1 U7855 ( .A1(n4734), .A2(n29153), .ZN(n14805) );
  OR2_X1 U7856 ( .A1(n13257), .A2(n14314), .ZN(n6307) );
  OR2_X1 U7857 ( .A1(n11237), .A2(n11236), .ZN(n2413) );
  OR2_X1 U7858 ( .A1(n7898), .A2(n7900), .ZN(n7596) );
  AND2_X1 U7859 ( .A1(n20319), .A2(n20323), .ZN(n2884) );
  AOI21_X1 U7860 ( .B1(n6376), .B2(n18344), .A(n18343), .ZN(n18345) );
  OR2_X1 U7861 ( .A1(n2717), .A2(n7340), .ZN(n2716) );
  INV_X1 U7862 ( .A(n2452), .ZN(n23415) );
  OR2_X1 U7863 ( .A1(n23416), .A2(n2452), .ZN(n2435) );
  OR2_X1 U7864 ( .A1(n15447), .A2(n15323), .ZN(n6521) );
  OR2_X1 U7865 ( .A1(n23535), .A2(n23531), .ZN(n4125) );
  XNOR2_X1 U7866 ( .A(n22698), .B(n22594), .ZN(n3092) );
  NOR2_X1 U7867 ( .A1(n17719), .A2(n18286), .ZN(n18525) );
  AND3_X1 U7868 ( .A1(n17858), .A2(n17719), .A3(n18081), .ZN(n5325) );
  AND2_X1 U7869 ( .A1(n17719), .A2(n17859), .ZN(n16980) );
  AND2_X1 U7870 ( .A1(n4046), .A2(n11430), .ZN(n11302) );
  NOR2_X1 U7872 ( .A1(n24484), .A2(n23968), .ZN(n24212) );
  OR2_X1 U7873 ( .A1(n20488), .A2(n20485), .ZN(n3532) );
  INV_X1 U7874 ( .A(n28620), .ZN(n20240) );
  OR2_X1 U7875 ( .A1(n28620), .A2(n20483), .ZN(n19092) );
  OR2_X1 U7876 ( .A1(n9530), .A2(n9531), .ZN(n3156) );
  NAND2_X1 U7877 ( .A1(n6892), .A2(n9530), .ZN(n7419) );
  INV_X1 U7879 ( .A(n27724), .ZN(n27714) );
  OR2_X1 U7880 ( .A1(n11135), .A2(n3829), .ZN(n3828) );
  XOR2_X1 U7881 ( .A(n10177), .B(n8863), .Z(n8885) );
  XNOR2_X1 U7882 ( .A(n19213), .B(n19214), .ZN(n20343) );
  OR2_X1 U7883 ( .A1(n20725), .A2(n21598), .ZN(n3530) );
  INV_X1 U7884 ( .A(n27773), .ZN(n6419) );
  OR2_X1 U7885 ( .A1(n29537), .A2(n27762), .ZN(n5776) );
  AND2_X1 U7886 ( .A1(n27904), .A2(n29536), .ZN(n27839) );
  INV_X1 U7887 ( .A(n26299), .ZN(n27060) );
  XNOR2_X1 U7888 ( .A(n25942), .B(n25940), .ZN(n5186) );
  XNOR2_X1 U7889 ( .A(n22302), .B(n2752), .ZN(n22235) );
  INV_X1 U7890 ( .A(n14304), .ZN(n5956) );
  AND2_X1 U7891 ( .A1(n11877), .A2(n10868), .ZN(n11879) );
  AND2_X1 U7892 ( .A1(n20636), .A2(n20639), .ZN(n2528) );
  XNOR2_X1 U7893 ( .A(n18900), .B(n28571), .ZN(n6468) );
  INV_X1 U7894 ( .A(n18900), .ZN(n19162) );
  OAI21_X1 U7895 ( .B1(n4667), .B2(n14278), .A(n14363), .ZN(n4666) );
  OAI21_X1 U7897 ( .B1(n27087), .B2(n26841), .A(n2877), .ZN(n27021) );
  OR2_X1 U7899 ( .A1(n17282), .A2(n17283), .ZN(n6380) );
  INV_X1 U7900 ( .A(n13725), .ZN(n5404) );
  MUX2_X1 U7901 ( .A(n8351), .B(n261), .S(n8353), .Z(n8356) );
  OR2_X1 U7902 ( .A1(n23235), .A2(n23716), .ZN(n23265) );
  NAND2_X1 U7903 ( .A1(n23537), .A2(n23541), .ZN(n2636) );
  AND2_X1 U7904 ( .A1(n29508), .A2(n20614), .ZN(n4684) );
  INV_X1 U7905 ( .A(n15727), .ZN(n16427) );
  OR2_X1 U7906 ( .A1(n8785), .A2(n8717), .ZN(n4320) );
  OR2_X1 U7907 ( .A1(n8047), .A2(n7127), .ZN(n7716) );
  INV_X1 U7908 ( .A(n16846), .ZN(n17009) );
  OR2_X1 U7909 ( .A1(n21322), .A2(n5983), .ZN(n21137) );
  NOR2_X1 U7910 ( .A1(n29569), .A2(n21322), .ZN(n20887) );
  XNOR2_X1 U7911 ( .A(n19272), .B(n19534), .ZN(n19598) );
  INV_X1 U7912 ( .A(n2728), .ZN(n5978) );
  INV_X1 U7913 ( .A(n12022), .ZN(n12353) );
  AND2_X1 U7914 ( .A1(n12022), .A2(n11901), .ZN(n10587) );
  INV_X1 U7915 ( .A(n7175), .ZN(n8730) );
  INV_X1 U7917 ( .A(n14008), .ZN(n4586) );
  NOR2_X1 U7918 ( .A1(n10114), .A2(n11120), .ZN(n4383) );
  OR2_X1 U7919 ( .A1(n13932), .A2(n14452), .ZN(n2327) );
  AND2_X1 U7921 ( .A1(n14451), .A2(n14452), .ZN(n3526) );
  OR2_X1 U7922 ( .A1(n12234), .A2(n375), .ZN(n6581) );
  OR2_X1 U7923 ( .A1(n11176), .A2(n434), .ZN(n11340) );
  AOI21_X1 U7924 ( .B1(n7273), .B2(n2104), .A(n9562), .ZN(n7274) );
  OR2_X1 U7925 ( .A1(n10853), .A2(n11163), .ZN(n11057) );
  INV_X1 U7926 ( .A(n15009), .ZN(n3784) );
  AND2_X1 U7927 ( .A1(n15371), .A2(n15009), .ZN(n3840) );
  XNOR2_X1 U7928 ( .A(n19251), .B(n5246), .ZN(n19473) );
  INV_X1 U7929 ( .A(n18799), .ZN(n5246) );
  OR2_X1 U7930 ( .A1(n29152), .A2(n6002), .ZN(n16964) );
  XNOR2_X1 U7931 ( .A(n12787), .B(n13159), .ZN(n12421) );
  AND2_X1 U7932 ( .A1(n29058), .A2(n25676), .ZN(n27003) );
  INV_X1 U7933 ( .A(n25676), .ZN(n27045) );
  XNOR2_X1 U7934 ( .A(n25545), .B(n25544), .ZN(n25676) );
  OR2_X1 U7935 ( .A1(n19761), .A2(n20066), .ZN(n3436) );
  NOR2_X1 U7936 ( .A1(n23233), .A2(n22174), .ZN(n6728) );
  OR2_X1 U7937 ( .A1(n21432), .A2(n21431), .ZN(n4312) );
  OAI21_X1 U7938 ( .B1(n1916), .B2(n20601), .A(n20599), .ZN(n5357) );
  AOI21_X1 U7940 ( .B1(n7362), .B2(n7363), .A(n8205), .ZN(n3429) );
  OR2_X1 U7941 ( .A1(n7886), .A2(n7071), .ZN(n2882) );
  NOR2_X1 U7942 ( .A1(n7585), .A2(n7886), .ZN(n2226) );
  OR2_X1 U7943 ( .A1(n6617), .A2(n27363), .ZN(n6616) );
  NOR2_X1 U7944 ( .A1(n27908), .A2(n27913), .ZN(n27889) );
  OR3_X1 U7945 ( .A1(n27010), .A2(n27013), .A3(n27052), .ZN(n5686) );
  INV_X1 U7946 ( .A(n7967), .ZN(n4697) );
  AND3_X1 U7947 ( .A1(n7965), .A2(n29302), .A3(n7967), .ZN(n5255) );
  OR2_X1 U7948 ( .A1(n7966), .A2(n7967), .ZN(n3226) );
  AOI21_X1 U7949 ( .B1(n27357), .B2(n27356), .A(n6287), .ZN(n2426) );
  OR2_X1 U7950 ( .A1(n20383), .A2(n19836), .ZN(n6237) );
  OR2_X1 U7951 ( .A1(n526), .A2(n18136), .ZN(n18143) );
  OR2_X1 U7952 ( .A1(n14192), .A2(n13953), .ZN(n5378) );
  NAND2_X1 U7953 ( .A1(n10532), .A2(n11294), .ZN(n5563) );
  OR2_X1 U7954 ( .A1(n10891), .A2(n11294), .ZN(n10892) );
  OR2_X1 U7955 ( .A1(n23800), .A2(n4726), .ZN(n5193) );
  OR2_X1 U7956 ( .A1(n4193), .A2(n21459), .ZN(n20754) );
  NAND3_X1 U7957 ( .A1(n2210), .A2(n10951), .A3(n10950), .ZN(n11859) );
  NAND2_X1 U7958 ( .A1(n2211), .A2(n10972), .ZN(n10949) );
  NAND2_X1 U7959 ( .A1(n10971), .A2(n10970), .ZN(n2211) );
  OAI211_X1 U7960 ( .C1(n18599), .C2(n28142), .A(n2213), .B(n6526), .ZN(n2212)
         );
  NAND2_X1 U7961 ( .A1(n17989), .A2(n28142), .ZN(n2213) );
  NAND2_X1 U7962 ( .A1(n28142), .A2(n6927), .ZN(n2215) );
  NAND2_X1 U7964 ( .A1(n2218), .A2(n2217), .ZN(n13036) );
  NAND3_X1 U7965 ( .A1(n2219), .A2(n10700), .A3(n11363), .ZN(n2218) );
  NAND2_X1 U7966 ( .A1(n2220), .A2(n4712), .ZN(n10515) );
  NAND2_X1 U7967 ( .A1(n6075), .A2(n11870), .ZN(n2220) );
  AND2_X1 U7968 ( .A1(n8658), .A2(n8502), .ZN(n8634) );
  NAND2_X1 U7969 ( .A1(n2226), .A2(n2225), .ZN(n2221) );
  NAND2_X1 U7970 ( .A1(n2224), .A2(n2223), .ZN(n2222) );
  INV_X1 U7971 ( .A(n7885), .ZN(n2225) );
  NAND3_X1 U7972 ( .A1(n591), .A2(n10972), .A3(n28608), .ZN(n4045) );
  INV_X1 U7974 ( .A(n2232), .ZN(n12015) );
  NAND3_X1 U7975 ( .A1(n11887), .A2(n11886), .A3(n12332), .ZN(n2232) );
  NAND2_X1 U7976 ( .A1(n10535), .A2(n10878), .ZN(n2227) );
  AOI21_X1 U7977 ( .B1(n11222), .B2(n435), .A(n11219), .ZN(n2228) );
  AOI21_X1 U7978 ( .B1(n7410), .B2(n9340), .A(n2230), .ZN(n2229) );
  OAI21_X1 U7979 ( .B1(n9132), .B2(n9340), .A(n8342), .ZN(n2230) );
  OAI21_X1 U7980 ( .B1(n601), .B2(n9131), .A(n2231), .ZN(n9341) );
  NAND3_X1 U7981 ( .A1(n7410), .A2(n8753), .A3(n600), .ZN(n2231) );
  NAND3_X1 U7984 ( .A1(n1166), .A2(n17229), .A3(n17038), .ZN(n2234) );
  NAND3_X1 U7986 ( .A1(n7585), .A2(n7886), .A3(n7071), .ZN(n2236) );
  INV_X2 U7987 ( .A(n7887), .ZN(n7585) );
  NAND3_X1 U7988 ( .A1(n7580), .A2(n7885), .A3(n7583), .ZN(n2237) );
  NAND2_X1 U7989 ( .A1(n2238), .A2(n8521), .ZN(n8524) );
  NAND2_X1 U7990 ( .A1(n2238), .A2(n8811), .ZN(n8813) );
  NAND3_X1 U7991 ( .A1(n2238), .A2(n8521), .A3(n8809), .ZN(n8252) );
  AOI21_X1 U7992 ( .B1(n8460), .B2(n8681), .A(n2238), .ZN(n8461) );
  MUX2_X1 U7993 ( .A(n20444), .B(n20443), .S(n6843), .Z(n19926) );
  OAI22_X1 U7994 ( .A1(n23747), .A2(n2239), .B1(n22978), .B2(n409), .ZN(n22983) );
  OAI21_X1 U7995 ( .B1(n23404), .B2(n23746), .A(n2239), .ZN(n5971) );
  NAND2_X1 U7996 ( .A1(n2240), .A2(n24435), .ZN(n24348) );
  NAND2_X1 U7997 ( .A1(n403), .A2(n2240), .ZN(n5348) );
  NAND2_X1 U7998 ( .A1(n24433), .A2(n24434), .ZN(n24188) );
  NAND2_X1 U7999 ( .A1(n18588), .A2(n18595), .ZN(n17837) );
  NAND2_X1 U8000 ( .A1(n17840), .A2(n17835), .ZN(n2241) );
  NAND2_X1 U8001 ( .A1(n17208), .A2(n18129), .ZN(n2243) );
  OAI21_X1 U8003 ( .B1(n14958), .B2(n13865), .A(n2244), .ZN(n13866) );
  NAND2_X1 U8004 ( .A1(n13861), .A2(n14958), .ZN(n2244) );
  NAND2_X1 U8006 ( .A1(n2246), .A2(n24810), .ZN(n3001) );
  NOR2_X1 U8007 ( .A1(n2251), .A2(n9009), .ZN(n2248) );
  INV_X1 U8009 ( .A(n9009), .ZN(n9191) );
  INV_X1 U8010 ( .A(n9184), .ZN(n2251) );
  OR2_X1 U8012 ( .A1(n7362), .A2(n7363), .ZN(n8200) );
  NAND2_X1 U8013 ( .A1(n10110), .A2(n10592), .ZN(n2255) );
  NAND2_X1 U8014 ( .A1(n9281), .A2(n10705), .ZN(n2256) );
  NAND2_X1 U8015 ( .A1(n2688), .A2(n2689), .ZN(n11024) );
  XNOR2_X1 U8017 ( .A(n4042), .B(n4043), .ZN(n2257) );
  NAND2_X1 U8020 ( .A1(n20980), .A2(n21811), .ZN(n2258) );
  MUX2_X1 U8022 ( .A(n24736), .B(n24735), .S(n24734), .Z(n24743) );
  NAND2_X1 U8023 ( .A1(n6118), .A2(n2260), .ZN(n6117) );
  NAND2_X1 U8024 ( .A1(n20726), .A2(n20986), .ZN(n2260) );
  NAND2_X1 U8025 ( .A1(n20177), .A2(n20173), .ZN(n19058) );
  XNOR2_X1 U8026 ( .A(n19606), .B(n19103), .ZN(n18746) );
  NAND3_X1 U8028 ( .A1(n18524), .A2(n18523), .A3(n17858), .ZN(n17722) );
  XNOR2_X1 U8030 ( .A(n15007), .B(n15452), .ZN(n4990) );
  AND3_X2 U8031 ( .A1(n2796), .A2(n2799), .A3(n2798), .ZN(n21655) );
  INV_X1 U8032 ( .A(n7525), .ZN(n7531) );
  NAND2_X1 U8033 ( .A1(n8014), .A2(n7533), .ZN(n7525) );
  NAND2_X1 U8035 ( .A1(n14776), .A2(n14777), .ZN(n16012) );
  NAND2_X1 U8036 ( .A1(n18488), .A2(n18489), .ZN(n15734) );
  NAND2_X1 U8037 ( .A1(n17146), .A2(n17076), .ZN(n16734) );
  NAND2_X1 U8038 ( .A1(n1831), .A2(n11755), .ZN(n11760) );
  OR2_X1 U8039 ( .A1(n29114), .A2(n28820), .ZN(n18790) );
  INV_X1 U8040 ( .A(n17235), .ZN(n2701) );
  NAND3_X1 U8043 ( .A1(n28068), .A2(n28067), .A3(n28069), .ZN(n3262) );
  NAND2_X1 U8044 ( .A1(n2263), .A2(n2262), .ZN(n26725) );
  NAND2_X1 U8045 ( .A1(n26720), .A2(n26215), .ZN(n2262) );
  NAND2_X1 U8046 ( .A1(n26719), .A2(n26718), .ZN(n2263) );
  NAND2_X1 U8049 ( .A1(n23894), .A2(n24322), .ZN(n2265) );
  OR2_X1 U8050 ( .A1(n23896), .A2(n24678), .ZN(n2266) );
  NAND2_X1 U8051 ( .A1(n27568), .A2(n2268), .ZN(n2267) );
  MUX2_X1 U8053 ( .A(n25833), .B(n25832), .S(n26842), .Z(n25834) );
  NAND3_X1 U8054 ( .A1(n2332), .A2(n2333), .A3(n811), .ZN(n24080) );
  NAND2_X1 U8056 ( .A1(n26333), .A2(n26836), .ZN(n2269) );
  NAND2_X1 U8057 ( .A1(n9197), .A2(n9206), .ZN(n9000) );
  NAND2_X1 U8058 ( .A1(n7637), .A2(n3428), .ZN(n9197) );
  NAND2_X1 U8059 ( .A1(n7362), .A2(n7634), .ZN(n7636) );
  NAND2_X1 U8061 ( .A1(n6685), .A2(n28908), .ZN(n24362) );
  NAND2_X1 U8062 ( .A1(n24827), .A2(n24828), .ZN(n24829) );
  NAND2_X1 U8063 ( .A1(n20027), .A2(n20273), .ZN(n20030) );
  NAND2_X1 U8065 ( .A1(n10447), .A2(n10446), .ZN(n2271) );
  NAND2_X1 U8067 ( .A1(n7813), .A2(n28627), .ZN(n2273) );
  NAND2_X1 U8069 ( .A1(n27827), .A2(n2275), .ZN(n5336) );
  NAND2_X1 U8070 ( .A1(n27841), .A2(n27101), .ZN(n2275) );
  NAND3_X1 U8071 ( .A1(n2276), .A2(n27765), .A3(n27764), .ZN(n27767) );
  NAND2_X1 U8072 ( .A1(n27785), .A2(n6419), .ZN(n2276) );
  OAI21_X1 U8075 ( .B1(n15055), .B2(n15259), .A(n2278), .ZN(n4418) );
  NAND2_X1 U8076 ( .A1(n15259), .A2(n14761), .ZN(n2278) );
  NAND2_X1 U8077 ( .A1(n5684), .A2(n21322), .ZN(n21588) );
  NAND3_X2 U8078 ( .A1(n3194), .A2(n3193), .A3(n20555), .ZN(n21322) );
  NAND2_X1 U8081 ( .A1(n19561), .A2(n19562), .ZN(n17797) );
  NAND2_X1 U8083 ( .A1(n3552), .A2(n12255), .ZN(n2709) );
  NAND3_X1 U8084 ( .A1(n7769), .A2(n7768), .A3(n7767), .ZN(n3183) );
  XOR2_X1 U8086 ( .A(n9619), .B(n629), .Z(n5896) );
  AOI21_X2 U8087 ( .B1(n2281), .B2(n2282), .A(n22862), .ZN(n4917) );
  INV_X1 U8088 ( .A(n22861), .ZN(n2282) );
  INV_X1 U8089 ( .A(n10657), .ZN(n11222) );
  XNOR2_X1 U8090 ( .A(n4493), .B(n16283), .ZN(n15965) );
  INV_X1 U8091 ( .A(n7496), .ZN(n3594) );
  AND2_X1 U8092 ( .A1(n4320), .A2(n8367), .ZN(n2340) );
  XNOR2_X1 U8093 ( .A(n10063), .B(n10062), .ZN(n5150) );
  NAND2_X1 U8097 ( .A1(n8993), .A2(n9434), .ZN(n3056) );
  XNOR2_X1 U8098 ( .A(n2285), .B(n25054), .ZN(n25058) );
  XNOR2_X1 U8099 ( .A(n25053), .B(n26108), .ZN(n2285) );
  NAND2_X1 U8100 ( .A1(n26781), .A2(n26919), .ZN(n3390) );
  NAND2_X1 U8102 ( .A1(n4672), .A2(n22863), .ZN(n6338) );
  NOR2_X1 U8105 ( .A1(n23067), .A2(n28164), .ZN(n2286) );
  INV_X1 U8107 ( .A(n23137), .ZN(n23136) );
  NAND2_X1 U8108 ( .A1(n23067), .A2(n28164), .ZN(n23137) );
  NAND2_X1 U8109 ( .A1(n2289), .A2(n9169), .ZN(n9172) );
  OR2_X1 U8113 ( .A1(n7654), .A2(n7653), .ZN(n7679) );
  AND2_X1 U8114 ( .A1(n10856), .A2(n5835), .ZN(n11313) );
  XNOR2_X1 U8115 ( .A(n2291), .B(n9770), .ZN(n9343) );
  XNOR2_X1 U8116 ( .A(n9339), .B(n10385), .ZN(n2291) );
  INV_X1 U8117 ( .A(n18273), .ZN(n2292) );
  NOR2_X1 U8118 ( .A1(n4211), .A2(n18516), .ZN(n18273) );
  NAND2_X1 U8119 ( .A1(n8178), .A2(n8179), .ZN(n8180) );
  NAND2_X1 U8120 ( .A1(n29631), .A2(n26950), .ZN(n26442) );
  AND2_X1 U8121 ( .A1(n2748), .A2(n6482), .ZN(n11789) );
  OR2_X1 U8122 ( .A1(n20333), .A2(n20630), .ZN(n19328) );
  INV_X1 U8124 ( .A(n14807), .ZN(n14715) );
  INV_X1 U8125 ( .A(n4105), .ZN(n12408) );
  XNOR2_X1 U8126 ( .A(n19183), .B(n18649), .ZN(n20563) );
  XNOR2_X1 U8127 ( .A(n12831), .B(n12828), .ZN(n2293) );
  OR2_X1 U8128 ( .A1(n10318), .A2(n11287), .ZN(n10664) );
  OR2_X1 U8129 ( .A1(n9364), .A2(n3274), .ZN(n3272) );
  INV_X1 U8130 ( .A(n21714), .ZN(n20976) );
  NAND2_X1 U8132 ( .A1(n17004), .A2(n15981), .ZN(n4614) );
  NAND2_X1 U8133 ( .A1(n15423), .A2(n15102), .ZN(n15421) );
  NAND2_X1 U8135 ( .A1(n12888), .A2(n14438), .ZN(n2294) );
  OAI22_X1 U8136 ( .A1(n24674), .A2(n29555), .B1(n24322), .B2(n24397), .ZN(
        n2379) );
  OR2_X1 U8137 ( .A1(n4854), .A2(n18159), .ZN(n17326) );
  NAND2_X1 U8138 ( .A1(n20955), .A2(n21090), .ZN(n2296) );
  XNOR2_X2 U8139 ( .A(n2297), .B(Key[15]), .ZN(n8177) );
  INV_X1 U8140 ( .A(Plaintext[15]), .ZN(n2297) );
  NOR2_X2 U8142 ( .A1(n23491), .A2(n23490), .ZN(n23946) );
  XNOR2_X1 U8145 ( .A(n25772), .B(n2300), .ZN(n25259) );
  XNOR2_X1 U8146 ( .A(n25257), .B(n25546), .ZN(n2300) );
  OAI21_X1 U8147 ( .B1(n21515), .B2(n21516), .A(n2301), .ZN(n21517) );
  NAND3_X1 U8148 ( .A1(n21532), .A2(n21514), .A3(n21513), .ZN(n2301) );
  NAND3_X1 U8150 ( .A1(n3740), .A2(n2832), .A3(n7590), .ZN(n6802) );
  NAND2_X1 U8152 ( .A1(n2335), .A2(n8560), .ZN(n2334) );
  AND2_X1 U8153 ( .A1(n11473), .A2(n12337), .ZN(n5466) );
  NAND2_X1 U8154 ( .A1(n13850), .A2(n14176), .ZN(n2304) );
  OAI211_X1 U8155 ( .C1(n20157), .C2(n20160), .A(n19985), .B(n2305), .ZN(n4235) );
  NAND2_X1 U8156 ( .A1(n20157), .A2(n29066), .ZN(n2305) );
  NAND2_X1 U8157 ( .A1(n21608), .A2(n2307), .ZN(n21335) );
  NAND3_X2 U8158 ( .A1(n2308), .A2(n8450), .A3(n8449), .ZN(n10038) );
  OAI211_X1 U8159 ( .C1(n9195), .C2(n9201), .A(n2309), .B(n8779), .ZN(n2308)
         );
  INV_X1 U8160 ( .A(n8451), .ZN(n2309) );
  INV_X1 U8161 ( .A(n2311), .ZN(n2310) );
  OAI21_X1 U8162 ( .B1(n7347), .B2(n7759), .A(n7763), .ZN(n2311) );
  NAND2_X1 U8163 ( .A1(n21367), .A2(n21366), .ZN(n2312) );
  XOR2_X1 U8165 ( .A(n9678), .B(n9619), .Z(n6796) );
  AOI22_X2 U8166 ( .A1(n4176), .A2(n24408), .B1(n24407), .B2(n24406), .ZN(
        n25345) );
  NOR2_X1 U8167 ( .A1(n17249), .A2(n16977), .ZN(n4863) );
  NAND2_X1 U8168 ( .A1(n2313), .A2(n6699), .ZN(n5577) );
  NAND4_X1 U8169 ( .A1(n14705), .A2(n14447), .A3(n14448), .A4(n14449), .ZN(
        n2313) );
  XNOR2_X1 U8170 ( .A(n15914), .B(n16296), .ZN(n16103) );
  AOI21_X2 U8171 ( .B1(n6262), .B2(n15405), .A(n15404), .ZN(n15914) );
  AOI22_X1 U8172 ( .A1(n421), .A2(n17119), .B1(n17121), .B2(n17120), .ZN(n2314) );
  NAND2_X1 U8173 ( .A1(n15462), .A2(n15464), .ZN(n4513) );
  AND3_X2 U8174 ( .A1(n13883), .A2(n13882), .A3(n13881), .ZN(n15462) );
  NAND2_X1 U8175 ( .A1(n16925), .A2(n16926), .ZN(n16927) );
  NAND2_X1 U8176 ( .A1(n24046), .A2(n24484), .ZN(n24047) );
  NAND3_X1 U8178 ( .A1(n11999), .A2(n11998), .A3(n11997), .ZN(n2604) );
  AOI21_X1 U8179 ( .B1(n21625), .B2(n22145), .A(n22143), .ZN(n21109) );
  OAI21_X1 U8181 ( .B1(n8501), .B2(n8502), .A(n8115), .ZN(n8118) );
  OR2_X2 U8182 ( .A1(n2315), .A2(n9476), .ZN(n13081) );
  AOI21_X1 U8183 ( .B1(n9467), .B2(n10108), .A(n588), .ZN(n2315) );
  NAND2_X1 U8184 ( .A1(n524), .A2(n2316), .ZN(n17578) );
  NAND2_X1 U8185 ( .A1(n2837), .A2(n2836), .ZN(n2318) );
  INV_X1 U8186 ( .A(n10834), .ZN(n3820) );
  INV_X1 U8189 ( .A(n9793), .ZN(n9515) );
  XNOR2_X1 U8190 ( .A(n5818), .B(n9514), .ZN(n9793) );
  XNOR2_X2 U8191 ( .A(n7087), .B(Key[5]), .ZN(n7775) );
  AOI22_X1 U8192 ( .A1(n4433), .A2(n1959), .B1(n13951), .B2(n4049), .ZN(n4050)
         );
  NAND2_X1 U8194 ( .A1(n8767), .A2(n604), .ZN(n8580) );
  NAND2_X1 U8195 ( .A1(n2496), .A2(n15098), .ZN(n2495) );
  NAND2_X1 U8197 ( .A1(n6069), .A2(n29610), .ZN(n6068) );
  NAND2_X1 U8199 ( .A1(n10682), .A2(n5265), .ZN(n11493) );
  OR2_X1 U8200 ( .A1(n20916), .A2(n18934), .ZN(n18933) );
  INV_X1 U8201 ( .A(n7770), .ZN(n7767) );
  AND2_X1 U8202 ( .A1(n14958), .A2(n15476), .ZN(n15169) );
  OR2_X1 U8205 ( .A1(n12228), .A2(n13081), .ZN(n11688) );
  INV_X1 U8206 ( .A(n18193), .ZN(n6663) );
  INV_X1 U8207 ( .A(n23433), .ZN(n5530) );
  INV_X1 U8208 ( .A(n1938), .ZN(n7964) );
  NOR2_X1 U8209 ( .A1(n14158), .A2(n14475), .ZN(n3867) );
  OAI211_X1 U8210 ( .C1(n27508), .C2(n27520), .A(n4165), .B(n4164), .ZN(n27519) );
  XNOR2_X1 U8211 ( .A(n10070), .B(n10069), .ZN(n10752) );
  AND2_X1 U8212 ( .A1(n28776), .A2(n17379), .ZN(n6501) );
  XNOR2_X1 U8213 ( .A(n4298), .B(n12559), .ZN(n12775) );
  XNOR2_X1 U8214 ( .A(n19500), .B(n1923), .ZN(n4221) );
  NAND2_X1 U8215 ( .A1(n11846), .A2(n11515), .ZN(n2319) );
  NAND2_X1 U8216 ( .A1(n8155), .A2(n7785), .ZN(n7171) );
  NAND2_X1 U8217 ( .A1(n7168), .A2(n7167), .ZN(n8155) );
  AND3_X2 U8218 ( .A1(n4398), .A2(n14011), .A3(n14012), .ZN(n14821) );
  NOR2_X1 U8219 ( .A1(n18261), .A2(n18326), .ZN(n17713) );
  INV_X1 U8220 ( .A(n2779), .ZN(n23470) );
  NOR2_X1 U8221 ( .A1(n2735), .A2(n20088), .ZN(n20040) );
  NAND2_X1 U8222 ( .A1(n2128), .A2(n8726), .ZN(n8852) );
  NAND2_X1 U8224 ( .A1(n28210), .A2(n9029), .ZN(n8795) );
  NAND2_X1 U8226 ( .A1(n2324), .A2(n2323), .ZN(n27304) );
  NAND2_X1 U8227 ( .A1(n26421), .A2(n28471), .ZN(n2324) );
  NAND3_X1 U8228 ( .A1(n11856), .A2(n12155), .A3(n12088), .ZN(n3008) );
  NAND2_X1 U8230 ( .A1(n29241), .A2(n8251), .ZN(n3224) );
  OR2_X1 U8231 ( .A1(n7890), .A2(n7891), .ZN(n7275) );
  NAND2_X1 U8232 ( .A1(n25406), .A2(n26191), .ZN(n25618) );
  OR2_X2 U8233 ( .A1(n11200), .A2(n5660), .ZN(n13118) );
  INV_X1 U8234 ( .A(Plaintext[156]), .ZN(n7046) );
  NAND3_X1 U8235 ( .A1(n23538), .A2(n23536), .A3(n23689), .ZN(n2326) );
  NAND2_X1 U8236 ( .A1(n5567), .A2(n9232), .ZN(n9049) );
  NAND2_X1 U8237 ( .A1(n15022), .A2(n15303), .ZN(n15025) );
  NAND2_X1 U8238 ( .A1(n13931), .A2(n2327), .ZN(n15303) );
  NAND2_X1 U8240 ( .A1(n18172), .A2(n18170), .ZN(n2329) );
  NAND2_X1 U8241 ( .A1(n17783), .A2(n18173), .ZN(n2330) );
  NAND2_X1 U8242 ( .A1(n5272), .A2(n5728), .ZN(n2332) );
  NAND2_X1 U8243 ( .A1(n5272), .A2(n24079), .ZN(n2333) );
  NAND2_X1 U8244 ( .A1(n4193), .A2(n21457), .ZN(n6803) );
  OR2_X1 U8245 ( .A1(n13646), .A2(n13816), .ZN(n5180) );
  XNOR2_X1 U8246 ( .A(n12069), .B(n12699), .ZN(n13438) );
  OR2_X1 U8247 ( .A1(n3936), .A2(n28580), .ZN(n3619) );
  NOR2_X1 U8248 ( .A1(n11449), .A2(n12328), .ZN(n12014) );
  INV_X1 U8249 ( .A(n13646), .ZN(n14299) );
  INV_X1 U8250 ( .A(n9913), .ZN(n11127) );
  XNOR2_X1 U8251 ( .A(n19520), .B(n18691), .ZN(n19066) );
  NAND3_X1 U8252 ( .A1(n10586), .A2(n12354), .A3(n11467), .ZN(n11469) );
  NAND2_X1 U8253 ( .A1(n5001), .A2(n17018), .ZN(n17254) );
  NAND2_X1 U8254 ( .A1(n7980), .A2(n7641), .ZN(n7193) );
  NAND2_X1 U8255 ( .A1(n29077), .A2(n10912), .ZN(n10688) );
  NAND3_X1 U8256 ( .A1(n21614), .A2(n28791), .A3(n2337), .ZN(n21616) );
  NAND2_X1 U8257 ( .A1(n21609), .A2(n2338), .ZN(n2337) );
  NAND3_X1 U8258 ( .A1(n6293), .A2(n15512), .A3(n15514), .ZN(n15517) );
  NAND2_X1 U8259 ( .A1(n4318), .A2(n2340), .ZN(n9823) );
  OAI21_X1 U8260 ( .B1(n10476), .B2(n11347), .A(n2342), .ZN(n11356) );
  NAND2_X1 U8261 ( .A1(n11347), .A2(n11350), .ZN(n2342) );
  NAND2_X1 U8263 ( .A1(n6210), .A2(n7507), .ZN(n2789) );
  NAND2_X1 U8265 ( .A1(n2345), .A2(n14400), .ZN(n2344) );
  INV_X1 U8266 ( .A(n13877), .ZN(n2345) );
  OR2_X1 U8267 ( .A1(n14398), .A2(n14400), .ZN(n2346) );
  NAND2_X1 U8268 ( .A1(n15514), .A2(n14697), .ZN(n2347) );
  XNOR2_X1 U8270 ( .A(n15642), .B(n16421), .ZN(n15644) );
  NAND2_X2 U8271 ( .A1(n4708), .A2(n14699), .ZN(n16421) );
  NAND2_X1 U8272 ( .A1(n11880), .A2(n11881), .ZN(n2348) );
  NAND2_X1 U8273 ( .A1(n11879), .A2(n287), .ZN(n2349) );
  NAND2_X1 U8274 ( .A1(n21661), .A2(n20833), .ZN(n21073) );
  NAND2_X1 U8275 ( .A1(n7746), .A2(n7533), .ZN(n7143) );
  NAND2_X1 U8277 ( .A1(n2614), .A2(n10712), .ZN(n11774) );
  NAND3_X1 U8278 ( .A1(n6738), .A2(n27427), .A3(n29542), .ZN(n26968) );
  NAND2_X1 U8279 ( .A1(n17116), .A2(n29539), .ZN(n3100) );
  OAI211_X2 U8280 ( .C1(n24045), .C2(n24044), .A(n2828), .B(n2829), .ZN(n26053) );
  NAND2_X1 U8281 ( .A1(n5888), .A2(n2352), .ZN(n9226) );
  NAND3_X1 U8283 ( .A1(n2794), .A2(n27746), .A3(n2795), .ZN(n2793) );
  NAND2_X1 U8287 ( .A1(n15315), .A2(n15319), .ZN(n15316) );
  MUX2_X1 U8288 ( .A(n18337), .B(n18331), .S(n18332), .Z(n17651) );
  NAND3_X1 U8292 ( .A1(n11196), .A2(n10751), .A3(n28207), .ZN(n2431) );
  AOI21_X1 U8294 ( .B1(n14924), .B2(n14923), .A(n15497), .ZN(n14925) );
  NAND2_X1 U8296 ( .A1(n10646), .A2(n12027), .ZN(n10647) );
  NAND3_X1 U8299 ( .A1(n1931), .A2(n12162), .A3(n2357), .ZN(n11380) );
  INV_X1 U8300 ( .A(n12103), .ZN(n2357) );
  XOR2_X1 U8301 ( .A(n19699), .B(n19698), .Z(n5006) );
  OR2_X1 U8302 ( .A1(n17269), .A2(n29299), .ZN(n3038) );
  OAI22_X1 U8303 ( .A1(n6034), .A2(n23686), .B1(n23168), .B2(n23679), .ZN(
        n23134) );
  NAND3_X2 U8304 ( .A1(n2359), .A2(n2780), .A3(n2358), .ZN(n9184) );
  NAND2_X1 U8305 ( .A1(n2781), .A2(n7141), .ZN(n2359) );
  NAND3_X1 U8306 ( .A1(n11790), .A2(n11791), .A3(n2360), .ZN(n11792) );
  NAND2_X1 U8307 ( .A1(n2361), .A2(n26729), .ZN(n25628) );
  OAI21_X1 U8308 ( .B1(n2361), .B2(n26729), .A(n26728), .ZN(n26730) );
  INV_X1 U8309 ( .A(n26481), .ZN(n2361) );
  MUX2_X1 U8310 ( .A(n10912), .B(n29078), .S(n10911), .Z(n10917) );
  OAI21_X1 U8311 ( .B1(n10689), .B2(n10911), .A(n29078), .ZN(n10690) );
  AOI21_X1 U8312 ( .B1(n10914), .B2(n10605), .A(n29077), .ZN(n10452) );
  NAND2_X1 U8313 ( .A1(n10915), .A2(n29077), .ZN(n10606) );
  AND2_X1 U8315 ( .A1(n2363), .A2(n18215), .ZN(n18502) );
  INV_X1 U8316 ( .A(n18216), .ZN(n2363) );
  NAND2_X1 U8317 ( .A1(n5692), .A2(n2364), .ZN(n5691) );
  INV_X1 U8318 ( .A(n18215), .ZN(n2364) );
  NAND2_X1 U8319 ( .A1(n5154), .A2(n2365), .ZN(n17727) );
  NAND2_X1 U8320 ( .A1(n5690), .A2(n18215), .ZN(n2365) );
  NAND2_X1 U8321 ( .A1(n14634), .A2(n14635), .ZN(n16567) );
  OR2_X2 U8322 ( .A1(n13845), .A2(n13846), .ZN(n15738) );
  INV_X1 U8324 ( .A(n10985), .ZN(n3802) );
  AOI22_X2 U8325 ( .A1(n23933), .A2(n24291), .B1(n23934), .B2(n24730), .ZN(
        n25808) );
  XNOR2_X1 U8327 ( .A(n12753), .B(n13136), .ZN(n13328) );
  NAND3_X1 U8328 ( .A1(n5659), .A2(n514), .A3(n17906), .ZN(n4076) );
  NAND2_X1 U8329 ( .A1(n2366), .A2(n23830), .ZN(n24095) );
  NAND2_X1 U8330 ( .A1(n481), .A2(n23833), .ZN(n23830) );
  INV_X1 U8331 ( .A(n2367), .ZN(n2366) );
  NAND3_X1 U8332 ( .A1(n2368), .A2(n8977), .A3(n8818), .ZN(n8822) );
  NAND2_X1 U8333 ( .A1(n8974), .A2(n8817), .ZN(n2368) );
  XNOR2_X1 U8334 ( .A(n9977), .B(n2034), .ZN(n6916) );
  NAND2_X1 U8335 ( .A1(n2369), .A2(n4554), .ZN(n10102) );
  NAND2_X1 U8336 ( .A1(n4553), .A2(n4555), .ZN(n2369) );
  NAND2_X1 U8337 ( .A1(n20579), .A2(n20417), .ZN(n2371) );
  NAND2_X1 U8338 ( .A1(n20578), .A2(n20577), .ZN(n2372) );
  OAI22_X1 U8340 ( .A1(n5064), .A2(n6011), .B1(n13909), .B2(n14043), .ZN(n2373) );
  XNOR2_X2 U8341 ( .A(n2374), .B(Key[108]), .ZN(n8217) );
  INV_X1 U8342 ( .A(Plaintext[108]), .ZN(n2374) );
  NAND2_X1 U8344 ( .A1(n2377), .A2(n2376), .ZN(n26873) );
  OAI21_X1 U8345 ( .B1(n3236), .B2(n26902), .A(n2378), .ZN(n2377) );
  NOR2_X2 U8346 ( .A1(n24069), .A2(n2379), .ZN(n25809) );
  OAI211_X1 U8347 ( .C1(n27478), .C2(n27492), .A(n2380), .B(n5606), .ZN(n26704) );
  NAND2_X1 U8348 ( .A1(n2882), .A2(n2883), .ZN(n2382) );
  NAND2_X1 U8352 ( .A1(n3005), .A2(n20481), .ZN(n2383) );
  NAND2_X1 U8354 ( .A1(n5147), .A2(n7604), .ZN(n8735) );
  XNOR2_X1 U8355 ( .A(n2384), .B(n9932), .ZN(n4600) );
  XNOR2_X1 U8356 ( .A(n9928), .B(n9929), .ZN(n2384) );
  AND2_X1 U8357 ( .A1(n14336), .A2(n14408), .ZN(n13813) );
  OR2_X1 U8358 ( .A1(n17304), .A2(n5714), .ZN(n16788) );
  OR2_X1 U8359 ( .A1(n18456), .A2(n4230), .ZN(n16793) );
  INV_X1 U8360 ( .A(n20090), .ZN(n20091) );
  NAND2_X1 U8361 ( .A1(n2386), .A2(n1568), .ZN(n4695) );
  OAI21_X1 U8362 ( .B1(n4696), .B2(n29301), .A(n3642), .ZN(n2386) );
  OAI21_X1 U8363 ( .B1(n12232), .B2(n776), .A(n2412), .ZN(n12039) );
  INV_X1 U8365 ( .A(Plaintext[164]), .ZN(n2387) );
  NAND2_X1 U8366 ( .A1(n2917), .A2(n3331), .ZN(n2388) );
  NAND2_X1 U8368 ( .A1(n6843), .A2(n20133), .ZN(n2390) );
  NAND2_X1 U8369 ( .A1(n2391), .A2(n8168), .ZN(n2942) );
  NAND2_X1 U8370 ( .A1(n7536), .A2(n7352), .ZN(n2391) );
  XNOR2_X1 U8372 ( .A(n2392), .B(n3633), .ZN(Ciphertext[76]) );
  NOR2_X1 U8373 ( .A1(n27206), .A2(n27207), .ZN(n2392) );
  OR2_X1 U8374 ( .A1(n14197), .A2(n28199), .ZN(n14198) );
  XNOR2_X1 U8377 ( .A(n22275), .B(n22485), .ZN(n2393) );
  XNOR2_X1 U8378 ( .A(n2394), .B(n22170), .ZN(n22173) );
  XNOR2_X1 U8379 ( .A(n22171), .B(n28387), .ZN(n2394) );
  NAND2_X1 U8380 ( .A1(n21394), .A2(n2395), .ZN(n2409) );
  NAND2_X1 U8382 ( .A1(n2918), .A2(n20863), .ZN(n2396) );
  NAND3_X2 U8384 ( .A1(n2397), .A2(n3487), .A3(n13518), .ZN(n16312) );
  NAND2_X1 U8385 ( .A1(n6668), .A2(n14884), .ZN(n2397) );
  NAND3_X1 U8386 ( .A1(n15717), .A2(n17366), .A3(n15731), .ZN(n15733) );
  NOR2_X1 U8387 ( .A1(n8301), .A2(n7400), .ZN(n3203) );
  NAND2_X1 U8388 ( .A1(n11908), .A2(n12363), .ZN(n11446) );
  NAND2_X1 U8389 ( .A1(n14231), .A2(n14230), .ZN(n3645) );
  OR2_X1 U8390 ( .A1(n17374), .A2(n17379), .ZN(n4651) );
  NAND2_X1 U8391 ( .A1(n21328), .A2(n21330), .ZN(n21163) );
  NOR2_X1 U8392 ( .A1(n29526), .A2(n21373), .ZN(n21273) );
  NAND2_X1 U8393 ( .A1(n2399), .A2(n2398), .ZN(n3058) );
  AOI21_X1 U8394 ( .B1(n349), .B2(n12072), .A(n12251), .ZN(n2398) );
  NAND2_X1 U8395 ( .A1(n11933), .A2(n12249), .ZN(n2399) );
  OAI21_X1 U8396 ( .B1(n23417), .B2(n485), .A(n2400), .ZN(n23420) );
  XNOR2_X1 U8397 ( .A(n9811), .B(n2401), .ZN(n9813) );
  XNOR2_X1 U8398 ( .A(n9810), .B(n10071), .ZN(n2401) );
  INV_X1 U8400 ( .A(Plaintext[168]), .ZN(n6208) );
  INV_X1 U8401 ( .A(n18762), .ZN(n3913) );
  NAND3_X1 U8402 ( .A1(n9436), .A2(n9211), .A3(n9209), .ZN(n7682) );
  AOI21_X1 U8406 ( .B1(n2898), .B2(n8291), .A(n8287), .ZN(n2406) );
  OAI21_X1 U8407 ( .B1(n27791), .B2(n2407), .A(n27800), .ZN(n27792) );
  NOR2_X1 U8408 ( .A1(n27790), .A2(n27819), .ZN(n2407) );
  NAND2_X1 U8409 ( .A1(n17763), .A2(n17873), .ZN(n17764) );
  NAND2_X1 U8410 ( .A1(n19833), .A2(n20382), .ZN(n5943) );
  NAND2_X1 U8412 ( .A1(n11235), .A2(n11013), .ZN(n11016) );
  AOI21_X1 U8413 ( .B1(n3464), .B2(n7238), .A(n7885), .ZN(n5174) );
  INV_X1 U8414 ( .A(n8801), .ZN(n9160) );
  OAI21_X1 U8415 ( .B1(n2945), .B2(n13747), .A(n13763), .ZN(n2408) );
  OR2_X1 U8416 ( .A1(n9124), .A2(n284), .ZN(n4060) );
  NOR2_X1 U8417 ( .A1(n10706), .A2(n10942), .ZN(n10447) );
  INV_X1 U8418 ( .A(n8136), .ZN(n7127) );
  INV_X1 U8419 ( .A(n23448), .ZN(n4794) );
  INV_X1 U8420 ( .A(n14259), .ZN(n2681) );
  INV_X1 U8421 ( .A(n14981), .ZN(n5635) );
  NAND2_X1 U8422 ( .A1(n21398), .A2(n2409), .ZN(n22158) );
  XNOR2_X2 U8423 ( .A(n7108), .B(Key[188]), .ZN(n7900) );
  NAND2_X1 U8424 ( .A1(n7800), .A2(n7801), .ZN(n7802) );
  NAND2_X1 U8425 ( .A1(n7127), .A2(n29646), .ZN(n8052) );
  NAND2_X1 U8426 ( .A1(n14262), .A2(n14260), .ZN(n14098) );
  NAND2_X1 U8428 ( .A1(n23376), .A2(n23377), .ZN(n23381) );
  NAND2_X1 U8430 ( .A1(n23497), .A2(n23493), .ZN(n23796) );
  NAND3_X1 U8432 ( .A1(n8830), .A2(n1839), .A3(n8829), .ZN(n2410) );
  NOR2_X1 U8433 ( .A1(n18286), .A2(n18524), .ZN(n18082) );
  AND2_X2 U8434 ( .A1(n4427), .A2(n4428), .ZN(n17719) );
  INV_X1 U8435 ( .A(n2413), .ZN(n10629) );
  NAND2_X1 U8436 ( .A1(n12232), .A2(n12234), .ZN(n2412) );
  NAND2_X1 U8437 ( .A1(n14702), .A2(n14916), .ZN(n15495) );
  NAND2_X1 U8438 ( .A1(n27631), .A2(n27630), .ZN(n2415) );
  INV_X1 U8439 ( .A(n17415), .ZN(n15811) );
  NAND2_X1 U8440 ( .A1(n2417), .A2(n17415), .ZN(n2416) );
  INV_X1 U8441 ( .A(n17413), .ZN(n2417) );
  NAND2_X1 U8442 ( .A1(n2419), .A2(n9188), .ZN(n2418) );
  NAND2_X1 U8443 ( .A1(n9187), .A2(n9186), .ZN(n2419) );
  NAND2_X1 U8444 ( .A1(n9189), .A2(n8445), .ZN(n2420) );
  NAND2_X1 U8447 ( .A1(n10697), .A2(n10989), .ZN(n2423) );
  NAND2_X1 U8449 ( .A1(n4577), .A2(n7579), .ZN(n2424) );
  NAND2_X1 U8450 ( .A1(n3379), .A2(n14141), .ZN(n13717) );
  NOR2_X1 U8452 ( .A1(n8956), .A2(n8954), .ZN(n2425) );
  INV_X1 U8453 ( .A(n21364), .ZN(n5772) );
  XOR2_X1 U8454 ( .A(n13398), .B(n13397), .Z(n2875) );
  OAI21_X1 U8455 ( .B1(n27359), .B2(n27360), .A(n2426), .ZN(n27361) );
  NAND2_X1 U8456 ( .A1(n6766), .A2(n6767), .ZN(n6769) );
  NAND2_X1 U8457 ( .A1(n20853), .A2(n2427), .ZN(n20855) );
  NAND3_X1 U8460 ( .A1(n4560), .A2(n4562), .A3(n2036), .ZN(n24138) );
  NOR2_X1 U8461 ( .A1(n27230), .A2(n2428), .ZN(n27232) );
  OAI22_X1 U8462 ( .A1(n27229), .A2(n27757), .B1(n27228), .B2(n29049), .ZN(
        n2428) );
  OAI211_X2 U8463 ( .C1(n9194), .C2(n7639), .A(n7638), .B(n2429), .ZN(n9772)
         );
  NAND2_X1 U8464 ( .A1(n6897), .A2(n9202), .ZN(n2429) );
  NAND2_X1 U8466 ( .A1(n10869), .A2(n11453), .ZN(n2430) );
  NAND2_X1 U8467 ( .A1(n11595), .A2(n12251), .ZN(n2710) );
  XNOR2_X2 U8468 ( .A(n9432), .B(n5895), .ZN(n10936) );
  OR2_X1 U8469 ( .A1(n8762), .A2(n8553), .ZN(n8557) );
  NAND3_X1 U8472 ( .A1(n8488), .A2(n8899), .A3(n1793), .ZN(n6317) );
  NAND2_X1 U8474 ( .A1(n4941), .A2(n3148), .ZN(n8132) );
  NAND2_X1 U8476 ( .A1(n27217), .A2(n2433), .ZN(n2432) );
  INV_X1 U8477 ( .A(n27562), .ZN(n2433) );
  NAND2_X1 U8478 ( .A1(n27216), .A2(n27562), .ZN(n2434) );
  INV_X1 U8483 ( .A(n27277), .ZN(n2438) );
  NAND2_X1 U8484 ( .A1(n27290), .A2(n27286), .ZN(n2439) );
  INV_X1 U8485 ( .A(n21292), .ZN(n20985) );
  OR2_X1 U8486 ( .A1(n28626), .A2(n23099), .ZN(n2451) );
  NAND2_X1 U8489 ( .A1(n2442), .A2(n464), .ZN(n3713) );
  INV_X1 U8490 ( .A(n9116), .ZN(n8071) );
  NAND2_X1 U8492 ( .A1(n17796), .A2(n2445), .ZN(n2444) );
  INV_X1 U8493 ( .A(n18087), .ZN(n2445) );
  NAND2_X1 U8494 ( .A1(n13678), .A2(n12743), .ZN(n14182) );
  NAND2_X1 U8495 ( .A1(n4261), .A2(n1993), .ZN(n13133) );
  NAND2_X1 U8496 ( .A1(n13852), .A2(n13933), .ZN(n14187) );
  NAND2_X1 U8499 ( .A1(n15381), .A2(n15384), .ZN(n2448) );
  NAND2_X1 U8500 ( .A1(n4283), .A2(n17357), .ZN(n2450) );
  XOR2_X1 U8502 ( .A(n13482), .B(n27515), .Z(n6652) );
  NAND2_X1 U8503 ( .A1(n11072), .A2(n11075), .ZN(n10891) );
  NAND2_X1 U8504 ( .A1(n5352), .A2(n13827), .ZN(n5351) );
  OAI211_X1 U8505 ( .C1(n25954), .C2(n27317), .A(n2454), .B(n2453), .ZN(n25955) );
  NAND2_X1 U8506 ( .A1(n26594), .A2(n27317), .ZN(n2453) );
  NAND2_X1 U8507 ( .A1(n25897), .A2(n27873), .ZN(n2454) );
  INV_X1 U8508 ( .A(n10008), .ZN(n3073) );
  OR2_X1 U8509 ( .A1(n5775), .A2(n22284), .ZN(n23040) );
  XNOR2_X1 U8510 ( .A(n10138), .B(n9735), .ZN(n9918) );
  NAND2_X1 U8511 ( .A1(n15294), .A2(n2455), .ZN(n14836) );
  XNOR2_X1 U8512 ( .A(n6665), .B(n6666), .ZN(n10875) );
  XNOR2_X1 U8515 ( .A(n22439), .B(n22440), .ZN(n2779) );
  NAND2_X1 U8517 ( .A1(n2458), .A2(n3831), .ZN(n19277) );
  NAND3_X1 U8518 ( .A1(n17714), .A2(n3832), .A3(n18323), .ZN(n2458) );
  NAND2_X1 U8520 ( .A1(n11414), .A2(n11415), .ZN(n11418) );
  NAND3_X1 U8521 ( .A1(n7952), .A2(n28614), .A3(n2461), .ZN(n7951) );
  NAND2_X1 U8522 ( .A1(n7946), .A2(n7947), .ZN(n2461) );
  OAI21_X1 U8524 ( .B1(n14281), .B2(n14285), .A(n2462), .ZN(n13621) );
  NAND2_X1 U8525 ( .A1(n14285), .A2(n14287), .ZN(n2462) );
  NAND4_X2 U8526 ( .A1(n11624), .A2(n11625), .A3(n11627), .A4(n11626), .ZN(
        n13567) );
  OAI21_X1 U8527 ( .B1(n6386), .B2(n6385), .A(n10888), .ZN(n10889) );
  AND2_X2 U8530 ( .A1(n3304), .A2(n3305), .ZN(n22139) );
  XNOR2_X2 U8531 ( .A(n7166), .B(Key[20]), .ZN(n7291) );
  NAND3_X1 U8532 ( .A1(n5659), .A2(n17906), .A3(n17663), .ZN(n5701) );
  NAND2_X1 U8533 ( .A1(n28105), .A2(n29056), .ZN(n2463) );
  OAI21_X2 U8534 ( .B1(n17495), .B2(n16733), .A(n16732), .ZN(n18203) );
  OAI21_X1 U8535 ( .B1(n7954), .B2(n8670), .A(n7953), .ZN(n7955) );
  XOR2_X1 U8536 ( .A(n9672), .B(n9671), .Z(n4601) );
  NAND2_X1 U8537 ( .A1(n12265), .A2(n2466), .ZN(n11060) );
  OAI22_X1 U8539 ( .A1(n14119), .A2(n14369), .B1(n14093), .B2(n564), .ZN(
        n13835) );
  NAND2_X1 U8540 ( .A1(n559), .A2(n14366), .ZN(n14119) );
  NAND2_X1 U8542 ( .A1(n11688), .A2(n11689), .ZN(n11691) );
  OAI21_X1 U8543 ( .B1(n612), .B2(n7981), .A(n7642), .ZN(n7454) );
  NAND2_X1 U8545 ( .A1(n8724), .A2(n8605), .ZN(n2890) );
  XNOR2_X1 U8546 ( .A(n19412), .B(n18857), .ZN(n19097) );
  NAND2_X1 U8547 ( .A1(n17167), .A2(n2468), .ZN(n19412) );
  NAND2_X1 U8548 ( .A1(n9221), .A2(n8525), .ZN(n9224) );
  NAND4_X2 U8549 ( .A1(n6330), .A2(n6329), .A3(n6328), .A4(n10465), .ZN(n13097) );
  AOI21_X1 U8551 ( .B1(n8893), .B2(n8892), .A(n8891), .ZN(n8894) );
  NAND2_X1 U8552 ( .A1(n8504), .A2(n8009), .ZN(n8892) );
  NOR2_X1 U8553 ( .A1(n2469), .A2(n2016), .ZN(n23008) );
  OAI21_X1 U8554 ( .B1(n21896), .B2(n23663), .A(n23522), .ZN(n2469) );
  NAND3_X1 U8555 ( .A1(n3157), .A2(n3156), .A3(n9529), .ZN(n9536) );
  NAND3_X1 U8557 ( .A1(n7990), .A2(n2472), .A3(n2471), .ZN(n2470) );
  NAND2_X1 U8558 ( .A1(n29639), .A2(n341), .ZN(n2471) );
  NAND3_X1 U8559 ( .A1(n4647), .A2(n4646), .A3(n6206), .ZN(n22227) );
  NAND2_X1 U8560 ( .A1(n6526), .A2(n6927), .ZN(n2935) );
  OAI21_X1 U8562 ( .B1(n24496), .B2(n24497), .A(n24810), .ZN(n2473) );
  OR2_X1 U8563 ( .A1(n14491), .A2(n14498), .ZN(n2964) );
  NAND2_X1 U8564 ( .A1(n28651), .A2(n28467), .ZN(n25035) );
  INV_X1 U8565 ( .A(n20597), .ZN(n20603) );
  XNOR2_X1 U8566 ( .A(n12872), .B(n4375), .ZN(n12652) );
  OR2_X2 U8567 ( .A1(n5031), .A2(n3405), .ZN(n4364) );
  OR2_X1 U8568 ( .A1(n26679), .A2(n27821), .ZN(n3561) );
  OR2_X1 U8569 ( .A1(n14451), .A2(n13753), .ZN(n2970) );
  AND2_X1 U8570 ( .A1(n23599), .A2(n23467), .ZN(n24257) );
  NOR2_X1 U8571 ( .A1(n24257), .A2(n5548), .ZN(n2806) );
  INV_X1 U8572 ( .A(n15290), .ZN(n15294) );
  INV_X1 U8573 ( .A(n6080), .ZN(n6449) );
  AND2_X1 U8574 ( .A1(n3227), .A2(n21626), .ZN(n5338) );
  OR2_X1 U8576 ( .A1(n15027), .A2(n15431), .ZN(n15029) );
  INV_X1 U8577 ( .A(n18646), .ZN(n19668) );
  OR2_X1 U8579 ( .A1(n7786), .A2(n7787), .ZN(n7167) );
  INV_X1 U8580 ( .A(n18231), .ZN(n18400) );
  AND2_X1 U8581 ( .A1(n21625), .A2(n22141), .ZN(n2911) );
  OAI22_X1 U8582 ( .A1(n3992), .A2(n10031), .B1(n10718), .B2(n11137), .ZN(
        n3991) );
  XNOR2_X1 U8583 ( .A(n25836), .B(n25903), .ZN(n25207) );
  XNOR2_X1 U8584 ( .A(n25207), .B(n26038), .ZN(n25502) );
  OR2_X1 U8585 ( .A1(n15101), .A2(n15103), .ZN(n2576) );
  INV_X1 U8586 ( .A(n14893), .ZN(n15107) );
  INV_X1 U8588 ( .A(n22992), .ZN(n23643) );
  OAI21_X1 U8589 ( .B1(n2020), .B2(n14344), .A(n14341), .ZN(n6234) );
  NAND3_X2 U8590 ( .A1(n17329), .A2(n17330), .A3(n2720), .ZN(n19136) );
  NAND2_X1 U8591 ( .A1(n2475), .A2(n2474), .ZN(n27639) );
  OR2_X1 U8592 ( .A1(n26357), .A2(n28651), .ZN(n2474) );
  NAND3_X1 U8593 ( .A1(n25043), .A2(n26270), .A3(n25042), .ZN(n2475) );
  INV_X1 U8594 ( .A(n29565), .ZN(n14486) );
  INV_X1 U8595 ( .A(n17570), .ZN(n17573) );
  XNOR2_X1 U8596 ( .A(n429), .B(n13414), .ZN(n12087) );
  AOI22_X1 U8599 ( .A1(n28422), .A2(n27537), .B1(n28468), .B2(n27547), .ZN(
        n27543) );
  NOR2_X1 U8600 ( .A1(n24420), .A2(n24517), .ZN(n24513) );
  XNOR2_X1 U8601 ( .A(n19634), .B(n19599), .ZN(n6487) );
  NAND3_X1 U8602 ( .A1(n4332), .A2(n17560), .A3(n2061), .ZN(n5428) );
  NAND2_X1 U8607 ( .A1(n4774), .A2(n17980), .ZN(n17981) );
  NAND2_X1 U8611 ( .A1(n7421), .A2(n7420), .ZN(n2480) );
  NAND2_X1 U8612 ( .A1(n2482), .A2(n2481), .ZN(n23745) );
  NAND2_X1 U8614 ( .A1(n23737), .A2(n23228), .ZN(n2482) );
  OAI21_X1 U8615 ( .B1(n13410), .B2(n2874), .A(n2873), .ZN(n13411) );
  NAND2_X1 U8618 ( .A1(n20458), .A2(n4569), .ZN(n20600) );
  OAI211_X1 U8620 ( .C1(n14498), .C2(n14493), .A(n2488), .B(n13672), .ZN(
        n12804) );
  NAND2_X1 U8621 ( .A1(n2489), .A2(n17089), .ZN(n18695) );
  OAI21_X1 U8622 ( .B1(n17082), .B2(n18596), .A(n5476), .ZN(n2489) );
  XNOR2_X1 U8623 ( .A(n19101), .B(n2490), .ZN(n19006) );
  XNOR2_X1 U8624 ( .A(n19004), .B(n19003), .ZN(n2490) );
  AOI21_X1 U8625 ( .B1(n7407), .B2(n7408), .A(n7480), .ZN(n2491) );
  NAND2_X1 U8627 ( .A1(n5693), .A2(n14178), .ZN(n2493) );
  NOR2_X1 U8629 ( .A1(n14006), .A2(n14386), .ZN(n13573) );
  NAND2_X1 U8630 ( .A1(n13572), .A2(n14380), .ZN(n14006) );
  XNOR2_X1 U8633 ( .A(n15966), .B(n15989), .ZN(n15042) );
  OAI211_X1 U8634 ( .C1(n23636), .C2(n23557), .A(n2494), .B(n23556), .ZN(
        n23561) );
  NOR2_X1 U8635 ( .A1(n23555), .A2(n23554), .ZN(n2494) );
  NAND2_X1 U8636 ( .A1(n184), .A2(n15094), .ZN(n2496) );
  NAND2_X1 U8638 ( .A1(n2500), .A2(n2499), .ZN(n2498) );
  OR2_X1 U8639 ( .A1(n5837), .A2(n11955), .ZN(n12258) );
  NAND2_X1 U8641 ( .A1(n7619), .A2(n8232), .ZN(n7620) );
  NAND2_X1 U8644 ( .A1(n2504), .A2(n2503), .ZN(n11900) );
  NAND2_X1 U8645 ( .A1(n11898), .A2(n29461), .ZN(n2503) );
  NAND2_X1 U8646 ( .A1(n11897), .A2(n11896), .ZN(n2504) );
  OR2_X1 U8650 ( .A1(n18215), .A2(n5155), .ZN(n5154) );
  INV_X1 U8651 ( .A(n7554), .ZN(n8133) );
  INV_X1 U8652 ( .A(n10937), .ZN(n10999) );
  XNOR2_X1 U8653 ( .A(n5412), .B(n10392), .ZN(n5411) );
  AND3_X2 U8654 ( .A1(n2071), .A2(n2564), .A3(n2565), .ZN(n9062) );
  OR2_X1 U8655 ( .A1(n7079), .A2(n7092), .ZN(n2507) );
  XNOR2_X1 U8656 ( .A(n15536), .B(n16201), .ZN(n15540) );
  NAND2_X1 U8659 ( .A1(n23529), .A2(n23531), .ZN(n23135) );
  NAND2_X1 U8660 ( .A1(n18235), .A2(n17977), .ZN(n2508) );
  NAND2_X1 U8662 ( .A1(n7634), .A2(n7828), .ZN(n7832) );
  XNOR2_X1 U8664 ( .A(n15761), .B(n4767), .ZN(n4766) );
  NAND2_X1 U8666 ( .A1(n16946), .A2(n16945), .ZN(n6176) );
  OR2_X1 U8667 ( .A1(n11449), .A2(n11747), .ZN(n11450) );
  NOR2_X1 U8670 ( .A1(n18053), .A2(n18054), .ZN(n18055) );
  NAND2_X1 U8671 ( .A1(n4680), .A2(n16667), .ZN(n16685) );
  BUF_X1 U8672 ( .A(n16764), .Z(n17002) );
  NAND2_X1 U8673 ( .A1(n7194), .A2(n7985), .ZN(n2514) );
  NAND2_X1 U8674 ( .A1(n7193), .A2(n7644), .ZN(n2516) );
  NAND3_X1 U8676 ( .A1(n20710), .A2(n20816), .A3(n21268), .ZN(n6426) );
  NAND2_X1 U8677 ( .A1(n11492), .A2(n4404), .ZN(n11497) );
  NOR2_X1 U8680 ( .A1(n11086), .A2(n28624), .ZN(n2518) );
  INV_X1 U8681 ( .A(n19891), .ZN(n3421) );
  NAND2_X1 U8682 ( .A1(n8133), .A2(n8047), .ZN(n7718) );
  NAND2_X1 U8683 ( .A1(n2519), .A2(n20718), .ZN(n22759) );
  NAND2_X1 U8684 ( .A1(n5206), .A2(n5205), .ZN(n2519) );
  NAND2_X1 U8685 ( .A1(n20514), .A2(n20513), .ZN(n19241) );
  NAND2_X1 U8686 ( .A1(n20343), .A2(n20342), .ZN(n20514) );
  NAND2_X1 U8687 ( .A1(n2521), .A2(n2520), .ZN(n11632) );
  NAND2_X1 U8688 ( .A1(n10757), .A2(n11345), .ZN(n2520) );
  NAND2_X1 U8689 ( .A1(n1926), .A2(n15320), .ZN(n3627) );
  INV_X1 U8690 ( .A(n27248), .ZN(n5335) );
  OAI211_X2 U8691 ( .C1(n27167), .C2(n26369), .A(n2525), .B(n2524), .ZN(n27625) );
  NAND2_X1 U8692 ( .A1(n27171), .A2(n27169), .ZN(n2524) );
  NAND2_X1 U8693 ( .A1(n26368), .A2(n29487), .ZN(n2525) );
  INV_X1 U8694 ( .A(n13260), .ZN(n13485) );
  OR2_X1 U8695 ( .A1(n26819), .A2(n6568), .ZN(n4926) );
  NOR2_X1 U8696 ( .A1(n26447), .A2(n26449), .ZN(n4832) );
  OAI22_X1 U8698 ( .A1(n2526), .A2(n24220), .B1(n24219), .B2(n23956), .ZN(
        n24221) );
  NAND2_X1 U8699 ( .A1(n28509), .A2(n24760), .ZN(n2526) );
  NOR2_X1 U8700 ( .A1(n7708), .A2(n7382), .ZN(n2897) );
  XNOR2_X1 U8701 ( .A(n6569), .B(n19387), .ZN(n20248) );
  AOI21_X1 U8702 ( .B1(n3504), .B2(n3503), .A(n20636), .ZN(n2529) );
  NAND2_X1 U8703 ( .A1(n15119), .A2(n14743), .ZN(n13660) );
  NAND2_X1 U8704 ( .A1(n4179), .A2(n7497), .ZN(n7499) );
  NAND2_X1 U8705 ( .A1(n2718), .A2(n18405), .ZN(n5022) );
  NAND4_X2 U8706 ( .A1(n24763), .A2(n24762), .A3(n2531), .A4(n2530), .ZN(
        n25810) );
  NAND2_X1 U8707 ( .A1(n2866), .A2(n378), .ZN(n2530) );
  NAND2_X1 U8708 ( .A1(n2865), .A2(n23588), .ZN(n2531) );
  XNOR2_X1 U8709 ( .A(n22388), .B(n22523), .ZN(n2532) );
  OAI211_X1 U8711 ( .C1(n27199), .C2(n27198), .A(n3899), .B(n2618), .ZN(n3898)
         );
  NAND2_X1 U8712 ( .A1(n18009), .A2(n2533), .ZN(n18762) );
  OR2_X1 U8713 ( .A1(n18010), .A2(n6079), .ZN(n2533) );
  XNOR2_X2 U8715 ( .A(n13529), .B(n13528), .ZN(n14007) );
  OAI22_X1 U8718 ( .A1(n19752), .A2(n20083), .B1(n5126), .B2(n18837), .ZN(
        n2534) );
  NAND2_X1 U8721 ( .A1(n12180), .A2(n12181), .ZN(n11411) );
  NAND2_X1 U8722 ( .A1(n24416), .A2(n24709), .ZN(n6513) );
  OAI21_X1 U8723 ( .B1(n24707), .B2(n24417), .A(n5795), .ZN(n24416) );
  NAND3_X1 U8724 ( .A1(n27825), .A2(n27101), .A3(n26901), .ZN(n26875) );
  XNOR2_X1 U8725 ( .A(n10328), .B(n10184), .ZN(n10185) );
  AOI21_X1 U8727 ( .B1(n8180), .B2(n8181), .A(n4856), .ZN(n8182) );
  OAI21_X2 U8728 ( .B1(n7647), .B2(n7648), .A(n7646), .ZN(n9211) );
  NAND2_X1 U8729 ( .A1(n11584), .A2(n567), .ZN(n11587) );
  NAND2_X1 U8730 ( .A1(n8028), .A2(n8032), .ZN(n7736) );
  OAI211_X1 U8734 ( .C1(n10499), .C2(n1834), .A(n10715), .B(n2539), .ZN(n10455) );
  NAND2_X1 U8735 ( .A1(n5672), .A2(n10498), .ZN(n2539) );
  INV_X1 U8736 ( .A(n10022), .ZN(n3452) );
  AOI21_X1 U8737 ( .B1(n11456), .B2(n11455), .A(n2542), .ZN(n13017) );
  OAI21_X1 U8738 ( .B1(n8829), .B2(n8826), .A(n8462), .ZN(n3706) );
  NAND2_X1 U8739 ( .A1(n8192), .A2(n4675), .ZN(n8462) );
  XNOR2_X1 U8745 ( .A(n18166), .B(n18167), .ZN(n19820) );
  OR2_X1 U8746 ( .A1(n13639), .A2(n14944), .ZN(n13586) );
  XNOR2_X1 U8747 ( .A(n3403), .B(n18913), .ZN(n19604) );
  NOR2_X1 U8748 ( .A1(n18214), .A2(n4824), .ZN(n18218) );
  OAI21_X1 U8750 ( .B1(n2546), .B2(n8147), .A(n2545), .ZN(n7151) );
  OR2_X1 U8751 ( .A1(n17439), .A2(n336), .ZN(n16926) );
  NAND3_X2 U8752 ( .A1(n3140), .A2(n8184), .A3(n3139), .ZN(n10321) );
  XNOR2_X2 U8753 ( .A(n8318), .B(n8319), .ZN(n11168) );
  NAND2_X1 U8754 ( .A1(n7928), .A2(n7927), .ZN(n2547) );
  OAI21_X1 U8755 ( .B1(n14064), .B2(n14065), .A(n3393), .ZN(n13164) );
  XOR2_X1 U8756 ( .A(n16444), .B(n16519), .Z(n5858) );
  AOI21_X2 U8757 ( .B1(n18419), .B2(n18418), .A(n18417), .ZN(n19206) );
  XNOR2_X1 U8759 ( .A(n2551), .B(n21766), .ZN(n21768) );
  XNOR2_X1 U8760 ( .A(n21765), .B(n22757), .ZN(n2551) );
  NAND2_X1 U8761 ( .A1(n27021), .A2(n27018), .ZN(n2552) );
  NAND3_X1 U8763 ( .A1(n29718), .A2(n17202), .A3(n17203), .ZN(n6335) );
  XOR2_X1 U8764 ( .A(n25188), .B(n28496), .Z(n6789) );
  NAND2_X1 U8766 ( .A1(n2839), .A2(n2840), .ZN(n6718) );
  INV_X1 U8767 ( .A(n14419), .ZN(n14420) );
  NAND3_X1 U8768 ( .A1(n13924), .A2(n14775), .A3(n13923), .ZN(n5893) );
  INV_X1 U8769 ( .A(n11330), .ZN(n8422) );
  XNOR2_X1 U8770 ( .A(n10145), .B(n2403), .ZN(n9935) );
  NAND3_X1 U8774 ( .A1(n23144), .A2(n24630), .A3(n24629), .ZN(n4365) );
  NAND3_X1 U8776 ( .A1(n8218), .A2(n7624), .A3(n7625), .ZN(n2556) );
  INV_X1 U8777 ( .A(n28195), .ZN(n5025) );
  NAND2_X1 U8779 ( .A1(n7896), .A2(n7897), .ZN(n7899) );
  INV_X1 U8780 ( .A(Plaintext[47]), .ZN(n2638) );
  OR3_X2 U8781 ( .A1(n21701), .A2(n21700), .A3(n21699), .ZN(n21872) );
  OAI21_X1 U8782 ( .B1(n499), .B2(n20180), .A(n20217), .ZN(n3078) );
  XNOR2_X2 U8783 ( .A(n21840), .B(n21839), .ZN(n23772) );
  NAND2_X1 U8785 ( .A1(n4849), .A2(n2557), .ZN(n24769) );
  NOR2_X1 U8786 ( .A1(n4847), .A2(n4848), .ZN(n2557) );
  NAND2_X1 U8787 ( .A1(n3429), .A2(n3430), .ZN(n3428) );
  NAND2_X1 U8788 ( .A1(n18020), .A2(n18018), .ZN(n2558) );
  NAND3_X1 U8789 ( .A1(n18603), .A2(n6714), .A3(n6713), .ZN(n18812) );
  NOR2_X1 U8790 ( .A1(n17475), .A2(n17478), .ZN(n2559) );
  INV_X1 U8791 ( .A(n17480), .ZN(n2560) );
  AND2_X1 U8792 ( .A1(n10810), .A2(n10473), .ZN(n11324) );
  NAND2_X1 U8794 ( .A1(n13839), .A2(n13838), .ZN(n2562) );
  INV_X1 U8795 ( .A(n11795), .ZN(n3558) );
  NAND2_X1 U8796 ( .A1(n3124), .A2(n24793), .ZN(n3714) );
  INV_X1 U8797 ( .A(n18330), .ZN(n6403) );
  NAND2_X1 U8798 ( .A1(n2563), .A2(n2663), .ZN(n10728) );
  NAND2_X1 U8799 ( .A1(n2661), .A2(n10927), .ZN(n2563) );
  NAND2_X1 U8800 ( .A1(n7531), .A2(n7141), .ZN(n2564) );
  NAND2_X1 U8801 ( .A1(n7532), .A2(n7523), .ZN(n2565) );
  OAI211_X1 U8802 ( .C1(n18591), .C2(n17837), .A(n17836), .B(n2044), .ZN(n2566) );
  INV_X1 U8803 ( .A(n20437), .ZN(n20611) );
  INV_X1 U8805 ( .A(n5945), .ZN(n6590) );
  XNOR2_X1 U8807 ( .A(n2567), .B(n15641), .ZN(n17030) );
  XNOR2_X1 U8808 ( .A(n15645), .B(n15640), .ZN(n2567) );
  NOR2_X1 U8809 ( .A1(n5164), .A2(n17888), .ZN(n5162) );
  NAND2_X1 U8810 ( .A1(n14084), .A2(n14286), .ZN(n13770) );
  XNOR2_X2 U8811 ( .A(n16225), .B(n16226), .ZN(n17138) );
  NAND3_X1 U8812 ( .A1(n21496), .A2(n28789), .A3(n21495), .ZN(n6749) );
  NAND2_X1 U8813 ( .A1(n11549), .A2(n11851), .ZN(n11548) );
  NAND3_X1 U8814 ( .A1(n7917), .A2(n7915), .A3(n7916), .ZN(n2569) );
  NOR2_X2 U8815 ( .A1(n3197), .A2(n18152), .ZN(n19376) );
  OAI211_X1 U8816 ( .C1(n18016), .C2(n18493), .A(n1997), .B(n3768), .ZN(n2571)
         );
  AOI21_X1 U8817 ( .B1(n21478), .B2(n1930), .A(n2572), .ZN(n21391) );
  OR2_X1 U8818 ( .A1(n15248), .A2(n15137), .ZN(n14116) );
  NAND2_X1 U8819 ( .A1(n2573), .A2(n14970), .ZN(n14977) );
  NAND2_X1 U8820 ( .A1(n5813), .A2(n14969), .ZN(n2573) );
  XNOR2_X1 U8823 ( .A(n2574), .B(n13522), .ZN(n12683) );
  XNOR2_X1 U8824 ( .A(n12680), .B(n13171), .ZN(n2574) );
  NAND2_X1 U8825 ( .A1(n6022), .A2(n6286), .ZN(n15583) );
  NAND3_X1 U8827 ( .A1(n2575), .A2(n23363), .A3(n3902), .ZN(n3901) );
  NAND2_X1 U8828 ( .A1(n16728), .A2(n17484), .ZN(n2578) );
  NAND2_X1 U8829 ( .A1(n17830), .A2(n17829), .ZN(n2579) );
  OR2_X1 U8830 ( .A1(n9220), .A2(n9221), .ZN(n9024) );
  OAI21_X1 U8831 ( .B1(n14843), .B2(n14844), .A(n15284), .ZN(n14848) );
  INV_X1 U8832 ( .A(n20551), .ZN(n6086) );
  NAND2_X1 U8834 ( .A1(n2581), .A2(n11816), .ZN(n11433) );
  OAI21_X1 U8835 ( .B1(n11724), .B2(n11819), .A(n11818), .ZN(n2581) );
  NAND2_X1 U8836 ( .A1(n2583), .A2(n2582), .ZN(n13863) );
  NAND2_X1 U8837 ( .A1(n13862), .A2(n14460), .ZN(n2582) );
  NAND2_X1 U8838 ( .A1(n2584), .A2(n3580), .ZN(n2583) );
  NAND2_X1 U8839 ( .A1(n14204), .A2(n14200), .ZN(n2584) );
  NOR2_X1 U8841 ( .A1(n14194), .A2(n29604), .ZN(n4434) );
  NAND2_X1 U8842 ( .A1(n2634), .A2(n526), .ZN(n2633) );
  OAI21_X1 U8843 ( .B1(n8532), .B2(n8709), .A(n2585), .ZN(n7035) );
  NAND2_X1 U8844 ( .A1(n8407), .A2(n8876), .ZN(n2585) );
  NOR2_X1 U8845 ( .A1(n8699), .A2(n8881), .ZN(n8407) );
  XNOR2_X1 U8846 ( .A(n19167), .B(n1989), .ZN(n19168) );
  NAND3_X1 U8847 ( .A1(n2586), .A2(n24593), .A3(n4692), .ZN(n4691) );
  NAND2_X1 U8848 ( .A1(n404), .A2(n24397), .ZN(n24674) );
  NAND2_X1 U8850 ( .A1(n2589), .A2(n29735), .ZN(n2587) );
  NAND2_X1 U8852 ( .A1(n7004), .A2(n2590), .ZN(n7005) );
  NOR2_X1 U8853 ( .A1(n2591), .A2(n17689), .ZN(n5201) );
  NAND3_X2 U8854 ( .A1(n2593), .A2(n2592), .A3(n2009), .ZN(n16272) );
  NAND2_X1 U8855 ( .A1(n14640), .A2(n15082), .ZN(n2593) );
  NAND2_X1 U8857 ( .A1(n20006), .A2(n20258), .ZN(n2594) );
  XNOR2_X1 U8859 ( .A(n9601), .B(n10228), .ZN(n10285) );
  NAND2_X1 U8860 ( .A1(n8597), .A2(n8819), .ZN(n2596) );
  INV_X1 U8861 ( .A(n8596), .ZN(n2597) );
  NAND2_X1 U8863 ( .A1(n2599), .A2(n16799), .ZN(n3017) );
  NAND3_X1 U8864 ( .A1(n3672), .A2(n17129), .A3(n2600), .ZN(n2599) );
  INV_X1 U8865 ( .A(n17990), .ZN(n18598) );
  NAND2_X1 U8866 ( .A1(n2601), .A2(n6152), .ZN(n6151) );
  NAND2_X1 U8867 ( .A1(n11133), .A2(n10457), .ZN(n2601) );
  OR2_X2 U8868 ( .A1(n6044), .A2(n13835), .ZN(n15180) );
  NAND2_X1 U8869 ( .A1(n8303), .A2(n8296), .ZN(n8299) );
  NAND2_X1 U8870 ( .A1(n17834), .A2(n18595), .ZN(n18130) );
  MUX2_X1 U8871 ( .A(n2610), .B(n17110), .S(n17106), .Z(n2609) );
  AOI21_X1 U8872 ( .B1(n10401), .B2(n8763), .A(n2104), .ZN(n8646) );
  NAND2_X1 U8873 ( .A1(n2611), .A2(n22742), .ZN(n2613) );
  NAND2_X1 U8874 ( .A1(n3043), .A2(n23286), .ZN(n2611) );
  MUX2_X1 U8875 ( .A(n24405), .B(n24404), .S(n24403), .Z(n23506) );
  AND3_X2 U8876 ( .A1(n2613), .A2(n3042), .A3(n2612), .ZN(n24403) );
  OAI22_X1 U8877 ( .A1(n11131), .A2(n2646), .B1(n4555), .B2(n2614), .ZN(n2655)
         );
  NAND2_X1 U8878 ( .A1(n10713), .A2(n10502), .ZN(n2614) );
  NAND2_X1 U8879 ( .A1(n27130), .A2(n29293), .ZN(n2615) );
  NOR2_X1 U8880 ( .A1(n27548), .A2(n27202), .ZN(n27545) );
  NAND2_X1 U8881 ( .A1(n2617), .A2(n28422), .ZN(n2618) );
  INV_X1 U8882 ( .A(n24437), .ZN(n23886) );
  INV_X1 U8883 ( .A(n24347), .ZN(n2619) );
  INV_X1 U8884 ( .A(n2621), .ZN(n2620) );
  OAI21_X1 U8886 ( .B1(n22994), .B2(n22995), .A(n22993), .ZN(n2623) );
  NAND2_X1 U8887 ( .A1(n2624), .A2(n7766), .ZN(n2629) );
  NAND2_X1 U8888 ( .A1(n2630), .A2(n2631), .ZN(n2625) );
  NAND2_X1 U8889 ( .A1(n8177), .A2(n2630), .ZN(n2626) );
  NAND3_X1 U8890 ( .A1(n2628), .A2(n2627), .A3(n2629), .ZN(n8335) );
  NAND2_X1 U8891 ( .A1(n2630), .A2(n2631), .ZN(n2627) );
  NAND2_X1 U8892 ( .A1(n8177), .A2(n2630), .ZN(n2628) );
  NAND2_X1 U8893 ( .A1(n8179), .A2(n8176), .ZN(n7766) );
  INV_X1 U8895 ( .A(n7289), .ZN(n2631) );
  NAND2_X1 U8896 ( .A1(n2632), .A2(n2122), .ZN(n5399) );
  NOR2_X1 U8897 ( .A1(n2632), .A2(n29483), .ZN(n15688) );
  NAND3_X1 U8898 ( .A1(n14376), .A2(n29059), .A3(n2849), .ZN(n6613) );
  NOR2_X1 U8899 ( .A1(n17847), .A2(n17846), .ZN(n2634) );
  NAND3_X1 U8900 ( .A1(n23024), .A2(n23539), .A3(n2637), .ZN(n6764) );
  NAND2_X1 U8901 ( .A1(n23687), .A2(n23801), .ZN(n2637) );
  NAND2_X1 U8902 ( .A1(n2637), .A2(n4337), .ZN(n4336) );
  AND2_X1 U8903 ( .A1(n21894), .A2(n2636), .ZN(n21895) );
  NAND2_X1 U8904 ( .A1(n7129), .A2(n29119), .ZN(n3148) );
  NAND3_X1 U8908 ( .A1(n14851), .A2(n2644), .A3(n2643), .ZN(n2642) );
  NAND2_X1 U8909 ( .A1(n15312), .A2(n15310), .ZN(n2643) );
  NAND3_X2 U8910 ( .A1(n5949), .A2(n6794), .A3(n14316), .ZN(n15310) );
  NAND2_X1 U8911 ( .A1(n15309), .A2(n15306), .ZN(n2644) );
  NAND2_X1 U8912 ( .A1(n14854), .A2(n14852), .ZN(n2645) );
  XNOR2_X2 U8913 ( .A(n9975), .B(n9974), .ZN(n10713) );
  NAND2_X1 U8914 ( .A1(n2648), .A2(n2647), .ZN(n24314) );
  NAND2_X1 U8915 ( .A1(n2649), .A2(n24391), .ZN(n2647) );
  NAND3_X1 U8917 ( .A1(n490), .A2(n21410), .A3(n20663), .ZN(n2650) );
  NAND2_X1 U8918 ( .A1(n21047), .A2(n2652), .ZN(n2651) );
  NOR2_X1 U8919 ( .A1(n21410), .A2(n21171), .ZN(n2652) );
  INV_X1 U8923 ( .A(n17889), .ZN(n2656) );
  NAND2_X1 U8924 ( .A1(n2659), .A2(n2657), .ZN(n7114) );
  OAI21_X1 U8925 ( .B1(n2658), .B2(n2631), .A(n8179), .ZN(n2657) );
  INV_X1 U8926 ( .A(n7290), .ZN(n2658) );
  NAND2_X1 U8929 ( .A1(n7289), .A2(n8173), .ZN(n7347) );
  NAND2_X1 U8930 ( .A1(n10930), .A2(n10932), .ZN(n2661) );
  NAND2_X1 U8931 ( .A1(n10727), .A2(n10929), .ZN(n2663) );
  NAND2_X1 U8933 ( .A1(n2741), .A2(n2664), .ZN(n16938) );
  AND2_X1 U8935 ( .A1(n21665), .A2(n3666), .ZN(n2669) );
  NAND3_X1 U8936 ( .A1(n9142), .A2(n8564), .A3(n599), .ZN(n8565) );
  NAND2_X1 U8937 ( .A1(n2670), .A2(n7331), .ZN(n7335) );
  AND2_X1 U8942 ( .A1(n13827), .A2(n14278), .ZN(n4369) );
  OAI21_X1 U8943 ( .B1(n28507), .B2(n4166), .A(n29691), .ZN(n13618) );
  XNOR2_X2 U8945 ( .A(n2675), .B(Key[23]), .ZN(n7330) );
  INV_X1 U8946 ( .A(Plaintext[23]), .ZN(n2675) );
  XNOR2_X1 U8947 ( .A(n2677), .B(n27952), .ZN(n7415) );
  XNOR2_X1 U8948 ( .A(n2677), .B(n3114), .ZN(n9740) );
  XNOR2_X1 U8949 ( .A(n9639), .B(n2677), .ZN(n9403) );
  XNOR2_X1 U8950 ( .A(n9702), .B(n2677), .ZN(n10368) );
  INV_X1 U8951 ( .A(n11310), .ZN(n2680) );
  NAND2_X1 U8952 ( .A1(n11163), .A2(n29637), .ZN(n11310) );
  NOR2_X1 U8953 ( .A1(n2681), .A2(n14260), .ZN(n2945) );
  NAND2_X1 U8954 ( .A1(n13614), .A2(n2681), .ZN(n12369) );
  NAND2_X1 U8957 ( .A1(n28203), .A2(n12109), .ZN(n2684) );
  NAND2_X1 U8958 ( .A1(n9655), .A2(n12109), .ZN(n2685) );
  AND2_X1 U8960 ( .A1(n11258), .A2(n2690), .ZN(n4326) );
  NAND2_X1 U8961 ( .A1(n2689), .A2(n2687), .ZN(n11023) );
  AND2_X1 U8962 ( .A1(n2690), .A2(n11318), .ZN(n2687) );
  MUX2_X1 U8963 ( .A(n2690), .B(n11254), .S(n594), .Z(n9503) );
  NAND2_X1 U8964 ( .A1(n14929), .A2(n2691), .ZN(n15781) );
  NAND2_X1 U8965 ( .A1(n7163), .A2(n7164), .ZN(n7771) );
  AOI21_X1 U8966 ( .B1(n2694), .B2(n17719), .A(n18081), .ZN(n6229) );
  OAI22_X1 U8967 ( .A1(n2694), .A2(n18285), .B1(n373), .B2(n17719), .ZN(n3753)
         );
  OAI21_X1 U8968 ( .B1(n18525), .B2(n18523), .A(n2694), .ZN(n18287) );
  NAND2_X1 U8970 ( .A1(n2696), .A2(n7985), .ZN(n2695) );
  NAND2_X1 U8971 ( .A1(n7983), .A2(n7984), .ZN(n2696) );
  NAND2_X1 U8973 ( .A1(n23656), .A2(n4232), .ZN(n2697) );
  NOR2_X1 U8974 ( .A1(n11666), .A2(n3946), .ZN(n11667) );
  XNOR2_X1 U8975 ( .A(n2700), .B(n2996), .ZN(n14675) );
  XNOR2_X1 U8976 ( .A(n2700), .B(n1046), .ZN(n16034) );
  XNOR2_X1 U8977 ( .A(n2700), .B(n3323), .ZN(n16511) );
  XNOR2_X1 U8978 ( .A(n16470), .B(n2700), .ZN(n16375) );
  NAND2_X1 U8979 ( .A1(n535), .A2(n17368), .ZN(n17233) );
  NAND2_X1 U8980 ( .A1(n2701), .A2(n17046), .ZN(n15732) );
  NAND2_X1 U8981 ( .A1(n535), .A2(n17234), .ZN(n17235) );
  NAND2_X1 U8982 ( .A1(n17043), .A2(n535), .ZN(n3549) );
  NOR2_X1 U8985 ( .A1(n18530), .A2(n29476), .ZN(n2702) );
  NAND2_X1 U8988 ( .A1(n509), .A2(n18529), .ZN(n18259) );
  NAND2_X1 U8989 ( .A1(n22084), .A2(n2708), .ZN(n6220) );
  AOI21_X1 U8990 ( .B1(n28431), .B2(n2708), .A(n28622), .ZN(n22085) );
  INV_X1 U8991 ( .A(n23706), .ZN(n2708) );
  XNOR2_X1 U8992 ( .A(n10344), .B(n3067), .ZN(n2711) );
  XNOR2_X1 U8993 ( .A(n2711), .B(n9698), .ZN(n9301) );
  INV_X1 U8994 ( .A(n8506), .ZN(n2713) );
  NAND2_X1 U8995 ( .A1(n563), .A2(n2714), .ZN(n13767) );
  NAND2_X1 U8996 ( .A1(n2715), .A2(n20155), .ZN(n4410) );
  OAI22_X1 U8997 ( .A1(n2815), .A2(n2715), .B1(n20100), .B2(n20101), .ZN(
        n20533) );
  NAND2_X1 U8998 ( .A1(n2717), .A2(n614), .ZN(n7165) );
  NAND2_X1 U8999 ( .A1(n7321), .A2(n7770), .ZN(n2717) );
  AND2_X1 U9000 ( .A1(n2718), .A2(n4756), .ZN(n6264) );
  NAND2_X1 U9001 ( .A1(n5021), .A2(n5023), .ZN(n2718) );
  NOR2_X1 U9002 ( .A1(n5439), .A2(n18230), .ZN(n19024) );
  OAI211_X1 U9003 ( .C1(n5439), .C2(n2723), .A(n2722), .B(n2721), .ZN(n18767)
         );
  NAND2_X1 U9004 ( .A1(n18230), .A2(n1887), .ZN(n2721) );
  NAND2_X1 U9005 ( .A1(n5439), .A2(n1887), .ZN(n2722) );
  INV_X1 U9008 ( .A(n14744), .ZN(n2727) );
  NAND2_X1 U9009 ( .A1(n29604), .A2(n14393), .ZN(n4436) );
  NAND2_X1 U9010 ( .A1(n2728), .A2(n14194), .ZN(n14394) );
  NAND2_X1 U9011 ( .A1(n14395), .A2(n29604), .ZN(n4047) );
  NAND2_X1 U9012 ( .A1(n13951), .A2(n29604), .ZN(n13870) );
  OAI22_X1 U9013 ( .A1(n5745), .A2(n14393), .B1(n28805), .B2(n29604), .ZN(
        n6283) );
  NAND4_X1 U9014 ( .A1(n14597), .A2(n6921), .A3(n2729), .A4(n14258), .ZN(n2730) );
  NAND2_X1 U9016 ( .A1(n15105), .A2(n15423), .ZN(n14934) );
  NAND2_X1 U9017 ( .A1(n2002), .A2(n15105), .ZN(n2732) );
  NAND2_X1 U9018 ( .A1(n15423), .A2(n549), .ZN(n2733) );
  NAND2_X1 U9019 ( .A1(n29104), .A2(n2735), .ZN(n6409) );
  OAI21_X1 U9020 ( .B1(n20093), .B2(n20041), .A(n2734), .ZN(n18789) );
  NAND2_X1 U9021 ( .A1(n20041), .A2(n20088), .ZN(n2734) );
  OAI22_X1 U9022 ( .A1(n20087), .A2(n19757), .B1(n20092), .B2(n2735), .ZN(
        n19758) );
  NAND2_X1 U9023 ( .A1(n24705), .A2(n2736), .ZN(n24710) );
  NAND2_X1 U9024 ( .A1(n24709), .A2(n29043), .ZN(n2736) );
  NAND2_X1 U9025 ( .A1(n2737), .A2(n14761), .ZN(n15264) );
  NAND3_X2 U9026 ( .A1(n14245), .A2(n14247), .A3(n14246), .ZN(n14761) );
  INV_X1 U9027 ( .A(n14762), .ZN(n2737) );
  NAND2_X1 U9028 ( .A1(n4162), .A2(n15260), .ZN(n4097) );
  NAND2_X1 U9029 ( .A1(n8504), .A2(n8886), .ZN(n2739) );
  NAND3_X1 U9031 ( .A1(n8504), .A2(n8336), .A3(n8889), .ZN(n2740) );
  NAND2_X1 U9033 ( .A1(n17335), .A2(n28564), .ZN(n17203) );
  NAND3_X1 U9034 ( .A1(n15180), .A2(n28803), .A3(n14534), .ZN(n2744) );
  OR2_X1 U9036 ( .A1(n3954), .A2(n1908), .ZN(n2746) );
  NAND3_X1 U9037 ( .A1(n20455), .A2(n20454), .A3(n20632), .ZN(n20456) );
  NAND2_X1 U9038 ( .A1(n20033), .A2(n20634), .ZN(n20455) );
  NAND2_X1 U9040 ( .A1(n5172), .A2(n5171), .ZN(n2749) );
  AND2_X1 U9041 ( .A1(n23363), .A2(n23360), .ZN(n21302) );
  OAI211_X2 U9042 ( .C1(n486), .C2(n23069), .A(n2751), .B(n2750), .ZN(n24711)
         );
  NAND2_X1 U9043 ( .A1(n23674), .A2(n23363), .ZN(n2750) );
  NAND2_X1 U9044 ( .A1(n23068), .A2(n486), .ZN(n2751) );
  NAND3_X1 U9045 ( .A1(n29122), .A2(n11047), .A3(n2753), .ZN(n9653) );
  NAND3_X1 U9046 ( .A1(n11260), .A2(n11266), .A3(n2753), .ZN(n10669) );
  INV_X1 U9047 ( .A(n11267), .ZN(n2753) );
  NAND2_X1 U9050 ( .A1(n11260), .A2(n11045), .ZN(n2755) );
  NAND3_X1 U9051 ( .A1(n1954), .A2(n2757), .A3(n2756), .ZN(n17770) );
  NAND3_X1 U9052 ( .A1(n17764), .A2(n3597), .A3(n28073), .ZN(n2756) );
  NAND2_X1 U9053 ( .A1(n2758), .A2(n1133), .ZN(n2757) );
  XNOR2_X1 U9054 ( .A(n2759), .B(n3321), .ZN(n19341) );
  XNOR2_X1 U9055 ( .A(n2759), .B(n3643), .ZN(n19633) );
  XNOR2_X1 U9056 ( .A(n2759), .B(n2986), .ZN(n18662) );
  XNOR2_X1 U9057 ( .A(n19688), .B(n2759), .ZN(n18868) );
  XNOR2_X1 U9058 ( .A(n19111), .B(n2759), .ZN(n19112) );
  NAND2_X1 U9059 ( .A1(n2761), .A2(n2760), .ZN(n23909) );
  NAND3_X1 U9060 ( .A1(n24405), .A2(n24083), .A3(n24403), .ZN(n2760) );
  NAND3_X1 U9061 ( .A1(n24408), .A2(n24404), .A3(n2762), .ZN(n2761) );
  INV_X1 U9062 ( .A(n27846), .ZN(n2765) );
  NAND3_X1 U9063 ( .A1(n27843), .A2(n27826), .A3(n27825), .ZN(n2763) );
  NAND2_X1 U9064 ( .A1(n2767), .A2(n3542), .ZN(n2764) );
  INV_X1 U9066 ( .A(n17567), .ZN(n2769) );
  NAND2_X1 U9067 ( .A1(n17759), .A2(n17758), .ZN(n2770) );
  NAND2_X1 U9068 ( .A1(n17969), .A2(n18236), .ZN(n17756) );
  NAND2_X1 U9069 ( .A1(n2773), .A2(n1354), .ZN(n2772) );
  NAND2_X1 U9070 ( .A1(n7888), .A2(n7777), .ZN(n2773) );
  NAND2_X1 U9071 ( .A1(n7778), .A2(n7315), .ZN(n7888) );
  INV_X1 U9072 ( .A(n17818), .ZN(n18413) );
  INV_X1 U9073 ( .A(n18120), .ZN(n2777) );
  NOR2_X1 U9074 ( .A1(n18414), .A2(n18410), .ZN(n2778) );
  NOR2_X1 U9075 ( .A1(n18411), .A2(n17818), .ZN(n18120) );
  NAND2_X1 U9077 ( .A1(n23651), .A2(n2779), .ZN(n23194) );
  NAND2_X1 U9078 ( .A1(n23046), .A2(n23654), .ZN(n23652) );
  MUX2_X1 U9079 ( .A(n23649), .B(n23650), .S(n23470), .Z(n23653) );
  NAND2_X1 U9080 ( .A1(n8019), .A2(n7747), .ZN(n2780) );
  OAI22_X1 U9081 ( .A1(n7746), .A2(n7745), .B1(n7743), .B2(n7744), .ZN(n2781)
         );
  NAND2_X1 U9082 ( .A1(n2783), .A2(n13703), .ZN(n14424) );
  NAND2_X1 U9083 ( .A1(n2783), .A2(n14426), .ZN(n14305) );
  NAND2_X1 U9084 ( .A1(n4522), .A2(n2783), .ZN(n12532) );
  AND2_X1 U9086 ( .A1(n2783), .A2(n29558), .ZN(n2782) );
  INV_X1 U9087 ( .A(n12534), .ZN(n2783) );
  MUX2_X1 U9089 ( .A(n23657), .B(n23351), .S(n29583), .Z(n23143) );
  INV_X1 U9090 ( .A(n19354), .ZN(n19655) );
  NAND3_X1 U9091 ( .A1(n2786), .A2(n17844), .A3(n18243), .ZN(n2784) );
  NAND2_X1 U9092 ( .A1(n2787), .A2(n17843), .ZN(n2785) );
  INV_X1 U9093 ( .A(n7506), .ZN(n6210) );
  XNOR2_X2 U9094 ( .A(Key[57]), .B(Plaintext[57]), .ZN(n7506) );
  NAND2_X1 U9095 ( .A1(n7514), .A2(n7506), .ZN(n2788) );
  XNOR2_X1 U9096 ( .A(n15853), .B(n15852), .ZN(n2790) );
  NAND2_X1 U9097 ( .A1(n18062), .A2(n2791), .ZN(n4348) );
  OAI22_X1 U9099 ( .A1(n17929), .A2(n2791), .B1(n18061), .B2(n17928), .ZN(
        n17930) );
  NAND2_X1 U9100 ( .A1(n397), .A2(n27744), .ZN(n2795) );
  NAND2_X1 U9102 ( .A1(n2797), .A2(n5303), .ZN(n2796) );
  NAND2_X1 U9103 ( .A1(n15208), .A2(n14928), .ZN(n15206) );
  INV_X1 U9104 ( .A(n15206), .ZN(n2800) );
  OAI211_X1 U9105 ( .C1(n2803), .C2(n18788), .A(n2802), .B(n2801), .ZN(n22312)
         );
  NAND2_X1 U9106 ( .A1(n18788), .A2(n2804), .ZN(n2801) );
  NAND2_X1 U9107 ( .A1(n18787), .A2(n2804), .ZN(n2802) );
  INV_X1 U9108 ( .A(Key[15]), .ZN(n2804) );
  XNOR2_X1 U9109 ( .A(n2805), .B(n22295), .ZN(n21850) );
  XNOR2_X1 U9110 ( .A(n2805), .B(n22073), .ZN(n20680) );
  NOR2_X1 U9111 ( .A1(n2806), .A2(n24976), .ZN(n24512) );
  OAI21_X1 U9112 ( .B1(n24975), .B2(n2806), .A(n24259), .ZN(n25059) );
  OAI211_X2 U9113 ( .C1(n23804), .C2(n28919), .A(n1976), .B(n2807), .ZN(n26054) );
  NAND2_X1 U9114 ( .A1(n2808), .A2(n24653), .ZN(n24028) );
  INV_X1 U9115 ( .A(n24651), .ZN(n2808) );
  NAND2_X1 U9116 ( .A1(n24029), .A2(n2809), .ZN(n24031) );
  NOR2_X1 U9117 ( .A1(n28481), .A2(n24523), .ZN(n2809) );
  NOR2_X1 U9118 ( .A1(n24651), .A2(n629), .ZN(n2810) );
  INV_X1 U9119 ( .A(n17846), .ZN(n2811) );
  XNOR2_X1 U9120 ( .A(n25343), .B(n25340), .ZN(n2813) );
  NAND3_X1 U9121 ( .A1(n1888), .A2(n18020), .A3(n18251), .ZN(n3069) );
  NAND2_X1 U9122 ( .A1(n2814), .A2(n2834), .ZN(n3084) );
  INV_X1 U9123 ( .A(n20156), .ZN(n2815) );
  NAND2_X1 U9124 ( .A1(n24513), .A2(n24421), .ZN(n2816) );
  NAND2_X1 U9126 ( .A1(n23748), .A2(n23749), .ZN(n2817) );
  XNOR2_X2 U9127 ( .A(n15931), .B(n15930), .ZN(n17570) );
  AOI21_X2 U9128 ( .B1(n2821), .B2(n6868), .A(n2820), .ZN(n25903) );
  NOR2_X1 U9129 ( .A1(n23126), .A2(n24020), .ZN(n24160) );
  INV_X1 U9130 ( .A(n24538), .ZN(n2823) );
  NAND2_X1 U9131 ( .A1(n24159), .A2(n24542), .ZN(n2824) );
  NAND2_X1 U9132 ( .A1(n23126), .A2(n24001), .ZN(n24159) );
  INV_X1 U9133 ( .A(n17424), .ZN(n2826) );
  INV_X1 U9134 ( .A(n17424), .ZN(n2825) );
  NAND2_X1 U9135 ( .A1(n2825), .A2(n17425), .ZN(n17008) );
  NAND2_X1 U9137 ( .A1(n24450), .A2(n24757), .ZN(n2828) );
  NAND3_X1 U9138 ( .A1(n24761), .A2(n28509), .A3(n24758), .ZN(n2829) );
  OAI211_X2 U9139 ( .C1(n21522), .C2(n21550), .A(n21521), .B(n2830), .ZN(
        n22567) );
  AND2_X1 U9140 ( .A1(n17393), .A2(n17293), .ZN(n16958) );
  NAND2_X1 U9141 ( .A1(n5487), .A2(n533), .ZN(n17000) );
  NAND2_X1 U9142 ( .A1(n16961), .A2(n533), .ZN(n5326) );
  AOI22_X1 U9143 ( .A1(n2831), .A2(n15268), .B1(n14703), .B2(n15269), .ZN(
        n14704) );
  INV_X1 U9144 ( .A(n14618), .ZN(n2831) );
  OAI21_X1 U9145 ( .B1(n15269), .B2(n3748), .A(n2831), .ZN(n15270) );
  INV_X1 U9146 ( .A(n7233), .ZN(n2832) );
  INV_X1 U9148 ( .A(n7589), .ZN(n2833) );
  NOR3_X1 U9149 ( .A1(n18017), .A2(n2834), .A3(n18020), .ZN(n17960) );
  NAND2_X1 U9150 ( .A1(n18022), .A2(n2834), .ZN(n3068) );
  NOR2_X1 U9151 ( .A1(n18353), .A2(n18354), .ZN(n2836) );
  NAND2_X1 U9152 ( .A1(n18311), .A2(n518), .ZN(n2837) );
  NAND3_X1 U9153 ( .A1(n6719), .A2(n6905), .A3(n7926), .ZN(n2839) );
  NAND3_X1 U9154 ( .A1(n7398), .A2(n6719), .A3(n7625), .ZN(n2840) );
  NAND3_X1 U9156 ( .A1(n7514), .A2(n7506), .A3(n29629), .ZN(n2841) );
  NAND2_X1 U9157 ( .A1(n28182), .A2(n23289), .ZN(n2842) );
  NAND2_X1 U9158 ( .A1(n2842), .A2(n23816), .ZN(n4415) );
  NAND2_X1 U9159 ( .A1(n2027), .A2(n12132), .ZN(n5039) );
  MUX2_X1 U9160 ( .A(n29149), .B(n3820), .S(n11033), .Z(n2843) );
  NAND2_X1 U9161 ( .A1(n8898), .A2(n8900), .ZN(n2844) );
  NOR2_X1 U9162 ( .A1(n81), .A2(n9124), .ZN(n8900) );
  XNOR2_X1 U9163 ( .A(n10251), .B(n2845), .ZN(n9907) );
  XNOR2_X1 U9164 ( .A(n10151), .B(n2845), .ZN(n10152) );
  XNOR2_X1 U9165 ( .A(n2845), .B(n15576), .ZN(n9621) );
  NAND3_X1 U9167 ( .A1(n6163), .A2(n10638), .A3(n6165), .ZN(n2846) );
  NOR2_X1 U9168 ( .A1(n2846), .A2(n12042), .ZN(n12044) );
  INV_X1 U9170 ( .A(n14372), .ZN(n2849) );
  NAND2_X1 U9171 ( .A1(n16985), .A2(n19560), .ZN(n17639) );
  XNOR2_X1 U9172 ( .A(n2850), .B(n24906), .ZN(Ciphertext[13]) );
  OAI21_X1 U9173 ( .B1(n4090), .B2(n2852), .A(n2851), .ZN(n2850) );
  INV_X1 U9174 ( .A(n27376), .ZN(n2851) );
  NAND2_X1 U9175 ( .A1(n5372), .A2(n5374), .ZN(n2852) );
  INV_X1 U9176 ( .A(n2853), .ZN(n18045) );
  NAND2_X1 U9177 ( .A1(n17225), .A2(n17224), .ZN(n2853) );
  NAND2_X1 U9178 ( .A1(n2853), .A2(n18430), .ZN(n17610) );
  NAND2_X1 U9179 ( .A1(n1894), .A2(n2853), .ZN(n18146) );
  NAND2_X1 U9181 ( .A1(n18432), .A2(n2854), .ZN(n18435) );
  NOR2_X1 U9182 ( .A1(n2855), .A2(n18045), .ZN(n2854) );
  NAND2_X1 U9183 ( .A1(n17482), .A2(n4271), .ZN(n2857) );
  NAND2_X1 U9186 ( .A1(n2864), .A2(n9070), .ZN(n2859) );
  NAND2_X1 U9187 ( .A1(n602), .A2(n8819), .ZN(n8475) );
  NAND2_X1 U9188 ( .A1(n2024), .A2(n8594), .ZN(n2860) );
  NAND2_X1 U9189 ( .A1(n2862), .A2(n8977), .ZN(n2861) );
  NAND2_X1 U9190 ( .A1(n5962), .A2(n8593), .ZN(n2862) );
  NAND3_X1 U9191 ( .A1(n602), .A2(n8819), .A3(n8594), .ZN(n2863) );
  NAND2_X1 U9192 ( .A1(n9072), .A2(n8741), .ZN(n2864) );
  NAND2_X1 U9193 ( .A1(n378), .A2(n24447), .ZN(n5991) );
  AND2_X1 U9196 ( .A1(n28996), .A2(n14695), .ZN(n14846) );
  INV_X1 U9197 ( .A(n20152), .ZN(n20097) );
  NAND2_X1 U9198 ( .A1(n2871), .A2(n2870), .ZN(n18890) );
  NAND3_X1 U9199 ( .A1(n5053), .A2(n20096), .A3(n20152), .ZN(n2870) );
  XNOR2_X2 U9200 ( .A(n18819), .B(n18818), .ZN(n20152) );
  NAND3_X1 U9201 ( .A1(n28188), .A2(n20098), .A3(n20155), .ZN(n2871) );
  INV_X1 U9203 ( .A(n2872), .ZN(n20052) );
  NAND2_X1 U9204 ( .A1(n20066), .A2(n20064), .ZN(n2872) );
  NAND2_X1 U9205 ( .A1(n3436), .A2(n2872), .ZN(n20051) );
  NAND2_X1 U9206 ( .A1(n6924), .A2(n2874), .ZN(n2873) );
  NAND2_X1 U9207 ( .A1(n2876), .A2(n26840), .ZN(n2877) );
  INV_X1 U9208 ( .A(n25815), .ZN(n2876) );
  XNOR2_X1 U9209 ( .A(n25813), .B(n25812), .ZN(n26507) );
  NAND3_X1 U9210 ( .A1(n24747), .A2(n24745), .A3(n2879), .ZN(n2878) );
  NAND2_X1 U9211 ( .A1(n29545), .A2(n28550), .ZN(n4980) );
  AND2_X1 U9212 ( .A1(n21303), .A2(n24745), .ZN(n24746) );
  INV_X1 U9213 ( .A(n4675), .ZN(n8827) );
  NAND2_X1 U9214 ( .A1(n3004), .A2(n7886), .ZN(n2883) );
  NAND3_X1 U9215 ( .A1(n15008), .A2(n15369), .A3(n426), .ZN(n5093) );
  NAND2_X1 U9217 ( .A1(n15236), .A2(n15235), .ZN(n2885) );
  NAND2_X1 U9219 ( .A1(n26385), .A2(n26384), .ZN(n27166) );
  NAND2_X1 U9220 ( .A1(n2888), .A2(n2887), .ZN(n23132) );
  NAND2_X1 U9221 ( .A1(n23360), .A2(n23673), .ZN(n2887) );
  NAND2_X1 U9222 ( .A1(n18521), .A2(n17724), .ZN(n3544) );
  NAND2_X1 U9223 ( .A1(n18286), .A2(n17719), .ZN(n17724) );
  NAND2_X1 U9224 ( .A1(n1925), .A2(n21425), .ZN(n3238) );
  NAND2_X1 U9226 ( .A1(n3266), .A2(n6543), .ZN(n23491) );
  NAND2_X1 U9228 ( .A1(n10403), .A2(n10402), .ZN(n2892) );
  NAND3_X1 U9229 ( .A1(n432), .A2(n5258), .A3(n11094), .ZN(n11095) );
  NAND3_X1 U9230 ( .A1(n19837), .A2(n20381), .A3(n20383), .ZN(n4361) );
  OR2_X1 U9231 ( .A1(n10003), .A2(n10002), .ZN(n10004) );
  OAI21_X1 U9232 ( .B1(n19960), .B2(n19819), .A(n20545), .ZN(n3473) );
  NOR2_X1 U9233 ( .A1(n27551), .A2(n29578), .ZN(n27217) );
  MUX2_X1 U9234 ( .A(n12371), .B(n12370), .S(n3362), .Z(n2895) );
  NAND3_X2 U9235 ( .A1(n4160), .A2(n4159), .A3(n2896), .ZN(n9037) );
  NAND2_X1 U9236 ( .A1(n7853), .A2(n2897), .ZN(n2896) );
  OAI211_X2 U9239 ( .C1(n21319), .C2(n21320), .A(n21318), .B(n21317), .ZN(
        n22152) );
  NAND2_X1 U9240 ( .A1(n21674), .A2(n21448), .ZN(n4460) );
  NAND2_X1 U9242 ( .A1(n5779), .A2(n5780), .ZN(n21596) );
  INV_X1 U9243 ( .A(n10884), .ZN(n11284) );
  NAND2_X1 U9245 ( .A1(n18592), .A2(n3450), .ZN(n2901) );
  INV_X1 U9248 ( .A(n4504), .ZN(n16085) );
  AND2_X1 U9249 ( .A1(n12234), .A2(n375), .ZN(n6871) );
  XNOR2_X1 U9250 ( .A(n2902), .B(n26113), .ZN(n26125) );
  XNOR2_X1 U9251 ( .A(n2903), .B(n22545), .ZN(n22017) );
  XNOR2_X1 U9252 ( .A(n22016), .B(n6141), .ZN(n2903) );
  NOR2_X1 U9253 ( .A1(n2904), .A2(n10920), .ZN(n10921) );
  NAND2_X1 U9254 ( .A1(n10919), .A2(n11135), .ZN(n2904) );
  NAND2_X1 U9256 ( .A1(n24377), .A2(n24376), .ZN(n2905) );
  NAND2_X1 U9257 ( .A1(n24379), .A2(n24378), .ZN(n2906) );
  NAND2_X1 U9259 ( .A1(n2908), .A2(n9071), .ZN(n2907) );
  NOR2_X1 U9260 ( .A1(n18223), .A2(n18222), .ZN(n17499) );
  NAND2_X1 U9262 ( .A1(n11294), .A2(n10318), .ZN(n10309) );
  NAND2_X1 U9263 ( .A1(n7750), .A2(n7349), .ZN(n7751) );
  NAND2_X1 U9264 ( .A1(n5694), .A2(n17215), .ZN(n16751) );
  INV_X1 U9266 ( .A(n27065), .ZN(n3178) );
  NAND2_X1 U9267 ( .A1(n5016), .A2(n14652), .ZN(n4642) );
  NOR2_X1 U9268 ( .A1(n24244), .A2(n2913), .ZN(n25065) );
  AND2_X1 U9269 ( .A1(n24238), .A2(n24559), .ZN(n2913) );
  INV_X1 U9270 ( .A(n11819), .ZN(n12190) );
  INV_X1 U9271 ( .A(n24717), .ZN(n4136) );
  AND2_X1 U9272 ( .A1(n23474), .A2(n23761), .ZN(n23190) );
  OAI21_X1 U9273 ( .B1(n9868), .B2(n12186), .A(n9867), .ZN(n13396) );
  NAND2_X1 U9275 ( .A1(n435), .A2(n10534), .ZN(n11104) );
  INV_X1 U9276 ( .A(n24404), .ZN(n24085) );
  OR3_X1 U9277 ( .A1(n29602), .A2(n22531), .A3(n29020), .ZN(n5713) );
  MUX2_X1 U9278 ( .A(n20051), .B(n20050), .S(n20063), .Z(n21210) );
  INV_X1 U9280 ( .A(n24316), .ZN(n24667) );
  XNOR2_X1 U9281 ( .A(n13097), .B(n12377), .ZN(n13229) );
  OR2_X1 U9282 ( .A1(n14195), .A2(n5978), .ZN(n4435) );
  AND2_X1 U9283 ( .A1(n18410), .A2(n17818), .ZN(n4240) );
  INV_X1 U9284 ( .A(n13922), .ZN(n14775) );
  XNOR2_X1 U9285 ( .A(n22316), .B(n22317), .ZN(n4003) );
  INV_X1 U9286 ( .A(n17620), .ZN(n18159) );
  INV_X1 U9287 ( .A(n3315), .ZN(n15099) );
  XNOR2_X1 U9288 ( .A(n9763), .B(n10074), .ZN(n10277) );
  INV_X1 U9289 ( .A(n12110), .ZN(n12208) );
  INV_X1 U9290 ( .A(n6000), .ZN(n12976) );
  OAI21_X1 U9292 ( .B1(n14175), .B2(n14239), .A(n14174), .ZN(n3011) );
  XNOR2_X1 U9293 ( .A(n12490), .B(n11389), .ZN(n3687) );
  NAND2_X1 U9295 ( .A1(n8448), .A2(n8451), .ZN(n8449) );
  NAND2_X1 U9296 ( .A1(n3330), .A2(n3329), .ZN(n2917) );
  NAND2_X1 U9297 ( .A1(n6718), .A2(n9132), .ZN(n8550) );
  NOR2_X1 U9298 ( .A1(n24892), .A2(n24227), .ZN(n24229) );
  NAND2_X1 U9299 ( .A1(n23134), .A2(n6035), .ZN(n5884) );
  NAND2_X1 U9300 ( .A1(n7438), .A2(n7626), .ZN(n6719) );
  NAND2_X1 U9301 ( .A1(n24245), .A2(n24246), .ZN(n24247) );
  OR2_X1 U9302 ( .A1(n11168), .A2(n10820), .ZN(n10746) );
  NAND2_X1 U9303 ( .A1(n2920), .A2(n2919), .ZN(n23069) );
  NAND2_X1 U9304 ( .A1(n23366), .A2(n23131), .ZN(n2919) );
  NAND2_X1 U9305 ( .A1(n23364), .A2(n2921), .ZN(n2920) );
  INV_X1 U9306 ( .A(n23131), .ZN(n2921) );
  NAND2_X1 U9308 ( .A1(n20429), .A2(n20619), .ZN(n2922) );
  NAND2_X1 U9310 ( .A1(n2927), .A2(n2924), .ZN(n9392) );
  NAND2_X1 U9311 ( .A1(n2925), .A2(n8077), .ZN(n2924) );
  OAI21_X1 U9312 ( .B1(n8430), .B2(n8119), .A(n2926), .ZN(n2925) );
  NAND2_X1 U9313 ( .A1(n261), .A2(n8426), .ZN(n2926) );
  NAND2_X1 U9314 ( .A1(n8432), .A2(n8431), .ZN(n2927) );
  NAND2_X1 U9315 ( .A1(n8936), .A2(n2928), .ZN(n8938) );
  NAND2_X1 U9316 ( .A1(n3032), .A2(n377), .ZN(n2929) );
  NAND2_X1 U9317 ( .A1(n20574), .A2(n20568), .ZN(n2930) );
  NAND2_X1 U9318 ( .A1(n19836), .A2(n20573), .ZN(n2931) );
  OAI21_X1 U9325 ( .B1(n3072), .B2(n14261), .A(n2934), .ZN(n14270) );
  NAND2_X1 U9326 ( .A1(n3071), .A2(n14263), .ZN(n2934) );
  NAND2_X1 U9330 ( .A1(n24792), .A2(n24269), .ZN(n2938) );
  NAND2_X1 U9331 ( .A1(n466), .A2(n29567), .ZN(n2939) );
  NAND2_X1 U9332 ( .A1(n29471), .A2(n24310), .ZN(n2940) );
  NAND2_X1 U9333 ( .A1(n7350), .A2(n7351), .ZN(n2941) );
  NAND2_X1 U9334 ( .A1(n11101), .A2(n11896), .ZN(n2943) );
  XNOR2_X2 U9335 ( .A(n5066), .B(n22901), .ZN(n23456) );
  NOR2_X1 U9337 ( .A1(n5403), .A2(n14376), .ZN(n14377) );
  NOR2_X1 U9338 ( .A1(n1991), .A2(n3031), .ZN(n3030) );
  OAI211_X1 U9339 ( .C1(n20240), .C2(n20239), .A(n3532), .B(n29527), .ZN(
        n20361) );
  OAI21_X1 U9340 ( .B1(n15098), .B2(n14901), .A(n15099), .ZN(n3316) );
  NAND2_X1 U9342 ( .A1(n11982), .A2(n11980), .ZN(n12227) );
  OR2_X1 U9343 ( .A1(n13703), .A2(n12534), .ZN(n4665) );
  NAND2_X1 U9344 ( .A1(n7744), .A2(n8013), .ZN(n8016) );
  OR2_X1 U9346 ( .A1(n27119), .A2(n29016), .ZN(n3456) );
  NAND3_X1 U9347 ( .A1(n5771), .A2(n2950), .A3(n2949), .ZN(n18646) );
  NAND2_X1 U9348 ( .A1(n17907), .A2(n18343), .ZN(n2949) );
  NAND2_X1 U9349 ( .A1(n17909), .A2(n17908), .ZN(n2950) );
  AND2_X1 U9350 ( .A1(n19949), .A2(n20196), .ZN(n20590) );
  NAND2_X1 U9351 ( .A1(n21322), .A2(n20886), .ZN(n6042) );
  NAND2_X1 U9352 ( .A1(n23732), .A2(n2951), .ZN(n23737) );
  NAND2_X1 U9353 ( .A1(n2963), .A2(n2952), .ZN(n7385) );
  NAND3_X1 U9354 ( .A1(n7384), .A2(n7853), .A3(n7496), .ZN(n2952) );
  NAND3_X2 U9355 ( .A1(n6856), .A2(n6851), .A3(n6852), .ZN(n16365) );
  AOI21_X1 U9358 ( .B1(n7451), .B2(n7452), .A(n8297), .ZN(n3445) );
  OR2_X1 U9360 ( .A1(n10726), .A2(n10924), .ZN(n10459) );
  OR2_X1 U9361 ( .A1(n1899), .A2(n7291), .ZN(n7332) );
  NAND2_X1 U9364 ( .A1(n6729), .A2(n20324), .ZN(n2956) );
  XOR2_X1 U9365 ( .A(n12432), .B(n12433), .Z(n4510) );
  XNOR2_X1 U9366 ( .A(n4360), .B(n16480), .ZN(n15779) );
  OAI21_X2 U9368 ( .B1(n23582), .B2(n23583), .A(n23581), .ZN(n24757) );
  NAND2_X1 U9369 ( .A1(n2958), .A2(n2957), .ZN(n14990) );
  NAND2_X1 U9370 ( .A1(n13682), .A2(n28806), .ZN(n2957) );
  NAND2_X1 U9371 ( .A1(n13683), .A2(n2959), .ZN(n2958) );
  NOR2_X1 U9372 ( .A1(n6565), .A2(n20433), .ZN(n6564) );
  NAND2_X1 U9373 ( .A1(n23799), .A2(n23793), .ZN(n23495) );
  NOR2_X1 U9374 ( .A1(n1938), .A2(n7675), .ZN(n5256) );
  XNOR2_X1 U9375 ( .A(n22771), .B(n22297), .ZN(n6837) );
  NAND2_X1 U9376 ( .A1(n1926), .A2(n15012), .ZN(n6333) );
  NAND4_X2 U9377 ( .A1(n4234), .A2(n4233), .A3(n6154), .A4(n6153), .ZN(n24756)
         );
  XNOR2_X1 U9379 ( .A(n15796), .B(n3813), .ZN(n3937) );
  XNOR2_X1 U9380 ( .A(n13248), .B(n12850), .ZN(n2962) );
  NAND3_X1 U9381 ( .A1(n7384), .A2(n7708), .A3(n7382), .ZN(n2963) );
  NAND2_X1 U9382 ( .A1(n12049), .A2(n12053), .ZN(n12057) );
  OR3_X1 U9383 ( .A1(n11951), .A2(n11943), .A3(n3946), .ZN(n10952) );
  OR2_X1 U9385 ( .A1(n13677), .A2(n12743), .ZN(n14471) );
  NAND2_X1 U9386 ( .A1(n2965), .A2(n2964), .ZN(n14496) );
  NAND2_X1 U9387 ( .A1(n2967), .A2(n9531), .ZN(n6405) );
  OAI21_X1 U9388 ( .B1(n5396), .B2(n8320), .A(n8749), .ZN(n2967) );
  OAI21_X1 U9389 ( .B1(n14101), .B2(n14230), .A(n3645), .ZN(n14595) );
  INV_X1 U9391 ( .A(n11136), .ZN(n2968) );
  NAND2_X1 U9392 ( .A1(n11135), .A2(n11140), .ZN(n10918) );
  NAND3_X1 U9393 ( .A1(n18018), .A2(n17564), .A3(n18017), .ZN(n17773) );
  NAND2_X1 U9395 ( .A1(n7309), .A2(n7306), .ZN(n7307) );
  NAND2_X1 U9396 ( .A1(n18150), .A2(n1894), .ZN(n3468) );
  NAND2_X1 U9397 ( .A1(n11708), .A2(n11417), .ZN(n11415) );
  OAI211_X1 U9399 ( .C1(n14181), .C2(n2972), .A(n190), .B(n2970), .ZN(n2969)
         );
  INV_X1 U9400 ( .A(n10809), .ZN(n6347) );
  NOR2_X1 U9403 ( .A1(n7982), .A2(n7981), .ZN(n7648) );
  XNOR2_X1 U9404 ( .A(n9003), .B(n9094), .ZN(n5924) );
  NAND2_X1 U9406 ( .A1(n8492), .A2(n2977), .ZN(n8004) );
  NAND2_X1 U9407 ( .A1(n20304), .A2(n2978), .ZN(n20120) );
  OAI21_X2 U9408 ( .B1(n11388), .B2(n11387), .A(n11386), .ZN(n4253) );
  NOR2_X1 U9409 ( .A1(n20894), .A2(n20895), .ZN(n5830) );
  NAND2_X1 U9410 ( .A1(n8735), .A2(n2983), .ZN(n8736) );
  NAND2_X1 U9411 ( .A1(n8741), .A2(n9073), .ZN(n8617) );
  NAND2_X1 U9412 ( .A1(n3149), .A2(n3150), .ZN(n22948) );
  NAND4_X2 U9413 ( .A1(n11993), .A2(n11994), .A3(n11992), .A4(n11991), .ZN(
        n13028) );
  NAND3_X1 U9414 ( .A1(n24520), .A2(n24516), .A3(n24421), .ZN(n3359) );
  OAI21_X1 U9415 ( .B1(n5625), .B2(n28471), .A(n4751), .ZN(n4750) );
  OAI211_X1 U9416 ( .C1(n17265), .C2(n16992), .A(n16996), .B(n2985), .ZN(
        n16998) );
  XNOR2_X1 U9417 ( .A(n9952), .B(n9951), .ZN(n5316) );
  OR2_X1 U9418 ( .A1(n20612), .A2(n29508), .ZN(n4682) );
  INV_X1 U9419 ( .A(n11877), .ZN(n11453) );
  NAND2_X1 U9421 ( .A1(n7939), .A2(n7400), .ZN(n8298) );
  NAND2_X1 U9422 ( .A1(n21655), .A2(n2989), .ZN(n2988) );
  NAND3_X1 U9423 ( .A1(n21072), .A2(n21073), .A3(n2992), .ZN(n2991) );
  INV_X1 U9424 ( .A(n18242), .ZN(n4725) );
  OR2_X1 U9425 ( .A1(n22991), .A2(n23640), .ZN(n22256) );
  OAI21_X1 U9426 ( .B1(n29315), .B2(n29146), .A(n2994), .ZN(n18574) );
  NAND2_X1 U9427 ( .A1(n29146), .A2(n20081), .ZN(n2994) );
  XNOR2_X2 U9428 ( .A(n7037), .B(Key[150]), .ZN(n7456) );
  INV_X1 U9429 ( .A(n20658), .ZN(n21750) );
  INV_X1 U9430 ( .A(n24809), .ZN(n24499) );
  OAI211_X2 U9431 ( .C1(n19731), .C2(n20117), .A(n4682), .B(n4683), .ZN(n21811) );
  OR2_X1 U9432 ( .A1(n17565), .A2(n4316), .ZN(n17040) );
  INV_X1 U9433 ( .A(n21374), .ZN(n21375) );
  XNOR2_X1 U9434 ( .A(n28433), .B(n1119), .ZN(n24847) );
  NAND2_X1 U9436 ( .A1(n3001), .A2(n2999), .ZN(n24208) );
  NAND2_X1 U9437 ( .A1(n220), .A2(n24817), .ZN(n2999) );
  XNOR2_X1 U9438 ( .A(n6100), .B(n22056), .ZN(n23702) );
  NOR2_X1 U9439 ( .A1(n5706), .A2(n10777), .ZN(n5705) );
  OR2_X1 U9440 ( .A1(n7508), .A2(n7514), .ZN(n7132) );
  NOR2_X2 U9441 ( .A1(n17343), .A2(n3002), .ZN(n18707) );
  NAND2_X1 U9442 ( .A1(n2069), .A2(n17341), .ZN(n3002) );
  NAND2_X1 U9443 ( .A1(n21085), .A2(n20804), .ZN(n20805) );
  NAND2_X1 U9444 ( .A1(n24242), .A2(n24635), .ZN(n24192) );
  NAND3_X1 U9445 ( .A1(n23808), .A2(n22742), .A3(n28653), .ZN(n3337) );
  NOR2_X1 U9446 ( .A1(n384), .A2(n20239), .ZN(n3005) );
  OAI21_X1 U9448 ( .B1(n18539), .B2(n18535), .A(n3006), .ZN(n17700) );
  NAND2_X1 U9449 ( .A1(n18539), .A2(n17864), .ZN(n3006) );
  NAND2_X1 U9450 ( .A1(n5616), .A2(n14349), .ZN(n14015) );
  NOR2_X1 U9451 ( .A1(n19895), .A2(n19896), .ZN(n3009) );
  XNOR2_X1 U9452 ( .A(n4764), .B(n29154), .ZN(n24877) );
  INV_X1 U9454 ( .A(n14952), .ZN(n14949) );
  NAND2_X1 U9455 ( .A1(n15077), .A2(n14948), .ZN(n14952) );
  NAND3_X1 U9456 ( .A1(n3461), .A2(n3460), .A3(n9914), .ZN(n11390) );
  INV_X1 U9457 ( .A(n3011), .ZN(n3010) );
  MUX2_X1 U9458 ( .A(n11927), .B(n11392), .S(n11391), .Z(n11393) );
  NAND2_X1 U9459 ( .A1(n11921), .A2(n11853), .ZN(n11391) );
  NAND2_X1 U9460 ( .A1(n10726), .A2(n10924), .ZN(n10051) );
  NOR2_X2 U9461 ( .A1(n3014), .A2(n11089), .ZN(n12578) );
  AOI21_X1 U9462 ( .B1(n11081), .B2(n11082), .A(n433), .ZN(n3014) );
  OR2_X1 U9463 ( .A1(n8741), .A2(n9073), .ZN(n8859) );
  INV_X1 U9464 ( .A(n14863), .ZN(n15369) );
  XNOR2_X1 U9465 ( .A(n25508), .B(n25322), .ZN(n26107) );
  INV_X1 U9466 ( .A(n4166), .ZN(n13827) );
  XNOR2_X1 U9468 ( .A(n9779), .B(n9446), .ZN(n10148) );
  NAND2_X1 U9469 ( .A1(n3017), .A2(n4706), .ZN(n18171) );
  XNOR2_X1 U9470 ( .A(n4669), .B(n13260), .ZN(n12966) );
  NAND2_X1 U9472 ( .A1(n3019), .A2(n21599), .ZN(n21319) );
  NAND2_X1 U9473 ( .A1(n28442), .A2(n21601), .ZN(n3019) );
  NAND3_X1 U9474 ( .A1(n4443), .A2(n11512), .A3(n12035), .ZN(n3020) );
  OAI22_X1 U9475 ( .A1(n10933), .A2(n1879), .B1(n10932), .B2(n10931), .ZN(
        n5905) );
  NAND3_X1 U9476 ( .A1(n8187), .A2(n8186), .A3(n8562), .ZN(n8190) );
  NAND2_X1 U9477 ( .A1(n15089), .A2(n3022), .ZN(n15092) );
  NAND2_X1 U9478 ( .A1(n10725), .A2(n10724), .ZN(n3023) );
  OAI211_X2 U9479 ( .C1(n21415), .C2(n21414), .A(n3025), .B(n3024), .ZN(n22473) );
  NAND2_X1 U9480 ( .A1(n21413), .A2(n4937), .ZN(n3024) );
  NAND2_X1 U9481 ( .A1(n21411), .A2(n21412), .ZN(n3025) );
  NAND2_X1 U9483 ( .A1(n23159), .A2(n23512), .ZN(n3026) );
  NOR2_X1 U9484 ( .A1(n11108), .A2(n3027), .ZN(n11109) );
  INV_X1 U9485 ( .A(n11942), .ZN(n3027) );
  NAND2_X1 U9486 ( .A1(n12271), .A2(n28202), .ZN(n11942) );
  NAND2_X1 U9488 ( .A1(n3205), .A2(n4662), .ZN(n3028) );
  OAI21_X1 U9489 ( .B1(n13612), .B2(n13611), .A(n14261), .ZN(n3346) );
  OAI211_X2 U9493 ( .C1(n8352), .C2(n8431), .A(n8060), .B(n8059), .ZN(n10071)
         );
  NOR2_X1 U9494 ( .A1(n26560), .A2(n28578), .ZN(n3032) );
  NAND2_X1 U9495 ( .A1(n26460), .A2(n28578), .ZN(n3033) );
  NAND3_X1 U9496 ( .A1(n8018), .A2(n7744), .A3(n7745), .ZN(n7247) );
  NOR2_X1 U9498 ( .A1(n15462), .A2(n15464), .ZN(n13889) );
  NAND2_X1 U9500 ( .A1(n10745), .A2(n4945), .ZN(n11636) );
  XNOR2_X1 U9501 ( .A(n3037), .B(n22471), .ZN(n23391) );
  XNOR2_X1 U9502 ( .A(n22469), .B(n22470), .ZN(n3037) );
  NAND2_X1 U9503 ( .A1(n17508), .A2(n17505), .ZN(n16728) );
  BUF_X1 U9505 ( .A(n25268), .Z(n25513) );
  AND2_X1 U9506 ( .A1(n26682), .A2(n27433), .ZN(n26833) );
  OR2_X1 U9507 ( .A1(n24117), .A2(n24433), .ZN(n24118) );
  OR2_X1 U9508 ( .A1(n23261), .A2(n23712), .ZN(n22972) );
  INV_X1 U9509 ( .A(n17872), .ZN(n17937) );
  OR2_X1 U9510 ( .A1(n21412), .A2(n20663), .ZN(n21415) );
  NAND3_X1 U9511 ( .A1(n16970), .A2(n16969), .A3(n3038), .ZN(n16972) );
  NOR2_X1 U9512 ( .A1(n13693), .A2(n29607), .ZN(n4610) );
  INV_X1 U9513 ( .A(n23290), .ZN(n23441) );
  AND2_X1 U9515 ( .A1(n24583), .A2(n29026), .ZN(n6056) );
  INV_X1 U9517 ( .A(n17438), .ZN(n17434) );
  INV_X1 U9518 ( .A(n16980), .ZN(n4002) );
  XNOR2_X1 U9519 ( .A(n3092), .B(n3091), .ZN(n22598) );
  OAI211_X1 U9520 ( .C1(n20493), .C2(n20496), .A(n3040), .B(n5225), .ZN(n5305)
         );
  NAND2_X1 U9521 ( .A1(n3041), .A2(n29616), .ZN(n3040) );
  INV_X1 U9522 ( .A(n20494), .ZN(n3041) );
  INV_X1 U9523 ( .A(n13060), .ZN(n14127) );
  INV_X1 U9524 ( .A(n18285), .ZN(n17859) );
  NAND2_X1 U9525 ( .A1(n28653), .A2(n23284), .ZN(n3042) );
  OR2_X1 U9526 ( .A1(n23809), .A2(n23806), .ZN(n3043) );
  XNOR2_X1 U9529 ( .A(n3044), .B(n13441), .ZN(n12048) );
  XNOR2_X1 U9530 ( .A(n12034), .B(n13167), .ZN(n3044) );
  NAND2_X1 U9531 ( .A1(n7565), .A2(n7562), .ZN(n7124) );
  INV_X1 U9532 ( .A(n14414), .ZN(n14216) );
  NAND2_X1 U9534 ( .A1(n555), .A2(n14414), .ZN(n3045) );
  NAND2_X1 U9536 ( .A1(n585), .A2(n11284), .ZN(n3046) );
  NAND2_X1 U9537 ( .A1(n11029), .A2(n10884), .ZN(n3047) );
  OAI211_X2 U9538 ( .C1(n18002), .C2(n18337), .A(n1973), .B(n3048), .ZN(n19427) );
  NAND2_X1 U9539 ( .A1(n18001), .A2(n18337), .ZN(n3048) );
  OAI21_X1 U9540 ( .B1(n5870), .B2(n8523), .A(n8524), .ZN(n3679) );
  NAND2_X1 U9544 ( .A1(n8748), .A2(n8751), .ZN(n3051) );
  NAND2_X1 U9545 ( .A1(n3052), .A2(n23713), .ZN(n23237) );
  NAND2_X1 U9546 ( .A1(n23261), .A2(n23587), .ZN(n3052) );
  NAND2_X1 U9547 ( .A1(n3053), .A2(n23057), .ZN(n6439) );
  OAI22_X1 U9548 ( .A1(n23426), .A2(n28122), .B1(n23428), .B2(n29108), .ZN(
        n3053) );
  NOR2_X2 U9550 ( .A1(n4114), .A2(n11603), .ZN(n6683) );
  OAI22_X1 U9551 ( .A1(n11340), .A2(n11338), .B1(n11175), .B2(n11345), .ZN(
        n6289) );
  NAND2_X1 U9552 ( .A1(n3055), .A2(n29470), .ZN(n23509) );
  INV_X1 U9553 ( .A(n23507), .ZN(n3055) );
  NAND2_X1 U9554 ( .A1(n24388), .A2(n24387), .ZN(n23507) );
  INV_X1 U9555 ( .A(n12244), .ZN(n5839) );
  NAND3_X1 U9556 ( .A1(n10570), .A2(n11068), .A3(n10571), .ZN(n11901) );
  XNOR2_X1 U9558 ( .A(n12529), .B(n13563), .ZN(n10538) );
  INV_X1 U9559 ( .A(n5593), .ZN(n5592) );
  XNOR2_X1 U9560 ( .A(n19438), .B(n18988), .ZN(n3912) );
  NAND3_X1 U9561 ( .A1(n12360), .A2(n12358), .A3(n6552), .ZN(n6551) );
  NOR2_X2 U9562 ( .A1(n17112), .A2(n17111), .ZN(n17847) );
  NAND2_X1 U9563 ( .A1(n11021), .A2(n3058), .ZN(n13371) );
  NAND3_X1 U9564 ( .A1(n14221), .A2(n5777), .A3(n14222), .ZN(n16510) );
  NAND2_X1 U9565 ( .A1(n3061), .A2(n3060), .ZN(n3059) );
  INV_X1 U9566 ( .A(n24030), .ZN(n3060) );
  NAND2_X1 U9567 ( .A1(n6501), .A2(n4295), .ZN(n6500) );
  NAND2_X1 U9568 ( .A1(n13852), .A2(n14184), .ZN(n14470) );
  NAND3_X1 U9569 ( .A1(n8536), .A2(n8384), .A3(n8730), .ZN(n7187) );
  NAND2_X1 U9570 ( .A1(n6466), .A2(n14217), .ZN(n14417) );
  NAND2_X1 U9571 ( .A1(n26637), .A2(n29092), .ZN(n3063) );
  NAND2_X1 U9572 ( .A1(n27970), .A2(n26636), .ZN(n3064) );
  NAND2_X1 U9573 ( .A1(n7851), .A2(n7708), .ZN(n7856) );
  INV_X1 U9575 ( .A(n10717), .ZN(n6479) );
  INV_X1 U9576 ( .A(n21536), .ZN(n20793) );
  NAND2_X1 U9577 ( .A1(n21514), .A2(n21199), .ZN(n21536) );
  NAND2_X1 U9578 ( .A1(n3065), .A2(n27514), .ZN(n27518) );
  NOR2_X1 U9579 ( .A1(n27513), .A2(n27516), .ZN(n3065) );
  NAND3_X1 U9580 ( .A1(n6435), .A2(n26917), .A3(n3066), .ZN(n6437) );
  INV_X1 U9581 ( .A(n27520), .ZN(n27523) );
  XNOR2_X1 U9582 ( .A(n25521), .B(n25069), .ZN(n4810) );
  NAND2_X1 U9583 ( .A1(n21210), .A2(n21209), .ZN(n22026) );
  NAND2_X1 U9584 ( .A1(n11922), .A2(n11852), .ZN(n3410) );
  NAND2_X1 U9587 ( .A1(n14268), .A2(n14262), .ZN(n3072) );
  INV_X1 U9588 ( .A(n9577), .ZN(n10192) );
  XNOR2_X1 U9589 ( .A(n9577), .B(n3073), .ZN(n9818) );
  OR2_X1 U9590 ( .A1(n11819), .A2(n12198), .ZN(n12127) );
  NAND2_X1 U9591 ( .A1(n12041), .A2(n12042), .ZN(n10643) );
  NAND2_X1 U9593 ( .A1(n5498), .A2(n24364), .ZN(n5501) );
  OAI211_X1 U9594 ( .C1(n17902), .C2(n18111), .A(n18110), .B(n17798), .ZN(
        n3074) );
  OAI21_X1 U9595 ( .B1(n7321), .B2(n7116), .A(n7768), .ZN(n5244) );
  NAND3_X1 U9596 ( .A1(n27288), .A2(n27275), .A3(n27287), .ZN(n3146) );
  INV_X1 U9598 ( .A(n3078), .ZN(n3077) );
  OAI21_X1 U9599 ( .B1(n5635), .B2(n3080), .A(n3079), .ZN(n15181) );
  AOI21_X2 U9600 ( .B1(n11561), .B2(n11562), .A(n11560), .ZN(n13190) );
  XNOR2_X2 U9601 ( .A(n12903), .B(n12902), .ZN(n14084) );
  NAND3_X1 U9602 ( .A1(n2014), .A2(n6322), .A3(n6323), .ZN(n26652) );
  AOI22_X1 U9603 ( .A1(n26653), .A2(n27548), .B1(n27541), .B2(n27547), .ZN(
        n26654) );
  OAI22_X1 U9604 ( .A1(n19032), .A2(n20232), .B1(n383), .B2(n20231), .ZN(n5274) );
  NOR2_X1 U9605 ( .A1(n20956), .A2(n20957), .ZN(n3280) );
  NAND2_X1 U9606 ( .A1(n5207), .A2(n14243), .ZN(n3082) );
  NAND2_X1 U9608 ( .A1(n17577), .A2(n18251), .ZN(n3085) );
  INV_X1 U9610 ( .A(n4515), .ZN(n14802) );
  NAND3_X2 U9611 ( .A1(n13875), .A2(n13876), .A3(n5015), .ZN(n4515) );
  NAND2_X1 U9612 ( .A1(n25994), .A2(n27371), .ZN(n25995) );
  NAND2_X1 U9613 ( .A1(n14167), .A2(n14169), .ZN(n6744) );
  NAND2_X1 U9614 ( .A1(n8081), .A2(n8336), .ZN(n8506) );
  INV_X1 U9615 ( .A(n21645), .ZN(n4659) );
  NAND2_X1 U9616 ( .A1(n2057), .A2(n424), .ZN(n3090) );
  NAND3_X1 U9617 ( .A1(n8277), .A2(n8279), .A3(n8278), .ZN(n3094) );
  NAND2_X1 U9619 ( .A1(n21216), .A2(n21000), .ZN(n20998) );
  NAND2_X1 U9620 ( .A1(n3095), .A2(n7967), .ZN(n4698) );
  OAI21_X1 U9621 ( .B1(n7963), .B2(n1938), .A(n7236), .ZN(n3095) );
  AND3_X1 U9622 ( .A1(n3541), .A2(n3481), .A3(n24588), .ZN(n5863) );
  OR2_X1 U9623 ( .A1(n10093), .A2(n11152), .ZN(n3165) );
  NAND2_X1 U9624 ( .A1(n5332), .A2(n2205), .ZN(n24637) );
  NAND2_X1 U9625 ( .A1(n5576), .A2(n3583), .ZN(n15535) );
  NAND2_X1 U9626 ( .A1(n18034), .A2(n18154), .ZN(n4854) );
  XNOR2_X1 U9627 ( .A(n13505), .B(n13134), .ZN(n3097) );
  NAND3_X2 U9628 ( .A1(n3668), .A2(n5371), .A3(n3667), .ZN(n13451) );
  NOR2_X1 U9630 ( .A1(n6374), .A2(n10863), .ZN(n6372) );
  NAND2_X1 U9631 ( .A1(n3100), .A2(n3099), .ZN(n17122) );
  AOI21_X1 U9633 ( .B1(n10686), .B2(n9362), .A(n6775), .ZN(n6774) );
  INV_X1 U9634 ( .A(n4852), .ZN(n16654) );
  NOR2_X2 U9635 ( .A1(n17257), .A2(n17256), .ZN(n18240) );
  OR2_X2 U9636 ( .A1(n12091), .A2(n12092), .ZN(n11856) );
  NAND2_X1 U9637 ( .A1(n14310), .A2(n14309), .ZN(n13888) );
  NAND2_X1 U9639 ( .A1(n3106), .A2(n3105), .ZN(n10818) );
  NAND2_X1 U9640 ( .A1(n10815), .A2(n28207), .ZN(n3105) );
  NAND2_X1 U9641 ( .A1(n3107), .A2(n28157), .ZN(n3106) );
  OAI21_X1 U9642 ( .B1(n28638), .B2(n3585), .A(n3584), .ZN(n3107) );
  NOR2_X1 U9643 ( .A1(n24368), .A2(n24367), .ZN(n24303) );
  INV_X1 U9645 ( .A(n15175), .ZN(n15459) );
  OR2_X1 U9646 ( .A1(n572), .A2(n11754), .ZN(n11477) );
  OR2_X1 U9647 ( .A1(n21936), .A2(n21935), .ZN(n21937) );
  INV_X1 U9648 ( .A(n21424), .ZN(n5000) );
  AND2_X1 U9649 ( .A1(n3922), .A2(n14893), .ZN(n12011) );
  XNOR2_X1 U9650 ( .A(n12849), .B(n12554), .ZN(n13332) );
  INV_X1 U9651 ( .A(n6482), .ZN(n4744) );
  OAI21_X1 U9653 ( .B1(n15169), .B2(n6925), .A(n1850), .ZN(n14553) );
  INV_X1 U9654 ( .A(n23765), .ZN(n23766) );
  XNOR2_X1 U9655 ( .A(n6416), .B(n6415), .ZN(n17272) );
  INV_X1 U9656 ( .A(n24397), .ZN(n24323) );
  INV_X1 U9657 ( .A(n23655), .ZN(n24793) );
  XNOR2_X1 U9658 ( .A(n3913), .B(n19584), .ZN(n18988) );
  INV_X1 U9659 ( .A(n22735), .ZN(n6119) );
  AOI21_X1 U9660 ( .B1(n28916), .B2(n21089), .A(n21930), .ZN(n3560) );
  XNOR2_X1 U9661 ( .A(n29035), .B(n19323), .ZN(n19693) );
  NOR2_X1 U9662 ( .A1(n8521), .A2(n8811), .ZN(n5869) );
  AOI21_X1 U9663 ( .B1(n28638), .B2(n10563), .A(n11196), .ZN(n6272) );
  NAND3_X1 U9664 ( .A1(n12508), .A2(n3108), .A3(n10863), .ZN(n11835) );
  INV_X1 U9666 ( .A(n26769), .ZN(n6768) );
  NAND2_X1 U9667 ( .A1(n296), .A2(n18972), .ZN(n5106) );
  INV_X1 U9668 ( .A(n15642), .ZN(n16425) );
  NAND3_X1 U9669 ( .A1(n7673), .A2(n7481), .A3(n8281), .ZN(n7482) );
  OR2_X1 U9670 ( .A1(n7851), .A2(n7384), .ZN(n7383) );
  AND2_X1 U9671 ( .A1(n14435), .A2(n14207), .ZN(n13957) );
  XNOR2_X1 U9672 ( .A(n12847), .B(n12848), .ZN(n3110) );
  XNOR2_X1 U9674 ( .A(n19263), .B(n19639), .ZN(n3111) );
  XNOR2_X1 U9675 ( .A(n9491), .B(n9492), .ZN(n6135) );
  NAND2_X1 U9676 ( .A1(n11255), .A2(n11315), .ZN(n3113) );
  NAND2_X1 U9679 ( .A1(n3895), .A2(n3896), .ZN(n5682) );
  XNOR2_X2 U9680 ( .A(n19107), .B(n19106), .ZN(n20488) );
  NAND3_X1 U9681 ( .A1(n8890), .A2(n8507), .A3(n8886), .ZN(n8508) );
  NAND3_X1 U9683 ( .A1(n3118), .A2(n8210), .A3(n3117), .ZN(n8838) );
  NAND2_X1 U9684 ( .A1(n3159), .A2(n8209), .ZN(n3118) );
  INV_X1 U9689 ( .A(n9431), .ZN(n9678) );
  AND2_X1 U9690 ( .A1(n20786), .A2(n21097), .ZN(n20799) );
  AOI21_X1 U9691 ( .B1(n3123), .B2(n7829), .A(n8205), .ZN(n7435) );
  NAND2_X1 U9692 ( .A1(n8201), .A2(n7828), .ZN(n3123) );
  AND2_X1 U9693 ( .A1(n24794), .A2(n28512), .ZN(n3124) );
  NAND2_X1 U9694 ( .A1(n16806), .A2(n17259), .ZN(n16669) );
  INV_X1 U9695 ( .A(n26746), .ZN(n5760) );
  NAND2_X1 U9697 ( .A1(n3125), .A2(n14322), .ZN(n14066) );
  NAND3_X1 U9698 ( .A1(n15294), .A2(n15293), .A3(n15291), .ZN(n14838) );
  OR2_X1 U9699 ( .A1(n13909), .A2(n14047), .ZN(n5730) );
  NAND2_X1 U9700 ( .A1(n6661), .A2(n12004), .ZN(n11686) );
  NOR2_X2 U9701 ( .A1(n10567), .A2(n10566), .ZN(n12004) );
  XNOR2_X1 U9702 ( .A(n6453), .B(n15978), .ZN(n6455) );
  OR2_X1 U9703 ( .A1(n21736), .A2(n29314), .ZN(n21477) );
  NAND2_X1 U9704 ( .A1(n3375), .A2(n14359), .ZN(n13032) );
  NAND3_X1 U9705 ( .A1(n8286), .A2(n7913), .A3(n7914), .ZN(n7918) );
  INV_X1 U9706 ( .A(n23658), .ZN(n5773) );
  INV_X1 U9707 ( .A(n13902), .ZN(n4425) );
  AND2_X1 U9708 ( .A1(n15361), .A2(n4992), .ZN(n14753) );
  NAND3_X1 U9709 ( .A1(n9234), .A2(n9235), .A3(n9233), .ZN(n9236) );
  NAND2_X1 U9710 ( .A1(n20105), .A2(n3126), .ZN(n20933) );
  INV_X1 U9711 ( .A(n7426), .ZN(n6993) );
  INV_X1 U9712 ( .A(n17864), .ZN(n18536) );
  OR2_X1 U9713 ( .A1(n27056), .A2(n26850), .ZN(n27055) );
  OR2_X1 U9714 ( .A1(n14771), .A2(n14770), .ZN(n3638) );
  OR2_X1 U9715 ( .A1(n23010), .A2(n6227), .ZN(n23140) );
  INV_X1 U9716 ( .A(n17957), .ZN(n4905) );
  OAI21_X1 U9717 ( .B1(n8658), .B2(n8654), .A(n8503), .ZN(n3127) );
  INV_X1 U9718 ( .A(n581), .ZN(n5914) );
  NAND2_X1 U9720 ( .A1(n10750), .A2(n11198), .ZN(n3130) );
  NAND2_X1 U9721 ( .A1(n20832), .A2(n3131), .ZN(n22718) );
  OR2_X1 U9722 ( .A1(n7308), .A2(n7093), .ZN(n7863) );
  AND2_X1 U9723 ( .A1(n28197), .A2(n15361), .ZN(n14750) );
  INV_X1 U9724 ( .A(n14922), .ZN(n6699) );
  AND2_X1 U9725 ( .A1(n10797), .A2(n11225), .ZN(n10621) );
  INV_X1 U9726 ( .A(n19554), .ZN(n19927) );
  AND2_X1 U9727 ( .A1(n28207), .A2(n10814), .ZN(n6677) );
  NAND3_X1 U9728 ( .A1(n349), .A2(n12252), .A3(n12253), .ZN(n3553) );
  INV_X1 U9730 ( .A(n20148), .ZN(n20102) );
  INV_X1 U9733 ( .A(n18011), .ZN(n18477) );
  NAND3_X1 U9735 ( .A1(n3137), .A2(n5854), .A3(n4877), .ZN(n3136) );
  INV_X1 U9736 ( .A(n20038), .ZN(n3137) );
  NOR2_X1 U9738 ( .A1(n4044), .A2(n17780), .ZN(n17783) );
  XNOR2_X1 U9739 ( .A(n22173), .B(n22483), .ZN(n23261) );
  INV_X1 U9741 ( .A(n3441), .ZN(n5709) );
  INV_X1 U9742 ( .A(n15265), .ZN(n15499) );
  NOR2_X1 U9744 ( .A1(n5584), .A2(n14331), .ZN(n14410) );
  OAI21_X1 U9745 ( .B1(n14410), .B2(n14409), .A(n14408), .ZN(n4001) );
  NOR2_X1 U9746 ( .A1(n24293), .A2(n24533), .ZN(n24892) );
  XNOR2_X1 U9747 ( .A(n25711), .B(n25713), .ZN(n3168) );
  OAI21_X1 U9748 ( .B1(n12075), .B2(n5974), .A(n5973), .ZN(n5972) );
  XNOR2_X1 U9749 ( .A(n18779), .B(n18991), .ZN(n18499) );
  XNOR2_X1 U9750 ( .A(n16279), .B(n3138), .ZN(n16370) );
  NAND2_X1 U9751 ( .A1(n17547), .A2(n4624), .ZN(n4623) );
  NAND2_X1 U9752 ( .A1(n4626), .A2(n4625), .ZN(n17547) );
  NAND3_X1 U9753 ( .A1(n6875), .A2(n9176), .A3(n8983), .ZN(n3140) );
  OAI21_X2 U9755 ( .B1(n8917), .B2(n8674), .A(n8673), .ZN(n10257) );
  XNOR2_X1 U9757 ( .A(n9272), .B(n10148), .ZN(n3141) );
  INV_X1 U9758 ( .A(n28523), .ZN(n24027) );
  OAI211_X2 U9759 ( .C1(n11408), .C2(n11645), .A(n3143), .B(n3142), .ZN(n13405) );
  NAND2_X1 U9760 ( .A1(n12142), .A2(n11715), .ZN(n3142) );
  AOI21_X1 U9762 ( .B1(n20336), .B2(n20625), .A(n20623), .ZN(n3144) );
  INV_X1 U9763 ( .A(n20889), .ZN(n5205) );
  OAI22_X1 U9764 ( .A1(n20643), .A2(n20905), .B1(n21605), .B2(n21599), .ZN(
        n3145) );
  XNOR2_X2 U9765 ( .A(n16502), .B(n16501), .ZN(n16797) );
  NAND3_X1 U9766 ( .A1(n3998), .A2(n3999), .A3(n11750), .ZN(n4000) );
  OAI21_X1 U9767 ( .B1(n27285), .B2(n27291), .A(n3146), .ZN(n27252) );
  NOR2_X1 U9768 ( .A1(n23513), .A2(n339), .ZN(n3147) );
  NAND2_X1 U9770 ( .A1(n12037), .A2(n12158), .ZN(n4443) );
  NOR2_X1 U9771 ( .A1(n17927), .A2(n18301), .ZN(n17929) );
  NAND2_X1 U9772 ( .A1(n19764), .A2(n5424), .ZN(n18847) );
  OAI22_X1 U9773 ( .A1(n20048), .A2(n19761), .B1(n18892), .B2(n20049), .ZN(
        n5424) );
  NOR2_X1 U9775 ( .A1(n21291), .A2(n21290), .ZN(n20913) );
  NAND2_X1 U9776 ( .A1(n29564), .A2(n23827), .ZN(n22944) );
  NAND2_X1 U9777 ( .A1(n22945), .A2(n23741), .ZN(n3150) );
  XNOR2_X1 U9778 ( .A(n9685), .B(n6440), .ZN(n4590) );
  XNOR2_X1 U9779 ( .A(n3151), .B(n624), .ZN(Ciphertext[111]) );
  OAI211_X1 U9780 ( .C1(n26893), .C2(n26894), .A(n26891), .B(n26892), .ZN(
        n3151) );
  NAND2_X1 U9782 ( .A1(n14518), .A2(n15217), .ZN(n14837) );
  XNOR2_X2 U9783 ( .A(n16268), .B(n16267), .ZN(n17487) );
  NAND2_X1 U9785 ( .A1(n803), .A2(n24803), .ZN(n24261) );
  NAND2_X1 U9786 ( .A1(n14767), .A2(n14810), .ZN(n13924) );
  NAND4_X2 U9788 ( .A1(n8833), .A2(n8834), .A3(n8832), .A4(n8831), .ZN(n9941)
         );
  OAI21_X2 U9789 ( .B1(n29119), .B2(n8137), .A(n4940), .ZN(n8981) );
  NAND2_X1 U9790 ( .A1(n1834), .A2(n10713), .ZN(n6152) );
  OR3_X1 U9791 ( .A1(n29083), .A2(n16541), .A3(n17456), .ZN(n16542) );
  NOR2_X1 U9792 ( .A1(n30), .A2(n14400), .ZN(n4010) );
  NAND2_X1 U9795 ( .A1(n5724), .A2(n5726), .ZN(n5721) );
  INV_X1 U9796 ( .A(n18301), .ZN(n3153) );
  NAND2_X1 U9797 ( .A1(n17278), .A2(n17277), .ZN(n16767) );
  NAND2_X1 U9798 ( .A1(n10528), .A2(n11047), .ZN(n11264) );
  AOI21_X1 U9800 ( .B1(n7210), .B2(n7211), .A(n8264), .ZN(n3155) );
  NAND2_X1 U9801 ( .A1(n29395), .A2(n9530), .ZN(n3157) );
  OR2_X1 U9802 ( .A1(n18919), .A2(n21091), .ZN(n4876) );
  OR2_X1 U9803 ( .A1(n14398), .A2(n14401), .ZN(n14210) );
  NAND2_X1 U9804 ( .A1(n11112), .A2(n11111), .ZN(n3509) );
  NAND2_X1 U9805 ( .A1(n29546), .A2(n17355), .ZN(n17358) );
  OR2_X2 U9806 ( .A1(n11663), .A2(n11664), .ZN(n13444) );
  AOI21_X2 U9807 ( .B1(n23195), .B2(n23470), .A(n3158), .ZN(n24559) );
  NAND2_X1 U9808 ( .A1(n370), .A2(n8208), .ZN(n3159) );
  INV_X1 U9809 ( .A(n5316), .ZN(n11111) );
  INV_X1 U9810 ( .A(n22026), .ZN(n22288) );
  OR2_X1 U9811 ( .A1(n14045), .A2(n14046), .ZN(n5064) );
  NAND2_X1 U9812 ( .A1(n3162), .A2(n3160), .ZN(n11473) );
  NAND3_X1 U9813 ( .A1(n3636), .A2(n10477), .A3(n3161), .ZN(n3160) );
  NAND2_X1 U9814 ( .A1(n10479), .A2(n11350), .ZN(n3162) );
  INV_X1 U9816 ( .A(n23228), .ZN(n3432) );
  NOR2_X1 U9817 ( .A1(n14842), .A2(n14695), .ZN(n14060) );
  OAI22_X1 U9818 ( .A1(n1076), .A2(n26426), .B1(n26431), .B2(n26425), .ZN(
        n26276) );
  NAND2_X1 U9819 ( .A1(n10696), .A2(n10989), .ZN(n3801) );
  OAI21_X1 U9820 ( .B1(n27121), .B2(n27122), .A(n3456), .ZN(n27128) );
  NAND3_X1 U9821 ( .A1(n7706), .A2(n3163), .A3(n371), .ZN(n4159) );
  NAND2_X1 U9822 ( .A1(n7705), .A2(n7852), .ZN(n3163) );
  INV_X1 U9823 ( .A(n29647), .ZN(n18509) );
  NOR2_X1 U9824 ( .A1(n5265), .A2(n28608), .ZN(n5264) );
  NAND3_X2 U9825 ( .A1(n5082), .A2(n4629), .A3(n17668), .ZN(n19232) );
  NAND2_X1 U9826 ( .A1(n28188), .A2(n20152), .ZN(n20043) );
  NAND2_X1 U9827 ( .A1(n3166), .A2(n6027), .ZN(n4733) );
  NAND2_X1 U9830 ( .A1(n3171), .A2(n3170), .ZN(n3169) );
  NAND2_X1 U9831 ( .A1(n17124), .A2(n16723), .ZN(n3170) );
  INV_X1 U9832 ( .A(n16725), .ZN(n3172) );
  NAND2_X1 U9834 ( .A1(n6407), .A2(n23331), .ZN(n24397) );
  OAI21_X1 U9836 ( .B1(n11742), .B2(n11740), .A(n3176), .ZN(n11448) );
  NAND2_X1 U9837 ( .A1(n11742), .A2(n11907), .ZN(n3176) );
  NAND3_X1 U9838 ( .A1(n27066), .A2(n26616), .A3(n3178), .ZN(n3177) );
  XNOR2_X1 U9839 ( .A(n16204), .B(n16242), .ZN(n16206) );
  INV_X1 U9841 ( .A(n14178), .ZN(n14450) );
  NAND3_X1 U9843 ( .A1(n8439), .A2(n8785), .A3(n8719), .ZN(n8367) );
  NAND2_X1 U9844 ( .A1(n3806), .A2(n4290), .ZN(n14463) );
  NAND2_X1 U9845 ( .A1(n19927), .A2(n20266), .ZN(n19931) );
  OAI21_X1 U9846 ( .B1(n10876), .B2(n11220), .A(n11104), .ZN(n10535) );
  INV_X1 U9847 ( .A(n6779), .ZN(n5573) );
  NAND2_X1 U9849 ( .A1(n18590), .A2(n18591), .ZN(n18593) );
  NAND2_X1 U9850 ( .A1(n17065), .A2(n17450), .ZN(n17128) );
  AND3_X2 U9852 ( .A1(n24165), .A2(n6946), .A3(n24164), .ZN(n26039) );
  NAND2_X1 U9853 ( .A1(n587), .A2(n11204), .ZN(n11205) );
  NAND2_X1 U9854 ( .A1(n7612), .A2(n7611), .ZN(n3179) );
  NAND3_X1 U9855 ( .A1(n17542), .A2(n17217), .A3(n28454), .ZN(n6642) );
  OAI21_X1 U9856 ( .B1(n11653), .B2(n3603), .A(n12155), .ZN(n3795) );
  XNOR2_X2 U9859 ( .A(n16364), .B(n16363), .ZN(n17374) );
  NAND3_X1 U9860 ( .A1(n3184), .A2(n1840), .A3(n22401), .ZN(n21069) );
  NAND2_X1 U9861 ( .A1(n21068), .A2(n21664), .ZN(n3184) );
  NAND3_X1 U9862 ( .A1(n7883), .A2(n7585), .A3(n7882), .ZN(n3185) );
  NAND2_X1 U9863 ( .A1(n20334), .A2(n20625), .ZN(n3186) );
  NAND3_X1 U9864 ( .A1(n14370), .A2(n14120), .A3(n14366), .ZN(n12977) );
  NAND2_X1 U9866 ( .A1(n23679), .A2(n29544), .ZN(n3189) );
  NOR2_X1 U9867 ( .A1(n28535), .A2(n3190), .ZN(n26133) );
  NAND2_X1 U9868 ( .A1(n7521), .A2(n7266), .ZN(n7710) );
  NAND2_X1 U9869 ( .A1(n5611), .A2(n23761), .ZN(n3192) );
  NAND3_X1 U9870 ( .A1(n20550), .A2(n5982), .A3(n20551), .ZN(n3194) );
  NAND2_X1 U9871 ( .A1(n21321), .A2(n28584), .ZN(n4342) );
  NAND2_X1 U9872 ( .A1(n3797), .A2(n24403), .ZN(n4081) );
  OAI21_X1 U9873 ( .B1(n471), .B2(n24256), .A(n24012), .ZN(n6788) );
  NAND2_X1 U9875 ( .A1(n3716), .A2(n4053), .ZN(n21227) );
  NAND2_X1 U9876 ( .A1(n4540), .A2(n4541), .ZN(n9684) );
  INV_X1 U9877 ( .A(n24639), .ZN(n24196) );
  NOR2_X1 U9879 ( .A1(n20611), .A2(n3547), .ZN(n20442) );
  XNOR2_X1 U9880 ( .A(n16196), .B(n6159), .ZN(n6158) );
  NAND3_X1 U9881 ( .A1(n14446), .A2(n14421), .A3(n13954), .ZN(n13956) );
  NAND2_X1 U9882 ( .A1(n20119), .A2(n19947), .ZN(n20307) );
  NAND2_X1 U9885 ( .A1(n28721), .A2(n7821), .ZN(n6987) );
  NAND2_X1 U9886 ( .A1(n17880), .A2(n19828), .ZN(n17958) );
  NAND2_X1 U9887 ( .A1(n7669), .A2(n7670), .ZN(n7672) );
  OR2_X1 U9889 ( .A1(n12057), .A2(n12313), .ZN(n11772) );
  INV_X1 U9890 ( .A(n15583), .ZN(n16328) );
  NOR2_X1 U9891 ( .A1(n9018), .A2(n9016), .ZN(n8481) );
  OR2_X1 U9892 ( .A1(n14534), .A2(n15456), .ZN(n15177) );
  INV_X1 U9893 ( .A(n5150), .ZN(n10804) );
  AOI22_X1 U9894 ( .A1(n20691), .A2(n20690), .B1(n21366), .B2(n21713), .ZN(
        n21718) );
  INV_X1 U9895 ( .A(n26222), .ZN(n5035) );
  XNOR2_X1 U9896 ( .A(n6212), .B(n21728), .ZN(n22777) );
  NAND2_X1 U9897 ( .A1(n3466), .A2(n3468), .ZN(n3197) );
  NAND2_X1 U9898 ( .A1(n3198), .A2(n10993), .ZN(n3455) );
  NAND2_X1 U9899 ( .A1(n10991), .A2(n10992), .ZN(n3198) );
  NAND3_X1 U9900 ( .A1(n23391), .A2(n23392), .A3(n23839), .ZN(n3199) );
  NAND2_X1 U9901 ( .A1(n11926), .A2(n3201), .ZN(n3200) );
  NAND2_X1 U9902 ( .A1(n11925), .A2(n574), .ZN(n3202) );
  NAND2_X1 U9903 ( .A1(n3203), .A2(n8303), .ZN(n8306) );
  NAND2_X1 U9904 ( .A1(n23304), .A2(n4178), .ZN(n3204) );
  NOR2_X1 U9905 ( .A1(n11347), .A2(n10476), .ZN(n10849) );
  NAND2_X1 U9906 ( .A1(n15409), .A2(n14893), .ZN(n14940) );
  NAND2_X1 U9908 ( .A1(n14994), .A2(n14992), .ZN(n14993) );
  NAND2_X1 U9910 ( .A1(n14916), .A2(n15490), .ZN(n5645) );
  XNOR2_X1 U9911 ( .A(n25889), .B(n25927), .ZN(n24932) );
  AOI21_X1 U9913 ( .B1(n19870), .B2(n3213), .A(n20106), .ZN(n20736) );
  NAND2_X1 U9914 ( .A1(n20147), .A2(n20148), .ZN(n3213) );
  NAND2_X1 U9915 ( .A1(n3216), .A2(n3214), .ZN(n23671) );
  NAND2_X1 U9916 ( .A1(n23669), .A2(n29123), .ZN(n3214) );
  NAND2_X1 U9918 ( .A1(n23664), .A2(n23663), .ZN(n3216) );
  OAI21_X1 U9919 ( .B1(n13206), .B2(n12125), .A(n3217), .ZN(n10441) );
  NAND2_X1 U9920 ( .A1(n11730), .A2(n11824), .ZN(n3217) );
  XNOR2_X1 U9921 ( .A(n13246), .B(n13243), .ZN(n5166) );
  NAND2_X1 U9922 ( .A1(n3314), .A2(n3316), .ZN(n3218) );
  AND3_X1 U9923 ( .A1(n26317), .A2(n26313), .A3(n2441), .ZN(n26319) );
  OAI22_X1 U9925 ( .A1(n26309), .A2(n27155), .B1(n401), .B2(n3220), .ZN(n26312) );
  OR2_X1 U9926 ( .A1(n17303), .A2(n3221), .ZN(n17422) );
  NOR2_X1 U9927 ( .A1(n17421), .A2(n29152), .ZN(n3221) );
  NAND2_X1 U9928 ( .A1(n5714), .A2(n17304), .ZN(n17303) );
  INV_X1 U9929 ( .A(n17018), .ZN(n6539) );
  NAND2_X1 U9930 ( .A1(n15087), .A2(n14563), .ZN(n14878) );
  NAND2_X1 U9931 ( .A1(n7917), .A2(n7912), .ZN(n7630) );
  NAND2_X1 U9932 ( .A1(n5236), .A2(n23153), .ZN(n24642) );
  NAND2_X1 U9933 ( .A1(n8133), .A2(n8048), .ZN(n7556) );
  MUX2_X1 U9934 ( .A(n9064), .B(n8866), .S(n8872), .Z(n8601) );
  XNOR2_X1 U9936 ( .A(n4504), .B(n16589), .ZN(n15998) );
  OAI21_X1 U9937 ( .B1(n11121), .B2(n11123), .A(n6144), .ZN(n10540) );
  NOR2_X1 U9938 ( .A1(n7649), .A2(n7998), .ZN(n7059) );
  NAND3_X1 U9939 ( .A1(n7968), .A2(n7964), .A3(n3226), .ZN(n5470) );
  OR2_X1 U9940 ( .A1(n21109), .A2(n5939), .ZN(n5634) );
  NAND2_X1 U9941 ( .A1(n3595), .A2(n9565), .ZN(n8947) );
  AND2_X1 U9942 ( .A1(n23783), .A2(n23786), .ZN(n23484) );
  NAND2_X1 U9945 ( .A1(n26622), .A2(n27084), .ZN(n3230) );
  INV_X1 U9946 ( .A(n26621), .ZN(n3231) );
  NAND2_X1 U9948 ( .A1(n27327), .A2(n29504), .ZN(n26544) );
  NAND2_X1 U9949 ( .A1(n3235), .A2(n3233), .ZN(n17299) );
  NAND2_X1 U9950 ( .A1(n3234), .A2(n17298), .ZN(n3233) );
  INV_X1 U9951 ( .A(n17296), .ZN(n3234) );
  NAND2_X1 U9952 ( .A1(n17297), .A2(n29072), .ZN(n3235) );
  OAI21_X1 U9955 ( .B1(n25968), .B2(n27003), .A(n29524), .ZN(n25679) );
  OAI21_X1 U9956 ( .B1(n5929), .B2(n21084), .A(n3238), .ZN(n3237) );
  INV_X1 U9957 ( .A(n14192), .ZN(n3269) );
  OAI22_X1 U9958 ( .A1(n27825), .A2(n27828), .B1(n26901), .B2(n27100), .ZN(
        n27249) );
  AOI21_X1 U9959 ( .B1(n6220), .B2(n28428), .A(n28622), .ZN(n23224) );
  INV_X1 U9960 ( .A(n23612), .ZN(n4599) );
  OAI211_X1 U9962 ( .C1(n5129), .C2(n5594), .A(n9425), .B(n3609), .ZN(n5330)
         );
  OR2_X1 U9963 ( .A1(n11113), .A2(n10461), .ZN(n11116) );
  NAND2_X1 U9964 ( .A1(n3241), .A2(n3240), .ZN(n22960) );
  NAND2_X1 U9965 ( .A1(n23391), .A2(n22958), .ZN(n3240) );
  NAND2_X1 U9966 ( .A1(n22959), .A2(n6279), .ZN(n3241) );
  INV_X1 U9967 ( .A(n10856), .ZN(n4591) );
  INV_X1 U9968 ( .A(n19718), .ZN(n5161) );
  OR2_X1 U9969 ( .A1(n17454), .A2(n17455), .ZN(n6800) );
  OR2_X1 U9970 ( .A1(n23343), .A2(n23138), .ZN(n6294) );
  INV_X1 U9972 ( .A(n18538), .ZN(n18528) );
  INV_X1 U9973 ( .A(n26708), .ZN(n25417) );
  INV_X1 U9974 ( .A(n12337), .ZN(n11915) );
  INV_X1 U9976 ( .A(n19463), .ZN(n18675) );
  OAI211_X1 U9977 ( .C1(n25404), .C2(n28908), .A(n25618), .B(n280), .ZN(n5831)
         );
  OAI22_X1 U9978 ( .A1(n18509), .A2(n18078), .B1(n18510), .B2(n418), .ZN(
        n17861) );
  XNOR2_X1 U9979 ( .A(n22269), .B(n22268), .ZN(n22284) );
  XNOR2_X1 U9980 ( .A(n12794), .B(n12793), .ZN(n13674) );
  OAI211_X1 U9981 ( .C1(n10851), .C2(n11163), .A(n11308), .B(n9686), .ZN(n3935) );
  NAND2_X1 U9985 ( .A1(n23613), .A2(n28544), .ZN(n3245) );
  NAND2_X1 U9986 ( .A1(n20444), .A2(n6843), .ZN(n3246) );
  OAI211_X1 U9987 ( .C1(n17620), .C2(n18155), .A(n18156), .B(n3249), .ZN(n3248) );
  NAND2_X1 U9988 ( .A1(n17620), .A2(n18034), .ZN(n3249) );
  NOR2_X1 U9989 ( .A1(n24143), .A2(n24593), .ZN(n3251) );
  INV_X1 U9990 ( .A(n24507), .ZN(n3715) );
  NAND2_X1 U9991 ( .A1(n3254), .A2(n25556), .ZN(n28027) );
  NAND2_X1 U9992 ( .A1(n25555), .A2(n27043), .ZN(n3254) );
  NAND2_X1 U9993 ( .A1(n3259), .A2(n3258), .ZN(n21246) );
  NAND3_X1 U9994 ( .A1(n21242), .A2(n21346), .A3(n21692), .ZN(n3258) );
  NAND2_X1 U9995 ( .A1(n21245), .A2(n3260), .ZN(n3259) );
  OAI211_X1 U9996 ( .C1(n28072), .C2(n28071), .A(n3262), .B(n3261), .ZN(n28074) );
  OR2_X1 U9997 ( .A1(n28070), .A2(n28069), .ZN(n3261) );
  NAND2_X1 U9998 ( .A1(n15100), .A2(n3315), .ZN(n3314) );
  XNOR2_X1 U9999 ( .A(n3263), .B(n26821), .ZN(Ciphertext[33]) );
  INV_X1 U10000 ( .A(n526), .ZN(n3264) );
  NAND2_X1 U10001 ( .A1(n27526), .A2(n27520), .ZN(n27509) );
  NOR2_X2 U10002 ( .A1(n19887), .A2(n19888), .ZN(n21457) );
  NAND2_X1 U10003 ( .A1(n23488), .A2(n23487), .ZN(n3266) );
  NOR2_X1 U10005 ( .A1(n495), .A2(n22013), .ZN(n4380) );
  NAND2_X1 U10006 ( .A1(n17854), .A2(n28142), .ZN(n6716) );
  NAND2_X1 U10010 ( .A1(n21645), .A2(n21642), .ZN(n21399) );
  NAND3_X1 U10011 ( .A1(n8409), .A2(n8408), .A3(n9177), .ZN(n8410) );
  OAI21_X1 U10013 ( .B1(n21304), .B2(n21150), .A(n6602), .ZN(n6601) );
  INV_X1 U10014 ( .A(n26990), .ZN(n26323) );
  NAND2_X1 U10015 ( .A1(n26322), .A2(n5306), .ZN(n26990) );
  NAND2_X1 U10016 ( .A1(n3269), .A2(n14193), .ZN(n13868) );
  NAND3_X1 U10017 ( .A1(n3287), .A2(n4677), .A3(n4853), .ZN(n4852) );
  INV_X1 U10019 ( .A(n17822), .ZN(n3875) );
  NAND2_X1 U10021 ( .A1(n20983), .A2(n20982), .ZN(n21812) );
  NOR2_X1 U10022 ( .A1(n8014), .A2(n7742), .ZN(n8019) );
  INV_X1 U10023 ( .A(n12080), .ZN(n12288) );
  NAND2_X1 U10025 ( .A1(n4278), .A2(n2023), .ZN(n20289) );
  OAI21_X1 U10026 ( .B1(n23356), .B2(n22925), .A(n23461), .ZN(n5269) );
  INV_X1 U10027 ( .A(n4581), .ZN(n20283) );
  OAI21_X1 U10028 ( .B1(n29183), .B2(n6203), .A(n20266), .ZN(n21061) );
  NAND2_X1 U10029 ( .A1(n20451), .A2(n20647), .ZN(n20266) );
  NAND2_X1 U10031 ( .A1(n12164), .A2(n11656), .ZN(n4346) );
  OR2_X1 U10035 ( .A1(n9220), .A2(n8525), .ZN(n8526) );
  INV_X1 U10036 ( .A(n5817), .ZN(n20955) );
  OR2_X1 U10037 ( .A1(n28096), .A2(n28107), .ZN(n3469) );
  OAI21_X1 U10038 ( .B1(n3270), .B2(n27984), .A(n27983), .ZN(n27989) );
  NAND2_X1 U10039 ( .A1(n27981), .A2(n3271), .ZN(n3270) );
  INV_X1 U10040 ( .A(n1793), .ZN(n3274) );
  NAND2_X1 U10041 ( .A1(n586), .A2(n3275), .ZN(n5716) );
  AOI22_X2 U10042 ( .A1(n18190), .A2(n16841), .B1(n16843), .B2(n16842), .ZN(
        n19474) );
  INV_X1 U10043 ( .A(n26448), .ZN(n26452) );
  XNOR2_X1 U10044 ( .A(n16646), .B(n16645), .ZN(n4687) );
  INV_X1 U10045 ( .A(n13914), .ZN(n3798) );
  XNOR2_X1 U10046 ( .A(n10017), .B(n6257), .ZN(n11142) );
  INV_X1 U10047 ( .A(n15202), .ZN(n15201) );
  NOR2_X1 U10048 ( .A1(n27700), .A2(n28504), .ZN(n26351) );
  XNOR2_X2 U10049 ( .A(n24931), .B(n24930), .ZN(n27702) );
  NAND3_X1 U10050 ( .A1(n5494), .A2(n7890), .A3(n7774), .ZN(n5493) );
  NAND2_X1 U10051 ( .A1(n17259), .A2(n29574), .ZN(n4085) );
  NAND2_X1 U10052 ( .A1(n5133), .A2(n29209), .ZN(n12024) );
  NAND2_X1 U10053 ( .A1(n7645), .A2(n7644), .ZN(n3279) );
  NOR2_X1 U10054 ( .A1(n20587), .A2(n20585), .ZN(n3974) );
  NOR2_X1 U10055 ( .A1(n4973), .A2(n4610), .ZN(n4609) );
  NAND2_X1 U10056 ( .A1(n17797), .A2(n17639), .ZN(n16841) );
  AOI21_X1 U10057 ( .B1(n8846), .B2(n11174), .A(n6289), .ZN(n8847) );
  NAND3_X1 U10058 ( .A1(n23884), .A2(n23887), .A3(n23885), .ZN(n23889) );
  NAND4_X2 U10060 ( .A1(n4911), .A2(n4909), .A3(n4910), .A4(n4912), .ZN(n5953)
         );
  OR2_X2 U10064 ( .A1(n7134), .A2(n7135), .ZN(n8109) );
  NAND2_X1 U10065 ( .A1(n17403), .A2(n17404), .ZN(n17408) );
  XNOR2_X1 U10066 ( .A(n19606), .B(n3284), .ZN(n18955) );
  NAND4_X2 U10067 ( .A1(n8068), .A2(n8067), .A3(n8066), .A4(n8065), .ZN(n10144) );
  NAND2_X1 U10069 ( .A1(n3285), .A2(n18234), .ZN(n4371) );
  OR2_X1 U10071 ( .A1(n11260), .A2(n11045), .ZN(n3572) );
  INV_X1 U10072 ( .A(n5918), .ZN(n13720) );
  XNOR2_X2 U10073 ( .A(Key[110]), .B(Plaintext[110]), .ZN(n8216) );
  AOI22_X1 U10074 ( .A1(n3286), .A2(n555), .B1(n6466), .B2(n13687), .ZN(n14630) );
  NAND2_X1 U10075 ( .A1(n13685), .A2(n13893), .ZN(n3286) );
  OR2_X1 U10076 ( .A1(n11423), .A2(n11782), .ZN(n11424) );
  AND2_X1 U10078 ( .A1(n21291), .A2(n21288), .ZN(n20915) );
  NAND2_X1 U10080 ( .A1(n3290), .A2(n3289), .ZN(n17257) );
  NAND2_X1 U10081 ( .A1(n17253), .A2(n16977), .ZN(n3289) );
  NAND2_X1 U10082 ( .A1(n17252), .A2(n16774), .ZN(n3290) );
  AND2_X1 U10083 ( .A1(n1888), .A2(n18251), .ZN(n17774) );
  NAND2_X1 U10084 ( .A1(n24975), .A2(n24258), .ZN(n3291) );
  NAND2_X1 U10085 ( .A1(n23598), .A2(n23597), .ZN(n3292) );
  NAND2_X1 U10086 ( .A1(n3294), .A2(n3293), .ZN(n22176) );
  NAND2_X1 U10087 ( .A1(n380), .A2(n23716), .ZN(n3293) );
  NAND2_X1 U10088 ( .A1(n22163), .A2(n23262), .ZN(n3294) );
  INV_X1 U10089 ( .A(n18388), .ZN(n5233) );
  NOR2_X2 U10091 ( .A1(n12336), .A2(n12335), .ZN(n12644) );
  OR2_X1 U10093 ( .A1(n11113), .A2(n10490), .ZN(n6241) );
  NAND2_X1 U10094 ( .A1(n8268), .A2(n3298), .ZN(n7213) );
  NAND2_X1 U10095 ( .A1(n3299), .A2(n5888), .ZN(n7226) );
  NAND2_X1 U10096 ( .A1(n8686), .A2(n3300), .ZN(n3299) );
  NAND3_X1 U10097 ( .A1(n3302), .A2(n17458), .A3(n16810), .ZN(n17461) );
  OAI21_X1 U10098 ( .B1(n16805), .B2(n16806), .A(n3303), .ZN(n4914) );
  NAND2_X1 U10099 ( .A1(n17261), .A2(n17260), .ZN(n3303) );
  NAND3_X1 U10100 ( .A1(n11111), .A2(n10492), .A3(n10461), .ZN(n10462) );
  NAND2_X1 U10101 ( .A1(n18253), .A2(n18017), .ZN(n18252) );
  MUX2_X1 U10102 ( .A(n22143), .B(n22142), .S(n22139), .Z(n3892) );
  INV_X1 U10103 ( .A(n3893), .ZN(n3304) );
  NAND2_X1 U10104 ( .A1(n3894), .A2(n20580), .ZN(n3305) );
  NAND3_X1 U10105 ( .A1(n4623), .A2(n17550), .A3(n17551), .ZN(n17564) );
  AND2_X1 U10106 ( .A1(n11852), .A2(n11853), .ZN(n3306) );
  AOI21_X1 U10107 ( .B1(n10905), .B2(n11851), .A(n11852), .ZN(n3307) );
  OAI21_X1 U10108 ( .B1(n12232), .B2(n1986), .A(n5579), .ZN(n12040) );
  OAI22_X1 U10109 ( .A1(n5209), .A2(n18170), .B1(n18175), .B2(n28649), .ZN(
        n18176) );
  NAND2_X1 U10111 ( .A1(n7334), .A2(n7333), .ZN(n3308) );
  NAND2_X1 U10112 ( .A1(n27387), .A2(n27400), .ZN(n27241) );
  AND2_X1 U10113 ( .A1(n24256), .A2(n24509), .ZN(n5548) );
  INV_X1 U10114 ( .A(n13979), .ZN(n15113) );
  XNOR2_X1 U10115 ( .A(n1985), .B(n10266), .ZN(n6665) );
  NAND2_X1 U10116 ( .A1(n5454), .A2(n3309), .ZN(n24149) );
  NAND2_X1 U10117 ( .A1(n3310), .A2(n22356), .ZN(n3309) );
  OAI21_X2 U10118 ( .B1(n412), .B2(n21006), .A(n21005), .ZN(n22734) );
  XNOR2_X1 U10119 ( .A(n22299), .B(n22296), .ZN(n6836) );
  NAND2_X1 U10122 ( .A1(n7631), .A2(n29568), .ZN(n7473) );
  OAI211_X2 U10123 ( .C1(n19784), .C2(n21117), .A(n3312), .B(n3311), .ZN(
        n22784) );
  NAND2_X1 U10124 ( .A1(n19783), .A2(n21117), .ZN(n3311) );
  NAND2_X1 U10125 ( .A1(n19782), .A2(n21144), .ZN(n3312) );
  NAND3_X1 U10127 ( .A1(n21394), .A2(n21631), .A3(n21639), .ZN(n3313) );
  NAND2_X1 U10128 ( .A1(n3810), .A2(n7792), .ZN(n7281) );
  XOR2_X1 U10129 ( .A(n19132), .B(n19131), .Z(n6157) );
  NAND3_X1 U10130 ( .A1(n3320), .A2(n21716), .A3(n3319), .ZN(n3318) );
  INV_X1 U10131 ( .A(n21263), .ZN(n3320) );
  NAND2_X1 U10133 ( .A1(n12363), .A2(n12359), .ZN(n10611) );
  NAND2_X1 U10134 ( .A1(n14204), .A2(n427), .ZN(n13684) );
  NAND2_X1 U10136 ( .A1(n12144), .A2(n11712), .ZN(n11710) );
  NAND2_X1 U10137 ( .A1(n11715), .A2(n12146), .ZN(n12144) );
  NAND2_X1 U10138 ( .A1(n409), .A2(n23251), .ZN(n5322) );
  NAND2_X1 U10140 ( .A1(n11262), .A2(n11266), .ZN(n3325) );
  OAI21_X1 U10142 ( .B1(n10993), .B2(n10785), .A(n3328), .ZN(n10996) );
  NAND2_X1 U10143 ( .A1(n10993), .A2(n10992), .ZN(n3328) );
  NAND2_X1 U10144 ( .A1(n7630), .A2(n7633), .ZN(n3330) );
  NAND2_X1 U10145 ( .A1(n7632), .A2(n7914), .ZN(n3331) );
  NAND2_X1 U10146 ( .A1(n28660), .A2(n28545), .ZN(n3332) );
  MUX2_X1 U10148 ( .A(n20743), .B(n3335), .S(n20857), .Z(n20748) );
  NOR2_X1 U10149 ( .A1(n21155), .A2(n20744), .ZN(n3335) );
  XNOR2_X1 U10150 ( .A(n3338), .B(n22408), .ZN(n23049) );
  NAND2_X1 U10151 ( .A1(n3339), .A2(n20121), .ZN(n18118) );
  NAND2_X1 U10152 ( .A1(n20202), .A2(n20201), .ZN(n3339) );
  OAI21_X1 U10154 ( .B1(n8245), .B2(n7818), .A(n3340), .ZN(n7819) );
  NAND2_X1 U10155 ( .A1(n8245), .A2(n7817), .ZN(n3340) );
  MUX2_X1 U10156 ( .A(n29565), .B(n14166), .S(n29306), .Z(n6143) );
  INV_X1 U10158 ( .A(n12868), .ZN(n12396) );
  NOR2_X1 U10160 ( .A1(n23790), .A2(n23789), .ZN(n5770) );
  INV_X1 U10161 ( .A(n5887), .ZN(n5847) );
  AND2_X1 U10162 ( .A1(n17030), .A2(n17357), .ZN(n17031) );
  NAND2_X1 U10163 ( .A1(n14693), .A2(n16995), .ZN(n3342) );
  INV_X1 U10165 ( .A(n11288), .ZN(n10665) );
  XNOR2_X1 U10166 ( .A(n13054), .B(n13159), .ZN(n13353) );
  NAND2_X1 U10167 ( .A1(n3345), .A2(n14689), .ZN(n3344) );
  NAND2_X1 U10168 ( .A1(n13985), .A2(n551), .ZN(n3345) );
  NAND2_X1 U10169 ( .A1(n18588), .A2(n18589), .ZN(n18590) );
  NAND2_X1 U10170 ( .A1(n1835), .A2(n19955), .ZN(n20112) );
  OAI211_X1 U10171 ( .C1(n17948), .C2(n18342), .A(n18344), .B(n3347), .ZN(
        n5771) );
  NAND2_X1 U10172 ( .A1(n17663), .A2(n18342), .ZN(n3347) );
  OAI211_X2 U10173 ( .C1(n29227), .C2(n21281), .A(n20994), .B(n20993), .ZN(
        n22856) );
  OAI211_X1 U10174 ( .C1(n19032), .C2(n20476), .A(n20478), .B(n4556), .ZN(
        n6451) );
  AOI21_X1 U10175 ( .B1(n23682), .B2(n23679), .A(n5882), .ZN(n5881) );
  NAND2_X1 U10176 ( .A1(n20517), .A2(n21356), .ZN(n20262) );
  NAND2_X1 U10177 ( .A1(n14132), .A2(n14342), .ZN(n3348) );
  XNOR2_X1 U10179 ( .A(n19422), .B(n19420), .ZN(n5809) );
  XNOR2_X1 U10180 ( .A(n16229), .B(n4029), .ZN(n16231) );
  NAND2_X1 U10181 ( .A1(n5535), .A2(n28649), .ZN(n3350) );
  NAND2_X1 U10182 ( .A1(n27980), .A2(n28456), .ZN(n27981) );
  AND2_X2 U10183 ( .A1(n3352), .A2(n3351), .ZN(n27908) );
  NAND2_X1 U10184 ( .A1(n27054), .A2(n27053), .ZN(n3352) );
  OAI21_X1 U10186 ( .B1(n9031), .B2(n8433), .A(n3353), .ZN(n8435) );
  INV_X1 U10188 ( .A(n16960), .ZN(n5327) );
  NOR2_X1 U10189 ( .A1(n14763), .A2(n15054), .ZN(n6393) );
  OAI21_X1 U10191 ( .B1(n8651), .B2(n8635), .A(n3354), .ZN(n8660) );
  NAND2_X1 U10192 ( .A1(n8651), .A2(n8652), .ZN(n3354) );
  AND2_X1 U10194 ( .A1(n24772), .A2(n24697), .ZN(n24699) );
  NAND2_X1 U10196 ( .A1(n13620), .A2(n14082), .ZN(n3356) );
  NAND2_X1 U10197 ( .A1(n13621), .A2(n28625), .ZN(n3357) );
  NAND2_X1 U10202 ( .A1(n3362), .A2(n15407), .ZN(n3361) );
  XNOR2_X1 U10203 ( .A(n18998), .B(n19236), .ZN(n19001) );
  XNOR2_X1 U10204 ( .A(n19468), .B(n19555), .ZN(n19236) );
  OAI22_X1 U10205 ( .A1(n17757), .A2(n522), .B1(n17966), .B2(n18240), .ZN(
        n17537) );
  NAND2_X1 U10206 ( .A1(n11969), .A2(n12158), .ZN(n10861) );
  INV_X1 U10209 ( .A(n27632), .ZN(n3366) );
  NAND2_X1 U10210 ( .A1(n1912), .A2(n27625), .ZN(n3367) );
  OAI21_X1 U10211 ( .B1(n11322), .B2(n11321), .A(n29316), .ZN(n6722) );
  INV_X1 U10215 ( .A(n7705), .ZN(n3639) );
  NAND2_X1 U10216 ( .A1(n7959), .A2(n7958), .ZN(n3368) );
  NAND3_X1 U10217 ( .A1(n3370), .A2(n6273), .A3(n6274), .ZN(n22919) );
  OAI211_X1 U10218 ( .C1(n21012), .C2(n21442), .A(n3371), .B(n21656), .ZN(
        n3370) );
  NAND2_X1 U10219 ( .A1(n21660), .A2(n20833), .ZN(n3371) );
  INV_X1 U10220 ( .A(n14393), .ZN(n13951) );
  OAI211_X1 U10221 ( .C1(n28157), .C2(n581), .A(n10751), .B(n11197), .ZN(n3373) );
  NAND2_X1 U10222 ( .A1(n20587), .A2(n20585), .ZN(n17880) );
  AND2_X1 U10223 ( .A1(n14358), .A2(n4166), .ZN(n3375) );
  NAND2_X1 U10224 ( .A1(n6314), .A2(n29101), .ZN(n21697) );
  INV_X1 U10226 ( .A(n4364), .ZN(n24630) );
  INV_X1 U10227 ( .A(n17834), .ZN(n18588) );
  INV_X1 U10228 ( .A(n23535), .ZN(n23694) );
  MUX2_X1 U10229 ( .A(n26265), .B(n26264), .S(n28392), .Z(n3376) );
  OAI21_X1 U10230 ( .B1(n8765), .B2(n9561), .A(n3377), .ZN(n8332) );
  NAND2_X1 U10231 ( .A1(n8765), .A2(n8944), .ZN(n3377) );
  NAND2_X1 U10232 ( .A1(n4885), .A2(n4886), .ZN(n4888) );
  XNOR2_X1 U10233 ( .A(n12955), .B(n3382), .ZN(n6831) );
  OAI21_X2 U10234 ( .B1(n17292), .B2(n17291), .A(n17295), .ZN(n18033) );
  OAI21_X1 U10236 ( .B1(n11767), .B2(n4197), .A(n3383), .ZN(n5019) );
  NAND2_X1 U10237 ( .A1(n3384), .A2(n4197), .ZN(n3383) );
  INV_X1 U10238 ( .A(n12305), .ZN(n3384) );
  NAND2_X1 U10239 ( .A1(n7589), .A2(n7233), .ZN(n7869) );
  NAND2_X1 U10240 ( .A1(n12976), .A2(n14091), .ZN(n14092) );
  AND2_X1 U10241 ( .A1(n20178), .A2(n20173), .ZN(n19055) );
  NAND2_X1 U10242 ( .A1(n18344), .A2(n18341), .ZN(n18340) );
  NAND2_X1 U10243 ( .A1(n3387), .A2(n20091), .ZN(n20094) );
  NOR2_X1 U10244 ( .A1(n20041), .A2(n20093), .ZN(n3387) );
  XNOR2_X1 U10245 ( .A(n21756), .B(n1271), .ZN(n6074) );
  NAND2_X1 U10248 ( .A1(n7978), .A2(n7979), .ZN(n8073) );
  NAND3_X1 U10249 ( .A1(n8730), .A2(n8731), .A3(n8381), .ZN(n7186) );
  NAND2_X1 U10251 ( .A1(n4916), .A2(n23447), .ZN(n3391) );
  NAND2_X1 U10252 ( .A1(n4915), .A2(n23371), .ZN(n3392) );
  NAND2_X1 U10253 ( .A1(n14064), .A2(n13652), .ZN(n3393) );
  NAND2_X1 U10254 ( .A1(n16788), .A2(n6002), .ZN(n5068) );
  NAND2_X1 U10256 ( .A1(n3396), .A2(n14264), .ZN(n3395) );
  INV_X1 U10257 ( .A(n14259), .ZN(n3396) );
  NAND3_X1 U10258 ( .A1(n29132), .A2(n28536), .A3(n27177), .ZN(n3397) );
  OAI21_X2 U10260 ( .B1(n22741), .B2(n23445), .A(n22740), .ZN(n24552) );
  NAND2_X1 U10261 ( .A1(n6541), .A2(n26800), .ZN(n6323) );
  NAND3_X1 U10262 ( .A1(n21158), .A2(n20744), .A3(n3401), .ZN(n3400) );
  INV_X1 U10264 ( .A(n15895), .ZN(n5447) );
  NAND2_X2 U10265 ( .A1(n4239), .A2(n4238), .ZN(n25836) );
  AOI21_X1 U10266 ( .B1(n5028), .B2(n23137), .A(n23694), .ZN(n3405) );
  XNOR2_X1 U10267 ( .A(n3406), .B(n16343), .ZN(n15931) );
  XNOR2_X1 U10268 ( .A(n15926), .B(n15925), .ZN(n3406) );
  NAND2_X1 U10269 ( .A1(n3409), .A2(n3408), .ZN(n13743) );
  NAND2_X1 U10270 ( .A1(n13742), .A2(n29306), .ZN(n3409) );
  OAI21_X1 U10272 ( .B1(n11852), .B2(n574), .A(n3410), .ZN(n10908) );
  INV_X1 U10273 ( .A(n4460), .ZN(n20830) );
  NAND2_X1 U10274 ( .A1(n20068), .A2(n20065), .ZN(n3411) );
  OAI211_X1 U10275 ( .C1(n10780), .C2(n28173), .A(n3413), .B(n10959), .ZN(
        n6773) );
  AOI21_X1 U10276 ( .B1(n24706), .B2(n29043), .A(n6612), .ZN(n6611) );
  XOR2_X1 U10277 ( .A(n10295), .B(n9613), .Z(n5032) );
  XNOR2_X1 U10278 ( .A(n25790), .B(n25543), .ZN(n25260) );
  INV_X1 U10279 ( .A(n4180), .ZN(n4179) );
  OAI21_X1 U10280 ( .B1(n8924), .B2(n9132), .A(n9131), .ZN(n9136) );
  INV_X1 U10281 ( .A(n15535), .ZN(n16653) );
  INV_X1 U10282 ( .A(n17276), .ZN(n16844) );
  OR2_X1 U10284 ( .A1(n9024), .A2(n8687), .ZN(n5889) );
  XNOR2_X1 U10286 ( .A(n25937), .B(n25936), .ZN(n27056) );
  NAND2_X1 U10288 ( .A1(n16819), .A2(n387), .ZN(n3415) );
  NAND2_X1 U10289 ( .A1(n16820), .A2(n17463), .ZN(n3416) );
  NOR2_X1 U10290 ( .A1(n16673), .A2(n17464), .ZN(n16820) );
  AND2_X1 U10292 ( .A1(n18383), .A2(n18379), .ZN(n5670) );
  XNOR2_X1 U10293 ( .A(n12830), .B(n13371), .ZN(n13479) );
  NAND2_X1 U10295 ( .A1(n13411), .A2(n2075), .ZN(n14881) );
  NAND2_X1 U10297 ( .A1(n3417), .A2(n21394), .ZN(n21228) );
  NAND2_X1 U10298 ( .A1(n21226), .A2(n3418), .ZN(n3417) );
  OR2_X1 U10301 ( .A1(n20720), .A2(n21596), .ZN(n20723) );
  OAI21_X1 U10302 ( .B1(n3421), .B2(n19890), .A(n3420), .ZN(n19894) );
  NAND2_X1 U10303 ( .A1(n19890), .A2(n28894), .ZN(n3420) );
  INV_X1 U10304 ( .A(n14039), .ZN(n13997) );
  INV_X1 U10305 ( .A(n14971), .ZN(n5813) );
  NOR2_X1 U10306 ( .A1(n20700), .A2(n21691), .ZN(n6313) );
  NOR2_X1 U10307 ( .A1(n10818), .A2(n10817), .ZN(n11646) );
  INV_X1 U10308 ( .A(n14923), .ZN(n15498) );
  INV_X1 U10309 ( .A(n21227), .ZN(n21633) );
  XNOR2_X1 U10310 ( .A(n12421), .B(n12652), .ZN(n11866) );
  INV_X1 U10312 ( .A(n21632), .ZN(n21637) );
  XNOR2_X1 U10313 ( .A(n22657), .B(n6863), .ZN(n20277) );
  XNOR2_X1 U10314 ( .A(n19408), .B(n16990), .ZN(n19590) );
  NAND2_X1 U10315 ( .A1(n3427), .A2(n3424), .ZN(n27437) );
  NAND3_X1 U10316 ( .A1(n3426), .A2(n3425), .A3(n26710), .ZN(n3424) );
  NAND2_X1 U10317 ( .A1(n27442), .A2(n27433), .ZN(n3425) );
  INV_X1 U10318 ( .A(n27432), .ZN(n3426) );
  NAND2_X1 U10319 ( .A1(n27435), .A2(n27434), .ZN(n3427) );
  NAND2_X1 U10320 ( .A1(n8201), .A2(n3431), .ZN(n3430) );
  NAND3_X1 U10321 ( .A1(n3433), .A2(n3748), .A3(n14917), .ZN(n14503) );
  NAND2_X1 U10322 ( .A1(n14703), .A2(n15489), .ZN(n3433) );
  AOI22_X1 U10323 ( .A1(n17108), .A2(n17472), .B1(n17107), .B2(n17470), .ZN(
        n17112) );
  OAI21_X1 U10324 ( .B1(n23169), .B2(n23516), .A(n3434), .ZN(n23521) );
  NAND2_X1 U10326 ( .A1(n15308), .A2(n15309), .ZN(n15271) );
  NAND3_X1 U10328 ( .A1(n14086), .A2(n14088), .A3(n14087), .ZN(n14089) );
  AND2_X1 U10329 ( .A1(n12271), .A2(n12270), .ZN(n11103) );
  INV_X1 U10330 ( .A(n24460), .ZN(n5004) );
  OAI211_X2 U10332 ( .C1(n6671), .C2(n3849), .A(n6670), .B(n18457), .ZN(n19595) );
  XNOR2_X1 U10333 ( .A(n9351), .B(n10188), .ZN(n3437) );
  NAND2_X1 U10334 ( .A1(n3438), .A2(n11707), .ZN(n12495) );
  NAND2_X1 U10336 ( .A1(n29559), .A2(n17283), .ZN(n16066) );
  NAND2_X1 U10337 ( .A1(n20571), .A2(n20568), .ZN(n3443) );
  AND2_X2 U10338 ( .A1(n6215), .A2(n2065), .ZN(n24852) );
  NAND2_X1 U10339 ( .A1(n8206), .A2(n3446), .ZN(n8836) );
  OAI211_X1 U10340 ( .C1(n8199), .C2(n28605), .A(n3448), .B(n3447), .ZN(n3446)
         );
  NAND2_X1 U10341 ( .A1(n8199), .A2(n8201), .ZN(n3448) );
  NAND3_X1 U10343 ( .A1(n6359), .A2(n6360), .A3(n10742), .ZN(n3449) );
  NAND2_X1 U10344 ( .A1(n28205), .A2(n10461), .ZN(n10099) );
  MUX2_X2 U10345 ( .A(n14152), .B(n14151), .S(n14380), .Z(n15359) );
  NAND3_X1 U10346 ( .A1(n21589), .A2(n20714), .A3(n5683), .ZN(n5206) );
  INV_X1 U10348 ( .A(n11751), .ZN(n4712) );
  NAND2_X1 U10349 ( .A1(n6439), .A2(n23429), .ZN(n23599) );
  INV_X1 U10350 ( .A(n10971), .ZN(n5267) );
  XNOR2_X1 U10351 ( .A(n3452), .B(n9295), .ZN(n10338) );
  XNOR2_X1 U10352 ( .A(n18727), .B(n1981), .ZN(n5586) );
  NAND2_X1 U10353 ( .A1(n10994), .A2(n3454), .ZN(n3453) );
  OAI22_X1 U10354 ( .A1(n10501), .A2(n10497), .B1(n11132), .B2(n10500), .ZN(
        n3458) );
  NAND2_X1 U10355 ( .A1(n21193), .A2(n6936), .ZN(n21197) );
  NAND2_X1 U10356 ( .A1(n11677), .A2(n11676), .ZN(n11678) );
  NAND2_X1 U10357 ( .A1(n21551), .A2(n21519), .ZN(n21552) );
  NAND2_X1 U10358 ( .A1(n15265), .A2(n14923), .ZN(n15266) );
  MUX2_X2 U10361 ( .A(n18250), .B(n18249), .S(n28558), .Z(n19496) );
  NAND2_X1 U10362 ( .A1(n11403), .A2(n11118), .ZN(n3461) );
  NAND3_X2 U10363 ( .A1(n9777), .A2(n9778), .A3(n11234), .ZN(n12189) );
  MUX2_X2 U10364 ( .A(n19775), .B(n19774), .S(n20098), .Z(n21119) );
  NOR2_X2 U10365 ( .A1(n4393), .A2(n21147), .ZN(n22059) );
  INV_X1 U10366 ( .A(n14366), .ZN(n14094) );
  AOI22_X1 U10367 ( .A1(n28179), .A2(n28429), .B1(n27585), .B2(n27596), .ZN(
        n27598) );
  INV_X1 U10368 ( .A(n7641), .ZN(n7457) );
  XNOR2_X1 U10369 ( .A(n16203), .B(n16202), .ZN(n6870) );
  NAND2_X1 U10370 ( .A1(n7886), .A2(n7583), .ZN(n7882) );
  NAND2_X1 U10371 ( .A1(n7580), .A2(n7582), .ZN(n3464) );
  OR2_X1 U10372 ( .A1(n18688), .A2(n18687), .ZN(n18703) );
  NOR2_X1 U10373 ( .A1(n6077), .A2(n18473), .ZN(n6076) );
  NAND3_X1 U10375 ( .A1(n28489), .A2(n20511), .A3(n19785), .ZN(n4912) );
  INV_X1 U10376 ( .A(n26733), .ZN(n5389) );
  NAND2_X1 U10377 ( .A1(n23318), .A2(n23648), .ZN(n23192) );
  NAND2_X1 U10378 ( .A1(n18151), .A2(n3467), .ZN(n3466) );
  INV_X1 U10379 ( .A(n18149), .ZN(n3467) );
  INV_X1 U10380 ( .A(n23290), .ZN(n5591) );
  INV_X1 U10381 ( .A(n24380), .ZN(n23906) );
  NAND2_X1 U10382 ( .A1(n17097), .A2(n17098), .ZN(n17099) );
  NAND2_X1 U10383 ( .A1(n28094), .A2(n28107), .ZN(n3470) );
  NAND2_X1 U10384 ( .A1(n24737), .A2(n24738), .ZN(n24742) );
  NAND3_X1 U10386 ( .A1(n4391), .A2(n18135), .A3(n3471), .ZN(n17636) );
  NAND2_X1 U10387 ( .A1(n21668), .A2(n4312), .ZN(n3474) );
  NAND2_X1 U10388 ( .A1(n21667), .A2(n22404), .ZN(n3475) );
  NAND2_X1 U10389 ( .A1(n3477), .A2(n18430), .ZN(n18436) );
  NAND2_X1 U10390 ( .A1(n18429), .A2(n4762), .ZN(n3477) );
  NAND2_X1 U10391 ( .A1(n2855), .A2(n18433), .ZN(n18429) );
  XNOR2_X1 U10392 ( .A(n3478), .B(n27453), .ZN(Ciphertext[42]) );
  NAND4_X1 U10393 ( .A1(n27450), .A2(n27451), .A3(n27448), .A4(n27449), .ZN(
        n3478) );
  NAND2_X1 U10394 ( .A1(n10742), .A2(n10808), .ZN(n7814) );
  OAI22_X1 U10395 ( .A1(n18887), .A2(n20150), .B1(n20099), .B2(n20098), .ZN(
        n20156) );
  NAND2_X1 U10396 ( .A1(n3479), .A2(n5599), .ZN(n5596) );
  NAND2_X1 U10397 ( .A1(n5597), .A2(n14551), .ZN(n3479) );
  NAND2_X1 U10398 ( .A1(n11283), .A2(n1854), .ZN(n11285) );
  INV_X1 U10399 ( .A(n21425), .ZN(n21085) );
  INV_X1 U10400 ( .A(n21494), .ZN(n20867) );
  OAI22_X1 U10401 ( .A1(n4025), .A2(n3480), .B1(n6406), .B2(n24324), .ZN(
        n24326) );
  NAND2_X1 U10402 ( .A1(n18425), .A2(n18426), .ZN(n18427) );
  NOR2_X1 U10403 ( .A1(n15389), .A2(n6517), .ZN(n14631) );
  NAND2_X1 U10404 ( .A1(n5557), .A2(n17301), .ZN(n15812) );
  NOR2_X2 U10405 ( .A1(n14666), .A2(n14660), .ZN(n15444) );
  NAND2_X1 U10406 ( .A1(n17299), .A2(n17415), .ZN(n3484) );
  NAND2_X1 U10410 ( .A1(n20946), .A2(n20945), .ZN(n5879) );
  INV_X1 U10411 ( .A(n20557), .ZN(n20548) );
  NAND2_X1 U10412 ( .A1(n17172), .A2(n28501), .ZN(n20557) );
  NAND3_X1 U10413 ( .A1(n14069), .A2(n14070), .A3(n6351), .ZN(n3488) );
  NAND2_X1 U10414 ( .A1(n21258), .A2(n21714), .ZN(n20977) );
  NAND2_X1 U10415 ( .A1(n7466), .A2(n28615), .ZN(n3489) );
  NAND2_X1 U10416 ( .A1(n6782), .A2(n6783), .ZN(n3490) );
  NAND2_X1 U10417 ( .A1(n21716), .A2(n21368), .ZN(n3492) );
  NAND3_X1 U10419 ( .A1(n5072), .A2(n7519), .A3(n7518), .ZN(n8592) );
  NAND2_X1 U10420 ( .A1(n3496), .A2(n3495), .ZN(n24001) );
  OR2_X1 U10421 ( .A1(n22951), .A2(n23397), .ZN(n3495) );
  OAI21_X1 U10422 ( .B1(n23401), .B2(n22950), .A(n23227), .ZN(n3496) );
  OAI211_X1 U10423 ( .C1(n29467), .C2(n3498), .A(n26456), .B(n3497), .ZN(n6736) );
  NAND3_X1 U10425 ( .A1(n23512), .A2(n23772), .A3(n23487), .ZN(n3499) );
  NAND2_X1 U10426 ( .A1(n3500), .A2(n12205), .ZN(n11440) );
  NAND2_X1 U10427 ( .A1(n11438), .A2(n11599), .ZN(n3500) );
  OR3_X1 U10429 ( .A1(n15290), .A2(n15217), .A3(n15036), .ZN(n15219) );
  OR2_X1 U10430 ( .A1(n4451), .A2(n14085), .ZN(n14086) );
  OR2_X1 U10431 ( .A1(n25239), .A2(n27395), .ZN(n25241) );
  OR2_X1 U10432 ( .A1(n14688), .A2(n15004), .ZN(n4689) );
  NAND2_X1 U10433 ( .A1(n20635), .A2(n20247), .ZN(n3503) );
  NAND2_X1 U10434 ( .A1(n498), .A2(n20632), .ZN(n3504) );
  INV_X1 U10435 ( .A(n17772), .ZN(n18018) );
  NOR2_X1 U10436 ( .A1(n18120), .A2(n4240), .ZN(n17821) );
  NAND3_X1 U10437 ( .A1(n23263), .A2(n23713), .A3(n3505), .ZN(n23264) );
  OAI21_X1 U10438 ( .B1(n380), .B2(n23710), .A(n23262), .ZN(n3505) );
  NOR2_X1 U10439 ( .A1(n26463), .A2(n2015), .ZN(n26471) );
  NAND2_X1 U10440 ( .A1(n545), .A2(n15464), .ZN(n3506) );
  NAND2_X1 U10441 ( .A1(n15159), .A2(n29153), .ZN(n3507) );
  OAI21_X2 U10442 ( .B1(n19677), .B2(n19808), .A(n19676), .ZN(n19732) );
  NAND2_X1 U10443 ( .A1(n9095), .A2(n8666), .ZN(n8631) );
  AOI21_X1 U10444 ( .B1(n7231), .B2(n441), .A(n7957), .ZN(n7961) );
  AOI21_X1 U10445 ( .B1(n3511), .B2(n3510), .A(n7692), .ZN(n7694) );
  NAND2_X1 U10446 ( .A1(n24064), .A2(n28415), .ZN(n3512) );
  NAND2_X1 U10447 ( .A1(n23269), .A2(n24138), .ZN(n3514) );
  NAND2_X1 U10448 ( .A1(n4611), .A2(n15251), .ZN(n15253) );
  OAI21_X1 U10449 ( .B1(n21192), .B2(n28611), .A(n3515), .ZN(n21544) );
  NAND2_X1 U10450 ( .A1(n28611), .A2(n21539), .ZN(n3515) );
  NOR2_X1 U10451 ( .A1(n28088), .A2(n3517), .ZN(Ciphertext[188]) );
  INV_X1 U10453 ( .A(n18136), .ZN(n5623) );
  NOR2_X1 U10454 ( .A1(n14752), .A2(n14153), .ZN(n15358) );
  AOI21_X1 U10456 ( .B1(n407), .B2(n28609), .A(n23816), .ZN(n3518) );
  OAI21_X1 U10457 ( .B1(n17425), .B2(n2826), .A(n3520), .ZN(n17432) );
  NAND2_X1 U10458 ( .A1(n17425), .A2(n5891), .ZN(n3520) );
  INV_X1 U10459 ( .A(n23773), .ZN(n6424) );
  OAI21_X1 U10460 ( .B1(n11549), .B2(n574), .A(n3521), .ZN(n10094) );
  NAND2_X1 U10461 ( .A1(n17598), .A2(n28558), .ZN(n3523) );
  NAND2_X1 U10462 ( .A1(n17599), .A2(n5021), .ZN(n3524) );
  NAND2_X1 U10463 ( .A1(n17600), .A2(n18709), .ZN(n3525) );
  NAND2_X1 U10464 ( .A1(n1320), .A2(n3526), .ZN(n5642) );
  OR2_X1 U10465 ( .A1(n16878), .A2(n16700), .ZN(n17159) );
  INV_X1 U10466 ( .A(n14174), .ZN(n15195) );
  OAI21_X1 U10467 ( .B1(n20623), .B2(n20626), .A(n20628), .ZN(n5318) );
  INV_X1 U10468 ( .A(n8808), .ZN(n8681) );
  XNOR2_X1 U10469 ( .A(n5984), .B(n10150), .ZN(n10155) );
  XNOR2_X1 U10470 ( .A(n22500), .B(n26032), .ZN(n5718) );
  NAND2_X1 U10471 ( .A1(n5918), .A2(n14039), .ZN(n6032) );
  AOI22_X1 U10473 ( .A1(n17270), .A2(n17265), .B1(n17269), .B2(n17268), .ZN(
        n17534) );
  NAND2_X1 U10475 ( .A1(n10515), .A2(n10516), .ZN(n12529) );
  NAND4_X2 U10476 ( .A1(n11306), .A2(n11305), .A3(n11304), .A4(n11303), .ZN(
        n13075) );
  OR2_X1 U10479 ( .A1(n10585), .A2(n3802), .ZN(n3533) );
  NAND2_X1 U10480 ( .A1(n1941), .A2(n2026), .ZN(n3534) );
  NAND2_X1 U10481 ( .A1(n16701), .A2(n29045), .ZN(n3535) );
  NAND2_X1 U10482 ( .A1(n10823), .A2(n3536), .ZN(n10822) );
  NAND2_X1 U10483 ( .A1(n8688), .A2(n8687), .ZN(n9227) );
  NAND2_X1 U10484 ( .A1(n17730), .A2(n18455), .ZN(n3538) );
  NAND2_X1 U10485 ( .A1(n17731), .A2(n18107), .ZN(n3539) );
  AND2_X1 U10486 ( .A1(n29641), .A2(n23772), .ZN(n21862) );
  NAND2_X1 U10487 ( .A1(n3540), .A2(n17721), .ZN(n17723) );
  NAND2_X1 U10488 ( .A1(n4621), .A2(n14116), .ZN(n4620) );
  OR2_X2 U10491 ( .A1(n7356), .A2(n7355), .ZN(n10193) );
  XOR2_X1 U10492 ( .A(n9388), .B(n9387), .Z(n4716) );
  AND2_X2 U10493 ( .A1(n20776), .A2(n20777), .ZN(n21500) );
  NAND3_X2 U10494 ( .A1(n6660), .A2(n6659), .A3(n11539), .ZN(n12830) );
  XNOR2_X2 U10495 ( .A(n5924), .B(n5925), .ZN(n10808) );
  AOI21_X1 U10496 ( .B1(n3543), .B2(n11740), .A(n12363), .ZN(n10615) );
  NAND2_X1 U10497 ( .A1(n11739), .A2(n12356), .ZN(n3543) );
  NAND2_X1 U10498 ( .A1(n11708), .A2(n11648), .ZN(n11416) );
  NAND2_X1 U10499 ( .A1(n3546), .A2(n3545), .ZN(n14597) );
  NAND2_X1 U10500 ( .A1(n14256), .A2(n14255), .ZN(n3545) );
  NAND2_X1 U10501 ( .A1(n14257), .A2(n14254), .ZN(n3546) );
  NAND2_X1 U10502 ( .A1(n10553), .A2(n10554), .ZN(n10555) );
  NAND2_X1 U10503 ( .A1(n10804), .A2(n10752), .ZN(n10553) );
  NAND3_X1 U10505 ( .A1(n22291), .A2(n29364), .A3(n3548), .ZN(n21055) );
  NAND3_X1 U10507 ( .A1(n29624), .A2(n24769), .A3(n24768), .ZN(n24770) );
  XNOR2_X1 U10508 ( .A(n5452), .B(n5453), .ZN(n23353) );
  OR2_X1 U10509 ( .A1(n20300), .A2(n6843), .ZN(n3551) );
  NOR2_X1 U10510 ( .A1(n8932), .A2(n6072), .ZN(n8933) );
  OAI211_X1 U10511 ( .C1(n20552), .C2(n6086), .A(n20553), .B(n6085), .ZN(n6084) );
  INV_X1 U10512 ( .A(n349), .ZN(n3552) );
  OR2_X1 U10513 ( .A1(n17989), .A2(n28142), .ZN(n17014) );
  AND2_X1 U10514 ( .A1(n7864), .A2(n7092), .ZN(n5191) );
  INV_X1 U10515 ( .A(n4193), .ZN(n21458) );
  NOR2_X1 U10516 ( .A1(n23303), .A2(n5530), .ZN(n23105) );
  INV_X1 U10517 ( .A(n17568), .ZN(n4118) );
  OAI21_X1 U10520 ( .B1(n20844), .B2(n20843), .A(n4193), .ZN(n3555) );
  OR2_X1 U10522 ( .A1(n14517), .A2(n15292), .ZN(n15216) );
  NAND2_X1 U10523 ( .A1(n12062), .A2(n3557), .ZN(n3556) );
  NAND2_X1 U10524 ( .A1(n8553), .A2(n8762), .ZN(n8764) );
  NAND2_X1 U10525 ( .A1(n20955), .A2(n20802), .ZN(n3559) );
  XNOR2_X1 U10528 ( .A(n9927), .B(n9926), .ZN(n10097) );
  NOR2_X2 U10529 ( .A1(n7693), .A2(n7694), .ZN(n9030) );
  NAND2_X1 U10530 ( .A1(n23319), .A2(n23493), .ZN(n23323) );
  NAND2_X1 U10531 ( .A1(n21569), .A2(n21570), .ZN(n3563) );
  NAND2_X1 U10532 ( .A1(n20314), .A2(n20585), .ZN(n19828) );
  NAND2_X1 U10534 ( .A1(n4345), .A2(n12163), .ZN(n3566) );
  NAND2_X1 U10535 ( .A1(n14846), .A2(n14845), .ZN(n14847) );
  AOI21_X1 U10536 ( .B1(n24120), .B2(n24121), .A(n403), .ZN(n3567) );
  AOI22_X1 U10537 ( .A1(n11978), .A2(n11977), .B1(n6871), .B2(n28201), .ZN(
        n4261) );
  NAND2_X1 U10538 ( .A1(n28201), .A2(n12234), .ZN(n11977) );
  OR2_X1 U10539 ( .A1(n20047), .A2(n28187), .ZN(n19987) );
  INV_X1 U10543 ( .A(n15998), .ZN(n16177) );
  NAND2_X1 U10544 ( .A1(n23979), .A2(n28519), .ZN(n23980) );
  XNOR2_X1 U10545 ( .A(n21998), .B(n21728), .ZN(n22246) );
  NAND2_X1 U10547 ( .A1(n18224), .A2(n17532), .ZN(n18387) );
  XNOR2_X1 U10549 ( .A(n10030), .B(n10027), .ZN(n5400) );
  INV_X1 U10550 ( .A(n22256), .ZN(n6378) );
  INV_X1 U10551 ( .A(n21457), .ZN(n21125) );
  NAND2_X1 U10553 ( .A1(n28438), .A2(n27944), .ZN(n3571) );
  AOI21_X2 U10554 ( .B1(n18310), .B2(n18309), .A(n18308), .ZN(n19688) );
  MUX2_X2 U10555 ( .A(n15768), .B(n15767), .S(n17560), .Z(n18063) );
  NOR2_X1 U10556 ( .A1(n3572), .A2(n6515), .ZN(n6514) );
  NAND2_X1 U10557 ( .A1(n3573), .A2(n4995), .ZN(n23992) );
  NAND2_X1 U10558 ( .A1(n4993), .A2(n24634), .ZN(n3573) );
  XNOR2_X1 U10559 ( .A(n11805), .B(n11804), .ZN(n13744) );
  NAND2_X1 U10561 ( .A1(n14792), .A2(n14881), .ZN(n14584) );
  OAI21_X2 U10562 ( .B1(n22961), .B2(n28418), .A(n22960), .ZN(n24020) );
  INV_X1 U10563 ( .A(n3575), .ZN(n3574) );
  OAI21_X1 U10564 ( .B1(n14765), .B2(n15262), .A(n3576), .ZN(n3575) );
  NAND2_X1 U10565 ( .A1(n6393), .A2(n15053), .ZN(n3576) );
  NAND2_X1 U10566 ( .A1(n14764), .A2(n15056), .ZN(n3577) );
  OAI21_X1 U10569 ( .B1(n17067), .B2(n17066), .A(n17065), .ZN(n4831) );
  OR2_X1 U10570 ( .A1(n11188), .A2(n11187), .ZN(n3905) );
  NAND2_X1 U10571 ( .A1(n12714), .A2(n4290), .ZN(n3579) );
  INV_X1 U10572 ( .A(n14460), .ZN(n3580) );
  NAND2_X1 U10573 ( .A1(n12713), .A2(n14460), .ZN(n3581) );
  XNOR2_X1 U10574 ( .A(n15634), .B(n16131), .ZN(n15635) );
  XNOR2_X1 U10575 ( .A(n16166), .B(n16167), .ZN(n3582) );
  OR2_X1 U10576 ( .A1(n15420), .A2(n15101), .ZN(n4547) );
  INV_X1 U10577 ( .A(n14451), .ZN(n14181) );
  INV_X1 U10578 ( .A(n13118), .ZN(n12637) );
  INV_X1 U10579 ( .A(n29145), .ZN(n3735) );
  XNOR2_X1 U10581 ( .A(n13104), .B(n13552), .ZN(n6375) );
  NAND3_X1 U10582 ( .A1(n23286), .A2(n5763), .A3(n23075), .ZN(n23076) );
  AOI22_X1 U10583 ( .A1(n5575), .A2(n6699), .B1(n15499), .B2(n14431), .ZN(
        n3583) );
  NAND2_X1 U10584 ( .A1(n11197), .A2(n10814), .ZN(n3584) );
  NOR2_X1 U10585 ( .A1(n17475), .A2(n3883), .ZN(n4367) );
  NAND2_X1 U10588 ( .A1(n27446), .A2(n27472), .ZN(n26907) );
  NAND2_X1 U10589 ( .A1(n7254), .A2(n3593), .ZN(n7255) );
  NAND2_X1 U10590 ( .A1(n7383), .A2(n3594), .ZN(n3593) );
  XNOR2_X1 U10592 ( .A(n23961), .B(n25713), .ZN(n3596) );
  NAND2_X1 U10594 ( .A1(n11273), .A2(n10522), .ZN(n11039) );
  NAND2_X1 U10595 ( .A1(n4245), .A2(n20265), .ZN(n20644) );
  XNOR2_X2 U10596 ( .A(n19539), .B(n19538), .ZN(n4245) );
  NAND3_X1 U10597 ( .A1(n3600), .A2(n24096), .A3(n3599), .ZN(n24099) );
  NAND2_X1 U10598 ( .A1(n24470), .A2(n24092), .ZN(n3600) );
  OAI211_X1 U10599 ( .C1(n7773), .C2(n7315), .A(n3601), .B(n7775), .ZN(n7277)
         );
  NAND2_X1 U10600 ( .A1(n7773), .A2(n7089), .ZN(n3601) );
  OAI22_X1 U10603 ( .A1(n28126), .A2(n4167), .B1(n28133), .B2(n21359), .ZN(
        n20263) );
  NAND2_X1 U10605 ( .A1(n13885), .A2(n14319), .ZN(n3602) );
  NAND2_X1 U10606 ( .A1(n3964), .A2(n4844), .ZN(n3963) );
  OR2_X1 U10607 ( .A1(n17719), .A2(n17859), .ZN(n17721) );
  NAND2_X1 U10608 ( .A1(n17438), .A2(n17433), .ZN(n17436) );
  NAND2_X1 U10609 ( .A1(n13694), .A2(n14323), .ZN(n13695) );
  XNOR2_X1 U10610 ( .A(n13315), .B(n13220), .ZN(n13094) );
  INV_X1 U10611 ( .A(n23486), .ZN(n3700) );
  NOR2_X2 U10612 ( .A1(n22875), .A2(n22876), .ZN(n24592) );
  INV_X2 U10613 ( .A(n16822), .ZN(n17707) );
  NAND2_X1 U10614 ( .A1(n12183), .A2(n3604), .ZN(n11731) );
  MUX2_X2 U10615 ( .A(n14229), .B(n14228), .S(n14715), .Z(n16449) );
  NAND2_X1 U10617 ( .A1(n7176), .A2(n7900), .ZN(n7803) );
  NAND2_X1 U10618 ( .A1(n27822), .A2(n27791), .ZN(n26678) );
  XNOR2_X2 U10619 ( .A(n16452), .B(n16451), .ZN(n17829) );
  NAND2_X1 U10620 ( .A1(n14364), .A2(n15514), .ZN(n14389) );
  XNOR2_X1 U10621 ( .A(n3611), .B(n3610), .ZN(Ciphertext[34]) );
  NAND2_X1 U10622 ( .A1(n485), .A2(n23419), .ZN(n23096) );
  NOR2_X1 U10624 ( .A1(n4741), .A2(n26128), .ZN(n4739) );
  OAI21_X1 U10625 ( .B1(n21019), .B2(n22023), .A(n21020), .ZN(n21053) );
  XNOR2_X1 U10626 ( .A(n4579), .B(n19664), .ZN(n4581) );
  NAND3_X1 U10627 ( .A1(n21242), .A2(n21692), .A3(n6314), .ZN(n20961) );
  NAND2_X1 U10628 ( .A1(n13467), .A2(n14033), .ZN(n3613) );
  NAND3_X2 U10629 ( .A1(n3614), .A2(n4421), .A3(n4422), .ZN(n15402) );
  NAND2_X1 U10630 ( .A1(n4424), .A2(n4426), .ZN(n3614) );
  OAI21_X1 U10631 ( .B1(n15337), .B2(n694), .A(n3615), .ZN(n14528) );
  NAND2_X1 U10634 ( .A1(n3617), .A2(n3616), .ZN(n5553) );
  NAND2_X1 U10635 ( .A1(n23387), .A2(n23220), .ZN(n3617) );
  NOR2_X2 U10636 ( .A1(n4542), .A2(n20757), .ZN(n22778) );
  INV_X1 U10638 ( .A(n11198), .ZN(n5917) );
  NAND2_X1 U10639 ( .A1(n3860), .A2(n14373), .ZN(n6050) );
  NAND3_X1 U10640 ( .A1(n24422), .A2(n24420), .A3(n3618), .ZN(n6547) );
  XNOR2_X1 U10642 ( .A(n4990), .B(n16302), .ZN(n4989) );
  OAI21_X1 U10643 ( .B1(n14753), .B2(n15062), .A(n15355), .ZN(n5969) );
  INV_X1 U10644 ( .A(n18111), .ZN(n17729) );
  NAND2_X1 U10647 ( .A1(n24072), .A2(n24666), .ZN(n23914) );
  NAND3_X2 U10648 ( .A1(n3621), .A2(n3620), .A3(n21461), .ZN(n22605) );
  XNOR2_X1 U10651 ( .A(n10268), .B(n10267), .ZN(n6666) );
  INV_X1 U10652 ( .A(n6432), .ZN(n12013) );
  NAND2_X1 U10654 ( .A1(n26496), .A2(n27366), .ZN(n3623) );
  NAND2_X1 U10655 ( .A1(n12304), .A2(n11491), .ZN(n11767) );
  INV_X1 U10656 ( .A(n11003), .ZN(n6779) );
  XNOR2_X1 U10657 ( .A(n13554), .B(n13007), .ZN(n3624) );
  NOR2_X1 U10658 ( .A1(n27368), .A2(n27362), .ZN(n27363) );
  NAND2_X1 U10659 ( .A1(n7093), .A2(n7601), .ZN(n7868) );
  NOR2_X1 U10660 ( .A1(n27152), .A2(n27151), .ZN(n27160) );
  NAND2_X1 U10663 ( .A1(n16613), .A2(n17491), .ZN(n3629) );
  NAND2_X1 U10666 ( .A1(n23758), .A2(n23326), .ZN(n23189) );
  XNOR2_X2 U10667 ( .A(n22344), .B(n22345), .ZN(n23758) );
  NAND2_X1 U10668 ( .A1(n3630), .A2(n24700), .ZN(n3696) );
  NAND2_X1 U10669 ( .A1(n1856), .A2(n24765), .ZN(n24700) );
  NAND2_X1 U10671 ( .A1(n23746), .A2(n23408), .ZN(n3631) );
  AOI21_X1 U10672 ( .B1(n26501), .B2(n27069), .A(n28545), .ZN(n3632) );
  NAND3_X1 U10673 ( .A1(n18015), .A2(n28633), .A3(n17674), .ZN(n17675) );
  NAND2_X1 U10674 ( .A1(n8162), .A2(n7348), .ZN(n7536) );
  NAND2_X1 U10675 ( .A1(n7303), .A2(n7582), .ZN(n7883) );
  NAND2_X1 U10676 ( .A1(n12088), .A2(n11856), .ZN(n3958) );
  NAND3_X1 U10678 ( .A1(n458), .A2(n24455), .A3(n24456), .ZN(n3634) );
  NAND2_X1 U10679 ( .A1(n5170), .A2(n11550), .ZN(n6027) );
  NAND3_X1 U10680 ( .A1(n17563), .A2(n17562), .A3(n532), .ZN(n3839) );
  OR2_X1 U10681 ( .A1(n431), .A2(n12337), .ZN(n12341) );
  NAND2_X1 U10682 ( .A1(n11351), .A2(n10847), .ZN(n3636) );
  NAND3_X1 U10683 ( .A1(n5987), .A2(n5988), .A3(n17067), .ZN(n5986) );
  NAND3_X1 U10684 ( .A1(n14806), .A2(n14769), .A3(n3638), .ZN(n14772) );
  NOR2_X1 U10686 ( .A1(n8525), .A2(n9221), .ZN(n8098) );
  XOR2_X1 U10687 ( .A(n16532), .B(n16533), .Z(n6890) );
  AOI21_X1 U10689 ( .B1(n17589), .B2(n18506), .A(n5392), .ZN(n17590) );
  XNOR2_X1 U10690 ( .A(n25757), .B(n25758), .ZN(n26322) );
  XNOR2_X2 U10691 ( .A(n13571), .B(n13570), .ZN(n14380) );
  NAND3_X1 U10692 ( .A1(n3641), .A2(n5572), .A3(n3640), .ZN(n11944) );
  NAND2_X1 U10693 ( .A1(n10938), .A2(n10937), .ZN(n3641) );
  XNOR2_X2 U10694 ( .A(n16016), .B(n16015), .ZN(n17249) );
  NAND2_X1 U10695 ( .A1(n29301), .A2(n1938), .ZN(n3642) );
  NAND2_X1 U10696 ( .A1(n15107), .A2(n14937), .ZN(n12370) );
  INV_X1 U10698 ( .A(n24725), .ZN(n24730) );
  INV_X1 U10699 ( .A(n7675), .ZN(n7963) );
  OAI211_X1 U10701 ( .C1(n11836), .C2(n12510), .A(n11835), .B(n11834), .ZN(
        n3647) );
  XNOR2_X1 U10706 ( .A(n25429), .B(n25368), .ZN(n3649) );
  OR2_X1 U10707 ( .A1(n3978), .A2(n15259), .ZN(n3977) );
  XNOR2_X1 U10709 ( .A(n10042), .B(n10041), .ZN(n3829) );
  INV_X1 U10710 ( .A(n9037), .ZN(n9031) );
  INV_X1 U10712 ( .A(n10534), .ZN(n11219) );
  INV_X1 U10713 ( .A(n17540), .ZN(n16939) );
  INV_X1 U10714 ( .A(n14630), .ZN(n15387) );
  INV_X1 U10715 ( .A(n3946), .ZN(n11858) );
  OAI21_X1 U10716 ( .B1(n1865), .B2(n10445), .A(n3651), .ZN(n10947) );
  NAND2_X1 U10717 ( .A1(n10940), .A2(n28495), .ZN(n3651) );
  INV_X1 U10719 ( .A(n24768), .ZN(n24427) );
  INV_X1 U10720 ( .A(n17179), .ZN(n4295) );
  OAI21_X1 U10721 ( .B1(n12508), .B2(n3653), .A(n3652), .ZN(n10118) );
  NAND2_X1 U10722 ( .A1(n12508), .A2(n12512), .ZN(n3652) );
  OR2_X1 U10723 ( .A1(n14301), .A2(n13646), .ZN(n13817) );
  AOI21_X1 U10724 ( .B1(n7725), .B2(n7723), .A(n7721), .ZN(n7339) );
  NAND2_X1 U10725 ( .A1(n6727), .A2(n17137), .ZN(n17142) );
  INV_X1 U10726 ( .A(n23377), .ZN(n23202) );
  MUX2_X2 U10727 ( .A(n25197), .B(n25196), .S(n26775), .Z(n27547) );
  NAND2_X1 U10729 ( .A1(n3655), .A2(n7691), .ZN(n5910) );
  NAND3_X1 U10730 ( .A1(n3656), .A2(n7366), .A3(n8207), .ZN(n7365) );
  NAND2_X1 U10731 ( .A1(n8202), .A2(n7634), .ZN(n3656) );
  NOR3_X1 U10733 ( .A1(n21442), .A2(n21653), .A3(n21655), .ZN(n5764) );
  INV_X1 U10734 ( .A(n18972), .ZN(n19989) );
  NAND2_X1 U10735 ( .A1(n12201), .A2(n12200), .ZN(n11703) );
  OR2_X2 U10736 ( .A1(n9257), .A2(n9256), .ZN(n12201) );
  NAND3_X1 U10737 ( .A1(n8039), .A2(n6210), .A3(n7514), .ZN(n7024) );
  AOI21_X1 U10738 ( .B1(n26969), .B2(n3657), .A(n27429), .ZN(n26970) );
  NAND2_X1 U10739 ( .A1(n27420), .A2(n27428), .ZN(n3657) );
  NAND2_X1 U10740 ( .A1(n20789), .A2(n29586), .ZN(n3658) );
  XNOR2_X1 U10741 ( .A(n19130), .B(n18875), .ZN(n3659) );
  MUX2_X1 U10742 ( .A(n28065), .B(n28066), .S(n28064), .Z(n28059) );
  NAND2_X1 U10743 ( .A1(n11640), .A2(n11672), .ZN(n11676) );
  OR2_X1 U10744 ( .A1(n13795), .A2(n14029), .ZN(n4251) );
  AOI22_X2 U10745 ( .A1(n23958), .A2(n23957), .B1(n23959), .B2(n24758), .ZN(
        n25868) );
  INV_X1 U10746 ( .A(n17349), .ZN(n5420) );
  XOR2_X1 U10747 ( .A(n12911), .B(n12912), .Z(n4961) );
  XNOR2_X1 U10748 ( .A(n21996), .B(n21997), .ZN(n23227) );
  NAND2_X1 U10749 ( .A1(n29726), .A2(n24435), .ZN(n23887) );
  NAND2_X1 U10750 ( .A1(n10577), .A2(n432), .ZN(n5278) );
  INV_X1 U10752 ( .A(n11094), .ZN(n5279) );
  XNOR2_X1 U10754 ( .A(n16140), .B(n16139), .ZN(n16142) );
  NAND2_X1 U10755 ( .A1(n13699), .A2(n14292), .ZN(n14298) );
  OAI21_X2 U10756 ( .B1(n11313), .B2(n11312), .A(n11311), .ZN(n4105) );
  AOI22_X1 U10757 ( .A1(n20880), .A2(n21266), .B1(n20879), .B2(n20881), .ZN(
        n20882) );
  INV_X1 U10758 ( .A(n10853), .ZN(n5753) );
  XNOR2_X1 U10759 ( .A(n21994), .B(n4861), .ZN(n22918) );
  NAND2_X1 U10760 ( .A1(n26757), .A2(n26753), .ZN(n25649) );
  OAI22_X1 U10762 ( .A1(n23196), .A2(n23799), .B1(n23319), .B2(n23795), .ZN(
        n21929) );
  OAI21_X1 U10765 ( .B1(n24724), .B2(n24729), .A(n6377), .ZN(n3725) );
  XNOR2_X1 U10766 ( .A(n9618), .B(n9617), .ZN(n10668) );
  INV_X1 U10769 ( .A(n3738), .ZN(n3737) );
  AOI21_X1 U10770 ( .B1(n20799), .B2(n20800), .A(n28916), .ZN(n6346) );
  XNOR2_X1 U10771 ( .A(n9301), .B(n9596), .ZN(n3663) );
  XNOR2_X1 U10772 ( .A(n25512), .B(n25511), .ZN(n27010) );
  INV_X1 U10774 ( .A(n23776), .ZN(n23513) );
  AOI21_X1 U10775 ( .B1(n14013), .B2(n14126), .A(n13060), .ZN(n14014) );
  XNOR2_X1 U10776 ( .A(n19154), .B(n19153), .ZN(n4747) );
  NAND2_X1 U10777 ( .A1(n4868), .A2(n4869), .ZN(n4867) );
  NAND2_X1 U10778 ( .A1(n20532), .A2(n22013), .ZN(n20934) );
  NAND2_X1 U10779 ( .A1(n20086), .A2(n20085), .ZN(n20532) );
  NAND2_X1 U10780 ( .A1(n3665), .A2(n3664), .ZN(n7095) );
  NAND2_X1 U10781 ( .A1(n7093), .A2(n7092), .ZN(n3665) );
  NAND2_X1 U10782 ( .A1(n20935), .A2(n22012), .ZN(n4378) );
  NAND2_X1 U10783 ( .A1(n7363), .A2(n28605), .ZN(n7831) );
  XNOR2_X1 U10784 ( .A(n24330), .B(n26056), .ZN(n24345) );
  OR3_X1 U10786 ( .A1(n7867), .A2(n7092), .A3(n7093), .ZN(n4438) );
  NAND2_X1 U10787 ( .A1(n5838), .A2(n6687), .ZN(n3667) );
  NAND2_X1 U10788 ( .A1(n5370), .A2(n11955), .ZN(n3668) );
  NOR2_X1 U10790 ( .A1(n13654), .A2(n13799), .ZN(n4780) );
  XNOR2_X1 U10791 ( .A(n16119), .B(n16122), .ZN(n3677) );
  NAND2_X1 U10792 ( .A1(n6657), .A2(n11537), .ZN(n6660) );
  OAI21_X1 U10793 ( .B1(n10754), .B2(n11155), .A(n3669), .ZN(n4971) );
  NAND2_X1 U10794 ( .A1(n4972), .A2(n10804), .ZN(n3669) );
  NOR2_X1 U10795 ( .A1(n16820), .A2(n17463), .ZN(n17090) );
  NAND2_X1 U10796 ( .A1(n15458), .A2(n28462), .ZN(n14537) );
  NAND2_X1 U10798 ( .A1(n17067), .A2(n17450), .ZN(n3672) );
  INV_X1 U10799 ( .A(n22902), .ZN(n6818) );
  AOI21_X1 U10801 ( .B1(n3674), .B2(n20496), .A(n20495), .ZN(n21329) );
  NAND2_X1 U10802 ( .A1(n20494), .A2(n29616), .ZN(n3674) );
  NOR3_X1 U10803 ( .A1(n29090), .A2(n27663), .A3(n27671), .ZN(n27195) );
  OAI21_X2 U10804 ( .B1(n27160), .B2(n27159), .A(n27158), .ZN(n27663) );
  NAND2_X1 U10805 ( .A1(n8765), .A2(n8763), .ZN(n8943) );
  NAND2_X1 U10807 ( .A1(n7226), .A2(n7225), .ZN(n3676) );
  INV_X1 U10809 ( .A(n3679), .ZN(n3678) );
  NAND2_X1 U10810 ( .A1(n3680), .A2(n29063), .ZN(n27955) );
  OAI21_X1 U10811 ( .B1(n27970), .B2(n27997), .A(n28456), .ZN(n3680) );
  NAND2_X1 U10813 ( .A1(n27854), .A2(n26641), .ZN(n3681) );
  NAND2_X1 U10814 ( .A1(n14044), .A2(n14045), .ZN(n14049) );
  AOI22_X1 U10815 ( .A1(n15357), .A2(n6674), .B1(n15358), .B2(n15359), .ZN(
        n3682) );
  XNOR2_X1 U10816 ( .A(n2003), .B(n13430), .ZN(n5165) );
  NAND3_X1 U10817 ( .A1(n26643), .A2(n6954), .A3(n26644), .ZN(n26645) );
  NAND2_X1 U10819 ( .A1(n11373), .A2(n12211), .ZN(n3684) );
  NAND2_X1 U10820 ( .A1(n11374), .A2(n6281), .ZN(n3685) );
  INV_X1 U10822 ( .A(n20769), .ZN(n20771) );
  AOI21_X1 U10823 ( .B1(n17354), .B2(n2449), .A(n17031), .ZN(n17199) );
  OAI21_X1 U10824 ( .B1(n21313), .B2(n21312), .A(n5899), .ZN(n5898) );
  XNOR2_X1 U10825 ( .A(n3689), .B(n19193), .ZN(n19197) );
  XNOR2_X1 U10826 ( .A(n3730), .B(n5416), .ZN(n3689) );
  NOR2_X1 U10827 ( .A1(n18709), .A2(n18248), .ZN(n17598) );
  NAND2_X1 U10828 ( .A1(n3691), .A2(n28794), .ZN(n3690) );
  NAND2_X1 U10829 ( .A1(n3693), .A2(n3692), .ZN(n20812) );
  NAND2_X1 U10830 ( .A1(n3694), .A2(n21664), .ZN(n3693) );
  NAND2_X1 U10831 ( .A1(n21662), .A2(n21429), .ZN(n3694) );
  INV_X1 U10832 ( .A(n19765), .ZN(n3911) );
  AOI22_X1 U10833 ( .A1(n27312), .A2(n27873), .B1(n27313), .B2(n27314), .ZN(
        n27323) );
  NAND3_X1 U10834 ( .A1(n20972), .A2(n20703), .A3(n21217), .ZN(n19915) );
  OAI21_X1 U10835 ( .B1(n27041), .B2(n4497), .A(n4496), .ZN(n4495) );
  NAND2_X1 U10836 ( .A1(n23777), .A2(n23776), .ZN(n6423) );
  NOR2_X2 U10837 ( .A1(n3698), .A2(n23485), .ZN(n24777) );
  NAND2_X1 U10838 ( .A1(n23484), .A2(n23483), .ZN(n3699) );
  OAI21_X1 U10839 ( .B1(n18502), .B2(n18501), .A(n515), .ZN(n3701) );
  NAND2_X1 U10841 ( .A1(n17137), .A2(n17138), .ZN(n5471) );
  XOR2_X1 U10842 ( .A(n22055), .B(n22843), .Z(n6100) );
  NAND3_X2 U10843 ( .A1(n3705), .A2(n12889), .A3(n12890), .ZN(n16606) );
  INV_X1 U10844 ( .A(n4073), .ZN(n4072) );
  XNOR2_X1 U10845 ( .A(n13438), .B(n12410), .ZN(n4198) );
  NAND2_X1 U10846 ( .A1(n11351), .A2(n11192), .ZN(n10478) );
  NAND3_X1 U10847 ( .A1(n11914), .A2(n12030), .A3(n12340), .ZN(n11917) );
  NAND2_X1 U10848 ( .A1(n3706), .A2(n8828), .ZN(n8467) );
  OAI211_X2 U10849 ( .C1(n24108), .C2(n24107), .A(n3708), .B(n3707), .ZN(
        n25385) );
  NAND2_X1 U10850 ( .A1(n24105), .A2(n24104), .ZN(n3707) );
  NAND2_X1 U10851 ( .A1(n24106), .A2(n28416), .ZN(n3708) );
  INV_X1 U10853 ( .A(n23978), .ZN(n23981) );
  INV_X1 U10854 ( .A(n13816), .ZN(n14300) );
  INV_X1 U10855 ( .A(n3826), .ZN(n3824) );
  NAND2_X1 U10856 ( .A1(n18495), .A2(n28745), .ZN(n3709) );
  XNOR2_X1 U10857 ( .A(n16185), .B(n3083), .ZN(n16005) );
  NAND2_X1 U10858 ( .A1(n15031), .A2(n14824), .ZN(n15433) );
  OAI21_X1 U10860 ( .B1(n28142), .B2(n17989), .A(n3711), .ZN(n17892) );
  NAND2_X1 U10861 ( .A1(n17989), .A2(n18599), .ZN(n3711) );
  XNOR2_X2 U10863 ( .A(n15710), .B(n15709), .ZN(n17365) );
  INV_X1 U10865 ( .A(n16526), .ZN(n15706) );
  OAI21_X1 U10866 ( .B1(n2762), .B2(n24405), .A(n4081), .ZN(n4176) );
  NAND2_X1 U10867 ( .A1(n4931), .A2(n9209), .ZN(n3718) );
  XNOR2_X1 U10868 ( .A(n6536), .B(n6534), .ZN(n20284) );
  INV_X1 U10869 ( .A(n22919), .ZN(n22574) );
  NOR2_X1 U10870 ( .A1(n23145), .A2(n23460), .ZN(n23356) );
  NAND2_X1 U10871 ( .A1(n26169), .A2(n26786), .ZN(n3720) );
  XNOR2_X1 U10872 ( .A(n3721), .B(n26288), .ZN(Ciphertext[185]) );
  NAND2_X1 U10873 ( .A1(n5214), .A2(n5215), .ZN(n3721) );
  NAND2_X1 U10874 ( .A1(n4839), .A2(n7715), .ZN(n6192) );
  NAND2_X1 U10875 ( .A1(n4644), .A2(n26684), .ZN(n26685) );
  NAND2_X1 U10877 ( .A1(n28064), .A2(n28066), .ZN(n5213) );
  NAND3_X1 U10878 ( .A1(n23030), .A2(n23031), .A3(n23029), .ZN(n23032) );
  OAI22_X1 U10879 ( .A1(n18456), .A2(n18106), .B1(n18109), .B2(n18111), .ZN(
        n17730) );
  XNOR2_X1 U10880 ( .A(n3724), .B(n12892), .ZN(n12871) );
  XNOR2_X1 U10881 ( .A(n12865), .B(n12866), .ZN(n3724) );
  NAND2_X1 U10883 ( .A1(n18261), .A2(n18326), .ZN(n4059) );
  INV_X1 U10884 ( .A(n21183), .ZN(n21129) );
  INV_X1 U10886 ( .A(n3726), .ZN(n6407) );
  OAI21_X1 U10887 ( .B1(n23333), .B2(n6462), .A(n23332), .ZN(n3726) );
  NAND3_X1 U10890 ( .A1(n17417), .A2(n17418), .A3(n17419), .ZN(n18402) );
  NAND3_X1 U10891 ( .A1(n10850), .A2(n10848), .A3(n4123), .ZN(n12158) );
  NAND3_X1 U10894 ( .A1(n17489), .A2(n17148), .A3(n17078), .ZN(n4653) );
  NAND2_X1 U10896 ( .A1(n16008), .A2(n1880), .ZN(n3729) );
  NOR2_X1 U10897 ( .A1(n294), .A2(n27213), .ZN(n6809) );
  NAND2_X1 U10899 ( .A1(n24891), .A2(n24532), .ZN(n6865) );
  XNOR2_X1 U10900 ( .A(n19192), .B(n3598), .ZN(n3730) );
  INV_X1 U10901 ( .A(n11462), .ZN(n11461) );
  OAI22_X1 U10902 ( .A1(n10803), .A2(n28559), .B1(n10553), .B2(n11158), .ZN(
        n10496) );
  NOR2_X1 U10903 ( .A1(n11941), .A2(n11942), .ZN(n3732) );
  NAND2_X1 U10904 ( .A1(n29573), .A2(n26278), .ZN(n26392) );
  NAND2_X1 U10905 ( .A1(n5064), .A2(n13909), .ZN(n6813) );
  INV_X1 U10907 ( .A(n3734), .ZN(n3733) );
  OAI21_X1 U10908 ( .B1(n13992), .B2(n15692), .A(n13990), .ZN(n3734) );
  NAND2_X1 U10910 ( .A1(n3735), .A2(n28526), .ZN(n19752) );
  NOR2_X1 U10912 ( .A1(n27150), .A2(n6592), .ZN(n6591) );
  NAND2_X1 U10913 ( .A1(n7244), .A2(n7648), .ZN(n3736) );
  OAI21_X1 U10914 ( .B1(n1801), .B2(n16383), .A(n16382), .ZN(n3738) );
  NAND3_X1 U10915 ( .A1(n4652), .A2(n4651), .A3(n29294), .ZN(n3739) );
  INV_X1 U10916 ( .A(n20977), .ZN(n21367) );
  INV_X1 U10917 ( .A(n8395), .ZN(n8396) );
  NOR2_X1 U10918 ( .A1(n23067), .A2(n4429), .ZN(n4459) );
  XOR2_X1 U10919 ( .A(n20655), .B(n20654), .Z(n4430) );
  NAND3_X1 U10920 ( .A1(n5267), .A2(n5265), .A3(n10976), .ZN(n10978) );
  NAND2_X1 U10921 ( .A1(n18354), .A2(n18312), .ZN(n6030) );
  NOR2_X1 U10922 ( .A1(n580), .A2(n12350), .ZN(n5133) );
  OAI22_X1 U10923 ( .A1(n28183), .A2(n29157), .B1(n23722), .B2(n23843), .ZN(
        n22127) );
  OR2_X1 U10924 ( .A1(n18340), .A2(n514), .ZN(n4244) );
  NAND2_X1 U10926 ( .A1(n3741), .A2(n14142), .ZN(n14143) );
  AND2_X1 U10928 ( .A1(n20349), .A2(n20510), .ZN(n5853) );
  INV_X1 U10929 ( .A(n18520), .ZN(n19262) );
  INV_X1 U10930 ( .A(n5953), .ZN(n21561) );
  INV_X1 U10931 ( .A(n10502), .ZN(n5672) );
  INV_X1 U10932 ( .A(n12186), .ZN(n4028) );
  XNOR2_X1 U10934 ( .A(n19598), .B(n18720), .ZN(n5211) );
  NAND3_X1 U10935 ( .A1(n474), .A2(n29544), .A3(n23169), .ZN(n23170) );
  NAND2_X1 U10936 ( .A1(n8511), .A2(n8914), .ZN(n9105) );
  NAND2_X1 U10937 ( .A1(n11132), .A2(n10711), .ZN(n10501) );
  NAND2_X1 U10939 ( .A1(n12264), .A2(n575), .ZN(n3745) );
  NAND2_X1 U10940 ( .A1(n8800), .A2(n8802), .ZN(n8957) );
  INV_X1 U10941 ( .A(n14702), .ZN(n3748) );
  NAND2_X1 U10942 ( .A1(n14851), .A2(n15310), .ZN(n5948) );
  NAND2_X1 U10943 ( .A1(n5928), .A2(n21088), .ZN(n5926) );
  MUX2_X2 U10944 ( .A(n22051), .B(n22050), .S(n28796), .Z(n24584) );
  OR2_X1 U10945 ( .A1(n7614), .A2(n7393), .ZN(n7930) );
  OR2_X1 U10946 ( .A1(n20784), .A2(n21177), .ZN(n5087) );
  XOR2_X1 U10947 ( .A(n20797), .B(n22383), .Z(n5452) );
  NOR2_X1 U10948 ( .A1(n6530), .A2(n21031), .ZN(n6527) );
  XNOR2_X1 U10949 ( .A(n26103), .B(n26100), .ZN(n6018) );
  NAND2_X1 U10950 ( .A1(n27186), .A2(n26397), .ZN(n3754) );
  NAND2_X1 U10951 ( .A1(n15502), .A2(n15265), .ZN(n14924) );
  NAND3_X2 U10952 ( .A1(n3757), .A2(n6402), .A3(n3756), .ZN(n19726) );
  NAND2_X1 U10953 ( .A1(n18328), .A2(n18329), .ZN(n3756) );
  INV_X1 U10955 ( .A(n21563), .ZN(n3759) );
  NOR2_X1 U10956 ( .A1(n21564), .A2(n28155), .ZN(n3760) );
  OAI21_X1 U10957 ( .B1(n20500), .B2(n29601), .A(n20498), .ZN(n3761) );
  AOI21_X1 U10958 ( .B1(n21156), .B2(n3762), .A(n494), .ZN(n4755) );
  NAND2_X1 U10960 ( .A1(n3764), .A2(n3763), .ZN(n5899) );
  INV_X1 U10961 ( .A(n21311), .ZN(n3763) );
  NAND2_X1 U10962 ( .A1(n29530), .A2(n21309), .ZN(n3764) );
  NAND2_X1 U10963 ( .A1(n6132), .A2(n12286), .ZN(n3765) );
  XNOR2_X1 U10964 ( .A(n1895), .B(n10184), .ZN(n6136) );
  OAI21_X1 U10965 ( .B1(n18711), .B2(n18709), .A(n3766), .ZN(n18714) );
  OAI21_X1 U10971 ( .B1(n9232), .B2(n9229), .A(n3773), .ZN(n9046) );
  NAND2_X1 U10972 ( .A1(n9232), .A2(n9233), .ZN(n3773) );
  OAI21_X1 U10973 ( .B1(n7695), .B2(n8227), .A(n3774), .ZN(n6991) );
  NAND2_X1 U10974 ( .A1(n7695), .A2(n8222), .ZN(n3774) );
  OR2_X2 U10975 ( .A1(n10596), .A2(n10595), .ZN(n12359) );
  XNOR2_X1 U10976 ( .A(n3775), .B(n22504), .ZN(n22991) );
  XNOR2_X1 U10977 ( .A(n6388), .B(n6389), .ZN(n3775) );
  AOI21_X1 U10978 ( .B1(n11612), .B2(n11613), .A(n566), .ZN(n5465) );
  NOR2_X1 U10980 ( .A1(n11140), .A2(n3829), .ZN(n10721) );
  AOI21_X1 U10983 ( .B1(n15078), .B2(n5229), .A(n3778), .ZN(n3777) );
  NOR2_X1 U10984 ( .A1(n14876), .A2(n15082), .ZN(n3778) );
  NAND3_X1 U10985 ( .A1(n5546), .A2(n26768), .A3(n26771), .ZN(n25158) );
  NAND2_X1 U10986 ( .A1(n6556), .A2(n24020), .ZN(n24002) );
  XOR2_X1 U10987 ( .A(n25389), .B(n25388), .Z(n6071) );
  XNOR2_X1 U10988 ( .A(n3779), .B(n19175), .ZN(n18785) );
  XNOR2_X1 U10989 ( .A(n18783), .B(n19331), .ZN(n3779) );
  NAND2_X1 U10990 ( .A1(n6734), .A2(n6737), .ZN(n26495) );
  NAND2_X1 U10992 ( .A1(n26497), .A2(n27364), .ZN(n25997) );
  INV_X1 U10993 ( .A(n18170), .ZN(n5200) );
  NAND2_X1 U10994 ( .A1(n23364), .A2(n23672), .ZN(n23362) );
  NAND2_X2 U10995 ( .A1(n6115), .A2(n20685), .ZN(n22890) );
  XNOR2_X1 U10998 ( .A(n16059), .B(n16649), .ZN(n15608) );
  NAND3_X2 U10999 ( .A1(n14022), .A2(n14023), .A3(n3782), .ZN(n16059) );
  NAND2_X1 U11000 ( .A1(n27071), .A2(n26614), .ZN(n3785) );
  NAND2_X1 U11001 ( .A1(n27070), .A2(n29520), .ZN(n3786) );
  XNOR2_X1 U11003 ( .A(n16201), .B(n16200), .ZN(n6869) );
  XNOR2_X1 U11004 ( .A(n13355), .B(n4490), .ZN(n13356) );
  OAI22_X1 U11005 ( .A1(n20397), .A2(n20396), .B1(n20395), .B2(n20394), .ZN(
        n5871) );
  INV_X1 U11006 ( .A(n19277), .ZN(n18369) );
  NAND2_X1 U11007 ( .A1(n4429), .A2(n23067), .ZN(n23348) );
  NAND2_X1 U11008 ( .A1(n6450), .A2(n3788), .ZN(n10372) );
  NAND3_X1 U11009 ( .A1(n7659), .A2(n8305), .A3(n3790), .ZN(n7402) );
  NAND2_X1 U11010 ( .A1(n8302), .A2(n7657), .ZN(n3790) );
  AND3_X2 U11011 ( .A1(n3836), .A2(n24781), .A3(n24782), .ZN(n25191) );
  NAND2_X1 U11014 ( .A1(n17480), .A2(n17477), .ZN(n3884) );
  INV_X1 U11016 ( .A(n26682), .ZN(n26710) );
  INV_X1 U11017 ( .A(n28395), .ZN(n14890) );
  XNOR2_X1 U11018 ( .A(n3792), .B(n16024), .ZN(n16555) );
  XNOR2_X1 U11019 ( .A(n28395), .B(n16199), .ZN(n15673) );
  AND2_X1 U11020 ( .A1(n7792), .A2(n7793), .ZN(n7795) );
  OAI21_X1 U11021 ( .B1(n7797), .B2(n28149), .A(n3793), .ZN(n7798) );
  NAND3_X1 U11022 ( .A1(n7284), .A2(n7792), .A3(n7793), .ZN(n3793) );
  NAND3_X1 U11023 ( .A1(n12990), .A2(n12090), .A3(n3796), .ZN(n3794) );
  NAND2_X1 U11024 ( .A1(n3961), .A2(n12151), .ZN(n12090) );
  NAND2_X1 U11025 ( .A1(n3797), .A2(n24405), .ZN(n23503) );
  NAND2_X1 U11026 ( .A1(n24085), .A2(n3797), .ZN(n23880) );
  NAND2_X1 U11028 ( .A1(n3799), .A2(n3798), .ZN(n5834) );
  NAND2_X1 U11030 ( .A1(n10983), .A2(n10982), .ZN(n10696) );
  INV_X1 U11032 ( .A(n10980), .ZN(n3804) );
  INV_X1 U11033 ( .A(n10980), .ZN(n10783) );
  NAND2_X1 U11034 ( .A1(n10988), .A2(n10985), .ZN(n3805) );
  NAND2_X1 U11035 ( .A1(n13968), .A2(n3806), .ZN(n13969) );
  INV_X1 U11036 ( .A(n12711), .ZN(n3806) );
  MUX2_X1 U11037 ( .A(n14459), .B(n4290), .S(n12711), .Z(n13683) );
  NAND3_X1 U11039 ( .A1(n19947), .A2(n20200), .A3(n20305), .ZN(n3808) );
  NAND3_X1 U11040 ( .A1(n8147), .A2(n7793), .A3(n7796), .ZN(n7286) );
  NAND3_X1 U11041 ( .A1(n7541), .A2(n8148), .A3(n3810), .ZN(n7354) );
  NAND2_X1 U11044 ( .A1(n16611), .A2(n18356), .ZN(n17920) );
  XNOR2_X1 U11045 ( .A(n16170), .B(n16279), .ZN(n3813) );
  NOR2_X2 U11046 ( .A1(n15340), .A2(n15341), .ZN(n16170) );
  INV_X1 U11047 ( .A(n11252), .ZN(n3817) );
  NAND2_X1 U11048 ( .A1(n11251), .A2(n3816), .ZN(n3815) );
  NAND2_X1 U11049 ( .A1(n11033), .A2(n11252), .ZN(n3818) );
  NOR2_X1 U11050 ( .A1(n11033), .A2(n3820), .ZN(n3819) );
  NAND3_X1 U11053 ( .A1(n6203), .A2(n5783), .A3(n4245), .ZN(n21065) );
  NAND2_X1 U11055 ( .A1(n3824), .A2(n18486), .ZN(n3823) );
  NAND2_X1 U11056 ( .A1(n18490), .A2(n18489), .ZN(n3826) );
  AOI22_X1 U11057 ( .A1(n15289), .A2(n15291), .B1(n15290), .B2(n3827), .ZN(
        n15298) );
  NAND2_X1 U11058 ( .A1(n3827), .A2(n14517), .ZN(n15215) );
  OAI21_X1 U11059 ( .B1(n15217), .B2(n15290), .A(n3827), .ZN(n15041) );
  OAI211_X1 U11061 ( .C1(n15217), .C2(n3827), .A(n15293), .B(n15292), .ZN(
        n14110) );
  OAI21_X1 U11062 ( .B1(n15289), .B2(n3827), .A(n14097), .ZN(n4957) );
  NAND2_X1 U11063 ( .A1(n11138), .A2(n3828), .ZN(n10719) );
  NAND2_X1 U11064 ( .A1(n11139), .A2(n3829), .ZN(n10923) );
  NAND2_X1 U11065 ( .A1(n10103), .A2(n3829), .ZN(n10106) );
  NAND2_X1 U11066 ( .A1(n5531), .A2(n13914), .ZN(n3830) );
  NAND2_X1 U11067 ( .A1(n17713), .A2(n18329), .ZN(n3831) );
  MUX2_X1 U11068 ( .A(n27106), .B(n27701), .S(n27702), .Z(n27107) );
  MUX2_X1 U11069 ( .A(n27162), .B(n27163), .S(n27702), .Z(n27164) );
  INV_X1 U11071 ( .A(n25133), .ZN(n3837) );
  XNOR2_X1 U11072 ( .A(n25191), .B(n24897), .ZN(n24898) );
  NAND2_X1 U11073 ( .A1(n3838), .A2(n21124), .ZN(n21461) );
  NOR2_X1 U11074 ( .A1(n3838), .A2(n21459), .ZN(n21460) );
  NOR2_X1 U11075 ( .A1(n1814), .A2(n3838), .ZN(n20843) );
  NAND2_X1 U11076 ( .A1(n3784), .A2(n15008), .ZN(n14867) );
  INV_X1 U11077 ( .A(n15373), .ZN(n15008) );
  NOR2_X1 U11078 ( .A1(n15373), .A2(n15374), .ZN(n3841) );
  NAND2_X1 U11079 ( .A1(n12508), .A2(n11990), .ZN(n3842) );
  NAND2_X1 U11080 ( .A1(n3842), .A2(n12507), .ZN(n11521) );
  OAI21_X1 U11081 ( .B1(n15471), .B2(n14551), .A(n15472), .ZN(n3845) );
  NAND2_X1 U11082 ( .A1(n1848), .A2(n15168), .ZN(n15472) );
  INV_X1 U11085 ( .A(n13866), .ZN(n3846) );
  NAND2_X1 U11086 ( .A1(n522), .A2(n17969), .ZN(n3848) );
  OR2_X1 U11089 ( .A1(n14209), .A2(n3851), .ZN(n3850) );
  NAND2_X1 U11090 ( .A1(n3853), .A2(n3852), .ZN(n3855) );
  NAND2_X1 U11091 ( .A1(n20228), .A2(n20227), .ZN(n3853) );
  NAND2_X1 U11092 ( .A1(n3854), .A2(n21439), .ZN(n21441) );
  AND2_X1 U11093 ( .A1(n3855), .A2(n21438), .ZN(n3854) );
  XNOR2_X1 U11094 ( .A(n3856), .B(n16585), .ZN(n15631) );
  XNOR2_X1 U11095 ( .A(n3856), .B(n16085), .ZN(n16243) );
  OR2_X1 U11096 ( .A1(n13725), .A2(n3860), .ZN(n13724) );
  AND2_X1 U11097 ( .A1(n3860), .A2(n13725), .ZN(n13440) );
  NAND2_X1 U11098 ( .A1(n14146), .A2(n3860), .ZN(n4331) );
  NAND2_X1 U11099 ( .A1(n5404), .A2(n3860), .ZN(n5403) );
  NAND2_X1 U11100 ( .A1(n5405), .A2(n3859), .ZN(n14009) );
  OAI21_X1 U11102 ( .B1(n3862), .B2(n11135), .A(n3861), .ZN(n3863) );
  NAND2_X1 U11103 ( .A1(n11136), .A2(n11135), .ZN(n3861) );
  NOR2_X2 U11104 ( .A1(n10766), .A2(n10767), .ZN(n11881) );
  OR2_X1 U11106 ( .A1(n18109), .A2(n17902), .ZN(n3866) );
  OAI21_X1 U11108 ( .B1(n3868), .B2(n3867), .A(n14157), .ZN(n14550) );
  NAND2_X1 U11109 ( .A1(n3869), .A2(n14158), .ZN(n14549) );
  NAND2_X1 U11110 ( .A1(n13847), .A2(n13936), .ZN(n3869) );
  XNOR2_X1 U11111 ( .A(n13444), .B(n13493), .ZN(n3870) );
  XNOR2_X1 U11112 ( .A(n12699), .B(n3871), .ZN(n12701) );
  XNOR2_X1 U11113 ( .A(n3871), .B(n3232), .ZN(n13239) );
  NAND3_X1 U11115 ( .A1(n3873), .A2(n29517), .A3(n11207), .ZN(n11208) );
  NAND2_X1 U11116 ( .A1(n11090), .A2(n3873), .ZN(n10576) );
  NAND2_X1 U11117 ( .A1(n432), .A2(n3873), .ZN(n11092) );
  NAND3_X1 U11118 ( .A1(n10431), .A2(n6164), .A3(n3873), .ZN(n6163) );
  INV_X1 U11119 ( .A(n11094), .ZN(n3873) );
  NAND3_X1 U11120 ( .A1(n3875), .A2(n512), .A3(n17823), .ZN(n3874) );
  NAND2_X1 U11122 ( .A1(n1530), .A2(n29594), .ZN(n3877) );
  INV_X1 U11123 ( .A(n3880), .ZN(n17265) );
  NAND2_X1 U11125 ( .A1(n3880), .A2(n29299), .ZN(n17267) );
  NAND2_X1 U11126 ( .A1(n16864), .A2(n3880), .ZN(n3879) );
  NAND2_X1 U11128 ( .A1(n6045), .A2(n14368), .ZN(n3881) );
  NAND2_X1 U11130 ( .A1(n17479), .A2(n17478), .ZN(n3885) );
  INV_X1 U11131 ( .A(n3887), .ZN(n23656) );
  NAND2_X1 U11132 ( .A1(n4231), .A2(n3887), .ZN(n4851) );
  OR2_X1 U11133 ( .A1(n20840), .A2(n3887), .ZN(n4770) );
  OAI22_X1 U11134 ( .A1(n23352), .A2(n3887), .B1(n23545), .B2(n4232), .ZN(
        n4648) );
  NAND2_X1 U11135 ( .A1(n23142), .A2(n4772), .ZN(n3886) );
  NAND2_X1 U11136 ( .A1(n3888), .A2(n12231), .ZN(n12230) );
  NAND2_X1 U11137 ( .A1(n12227), .A2(n12226), .ZN(n3888) );
  NAND2_X1 U11138 ( .A1(n3890), .A2(n5339), .ZN(n3889) );
  INV_X1 U11139 ( .A(n21030), .ZN(n3890) );
  NAND2_X1 U11140 ( .A1(n3892), .A2(n22146), .ZN(n3891) );
  OAI21_X1 U11141 ( .B1(n20418), .B2(n20192), .A(n5334), .ZN(n3893) );
  NAND2_X1 U11142 ( .A1(n19748), .A2(n19749), .ZN(n3894) );
  OR2_X1 U11143 ( .A1(n308), .A2(n14366), .ZN(n4812) );
  NAND2_X1 U11144 ( .A1(n559), .A2(n6000), .ZN(n3895) );
  AOI21_X1 U11145 ( .B1(n308), .B2(n14123), .A(n14366), .ZN(n3896) );
  XNOR2_X2 U11146 ( .A(n12953), .B(n12952), .ZN(n14366) );
  XNOR2_X1 U11147 ( .A(n3898), .B(n3897), .ZN(Ciphertext[73]) );
  INV_X1 U11148 ( .A(n27546), .ZN(n3899) );
  AND2_X1 U11149 ( .A1(n27549), .A2(n27203), .ZN(n27199) );
  NAND2_X1 U11150 ( .A1(n28604), .A2(n23673), .ZN(n3902) );
  AOI22_X2 U11151 ( .A1(n3903), .A2(n21678), .B1(n21082), .B2(n21081), .ZN(
        n22199) );
  INV_X1 U11152 ( .A(n11322), .ZN(n11187) );
  INV_X1 U11153 ( .A(n5595), .ZN(n11181) );
  AOI21_X1 U11154 ( .B1(n11162), .B2(n6411), .A(n3904), .ZN(n3910) );
  AOI21_X1 U11155 ( .B1(n3909), .B2(n11053), .A(n1933), .ZN(n3908) );
  OAI211_X2 U11156 ( .C1(n3907), .C2(n11322), .A(n3906), .B(n3905), .ZN(n11195) );
  NAND2_X1 U11158 ( .A1(n11164), .A2(n11165), .ZN(n3909) );
  OR2_X1 U11159 ( .A1(n17199), .A2(n17198), .ZN(n3914) );
  NAND3_X1 U11160 ( .A1(n18413), .A2(n3915), .A3(n28688), .ZN(n6101) );
  NAND2_X1 U11162 ( .A1(n17340), .A2(n17336), .ZN(n6337) );
  NAND2_X1 U11163 ( .A1(n3918), .A2(n3921), .ZN(n3917) );
  NAND2_X1 U11164 ( .A1(n3922), .A2(n14893), .ZN(n3921) );
  INV_X1 U11165 ( .A(n14937), .ZN(n15409) );
  NOR2_X1 U11166 ( .A1(n15224), .A2(n15342), .ZN(n3924) );
  MUX2_X1 U11167 ( .A(n15222), .B(n15343), .S(n15046), .Z(n3926) );
  NAND3_X1 U11170 ( .A1(n14162), .A2(n14163), .A3(n14161), .ZN(n3927) );
  NAND2_X1 U11171 ( .A1(n14160), .A2(n14159), .ZN(n3928) );
  INV_X1 U11172 ( .A(n7696), .ZN(n3930) );
  NAND2_X1 U11173 ( .A1(n7424), .A2(n7822), .ZN(n7696) );
  NAND2_X1 U11174 ( .A1(n3930), .A2(n7827), .ZN(n3929) );
  NAND3_X1 U11175 ( .A1(n18416), .A2(n18413), .A3(n3932), .ZN(n3931) );
  XNOR2_X1 U11177 ( .A(n15698), .B(n5798), .ZN(n3938) );
  NAND2_X1 U11178 ( .A1(n3939), .A2(n2052), .ZN(n17343) );
  NAND2_X1 U11179 ( .A1(n17155), .A2(n17204), .ZN(n17156) );
  NAND2_X1 U11180 ( .A1(n17337), .A2(n17336), .ZN(n3939) );
  INV_X1 U11181 ( .A(n10945), .ZN(n3941) );
  NAND2_X1 U11182 ( .A1(n3946), .A2(n11944), .ZN(n11665) );
  NAND2_X1 U11183 ( .A1(n10947), .A2(n10946), .ZN(n3942) );
  NAND3_X1 U11184 ( .A1(n11948), .A2(n3946), .A3(n11945), .ZN(n11946) );
  NAND3_X1 U11185 ( .A1(n11947), .A2(n3946), .A3(n11948), .ZN(n11949) );
  NAND2_X1 U11186 ( .A1(n11857), .A2(n3943), .ZN(n10954) );
  AND2_X1 U11187 ( .A1(n11952), .A2(n3946), .ZN(n3943) );
  NAND2_X1 U11188 ( .A1(n11556), .A2(n3945), .ZN(n3944) );
  AND2_X1 U11189 ( .A1(n11943), .A2(n3946), .ZN(n3945) );
  INV_X1 U11190 ( .A(n14346), .ZN(n14136) );
  NAND2_X1 U11192 ( .A1(n14134), .A2(n3948), .ZN(n3947) );
  OR2_X1 U11193 ( .A1(n14346), .A2(n3949), .ZN(n3948) );
  NAND2_X1 U11194 ( .A1(n13842), .A2(n14010), .ZN(n3949) );
  INV_X1 U11195 ( .A(n13843), .ZN(n3950) );
  NAND2_X1 U11196 ( .A1(n20633), .A2(n28538), .ZN(n3954) );
  NAND2_X1 U11197 ( .A1(n20456), .A2(n1908), .ZN(n3951) );
  INV_X1 U11198 ( .A(n20453), .ZN(n20633) );
  XNOR2_X1 U11199 ( .A(n12420), .B(n13175), .ZN(n13287) );
  NAND2_X1 U11201 ( .A1(n3962), .A2(n12151), .ZN(n3955) );
  NAND2_X1 U11202 ( .A1(n3957), .A2(n12991), .ZN(n3956) );
  NAND2_X1 U11203 ( .A1(n12994), .A2(n3958), .ZN(n3957) );
  NAND2_X1 U11205 ( .A1(n430), .A2(n579), .ZN(n3960) );
  NOR2_X1 U11206 ( .A1(n12150), .A2(n3961), .ZN(n3962) );
  INV_X1 U11207 ( .A(n12088), .ZN(n3961) );
  NAND4_X1 U11208 ( .A1(n4843), .A2(n3966), .A3(n3965), .A4(n3963), .ZN(n4842)
         );
  NOR2_X1 U11209 ( .A1(n12200), .A2(n12201), .ZN(n3964) );
  NAND2_X1 U11210 ( .A1(n12202), .A2(n4844), .ZN(n3965) );
  NAND2_X1 U11211 ( .A1(n12201), .A2(n12203), .ZN(n3966) );
  INV_X1 U11212 ( .A(n3968), .ZN(n3967) );
  OAI21_X1 U11213 ( .B1(n19794), .B2(n20517), .A(n3969), .ZN(n3968) );
  INV_X1 U11216 ( .A(n20584), .ZN(n3973) );
  OAI21_X1 U11217 ( .B1(n20590), .B2(n3975), .A(n20589), .ZN(n21135) );
  NAND2_X1 U11218 ( .A1(n20590), .A2(n20589), .ZN(n3971) );
  NAND2_X1 U11219 ( .A1(n3975), .A2(n20589), .ZN(n3972) );
  INV_X1 U11220 ( .A(n19828), .ZN(n3975) );
  NAND2_X1 U11221 ( .A1(n14258), .A2(n6921), .ZN(n3976) );
  NAND2_X1 U11222 ( .A1(n14761), .A2(n15260), .ZN(n3978) );
  NAND3_X1 U11223 ( .A1(n29737), .A2(n4246), .A3(n1666), .ZN(n3980) );
  XNOR2_X1 U11225 ( .A(n22100), .B(n3984), .ZN(n3983) );
  INV_X1 U11226 ( .A(n22655), .ZN(n3984) );
  NAND2_X1 U11227 ( .A1(n23437), .A2(n23436), .ZN(n3985) );
  MUX2_X1 U11228 ( .A(n24972), .B(n24973), .S(n24509), .Z(n23600) );
  NAND3_X1 U11230 ( .A1(n574), .A2(n11922), .A3(n11549), .ZN(n3987) );
  AOI21_X1 U11231 ( .B1(n11547), .B2(n11922), .A(n11927), .ZN(n3989) );
  NAND2_X1 U11233 ( .A1(n2968), .A2(n10919), .ZN(n3992) );
  OAI21_X1 U11234 ( .B1(n18277), .B2(n3995), .A(n3993), .ZN(n3996) );
  NAND2_X1 U11235 ( .A1(n3994), .A2(n18277), .ZN(n3993) );
  INV_X1 U11236 ( .A(n18204), .ZN(n3994) );
  AOI22_X2 U11237 ( .A1(n18206), .A2(n3997), .B1(n3996), .B2(n18279), .ZN(
        n19194) );
  NAND2_X1 U11239 ( .A1(n18275), .A2(n17696), .ZN(n3997) );
  NAND2_X1 U11240 ( .A1(n578), .A2(n11869), .ZN(n3998) );
  NAND2_X1 U11241 ( .A1(n6181), .A2(n11500), .ZN(n11750) );
  NAND2_X1 U11242 ( .A1(n11868), .A2(n11867), .ZN(n3999) );
  NAND2_X1 U11244 ( .A1(n373), .A2(n4002), .ZN(n5328) );
  NAND2_X1 U11245 ( .A1(n29620), .A2(n23762), .ZN(n23476) );
  NAND2_X1 U11246 ( .A1(n23759), .A2(n29620), .ZN(n5743) );
  XNOR2_X1 U11247 ( .A(n15946), .B(n15945), .ZN(n17276) );
  NAND3_X1 U11249 ( .A1(n17271), .A2(n17275), .A3(n6465), .ZN(n4004) );
  OAI211_X1 U11250 ( .C1(n414), .C2(n20089), .A(n4007), .B(n4006), .ZN(n20095)
         );
  NAND2_X1 U11251 ( .A1(n4008), .A2(n29104), .ZN(n4007) );
  NAND2_X1 U11252 ( .A1(n20039), .A2(n29114), .ZN(n4008) );
  XNOR2_X2 U11254 ( .A(n18717), .B(n18716), .ZN(n20041) );
  AOI22_X1 U11255 ( .A1(n4012), .A2(n4010), .B1(n2549), .B2(n4009), .ZN(n13708) );
  NAND2_X1 U11256 ( .A1(n21078), .A2(n20933), .ZN(n21077) );
  NAND2_X1 U11257 ( .A1(n4015), .A2(n4014), .ZN(n4013) );
  NAND3_X1 U11258 ( .A1(n26450), .A2(n26179), .A3(n26447), .ZN(n4014) );
  NAND2_X1 U11259 ( .A1(n25625), .A2(n26456), .ZN(n4015) );
  AOI22_X2 U11260 ( .A1(n16956), .A2(n16955), .B1(n16957), .B2(n18259), .ZN(
        n19085) );
  NAND3_X1 U11261 ( .A1(n6706), .A2(n4341), .A3(n571), .ZN(n4016) );
  NAND2_X1 U11263 ( .A1(n11180), .A2(n11179), .ZN(n11955) );
  XNOR2_X1 U11264 ( .A(n6939), .B(n22667), .ZN(n23305) );
  INV_X1 U11265 ( .A(n11982), .ZN(n13083) );
  OAI21_X1 U11266 ( .B1(n11811), .B2(n4021), .A(n11810), .ZN(n11814) );
  MUX2_X1 U11269 ( .A(n7665), .B(n8264), .S(n8270), .Z(n4022) );
  XNOR2_X2 U11270 ( .A(Key[146]), .B(Plaintext[146]), .ZN(n8270) );
  AOI21_X1 U11271 ( .B1(n10507), .B2(n4023), .A(n11124), .ZN(n10508) );
  NAND2_X1 U11272 ( .A1(n4024), .A2(n11120), .ZN(n4023) );
  INV_X1 U11273 ( .A(n11123), .ZN(n4024) );
  XNOR2_X2 U11274 ( .A(n9885), .B(n9884), .ZN(n11123) );
  OR2_X1 U11275 ( .A1(n6095), .A2(n27525), .ZN(n27510) );
  OAI21_X1 U11277 ( .B1(n27510), .B2(n27531), .A(n3067), .ZN(n27511) );
  INV_X1 U11278 ( .A(n24677), .ZN(n24322) );
  NAND2_X1 U11279 ( .A1(n20324), .A2(n20109), .ZN(n20321) );
  XNOR2_X2 U11280 ( .A(n19589), .B(n19588), .ZN(n20109) );
  INV_X1 U11281 ( .A(n14487), .ZN(n12120) );
  OAI21_X1 U11282 ( .B1(n14167), .B2(n14164), .A(n4027), .ZN(n4026) );
  NAND3_X1 U11283 ( .A1(n12120), .A2(n14484), .A3(n29565), .ZN(n4027) );
  NAND2_X1 U11284 ( .A1(n4028), .A2(n2483), .ZN(n12195) );
  NAND2_X1 U11285 ( .A1(n4028), .A2(n12128), .ZN(n11727) );
  OR2_X1 U11287 ( .A1(n12127), .A2(n4028), .ZN(n4982) );
  XNOR2_X1 U11288 ( .A(n4031), .B(n2505), .ZN(n12848) );
  XNOR2_X1 U11289 ( .A(n4031), .B(n13414), .ZN(n12908) );
  XNOR2_X1 U11290 ( .A(n4031), .B(n13269), .ZN(n13412) );
  XNOR2_X1 U11291 ( .A(n12826), .B(n4031), .ZN(n12829) );
  XNOR2_X1 U11292 ( .A(n12780), .B(n4031), .ZN(n12117) );
  XNOR2_X1 U11293 ( .A(n12637), .B(n4031), .ZN(n12385) );
  OAI211_X2 U11294 ( .C1(n12115), .C2(n12114), .A(n12113), .B(n12112), .ZN(
        n4031) );
  NOR2_X1 U11297 ( .A1(n27380), .A2(n28394), .ZN(n4035) );
  INV_X1 U11298 ( .A(n26610), .ZN(n4036) );
  NOR2_X1 U11299 ( .A1(n4038), .A2(n12211), .ZN(n9655) );
  MUX2_X1 U11302 ( .A(n14808), .B(n14810), .S(n14775), .Z(n14229) );
  NAND2_X1 U11303 ( .A1(n11428), .A2(n11426), .ZN(n4046) );
  INV_X1 U11304 ( .A(n14192), .ZN(n14395) );
  OR2_X1 U11305 ( .A1(n14393), .A2(n14192), .ZN(n14195) );
  OAI211_X1 U11306 ( .C1(n28805), .C2(n14395), .A(n14393), .B(n4047), .ZN(
        n4048) );
  NOR2_X1 U11308 ( .A1(n14192), .A2(n14194), .ZN(n4049) );
  OR2_X1 U11309 ( .A1(n7116), .A2(n7320), .ZN(n4052) );
  NAND2_X1 U11310 ( .A1(n20252), .A2(n1951), .ZN(n4053) );
  NAND2_X1 U11311 ( .A1(n21631), .A2(n21036), .ZN(n21039) );
  INV_X1 U11312 ( .A(n14593), .ZN(n4054) );
  NAND2_X1 U11313 ( .A1(n13783), .A2(n4055), .ZN(n4151) );
  NOR2_X1 U11314 ( .A1(n14593), .A2(n4056), .ZN(n4055) );
  INV_X1 U11315 ( .A(n14105), .ZN(n4056) );
  NAND2_X1 U11316 ( .A1(n14594), .A2(n14593), .ZN(n14258) );
  NAND3_X2 U11317 ( .A1(n4057), .A2(n10536), .A3(n10537), .ZN(n13563) );
  NAND2_X1 U11318 ( .A1(n10531), .A2(n12333), .ZN(n4057) );
  INV_X1 U11319 ( .A(n13563), .ZN(n13178) );
  NAND2_X1 U11320 ( .A1(n464), .A2(n24507), .ZN(n4063) );
  INV_X1 U11321 ( .A(n24269), .ZN(n24789) );
  NAND2_X1 U11322 ( .A1(n1955), .A2(n4065), .ZN(n4064) );
  NAND2_X1 U11323 ( .A1(n4576), .A2(n4066), .ZN(n4065) );
  NAND2_X1 U11324 ( .A1(n23655), .A2(n24269), .ZN(n4066) );
  NAND2_X1 U11325 ( .A1(n1854), .A2(n4067), .ZN(n4068) );
  MUX2_X1 U11326 ( .A(n11282), .B(n10884), .S(n11281), .Z(n4067) );
  XNOR2_X2 U11327 ( .A(n10369), .B(n10370), .ZN(n10884) );
  XNOR2_X1 U11330 ( .A(n19681), .B(n4069), .ZN(n19432) );
  XNOR2_X1 U11331 ( .A(n18653), .B(n4070), .ZN(n4069) );
  NAND3_X1 U11332 ( .A1(n4071), .A2(n21040), .A3(n21748), .ZN(n5976) );
  AND2_X1 U11333 ( .A1(n15342), .A2(n15224), .ZN(n14757) );
  NAND3_X1 U11335 ( .A1(n26131), .A2(n4079), .A3(n4078), .ZN(n27724) );
  NAND3_X1 U11336 ( .A1(n27129), .A2(n28536), .A3(n27177), .ZN(n4078) );
  NAND2_X1 U11337 ( .A1(n27173), .A2(n4080), .ZN(n4079) );
  OAI21_X2 U11338 ( .B1(n23307), .B2(n23306), .A(n4081), .ZN(n25884) );
  XNOR2_X1 U11339 ( .A(n25347), .B(n4083), .ZN(n4082) );
  XNOR2_X1 U11340 ( .A(n25346), .B(n25345), .ZN(n4083) );
  XNOR2_X1 U11341 ( .A(n25348), .B(n25713), .ZN(n4084) );
  XNOR2_X2 U11342 ( .A(n16118), .B(n16117), .ZN(n17259) );
  AOI21_X1 U11344 ( .B1(n4086), .B2(n23531), .A(n28164), .ZN(n4124) );
  OAI21_X1 U11345 ( .B1(n484), .B2(n23067), .A(n4086), .ZN(n5402) );
  NAND2_X1 U11346 ( .A1(n28164), .A2(n4086), .ZN(n6903) );
  OAI22_X1 U11347 ( .A1(n5029), .A2(n4086), .B1(n23135), .B2(n23535), .ZN(
        n5031) );
  NAND2_X1 U11348 ( .A1(n10627), .A2(n11014), .ZN(n4087) );
  INV_X1 U11349 ( .A(n13824), .ZN(n4088) );
  XNOR2_X2 U11350 ( .A(n13053), .B(n13052), .ZN(n13060) );
  NAND2_X1 U11351 ( .A1(n29373), .A2(n17491), .ZN(n17063) );
  NAND2_X1 U11353 ( .A1(n17063), .A2(n16882), .ZN(n4089) );
  NAND2_X1 U11354 ( .A1(n4092), .A2(n4091), .ZN(n4090) );
  NAND3_X1 U11355 ( .A1(n27382), .A2(n28394), .A3(n27213), .ZN(n4092) );
  NAND2_X1 U11356 ( .A1(n4093), .A2(n21304), .ZN(n6733) );
  NAND2_X1 U11357 ( .A1(n21150), .A2(n4094), .ZN(n4093) );
  NAND2_X1 U11358 ( .A1(n21311), .A2(n20938), .ZN(n4094) );
  NAND2_X1 U11359 ( .A1(n11292), .A2(n11291), .ZN(n4095) );
  MUX2_X1 U11360 ( .A(n11795), .B(n12081), .S(n29498), .Z(n11799) );
  NAND2_X1 U11362 ( .A1(n17219), .A2(n17555), .ZN(n4100) );
  NAND3_X1 U11364 ( .A1(n4982), .A2(n12131), .A3(n4981), .ZN(n4102) );
  INV_X1 U11365 ( .A(n21493), .ZN(n4104) );
  OAI21_X1 U11366 ( .B1(n21183), .B2(n21495), .A(n4104), .ZN(n4103) );
  NAND3_X1 U11367 ( .A1(n21186), .A2(n6503), .A3(n4103), .ZN(n6504) );
  NAND2_X1 U11368 ( .A1(n4105), .A2(n12280), .ZN(n11359) );
  OR2_X1 U11369 ( .A1(n12408), .A2(n4106), .ZN(n11627) );
  NAND2_X1 U11370 ( .A1(n12281), .A2(n12402), .ZN(n4106) );
  NAND3_X1 U11371 ( .A1(n4105), .A2(n12400), .A3(n11801), .ZN(n11626) );
  NAND3_X1 U11372 ( .A1(n4105), .A2(n12400), .A3(n12407), .ZN(n12067) );
  OAI21_X1 U11373 ( .B1(n12286), .B2(n4105), .A(n12400), .ZN(n12405) );
  NOR2_X1 U11374 ( .A1(n11333), .A2(n4107), .ZN(n4461) );
  NAND2_X1 U11375 ( .A1(n10466), .A2(n4107), .ZN(n10469) );
  NAND3_X1 U11378 ( .A1(n27193), .A2(n4243), .A3(n4109), .ZN(n4108) );
  NAND2_X1 U11379 ( .A1(n8155), .A2(n8154), .ZN(n4111) );
  NAND2_X1 U11380 ( .A1(n2056), .A2(n17393), .ZN(n4113) );
  NAND2_X1 U11381 ( .A1(n4116), .A2(n4115), .ZN(n4114) );
  NAND3_X1 U11382 ( .A1(n4117), .A2(n12201), .A3(n12202), .ZN(n4115) );
  NAND2_X1 U11383 ( .A1(n11602), .A2(n5825), .ZN(n4116) );
  NAND2_X1 U11384 ( .A1(n1966), .A2(n2063), .ZN(n4117) );
  INV_X1 U11385 ( .A(n12202), .ZN(n6020) );
  NAND3_X1 U11386 ( .A1(n17986), .A2(n17985), .A3(n18268), .ZN(n4120) );
  MUX2_X1 U11387 ( .A(n13842), .B(n14010), .S(n14131), .Z(n4122) );
  NAND2_X1 U11389 ( .A1(n11348), .A2(n11192), .ZN(n4123) );
  AOI21_X1 U11390 ( .B1(n4123), .B2(n9219), .A(n9218), .ZN(n9257) );
  XNOR2_X2 U11391 ( .A(n19737), .B(n19738), .ZN(n23535) );
  INV_X1 U11392 ( .A(n10547), .ZN(n4126) );
  NAND3_X1 U11393 ( .A1(n11111), .A2(n242), .A3(n10492), .ZN(n4127) );
  NAND2_X1 U11394 ( .A1(n4056), .A2(n14107), .ZN(n13608) );
  NAND2_X1 U11395 ( .A1(n14230), .A2(n4056), .ZN(n14103) );
  MUX2_X1 U11396 ( .A(n14107), .B(n4056), .S(n14231), .Z(n11371) );
  NAND3_X1 U11397 ( .A1(n4150), .A2(n14231), .A3(n4056), .ZN(n4149) );
  NAND3_X1 U11398 ( .A1(n4129), .A2(n7728), .A3(n7727), .ZN(n7731) );
  NAND2_X1 U11399 ( .A1(n27033), .A2(n27032), .ZN(n4130) );
  NAND2_X1 U11400 ( .A1(n27030), .A2(n4133), .ZN(n4132) );
  INV_X1 U11401 ( .A(n28592), .ZN(n4133) );
  NAND2_X1 U11402 ( .A1(n24713), .A2(n24716), .ZN(n4135) );
  NAND2_X1 U11403 ( .A1(n23060), .A2(n23344), .ZN(n4137) );
  NAND2_X1 U11404 ( .A1(n23059), .A2(n29108), .ZN(n4138) );
  INV_X1 U11405 ( .A(n13552), .ZN(n4139) );
  XNOR2_X1 U11406 ( .A(n4139), .B(n12566), .ZN(n11684) );
  NAND3_X2 U11408 ( .A1(n21228), .A2(n4142), .A3(n2022), .ZN(n6141) );
  INV_X1 U11409 ( .A(n21639), .ZN(n4143) );
  NAND3_X1 U11410 ( .A1(n28797), .A2(n4143), .A3(n21638), .ZN(n4142) );
  INV_X1 U11411 ( .A(n12017), .ZN(n12016) );
  NAND2_X1 U11412 ( .A1(n11747), .A2(n12328), .ZN(n12017) );
  OAI211_X1 U11413 ( .C1(n10523), .C2(n11038), .A(n28612), .B(n11275), .ZN(
        n4145) );
  NAND2_X1 U11414 ( .A1(n10525), .A2(n29148), .ZN(n4146) );
  INV_X1 U11415 ( .A(n4148), .ZN(n21613) );
  OR2_X2 U11416 ( .A1(n20492), .A2(n21329), .ZN(n4148) );
  NAND2_X1 U11417 ( .A1(n4148), .A2(n21327), .ZN(n21618) );
  AND2_X1 U11418 ( .A1(n28791), .A2(n21613), .ZN(n20910) );
  NAND2_X1 U11419 ( .A1(n4148), .A2(n21326), .ZN(n20906) );
  NAND2_X1 U11420 ( .A1(n4147), .A2(n21163), .ZN(n20732) );
  AND2_X1 U11421 ( .A1(n28791), .A2(n4148), .ZN(n4147) );
  NAND3_X1 U11422 ( .A1(n4151), .A2(n4149), .A3(n13784), .ZN(n14928) );
  INV_X1 U11423 ( .A(n14107), .ZN(n13783) );
  INV_X1 U11424 ( .A(n4152), .ZN(n4153) );
  INV_X1 U11425 ( .A(n17771), .ZN(n17583) );
  NAND3_X1 U11427 ( .A1(n4157), .A2(n4158), .A3(n4156), .ZN(n4154) );
  MUX2_X1 U11428 ( .A(n17575), .B(n17574), .S(n17707), .Z(n4155) );
  NAND2_X1 U11429 ( .A1(n17707), .A2(n17570), .ZN(n4158) );
  XNOR2_X1 U11430 ( .A(n4161), .B(n25454), .ZN(n24948) );
  XNOR2_X1 U11431 ( .A(n4161), .B(n25855), .ZN(n25857) );
  XNOR2_X1 U11432 ( .A(n4161), .B(n4384), .ZN(n25479) );
  XNOR2_X1 U11433 ( .A(n25944), .B(n4161), .ZN(n25094) );
  OAI21_X1 U11435 ( .B1(n15055), .B2(n15054), .A(n4162), .ZN(n14764) );
  NAND2_X1 U11438 ( .A1(n27508), .A2(n29556), .ZN(n4165) );
  NAND2_X1 U11439 ( .A1(n4166), .A2(n14278), .ZN(n14274) );
  NAND2_X1 U11440 ( .A1(n14362), .A2(n4166), .ZN(n4667) );
  NAND2_X1 U11442 ( .A1(n6188), .A2(n9037), .ZN(n6190) );
  NAND3_X1 U11443 ( .A1(n424), .A2(n16878), .A3(n29045), .ZN(n4168) );
  NAND3_X1 U11444 ( .A1(n15072), .A2(n15071), .A3(n14571), .ZN(n4169) );
  NAND2_X1 U11445 ( .A1(n4172), .A2(n20125), .ZN(n18546) );
  OAI21_X1 U11446 ( .B1(n20294), .B2(n20293), .A(n4172), .ZN(n20296) );
  NAND2_X1 U11447 ( .A1(n20293), .A2(n19815), .ZN(n4172) );
  AOI21_X1 U11448 ( .B1(n26230), .B2(n26740), .A(n26229), .ZN(n26231) );
  NAND2_X1 U11449 ( .A1(n25598), .A2(n26740), .ZN(n25600) );
  NAND2_X1 U11450 ( .A1(n25349), .A2(n26740), .ZN(n4173) );
  NAND2_X1 U11451 ( .A1(n4174), .A2(n18198), .ZN(n16719) );
  NOR2_X1 U11452 ( .A1(n4174), .A2(n18449), .ZN(n6326) );
  INV_X1 U11453 ( .A(n23302), .ZN(n4178) );
  NAND2_X1 U11455 ( .A1(n7496), .A2(n7250), .ZN(n7254) );
  NAND2_X1 U11456 ( .A1(n7494), .A2(n7250), .ZN(n7251) );
  OAI21_X1 U11457 ( .B1(n7250), .B2(n7498), .A(n7496), .ZN(n4180) );
  NAND2_X1 U11458 ( .A1(n7705), .A2(n7250), .ZN(n7497) );
  NAND2_X1 U11460 ( .A1(n4186), .A2(n14841), .ZN(n4185) );
  NAND2_X1 U11461 ( .A1(n6048), .A2(n14842), .ZN(n4186) );
  NAND2_X1 U11463 ( .A1(n4188), .A2(n16805), .ZN(n16807) );
  INV_X1 U11464 ( .A(n17260), .ZN(n4188) );
  NAND2_X1 U11465 ( .A1(n6408), .A2(n414), .ZN(n4189) );
  NAND2_X1 U11466 ( .A1(n20040), .A2(n20039), .ZN(n4190) );
  NAND2_X1 U11467 ( .A1(n17958), .A2(n6914), .ZN(n4192) );
  OAI211_X2 U11468 ( .C1(n17473), .C2(n17472), .A(n17471), .B(n17515), .ZN(
        n18216) );
  NAND2_X1 U11469 ( .A1(n21567), .A2(n4193), .ZN(n21462) );
  NOR2_X1 U11470 ( .A1(n4193), .A2(n21567), .ZN(n21572) );
  AND2_X1 U11471 ( .A1(n4494), .A2(n4193), .ZN(n21568) );
  NAND2_X1 U11472 ( .A1(n5176), .A2(n4193), .ZN(n5175) );
  OAI21_X1 U11473 ( .B1(n24075), .B2(n4195), .A(n4194), .ZN(n24670) );
  INV_X1 U11475 ( .A(n12305), .ZN(n12299) );
  OAI21_X2 U11476 ( .B1(n6774), .B2(n10959), .A(n6773), .ZN(n12305) );
  NAND2_X1 U11479 ( .A1(n21183), .A2(n21497), .ZN(n4201) );
  NAND2_X1 U11480 ( .A1(n20751), .A2(n7), .ZN(n4202) );
  NAND2_X1 U11481 ( .A1(n20752), .A2(n4104), .ZN(n4206) );
  XNOR2_X2 U11482 ( .A(n13424), .B(n13423), .ZN(n13725) );
  NAND3_X1 U11483 ( .A1(n14372), .A2(n5404), .A3(n14373), .ZN(n6614) );
  INV_X1 U11484 ( .A(n17694), .ZN(n4209) );
  NAND2_X1 U11485 ( .A1(n17692), .A2(n18509), .ZN(n4210) );
  INV_X1 U11486 ( .A(n18512), .ZN(n4211) );
  NAND2_X1 U11487 ( .A1(n17691), .A2(n18512), .ZN(n4212) );
  NOR2_X1 U11488 ( .A1(n4213), .A2(n18333), .ZN(n4214) );
  XNOR2_X1 U11489 ( .A(n4216), .B(n1998), .ZN(n4215) );
  XNOR2_X1 U11490 ( .A(n15612), .B(n1967), .ZN(n4216) );
  OR2_X1 U11491 ( .A1(n17549), .A2(n4218), .ZN(n17241) );
  NOR2_X1 U11492 ( .A1(n17239), .A2(n4218), .ZN(n15685) );
  NAND3_X1 U11493 ( .A1(n2122), .A2(n17548), .A3(n4218), .ZN(n17550) );
  AOI21_X1 U11494 ( .B1(n5398), .B2(n4218), .A(n16762), .ZN(n17240) );
  OR2_X2 U11495 ( .A1(n12097), .A2(n10784), .ZN(n12151) );
  NAND4_X2 U11496 ( .A1(n6149), .A2(n4219), .A3(n26437), .A4(n6148), .ZN(
        n27301) );
  NAND3_X1 U11497 ( .A1(n456), .A2(n26944), .A3(n26768), .ZN(n4219) );
  XNOR2_X1 U11501 ( .A(n4221), .B(n19702), .ZN(n19454) );
  NAND2_X1 U11502 ( .A1(n21561), .A2(n21113), .ZN(n4223) );
  NAND2_X1 U11503 ( .A1(n6861), .A2(n1897), .ZN(n4225) );
  MUX2_X1 U11504 ( .A(n4227), .B(n26336), .S(n27123), .Z(n26337) );
  INV_X1 U11505 ( .A(n27191), .ZN(n4227) );
  NAND2_X1 U11507 ( .A1(n18107), .A2(n18106), .ZN(n4230) );
  NAND2_X1 U11508 ( .A1(n18789), .A2(n29114), .ZN(n6400) );
  INV_X1 U11511 ( .A(n19985), .ZN(n20164) );
  NOR2_X1 U11512 ( .A1(n24631), .A2(n24630), .ZN(n24294) );
  NAND2_X1 U11513 ( .A1(n27038), .A2(n5581), .ZN(n4236) );
  NOR2_X1 U11515 ( .A1(n5314), .A2(n27213), .ZN(n27380) );
  NAND2_X1 U11518 ( .A1(n24632), .A2(n6867), .ZN(n4239) );
  INV_X1 U11519 ( .A(n21388), .ZN(n4242) );
  INV_X1 U11520 ( .A(n27124), .ZN(n4243) );
  NAND2_X1 U11521 ( .A1(n20449), .A2(n4245), .ZN(n19573) );
  NAND2_X1 U11522 ( .A1(n5377), .A2(n4245), .ZN(n19899) );
  NOR2_X1 U11523 ( .A1(n19927), .A2(n4245), .ZN(n19930) );
  OAI21_X1 U11524 ( .B1(n6203), .B2(n4245), .A(n20451), .ZN(n5375) );
  XNOR2_X2 U11525 ( .A(n16175), .B(n16174), .ZN(n4246) );
  NAND2_X1 U11526 ( .A1(n4246), .A2(n17464), .ZN(n16675) );
  NOR2_X1 U11527 ( .A1(n17467), .A2(n4246), .ZN(n16819) );
  NAND2_X1 U11528 ( .A1(n17467), .A2(n4246), .ZN(n17093) );
  OAI21_X1 U11529 ( .B1(n29022), .B2(n29118), .A(n4247), .ZN(n6490) );
  NAND2_X1 U11530 ( .A1(n29022), .A2(n27772), .ZN(n4247) );
  NAND2_X1 U11531 ( .A1(n4247), .A2(n4248), .ZN(n27776) );
  NAND2_X1 U11533 ( .A1(n27784), .A2(n4250), .ZN(n27770) );
  NAND2_X1 U11534 ( .A1(n14033), .A2(n14030), .ZN(n13794) );
  NAND3_X1 U11535 ( .A1(n14033), .A2(n14030), .A3(n14029), .ZN(n4252) );
  XNOR2_X1 U11536 ( .A(n4253), .B(n12931), .ZN(n13457) );
  XNOR2_X1 U11537 ( .A(n4253), .B(n2894), .ZN(n11389) );
  XNOR2_X1 U11538 ( .A(n4253), .B(n6683), .ZN(n12705) );
  XNOR2_X1 U11539 ( .A(n4253), .B(n12960), .ZN(n12962) );
  XNOR2_X1 U11540 ( .A(n13222), .B(n4253), .ZN(n13223) );
  NAND2_X1 U11541 ( .A1(n21118), .A2(n29581), .ZN(n20650) );
  MUX2_X1 U11542 ( .A(n21145), .B(n21118), .S(n21144), .Z(n19784) );
  NOR2_X1 U11543 ( .A1(n13572), .A2(n14380), .ZN(n4258) );
  NAND2_X1 U11544 ( .A1(n556), .A2(n14004), .ZN(n14379) );
  XNOR2_X2 U11545 ( .A(n13560), .B(n13561), .ZN(n14004) );
  NAND2_X1 U11546 ( .A1(n8642), .A2(n8984), .ZN(n8456) );
  NAND3_X1 U11547 ( .A1(n8642), .A2(n8984), .A3(n8981), .ZN(n8987) );
  NAND2_X1 U11548 ( .A1(n13729), .A2(n13914), .ZN(n4260) );
  XNOR2_X1 U11549 ( .A(n4263), .B(n25515), .ZN(n24923) );
  XNOR2_X1 U11550 ( .A(n4263), .B(n26108), .ZN(n25877) );
  NAND2_X1 U11551 ( .A1(n11677), .A2(n11515), .ZN(n11517) );
  AOI21_X1 U11552 ( .B1(n10746), .B2(n10819), .A(n28208), .ZN(n11633) );
  NAND3_X1 U11553 ( .A1(n10976), .A2(n4264), .A3(n28608), .ZN(n6896) );
  INV_X1 U11554 ( .A(n10972), .ZN(n4264) );
  INV_X1 U11555 ( .A(n19732), .ZN(n4266) );
  OAI21_X1 U11556 ( .B1(n21379), .B2(n21810), .A(n4266), .ZN(n21381) );
  NAND2_X1 U11557 ( .A1(n4270), .A2(n17484), .ZN(n4269) );
  AOI21_X1 U11558 ( .B1(n17831), .B2(n17830), .A(n4272), .ZN(n17832) );
  NAND3_X1 U11562 ( .A1(n11146), .A2(n28206), .A3(n10544), .ZN(n4275) );
  NAND2_X1 U11563 ( .A1(n12071), .A2(n12070), .ZN(n4276) );
  NAND2_X1 U11564 ( .A1(n19808), .A2(n20137), .ZN(n4278) );
  OAI21_X1 U11565 ( .B1(n4283), .B2(n16953), .A(n4279), .ZN(n4282) );
  NAND2_X1 U11567 ( .A1(n4282), .A2(n28793), .ZN(n4280) );
  NAND2_X1 U11568 ( .A1(n18539), .A2(n18260), .ZN(n16955) );
  NAND2_X1 U11569 ( .A1(n16952), .A2(n17354), .ZN(n4281) );
  INV_X1 U11570 ( .A(n14376), .ZN(n13594) );
  NAND2_X1 U11571 ( .A1(n14533), .A2(n15190), .ZN(n14531) );
  NAND2_X1 U11572 ( .A1(n13814), .A2(n4284), .ZN(n14784) );
  NAND3_X1 U11573 ( .A1(n29737), .A2(n387), .A3(n17467), .ZN(n4285) );
  XNOR2_X1 U11574 ( .A(n6080), .B(n16414), .ZN(n16454) );
  NAND2_X1 U11575 ( .A1(n14577), .A2(n14936), .ZN(n4287) );
  NAND2_X1 U11576 ( .A1(n14576), .A2(n549), .ZN(n4288) );
  AND2_X1 U11577 ( .A1(n28806), .A2(n14460), .ZN(n14458) );
  MUX2_X1 U11578 ( .A(n4290), .B(n14204), .S(n28806), .Z(n13864) );
  INV_X1 U11580 ( .A(n12712), .ZN(n4290) );
  NAND2_X1 U11581 ( .A1(n380), .A2(n23712), .ZN(n6153) );
  NAND2_X2 U11582 ( .A1(n4291), .A2(n4293), .ZN(n18382) );
  OAI21_X1 U11584 ( .B1(n18351), .B2(n18383), .A(n18350), .ZN(n5920) );
  NAND2_X1 U11585 ( .A1(n4295), .A2(n16712), .ZN(n4294) );
  INV_X1 U11586 ( .A(n11317), .ZN(n4815) );
  NAND2_X1 U11587 ( .A1(n4296), .A2(n11253), .ZN(n11317) );
  XNOR2_X1 U11588 ( .A(n4298), .B(n13433), .ZN(n13362) );
  XNOR2_X1 U11589 ( .A(n12064), .B(n4297), .ZN(n12972) );
  XNOR2_X1 U11590 ( .A(n12808), .B(n4298), .ZN(n11563) );
  NAND2_X1 U11591 ( .A1(n23261), .A2(n23712), .ZN(n23235) );
  OAI21_X2 U11592 ( .B1(n4299), .B2(n14994), .A(n14993), .ZN(n16444) );
  NAND2_X1 U11594 ( .A1(n4303), .A2(n9202), .ZN(n4302) );
  NAND2_X1 U11596 ( .A1(n8994), .A2(n4305), .ZN(n4304) );
  INV_X1 U11597 ( .A(n8995), .ZN(n4305) );
  NAND2_X1 U11598 ( .A1(n3900), .A2(n11553), .ZN(n6742) );
  NAND2_X1 U11599 ( .A1(n20458), .A2(n4306), .ZN(n20459) );
  NOR2_X1 U11600 ( .A1(n20458), .A2(n4306), .ZN(n20027) );
  INV_X1 U11603 ( .A(n22401), .ZN(n22398) );
  OR2_X2 U11604 ( .A1(n20264), .A2(n20263), .ZN(n22401) );
  NAND2_X1 U11605 ( .A1(n4310), .A2(n4308), .ZN(n4311) );
  NAND2_X1 U11606 ( .A1(n5151), .A2(n22401), .ZN(n4309) );
  NAND2_X1 U11607 ( .A1(n22396), .A2(n22398), .ZN(n4310) );
  NAND2_X1 U11608 ( .A1(n17064), .A2(n538), .ZN(n4315) );
  NAND2_X1 U11609 ( .A1(n4315), .A2(n4313), .ZN(n17206) );
  AOI21_X1 U11610 ( .B1(n2549), .B2(n4509), .A(n14402), .ZN(n13965) );
  NAND2_X1 U11611 ( .A1(n17566), .A2(n4316), .ZN(n17227) );
  NAND2_X1 U11612 ( .A1(n17568), .A2(n4316), .ZN(n6306) );
  XNOR2_X1 U11613 ( .A(n9823), .B(n9824), .ZN(n10229) );
  NAND2_X1 U11614 ( .A1(n4319), .A2(n28743), .ZN(n4318) );
  NAND2_X1 U11615 ( .A1(n4322), .A2(n8366), .ZN(n4319) );
  XNOR2_X1 U11616 ( .A(n4323), .B(n3378), .ZN(n14868) );
  XNOR2_X1 U11617 ( .A(n16606), .B(n4323), .ZN(n16609) );
  XNOR2_X1 U11618 ( .A(n3661), .B(n4323), .ZN(n16347) );
  XNOR2_X1 U11619 ( .A(n15780), .B(n4323), .ZN(n15649) );
  AOI22_X1 U11620 ( .A1(n4296), .A2(n11318), .B1(n11314), .B2(n4326), .ZN(
        n4325) );
  NAND2_X1 U11621 ( .A1(n4296), .A2(n11315), .ZN(n4327) );
  NAND2_X1 U11622 ( .A1(n4329), .A2(n11253), .ZN(n4328) );
  NAND2_X1 U11623 ( .A1(n29059), .A2(n14372), .ZN(n14374) );
  NAND2_X1 U11624 ( .A1(n16918), .A2(n29550), .ZN(n4332) );
  NAND2_X1 U11625 ( .A1(n4335), .A2(n24804), .ZN(n4333) );
  NAND2_X1 U11626 ( .A1(n24805), .A2(n24806), .ZN(n4334) );
  NAND2_X1 U11627 ( .A1(n23689), .A2(n1914), .ZN(n23803) );
  OR2_X1 U11629 ( .A1(n23800), .A2(n23801), .ZN(n4337) );
  OAI211_X1 U11630 ( .C1(n416), .C2(n4340), .A(n5436), .B(n4338), .ZN(n20890)
         );
  NAND2_X1 U11631 ( .A1(n4340), .A2(n20302), .ZN(n18117) );
  NAND2_X1 U11632 ( .A1(n20303), .A2(n4340), .ZN(n20204) );
  NAND2_X1 U11633 ( .A1(n4341), .A2(n11194), .ZN(n11956) );
  OAI21_X1 U11635 ( .B1(n21590), .B2(n28584), .A(n4342), .ZN(n4343) );
  NOR2_X1 U11636 ( .A1(n21586), .A2(n21585), .ZN(n4344) );
  NAND2_X1 U11638 ( .A1(n11843), .A2(n4346), .ZN(n4345) );
  NAND2_X1 U11639 ( .A1(n373), .A2(n17858), .ZN(n6230) );
  NAND2_X1 U11640 ( .A1(n12232), .A2(n776), .ZN(n11680) );
  NAND3_X1 U11641 ( .A1(n12232), .A2(n776), .A3(n12236), .ZN(n4349) );
  INV_X1 U11642 ( .A(n10662), .ZN(n4350) );
  INV_X1 U11643 ( .A(n10658), .ZN(n4351) );
  AND2_X2 U11644 ( .A1(n4353), .A2(n2078), .ZN(n27855) );
  NAND2_X1 U11645 ( .A1(n26990), .A2(n26321), .ZN(n4354) );
  NAND2_X1 U11646 ( .A1(n27079), .A2(n27074), .ZN(n4355) );
  OAI211_X1 U11647 ( .C1(n4358), .C2(n14840), .A(n4357), .B(n4356), .ZN(n4360)
         );
  NAND2_X1 U11648 ( .A1(n14840), .A2(n4359), .ZN(n4356) );
  NAND2_X1 U11649 ( .A1(n14839), .A2(n4359), .ZN(n4357) );
  INV_X1 U11650 ( .A(n15887), .ZN(n16436) );
  NOR2_X1 U11651 ( .A1(n21028), .A2(n21627), .ZN(n6530) );
  INV_X1 U11652 ( .A(n24629), .ZN(n24293) );
  NAND2_X1 U11653 ( .A1(n4365), .A2(n4363), .ZN(n6198) );
  NAND3_X1 U11654 ( .A1(n6867), .A2(n24891), .A3(n4364), .ZN(n4363) );
  INV_X1 U11655 ( .A(n4364), .ZN(n4366) );
  NAND2_X1 U11657 ( .A1(n4369), .A2(n14075), .ZN(n14830) );
  INV_X1 U11659 ( .A(n7199), .ZN(n4370) );
  NAND2_X1 U11660 ( .A1(n7406), .A2(n8280), .ZN(n7199) );
  OR2_X1 U11661 ( .A1(n17979), .A2(n18234), .ZN(n4372) );
  INV_X1 U11662 ( .A(n17979), .ZN(n4373) );
  NAND2_X1 U11663 ( .A1(n18233), .A2(n18398), .ZN(n17979) );
  OAI21_X1 U11664 ( .B1(n18400), .B2(n18398), .A(n18401), .ZN(n4374) );
  NAND3_X1 U11665 ( .A1(n4376), .A2(n13938), .A3(n14237), .ZN(n13940) );
  OR2_X1 U11666 ( .A1(n491), .A2(n4382), .ZN(n4377) );
  INV_X1 U11667 ( .A(n22000), .ZN(n22897) );
  OAI211_X2 U11668 ( .C1(n4380), .C2(n4379), .A(n4378), .B(n4377), .ZN(n22000)
         );
  NAND2_X1 U11669 ( .A1(n4381), .A2(n21823), .ZN(n4379) );
  NAND2_X1 U11670 ( .A1(n495), .A2(n21078), .ZN(n4381) );
  OR2_X1 U11671 ( .A1(n20933), .A2(n22013), .ZN(n4382) );
  AND2_X1 U11672 ( .A1(n10114), .A2(n11124), .ZN(n10505) );
  XNOR2_X1 U11673 ( .A(n4384), .B(n24060), .ZN(n24061) );
  XNOR2_X1 U11674 ( .A(n4384), .B(n3334), .ZN(n24873) );
  XNOR2_X1 U11675 ( .A(n4384), .B(n25947), .ZN(n25950) );
  XNOR2_X1 U11676 ( .A(n25149), .B(n4384), .ZN(n5432) );
  INV_X1 U11678 ( .A(n29102), .ZN(n4385) );
  AND2_X1 U11679 ( .A1(n20041), .A2(n29104), .ZN(n6408) );
  XNOR2_X1 U11680 ( .A(n13180), .B(n4387), .ZN(n12530) );
  INV_X1 U11681 ( .A(n13284), .ZN(n4387) );
  XNOR2_X1 U11682 ( .A(n4388), .B(n13449), .ZN(n13455) );
  INV_X1 U11683 ( .A(n13180), .ZN(n4388) );
  NAND2_X1 U11684 ( .A1(n28206), .A2(n10808), .ZN(n10740) );
  INV_X1 U11686 ( .A(n17125), .ZN(n4391) );
  NAND2_X1 U11687 ( .A1(n4392), .A2(n17627), .ZN(n6654) );
  NAND2_X1 U11688 ( .A1(n17626), .A2(n17636), .ZN(n4392) );
  NAND2_X1 U11689 ( .A1(n21146), .A2(n4394), .ZN(n4393) );
  NAND2_X1 U11690 ( .A1(n21144), .A2(n21145), .ZN(n4395) );
  OAI211_X1 U11692 ( .C1(n14341), .C2(n14131), .A(n14010), .B(n4396), .ZN(
        n4398) );
  NAND2_X1 U11693 ( .A1(n14136), .A2(n14131), .ZN(n4396) );
  AOI21_X1 U11694 ( .B1(n20049), .B2(n20067), .A(n6477), .ZN(n4403) );
  OAI21_X1 U11695 ( .B1(n4403), .B2(n20068), .A(n6476), .ZN(n20425) );
  AOI21_X1 U11696 ( .B1(n21076), .B2(n20933), .A(n21823), .ZN(n20428) );
  NAND2_X1 U11697 ( .A1(n12300), .A2(n12305), .ZN(n4404) );
  NAND3_X1 U11698 ( .A1(n11493), .A2(n12307), .A3(n11495), .ZN(n11768) );
  NAND2_X1 U11700 ( .A1(n10737), .A2(n10914), .ZN(n4405) );
  NAND3_X1 U11701 ( .A1(n18125), .A2(n18588), .A3(n18126), .ZN(n4406) );
  OAI21_X1 U11702 ( .B1(n18129), .B2(n18127), .A(n4406), .ZN(n18133) );
  OAI21_X1 U11703 ( .B1(n18593), .B2(n18592), .A(n4406), .ZN(n18594) );
  OAI21_X2 U11704 ( .B1(n6813), .B2(n13256), .A(n6812), .ZN(n15691) );
  INV_X1 U11706 ( .A(n29058), .ZN(n4411) );
  AOI21_X1 U11707 ( .B1(n28783), .B2(n4411), .A(n29570), .ZN(n4486) );
  NAND2_X1 U11708 ( .A1(n2007), .A2(n28448), .ZN(n6476) );
  INV_X1 U11709 ( .A(n20064), .ZN(n18765) );
  INV_X1 U11710 ( .A(n17505), .ZN(n17073) );
  INV_X1 U11711 ( .A(n17484), .ZN(n17074) );
  NAND2_X1 U11712 ( .A1(n17073), .A2(n17830), .ZN(n4413) );
  NAND2_X1 U11713 ( .A1(n4415), .A2(n407), .ZN(n23439) );
  NAND2_X1 U11714 ( .A1(n4418), .A2(n6207), .ZN(n4417) );
  INV_X1 U11715 ( .A(n15260), .ZN(n15055) );
  NAND2_X1 U11717 ( .A1(n17891), .A2(n18600), .ZN(n4420) );
  NAND2_X1 U11718 ( .A1(n13581), .A2(n13900), .ZN(n4422) );
  INV_X1 U11719 ( .A(n14144), .ZN(n4423) );
  AOI21_X1 U11720 ( .B1(n4423), .B2(n4425), .A(n2974), .ZN(n4424) );
  NAND2_X1 U11721 ( .A1(n389), .A2(n13902), .ZN(n4426) );
  NAND2_X1 U11722 ( .A1(n12202), .A2(n12203), .ZN(n11438) );
  XNOR2_X2 U11725 ( .A(n12838), .B(n12837), .ZN(n14192) );
  NAND2_X1 U11727 ( .A1(n8326), .A2(n9425), .ZN(n5132) );
  NAND2_X1 U11730 ( .A1(n7310), .A2(n7092), .ZN(n4439) );
  NAND3_X1 U11732 ( .A1(n4442), .A2(n4441), .A3(n7419), .ZN(n4440) );
  NAND2_X1 U11733 ( .A1(n8609), .A2(n8751), .ZN(n4441) );
  OAI21_X1 U11734 ( .B1(n29395), .B2(n9532), .A(n9531), .ZN(n4442) );
  XNOR2_X1 U11735 ( .A(n12787), .B(n12788), .ZN(n12949) );
  NAND2_X1 U11737 ( .A1(n4449), .A2(n4037), .ZN(n4447) );
  NAND2_X1 U11738 ( .A1(n12211), .A2(n12110), .ZN(n4448) );
  NAND2_X1 U11739 ( .A1(n24078), .A2(n24081), .ZN(n5272) );
  OR2_X2 U11740 ( .A1(n6277), .A2(n6278), .ZN(n24078) );
  INV_X1 U11741 ( .A(n4450), .ZN(n5857) );
  NOR2_X1 U11742 ( .A1(n18504), .A2(n4450), .ZN(n18505) );
  NAND3_X1 U11743 ( .A1(n4685), .A2(n24809), .A3(n24808), .ZN(n24500) );
  NOR2_X1 U11744 ( .A1(n29500), .A2(n27069), .ZN(n25720) );
  NAND2_X1 U11745 ( .A1(n27063), .A2(n27069), .ZN(n26616) );
  AOI21_X1 U11746 ( .B1(n14288), .B2(n4451), .A(n14287), .ZN(n14289) );
  XNOR2_X1 U11747 ( .A(n15973), .B(n15972), .ZN(n4452) );
  XNOR2_X1 U11748 ( .A(n15975), .B(n16198), .ZN(n4453) );
  XNOR2_X1 U11750 ( .A(n16294), .B(n3457), .ZN(n15558) );
  NAND4_X2 U11751 ( .A1(n14651), .A2(n4458), .A3(n4457), .A4(n4456), .ZN(
        n16294) );
  NAND2_X1 U11752 ( .A1(n14650), .A2(n6879), .ZN(n4456) );
  NAND2_X1 U11753 ( .A1(n15373), .A2(n14863), .ZN(n4457) );
  NAND2_X1 U11754 ( .A1(n4459), .A2(n23529), .ZN(n6442) );
  NAND2_X1 U11755 ( .A1(n21004), .A2(n4460), .ZN(n20213) );
  NOR2_X1 U11756 ( .A1(n23545), .A2(n4231), .ZN(n4847) );
  NAND2_X1 U11757 ( .A1(n5773), .A2(n23351), .ZN(n23545) );
  AOI21_X1 U11758 ( .B1(n20847), .B2(n4464), .A(n5142), .ZN(n4465) );
  NAND2_X1 U11759 ( .A1(n21576), .A2(n21577), .ZN(n4464) );
  NOR2_X1 U11760 ( .A1(n21487), .A2(n21580), .ZN(n4467) );
  XNOR2_X1 U11762 ( .A(n4468), .B(n27850), .ZN(Ciphertext[139]) );
  OAI211_X1 U11763 ( .C1(n27848), .C2(n27849), .A(n4470), .B(n4469), .ZN(n4468) );
  NAND2_X1 U11764 ( .A1(n27847), .A2(n2010), .ZN(n4469) );
  NAND2_X1 U11765 ( .A1(n27852), .A2(n27859), .ZN(n4470) );
  NOR2_X1 U11769 ( .A1(n28183), .A2(n23726), .ZN(n23848) );
  XNOR2_X1 U11770 ( .A(n4474), .B(n12608), .ZN(n13510) );
  INV_X1 U11771 ( .A(n13510), .ZN(n13038) );
  NAND2_X1 U11772 ( .A1(n16759), .A2(n17232), .ZN(n4476) );
  NAND2_X1 U11773 ( .A1(n16760), .A2(n4478), .ZN(n4477) );
  XNOR2_X1 U11774 ( .A(n4479), .B(n3385), .ZN(n9955) );
  XNOR2_X1 U11775 ( .A(n4479), .B(n10356), .ZN(n10015) );
  XNOR2_X1 U11776 ( .A(n4479), .B(n10208), .ZN(n9631) );
  NAND3_X1 U11777 ( .A1(n28497), .A2(n17389), .A3(n16879), .ZN(n4480) );
  XNOR2_X1 U11778 ( .A(n4482), .B(n29548), .ZN(n22581) );
  XNOR2_X1 U11779 ( .A(n22407), .B(n22668), .ZN(n4482) );
  NAND2_X1 U11780 ( .A1(n24489), .A2(n24471), .ZN(n24493) );
  NAND2_X1 U11781 ( .A1(n23848), .A2(n23849), .ZN(n24093) );
  OAI211_X1 U11782 ( .C1(n28183), .C2(n23849), .A(n23846), .B(n23843), .ZN(
        n4484) );
  NAND2_X1 U11784 ( .A1(n4487), .A2(n4486), .ZN(n4485) );
  OAI21_X1 U11785 ( .B1(n1530), .B2(n18042), .A(n17802), .ZN(n16866) );
  XNOR2_X1 U11786 ( .A(n4489), .B(n12833), .ZN(n12838) );
  INV_X1 U11787 ( .A(n12834), .ZN(n4489) );
  INV_X1 U11788 ( .A(n12833), .ZN(n4490) );
  NAND3_X1 U11789 ( .A1(n15024), .A2(n15023), .A3(n4491), .ZN(n4493) );
  XNOR2_X1 U11790 ( .A(n15862), .B(n4492), .ZN(n5798) );
  XNOR2_X1 U11791 ( .A(n15862), .B(n630), .ZN(n16505) );
  INV_X1 U11792 ( .A(n21457), .ZN(n4494) );
  NOR2_X2 U11793 ( .A1(n4495), .A2(n4498), .ZN(n27996) );
  NAND2_X1 U11794 ( .A1(n26633), .A2(n29058), .ZN(n4496) );
  MUX2_X1 U11795 ( .A(n27997), .B(n27977), .S(n27996), .Z(n26636) );
  MUX2_X1 U11796 ( .A(n27045), .B(n28130), .S(n29058), .Z(n4499) );
  XNOR2_X1 U11798 ( .A(n13273), .B(n4502), .ZN(n12499) );
  XNOR2_X1 U11799 ( .A(n13273), .B(n4503), .ZN(n12384) );
  INV_X1 U11800 ( .A(n1248), .ZN(n4503) );
  XNOR2_X1 U11801 ( .A(n10143), .B(n301), .ZN(n4508) );
  XNOR2_X1 U11802 ( .A(n10147), .B(n10148), .ZN(n4506) );
  MUX2_X1 U11803 ( .A(n28804), .B(n14400), .S(n13877), .Z(n14213) );
  NAND2_X1 U11804 ( .A1(n13707), .A2(n4509), .ZN(n13709) );
  OAI21_X1 U11805 ( .B1(n4801), .B2(n29148), .A(n4511), .ZN(n10480) );
  NAND2_X1 U11806 ( .A1(n3820), .A2(n29149), .ZN(n4511) );
  OAI211_X1 U11807 ( .C1(n15462), .C2(n4515), .A(n4513), .B(n15160), .ZN(n4512) );
  NAND2_X1 U11808 ( .A1(n15462), .A2(n15463), .ZN(n4514) );
  NAND2_X1 U11809 ( .A1(n4517), .A2(n17696), .ZN(n4516) );
  MUX2_X1 U11810 ( .A(n17695), .B(n18275), .S(n18203), .Z(n4517) );
  NAND3_X1 U11812 ( .A1(n14705), .A2(n15265), .A3(n15506), .ZN(n6217) );
  NAND2_X1 U11813 ( .A1(n29558), .A2(n4520), .ZN(n4519) );
  NOR2_X1 U11814 ( .A1(n28199), .A2(n14426), .ZN(n4520) );
  NAND2_X1 U11815 ( .A1(n4523), .A2(n4522), .ZN(n4521) );
  INV_X1 U11816 ( .A(n13874), .ZN(n4522) );
  OAI211_X1 U11817 ( .C1(n4526), .C2(n27224), .A(n4525), .B(n4524), .ZN(
        Ciphertext[54]) );
  NAND2_X1 U11818 ( .A1(n27224), .A2(n4527), .ZN(n4524) );
  OAI21_X1 U11819 ( .B1(n27223), .B2(n4528), .A(n4527), .ZN(n4525) );
  INV_X1 U11821 ( .A(n27225), .ZN(n4527) );
  AOI21_X1 U11822 ( .B1(n27222), .B2(n27221), .A(n27520), .ZN(n4528) );
  NAND2_X1 U11823 ( .A1(n27525), .A2(n6095), .ZN(n27221) );
  XNOR2_X1 U11824 ( .A(n5621), .B(n4529), .ZN(n4531) );
  XNOR2_X1 U11825 ( .A(n16005), .B(n4530), .ZN(n4529) );
  INV_X1 U11826 ( .A(n16649), .ZN(n4530) );
  NAND2_X1 U11827 ( .A1(n24094), .A2(n24470), .ZN(n24096) );
  NAND2_X1 U11828 ( .A1(n4536), .A2(n27854), .ZN(n4533) );
  XNOR2_X1 U11829 ( .A(n4535), .B(n2116), .ZN(Ciphertext[143]) );
  NAND2_X1 U11830 ( .A1(n10785), .A2(n10993), .ZN(n10691) );
  NOR2_X1 U11831 ( .A1(n3454), .A2(n10991), .ZN(n4539) );
  XNOR2_X2 U11832 ( .A(n9798), .B(n9793), .ZN(n10993) );
  NAND2_X1 U11833 ( .A1(n9179), .A2(n6828), .ZN(n4540) );
  NAND2_X1 U11834 ( .A1(n9178), .A2(n9177), .ZN(n4541) );
  XNOR2_X1 U11835 ( .A(n10146), .B(n9779), .ZN(n10080) );
  NAND3_X1 U11836 ( .A1(n9581), .A2(n9582), .A3(n9580), .ZN(n9779) );
  OAI21_X1 U11839 ( .B1(n18400), .B2(n18233), .A(n17976), .ZN(n4545) );
  INV_X1 U11840 ( .A(n18232), .ZN(n4546) );
  NAND2_X1 U11841 ( .A1(n29074), .A2(n23177), .ZN(n23564) );
  NAND2_X1 U11842 ( .A1(n4549), .A2(n15420), .ZN(n4548) );
  INV_X1 U11843 ( .A(n15103), .ZN(n4549) );
  NAND3_X1 U11844 ( .A1(n7823), .A2(n8222), .A3(n1842), .ZN(n4551) );
  NAND2_X1 U11845 ( .A1(n7821), .A2(n7424), .ZN(n4552) );
  NAND2_X1 U11846 ( .A1(n10101), .A2(n11132), .ZN(n4554) );
  INV_X1 U11847 ( .A(n10713), .ZN(n10499) );
  INV_X1 U11848 ( .A(n10711), .ZN(n4555) );
  INV_X1 U11849 ( .A(n20480), .ZN(n20476) );
  INV_X1 U11850 ( .A(n20479), .ZN(n4557) );
  NOR2_X2 U11851 ( .A1(n4558), .A2(n23898), .ZN(n25855) );
  AOI21_X1 U11852 ( .B1(n24368), .B2(n24367), .A(n24369), .ZN(n4559) );
  NAND2_X1 U11853 ( .A1(n379), .A2(n28581), .ZN(n4561) );
  NAND2_X1 U11854 ( .A1(n23268), .A2(n23611), .ZN(n4562) );
  NAND2_X1 U11855 ( .A1(n16541), .A2(n16812), .ZN(n17117) );
  NAND2_X1 U11856 ( .A1(n421), .A2(n4563), .ZN(n17460) );
  AND2_X1 U11857 ( .A1(n29539), .A2(n17459), .ZN(n4563) );
  NOR2_X1 U11858 ( .A1(n421), .A2(n29539), .ZN(n16101) );
  OR2_X1 U11859 ( .A1(n16813), .A2(n29539), .ZN(n4564) );
  NAND2_X1 U11860 ( .A1(n5295), .A2(n27855), .ZN(n27848) );
  NAND2_X1 U11861 ( .A1(n1916), .A2(n20601), .ZN(n4567) );
  NAND2_X1 U11862 ( .A1(n20457), .A2(n4567), .ZN(n20460) );
  NAND2_X1 U11863 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  MUX2_X1 U11864 ( .A(n18305), .B(n18306), .S(n18476), .Z(n15524) );
  NAND2_X1 U11865 ( .A1(n24795), .A2(n24796), .ZN(n4572) );
  NAND2_X1 U11866 ( .A1(n4574), .A2(n1955), .ZN(n4573) );
  NAND2_X1 U11867 ( .A1(n4576), .A2(n28455), .ZN(n4574) );
  OR2_X1 U11868 ( .A1(n7993), .A2(n7995), .ZN(n4578) );
  NAND2_X1 U11869 ( .A1(n7650), .A2(n4578), .ZN(n4577) );
  XNOR2_X1 U11870 ( .A(n4580), .B(n19652), .ZN(n4579) );
  INV_X1 U11871 ( .A(n19651), .ZN(n4580) );
  OAI211_X1 U11872 ( .C1(n17192), .C2(n17025), .A(n17346), .B(n4582), .ZN(
        n4583) );
  NAND2_X1 U11873 ( .A1(n17192), .A2(n17344), .ZN(n4582) );
  INV_X1 U11877 ( .A(n9074), .ZN(n4585) );
  XNOR2_X1 U11878 ( .A(n10005), .B(n9658), .ZN(n4592) );
  OAI21_X1 U11879 ( .B1(n23611), .B2(n28582), .A(n4593), .ZN(n4598) );
  NAND2_X1 U11880 ( .A1(n23611), .A2(n29115), .ZN(n4593) );
  NOR2_X1 U11881 ( .A1(n23217), .A2(n406), .ZN(n4596) );
  NOR2_X1 U11882 ( .A1(n23955), .A2(n4596), .ZN(n4594) );
  NAND2_X1 U11883 ( .A1(n4598), .A2(n4599), .ZN(n4597) );
  NAND2_X1 U11884 ( .A1(n4597), .A2(n4595), .ZN(n23956) );
  MUX2_X1 U11885 ( .A(n11052), .B(n10856), .S(n11163), .Z(n11055) );
  NAND3_X1 U11886 ( .A1(n4604), .A2(n24667), .A3(n24666), .ZN(n4603) );
  NAND2_X1 U11887 ( .A1(n24668), .A2(n4605), .ZN(n4604) );
  XNOR2_X1 U11888 ( .A(n16536), .B(n4606), .ZN(n15945) );
  XNOR2_X1 U11889 ( .A(n15727), .B(n4607), .ZN(n4606) );
  NOR2_X2 U11890 ( .A1(n15254), .A2(n15255), .ZN(n15727) );
  NAND2_X1 U11891 ( .A1(n13692), .A2(n5584), .ZN(n4608) );
  NOR2_X1 U11892 ( .A1(n15138), .A2(n14733), .ZN(n4611) );
  INV_X1 U11893 ( .A(n14733), .ZN(n15249) );
  NAND3_X1 U11894 ( .A1(n17001), .A2(n539), .A3(n16844), .ZN(n4612) );
  NAND2_X1 U11895 ( .A1(n4615), .A2(n4616), .ZN(n12868) );
  INV_X1 U11896 ( .A(n12241), .ZN(n12035) );
  INV_X1 U11897 ( .A(n14729), .ZN(n4621) );
  NAND2_X1 U11898 ( .A1(n17242), .A2(n16944), .ZN(n4625) );
  NAND2_X1 U11899 ( .A1(n29483), .A2(n17548), .ZN(n4626) );
  NAND2_X1 U11901 ( .A1(n28199), .A2(n13872), .ZN(n4627) );
  NAND2_X1 U11903 ( .A1(n6933), .A2(n21414), .ZN(n4631) );
  OAI21_X1 U11904 ( .B1(n490), .B2(n20663), .A(n21410), .ZN(n4633) );
  NAND2_X1 U11905 ( .A1(n4635), .A2(n4828), .ZN(n4634) );
  OAI21_X1 U11906 ( .B1(n21823), .B2(n20532), .A(n4636), .ZN(n4635) );
  NAND2_X1 U11907 ( .A1(n21823), .A2(n21078), .ZN(n4636) );
  NAND2_X1 U11909 ( .A1(n21819), .A2(n22013), .ZN(n4638) );
  INV_X1 U11910 ( .A(n4639), .ZN(n6835) );
  NAND2_X1 U11911 ( .A1(n4642), .A2(n4641), .ZN(n14547) );
  NAND3_X1 U11912 ( .A1(n4515), .A2(n15466), .A3(n29153), .ZN(n4641) );
  NAND2_X1 U11913 ( .A1(n4515), .A2(n15466), .ZN(n5016) );
  OAI21_X1 U11914 ( .B1(n4645), .B2(n26833), .A(n27442), .ZN(n4644) );
  AND2_X1 U11915 ( .A1(n27438), .A2(n26829), .ZN(n4645) );
  OAI21_X2 U11916 ( .B1(n25363), .B2(n26560), .A(n25362), .ZN(n27433) );
  NAND3_X1 U11917 ( .A1(n21750), .A2(n21237), .A3(n21399), .ZN(n4646) );
  NAND2_X1 U11918 ( .A1(n11316), .A2(n594), .ZN(n4650) );
  NAND2_X1 U11919 ( .A1(n17151), .A2(n17146), .ZN(n4654) );
  INV_X1 U11920 ( .A(n17489), .ZN(n4655) );
  AND2_X1 U11921 ( .A1(n20658), .A2(n4659), .ZN(n20659) );
  OR2_X1 U11922 ( .A1(n19921), .A2(n19920), .ZN(n4658) );
  XNOR2_X1 U11923 ( .A(n16494), .B(n16039), .ZN(n16351) );
  NAND2_X1 U11925 ( .A1(n6681), .A2(n15094), .ZN(n4661) );
  NAND2_X1 U11926 ( .A1(n4663), .A2(n24378), .ZN(n4662) );
  NOR2_X1 U11927 ( .A1(n24373), .A2(n24374), .ZN(n4663) );
  NAND2_X1 U11928 ( .A1(n24373), .A2(n24380), .ZN(n4664) );
  OAI21_X1 U11929 ( .B1(n14429), .B2(n28199), .A(n4665), .ZN(n12533) );
  XNOR2_X1 U11930 ( .A(n18991), .B(n19347), .ZN(n19353) );
  INV_X1 U11931 ( .A(n13008), .ZN(n4670) );
  INV_X1 U11932 ( .A(n13244), .ZN(n4669) );
  XNOR2_X1 U11933 ( .A(n4669), .B(n12686), .ZN(n12688) );
  XNOR2_X1 U11934 ( .A(n4670), .B(n12686), .ZN(n13010) );
  AOI21_X1 U11935 ( .B1(n5120), .B2(n7875), .A(n7958), .ZN(n4671) );
  OR2_X1 U11937 ( .A1(n4672), .A2(n23298), .ZN(n5940) );
  INV_X1 U11938 ( .A(n8192), .ZN(n4676) );
  NAND2_X1 U11939 ( .A1(n7095), .A2(n7868), .ZN(n4673) );
  NAND2_X1 U11940 ( .A1(n7861), .A2(n7094), .ZN(n4674) );
  NOR3_X1 U11941 ( .A1(n8828), .A2(n4676), .A3(n8586), .ZN(n8587) );
  NAND3_X1 U11942 ( .A1(n8826), .A2(n8827), .A3(n4676), .ZN(n8832) );
  NAND2_X1 U11943 ( .A1(n1839), .A2(n4676), .ZN(n8196) );
  OAI21_X1 U11944 ( .B1(n26431), .B2(n26382), .A(n26378), .ZN(n4678) );
  INV_X1 U11945 ( .A(n26275), .ZN(n4679) );
  INV_X1 U11946 ( .A(n17279), .ZN(n5968) );
  NAND2_X1 U11947 ( .A1(n539), .A2(n17272), .ZN(n17279) );
  OAI21_X1 U11948 ( .B1(n16665), .B2(n5968), .A(n4681), .ZN(n4680) );
  INV_X1 U11949 ( .A(n17271), .ZN(n4681) );
  NAND2_X1 U11950 ( .A1(n21253), .A2(n21811), .ZN(n21808) );
  NAND2_X1 U11951 ( .A1(n20117), .A2(n4684), .ZN(n4683) );
  AND2_X1 U11952 ( .A1(n4685), .A2(n24810), .ZN(n23692) );
  INV_X1 U11953 ( .A(n24812), .ZN(n4685) );
  AND2_X1 U11954 ( .A1(n17478), .A2(n4687), .ZN(n6560) );
  NAND2_X1 U11955 ( .A1(n17481), .A2(n1816), .ZN(n16690) );
  XNOR2_X1 U11956 ( .A(n4688), .B(n16579), .ZN(n6753) );
  XNOR2_X1 U11957 ( .A(n4688), .B(n1193), .ZN(n13670) );
  XNOR2_X1 U11958 ( .A(n16574), .B(n4688), .ZN(n15597) );
  XNOR2_X1 U11959 ( .A(n16318), .B(n4688), .ZN(n15703) );
  XNOR2_X1 U11960 ( .A(n16012), .B(n4688), .ZN(n15764) );
  XNOR2_X1 U11961 ( .A(n16255), .B(n4688), .ZN(n15825) );
  XNOR2_X1 U11962 ( .A(n16455), .B(n4688), .ZN(n16458) );
  NAND2_X1 U11964 ( .A1(n4693), .A2(n24279), .ZN(n4694) );
  INV_X1 U11965 ( .A(n7966), .ZN(n4696) );
  NAND2_X1 U11967 ( .A1(n16721), .A2(n17455), .ZN(n4699) );
  NAND3_X1 U11968 ( .A1(n4701), .A2(n4706), .A3(n28801), .ZN(n4700) );
  NAND2_X1 U11969 ( .A1(n4703), .A2(n17450), .ZN(n4701) );
  INV_X1 U11970 ( .A(n17065), .ZN(n4703) );
  NAND2_X1 U11972 ( .A1(n17065), .A2(n17452), .ZN(n4706) );
  NAND3_X1 U11973 ( .A1(n390), .A2(n4712), .A3(n11458), .ZN(n4711) );
  NOR2_X2 U11974 ( .A1(n10509), .A2(n10508), .ZN(n11458) );
  XNOR2_X1 U11976 ( .A(n4713), .B(n10263), .ZN(n9706) );
  XNOR2_X1 U11977 ( .A(n10191), .B(n4713), .ZN(n7329) );
  XNOR2_X1 U11978 ( .A(n4713), .B(n9318), .ZN(n9962) );
  XNOR2_X1 U11979 ( .A(n4714), .B(n10363), .ZN(n10086) );
  XNOR2_X1 U11980 ( .A(n4714), .B(n2325), .ZN(n9703) );
  XNOR2_X1 U11981 ( .A(n9266), .B(n4714), .ZN(n9268) );
  NOR2_X1 U11982 ( .A1(n10964), .A2(n4715), .ZN(n10967) );
  INV_X1 U11984 ( .A(n17569), .ZN(n4717) );
  OAI22_X1 U11985 ( .A1(n4719), .A2(n14998), .B1(n14747), .B2(n15132), .ZN(
        n4718) );
  NAND2_X1 U11986 ( .A1(n15132), .A2(n551), .ZN(n4719) );
  NAND2_X1 U11987 ( .A1(n14119), .A2(n4721), .ZN(n13625) );
  XNOR2_X2 U11988 ( .A(n12947), .B(n12946), .ZN(n6000) );
  INV_X1 U11989 ( .A(n23642), .ZN(n23641) );
  OAI21_X1 U11990 ( .B1(n21002), .B2(n21220), .A(n21001), .ZN(n4723) );
  NOR2_X2 U11991 ( .A1(n20702), .A2(n18753), .ZN(n21220) );
  NAND2_X1 U11992 ( .A1(n4722), .A2(n4724), .ZN(n20702) );
  NAND2_X1 U11993 ( .A1(n18574), .A2(n19844), .ZN(n4722) );
  AOI21_X2 U11994 ( .B1(n21003), .B2(n21220), .A(n4723), .ZN(n22912) );
  NAND2_X1 U11995 ( .A1(n18573), .A2(n29551), .ZN(n4724) );
  NAND2_X1 U11996 ( .A1(n6379), .A2(n17286), .ZN(n18236) );
  AND2_X1 U11997 ( .A1(n1914), .A2(n23802), .ZN(n5192) );
  NOR2_X1 U11998 ( .A1(n1914), .A2(n23689), .ZN(n23540) );
  AOI21_X1 U11999 ( .B1(n23689), .B2(n23802), .A(n1914), .ZN(n23175) );
  NAND2_X1 U12000 ( .A1(n29598), .A2(n16811), .ZN(n17118) );
  NAND2_X1 U12002 ( .A1(n4729), .A2(n597), .ZN(n4728) );
  INV_X1 U12003 ( .A(n9825), .ZN(n9603) );
  NAND2_X1 U12004 ( .A1(n5569), .A2(n5160), .ZN(n4731) );
  NAND2_X1 U12006 ( .A1(n17846), .A2(n17847), .ZN(n4732) );
  NAND2_X1 U12007 ( .A1(n21574), .A2(n21575), .ZN(n20848) );
  NAND2_X1 U12009 ( .A1(n13891), .A2(n14444), .ZN(n13685) );
  NOR2_X1 U12010 ( .A1(n28647), .A2(n14414), .ZN(n6232) );
  NAND2_X1 U12011 ( .A1(n14419), .A2(n28648), .ZN(n13687) );
  XNOR2_X1 U12013 ( .A(n8648), .B(n8647), .ZN(n10334) );
  NAND2_X1 U12014 ( .A1(n4836), .A2(n13894), .ZN(n15463) );
  NOR2_X2 U12015 ( .A1(n21776), .A2(n4735), .ZN(n24596) );
  NAND2_X1 U12016 ( .A1(n4737), .A2(n4736), .ZN(n4735) );
  NAND3_X1 U12017 ( .A1(n23788), .A2(n23036), .A3(n473), .ZN(n4736) );
  NAND2_X1 U12018 ( .A1(n21769), .A2(n23482), .ZN(n4737) );
  XNOR2_X1 U12019 ( .A(n21994), .B(n20885), .ZN(n4738) );
  XNOR2_X1 U12020 ( .A(n21761), .B(n4738), .ZN(n21764) );
  INV_X1 U12021 ( .A(n4738), .ZN(n21760) );
  AND2_X1 U12022 ( .A1(n455), .A2(n27701), .ZN(n4741) );
  AOI21_X1 U12024 ( .B1(n27175), .B2(n26263), .A(n28480), .ZN(n26265) );
  OAI21_X1 U12027 ( .B1(n10717), .B2(n28436), .A(n4744), .ZN(n11791) );
  AOI22_X1 U12028 ( .A1(n11720), .A2(n10717), .B1(n11719), .B2(n4744), .ZN(
        n11721) );
  NAND2_X1 U12030 ( .A1(n24596), .A2(n24597), .ZN(n4748) );
  NAND2_X1 U12031 ( .A1(n4752), .A2(n4750), .ZN(n26571) );
  NAND2_X1 U12032 ( .A1(n26566), .A2(n29610), .ZN(n4752) );
  NAND2_X1 U12033 ( .A1(n28775), .A2(n17179), .ZN(n17377) );
  XNOR2_X1 U12035 ( .A(n16340), .B(n1979), .ZN(n4753) );
  NAND2_X1 U12036 ( .A1(n23968), .A2(n24484), .ZN(n24486) );
  NAND3_X1 U12039 ( .A1(n4757), .A2(n17353), .A3(n28558), .ZN(n4756) );
  INV_X1 U12040 ( .A(n18404), .ZN(n4757) );
  XNOR2_X1 U12044 ( .A(n22008), .B(n21804), .ZN(n4760) );
  INV_X1 U12045 ( .A(n18431), .ZN(n4762) );
  XNOR2_X1 U12047 ( .A(n4764), .B(n25890), .ZN(n25072) );
  XNOR2_X1 U12048 ( .A(n4764), .B(n25381), .ZN(n25817) );
  XNOR2_X1 U12049 ( .A(n16510), .B(n16176), .ZN(n4811) );
  XNOR2_X1 U12050 ( .A(n15909), .B(n16000), .ZN(n4767) );
  XNOR2_X1 U12051 ( .A(n16031), .B(n4811), .ZN(n4765) );
  NAND2_X1 U12052 ( .A1(n23011), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U12054 ( .A1(n5774), .A2(n23010), .ZN(n23546) );
  NAND2_X1 U12055 ( .A1(n6227), .A2(n23351), .ZN(n4773) );
  NAND2_X1 U12056 ( .A1(n18710), .A2(n18404), .ZN(n4774) );
  OR2_X1 U12057 ( .A1(n18248), .A2(n18708), .ZN(n18710) );
  NAND2_X1 U12058 ( .A1(n20339), .A2(n20504), .ZN(n20226) );
  INV_X1 U12059 ( .A(n4776), .ZN(n20909) );
  XNOR2_X1 U12061 ( .A(n16443), .B(n16262), .ZN(n4777) );
  XNOR2_X1 U12062 ( .A(n4777), .B(n15592), .ZN(n15593) );
  INV_X1 U12063 ( .A(n4777), .ZN(n15720) );
  NAND2_X1 U12064 ( .A1(n4780), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U12065 ( .A1(n14325), .A2(n14323), .ZN(n4779) );
  INV_X1 U12066 ( .A(n24578), .ZN(n4784) );
  NAND3_X1 U12067 ( .A1(n4784), .A2(n29025), .A3(n24581), .ZN(n4783) );
  NAND2_X1 U12068 ( .A1(n24581), .A2(n29025), .ZN(n24055) );
  NOR2_X1 U12069 ( .A1(n4786), .A2(n4953), .ZN(n4785) );
  NOR2_X2 U12070 ( .A1(n20318), .A2(n20317), .ZN(n21306) );
  OAI21_X1 U12071 ( .B1(n10804), .B2(n4788), .A(n6745), .ZN(n4789) );
  NAND2_X1 U12072 ( .A1(n593), .A2(n5150), .ZN(n6745) );
  NAND2_X1 U12073 ( .A1(n11153), .A2(n11158), .ZN(n4788) );
  NAND2_X1 U12074 ( .A1(n11158), .A2(n11154), .ZN(n10803) );
  XNOR2_X2 U12075 ( .A(n6184), .B(n6183), .ZN(n11158) );
  INV_X1 U12077 ( .A(n6745), .ZN(n11159) );
  AOI21_X1 U12078 ( .B1(n10802), .B2(n10803), .A(n11153), .ZN(n4790) );
  NAND2_X1 U12079 ( .A1(n4791), .A2(n14824), .ZN(n14779) );
  NAND2_X1 U12080 ( .A1(n15433), .A2(n4791), .ZN(n15894) );
  NAND2_X1 U12081 ( .A1(n15027), .A2(n15431), .ZN(n4791) );
  NAND2_X1 U12082 ( .A1(n20242), .A2(n20241), .ZN(n4793) );
  OAI21_X1 U12084 ( .B1(n18441), .B2(n4929), .A(n4796), .ZN(n18185) );
  NAND2_X1 U12085 ( .A1(n4929), .A2(n18178), .ZN(n4796) );
  AND2_X1 U12086 ( .A1(n5973), .A2(n12075), .ZN(n4797) );
  OAI21_X2 U12087 ( .B1(n4797), .B2(n5947), .A(n4798), .ZN(n12677) );
  NAND2_X1 U12088 ( .A1(n12076), .A2(n12575), .ZN(n4798) );
  INV_X1 U12089 ( .A(n12578), .ZN(n12575) );
  AND3_X2 U12090 ( .A1(n6438), .A2(n1996), .A3(n6437), .ZN(n27520) );
  NAND2_X1 U12091 ( .A1(n4801), .A2(n29149), .ZN(n4800) );
  XNOR2_X1 U12092 ( .A(n4806), .B(n9590), .ZN(n9595) );
  INV_X1 U12093 ( .A(n9591), .ZN(n4806) );
  XNOR2_X1 U12094 ( .A(n4807), .B(n9940), .ZN(n9945) );
  NOR2_X1 U12095 ( .A1(n27502), .A2(n4808), .ZN(n27223) );
  NAND2_X1 U12096 ( .A1(n4809), .A2(n27520), .ZN(n4808) );
  AOI22_X2 U12097 ( .A1(n23931), .A2(n24591), .B1(n23930), .B2(n23929), .ZN(
        n25249) );
  XNOR2_X1 U12098 ( .A(n4811), .B(n14223), .ZN(n14224) );
  INV_X1 U12099 ( .A(n16510), .ZN(n16642) );
  OAI21_X1 U12100 ( .B1(n564), .B2(n4812), .A(n14367), .ZN(n14371) );
  NAND2_X1 U12102 ( .A1(n4814), .A2(n20373), .ZN(n4813) );
  NAND2_X1 U12103 ( .A1(n20070), .A2(n20071), .ZN(n4814) );
  NAND2_X1 U12104 ( .A1(n18843), .A2(n18699), .ZN(n20071) );
  NOR2_X2 U12106 ( .A1(n4817), .A2(n4816), .ZN(n27447) );
  NAND2_X1 U12107 ( .A1(n4820), .A2(n26172), .ZN(n4819) );
  XNOR2_X1 U12108 ( .A(n4821), .B(n26176), .ZN(Ciphertext[47]) );
  NAND2_X1 U12109 ( .A1(n26175), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U12110 ( .A1(n26606), .A2(n4823), .ZN(n4822) );
  NAND2_X1 U12112 ( .A1(n7643), .A2(n7981), .ZN(n4826) );
  NAND2_X1 U12114 ( .A1(n4831), .A2(n28801), .ZN(n4829) );
  NAND2_X1 U12115 ( .A1(n17069), .A2(n17068), .ZN(n4830) );
  OAI21_X1 U12116 ( .B1(n4832), .B2(n26450), .A(n26179), .ZN(n6124) );
  AOI21_X1 U12117 ( .B1(n25622), .B2(n29105), .A(n4832), .ZN(n24039) );
  NAND3_X1 U12118 ( .A1(n7982), .A2(n7644), .A3(n7980), .ZN(n4833) );
  NAND3_X1 U12119 ( .A1(n7642), .A2(n7644), .A3(n7641), .ZN(n4834) );
  MUX2_X1 U12122 ( .A(n4515), .B(n29153), .S(n15463), .Z(n4835) );
  XNOR2_X1 U12124 ( .A(n19668), .B(n18927), .ZN(n4838) );
  XNOR2_X1 U12125 ( .A(n12726), .B(n12725), .ZN(n14469) );
  INV_X1 U12126 ( .A(n12743), .ZN(n4840) );
  NAND2_X1 U12127 ( .A1(n4842), .A2(n4841), .ZN(n12799) );
  NAND2_X1 U12128 ( .A1(n11702), .A2(n12201), .ZN(n4841) );
  NAND2_X1 U12129 ( .A1(n16889), .A2(n16888), .ZN(n4845) );
  NAND2_X1 U12130 ( .A1(n17088), .A2(n17137), .ZN(n4846) );
  OAI21_X1 U12131 ( .B1(n23546), .B2(n4232), .A(n4851), .ZN(n4850) );
  INV_X1 U12132 ( .A(n4850), .ZN(n4849) );
  NAND2_X1 U12133 ( .A1(n15162), .A2(n4515), .ZN(n4853) );
  NAND3_X1 U12135 ( .A1(n7758), .A2(n8176), .A3(n4856), .ZN(n7180) );
  OR2_X1 U12136 ( .A1(n8175), .A2(n4856), .ZN(n7182) );
  INV_X1 U12137 ( .A(n7759), .ZN(n4856) );
  MUX2_X1 U12138 ( .A(n24081), .B(n24079), .S(n24078), .Z(n4857) );
  NAND2_X1 U12139 ( .A1(n4859), .A2(n29470), .ZN(n4858) );
  NAND2_X1 U12140 ( .A1(n5728), .A2(n24388), .ZN(n4859) );
  INV_X1 U12141 ( .A(Key[101]), .ZN(n4861) );
  XNOR2_X1 U12142 ( .A(n21994), .B(n4862), .ZN(n21384) );
  OAI21_X1 U12143 ( .B1(n17017), .B2(n17249), .A(n17251), .ZN(n4865) );
  NAND2_X1 U12144 ( .A1(n17016), .A2(n4863), .ZN(n4864) );
  AOI21_X1 U12145 ( .B1(n12272), .B2(n12578), .A(n11940), .ZN(n4868) );
  NAND2_X1 U12146 ( .A1(n4867), .A2(n4870), .ZN(n12453) );
  NAND2_X1 U12147 ( .A1(n12274), .A2(n11940), .ZN(n4870) );
  NAND2_X1 U12152 ( .A1(n20147), .A2(n4875), .ZN(n4874) );
  OAI21_X1 U12153 ( .B1(n29134), .B2(n4877), .A(n4876), .ZN(n4875) );
  NAND2_X1 U12154 ( .A1(n28479), .A2(n21096), .ZN(n4878) );
  XNOR2_X1 U12156 ( .A(n4880), .B(n19025), .ZN(n18581) );
  XNOR2_X1 U12157 ( .A(n19025), .B(n4881), .ZN(n17850) );
  XNOR2_X1 U12158 ( .A(n19025), .B(n4882), .ZN(n18640) );
  INV_X1 U12159 ( .A(n1119), .ZN(n4882) );
  NOR2_X1 U12160 ( .A1(n20054), .A2(n6114), .ZN(n4885) );
  INV_X1 U12161 ( .A(n20172), .ZN(n4886) );
  NAND2_X1 U12162 ( .A1(n4888), .A2(n4889), .ZN(n4887) );
  NAND2_X1 U12165 ( .A1(n23150), .A2(n23459), .ZN(n4891) );
  MUX2_X1 U12166 ( .A(n4364), .B(n24629), .S(n24533), .Z(n23984) );
  OAI21_X1 U12167 ( .B1(n13826), .B2(n13060), .A(n4893), .ZN(n4895) );
  NAND2_X1 U12168 ( .A1(n6872), .A2(n14127), .ZN(n4894) );
  NAND2_X1 U12170 ( .A1(n17382), .A2(n16878), .ZN(n4900) );
  NAND2_X1 U12171 ( .A1(n17388), .A2(n17389), .ZN(n4901) );
  NAND2_X1 U12172 ( .A1(n5532), .A2(n10847), .ZN(n4904) );
  MUX2_X1 U12173 ( .A(n21698), .B(n29101), .S(n6314), .Z(n18549) );
  MUX2_X1 U12174 ( .A(n21243), .B(n21244), .S(n6314), .Z(n21247) );
  NAND2_X1 U12175 ( .A1(n11090), .A2(n10431), .ZN(n4908) );
  NAND2_X1 U12176 ( .A1(n4908), .A2(n29517), .ZN(n4907) );
  NAND2_X1 U12177 ( .A1(n20345), .A2(n19786), .ZN(n4910) );
  NAND2_X1 U12178 ( .A1(n5853), .A2(n20014), .ZN(n4911) );
  OAI21_X1 U12179 ( .B1(n21560), .B2(n21561), .A(n21113), .ZN(n21114) );
  INV_X1 U12180 ( .A(n28578), .ZN(n4913) );
  MUX2_X1 U12181 ( .A(n28434), .B(n28385), .S(n28578), .Z(n25363) );
  OAI22_X1 U12183 ( .A1(n23447), .A2(n23445), .B1(n23446), .B2(n292), .ZN(
        n4915) );
  INV_X1 U12184 ( .A(n14797), .ZN(n14980) );
  NAND2_X1 U12185 ( .A1(n4917), .A2(n24552), .ZN(n24553) );
  MUX2_X1 U12186 ( .A(n4917), .B(n28519), .S(n24552), .Z(n22868) );
  OAI22_X1 U12187 ( .A1(n23205), .A2(n4917), .B1(n24551), .B2(n24173), .ZN(
        n23936) );
  NAND2_X1 U12188 ( .A1(n23937), .A2(n4917), .ZN(n6121) );
  MUX2_X1 U12189 ( .A(n23976), .B(n23977), .S(n22869), .Z(n23978) );
  XNOR2_X1 U12190 ( .A(n4918), .B(n4923), .ZN(Ciphertext[21]) );
  NAND2_X1 U12191 ( .A1(n4921), .A2(n4922), .ZN(n4919) );
  NAND3_X1 U12193 ( .A1(n27242), .A2(n27386), .A3(n28177), .ZN(n4924) );
  AND2_X1 U12194 ( .A1(n29138), .A2(n17229), .ZN(n6292) );
  OR2_X1 U12195 ( .A1(n18442), .A2(n18181), .ZN(n4927) );
  INV_X1 U12196 ( .A(n19252), .ZN(n19383) );
  NAND2_X1 U12197 ( .A1(n2039), .A2(n16763), .ZN(n4930) );
  AOI21_X1 U12198 ( .B1(n8998), .B2(n9438), .A(n9211), .ZN(n4931) );
  NAND2_X1 U12199 ( .A1(n8776), .A2(n8996), .ZN(n4932) );
  INV_X1 U12200 ( .A(n9434), .ZN(n8998) );
  NAND2_X1 U12202 ( .A1(n5742), .A2(n5741), .ZN(n4934) );
  NAND2_X1 U12203 ( .A1(n23033), .A2(n4936), .ZN(n4935) );
  NOR2_X1 U12204 ( .A1(n23758), .A2(n29131), .ZN(n4936) );
  INV_X1 U12205 ( .A(n4937), .ZN(n21414) );
  NOR2_X1 U12206 ( .A1(n28184), .A2(n4937), .ZN(n21052) );
  NAND2_X1 U12207 ( .A1(n21230), .A2(n4937), .ZN(n21176) );
  NAND2_X1 U12208 ( .A1(n7774), .A2(n7889), .ZN(n4939) );
  INV_X1 U12209 ( .A(n8048), .ZN(n4942) );
  NAND2_X1 U12210 ( .A1(n8132), .A2(n8131), .ZN(n4940) );
  NAND2_X1 U12211 ( .A1(n4942), .A2(n7554), .ZN(n4941) );
  NAND2_X1 U12212 ( .A1(n26426), .A2(n26378), .ZN(n4944) );
  NAND2_X1 U12214 ( .A1(n17555), .A2(n16913), .ZN(n16917) );
  XNOR2_X1 U12215 ( .A(n4946), .B(n27550), .ZN(Ciphertext[77]) );
  NAND2_X1 U12216 ( .A1(n4948), .A2(n4947), .ZN(n4946) );
  OAI21_X1 U12217 ( .B1(n5540), .B2(n27548), .A(n27547), .ZN(n4947) );
  NOR2_X1 U12218 ( .A1(n27537), .A2(n27202), .ZN(n5540) );
  OAI21_X1 U12219 ( .B1(n27545), .B2(n27546), .A(n394), .ZN(n4948) );
  NAND2_X1 U12223 ( .A1(n22851), .A2(n28182), .ZN(n4951) );
  NOR2_X1 U12224 ( .A1(n17792), .A2(n17793), .ZN(n4953) );
  INV_X1 U12225 ( .A(n16332), .ZN(n4956) );
  XNOR2_X1 U12226 ( .A(n4956), .B(n15545), .ZN(n16376) );
  OR2_X2 U12229 ( .A1(n14089), .A2(n14090), .ZN(n15290) );
  INV_X1 U12230 ( .A(n14285), .ZN(n14282) );
  AOI21_X1 U12233 ( .B1(n17502), .B2(n6727), .A(n17501), .ZN(n4963) );
  NAND2_X1 U12234 ( .A1(n24378), .A2(n24380), .ZN(n23377) );
  XNOR2_X1 U12235 ( .A(n16596), .B(n15989), .ZN(n4965) );
  XNOR2_X1 U12236 ( .A(n4965), .B(n16193), .ZN(n16194) );
  INV_X1 U12237 ( .A(n4965), .ZN(n15561) );
  NAND2_X1 U12238 ( .A1(n24592), .A2(n24591), .ZN(n4966) );
  NAND3_X1 U12239 ( .A1(n24143), .A2(n24144), .A3(n4693), .ZN(n24145) );
  XNOR2_X1 U12240 ( .A(n22008), .B(n22238), .ZN(n4967) );
  INV_X1 U12241 ( .A(n4971), .ZN(n4970) );
  NOR2_X1 U12242 ( .A1(n11154), .A2(n11158), .ZN(n4972) );
  NOR2_X1 U12243 ( .A1(n14336), .A2(n5584), .ZN(n4975) );
  NOR2_X1 U12244 ( .A1(n1830), .A2(n4974), .ZN(n4973) );
  NAND2_X1 U12245 ( .A1(n4975), .A2(n14408), .ZN(n13882) );
  XNOR2_X1 U12246 ( .A(n19305), .B(n19306), .ZN(n19308) );
  XNOR2_X1 U12247 ( .A(n15727), .B(n4978), .ZN(n4977) );
  NAND2_X1 U12248 ( .A1(n16430), .A2(n4979), .ZN(n17185) );
  NAND2_X1 U12249 ( .A1(n2483), .A2(n12127), .ZN(n4981) );
  NAND2_X1 U12250 ( .A1(n8670), .A2(n9107), .ZN(n8672) );
  NAND3_X1 U12251 ( .A1(n8670), .A2(n8914), .A3(n9107), .ZN(n8514) );
  NAND2_X1 U12252 ( .A1(n9106), .A2(n8670), .ZN(n9121) );
  OAI21_X2 U12253 ( .B1(n28186), .B2(n4984), .A(n19329), .ZN(n21714) );
  OAI21_X1 U12254 ( .B1(n20334), .B2(n20626), .A(n4985), .ZN(n4984) );
  NAND2_X1 U12255 ( .A1(n20623), .A2(n20626), .ZN(n4985) );
  NAND2_X1 U12256 ( .A1(n4986), .A2(n18398), .ZN(n5757) );
  NAND2_X1 U12257 ( .A1(n18233), .A2(n18231), .ZN(n4986) );
  NAND2_X1 U12259 ( .A1(n5460), .A2(n17434), .ZN(n4987) );
  NAND2_X1 U12261 ( .A1(n6605), .A2(n20498), .ZN(n4991) );
  AND2_X2 U12262 ( .A1(n20010), .A2(n20011), .ZN(n21638) );
  MUX2_X1 U12263 ( .A(n4992), .B(n15243), .S(n15359), .Z(n14508) );
  AOI22_X1 U12264 ( .A1(n15061), .A2(n4992), .B1(n15359), .B2(n15062), .ZN(
        n15063) );
  OAI21_X1 U12265 ( .B1(n15358), .B2(n28197), .A(n4992), .ZN(n6003) );
  MUX2_X1 U12266 ( .A(n24240), .B(n24559), .S(n24633), .Z(n4993) );
  NAND2_X1 U12267 ( .A1(n23558), .A2(n23188), .ZN(n4994) );
  NAND2_X1 U12268 ( .A1(n23989), .A2(n24557), .ZN(n4995) );
  NAND2_X1 U12269 ( .A1(n5966), .A2(n11435), .ZN(n4996) );
  INV_X1 U12270 ( .A(n27938), .ZN(n4998) );
  OAI211_X1 U12271 ( .C1(n27942), .C2(n27941), .A(n27940), .B(n4999), .ZN(
        n27943) );
  NAND2_X1 U12272 ( .A1(n5000), .A2(n20899), .ZN(n20141) );
  NOR2_X1 U12273 ( .A1(n1925), .A2(n5000), .ZN(n20143) );
  NOR2_X1 U12274 ( .A1(n17254), .A2(n1880), .ZN(n17256) );
  INV_X1 U12275 ( .A(n17249), .ZN(n5001) );
  XNOR2_X1 U12276 ( .A(n13474), .B(n12473), .ZN(n5002) );
  XNOR2_X1 U12277 ( .A(n12474), .B(n12471), .ZN(n5003) );
  NAND3_X1 U12278 ( .A1(n28441), .A2(n28438), .A3(n27944), .ZN(n27940) );
  NAND3_X1 U12279 ( .A1(n4998), .A2(n28439), .A3(n27941), .ZN(n27928) );
  MUX2_X1 U12280 ( .A(n28438), .B(n27941), .S(n27925), .Z(n27245) );
  MUX2_X1 U12281 ( .A(n27244), .B(n27925), .S(n28439), .Z(n27023) );
  NAND2_X1 U12282 ( .A1(n27932), .A2(n2060), .ZN(n27933) );
  XNOR2_X1 U12283 ( .A(n19693), .B(n19694), .ZN(n5005) );
  AND3_X1 U12284 ( .A1(n12234), .A2(n12236), .A3(n12233), .ZN(n5007) );
  NAND2_X1 U12285 ( .A1(n12234), .A2(n12233), .ZN(n12235) );
  AOI21_X1 U12286 ( .B1(n5009), .B2(n5008), .A(n5007), .ZN(n5012) );
  INV_X1 U12287 ( .A(n1986), .ZN(n5009) );
  NAND2_X1 U12288 ( .A1(n5012), .A2(n5010), .ZN(n12472) );
  NAND2_X1 U12289 ( .A1(n5011), .A2(n1986), .ZN(n5010) );
  OAI21_X1 U12290 ( .B1(n776), .B2(n12232), .A(n12234), .ZN(n5011) );
  NAND2_X1 U12291 ( .A1(n20900), .A2(n21084), .ZN(n5013) );
  INV_X1 U12292 ( .A(n15463), .ZN(n15161) );
  INV_X1 U12293 ( .A(n15464), .ZN(n14652) );
  INV_X1 U12294 ( .A(n28024), .ZN(n28034) );
  NOR2_X1 U12295 ( .A1(n28026), .A2(n5017), .ZN(n28031) );
  INV_X1 U12297 ( .A(n20865), .ZN(n21185) );
  INV_X1 U12298 ( .A(n22132), .ZN(n22723) );
  OR2_X1 U12299 ( .A1(n20187), .A2(n20186), .ZN(n5018) );
  AOI22_X2 U12300 ( .A1(n5020), .A2(n10701), .B1(n5019), .B2(n11768), .ZN(
        n13014) );
  INV_X1 U12301 ( .A(n18708), .ZN(n5021) );
  NAND2_X1 U12302 ( .A1(n5025), .A2(n15404), .ZN(n5024) );
  NAND2_X1 U12304 ( .A1(n28195), .A2(n15402), .ZN(n15398) );
  INV_X1 U12306 ( .A(n23067), .ZN(n23693) );
  NAND2_X1 U12307 ( .A1(n23693), .A2(n23531), .ZN(n5028) );
  INV_X1 U12308 ( .A(n23531), .ZN(n5030) );
  INV_X1 U12310 ( .A(n23531), .ZN(n23696) );
  XNOR2_X1 U12311 ( .A(n10421), .B(n2035), .ZN(n9617) );
  XNOR2_X1 U12312 ( .A(n10421), .B(n5032), .ZN(n9386) );
  NAND2_X1 U12313 ( .A1(n20156), .A2(n20155), .ZN(n5033) );
  AOI21_X1 U12314 ( .B1(n1121), .B2(n17347), .A(n542), .ZN(n16951) );
  NAND2_X1 U12315 ( .A1(n29100), .A2(n26748), .ZN(n5036) );
  NAND3_X1 U12316 ( .A1(n12134), .A2(n12265), .A3(n12133), .ZN(n5038) );
  MUX2_X1 U12317 ( .A(n12267), .B(n12132), .S(n11574), .Z(n5040) );
  NAND2_X1 U12320 ( .A1(n5042), .A2(n23405), .ZN(n5041) );
  XNOR2_X1 U12321 ( .A(n5043), .B(n22584), .ZN(n22032) );
  NAND3_X1 U12322 ( .A1(n5046), .A2(n22029), .A3(n5044), .ZN(n5043) );
  NAND2_X1 U12323 ( .A1(n5045), .A2(n28108), .ZN(n5044) );
  INV_X1 U12324 ( .A(n22030), .ZN(n5045) );
  NAND4_X1 U12325 ( .A1(n22294), .A2(n1927), .A3(n22030), .A4(n5047), .ZN(
        n5046) );
  INV_X1 U12326 ( .A(n22028), .ZN(n5047) );
  NAND3_X1 U12328 ( .A1(n15512), .A2(n15514), .A3(n15515), .ZN(n5051) );
  INV_X1 U12329 ( .A(n15275), .ZN(n5049) );
  NAND2_X1 U12330 ( .A1(n15274), .A2(n15275), .ZN(n14920) );
  NAND2_X1 U12331 ( .A1(n5048), .A2(n15274), .ZN(n5050) );
  NOR2_X1 U12332 ( .A1(n5049), .A2(n15514), .ZN(n5048) );
  NAND2_X1 U12333 ( .A1(n15279), .A2(n15512), .ZN(n5052) );
  OAI21_X1 U12334 ( .B1(n20152), .B2(n5053), .A(n20098), .ZN(n5054) );
  INV_X1 U12335 ( .A(n20150), .ZN(n5053) );
  NAND2_X1 U12336 ( .A1(n20042), .A2(n20096), .ZN(n5055) );
  INV_X1 U12337 ( .A(n20098), .ZN(n5056) );
  AOI21_X1 U12338 ( .B1(n14375), .B2(n14374), .A(n5057), .ZN(n14378) );
  INV_X1 U12339 ( .A(n13725), .ZN(n5058) );
  NAND2_X1 U12340 ( .A1(n16852), .A2(n16853), .ZN(n16854) );
  INV_X1 U12341 ( .A(n18761), .ZN(n18949) );
  OAI211_X1 U12342 ( .C1(n16868), .C2(n5059), .A(n5061), .B(n5060), .ZN(n5062)
         );
  NAND3_X1 U12343 ( .A1(n16868), .A2(n16867), .A3(n5059), .ZN(n5061) );
  XNOR2_X1 U12344 ( .A(n29136), .B(n5067), .ZN(n5066) );
  XNOR2_X1 U12345 ( .A(n22000), .B(n22896), .ZN(n5067) );
  NAND2_X1 U12346 ( .A1(n5068), .A2(n16968), .ZN(n16792) );
  XNOR2_X2 U12347 ( .A(n15111), .B(n15112), .ZN(n17304) );
  XNOR2_X1 U12348 ( .A(n5069), .B(n13055), .ZN(n12833) );
  XNOR2_X1 U12350 ( .A(n12593), .B(n5070), .ZN(n13569) );
  INV_X1 U12351 ( .A(n13566), .ZN(n5070) );
  NAND2_X1 U12352 ( .A1(n7515), .A2(n29321), .ZN(n7261) );
  OAI22_X1 U12353 ( .A1(n29201), .A2(n1959), .B1(n3269), .B2(n14394), .ZN(
        n5073) );
  NAND2_X1 U12354 ( .A1(n1952), .A2(n29104), .ZN(n5074) );
  NAND3_X1 U12355 ( .A1(n28820), .A2(n20091), .A3(n20039), .ZN(n5075) );
  NAND2_X1 U12356 ( .A1(n5078), .A2(n5077), .ZN(n5076) );
  NAND3_X1 U12357 ( .A1(n11515), .A2(n11671), .A3(n29139), .ZN(n5077) );
  NAND2_X1 U12358 ( .A1(n11632), .A2(n11634), .ZN(n11515) );
  NAND2_X1 U12359 ( .A1(n11406), .A2(n5079), .ZN(n5078) );
  NAND3_X1 U12360 ( .A1(n5080), .A2(n24093), .A3(n24091), .ZN(n24097) );
  NAND2_X1 U12361 ( .A1(n17798), .A2(n18106), .ZN(n18457) );
  MUX2_X1 U12362 ( .A(n23862), .B(n26572), .S(n25418), .Z(n26573) );
  NAND2_X1 U12364 ( .A1(n518), .A2(n18354), .ZN(n5083) );
  INV_X1 U12365 ( .A(n18353), .ZN(n6225) );
  NAND3_X1 U12367 ( .A1(n21180), .A2(n21551), .A3(n20351), .ZN(n5086) );
  NAND3_X1 U12368 ( .A1(n5088), .A2(n5087), .A3(n5086), .ZN(n22792) );
  NAND2_X1 U12369 ( .A1(n2067), .A2(n21553), .ZN(n5088) );
  OR2_X1 U12370 ( .A1(n10116), .A2(n11127), .ZN(n5089) );
  NAND2_X1 U12371 ( .A1(n6833), .A2(n5090), .ZN(n6832) );
  NAND2_X1 U12372 ( .A1(n15374), .A2(n15376), .ZN(n5092) );
  INV_X1 U12373 ( .A(n18034), .ZN(n18158) );
  MUX2_X1 U12375 ( .A(n11970), .B(n5097), .S(n12159), .Z(n5095) );
  NAND2_X1 U12376 ( .A1(n5098), .A2(n4617), .ZN(n5096) );
  NAND2_X1 U12377 ( .A1(n12244), .A2(n12158), .ZN(n5097) );
  MUX2_X1 U12378 ( .A(n12156), .B(n12241), .S(n12244), .Z(n5098) );
  NAND3_X1 U12379 ( .A1(n97), .A2(n28637), .A3(n20383), .ZN(n5099) );
  NAND2_X1 U12380 ( .A1(n5103), .A2(n5102), .ZN(n5101) );
  NAND2_X1 U12381 ( .A1(n24631), .A2(n23144), .ZN(n5102) );
  INV_X1 U12382 ( .A(n24531), .ZN(n5103) );
  NOR2_X1 U12383 ( .A1(n24530), .A2(n24533), .ZN(n5105) );
  XNOR2_X1 U12384 ( .A(n18321), .B(n18320), .ZN(n20539) );
  INV_X1 U12385 ( .A(n20539), .ZN(n20389) );
  INV_X1 U12386 ( .A(n19959), .ZN(n20188) );
  NAND2_X1 U12387 ( .A1(n20223), .A2(n5106), .ZN(n19861) );
  INV_X1 U12388 ( .A(n17989), .ZN(n18367) );
  NAND2_X1 U12391 ( .A1(n27077), .A2(n5113), .ZN(n5112) );
  NOR2_X1 U12392 ( .A1(n26991), .A2(n5263), .ZN(n5113) );
  INV_X1 U12393 ( .A(n26994), .ZN(n5114) );
  NOR2_X1 U12395 ( .A1(n24277), .A2(n24591), .ZN(n5116) );
  NAND2_X1 U12396 ( .A1(n24593), .A2(n5116), .ZN(n5115) );
  INV_X1 U12398 ( .A(n12929), .ZN(n5121) );
  XNOR2_X1 U12399 ( .A(n12882), .B(n5121), .ZN(n5122) );
  OAI21_X1 U12400 ( .B1(n1876), .B2(n14440), .A(n14433), .ZN(n14436) );
  NAND2_X1 U12401 ( .A1(n21823), .A2(n22013), .ZN(n5123) );
  NAND2_X1 U12402 ( .A1(n4828), .A2(n5125), .ZN(n5124) );
  NAND2_X1 U12403 ( .A1(n6495), .A2(n29551), .ZN(n5126) );
  MUX2_X1 U12404 ( .A(n5053), .B(n20151), .S(n20152), .Z(n19775) );
  MUX2_X1 U12405 ( .A(n20152), .B(n20151), .S(n20150), .Z(n18888) );
  AOI21_X1 U12406 ( .B1(n20096), .B2(n20155), .A(n5053), .ZN(n18833) );
  XNOR2_X1 U12407 ( .A(n17597), .B(n5127), .ZN(n17606) );
  INV_X1 U12408 ( .A(n18556), .ZN(n5127) );
  XNOR2_X1 U12409 ( .A(n18725), .B(n19139), .ZN(n18556) );
  NAND3_X1 U12410 ( .A1(n21143), .A2(n21119), .A3(n21140), .ZN(n5128) );
  INV_X1 U12411 ( .A(n7569), .ZN(n5129) );
  NAND2_X1 U12412 ( .A1(n5131), .A2(n603), .ZN(n5130) );
  OAI21_X1 U12413 ( .B1(n9425), .B2(n7569), .A(n5132), .ZN(n5131) );
  NAND3_X1 U12414 ( .A1(n11902), .A2(n12428), .A3(n5134), .ZN(n11905) );
  XNOR2_X1 U12415 ( .A(n25876), .B(n25165), .ZN(n25517) );
  XNOR2_X1 U12416 ( .A(n25517), .B(n25056), .ZN(n24624) );
  NAND2_X1 U12420 ( .A1(n5142), .A2(n21481), .ZN(n5140) );
  NAND3_X1 U12421 ( .A1(n21575), .A2(n20749), .A3(n21580), .ZN(n5141) );
  INV_X1 U12422 ( .A(n20749), .ZN(n21576) );
  INV_X1 U12423 ( .A(n21483), .ZN(n21484) );
  MUX2_X1 U12424 ( .A(n10696), .B(n10984), .S(n10989), .Z(n10584) );
  NAND2_X1 U12425 ( .A1(n23629), .A2(n23308), .ZN(n5143) );
  XNOR2_X1 U12428 ( .A(n5146), .B(n28327), .ZN(n24703) );
  NAND2_X1 U12430 ( .A1(n11152), .A2(n5150), .ZN(n10554) );
  AOI22_X1 U12431 ( .A1(n593), .A2(n11153), .B1(n11154), .B2(n5150), .ZN(
        n10093) );
  NAND2_X1 U12432 ( .A1(n22401), .A2(n5151), .ZN(n21018) );
  NOR2_X1 U12433 ( .A1(n22401), .A2(n5151), .ZN(n21067) );
  NAND3_X1 U12434 ( .A1(n21665), .A2(n21429), .A3(n5151), .ZN(n21017) );
  NAND2_X1 U12438 ( .A1(n28802), .A2(n15334), .ZN(n14781) );
  MUX2_X1 U12440 ( .A(n15047), .B(n15233), .S(n28802), .Z(n15051) );
  NAND2_X1 U12442 ( .A1(n18213), .A2(n18216), .ZN(n5155) );
  NAND2_X1 U12443 ( .A1(n5157), .A2(n28763), .ZN(n18219) );
  INV_X1 U12445 ( .A(n9045), .ZN(n9235) );
  OAI21_X1 U12446 ( .B1(n6590), .B2(n5159), .A(n5158), .ZN(n9240) );
  INV_X1 U12447 ( .A(n9230), .ZN(n5160) );
  XNOR2_X1 U12448 ( .A(n19315), .B(n19314), .ZN(n19319) );
  AND3_X2 U12450 ( .A1(n17886), .A2(n17885), .A3(n17884), .ZN(n19718) );
  INV_X1 U12451 ( .A(n19718), .ZN(n18937) );
  NAND2_X1 U12452 ( .A1(n17887), .A2(n18334), .ZN(n5163) );
  INV_X1 U12453 ( .A(n13661), .ZN(n14044) );
  XNOR2_X1 U12454 ( .A(n5166), .B(n5165), .ZN(n13661) );
  INV_X1 U12455 ( .A(n23924), .ZN(n6321) );
  NAND2_X1 U12456 ( .A1(n5167), .A2(n6746), .ZN(n23924) );
  NAND2_X1 U12457 ( .A1(n5168), .A2(n24612), .ZN(n5167) );
  NAND2_X1 U12458 ( .A1(n11159), .A2(n11158), .ZN(n11783) );
  NAND2_X1 U12459 ( .A1(n11156), .A2(n11155), .ZN(n5171) );
  NAND2_X1 U12460 ( .A1(n11157), .A2(n11154), .ZN(n5172) );
  INV_X1 U12461 ( .A(n23651), .ZN(n23318) );
  INV_X1 U12462 ( .A(n23261), .ZN(n23584) );
  OR2_X2 U12464 ( .A1(n5174), .A2(n5173), .ZN(n9530) );
  XNOR2_X1 U12466 ( .A(n13405), .B(n13461), .ZN(n5177) );
  XNOR2_X1 U12467 ( .A(n13501), .B(n5177), .ZN(n12963) );
  INV_X1 U12468 ( .A(n5177), .ZN(n13131) );
  NAND2_X1 U12469 ( .A1(n5180), .A2(n29611), .ZN(n5344) );
  NAND2_X1 U12470 ( .A1(n5180), .A2(n14304), .ZN(n5343) );
  OAI21_X1 U12472 ( .B1(n20145), .B2(n20148), .A(n5182), .ZN(n5181) );
  OR2_X1 U12473 ( .A1(n21095), .A2(n21092), .ZN(n5182) );
  XNOR2_X1 U12475 ( .A(n22555), .B(n22714), .ZN(n5184) );
  XNOR2_X1 U12476 ( .A(n10135), .B(n10055), .ZN(n5185) );
  INV_X1 U12478 ( .A(n11869), .ZN(n11868) );
  INV_X1 U12480 ( .A(n27771), .ZN(n5188) );
  NAND2_X1 U12481 ( .A1(n15309), .A2(n15310), .ZN(n5190) );
  NOR2_X1 U12486 ( .A1(n11501), .A2(n11874), .ZN(n6305) );
  XNOR2_X2 U12487 ( .A(n8746), .B(n8745), .ZN(n11176) );
  OAI21_X1 U12489 ( .B1(n23151), .B2(n5237), .A(n23767), .ZN(n5236) );
  XNOR2_X2 U12490 ( .A(n9776), .B(n9775), .ZN(n11235) );
  OR2_X1 U12491 ( .A1(n16922), .A2(n5429), .ZN(n5365) );
  XNOR2_X1 U12492 ( .A(n5996), .B(n9843), .ZN(n8884) );
  XNOR2_X2 U12493 ( .A(n13003), .B(n13004), .ZN(n14278) );
  INV_X1 U12494 ( .A(n6886), .ZN(n19510) );
  OAI211_X2 U12495 ( .C1(n28666), .C2(n15084), .A(n14672), .B(n14671), .ZN(
        n16641) );
  XNOR2_X1 U12496 ( .A(n19597), .B(n6193), .ZN(n19344) );
  INV_X1 U12497 ( .A(n15056), .ZN(n6207) );
  XNOR2_X1 U12498 ( .A(n16397), .B(n13926), .ZN(n6707) );
  AOI21_X2 U12499 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(n16603) );
  INV_X1 U12500 ( .A(n27352), .ZN(n5421) );
  OAI21_X2 U12502 ( .B1(n11828), .B2(n11827), .A(n11826), .ZN(n13360) );
  OAI21_X1 U12503 ( .B1(n27771), .B2(n6419), .A(n6418), .ZN(n6498) );
  NOR2_X2 U12507 ( .A1(n14718), .A2(n14717), .ZN(n16422) );
  OAI21_X1 U12508 ( .B1(n6706), .B2(n11622), .A(n6705), .ZN(n11570) );
  OAI21_X1 U12509 ( .B1(n17451), .B2(n28801), .A(n17128), .ZN(n17069) );
  INV_X1 U12511 ( .A(n29044), .ZN(n18187) );
  OAI21_X1 U12516 ( .B1(n23282), .B2(n1893), .A(n23283), .ZN(n5619) );
  XNOR2_X1 U12521 ( .A(n25557), .B(n25933), .ZN(n25559) );
  NAND2_X1 U12522 ( .A1(n5191), .A2(n5149), .ZN(n7602) );
  NAND3_X1 U12523 ( .A1(n7863), .A2(n7092), .A3(n6162), .ZN(n5362) );
  INV_X1 U12526 ( .A(n10079), .ZN(n5195) );
  NAND2_X1 U12528 ( .A1(n15150), .A2(n15151), .ZN(n5199) );
  OAI22_X1 U12529 ( .A1(n21333), .A2(n21332), .B1(n21613), .B2(n21612), .ZN(
        n21336) );
  INV_X1 U12530 ( .A(n21329), .ZN(n20497) );
  INV_X1 U12531 ( .A(n20492), .ZN(n21331) );
  NAND3_X1 U12532 ( .A1(n10739), .A2(n10738), .A3(n5204), .ZN(n12919) );
  NAND2_X1 U12533 ( .A1(n11489), .A2(n11431), .ZN(n5204) );
  NAND2_X1 U12534 ( .A1(n14240), .A2(n29097), .ZN(n13739) );
  NOR2_X1 U12535 ( .A1(n14240), .A2(n29097), .ZN(n14173) );
  OR2_X1 U12536 ( .A1(n14240), .A2(n15194), .ZN(n5207) );
  NAND2_X1 U12537 ( .A1(n19791), .A2(n20481), .ZN(n5208) );
  NAND2_X1 U12538 ( .A1(n18173), .A2(n18172), .ZN(n5209) );
  NAND2_X1 U12539 ( .A1(n24064), .A2(n23897), .ZN(n5210) );
  AOI21_X1 U12540 ( .B1(n28047), .B2(n28069), .A(n5212), .ZN(n5214) );
  AOI21_X1 U12541 ( .B1(n5213), .B2(n28065), .A(n28069), .ZN(n5212) );
  INV_X1 U12542 ( .A(n28065), .ZN(n28071) );
  NAND2_X1 U12543 ( .A1(n28052), .A2(n28067), .ZN(n5215) );
  NAND2_X1 U12544 ( .A1(n5218), .A2(n5216), .ZN(n5289) );
  NAND2_X1 U12545 ( .A1(n5137), .A2(n5217), .ZN(n5216) );
  NAND2_X1 U12547 ( .A1(n22593), .A2(n23829), .ZN(n5219) );
  INV_X1 U12549 ( .A(n26246), .ZN(n5221) );
  AND2_X1 U12550 ( .A1(n18172), .A2(n18174), .ZN(n5222) );
  XNOR2_X1 U12552 ( .A(n19590), .B(n19628), .ZN(n5224) );
  NAND2_X1 U12553 ( .A1(n20495), .A2(n5225), .ZN(n20491) );
  NAND2_X1 U12554 ( .A1(n29616), .A2(n5225), .ZN(n20180) );
  NOR2_X1 U12555 ( .A1(n29616), .A2(n5225), .ZN(n19179) );
  NOR2_X1 U12556 ( .A1(n19863), .A2(n5225), .ZN(n19865) );
  NAND2_X1 U12557 ( .A1(n6834), .A2(n5225), .ZN(n20183) );
  NAND2_X1 U12559 ( .A1(n5229), .A2(n14874), .ZN(n13128) );
  OAI21_X1 U12560 ( .B1(n12053), .B2(n12320), .A(n5230), .ZN(n6679) );
  NAND2_X1 U12561 ( .A1(n12320), .A2(n12051), .ZN(n5230) );
  INV_X1 U12563 ( .A(n18393), .ZN(n17767) );
  NAND2_X1 U12564 ( .A1(n5234), .A2(n17766), .ZN(n5231) );
  OR2_X1 U12565 ( .A1(n17769), .A2(n18388), .ZN(n5235) );
  NAND2_X1 U12566 ( .A1(n15046), .A2(n15225), .ZN(n15353) );
  INV_X1 U12567 ( .A(n7116), .ZN(n7340) );
  NAND2_X1 U12569 ( .A1(n7118), .A2(n5240), .ZN(n5239) );
  NAND2_X1 U12570 ( .A1(n5241), .A2(n7767), .ZN(n5240) );
  NAND2_X1 U12571 ( .A1(n7116), .A2(n5242), .ZN(n5241) );
  NAND2_X1 U12572 ( .A1(n5244), .A2(n7164), .ZN(n5243) );
  XNOR2_X1 U12573 ( .A(n5245), .B(n18799), .ZN(n19290) );
  NAND2_X1 U12575 ( .A1(n28506), .A2(n23800), .ZN(n23538) );
  OAI21_X1 U12576 ( .B1(n23172), .B2(n23540), .A(n28506), .ZN(n23173) );
  NAND2_X1 U12577 ( .A1(n20417), .A2(n20578), .ZN(n6508) );
  AND2_X1 U12578 ( .A1(n5248), .A2(n24768), .ZN(n23548) );
  INV_X1 U12579 ( .A(n24697), .ZN(n5248) );
  NAND2_X1 U12581 ( .A1(n6830), .A2(n5251), .ZN(n5250) );
  NAND2_X1 U12582 ( .A1(n11812), .A2(n12231), .ZN(n5488) );
  OAI22_X1 U12583 ( .A1(n21590), .A2(n21591), .B1(n5684), .B2(n21589), .ZN(
        n21592) );
  NAND3_X1 U12586 ( .A1(n386), .A2(n20275), .A3(n20597), .ZN(n5253) );
  XNOR2_X2 U12587 ( .A(n7047), .B(Key[161]), .ZN(n7967) );
  NAND2_X1 U12588 ( .A1(n7967), .A2(n29300), .ZN(n7962) );
  OAI21_X2 U12589 ( .B1(n10578), .B2(n5258), .A(n5257), .ZN(n12428) );
  NAND3_X1 U12590 ( .A1(n11092), .A2(n10577), .A3(n5258), .ZN(n5257) );
  OAI21_X1 U12591 ( .B1(n17192), .B2(n17347), .A(n5259), .ZN(n5260) );
  NAND2_X1 U12592 ( .A1(n17192), .A2(n17346), .ZN(n5259) );
  NAND2_X1 U12593 ( .A1(n14146), .A2(n13725), .ZN(n5261) );
  OAI21_X1 U12594 ( .B1(n29059), .B2(n13725), .A(n5261), .ZN(n13593) );
  NOR2_X1 U12595 ( .A1(n28521), .A2(n5263), .ZN(n27075) );
  NAND2_X1 U12596 ( .A1(n28521), .A2(n5263), .ZN(n26862) );
  INV_X1 U12597 ( .A(n10973), .ZN(n5265) );
  INV_X1 U12598 ( .A(n10972), .ZN(n10681) );
  NOR2_X1 U12600 ( .A1(n5267), .A2(n10970), .ZN(n5266) );
  XNOR2_X2 U12601 ( .A(n5268), .B(n9297), .ZN(n10970) );
  INV_X1 U12602 ( .A(n337), .ZN(n17309) );
  NAND2_X1 U12603 ( .A1(n15307), .A2(n15311), .ZN(n15272) );
  NAND2_X1 U12606 ( .A1(n1921), .A2(n29569), .ZN(n20888) );
  OAI21_X1 U12607 ( .B1(n5728), .B2(n24079), .A(n5272), .ZN(n5307) );
  OAI22_X1 U12608 ( .A1(n20230), .A2(n4557), .B1(n20353), .B2(n20475), .ZN(
        n21437) );
  XNOR2_X1 U12609 ( .A(n5275), .B(n25869), .ZN(n25215) );
  XNOR2_X1 U12610 ( .A(n25868), .B(n5275), .ZN(n25145) );
  XNOR2_X1 U12611 ( .A(n5275), .B(n25922), .ZN(n25923) );
  XNOR2_X1 U12612 ( .A(n5275), .B(n2523), .ZN(n24137) );
  XNOR2_X1 U12613 ( .A(n26095), .B(n5275), .ZN(n25475) );
  NAND3_X1 U12614 ( .A1(n7340), .A2(n7770), .A3(n7320), .ZN(n5282) );
  NAND2_X1 U12615 ( .A1(n2017), .A2(n5956), .ZN(n5284) );
  MUX2_X1 U12616 ( .A(n14300), .B(n28478), .S(n14299), .Z(n5285) );
  INV_X1 U12617 ( .A(n15069), .ZN(n5287) );
  NAND3_X1 U12619 ( .A1(n16962), .A2(n17309), .A3(n17440), .ZN(n5288) );
  NAND2_X1 U12621 ( .A1(n23078), .A2(n28460), .ZN(n23283) );
  NAND2_X1 U12622 ( .A1(n23839), .A2(n23390), .ZN(n5291) );
  OR2_X1 U12623 ( .A1(n29536), .A2(n29497), .ZN(n5297) );
  NAND2_X1 U12624 ( .A1(n5295), .A2(n5294), .ZN(n27856) );
  NAND2_X1 U12626 ( .A1(n27902), .A2(n29575), .ZN(n5301) );
  NAND2_X1 U12627 ( .A1(n5304), .A2(n5303), .ZN(n5302) );
  MUX2_X1 U12628 ( .A(n20182), .B(n20493), .S(n20495), .Z(n5304) );
  INV_X1 U12629 ( .A(n17313), .ZN(n17317) );
  NAND2_X1 U12630 ( .A1(n13060), .A2(n14354), .ZN(n14356) );
  NAND2_X1 U12631 ( .A1(n13060), .A2(n13824), .ZN(n14349) );
  NAND3_X1 U12632 ( .A1(n4088), .A2(n13060), .A3(n14351), .ZN(n14128) );
  NAND2_X1 U12633 ( .A1(n13825), .A2(n13060), .ZN(n13627) );
  INV_X2 U12635 ( .A(n5306), .ZN(n27076) );
  NAND2_X1 U12636 ( .A1(n26178), .A2(n26177), .ZN(n6125) );
  OAI22_X1 U12637 ( .A1(n6947), .A2(n26447), .B1(n26452), .B2(n26179), .ZN(
        n26178) );
  AOI21_X1 U12638 ( .B1(n6828), .B2(n8643), .A(n9396), .ZN(n5308) );
  NAND2_X1 U12639 ( .A1(n436), .A2(n8981), .ZN(n6828) );
  NAND2_X1 U12640 ( .A1(n409), .A2(n23405), .ZN(n5310) );
  NAND2_X1 U12643 ( .A1(n27209), .A2(n446), .ZN(n5312) );
  NAND2_X1 U12644 ( .A1(n5313), .A2(n295), .ZN(n27212) );
  INV_X1 U12645 ( .A(n27208), .ZN(n5313) );
  OAI21_X1 U12646 ( .B1(n12049), .B2(n12050), .A(n5315), .ZN(n11770) );
  NAND2_X1 U12647 ( .A1(n12049), .A2(n12320), .ZN(n5315) );
  NAND2_X1 U12648 ( .A1(n10490), .A2(n29627), .ZN(n10098) );
  NAND2_X1 U12649 ( .A1(n10549), .A2(n29627), .ZN(n10548) );
  AOI21_X1 U12650 ( .B1(n11114), .B2(n11115), .A(n29627), .ZN(n6250) );
  OAI211_X2 U12651 ( .C1(n1881), .C2(n20631), .A(n20629), .B(n5317), .ZN(
        n21601) );
  NAND2_X1 U12652 ( .A1(n5318), .A2(n28186), .ZN(n5317) );
  NAND2_X1 U12653 ( .A1(n5322), .A2(n5321), .ZN(n5320) );
  NAND2_X1 U12654 ( .A1(n23254), .A2(n28796), .ZN(n5321) );
  AND2_X1 U12655 ( .A1(n11685), .A2(n11996), .ZN(n5323) );
  OAI21_X2 U12657 ( .B1(n5323), .B2(n11757), .A(n11687), .ZN(n12686) );
  OAI21_X2 U12658 ( .B1(n5328), .B2(n18521), .A(n5324), .ZN(n19577) );
  NAND3_X1 U12659 ( .A1(n27287), .A2(n27282), .A3(n27286), .ZN(n5331) );
  MUX2_X1 U12660 ( .A(n5332), .B(n24558), .S(n25794), .Z(n24563) );
  NAND2_X1 U12661 ( .A1(n20577), .A2(n20413), .ZN(n5334) );
  OAI211_X1 U12662 ( .C1(n5336), .C2(n5335), .A(n27103), .B(n27104), .ZN(n5337) );
  XNOR2_X1 U12663 ( .A(n5337), .B(n27105), .ZN(Ciphertext[134]) );
  OAI21_X2 U12664 ( .B1(n21628), .B2(n22141), .A(n5338), .ZN(n22606) );
  NAND3_X1 U12666 ( .A1(n5344), .A2(n5343), .A3(n14302), .ZN(n5342) );
  OAI21_X1 U12667 ( .B1(n23603), .B2(n23247), .A(n5347), .ZN(n5346) );
  NAND2_X1 U12668 ( .A1(n21512), .A2(n21530), .ZN(n21515) );
  NOR2_X1 U12669 ( .A1(n14278), .A2(n14362), .ZN(n5352) );
  NAND2_X1 U12670 ( .A1(n5355), .A2(n23329), .ZN(n5353) );
  NAND2_X1 U12671 ( .A1(n5358), .A2(n5356), .ZN(n21432) );
  NAND2_X1 U12672 ( .A1(n5357), .A2(n4569), .ZN(n5356) );
  NOR2_X1 U12674 ( .A1(n6507), .A2(n29541), .ZN(n26496) );
  INV_X1 U12676 ( .A(n7871), .ZN(n5360) );
  NAND3_X1 U12677 ( .A1(n5362), .A2(n7866), .A3(n5361), .ZN(n8499) );
  OAI21_X1 U12679 ( .B1(n8656), .B2(n8116), .A(n8500), .ZN(n8117) );
  NAND2_X1 U12680 ( .A1(n7880), .A2(n5364), .ZN(n5363) );
  OAI21_X1 U12681 ( .B1(n7879), .B2(n7999), .A(n7878), .ZN(n5364) );
  XNOR2_X1 U12682 ( .A(n19568), .B(n1246), .ZN(n19569) );
  OR2_X1 U12683 ( .A1(n10467), .A2(n5366), .ZN(n6885) );
  AND2_X1 U12684 ( .A1(n5377), .A2(n20644), .ZN(n20646) );
  NAND3_X1 U12685 ( .A1(n5368), .A2(n27497), .A3(n29523), .ZN(n5367) );
  INV_X1 U12686 ( .A(n27492), .ZN(n5368) );
  INV_X1 U12687 ( .A(n27497), .ZN(n27480) );
  NAND2_X1 U12688 ( .A1(n29522), .A2(n27496), .ZN(n5369) );
  OAI22_X1 U12689 ( .A1(n6706), .A2(n11194), .B1(n6687), .B2(n11622), .ZN(
        n5370) );
  NAND2_X1 U12690 ( .A1(n5603), .A2(n11953), .ZN(n5371) );
  NAND2_X1 U12691 ( .A1(n8320), .A2(n9531), .ZN(n8576) );
  OAI21_X1 U12692 ( .B1(n8320), .B2(n8610), .A(n9529), .ZN(n8611) );
  OAI21_X1 U12693 ( .B1(n29662), .B2(n8320), .A(n8747), .ZN(n8748) );
  NAND2_X1 U12694 ( .A1(n27038), .A2(n27213), .ZN(n5372) );
  NAND2_X1 U12695 ( .A1(n20452), .A2(n5377), .ZN(n5376) );
  AOI21_X1 U12696 ( .B1(n14394), .B2(n5378), .A(n14193), .ZN(n12846) );
  MUX2_X1 U12698 ( .A(n15423), .B(n15101), .S(n15102), .Z(n5382) );
  AND2_X2 U12699 ( .A1(n12805), .A2(n12804), .ZN(n15102) );
  INV_X1 U12700 ( .A(n18379), .ZN(n17647) );
  OAI21_X2 U12701 ( .B1(n17154), .B2(n17153), .A(n17152), .ZN(n18379) );
  NOR2_X1 U12702 ( .A1(n28791), .A2(n21326), .ZN(n20907) );
  NAND3_X1 U12703 ( .A1(n13907), .A2(n13906), .A3(n14051), .ZN(n5386) );
  NAND3_X1 U12704 ( .A1(n23487), .A2(n6424), .A3(n23776), .ZN(n5387) );
  XNOR2_X1 U12706 ( .A(n19124), .B(n5393), .ZN(n19128) );
  XNOR2_X1 U12707 ( .A(n19123), .B(n19122), .ZN(n5393) );
  INV_X1 U12709 ( .A(n8608), .ZN(n5396) );
  NAND2_X1 U12710 ( .A1(n17548), .A2(n5398), .ZN(n5397) );
  XNOR2_X1 U12711 ( .A(n10393), .B(n10081), .ZN(n5401) );
  NAND2_X1 U12712 ( .A1(n23694), .A2(n5402), .ZN(n6441) );
  NAND2_X1 U12713 ( .A1(n29059), .A2(n14146), .ZN(n5405) );
  NAND2_X1 U12715 ( .A1(n13958), .A2(n5409), .ZN(n13961) );
  NAND2_X1 U12716 ( .A1(n562), .A2(n14433), .ZN(n5409) );
  XNOR2_X1 U12717 ( .A(n5416), .B(n1046), .ZN(n19543) );
  XNOR2_X1 U12718 ( .A(n5416), .B(n891), .ZN(n19003) );
  XNOR2_X1 U12719 ( .A(n5416), .B(n2916), .ZN(n18256) );
  XNOR2_X1 U12720 ( .A(n19403), .B(n5416), .ZN(n19607) );
  OR2_X1 U12721 ( .A1(n18706), .A2(n18404), .ZN(n18405) );
  NAND2_X1 U12722 ( .A1(n6693), .A2(n8819), .ZN(n6692) );
  NAND3_X1 U12723 ( .A1(n17352), .A2(n17351), .A3(n5418), .ZN(n17353) );
  NAND3_X1 U12724 ( .A1(n17348), .A2(n17347), .A3(n5419), .ZN(n5418) );
  NAND2_X1 U12725 ( .A1(n5420), .A2(n17344), .ZN(n5419) );
  AND3_X1 U12727 ( .A1(n5421), .A2(n27358), .A3(n27355), .ZN(n6287) );
  INV_X1 U12728 ( .A(n14362), .ZN(n14359) );
  NAND2_X1 U12729 ( .A1(n27259), .A2(n5425), .ZN(n26881) );
  INV_X1 U12730 ( .A(n27255), .ZN(n5425) );
  AOI22_X1 U12731 ( .A1(n26887), .A2(n5426), .B1(n26885), .B2(n26886), .ZN(
        n26888) );
  NAND2_X1 U12732 ( .A1(n24028), .A2(n6664), .ZN(n5427) );
  NOR2_X1 U12733 ( .A1(n17297), .A2(n17414), .ZN(n16922) );
  NAND2_X1 U12734 ( .A1(n5430), .A2(n3234), .ZN(n5429) );
  XNOR2_X1 U12735 ( .A(n25336), .B(n5431), .ZN(n5433) );
  XNOR2_X1 U12736 ( .A(n25150), .B(n5432), .ZN(n5434) );
  NAND2_X1 U12738 ( .A1(n19807), .A2(n5436), .ZN(n5435) );
  NAND2_X1 U12739 ( .A1(n19806), .A2(n20302), .ZN(n5437) );
  NAND2_X1 U12741 ( .A1(n5234), .A2(n18227), .ZN(n18389) );
  NOR2_X1 U12742 ( .A1(n5234), .A2(n17592), .ZN(n18220) );
  XNOR2_X1 U12743 ( .A(n22334), .B(n22896), .ZN(n22362) );
  AOI21_X1 U12744 ( .B1(n21311), .B2(n21309), .A(n21308), .ZN(n5443) );
  XNOR2_X1 U12745 ( .A(n15828), .B(n16071), .ZN(n6637) );
  OAI21_X2 U12746 ( .B1(n5447), .B2(n15434), .A(n5446), .ZN(n16071) );
  NAND2_X1 U12747 ( .A1(n15894), .A2(n15434), .ZN(n5446) );
  MUX2_X1 U12748 ( .A(n15431), .B(n15432), .S(n14826), .Z(n15895) );
  NOR2_X1 U12749 ( .A1(n23474), .A2(n23762), .ZN(n5448) );
  NAND2_X1 U12750 ( .A1(n2042), .A2(n8354), .ZN(n5449) );
  NAND3_X1 U12751 ( .A1(n5450), .A2(n279), .A3(n11272), .ZN(n10842) );
  MUX2_X1 U12752 ( .A(n279), .B(n10523), .S(n5450), .Z(n9555) );
  INV_X1 U12753 ( .A(n11275), .ZN(n5450) );
  MUX2_X1 U12754 ( .A(n29131), .B(n23762), .S(n23761), .Z(n23328) );
  NAND3_X1 U12755 ( .A1(n4617), .A2(n11969), .A3(n12156), .ZN(n11973) );
  NAND2_X1 U12756 ( .A1(n12241), .A2(n4617), .ZN(n11514) );
  NOR2_X1 U12757 ( .A1(n5839), .A2(n4617), .ZN(n10862) );
  NAND2_X1 U12758 ( .A1(n5693), .A2(n14452), .ZN(n5451) );
  XNOR2_X1 U12760 ( .A(n22461), .B(n21856), .ZN(n5453) );
  INV_X1 U12761 ( .A(n24602), .ZN(n24738) );
  NAND2_X1 U12763 ( .A1(n22355), .A2(n22354), .ZN(n5456) );
  NAND2_X1 U12764 ( .A1(n22310), .A2(n23636), .ZN(n5457) );
  AND2_X1 U12765 ( .A1(n29566), .A2(n17435), .ZN(n5460) );
  NAND2_X1 U12766 ( .A1(n5461), .A2(n17440), .ZN(n5459) );
  AND2_X1 U12767 ( .A1(n336), .A2(n17439), .ZN(n5461) );
  INV_X1 U12768 ( .A(n21306), .ZN(n21307) );
  NAND2_X1 U12769 ( .A1(n20768), .A2(n29530), .ZN(n20774) );
  XNOR2_X1 U12770 ( .A(n13054), .B(n5463), .ZN(n12551) );
  NAND2_X1 U12771 ( .A1(n12239), .A2(n5839), .ZN(n5462) );
  NAND2_X1 U12772 ( .A1(n11612), .A2(n11613), .ZN(n5464) );
  NAND2_X1 U12773 ( .A1(n12316), .A2(n12049), .ZN(n11612) );
  INV_X1 U12774 ( .A(n13054), .ZN(n12790) );
  OAI21_X1 U12775 ( .B1(n12028), .B2(n5466), .A(n12026), .ZN(n5467) );
  NAND2_X1 U12776 ( .A1(n10489), .A2(n431), .ZN(n5468) );
  NAND2_X1 U12777 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  NAND2_X1 U12778 ( .A1(n18130), .A2(n18591), .ZN(n5472) );
  NAND3_X1 U12779 ( .A1(n5475), .A2(n17835), .A3(n18129), .ZN(n5473) );
  OAI21_X2 U12780 ( .B1(n5476), .B2(n17632), .A(n5474), .ZN(n19256) );
  NAND2_X1 U12781 ( .A1(n17835), .A2(n18589), .ZN(n17632) );
  NAND2_X1 U12783 ( .A1(n24814), .A2(n24809), .ZN(n5478) );
  OAI21_X2 U12784 ( .B1(n14052), .B2(n14051), .A(n14050), .ZN(n14695) );
  NAND2_X1 U12785 ( .A1(n7869), .A2(n5483), .ZN(n7959) );
  NAND3_X1 U12787 ( .A1(n5486), .A2(n5484), .A3(n29585), .ZN(n5485) );
  NAND2_X1 U12788 ( .A1(n27193), .A2(n27124), .ZN(n5484) );
  OAI211_X1 U12789 ( .C1(n17394), .C2(n17393), .A(n5487), .B(n17400), .ZN(
        n17399) );
  NAND3_X2 U12790 ( .A1(n11530), .A2(n11531), .A3(n5488), .ZN(n13533) );
  NAND3_X1 U12791 ( .A1(n12230), .A2(n12229), .A3(n5489), .ZN(n13448) );
  NAND2_X1 U12792 ( .A1(n11812), .A2(n13087), .ZN(n5489) );
  NAND2_X1 U12794 ( .A1(n18043), .A2(n18042), .ZN(n5496) );
  OAI21_X1 U12796 ( .B1(n27025), .B2(n28592), .A(n5497), .ZN(n5498) );
  NAND2_X1 U12797 ( .A1(n393), .A2(n27029), .ZN(n5497) );
  NAND2_X1 U12798 ( .A1(n5501), .A2(n5499), .ZN(n26593) );
  NAND2_X1 U12799 ( .A1(n5500), .A2(n306), .ZN(n5499) );
  MUX2_X1 U12800 ( .A(n29588), .B(n27032), .S(n27025), .Z(n5500) );
  NAND2_X1 U12801 ( .A1(n24576), .A2(n28482), .ZN(n5502) );
  NAND2_X1 U12802 ( .A1(n26933), .A2(n5505), .ZN(n26166) );
  INV_X1 U12803 ( .A(n26579), .ZN(n5505) );
  INV_X1 U12805 ( .A(n26581), .ZN(n26930) );
  INV_X1 U12806 ( .A(n24916), .ZN(n5873) );
  NAND2_X1 U12807 ( .A1(n5511), .A2(n5512), .ZN(n5507) );
  XNOR2_X1 U12808 ( .A(n5873), .B(n26083), .ZN(n24753) );
  NAND3_X1 U12809 ( .A1(n24550), .A2(n5509), .A3(n22869), .ZN(n5508) );
  NAND2_X1 U12810 ( .A1(n24554), .A2(n24555), .ZN(n5510) );
  NAND2_X1 U12811 ( .A1(n24052), .A2(n24468), .ZN(n5511) );
  NAND2_X1 U12812 ( .A1(n24467), .A2(n24053), .ZN(n5512) );
  INV_X1 U12813 ( .A(n12891), .ZN(n5514) );
  OAI21_X1 U12814 ( .B1(n15209), .B2(n14960), .A(n5515), .ZN(n14927) );
  NAND2_X1 U12815 ( .A1(n11608), .A2(n4197), .ZN(n11492) );
  NAND2_X1 U12816 ( .A1(n18397), .A2(n18396), .ZN(n18403) );
  NAND2_X1 U12817 ( .A1(n18232), .A2(n17977), .ZN(n18396) );
  NAND2_X1 U12818 ( .A1(n17407), .A2(n423), .ZN(n5517) );
  NAND2_X1 U12819 ( .A1(n17408), .A2(n17570), .ZN(n5518) );
  AND2_X2 U12820 ( .A1(n6765), .A2(n6900), .ZN(n18232) );
  INV_X1 U12821 ( .A(n14494), .ZN(n14154) );
  NAND3_X1 U12823 ( .A1(n14154), .A2(n14498), .A3(n14493), .ZN(n5519) );
  XNOR2_X1 U12824 ( .A(n18802), .B(n1248), .ZN(n5521) );
  XNOR2_X1 U12825 ( .A(n18761), .B(n5759), .ZN(n5522) );
  XNOR2_X1 U12826 ( .A(n18409), .B(n18987), .ZN(n5523) );
  NAND2_X1 U12827 ( .A1(n11599), .A2(n12202), .ZN(n5526) );
  NOR2_X1 U12828 ( .A1(n10988), .A2(n10983), .ZN(n10697) );
  NAND2_X1 U12829 ( .A1(n10630), .A2(n10983), .ZN(n10634) );
  OAI21_X1 U12830 ( .B1(n16888), .B2(n17143), .A(n5527), .ZN(n16228) );
  NAND2_X1 U12831 ( .A1(n17143), .A2(n17137), .ZN(n5527) );
  NAND2_X1 U12833 ( .A1(n5408), .A2(n383), .ZN(n5529) );
  XNOR2_X2 U12834 ( .A(n13321), .B(n13320), .ZN(n5531) );
  NAND3_X1 U12835 ( .A1(n13910), .A2(n13729), .A3(n5531), .ZN(n5886) );
  NOR2_X1 U12836 ( .A1(n28171), .A2(n5531), .ZN(n13915) );
  NAND3_X1 U12837 ( .A1(n3798), .A2(n13730), .A3(n5531), .ZN(n6352) );
  AOI21_X1 U12838 ( .B1(n13643), .B2(n13912), .A(n5531), .ZN(n13644) );
  NAND2_X1 U12839 ( .A1(n5534), .A2(n11190), .ZN(n5532) );
  NAND3_X1 U12840 ( .A1(n11191), .A2(n11355), .A3(n11352), .ZN(n5533) );
  NAND2_X1 U12841 ( .A1(n11355), .A2(n11351), .ZN(n5534) );
  NOR2_X1 U12842 ( .A1(n18172), .A2(n18168), .ZN(n5535) );
  XNOR2_X1 U12844 ( .A(n19590), .B(n19269), .ZN(n5539) );
  XNOR2_X1 U12845 ( .A(n19591), .B(n19593), .ZN(n5538) );
  INV_X1 U12846 ( .A(n17255), .ZN(n17251) );
  NAND2_X1 U12850 ( .A1(n12399), .A2(n14411), .ZN(n5542) );
  XNOR2_X1 U12851 ( .A(n13447), .B(n13227), .ZN(n12834) );
  OAI22_X1 U12852 ( .A1(n5544), .A2(n28155), .B1(n21563), .B2(n21560), .ZN(
        n20757) );
  NAND2_X1 U12853 ( .A1(n20418), .A2(n5545), .ZN(n20419) );
  OAI22_X1 U12854 ( .A1(n25152), .A2(n5546), .B1(n26936), .B2(n26944), .ZN(
        n25159) );
  NAND2_X1 U12855 ( .A1(n23420), .A2(n483), .ZN(n5547) );
  NAND2_X1 U12856 ( .A1(n29507), .A2(n17802), .ZN(n18426) );
  INV_X1 U12857 ( .A(n5551), .ZN(n5550) );
  NAND2_X1 U12859 ( .A1(n23625), .A2(n23624), .ZN(n5554) );
  NAND2_X1 U12860 ( .A1(n23623), .A2(n23622), .ZN(n5556) );
  OR2_X1 U12861 ( .A1(n17298), .A2(n3234), .ZN(n5557) );
  NAND2_X1 U12862 ( .A1(n7885), .A2(n7886), .ZN(n5559) );
  NAND2_X1 U12863 ( .A1(n28479), .A2(n21091), .ZN(n5560) );
  NAND2_X1 U12865 ( .A1(n17933), .A2(n18480), .ZN(n5561) );
  XNOR2_X1 U12867 ( .A(n22705), .B(n27534), .ZN(n22769) );
  NAND2_X1 U12868 ( .A1(n20985), .A2(n19013), .ZN(n5564) );
  NAND2_X1 U12869 ( .A1(n20913), .A2(n19014), .ZN(n5565) );
  XNOR2_X1 U12870 ( .A(n15893), .B(n14523), .ZN(n5566) );
  INV_X1 U12871 ( .A(n9045), .ZN(n5568) );
  INV_X1 U12872 ( .A(n9233), .ZN(n5567) );
  NOR2_X1 U12873 ( .A1(n9235), .A2(n9233), .ZN(n5569) );
  OAI21_X1 U12874 ( .B1(n9233), .B2(n5945), .A(n5570), .ZN(n7001) );
  NAND2_X1 U12875 ( .A1(n5160), .A2(n5945), .ZN(n5570) );
  INV_X1 U12876 ( .A(n24704), .ZN(n24708) );
  OAI211_X1 U12877 ( .C1(n592), .C2(n28405), .A(n5574), .B(n5573), .ZN(n5572)
         );
  NAND2_X1 U12878 ( .A1(n592), .A2(n10936), .ZN(n5574) );
  OAI21_X1 U12879 ( .B1(n14622), .B2(n15500), .A(n5577), .ZN(n5576) );
  AND2_X1 U12880 ( .A1(n14705), .A2(n15498), .ZN(n14622) );
  NAND2_X1 U12881 ( .A1(n12236), .A2(n375), .ZN(n5578) );
  NAND2_X1 U12882 ( .A1(n1986), .A2(n12236), .ZN(n5579) );
  INV_X1 U12883 ( .A(n294), .ZN(n5581) );
  NAND2_X1 U12884 ( .A1(n11077), .A2(n11076), .ZN(n10663) );
  INV_X1 U12885 ( .A(n11294), .ZN(n11077) );
  NAND2_X1 U12886 ( .A1(n1830), .A2(n5584), .ZN(n13815) );
  NAND2_X1 U12887 ( .A1(n13880), .A2(n5584), .ZN(n13883) );
  NAND2_X1 U12888 ( .A1(n16722), .A2(n16803), .ZN(n5585) );
  NAND2_X1 U12889 ( .A1(n16725), .A2(n3883), .ZN(n16802) );
  NAND2_X1 U12891 ( .A1(n11335), .A2(n11176), .ZN(n11175) );
  NAND2_X1 U12894 ( .A1(n6849), .A2(n5590), .ZN(n6848) );
  NAND3_X1 U12895 ( .A1(n571), .A2(n6687), .A3(n5838), .ZN(n5590) );
  INV_X1 U12896 ( .A(n14972), .ZN(n14583) );
  NOR2_X1 U12897 ( .A1(n8575), .A2(n5594), .ZN(n9420) );
  MUX2_X1 U12898 ( .A(n606), .B(n5594), .S(n7569), .Z(n8582) );
  NAND3_X1 U12899 ( .A1(n5129), .A2(n5594), .A3(n603), .ZN(n8768) );
  OAI21_X1 U12900 ( .B1(n5129), .B2(n5594), .A(n5592), .ZN(n9422) );
  OAI21_X1 U12901 ( .B1(n8327), .B2(n606), .A(n9425), .ZN(n5593) );
  NAND2_X1 U12903 ( .A1(n11184), .A2(n29316), .ZN(n11185) );
  OAI211_X1 U12904 ( .C1(n11321), .C2(n29316), .A(n10473), .B(n11183), .ZN(
        n10475) );
  MUX2_X1 U12906 ( .A(n15167), .B(n15166), .S(n15165), .Z(n5597) );
  NAND2_X1 U12907 ( .A1(n15169), .A2(n15168), .ZN(n5599) );
  NOR2_X1 U12908 ( .A1(n27409), .A2(n1175), .ZN(n5601) );
  INV_X1 U12909 ( .A(n27403), .ZN(n5600) );
  NAND2_X1 U12910 ( .A1(n5601), .A2(n5600), .ZN(n25638) );
  NOR2_X1 U12911 ( .A1(n27403), .A2(n27409), .ZN(n5602) );
  NOR2_X1 U12912 ( .A1(n25634), .A2(n5602), .ZN(n25640) );
  XNOR2_X1 U12913 ( .A(n13226), .B(n13451), .ZN(n11629) );
  INV_X1 U12914 ( .A(n27496), .ZN(n5607) );
  INV_X1 U12915 ( .A(n5605), .ZN(n27476) );
  INV_X1 U12916 ( .A(n27494), .ZN(n5604) );
  NAND2_X1 U12917 ( .A1(n5608), .A2(n5607), .ZN(n5606) );
  NOR2_X1 U12918 ( .A1(n29523), .A2(n27497), .ZN(n5608) );
  NAND2_X1 U12919 ( .A1(n16953), .A2(n17359), .ZN(n16714) );
  OAI21_X1 U12920 ( .B1(n23759), .B2(n23760), .A(n23758), .ZN(n5611) );
  XNOR2_X2 U12922 ( .A(n5613), .B(n5612), .ZN(n6114) );
  XNOR2_X1 U12923 ( .A(n18989), .B(n18990), .ZN(n5612) );
  XNOR2_X1 U12924 ( .A(n18987), .B(n18988), .ZN(n5613) );
  NAND2_X1 U12925 ( .A1(n14127), .A2(n5615), .ZN(n14129) );
  NOR2_X1 U12926 ( .A1(n14353), .A2(n14126), .ZN(n5615) );
  NAND2_X1 U12927 ( .A1(n5617), .A2(n14126), .ZN(n5616) );
  INV_X1 U12928 ( .A(n14354), .ZN(n5617) );
  NAND2_X1 U12930 ( .A1(n16601), .A2(n17109), .ZN(n5620) );
  XNOR2_X1 U12931 ( .A(n14983), .B(n5621), .ZN(n14984) );
  XNOR2_X1 U12932 ( .A(n16650), .B(n5621), .ZN(n16651) );
  OAI211_X2 U12933 ( .C1(n24524), .C2(n24525), .A(n24528), .B(n6223), .ZN(
        n25948) );
  OAI21_X2 U12934 ( .B1(n5622), .B2(n20143), .A(n20142), .ZN(n22270) );
  NAND2_X1 U12936 ( .A1(n6656), .A2(n5623), .ZN(n6655) );
  INV_X1 U12937 ( .A(n27433), .ZN(n27441) );
  NAND2_X1 U12939 ( .A1(n437), .A2(n7993), .ZN(n7241) );
  XNOR2_X2 U12940 ( .A(n7056), .B(Key[165]), .ZN(n7993) );
  OAI21_X1 U12941 ( .B1(n23171), .B2(n23516), .A(n23170), .ZN(n5626) );
  AOI21_X1 U12942 ( .B1(n23681), .B2(n5883), .A(n29544), .ZN(n5627) );
  OAI211_X1 U12943 ( .C1(n5632), .C2(n6420), .A(n5631), .B(n5628), .ZN(n5629)
         );
  NAND2_X1 U12944 ( .A1(n6420), .A2(n5633), .ZN(n5628) );
  XNOR2_X1 U12945 ( .A(n25820), .B(n5629), .ZN(n5630) );
  XNOR2_X1 U12946 ( .A(n25071), .B(n5630), .ZN(n25073) );
  NAND2_X1 U12948 ( .A1(n6422), .A2(n5633), .ZN(n5631) );
  XNOR2_X2 U12950 ( .A(n13356), .B(n13357), .ZN(n13914) );
  NAND2_X1 U12951 ( .A1(n5637), .A2(n12512), .ZN(n11837) );
  NAND3_X1 U12953 ( .A1(n15892), .A2(n18299), .A3(n18298), .ZN(n18300) );
  AOI21_X1 U12954 ( .B1(n5645), .B2(n5644), .A(n15494), .ZN(n5640) );
  NAND2_X1 U12956 ( .A1(n22955), .A2(n28484), .ZN(n5646) );
  NAND2_X1 U12957 ( .A1(n22956), .A2(n28183), .ZN(n5647) );
  XNOR2_X1 U12958 ( .A(n5650), .B(n5649), .ZN(Ciphertext[16]) );
  NAND2_X1 U12961 ( .A1(n26612), .A2(n26613), .ZN(n5652) );
  NAND2_X1 U12963 ( .A1(n24729), .A2(n24598), .ZN(n5653) );
  NAND2_X1 U12965 ( .A1(n5656), .A2(n460), .ZN(n5655) );
  NOR2_X1 U12966 ( .A1(n24730), .A2(n24726), .ZN(n5656) );
  NAND2_X1 U12967 ( .A1(n19832), .A2(n5657), .ZN(n21758) );
  MUX2_X1 U12968 ( .A(n20864), .B(n21497), .S(n21493), .Z(n5658) );
  INV_X1 U12969 ( .A(n18344), .ZN(n5659) );
  OAI21_X1 U12970 ( .B1(n11954), .B2(n11580), .A(n5661), .ZN(n5660) );
  AOI22_X1 U12971 ( .A1(n1924), .A2(n21420), .B1(n5664), .B2(n21087), .ZN(
        n5663) );
  NOR2_X1 U12972 ( .A1(n21425), .A2(n21424), .ZN(n5664) );
  NAND2_X1 U12973 ( .A1(n21427), .A2(n28602), .ZN(n5665) );
  NOR2_X1 U12974 ( .A1(n7114), .A2(n8828), .ZN(n7447) );
  INV_X1 U12975 ( .A(n8828), .ZN(n8193) );
  NAND2_X1 U12976 ( .A1(n5667), .A2(n14177), .ZN(n5666) );
  OAI21_X1 U12977 ( .B1(n14451), .B2(n13753), .A(n14450), .ZN(n5667) );
  OR2_X1 U12978 ( .A1(n20181), .A2(n20182), .ZN(n5668) );
  NAND2_X1 U12979 ( .A1(n20163), .A2(n20162), .ZN(n5669) );
  AND2_X1 U12980 ( .A1(n17883), .A2(n18379), .ZN(n5671) );
  NAND2_X1 U12981 ( .A1(n3283), .A2(n5671), .ZN(n17884) );
  NAND2_X1 U12984 ( .A1(n8661), .A2(n8910), .ZN(n5677) );
  NAND2_X1 U12985 ( .A1(n9015), .A2(n8908), .ZN(n8661) );
  INV_X1 U12986 ( .A(n14916), .ZN(n5679) );
  NAND2_X1 U12987 ( .A1(n14500), .A2(n14501), .ZN(n5678) );
  NAND3_X1 U12988 ( .A1(n15488), .A2(n15487), .A3(n5679), .ZN(n15493) );
  NAND2_X1 U12989 ( .A1(n21495), .A2(n21493), .ZN(n21126) );
  NAND2_X1 U12990 ( .A1(n19850), .A2(n19851), .ZN(n5680) );
  NAND3_X1 U12991 ( .A1(n5680), .A2(n20394), .A3(n20560), .ZN(n19853) );
  NAND2_X1 U12992 ( .A1(n14657), .A2(n548), .ZN(n5681) );
  NAND2_X1 U12994 ( .A1(n12977), .A2(n5682), .ZN(n14874) );
  NOR2_X1 U12995 ( .A1(n21322), .A2(n5684), .ZN(n20575) );
  NAND2_X1 U12996 ( .A1(n28584), .A2(n5684), .ZN(n6043) );
  NAND2_X1 U13000 ( .A1(n26625), .A2(n27013), .ZN(n5687) );
  NAND2_X1 U13001 ( .A1(n5691), .A2(n5689), .ZN(n5688) );
  NAND3_X1 U13002 ( .A1(n5690), .A2(n18216), .A3(n18500), .ZN(n5689) );
  INV_X1 U13003 ( .A(n13753), .ZN(n5693) );
  INV_X1 U13004 ( .A(n17543), .ZN(n5695) );
  INV_X1 U13005 ( .A(n17543), .ZN(n17217) );
  XNOR2_X2 U13006 ( .A(n15800), .B(n15799), .ZN(n17540) );
  NAND2_X1 U13007 ( .A1(n22676), .A2(n5699), .ZN(n5698) );
  NAND3_X1 U13008 ( .A1(n18346), .A2(n17948), .A3(n514), .ZN(n5700) );
  XNOR2_X1 U13009 ( .A(n21876), .B(n22809), .ZN(n5702) );
  XNOR2_X1 U13010 ( .A(n21877), .B(n21878), .ZN(n5703) );
  OR2_X1 U13012 ( .A1(n11237), .A2(n11235), .ZN(n5707) );
  XNOR2_X2 U13014 ( .A(n9738), .B(n9739), .ZN(n11237) );
  NAND2_X1 U13015 ( .A1(n23296), .A2(n22864), .ZN(n23298) );
  OAI211_X1 U13019 ( .C1(n12288), .C2(n12289), .A(n3558), .B(n5715), .ZN(
        n12295) );
  XNOR2_X1 U13020 ( .A(n5718), .B(n22501), .ZN(n22503) );
  NAND2_X1 U13022 ( .A1(n5725), .A2(n5726), .ZN(n5723) );
  INV_X1 U13023 ( .A(n15502), .ZN(n5726) );
  NOR2_X1 U13024 ( .A1(n15506), .A2(n15265), .ZN(n5724) );
  NOR2_X1 U13025 ( .A1(n15500), .A2(n15265), .ZN(n5725) );
  INV_X1 U13026 ( .A(n24077), .ZN(n5728) );
  NAND2_X1 U13027 ( .A1(n5729), .A2(n28401), .ZN(n23508) );
  AND2_X1 U13028 ( .A1(n24081), .A2(n24133), .ZN(n5729) );
  NAND3_X1 U13029 ( .A1(n23911), .A2(n24079), .A3(n28401), .ZN(n23912) );
  OAI211_X1 U13030 ( .C1(n14774), .C2(n14775), .A(n14773), .B(n14812), .ZN(
        n14776) );
  NAND2_X1 U13031 ( .A1(n14772), .A2(n14807), .ZN(n14812) );
  INV_X1 U13032 ( .A(n14051), .ZN(n5731) );
  NAND2_X1 U13035 ( .A1(n16538), .A2(n4703), .ZN(n5734) );
  NOR2_X1 U13036 ( .A1(n393), .A2(n306), .ZN(n24826) );
  AOI21_X1 U13037 ( .B1(n393), .B2(n306), .A(n27032), .ZN(n26692) );
  AOI21_X1 U13038 ( .B1(n26691), .B2(n26819), .A(n393), .ZN(n26694) );
  NOR2_X1 U13040 ( .A1(n24823), .A2(n1978), .ZN(n5735) );
  OAI211_X1 U13041 ( .C1(n17078), .C2(n5738), .A(n4655), .B(n5736), .ZN(n5739)
         );
  INV_X1 U13042 ( .A(n17148), .ZN(n5737) );
  INV_X1 U13043 ( .A(n17485), .ZN(n5738) );
  NAND2_X1 U13044 ( .A1(n17490), .A2(n17489), .ZN(n5740) );
  NAND2_X1 U13045 ( .A1(n23759), .A2(n23760), .ZN(n5741) );
  NAND2_X1 U13047 ( .A1(n13953), .A2(n14194), .ZN(n5745) );
  XNOR2_X1 U13048 ( .A(n19520), .B(n5746), .ZN(n18929) );
  AND3_X2 U13049 ( .A1(n5747), .A2(n17594), .A3(n17595), .ZN(n19139) );
  XNOR2_X1 U13050 ( .A(n25440), .B(n25819), .ZN(n25113) );
  NAND2_X1 U13052 ( .A1(n5751), .A2(n5752), .ZN(n5748) );
  NAND2_X1 U13053 ( .A1(n5753), .A2(n11308), .ZN(n5835) );
  MUX2_X1 U13054 ( .A(n11309), .B(n11310), .S(n1933), .Z(n11311) );
  MUX2_X1 U13055 ( .A(n23445), .B(n23442), .S(n23448), .Z(n23111) );
  XNOR2_X1 U13056 ( .A(n24924), .B(n24926), .ZN(n5755) );
  XNOR2_X1 U13058 ( .A(n19289), .B(n19290), .ZN(n19295) );
  NAND2_X1 U13060 ( .A1(n5757), .A2(n18401), .ZN(n5756) );
  NAND2_X1 U13061 ( .A1(n18403), .A2(n18402), .ZN(n5758) );
  OR2_X1 U13062 ( .A1(n5760), .A2(n26748), .ZN(n25644) );
  AND2_X1 U13063 ( .A1(n26748), .A2(n5760), .ZN(n25979) );
  NAND2_X1 U13064 ( .A1(n29099), .A2(n28563), .ZN(n5761) );
  NOR2_X1 U13065 ( .A1(n28583), .A2(n5760), .ZN(n25978) );
  MUX2_X1 U13066 ( .A(n28583), .B(n26224), .S(n28563), .Z(n26225) );
  NAND2_X1 U13071 ( .A1(n7116), .A2(n7320), .ZN(n7768) );
  NAND2_X1 U13072 ( .A1(n7321), .A2(n7116), .ZN(n7322) );
  AOI21_X1 U13073 ( .B1(n7769), .B2(n7116), .A(n614), .ZN(n7325) );
  NAND2_X1 U13074 ( .A1(n24729), .A2(n5767), .ZN(n24290) );
  NAND2_X1 U13075 ( .A1(n460), .A2(n5768), .ZN(n24147) );
  INV_X1 U13076 ( .A(n5769), .ZN(n6310) );
  OAI21_X1 U13077 ( .B1(n5770), .B2(n23492), .A(n23799), .ZN(n5769) );
  OAI22_X1 U13078 ( .A1(n23011), .A2(n23351), .B1(n5773), .B2(n23657), .ZN(
        n23659) );
  INV_X1 U13079 ( .A(n23351), .ZN(n5774) );
  NAND2_X1 U13080 ( .A1(n11377), .A2(n12166), .ZN(n11843) );
  INV_X1 U13081 ( .A(n22284), .ZN(n23628) );
  NAND2_X1 U13082 ( .A1(n23040), .A2(n23309), .ZN(n23041) );
  INV_X1 U13083 ( .A(n23633), .ZN(n5775) );
  OR2_X1 U13084 ( .A1(n27771), .A2(n5776), .ZN(n27775) );
  NAND2_X1 U13085 ( .A1(n15047), .A2(n15238), .ZN(n5777) );
  INV_X1 U13087 ( .A(n20041), .ZN(n5778) );
  NAND2_X1 U13088 ( .A1(n5781), .A2(n20646), .ZN(n5779) );
  XNOR2_X1 U13090 ( .A(n16481), .B(n16479), .ZN(n5784) );
  XNOR2_X1 U13091 ( .A(n16399), .B(n16398), .ZN(n16488) );
  OAI211_X2 U13092 ( .C1(n3362), .C2(n5788), .A(n5786), .B(n5785), .ZN(n16398)
         );
  NAND3_X1 U13093 ( .A1(n3362), .A2(n15407), .A3(n15406), .ZN(n5786) );
  NAND2_X1 U13095 ( .A1(n29312), .A2(n14250), .ZN(n5936) );
  NAND2_X1 U13096 ( .A1(n5789), .A2(n29312), .ZN(n5790) );
  NAND2_X1 U13097 ( .A1(n16491), .A2(n17829), .ZN(n5792) );
  NAND2_X1 U13098 ( .A1(n17073), .A2(n17506), .ZN(n16550) );
  NAND2_X1 U13099 ( .A1(n19768), .A2(n5793), .ZN(n21145) );
  NAND3_X1 U13100 ( .A1(n18919), .A2(n5794), .A3(n20106), .ZN(n5793) );
  NOR2_X1 U13101 ( .A1(n20704), .A2(n20967), .ZN(n20705) );
  NAND2_X1 U13102 ( .A1(n381), .A2(n20972), .ZN(n20704) );
  AND2_X1 U13103 ( .A1(n14697), .A2(n15513), .ZN(n15276) );
  NAND2_X1 U13104 ( .A1(n5168), .A2(n24017), .ZN(n5799) );
  XNOR2_X1 U13105 ( .A(n5801), .B(n21903), .ZN(n22620) );
  INV_X1 U13106 ( .A(n21987), .ZN(n5801) );
  XNOR2_X1 U13107 ( .A(n21903), .B(n5802), .ZN(n22101) );
  INV_X1 U13108 ( .A(n21903), .ZN(n5803) );
  NAND2_X1 U13109 ( .A1(n558), .A2(n14158), .ZN(n14159) );
  NOR2_X1 U13111 ( .A1(n29320), .A2(n14479), .ZN(n5804) );
  NAND2_X1 U13113 ( .A1(n17070), .A2(n17830), .ZN(n17513) );
  NAND2_X1 U13114 ( .A1(n5808), .A2(n17070), .ZN(n5807) );
  NAND2_X1 U13115 ( .A1(n5812), .A2(n5810), .ZN(n13791) );
  INV_X1 U13117 ( .A(n14882), .ZN(n5811) );
  NAND2_X1 U13118 ( .A1(n13790), .A2(n5813), .ZN(n5812) );
  NAND2_X1 U13119 ( .A1(n1896), .A2(n14044), .ZN(n6010) );
  NOR2_X1 U13120 ( .A1(n28626), .A2(n23416), .ZN(n22928) );
  MUX2_X1 U13121 ( .A(n23417), .B(n28626), .S(n23416), .Z(n6091) );
  MUX2_X1 U13122 ( .A(n23419), .B(n28626), .S(n5856), .Z(n22808) );
  XNOR2_X1 U13123 ( .A(n22459), .B(n22123), .ZN(n20923) );
  OAI21_X1 U13126 ( .B1(n20802), .B2(n5817), .A(n20801), .ZN(n20803) );
  OAI21_X1 U13127 ( .B1(n20955), .B2(n29586), .A(n5816), .ZN(n21101) );
  NAND2_X1 U13128 ( .A1(n21930), .A2(n21099), .ZN(n5816) );
  OR2_X1 U13129 ( .A1(n21934), .A2(n5817), .ZN(n6345) );
  XOR2_X1 U13131 ( .A(n10087), .B(n10426), .Z(n5818) );
  AND2_X1 U13132 ( .A1(n8117), .A2(n8502), .ZN(n5819) );
  NAND2_X1 U13134 ( .A1(n13757), .A2(n14158), .ZN(n5822) );
  NAND2_X1 U13135 ( .A1(n14162), .A2(n13756), .ZN(n5823) );
  NAND2_X1 U13136 ( .A1(n14474), .A2(n13754), .ZN(n14162) );
  XNOR2_X1 U13137 ( .A(n9924), .B(n5824), .ZN(n8520) );
  INV_X1 U13138 ( .A(n5824), .ZN(n10320) );
  XNOR2_X1 U13139 ( .A(n10250), .B(n10386), .ZN(n5824) );
  NAND2_X1 U13140 ( .A1(n5825), .A2(n12203), .ZN(n6073) );
  NAND2_X1 U13141 ( .A1(n20587), .A2(n20584), .ZN(n6914) );
  NAND2_X1 U13144 ( .A1(n5827), .A2(n21424), .ZN(n21422) );
  NAND2_X1 U13145 ( .A1(n5827), .A2(n20899), .ZN(n20804) );
  NOR2_X1 U13146 ( .A1(n21425), .A2(n5827), .ZN(n20140) );
  INV_X1 U13147 ( .A(n16588), .ZN(n5828) );
  NAND3_X1 U13149 ( .A1(n5832), .A2(n25405), .A3(n5831), .ZN(n26708) );
  NAND2_X1 U13150 ( .A1(n26463), .A2(n26469), .ZN(n5832) );
  NAND2_X1 U13151 ( .A1(n25008), .A2(n25005), .ZN(n24305) );
  NOR2_X1 U13152 ( .A1(n388), .A2(n14882), .ZN(n6061) );
  NAND2_X1 U13154 ( .A1(n24338), .A2(n24341), .ZN(n24128) );
  NAND3_X1 U13155 ( .A1(n24708), .A2(n24338), .A3(n24707), .ZN(n24342) );
  OAI21_X1 U13156 ( .B1(n6611), .B2(n24338), .A(n5836), .ZN(n25543) );
  XNOR2_X1 U13157 ( .A(n5841), .B(n5840), .ZN(n22283) );
  NAND2_X1 U13158 ( .A1(n16615), .A2(n5844), .ZN(n5843) );
  NAND2_X1 U13159 ( .A1(n518), .A2(n18356), .ZN(n5844) );
  NAND2_X1 U13160 ( .A1(n5847), .A2(n5846), .ZN(n5845) );
  NOR2_X1 U13161 ( .A1(n13912), .A2(n13914), .ZN(n5846) );
  NAND2_X1 U13162 ( .A1(n13914), .A2(n13915), .ZN(n5848) );
  XNOR2_X1 U13163 ( .A(n5849), .B(n26409), .ZN(Ciphertext[178]) );
  OAI211_X1 U13164 ( .C1(n26408), .C2(n29031), .A(n5851), .B(n5850), .ZN(n5849) );
  OAI21_X1 U13165 ( .B1(n5852), .B2(n28040), .A(n6859), .ZN(n5851) );
  AND2_X1 U13166 ( .A1(n28024), .A2(n28027), .ZN(n28040) );
  AND2_X1 U13167 ( .A1(n28025), .A2(n29031), .ZN(n5852) );
  NOR2_X1 U13168 ( .A1(n21213), .A2(n21211), .ZN(n5855) );
  MUX2_X1 U13169 ( .A(n25750), .B(n27074), .S(n27076), .Z(n25770) );
  MUX2_X1 U13170 ( .A(n27074), .B(n27075), .S(n27076), .Z(n27900) );
  MUX2_X1 U13171 ( .A(n25767), .B(n25768), .S(n27076), .Z(n25769) );
  INV_X1 U13172 ( .A(n23073), .ZN(n5856) );
  XNOR2_X1 U13173 ( .A(n14997), .B(n5858), .ZN(n5859) );
  NAND2_X1 U13176 ( .A1(n20340), .A2(n20504), .ZN(n5865) );
  NAND2_X1 U13177 ( .A1(n15006), .A2(n5866), .ZN(n15772) );
  INV_X1 U13178 ( .A(n8521), .ZN(n8812) );
  NOR2_X1 U13181 ( .A1(n5869), .A2(n8810), .ZN(n5868) );
  OR2_X1 U13182 ( .A1(n8808), .A2(n8521), .ZN(n5870) );
  XNOR2_X1 U13183 ( .A(n5872), .B(n24916), .ZN(n25722) );
  INV_X1 U13184 ( .A(n24949), .ZN(n5872) );
  XNOR2_X1 U13185 ( .A(n25244), .B(n5873), .ZN(n25245) );
  NAND3_X1 U13186 ( .A1(n5877), .A2(n27653), .A3(n5874), .ZN(n27654) );
  MUX2_X1 U13190 ( .A(n29090), .B(n27663), .S(n27672), .Z(n27196) );
  XNOR2_X1 U13191 ( .A(n22481), .B(n22502), .ZN(n22022) );
  NAND4_X2 U13192 ( .A1(n5880), .A2(n5878), .A3(n20949), .A4(n5879), .ZN(
        n22692) );
  NAND2_X1 U13193 ( .A1(n20947), .A2(n28185), .ZN(n5880) );
  INV_X1 U13194 ( .A(n28457), .ZN(n5882) );
  NAND2_X1 U13195 ( .A1(n23517), .A2(n474), .ZN(n23518) );
  INV_X1 U13197 ( .A(n23682), .ZN(n5883) );
  INV_X1 U13198 ( .A(n13912), .ZN(n14068) );
  INV_X1 U13199 ( .A(n13913), .ZN(n5887) );
  NAND2_X1 U13200 ( .A1(n8526), .A2(n5888), .ZN(n5961) );
  INV_X1 U13201 ( .A(n8687), .ZN(n5888) );
  NAND2_X1 U13204 ( .A1(n17005), .A2(n5891), .ZN(n16974) );
  OAI21_X1 U13205 ( .B1(n17720), .B2(n17425), .A(n5891), .ZN(n14227) );
  NAND2_X1 U13206 ( .A1(n14712), .A2(n13922), .ZN(n5894) );
  XNOR2_X1 U13207 ( .A(n21982), .B(n22152), .ZN(n22596) );
  NAND2_X1 U13208 ( .A1(n21304), .A2(n21305), .ZN(n5897) );
  NAND3_X1 U13209 ( .A1(n11947), .A2(n11952), .A3(n11951), .ZN(n5901) );
  NAND2_X1 U13210 ( .A1(n10917), .A2(n10605), .ZN(n5902) );
  NAND2_X1 U13211 ( .A1(n10914), .A2(n10913), .ZN(n5903) );
  XNOR2_X1 U13212 ( .A(n19472), .B(n19473), .ZN(n19479) );
  NAND2_X1 U13214 ( .A1(n17860), .A2(n17859), .ZN(n5906) );
  NAND2_X1 U13215 ( .A1(n18526), .A2(n18081), .ZN(n5907) );
  NAND2_X1 U13216 ( .A1(n18525), .A2(n5909), .ZN(n5908) );
  NAND3_X1 U13217 ( .A1(n5913), .A2(n5915), .A3(n5912), .ZN(n12257) );
  NAND2_X1 U13218 ( .A1(n5914), .A2(n5916), .ZN(n5912) );
  NAND3_X1 U13219 ( .A1(n5917), .A2(n28157), .A3(n5914), .ZN(n5913) );
  OAI21_X1 U13220 ( .B1(n10749), .B2(n3585), .A(n28638), .ZN(n5915) );
  NOR2_X1 U13221 ( .A1(n28569), .A2(n5918), .ZN(n13718) );
  NAND2_X1 U13222 ( .A1(n13587), .A2(n5918), .ZN(n14037) );
  NAND2_X1 U13223 ( .A1(n13997), .A2(n5918), .ZN(n13998) );
  NAND2_X1 U13224 ( .A1(n17182), .A2(n17183), .ZN(n5921) );
  XNOR2_X1 U13225 ( .A(n25436), .B(n26007), .ZN(n25395) );
  NAND2_X1 U13226 ( .A1(n24149), .A2(n5923), .ZN(n5922) );
  INV_X1 U13227 ( .A(n24740), .ZN(n5923) );
  XNOR2_X1 U13228 ( .A(n7415), .B(n7329), .ZN(n5925) );
  INV_X1 U13229 ( .A(n21084), .ZN(n5927) );
  INV_X1 U13230 ( .A(n20141), .ZN(n5929) );
  INV_X1 U13231 ( .A(n16575), .ZN(n15701) );
  NAND2_X1 U13235 ( .A1(n14237), .A2(n5936), .ZN(n13939) );
  NAND2_X1 U13236 ( .A1(n18838), .A2(n20077), .ZN(n5937) );
  NAND3_X1 U13238 ( .A1(n21028), .A2(n21029), .A3(n22142), .ZN(n5938) );
  INV_X1 U13239 ( .A(n22140), .ZN(n5939) );
  XNOR2_X1 U13240 ( .A(n16526), .B(n16605), .ZN(n16138) );
  INV_X1 U13241 ( .A(n16138), .ZN(n16139) );
  XNOR2_X1 U13242 ( .A(n14850), .B(n16138), .ZN(n14870) );
  INV_X1 U13243 ( .A(n17847), .ZN(n18138) );
  OAI211_X2 U13244 ( .C1(n21579), .C2(n5142), .A(n5942), .B(n5941), .ZN(n22033) );
  NAND2_X1 U13245 ( .A1(n20849), .A2(n5142), .ZN(n5941) );
  INV_X1 U13246 ( .A(n23126), .ZN(n6556) );
  NAND2_X1 U13247 ( .A1(n9045), .A2(n9230), .ZN(n5944) );
  NAND2_X1 U13248 ( .A1(n14315), .A2(n14320), .ZN(n5949) );
  XNOR2_X1 U13249 ( .A(n5950), .B(n17779), .ZN(n19949) );
  XNOR2_X1 U13250 ( .A(n5951), .B(n18670), .ZN(n5950) );
  XNOR2_X1 U13251 ( .A(n17770), .B(n5952), .ZN(n5951) );
  OAI21_X1 U13253 ( .B1(n21463), .B2(n5953), .A(n6636), .ZN(n20863) );
  NAND2_X1 U13254 ( .A1(n5955), .A2(n5954), .ZN(n21469) );
  OR2_X1 U13255 ( .A1(n21465), .A2(n21561), .ZN(n5954) );
  NAND2_X1 U13256 ( .A1(n29236), .A2(n21465), .ZN(n5955) );
  NAND2_X1 U13257 ( .A1(n6072), .A2(n9146), .ZN(n9373) );
  NAND3_X1 U13258 ( .A1(n6072), .A2(n9146), .A3(n5958), .ZN(n5957) );
  NAND2_X1 U13260 ( .A1(n8592), .A2(n8817), .ZN(n5962) );
  OAI21_X1 U13261 ( .B1(n12133), .B2(n11574), .A(n5963), .ZN(n5966) );
  OR2_X1 U13263 ( .A1(n16768), .A2(n5968), .ZN(n5967) );
  AND2_X2 U13264 ( .A1(n6252), .A2(n6254), .ZN(n15361) );
  NAND2_X1 U13265 ( .A1(n14508), .A2(n15360), .ZN(n5970) );
  NAND2_X1 U13266 ( .A1(n23407), .A2(n5971), .ZN(n24387) );
  INV_X1 U13267 ( .A(n12516), .ZN(n5974) );
  NAND2_X1 U13268 ( .A1(n5974), .A2(n12578), .ZN(n5973) );
  NAND3_X1 U13269 ( .A1(n5978), .A2(n14393), .A3(n14192), .ZN(n5977) );
  NAND2_X1 U13270 ( .A1(n13952), .A2(n13953), .ZN(n5979) );
  NAND2_X1 U13271 ( .A1(n14192), .A2(n14194), .ZN(n5980) );
  INV_X1 U13272 ( .A(n14194), .ZN(n5981) );
  NAND2_X1 U13273 ( .A1(n17266), .A2(n17267), .ZN(n17268) );
  INV_X1 U13274 ( .A(n5984), .ZN(n6644) );
  XNOR2_X1 U13275 ( .A(n5984), .B(n9242), .ZN(n10063) );
  XNOR2_X1 U13276 ( .A(n29136), .B(n1984), .ZN(n22637) );
  NAND2_X1 U13277 ( .A1(n17065), .A2(n16797), .ZN(n5988) );
  NAND2_X1 U13278 ( .A1(n7700), .A2(n5990), .ZN(n5989) );
  NAND2_X1 U13279 ( .A1(n7368), .A2(n7367), .ZN(n5990) );
  NAND2_X1 U13280 ( .A1(n5991), .A2(n28509), .ZN(n23958) );
  NAND2_X1 U13281 ( .A1(n17987), .A2(n29603), .ZN(n5992) );
  XNOR2_X1 U13282 ( .A(n19568), .B(n27298), .ZN(n19017) );
  NAND2_X1 U13283 ( .A1(n27673), .A2(n27671), .ZN(n27664) );
  NAND2_X1 U13284 ( .A1(n2011), .A2(n5994), .ZN(n5993) );
  XNOR2_X1 U13285 ( .A(n5995), .B(n1853), .ZN(n9843) );
  INV_X1 U13286 ( .A(n8883), .ZN(n5996) );
  INV_X1 U13287 ( .A(n12151), .ZN(n12149) );
  NAND2_X1 U13291 ( .A1(n6000), .A2(n14091), .ZN(n14120) );
  NOR2_X1 U13292 ( .A1(n14366), .A2(n6000), .ZN(n6045) );
  NAND3_X1 U13293 ( .A1(n14366), .A2(n6000), .A3(n14365), .ZN(n14367) );
  NAND2_X1 U13294 ( .A1(n13834), .A2(n6000), .ZN(n6046) );
  NAND2_X1 U13295 ( .A1(n17304), .A2(n6002), .ZN(n17013) );
  NAND3_X1 U13297 ( .A1(n15361), .A2(n14752), .A3(n6674), .ZN(n6004) );
  NAND2_X1 U13298 ( .A1(n6007), .A2(n6005), .ZN(n27691) );
  NAND2_X1 U13299 ( .A1(n6009), .A2(n6006), .ZN(n6005) );
  NAND2_X1 U13300 ( .A1(n6008), .A2(n455), .ZN(n6006) );
  NAND2_X1 U13301 ( .A1(n26127), .A2(n27702), .ZN(n6007) );
  AOI21_X1 U13302 ( .B1(n27700), .B2(n27701), .A(n27702), .ZN(n6009) );
  MUX2_X1 U13303 ( .A(n14044), .B(n14046), .S(n14047), .Z(n13908) );
  NAND2_X1 U13304 ( .A1(n13468), .A2(n6010), .ZN(n13470) );
  MUX2_X1 U13305 ( .A(n14046), .B(n13576), .S(n1896), .Z(n13580) );
  OAI21_X1 U13306 ( .B1(n17008), .B2(n17431), .A(n6012), .ZN(n17010) );
  NAND2_X1 U13307 ( .A1(n16846), .A2(n17426), .ZN(n6012) );
  INV_X1 U13308 ( .A(n17716), .ZN(n6013) );
  XNOR2_X1 U13309 ( .A(n6018), .B(n26101), .ZN(n26105) );
  NOR2_X1 U13310 ( .A1(n2656), .A2(n6526), .ZN(n6019) );
  NAND2_X1 U13311 ( .A1(n11053), .A2(n11165), .ZN(n6411) );
  OR2_X1 U13312 ( .A1(n12202), .A2(n2063), .ZN(n8650) );
  NAND2_X1 U13313 ( .A1(n11599), .A2(n6020), .ZN(n11601) );
  OAI21_X1 U13314 ( .B1(n11127), .B2(n11119), .A(n11118), .ZN(n6021) );
  NAND2_X1 U13315 ( .A1(n15102), .A2(n14575), .ZN(n6023) );
  OAI21_X1 U13316 ( .B1(n26296), .B2(n26351), .A(n26295), .ZN(n6025) );
  AOI22_X1 U13318 ( .A1(n26326), .A2(n27142), .B1(n26519), .B2(n29633), .ZN(
        n6026) );
  AND2_X1 U13319 ( .A1(n29070), .A2(n27772), .ZN(n26298) );
  NAND2_X1 U13320 ( .A1(n19999), .A2(n20353), .ZN(n6028) );
  NAND2_X1 U13321 ( .A1(n19997), .A2(n20480), .ZN(n20353) );
  NAND2_X1 U13323 ( .A1(n6029), .A2(n18357), .ZN(n18358) );
  OAI21_X1 U13324 ( .B1(n518), .B2(n18356), .A(n6030), .ZN(n6029) );
  NAND3_X1 U13325 ( .A1(n6033), .A2(n29544), .A3(n23679), .ZN(n23017) );
  NAND2_X1 U13326 ( .A1(n23167), .A2(n23680), .ZN(n6033) );
  INV_X1 U13327 ( .A(n23016), .ZN(n6034) );
  INV_X1 U13328 ( .A(n23167), .ZN(n6035) );
  AOI22_X1 U13329 ( .A1(n29120), .A2(n24800), .B1(n24804), .B2(n24806), .ZN(
        n24506) );
  NAND3_X1 U13330 ( .A1(n6038), .A2(n6037), .A3(n18457), .ZN(n6036) );
  OAI21_X1 U13331 ( .B1(n17902), .B2(n18111), .A(n18456), .ZN(n6037) );
  NAND2_X1 U13332 ( .A1(n20887), .A2(n21591), .ZN(n6040) );
  MUX2_X1 U13333 ( .A(n6043), .B(n6042), .S(n21591), .Z(n6041) );
  OAI21_X1 U13334 ( .B1(n20580), .B2(n28779), .A(n20941), .ZN(n20582) );
  OAI21_X1 U13335 ( .B1(n14146), .B2(n14008), .A(n6050), .ZN(n14148) );
  XNOR2_X1 U13336 ( .A(n13426), .B(n13427), .ZN(n6051) );
  NAND2_X1 U13337 ( .A1(n20755), .A2(n21463), .ZN(n6053) );
  INV_X1 U13338 ( .A(n23735), .ZN(n22949) );
  NAND2_X1 U13339 ( .A1(n23733), .A2(n23736), .ZN(n6054) );
  NAND2_X1 U13341 ( .A1(n24467), .A2(n29025), .ZN(n24579) );
  INV_X1 U13342 ( .A(n20334), .ZN(n6057) );
  NAND2_X1 U13343 ( .A1(n6057), .A2(n1881), .ZN(n20012) );
  INV_X1 U13344 ( .A(n9073), .ZN(n9071) );
  OAI21_X1 U13347 ( .B1(n6066), .B2(n14031), .A(n6062), .ZN(n6065) );
  NAND2_X1 U13348 ( .A1(n6063), .A2(n29107), .ZN(n6062) );
  INV_X1 U13349 ( .A(n13917), .ZN(n6063) );
  NAND2_X1 U13350 ( .A1(n6064), .A2(n13667), .ZN(n13979) );
  MUX2_X1 U13351 ( .A(n6065), .B(n13794), .S(n13921), .Z(n6064) );
  INV_X1 U13352 ( .A(n13917), .ZN(n6066) );
  OAI21_X1 U13353 ( .B1(n26567), .B2(n29610), .A(n6068), .ZN(n26915) );
  INV_X1 U13354 ( .A(n26565), .ZN(n6069) );
  NOR2_X1 U13355 ( .A1(n1872), .A2(n26568), .ZN(n6070) );
  INV_X1 U13356 ( .A(n9148), .ZN(n6072) );
  NAND2_X1 U13357 ( .A1(n578), .A2(n11867), .ZN(n6075) );
  NAND2_X1 U13358 ( .A1(n18470), .A2(n6079), .ZN(n6078) );
  NAND3_X1 U13359 ( .A1(n20206), .A2(n6083), .A3(n28501), .ZN(n6082) );
  NAND2_X1 U13360 ( .A1(n20552), .A2(n20404), .ZN(n6083) );
  NAND2_X1 U13362 ( .A1(n505), .A2(n20549), .ZN(n20206) );
  OAI21_X1 U13363 ( .B1(n28642), .B2(n26387), .A(n28572), .ZN(n6087) );
  XNOR2_X1 U13364 ( .A(n16505), .B(n16506), .ZN(n16507) );
  XNOR2_X1 U13365 ( .A(n15618), .B(n15992), .ZN(n16506) );
  NAND2_X1 U13366 ( .A1(n14742), .A2(n544), .ZN(n6088) );
  NAND3_X1 U13367 ( .A1(n14745), .A2(n15117), .A3(n14744), .ZN(n6089) );
  NAND2_X1 U13368 ( .A1(n14741), .A2(n15115), .ZN(n6090) );
  NAND2_X1 U13369 ( .A1(n6973), .A2(n7358), .ZN(n7357) );
  MUX2_X1 U13370 ( .A(n6973), .B(n29110), .S(n8231), .Z(n8233) );
  MUX2_X1 U13371 ( .A(n7620), .B(n29110), .S(n6973), .Z(n7623) );
  MUX2_X1 U13372 ( .A(n7431), .B(n6974), .S(n6973), .Z(n6975) );
  INV_X1 U13373 ( .A(n11350), .ZN(n11348) );
  XNOR2_X2 U13374 ( .A(n9130), .B(n9129), .ZN(n11350) );
  INV_X1 U13375 ( .A(n14484), .ZN(n14170) );
  INV_X1 U13377 ( .A(n14483), .ZN(n12122) );
  NAND2_X1 U13380 ( .A1(n8795), .A2(n8794), .ZN(n6092) );
  NAND2_X1 U13381 ( .A1(n7689), .A2(n7688), .ZN(n6093) );
  NAND2_X1 U13382 ( .A1(n7686), .A2(n7687), .ZN(n6094) );
  NAND2_X1 U13383 ( .A1(n6095), .A2(n27528), .ZN(n27096) );
  NOR2_X1 U13384 ( .A1(n6095), .A2(n27531), .ZN(n27508) );
  NAND2_X1 U13387 ( .A1(n24489), .A2(n29051), .ZN(n6098) );
  INV_X1 U13388 ( .A(n24100), .ZN(n6097) );
  NOR2_X1 U13389 ( .A1(n6099), .A2(n23706), .ZN(n23707) );
  NOR2_X1 U13390 ( .A1(n23220), .A2(n6099), .ZN(n6582) );
  OAI21_X1 U13391 ( .B1(n22451), .B2(n22452), .A(n6099), .ZN(n22454) );
  NAND2_X1 U13393 ( .A1(n17625), .A2(n18411), .ZN(n6103) );
  NAND2_X1 U13394 ( .A1(n6104), .A2(n21702), .ZN(n20994) );
  INV_X1 U13399 ( .A(n10919), .ZN(n11138) );
  INV_X1 U13401 ( .A(n10415), .ZN(n6107) );
  NAND2_X1 U13402 ( .A1(n6111), .A2(n24078), .ZN(n6109) );
  XNOR2_X1 U13403 ( .A(n6110), .B(n12503), .ZN(n25180) );
  NAND2_X1 U13404 ( .A1(n29584), .A2(n6114), .ZN(n19977) );
  OAI21_X1 U13405 ( .B1(n20178), .B2(n20173), .A(n6112), .ZN(n19868) );
  NAND2_X1 U13406 ( .A1(n6114), .A2(n20173), .ZN(n6112) );
  INV_X1 U13407 ( .A(n504), .ZN(n6113) );
  MUX2_X1 U13408 ( .A(n20177), .B(n20171), .S(n6114), .Z(n6341) );
  NAND2_X1 U13410 ( .A1(n6117), .A2(n6116), .ZN(n6115) );
  NAND2_X1 U13411 ( .A1(n21289), .A2(n21288), .ZN(n6118) );
  XNOR2_X1 U13412 ( .A(n22845), .B(n21872), .ZN(n22599) );
  XNOR2_X1 U13413 ( .A(n22845), .B(n6119), .ZN(n21786) );
  XNOR2_X1 U13414 ( .A(n25807), .B(n24890), .ZN(n6122) );
  NAND2_X1 U13415 ( .A1(n23936), .A2(n24556), .ZN(n6120) );
  NAND2_X1 U13416 ( .A1(n6123), .A2(n6097), .ZN(n23944) );
  OR2_X1 U13420 ( .A1(n17304), .A2(n28768), .ZN(n6128) );
  OAI211_X2 U13422 ( .C1(n6132), .C2(n11507), .A(n12283), .B(n11506), .ZN(
        n13150) );
  XNOR2_X1 U13423 ( .A(n9601), .B(n10231), .ZN(n9985) );
  XNOR2_X1 U13424 ( .A(n6134), .B(n6136), .ZN(n6133) );
  INV_X1 U13425 ( .A(n9985), .ZN(n6134) );
  NAND2_X1 U13426 ( .A1(n6140), .A2(n6139), .ZN(n17856) );
  OR2_X1 U13427 ( .A1(n6927), .A2(n17989), .ZN(n6139) );
  NAND2_X1 U13428 ( .A1(n17990), .A2(n6927), .ZN(n6140) );
  XNOR2_X1 U13429 ( .A(n22919), .B(n6141), .ZN(n22838) );
  XNOR2_X1 U13430 ( .A(n6141), .B(n22441), .ZN(n22443) );
  NAND2_X1 U13432 ( .A1(n13948), .A2(n14170), .ZN(n6142) );
  NAND2_X1 U13433 ( .A1(n10114), .A2(n11120), .ZN(n6144) );
  NAND2_X1 U13434 ( .A1(n11477), .A2(n11998), .ZN(n6145) );
  NAND2_X1 U13435 ( .A1(n12000), .A2(n11755), .ZN(n11540) );
  INV_X1 U13436 ( .A(n8908), .ZN(n6147) );
  INV_X1 U13437 ( .A(n27300), .ZN(n6150) );
  NAND2_X1 U13438 ( .A1(n6948), .A2(n26935), .ZN(n6148) );
  NAND2_X1 U13439 ( .A1(n26558), .A2(n26940), .ZN(n6149) );
  MUX2_X1 U13440 ( .A(n24760), .B(n24215), .S(n24756), .Z(n24216) );
  NAND2_X1 U13443 ( .A1(n20500), .A2(n29601), .ZN(n6156) );
  INV_X1 U13444 ( .A(n22139), .ZN(n21624) );
  XNOR2_X1 U13445 ( .A(n16198), .B(n16197), .ZN(n6160) );
  MUX2_X1 U13446 ( .A(n16706), .B(n16884), .S(n17526), .Z(n16885) );
  INV_X1 U13447 ( .A(n6162), .ZN(n7861) );
  NAND2_X1 U13448 ( .A1(n7308), .A2(n7172), .ZN(n6162) );
  NAND2_X1 U13449 ( .A1(n587), .A2(n29517), .ZN(n6164) );
  INV_X1 U13450 ( .A(n18856), .ZN(n18922) );
  OAI21_X1 U13451 ( .B1(n14334), .B2(n14410), .A(n14333), .ZN(n14335) );
  NAND2_X1 U13452 ( .A1(n6166), .A2(n29607), .ZN(n14333) );
  INV_X1 U13454 ( .A(n14408), .ZN(n6166) );
  OR2_X1 U13455 ( .A1(n24430), .A2(n19041), .ZN(n6171) );
  XNOR2_X1 U13456 ( .A(n25145), .B(n6167), .ZN(n25148) );
  XNOR2_X1 U13457 ( .A(n6168), .B(n365), .ZN(n6167) );
  OAI211_X1 U13458 ( .C1(n6171), .C2(n24429), .A(n6169), .B(n6170), .ZN(n6168)
         );
  NAND2_X1 U13459 ( .A1(n24429), .A2(n19041), .ZN(n6169) );
  NAND2_X1 U13460 ( .A1(n24430), .A2(n19041), .ZN(n6170) );
  NOR2_X2 U13461 ( .A1(n24429), .A2(n24430), .ZN(n25867) );
  XNOR2_X1 U13462 ( .A(n15575), .B(n26656), .ZN(n15763) );
  INV_X1 U13463 ( .A(n16579), .ZN(n6173) );
  XNOR2_X1 U13464 ( .A(n15575), .B(n6173), .ZN(n15658) );
  XNOR2_X1 U13465 ( .A(n15575), .B(n6174), .ZN(n15904) );
  NAND2_X1 U13467 ( .A1(n17547), .A2(n16947), .ZN(n6175) );
  NAND2_X1 U13468 ( .A1(n18529), .A2(n17864), .ZN(n6177) );
  AND2_X2 U13469 ( .A1(n6179), .A2(n6178), .ZN(n17864) );
  NAND2_X1 U13470 ( .A1(n16933), .A2(n17046), .ZN(n6178) );
  NAND2_X1 U13471 ( .A1(n16934), .A2(n6180), .ZN(n6179) );
  INV_X1 U13472 ( .A(n11458), .ZN(n6181) );
  INV_X1 U13473 ( .A(n11457), .ZN(n11460) );
  INV_X1 U13474 ( .A(n11152), .ZN(n6182) );
  NAND2_X1 U13475 ( .A1(n6182), .A2(n11158), .ZN(n10494) );
  OAI21_X2 U13476 ( .B1(n27171), .B2(n6185), .A(n27170), .ZN(n27672) );
  NAND2_X1 U13477 ( .A1(n6567), .A2(n20618), .ZN(n19921) );
  INV_X1 U13478 ( .A(n9030), .ZN(n8433) );
  NOR2_X1 U13479 ( .A1(n28210), .A2(n9030), .ZN(n6188) );
  NAND3_X1 U13480 ( .A1(n9027), .A2(n9030), .A3(n7714), .ZN(n6191) );
  INV_X1 U13481 ( .A(n6193), .ZN(n19338) );
  XNOR2_X1 U13482 ( .A(n19220), .B(n19111), .ZN(n6193) );
  NOR2_X1 U13483 ( .A1(n6294), .A2(n28122), .ZN(n6196) );
  INV_X1 U13484 ( .A(n23139), .ZN(n6194) );
  NAND2_X1 U13485 ( .A1(n23427), .A2(n23138), .ZN(n23139) );
  INV_X1 U13487 ( .A(n6200), .ZN(n6199) );
  OAI22_X1 U13488 ( .A1(n7241), .A2(n7995), .B1(n7993), .B2(n6201), .ZN(n6200)
         );
  OR2_X1 U13489 ( .A1(n7992), .A2(n7876), .ZN(n6201) );
  MUX2_X1 U13490 ( .A(n27300), .B(n5425), .S(n27301), .Z(n26689) );
  NAND2_X1 U13492 ( .A1(n6203), .A2(n28417), .ZN(n6202) );
  INV_X1 U13493 ( .A(n19928), .ZN(n6203) );
  NAND2_X1 U13494 ( .A1(n20451), .A2(n20449), .ZN(n6204) );
  AND2_X1 U13495 ( .A1(n28417), .A2(n20265), .ZN(n6205) );
  MUX2_X1 U13496 ( .A(n20449), .B(n28552), .S(n28417), .Z(n20452) );
  INV_X1 U13497 ( .A(n21749), .ZN(n21643) );
  NAND2_X1 U13498 ( .A1(n20659), .A2(n21748), .ZN(n6206) );
  XOR2_X1 U13499 ( .A(n16090), .B(n16233), .Z(n15366) );
  NAND2_X1 U13500 ( .A1(n7231), .A2(n7591), .ZN(n7318) );
  NAND2_X1 U13501 ( .A1(n6210), .A2(n29629), .ZN(n7727) );
  NAND2_X1 U13502 ( .A1(n6211), .A2(n22944), .ZN(n22593) );
  NAND2_X1 U13503 ( .A1(n28181), .A2(n23738), .ZN(n6211) );
  INV_X1 U13504 ( .A(n21738), .ZN(n6212) );
  NAND3_X1 U13505 ( .A1(n1814), .A2(n20841), .A3(n21458), .ZN(n6213) );
  XNOR2_X1 U13506 ( .A(n24852), .B(n2306), .ZN(n24453) );
  NAND2_X1 U13508 ( .A1(n28552), .A2(n21063), .ZN(n6219) );
  AOI21_X1 U13509 ( .B1(n9686), .B2(n1933), .A(n29637), .ZN(n10485) );
  AOI22_X1 U13510 ( .A1(n10486), .A2(n29637), .B1(n10487), .B2(n1933), .ZN(
        n10488) );
  OAI21_X1 U13511 ( .B1(n9248), .B2(n9245), .A(n28211), .ZN(n7161) );
  XNOR2_X1 U13512 ( .A(n16588), .B(n1980), .ZN(n15280) );
  AOI211_X1 U13514 ( .C1(n28482), .C2(n377), .A(n6222), .B(n26461), .ZN(n6221)
         );
  AND2_X1 U13515 ( .A1(n28476), .A2(n26559), .ZN(n6222) );
  NAND2_X1 U13517 ( .A1(n6225), .A2(n18354), .ZN(n17919) );
  NAND2_X1 U13518 ( .A1(n17666), .A2(n6225), .ZN(n17668) );
  INV_X1 U13519 ( .A(n13458), .ZN(n13460) );
  NAND3_X1 U13520 ( .A1(n2012), .A2(n11592), .A3(n12581), .ZN(n13458) );
  NAND4_X1 U13521 ( .A1(n1864), .A2(n6226), .A3(n27302), .A4(n27301), .ZN(
        n27307) );
  XNOR2_X1 U13522 ( .A(n20735), .B(n20734), .ZN(n6227) );
  XNOR2_X1 U13523 ( .A(n19717), .B(n19668), .ZN(n19399) );
  NAND2_X1 U13525 ( .A1(n13728), .A2(n14135), .ZN(n6233) );
  NAND2_X1 U13526 ( .A1(n20381), .A2(n28637), .ZN(n6236) );
  NAND2_X1 U13527 ( .A1(n20779), .A2(n20778), .ZN(n6240) );
  OAI211_X1 U13528 ( .C1(n10549), .C2(n10492), .A(n11115), .B(n6241), .ZN(
        n6242) );
  NOR2_X1 U13529 ( .A1(n17854), .A2(n6526), .ZN(n17988) );
  NAND2_X1 U13530 ( .A1(n17988), .A2(n18367), .ZN(n6243) );
  XNOR2_X1 U13531 ( .A(n16291), .B(n14709), .ZN(n16270) );
  NAND2_X1 U13532 ( .A1(n14704), .A2(n6244), .ZN(n16291) );
  NAND3_X1 U13533 ( .A1(n6245), .A2(n6246), .A3(n15268), .ZN(n6244) );
  NAND2_X1 U13534 ( .A1(n6250), .A2(n6249), .ZN(n6248) );
  NAND2_X1 U13535 ( .A1(n242), .A2(n10549), .ZN(n6249) );
  NAND2_X1 U13536 ( .A1(n6253), .A2(n13724), .ZN(n6252) );
  NAND2_X1 U13537 ( .A1(n14148), .A2(n14374), .ZN(n6253) );
  XNOR2_X1 U13540 ( .A(n10018), .B(n10016), .ZN(n6257) );
  NAND2_X1 U13541 ( .A1(n11136), .A2(n11142), .ZN(n11139) );
  INV_X1 U13542 ( .A(n11139), .ZN(n10463) );
  NAND2_X1 U13544 ( .A1(n20190), .A2(n20547), .ZN(n6259) );
  INV_X1 U13549 ( .A(n24408), .ZN(n6265) );
  INV_X1 U13550 ( .A(n24404), .ZN(n6266) );
  OAI21_X1 U13551 ( .B1(n27539), .B2(n27548), .A(n27538), .ZN(n6268) );
  XNOR2_X1 U13552 ( .A(n6647), .B(n13208), .ZN(n13542) );
  NAND2_X1 U13553 ( .A1(n10749), .A2(n11198), .ZN(n6271) );
  NAND2_X1 U13554 ( .A1(n21658), .A2(n21657), .ZN(n6273) );
  NAND2_X1 U13555 ( .A1(n21659), .A2(n6275), .ZN(n6274) );
  INV_X1 U13556 ( .A(n6276), .ZN(n19144) );
  XNOR2_X1 U13557 ( .A(n19145), .B(n6276), .ZN(n6606) );
  INV_X1 U13558 ( .A(n18948), .ZN(n19199) );
  NOR2_X1 U13559 ( .A1(n23393), .A2(n23392), .ZN(n6277) );
  AOI21_X1 U13560 ( .B1(n23838), .B2(n6610), .A(n6279), .ZN(n6278) );
  INV_X1 U13561 ( .A(n23391), .ZN(n6279) );
  NAND2_X1 U13562 ( .A1(n7662), .A2(n8265), .ZN(n9084) );
  OR2_X2 U13563 ( .A1(n12846), .A2(n6283), .ZN(n14575) );
  NAND2_X1 U13564 ( .A1(n18540), .A2(n18539), .ZN(n6284) );
  NAND2_X1 U13565 ( .A1(n18541), .A2(n18529), .ZN(n6285) );
  NAND2_X1 U13566 ( .A1(n7233), .A2(n7231), .ZN(n7594) );
  INV_X1 U13568 ( .A(n28549), .ZN(n27353) );
  INV_X1 U13569 ( .A(n11176), .ZN(n11334) );
  NOR2_X1 U13570 ( .A1(n6292), .A2(n6290), .ZN(n16755) );
  NOR2_X1 U13571 ( .A1(n17229), .A2(n6291), .ZN(n6290) );
  NAND2_X1 U13572 ( .A1(n17567), .A2(n17568), .ZN(n6291) );
  NAND2_X1 U13573 ( .A1(n15279), .A2(n6293), .ZN(n6493) );
  XNOR2_X1 U13574 ( .A(n15545), .B(n6296), .ZN(n15836) );
  INV_X1 U13575 ( .A(n13456), .ZN(n6297) );
  AOI21_X1 U13576 ( .B1(n6299), .B2(n8024), .A(n29130), .ZN(n8025) );
  NAND2_X1 U13578 ( .A1(n26860), .A2(n29633), .ZN(n6300) );
  NAND3_X1 U13579 ( .A1(n26855), .A2(n27142), .A3(n28487), .ZN(n6301) );
  NAND2_X1 U13580 ( .A1(n26325), .A2(n27139), .ZN(n6302) );
  INV_X1 U13581 ( .A(n27141), .ZN(n27139) );
  OAI21_X1 U13585 ( .B1(n24288), .B2(n24597), .A(n24148), .ZN(n23933) );
  XNOR2_X1 U13586 ( .A(n22248), .B(n2350), .ZN(n21902) );
  OAI21_X2 U13587 ( .B1(n6321), .B2(n6835), .A(n23954), .ZN(n25773) );
  NAND3_X1 U13588 ( .A1(n6325), .A2(n16711), .A3(n6324), .ZN(n16718) );
  NAND2_X1 U13589 ( .A1(n16709), .A2(n17335), .ZN(n6324) );
  NAND2_X1 U13590 ( .A1(n16710), .A2(n17342), .ZN(n6325) );
  INV_X1 U13591 ( .A(n19534), .ZN(n6327) );
  XNOR2_X1 U13592 ( .A(n6327), .B(n19220), .ZN(n18984) );
  NAND2_X1 U13593 ( .A1(n12240), .A2(n11969), .ZN(n12242) );
  NAND2_X1 U13594 ( .A1(n12156), .A2(n12158), .ZN(n12240) );
  NAND2_X1 U13595 ( .A1(n10453), .A2(n11876), .ZN(n10869) );
  NAND2_X1 U13596 ( .A1(n11879), .A2(n567), .ZN(n6329) );
  NAND3_X1 U13597 ( .A1(n1926), .A2(n15013), .A3(n15014), .ZN(n6332) );
  NAND2_X1 U13600 ( .A1(n6338), .A2(n23830), .ZN(n6579) );
  INV_X1 U13602 ( .A(n20053), .ZN(n20172) );
  XNOR2_X1 U13603 ( .A(n13350), .B(n12822), .ZN(n6343) );
  NAND2_X1 U13604 ( .A1(n6348), .A2(n23842), .ZN(n24492) );
  NAND2_X1 U13605 ( .A1(n6348), .A2(n24471), .ZN(n23850) );
  NOR2_X1 U13606 ( .A1(n29033), .A2(n6348), .ZN(n24473) );
  NAND3_X1 U13607 ( .A1(n24100), .A2(n29033), .A3(n6348), .ZN(n24101) );
  AOI21_X1 U13608 ( .B1(n24490), .B2(n24489), .A(n6348), .ZN(n24495) );
  OAI211_X1 U13609 ( .C1(n21442), .C2(n6275), .A(n21441), .B(n21440), .ZN(
        n6350) );
  NAND2_X1 U13610 ( .A1(n13729), .A2(n13912), .ZN(n14070) );
  NAND3_X1 U13611 ( .A1(n6462), .A2(n6354), .A3(n6353), .ZN(n6356) );
  NAND2_X1 U13612 ( .A1(n28554), .A2(n23765), .ZN(n6353) );
  NAND2_X1 U13613 ( .A1(n23764), .A2(n23763), .ZN(n6354) );
  NAND3_X1 U13614 ( .A1(n6356), .A2(n6357), .A3(n6355), .ZN(n24502) );
  NAND2_X1 U13615 ( .A1(n23766), .A2(n6358), .ZN(n6357) );
  NAND2_X1 U13616 ( .A1(n7813), .A2(n10806), .ZN(n6359) );
  NAND2_X1 U13617 ( .A1(n10512), .A2(n10544), .ZN(n6361) );
  INV_X1 U13618 ( .A(n21304), .ZN(n6362) );
  INV_X1 U13619 ( .A(n22301), .ZN(n22757) );
  NAND2_X1 U13620 ( .A1(n6363), .A2(n20327), .ZN(n22301) );
  NAND2_X1 U13621 ( .A1(n8825), .A2(n29147), .ZN(n8584) );
  NAND3_X1 U13622 ( .A1(n8825), .A2(n8586), .A3(n8824), .ZN(n8834) );
  NAND2_X1 U13623 ( .A1(n6365), .A2(n6086), .ZN(n19856) );
  NAND2_X1 U13624 ( .A1(n20206), .A2(n20404), .ZN(n6365) );
  NAND2_X1 U13625 ( .A1(n10972), .A2(n10976), .ZN(n6367) );
  NAND3_X1 U13626 ( .A1(n21484), .A2(n21581), .A3(n21481), .ZN(n6369) );
  NAND2_X1 U13627 ( .A1(n6371), .A2(n16814), .ZN(n16817) );
  OR2_X1 U13628 ( .A1(n17097), .A2(n16815), .ZN(n17104) );
  NAND3_X1 U13629 ( .A1(n6371), .A2(n1466), .A3(n16860), .ZN(n16680) );
  INV_X1 U13630 ( .A(n17097), .ZN(n6371) );
  NAND2_X1 U13631 ( .A1(n12510), .A2(n6372), .ZN(n11993) );
  INV_X1 U13633 ( .A(n6375), .ZN(n12685) );
  XNOR2_X1 U13634 ( .A(n6375), .B(n12389), .ZN(n12393) );
  NAND2_X1 U13635 ( .A1(n18341), .A2(n18342), .ZN(n6376) );
  NAND2_X1 U13636 ( .A1(n24727), .A2(n29695), .ZN(n6377) );
  NAND2_X1 U13637 ( .A1(n24596), .A2(n24288), .ZN(n24724) );
  XNOR2_X1 U13638 ( .A(n22691), .B(n22437), .ZN(n21739) );
  NAND2_X1 U13639 ( .A1(n7234), .A2(n7591), .ZN(n6381) );
  NOR2_X1 U13640 ( .A1(n11048), .A2(n11266), .ZN(n6385) );
  INV_X1 U13641 ( .A(n29122), .ZN(n11044) );
  NAND3_X1 U13642 ( .A1(n17906), .A2(n17947), .A3(n18341), .ZN(n6387) );
  XNOR2_X1 U13643 ( .A(n22246), .B(n22265), .ZN(n6388) );
  NAND2_X1 U13644 ( .A1(n6392), .A2(n6390), .ZN(n16388) );
  NAND2_X1 U13645 ( .A1(n15263), .A2(n6391), .ZN(n6390) );
  OAI21_X1 U13646 ( .B1(n6393), .B2(n14761), .A(n15264), .ZN(n6392) );
  NAND2_X1 U13648 ( .A1(n21270), .A2(n21271), .ZN(n6394) );
  NAND2_X1 U13650 ( .A1(n20815), .A2(n21269), .ZN(n21272) );
  NAND2_X1 U13651 ( .A1(n6398), .A2(n29488), .ZN(n6397) );
  NAND2_X1 U13652 ( .A1(n21267), .A2(n21268), .ZN(n6398) );
  NAND2_X1 U13653 ( .A1(n16930), .A2(n6403), .ZN(n6402) );
  NAND3_X1 U13654 ( .A1(n8610), .A2(n8749), .A3(n9533), .ZN(n6404) );
  NAND2_X1 U13655 ( .A1(n6413), .A2(n694), .ZN(n6412) );
  NAND2_X1 U13656 ( .A1(n14781), .A2(n15338), .ZN(n6413) );
  XNOR2_X1 U13657 ( .A(n21791), .B(n21792), .ZN(n6414) );
  XNOR2_X2 U13658 ( .A(n6414), .B(n21795), .ZN(n23764) );
  XNOR2_X1 U13659 ( .A(n16518), .B(n15941), .ZN(n6415) );
  XNOR2_X1 U13660 ( .A(n15942), .B(n5858), .ZN(n6416) );
  AOI21_X1 U13661 ( .B1(n17037), .B2(n6417), .A(n17569), .ZN(n17042) );
  OAI21_X1 U13662 ( .B1(n4784), .B2(n24466), .A(n6421), .ZN(n6420) );
  NAND2_X1 U13665 ( .A1(n12481), .A2(n14215), .ZN(n14214) );
  NAND2_X1 U13666 ( .A1(n555), .A2(n12481), .ZN(n12470) );
  NAND3_X1 U13670 ( .A1(n6432), .A2(n12332), .A3(n12327), .ZN(n10537) );
  NAND2_X1 U13671 ( .A1(n12018), .A2(n6432), .ZN(n12334) );
  NAND2_X1 U13672 ( .A1(n12016), .A2(n6432), .ZN(n10536) );
  NAND2_X1 U13673 ( .A1(n12015), .A2(n6432), .ZN(n11890) );
  NAND3_X1 U13674 ( .A1(n11449), .A2(n12332), .A3(n6432), .ZN(n6431) );
  NAND3_X1 U13675 ( .A1(n4118), .A2(n17569), .A3(n17227), .ZN(n16756) );
  NAND2_X1 U13677 ( .A1(n14313), .A2(n14314), .ZN(n6434) );
  XNOR2_X1 U13679 ( .A(n25061), .B(n25060), .ZN(n6436) );
  NAND2_X1 U13680 ( .A1(n26918), .A2(n457), .ZN(n6438) );
  XNOR2_X1 U13681 ( .A(n10146), .B(n9934), .ZN(n6440) );
  XNOR2_X1 U13683 ( .A(n16076), .B(n6448), .ZN(n6447) );
  XNOR2_X1 U13684 ( .A(n6449), .B(n29319), .ZN(n6448) );
  NAND2_X1 U13685 ( .A1(n8871), .A2(n7568), .ZN(n6450) );
  NAND2_X1 U13686 ( .A1(n9059), .A2(n9064), .ZN(n8868) );
  INV_X1 U13687 ( .A(n16323), .ZN(n6454) );
  INV_X1 U13688 ( .A(n16323), .ZN(n16455) );
  OR2_X1 U13689 ( .A1(n15318), .A2(n15319), .ZN(n6457) );
  XNOR2_X1 U13690 ( .A(n6458), .B(n1928), .ZN(n20837) );
  XNOR2_X1 U13691 ( .A(n6458), .B(n3369), .ZN(n22368) );
  XNOR2_X1 U13692 ( .A(n21805), .B(n6458), .ZN(n21816) );
  XNOR2_X1 U13693 ( .A(n22180), .B(n6458), .ZN(n22902) );
  XNOR2_X1 U13694 ( .A(n22609), .B(n6458), .ZN(n22612) );
  NAND2_X1 U13697 ( .A1(n21829), .A2(n6462), .ZN(n6461) );
  XNOR2_X2 U13698 ( .A(n8991), .B(n8990), .ZN(n11322) );
  OAI21_X1 U13701 ( .B1(n27592), .B2(n26285), .A(n27597), .ZN(n6464) );
  INV_X1 U13702 ( .A(n17272), .ZN(n6465) );
  INV_X1 U13703 ( .A(n14416), .ZN(n6466) );
  NAND2_X1 U13705 ( .A1(n14420), .A2(n14421), .ZN(n14448) );
  OR2_X1 U13706 ( .A1(n14416), .A2(n14414), .ZN(n14421) );
  XNOR2_X1 U13707 ( .A(n19290), .B(n6468), .ZN(n6467) );
  NAND2_X1 U13711 ( .A1(n885), .A2(n29564), .ZN(n6474) );
  NAND2_X1 U13714 ( .A1(n6480), .A2(n6479), .ZN(n6478) );
  NOR2_X1 U13715 ( .A1(n16539), .A2(n28801), .ZN(n6485) );
  NAND2_X1 U13716 ( .A1(n17899), .A2(n6484), .ZN(n6483) );
  INV_X1 U13717 ( .A(n18356), .ZN(n6484) );
  XNOR2_X1 U13720 ( .A(n6487), .B(n19276), .ZN(n20597) );
  INV_X2 U13721 ( .A(n6488), .ZN(n19487) );
  XNOR2_X1 U13722 ( .A(n19313), .B(n19487), .ZN(n18210) );
  NAND3_X1 U13723 ( .A1(n27772), .A2(n29537), .A3(n29022), .ZN(n27774) );
  OAI22_X1 U13724 ( .A1(n27233), .A2(n6490), .B1(n27762), .B2(n29022), .ZN(
        n27234) );
  OR2_X1 U13725 ( .A1(n26289), .A2(n29633), .ZN(n6492) );
  INV_X1 U13727 ( .A(n20081), .ZN(n6495) );
  NAND2_X1 U13728 ( .A1(n19846), .A2(n29145), .ZN(n6494) );
  XNOR2_X1 U13730 ( .A(n6496), .B(n15576), .ZN(Ciphertext[123]) );
  NAND3_X1 U13731 ( .A1(n6498), .A2(n27770), .A3(n6497), .ZN(n6496) );
  NAND2_X1 U13732 ( .A1(n29117), .A2(n27769), .ZN(n6497) );
  XNOR2_X1 U13733 ( .A(n16379), .B(n16378), .ZN(n6502) );
  NAND3_X1 U13734 ( .A1(n21493), .A2(n21185), .A3(n21496), .ZN(n6503) );
  NAND2_X1 U13735 ( .A1(n9042), .A2(n9247), .ZN(n6505) );
  NAND2_X1 U13736 ( .A1(n24417), .A2(n24341), .ZN(n6506) );
  INV_X1 U13737 ( .A(n25998), .ZN(n6507) );
  NAND2_X1 U13738 ( .A1(n19858), .A2(n20412), .ZN(n6509) );
  OAI21_X1 U13739 ( .B1(n11188), .B2(n11322), .A(n6510), .ZN(n10813) );
  INV_X1 U13741 ( .A(n15274), .ZN(n14698) );
  NAND2_X1 U13742 ( .A1(n20481), .A2(n20485), .ZN(n6512) );
  NAND2_X1 U13743 ( .A1(n10669), .A2(n10670), .ZN(n6516) );
  XNOR2_X1 U13744 ( .A(n13482), .B(n13273), .ZN(n12944) );
  NAND3_X1 U13745 ( .A1(n11680), .A2(n5009), .A3(n11541), .ZN(n6518) );
  XNOR2_X1 U13746 ( .A(n6520), .B(n29549), .ZN(n21884) );
  XNOR2_X1 U13747 ( .A(n6520), .B(n22110), .ZN(n22111) );
  NAND2_X1 U13749 ( .A1(n6522), .A2(n6521), .ZN(n15449) );
  OAI21_X1 U13750 ( .B1(n15327), .B2(n15322), .A(n6522), .ZN(n13978) );
  NAND2_X1 U13751 ( .A1(n15327), .A2(n15323), .ZN(n6522) );
  AND2_X1 U13752 ( .A1(n23290), .A2(n23816), .ZN(n23821) );
  INV_X1 U13754 ( .A(n12775), .ZN(n12476) );
  NAND2_X1 U13755 ( .A1(n17000), .A2(n17402), .ZN(n6524) );
  XNOR2_X1 U13757 ( .A(n22271), .B(n22248), .ZN(n22728) );
  XNOR2_X1 U13758 ( .A(n22728), .B(n22727), .ZN(n22729) );
  XNOR2_X1 U13759 ( .A(n19631), .B(n19632), .ZN(n6535) );
  XNOR2_X1 U13760 ( .A(n19634), .B(n19635), .ZN(n6536) );
  NAND3_X1 U13761 ( .A1(n24712), .A2(n28524), .A3(n24713), .ZN(n24352) );
  NAND2_X1 U13762 ( .A1(n23055), .A2(n23054), .ZN(n6537) );
  MUX2_X1 U13763 ( .A(n29573), .B(n26799), .S(n26278), .Z(n6541) );
  OAI22_X1 U13765 ( .A1(n6542), .A2(n10593), .B1(n10705), .B2(n10944), .ZN(
        n10596) );
  NAND2_X1 U13767 ( .A1(n9581), .A2(n9580), .ZN(n9579) );
  OAI211_X2 U13768 ( .C1(n7314), .C2(n7900), .A(n6546), .B(n6545), .ZN(n7569)
         );
  NAND3_X1 U13769 ( .A1(n7804), .A2(n7800), .A3(n7898), .ZN(n6546) );
  NAND2_X1 U13770 ( .A1(n24423), .A2(n24422), .ZN(n6548) );
  INV_X1 U13771 ( .A(n12359), .ZN(n12361) );
  NAND2_X1 U13772 ( .A1(n11739), .A2(n11740), .ZN(n12360) );
  NAND3_X1 U13773 ( .A1(n11742), .A2(n11740), .A3(n12359), .ZN(n6549) );
  NAND3_X1 U13774 ( .A1(n12363), .A2(n12362), .A3(n12361), .ZN(n6550) );
  NAND2_X1 U13775 ( .A1(n12357), .A2(n12356), .ZN(n6552) );
  NAND2_X1 U13776 ( .A1(n17544), .A2(n17543), .ZN(n6553) );
  NAND2_X1 U13777 ( .A1(n6555), .A2(n17217), .ZN(n6554) );
  MUX2_X1 U13778 ( .A(n17540), .B(n17539), .S(n17545), .Z(n6555) );
  NAND2_X1 U13779 ( .A1(n16939), .A2(n28454), .ZN(n17546) );
  NAND2_X1 U13782 ( .A1(n24547), .A2(n6556), .ZN(n6868) );
  NOR2_X1 U13783 ( .A1(n24547), .A2(n6556), .ZN(n23129) );
  AOI21_X1 U13784 ( .B1(n24543), .B2(n24544), .A(n6556), .ZN(n24545) );
  NAND2_X1 U13785 ( .A1(n22965), .A2(n29020), .ZN(n6558) );
  NOR2_X1 U13786 ( .A1(n6559), .A2(n16723), .ZN(n16726) );
  NAND2_X1 U13787 ( .A1(n17476), .A2(n6560), .ZN(n16801) );
  OR2_X1 U13788 ( .A1(n14107), .A2(n6563), .ZN(n6562) );
  INV_X1 U13790 ( .A(n20617), .ZN(n20432) );
  NOR2_X2 U13791 ( .A1(n20434), .A2(n6564), .ZN(n21514) );
  OAI21_X1 U13792 ( .B1(n20617), .B2(n6567), .A(n6566), .ZN(n6565) );
  NAND2_X1 U13793 ( .A1(n6567), .A2(n20619), .ZN(n6566) );
  INV_X1 U13794 ( .A(n20431), .ZN(n6567) );
  NOR2_X1 U13795 ( .A1(n20635), .A2(n20248), .ZN(n20032) );
  NAND2_X1 U13797 ( .A1(n13943), .A2(n15194), .ZN(n14175) );
  NAND2_X1 U13798 ( .A1(n6571), .A2(n13943), .ZN(n6572) );
  INV_X1 U13799 ( .A(n15415), .ZN(n15410) );
  XNOR2_X1 U13800 ( .A(n18802), .B(n19643), .ZN(n19039) );
  NAND2_X1 U13801 ( .A1(n18479), .A2(n18011), .ZN(n6574) );
  NAND2_X1 U13802 ( .A1(n6576), .A2(n18475), .ZN(n6575) );
  INV_X1 U13803 ( .A(n20219), .ZN(n19992) );
  INV_X1 U13804 ( .A(n18972), .ZN(n6578) );
  NOR2_X1 U13806 ( .A1(n28551), .A2(n23281), .ZN(n6580) );
  NAND3_X1 U13807 ( .A1(n27433), .A2(n25417), .A3(n26830), .ZN(n25424) );
  NAND2_X1 U13808 ( .A1(n28622), .A2(n6582), .ZN(n6584) );
  NAND2_X1 U13809 ( .A1(n22084), .A2(n23700), .ZN(n6587) );
  NAND2_X1 U13811 ( .A1(n22085), .A2(n6587), .ZN(n6586) );
  NAND2_X1 U13812 ( .A1(n17717), .A2(n17720), .ZN(n6588) );
  NAND3_X1 U13813 ( .A1(n9235), .A2(n9047), .A3(n6590), .ZN(n9048) );
  XNOR2_X1 U13814 ( .A(n6591), .B(n3654), .ZN(Ciphertext[81]) );
  NAND2_X1 U13815 ( .A1(n6594), .A2(n6593), .ZN(n6592) );
  NAND2_X1 U13816 ( .A1(n27554), .A2(n29085), .ZN(n6593) );
  NAND2_X1 U13817 ( .A1(n27149), .A2(n29578), .ZN(n6594) );
  NAND2_X1 U13818 ( .A1(n24503), .A2(n6596), .ZN(n6595) );
  OAI21_X1 U13820 ( .B1(n10572), .B2(n10883), .A(n6603), .ZN(n10655) );
  NAND2_X1 U13821 ( .A1(n11212), .A2(n10883), .ZN(n6603) );
  AND2_X1 U13822 ( .A1(n6605), .A2(n20504), .ZN(n19799) );
  XNOR2_X2 U13823 ( .A(n19148), .B(n6606), .ZN(n20504) );
  INV_X1 U13824 ( .A(n20339), .ZN(n6605) );
  NAND2_X1 U13825 ( .A1(n23791), .A2(n23789), .ZN(n6607) );
  INV_X1 U13826 ( .A(n23280), .ZN(n6610) );
  INV_X1 U13827 ( .A(n24707), .ZN(n24124) );
  NOR2_X1 U13828 ( .A1(n24704), .A2(n24707), .ZN(n6612) );
  INV_X1 U13829 ( .A(n7997), .ZN(n7998) );
  OAI211_X1 U13830 ( .C1(n6623), .C2(n6622), .A(n6616), .B(n6618), .ZN(
        Ciphertext[9]) );
  INV_X1 U13831 ( .A(n27367), .ZN(n6617) );
  INV_X1 U13832 ( .A(n6619), .ZN(n6618) );
  OAI21_X1 U13833 ( .B1(n3751), .B2(n27375), .A(n6620), .ZN(n6619) );
  NAND3_X1 U13834 ( .A1(n27375), .A2(n27374), .A3(n3751), .ZN(n6622) );
  AOI21_X1 U13835 ( .B1(n27369), .B2(n6624), .A(n27364), .ZN(n6623) );
  OR2_X1 U13836 ( .A1(n27370), .A2(n29541), .ZN(n6624) );
  NAND2_X1 U13837 ( .A1(n26237), .A2(n26757), .ZN(n26760) );
  NAND2_X1 U13838 ( .A1(n6625), .A2(n26237), .ZN(n6626) );
  NAND2_X1 U13839 ( .A1(n26756), .A2(n26241), .ZN(n6627) );
  OAI21_X1 U13841 ( .B1(n23458), .B2(n23461), .A(n23357), .ZN(n6628) );
  INV_X1 U13842 ( .A(n23148), .ZN(n23455) );
  NAND2_X1 U13843 ( .A1(n11266), .A2(n29122), .ZN(n6631) );
  NAND2_X1 U13845 ( .A1(n25079), .A2(n26422), .ZN(n6634) );
  INV_X1 U13846 ( .A(n21565), .ZN(n6636) );
  XNOR2_X1 U13847 ( .A(n15635), .B(n6637), .ZN(n15638) );
  INV_X1 U13848 ( .A(n6637), .ZN(n16266) );
  NAND2_X1 U13849 ( .A1(n17273), .A2(n539), .ZN(n6638) );
  NAND2_X1 U13850 ( .A1(n13916), .A2(n6066), .ZN(n6639) );
  XNOR2_X1 U13851 ( .A(n6644), .B(n9787), .ZN(n9792) );
  NAND2_X1 U13852 ( .A1(n11361), .A2(n15576), .ZN(n6646) );
  XNOR2_X1 U13853 ( .A(n13061), .B(n6647), .ZN(n12349) );
  XNOR2_X1 U13854 ( .A(n12746), .B(n6647), .ZN(n11368) );
  XNOR2_X1 U13855 ( .A(n15779), .B(n16617), .ZN(n6650) );
  NAND2_X1 U13856 ( .A1(n15402), .A2(n13639), .ZN(n13602) );
  NAND2_X1 U13857 ( .A1(n13579), .A2(n13580), .ZN(n13639) );
  XNOR2_X1 U13858 ( .A(n13481), .B(n6652), .ZN(n6651) );
  NAND2_X1 U13859 ( .A1(n17848), .A2(n17847), .ZN(n6656) );
  INV_X1 U13860 ( .A(n17269), .ZN(n16863) );
  NAND2_X1 U13861 ( .A1(n2985), .A2(n29299), .ZN(n16773) );
  INV_X1 U13862 ( .A(n12000), .ZN(n6658) );
  OAI21_X1 U13863 ( .B1(n12004), .B2(n11996), .A(n6658), .ZN(n6657) );
  INV_X1 U13864 ( .A(n12004), .ZN(n11538) );
  INV_X1 U13865 ( .A(n11755), .ZN(n6661) );
  NAND2_X1 U13866 ( .A1(n8957), .A2(n6662), .ZN(n8959) );
  OR2_X1 U13867 ( .A1(n18195), .A2(n6663), .ZN(n18103) );
  NAND2_X1 U13868 ( .A1(n10876), .A2(n29593), .ZN(n11217) );
  INV_X1 U13869 ( .A(n18774), .ZN(n19154) );
  XNOR2_X1 U13870 ( .A(n18774), .B(n1982), .ZN(n6667) );
  AND2_X1 U13872 ( .A1(n29537), .A2(n27777), .ZN(n27784) );
  INV_X1 U13873 ( .A(n15361), .ZN(n6675) );
  NOR2_X1 U13877 ( .A1(n10815), .A2(n6677), .ZN(n10565) );
  NAND2_X1 U13878 ( .A1(n11246), .A2(n12316), .ZN(n6680) );
  INV_X1 U13880 ( .A(n16797), .ZN(n17451) );
  XNOR2_X1 U13883 ( .A(n6683), .B(n13543), .ZN(n13456) );
  XNOR2_X1 U13884 ( .A(n6683), .B(n5490), .ZN(n11604) );
  XNOR2_X1 U13885 ( .A(n6683), .B(n13459), .ZN(n13296) );
  XNOR2_X1 U13886 ( .A(n6683), .B(n13133), .ZN(n12417) );
  OAI211_X1 U13887 ( .C1(n28648), .C2(n14215), .A(n14413), .B(n6466), .ZN(
        n13955) );
  NAND2_X1 U13889 ( .A1(n24020), .A2(n23126), .ZN(n24019) );
  AND2_X1 U13890 ( .A1(n24020), .A2(n2054), .ZN(n24543) );
  INV_X1 U13891 ( .A(n24020), .ZN(n6686) );
  NAND2_X1 U13892 ( .A1(n6693), .A2(n8977), .ZN(n6691) );
  NAND2_X1 U13893 ( .A1(n8978), .A2(n8976), .ZN(n6693) );
  XNOR2_X1 U13894 ( .A(n22437), .B(n22501), .ZN(n22172) );
  NAND3_X1 U13895 ( .A1(n6698), .A2(n5142), .A3(n6697), .ZN(n6695) );
  NAND2_X1 U13896 ( .A1(n20849), .A2(n21576), .ZN(n6696) );
  NAND2_X1 U13897 ( .A1(n21577), .A2(n21485), .ZN(n6697) );
  NAND2_X1 U13899 ( .A1(n17278), .A2(n539), .ZN(n16766) );
  XNOR2_X1 U13901 ( .A(n18929), .B(n19181), .ZN(n6702) );
  XNOR2_X2 U13902 ( .A(n6702), .B(n6701), .ZN(n20148) );
  NAND2_X1 U13903 ( .A1(n8427), .A2(n8351), .ZN(n7809) );
  NAND2_X1 U13904 ( .A1(n11195), .A2(n6687), .ZN(n11568) );
  XNOR2_X1 U13905 ( .A(n6708), .B(n26910), .ZN(Ciphertext[46]) );
  OR2_X1 U13906 ( .A1(n26908), .A2(n27458), .ZN(n6709) );
  OAI21_X1 U13907 ( .B1(n6712), .B2(n6711), .A(n27458), .ZN(n6710) );
  NOR2_X1 U13908 ( .A1(n28435), .A2(n29468), .ZN(n6711) );
  NAND2_X1 U13909 ( .A1(n23862), .A2(n25418), .ZN(n26151) );
  NOR2_X1 U13910 ( .A1(n17988), .A2(n17890), .ZN(n6715) );
  NAND2_X1 U13911 ( .A1(n6716), .A2(n6715), .ZN(n6714) );
  XNOR2_X1 U13912 ( .A(n20761), .B(n20760), .ZN(n23010) );
  INV_X1 U13913 ( .A(n23010), .ZN(n23657) );
  INV_X1 U13914 ( .A(n23140), .ZN(n23141) );
  XNOR2_X1 U13915 ( .A(n19015), .B(n19016), .ZN(n6717) );
  INV_X1 U13916 ( .A(n28142), .ZN(n18366) );
  XNOR2_X1 U13918 ( .A(n22363), .B(n22434), .ZN(n21620) );
  OAI21_X1 U13919 ( .B1(n11328), .B2(n10858), .A(n6721), .ZN(n6720) );
  INV_X1 U13920 ( .A(n6722), .ZN(n6721) );
  NAND2_X1 U13921 ( .A1(n26940), .A2(n26943), .ZN(n6724) );
  NAND2_X1 U13922 ( .A1(n15407), .A2(n15108), .ZN(n12371) );
  NAND2_X1 U13924 ( .A1(n17500), .A2(n6727), .ZN(n17503) );
  NOR2_X1 U13926 ( .A1(n1835), .A2(n19956), .ZN(n6729) );
  INV_X1 U13927 ( .A(n20321), .ZN(n6730) );
  NOR2_X1 U13928 ( .A1(n21248), .A2(n6730), .ZN(n21249) );
  NOR2_X1 U13929 ( .A1(n20695), .A2(n6730), .ZN(n21254) );
  OR3_X1 U13930 ( .A1(n21304), .A2(n21311), .A3(n29328), .ZN(n6731) );
  NAND2_X1 U13932 ( .A1(n6735), .A2(n27425), .ZN(n6734) );
  MUX2_X1 U13933 ( .A(n27428), .B(n27427), .S(n29542), .Z(n6735) );
  NAND2_X1 U13934 ( .A1(n26494), .A2(n29515), .ZN(n6737) );
  NAND2_X1 U13937 ( .A1(n6741), .A2(n24582), .ZN(n6740) );
  NAND2_X1 U13938 ( .A1(n11554), .A2(n6742), .ZN(n6743) );
  OAI21_X1 U13939 ( .B1(n11152), .B2(n593), .A(n6745), .ZN(n11157) );
  INV_X1 U13940 ( .A(n9146), .ZN(n6747) );
  INV_X1 U13941 ( .A(n9146), .ZN(n9150) );
  OAI211_X2 U13942 ( .C1(n4104), .C2(n6751), .A(n6750), .B(n6749), .ZN(n22619)
         );
  NAND2_X1 U13943 ( .A1(n21494), .A2(n6752), .ZN(n6751) );
  INV_X1 U13944 ( .A(n21496), .ZN(n6752) );
  XNOR2_X1 U13945 ( .A(n6753), .B(n16041), .ZN(n6754) );
  XNOR2_X1 U13946 ( .A(n6754), .B(n16042), .ZN(n16679) );
  NAND2_X1 U13947 ( .A1(n8227), .A2(n7424), .ZN(n8224) );
  NAND2_X1 U13948 ( .A1(n6756), .A2(n26995), .ZN(n6755) );
  NAND2_X1 U13949 ( .A1(n6757), .A2(n26632), .ZN(n6756) );
  INV_X1 U13950 ( .A(n26632), .ZN(n26996) );
  NAND2_X1 U13951 ( .A1(n26997), .A2(n26998), .ZN(n6757) );
  NAND2_X1 U13953 ( .A1(n6759), .A2(n14796), .ZN(n6758) );
  NAND2_X1 U13954 ( .A1(n15204), .A2(n14961), .ZN(n6759) );
  NAND2_X1 U13955 ( .A1(n14927), .A2(n14968), .ZN(n6760) );
  INV_X1 U13956 ( .A(n14961), .ZN(n14967) );
  NAND2_X1 U13957 ( .A1(n6762), .A2(n29531), .ZN(n6761) );
  INV_X1 U13958 ( .A(n21308), .ZN(n6762) );
  NAND2_X1 U13959 ( .A1(n17399), .A2(n17398), .ZN(n6765) );
  NAND2_X1 U13960 ( .A1(n14238), .A2(n14171), .ZN(n14174) );
  NAND2_X1 U13961 ( .A1(n26435), .A2(n6768), .ZN(n6767) );
  XNOR2_X1 U13962 ( .A(n22270), .B(n22418), .ZN(n22100) );
  INV_X1 U13963 ( .A(n16797), .ZN(n6772) );
  NAND2_X1 U13964 ( .A1(n6772), .A2(n17129), .ZN(n17454) );
  NAND2_X1 U13966 ( .A1(n10683), .A2(n5573), .ZN(n6777) );
  NAND2_X1 U13967 ( .A1(n10684), .A2(n6779), .ZN(n6778) );
  NOR2_X1 U13968 ( .A1(n8258), .A2(n28615), .ZN(n6783) );
  AOI22_X1 U13972 ( .A1(n8257), .A2(n6782), .B1(n28614), .B2(n28618), .ZN(
        n6785) );
  NAND2_X1 U13974 ( .A1(n24976), .A2(n23467), .ZN(n6786) );
  NAND2_X1 U13975 ( .A1(n24256), .A2(n24972), .ZN(n24012) );
  OAI21_X1 U13978 ( .B1(n26723), .B2(n26716), .A(n6790), .ZN(n25316) );
  NAND2_X1 U13979 ( .A1(n26716), .A2(n283), .ZN(n6790) );
  OAI21_X1 U13983 ( .B1(n26216), .B2(n26217), .A(n6793), .ZN(n26218) );
  INV_X1 U13984 ( .A(n26723), .ZN(n6793) );
  XNOR2_X2 U13985 ( .A(n6795), .B(n9623), .ZN(n11045) );
  XNOR2_X1 U13986 ( .A(n29509), .B(n6796), .ZN(n6795) );
  NAND2_X1 U13987 ( .A1(n17453), .A2(n28193), .ZN(n6799) );
  OAI21_X1 U13988 ( .B1(n1814), .B2(n21459), .A(n6803), .ZN(n21570) );
  XNOR2_X1 U13989 ( .A(n19724), .B(n19723), .ZN(n6804) );
  MUX2_X1 U13991 ( .A(n20440), .B(n20609), .S(n20437), .Z(n19886) );
  AOI22_X1 U13993 ( .A1(n27372), .A2(n27366), .B1(n25360), .B2(n25359), .ZN(
        n6806) );
  NOR2_X1 U13994 ( .A1(n295), .A2(n28394), .ZN(n27376) );
  OAI21_X1 U13995 ( .B1(n27212), .B2(n27382), .A(n6808), .ZN(n6810) );
  NAND2_X1 U13996 ( .A1(n6809), .A2(n5313), .ZN(n6808) );
  NOR2_X1 U13997 ( .A1(n27214), .A2(n6810), .ZN(n27215) );
  OAI211_X1 U13998 ( .C1(n524), .C2(n17771), .A(n18254), .B(n18252), .ZN(n6811) );
  NAND2_X1 U13999 ( .A1(n11867), .A2(n11869), .ZN(n11462) );
  NOR2_X1 U14002 ( .A1(n6814), .A2(n333), .ZN(n10568) );
  INV_X1 U14003 ( .A(n10797), .ZN(n6814) );
  NAND2_X1 U14004 ( .A1(n11227), .A2(n11225), .ZN(n6815) );
  NAND2_X1 U14005 ( .A1(n11232), .A2(n6816), .ZN(n11894) );
  XNOR2_X1 U14006 ( .A(n6817), .B(n22238), .ZN(n22244) );
  INV_X1 U14007 ( .A(n22748), .ZN(n6817) );
  XNOR2_X1 U14008 ( .A(n22238), .B(n6818), .ZN(n22907) );
  XNOR2_X1 U14009 ( .A(n13221), .B(n13220), .ZN(n6820) );
  XNOR2_X2 U14010 ( .A(n6820), .B(n6819), .ZN(n14045) );
  NAND2_X1 U14011 ( .A1(n23644), .A2(n23180), .ZN(n6822) );
  NAND2_X1 U14012 ( .A1(n6827), .A2(n26793), .ZN(n6823) );
  NAND2_X1 U14013 ( .A1(n25419), .A2(n6826), .ZN(n6825) );
  INV_X1 U14014 ( .A(n26793), .ZN(n6826) );
  NAND2_X1 U14015 ( .A1(n26792), .A2(n26789), .ZN(n6827) );
  INV_X1 U14016 ( .A(n16973), .ZN(n6829) );
  INV_X1 U14017 ( .A(n12955), .ZN(n12514) );
  INV_X1 U14018 ( .A(n13014), .ZN(n13524) );
  XNOR2_X1 U14019 ( .A(n6831), .B(n13014), .ZN(n13442) );
  INV_X1 U14020 ( .A(n20495), .ZN(n6834) );
  INV_X1 U14021 ( .A(n20494), .ZN(n20218) );
  NAND2_X1 U14022 ( .A1(n6841), .A2(n6838), .ZN(n21251) );
  NAND2_X1 U14023 ( .A1(n19506), .A2(n6843), .ZN(n6841) );
  OAI22_X2 U14024 ( .A1(n6841), .A2(n21248), .B1(n6839), .B2(n6842), .ZN(
        n21809) );
  NAND2_X1 U14025 ( .A1(n21251), .A2(n6840), .ZN(n21807) );
  NAND4_X1 U14026 ( .A1(n27500), .A2(n27499), .A3(n6845), .A4(n6844), .ZN(
        n27501) );
  NAND3_X1 U14027 ( .A1(n27487), .A2(n29093), .A3(n27496), .ZN(n6844) );
  NAND2_X1 U14028 ( .A1(n27495), .A2(n29093), .ZN(n6845) );
  NAND3_X1 U14029 ( .A1(n5811), .A2(n14969), .A3(n13789), .ZN(n13788) );
  XNOR2_X1 U14030 ( .A(n22495), .B(n22497), .ZN(n6846) );
  XNOR2_X1 U14031 ( .A(n22498), .B(n22496), .ZN(n6847) );
  NAND2_X1 U14032 ( .A1(n6850), .A2(n12257), .ZN(n6849) );
  NAND2_X1 U14033 ( .A1(n6855), .A2(n6853), .ZN(n6852) );
  NAND2_X1 U14034 ( .A1(n14943), .A2(n14944), .ZN(n6855) );
  NAND2_X1 U14035 ( .A1(n25506), .A2(n25505), .ZN(n27054) );
  XNOR2_X1 U14036 ( .A(n6858), .B(n26604), .ZN(Ciphertext[177]) );
  NAND2_X1 U14037 ( .A1(n9028), .A2(n9030), .ZN(n7715) );
  NOR2_X1 U14038 ( .A1(n6636), .A2(n21465), .ZN(n20755) );
  NOR2_X1 U14039 ( .A1(n28155), .A2(n29236), .ZN(n6861) );
  INV_X1 U14041 ( .A(n20277), .ZN(n22041) );
  INV_X1 U14042 ( .A(n24631), .ZN(n6867) );
  NOR2_X1 U14043 ( .A1(n6866), .A2(n6867), .ZN(n6864) );
  NOR2_X1 U14044 ( .A1(n4366), .A2(n24532), .ZN(n6866) );
  XNOR2_X1 U14045 ( .A(n13133), .B(n12768), .ZN(n13325) );
  INV_X1 U14046 ( .A(n14351), .ZN(n13825) );
  NOR2_X1 U14047 ( .A1(n13826), .A2(n14351), .ZN(n6872) );
  NAND2_X1 U14048 ( .A1(n596), .A2(n8642), .ZN(n6875) );
  MUX2_X1 U14049 ( .A(n23849), .B(n23721), .S(n23726), .Z(n22956) );
  NAND2_X1 U14050 ( .A1(n23723), .A2(n29157), .ZN(n23731) );
  NAND3_X1 U14051 ( .A1(n6880), .A2(n6878), .A3(n6877), .ZN(n15940) );
  NAND3_X1 U14052 ( .A1(n6879), .A2(n3784), .A3(n426), .ZN(n6878) );
  INV_X1 U14053 ( .A(n15371), .ZN(n6879) );
  NAND3_X1 U14054 ( .A1(n20628), .A2(n20334), .A3(n20258), .ZN(n6882) );
  NAND2_X1 U14055 ( .A1(n6884), .A2(n28186), .ZN(n6881) );
  AND2_X1 U14056 ( .A1(n20625), .A2(n20626), .ZN(n6884) );
  XNOR2_X1 U14057 ( .A(n19322), .B(n6886), .ZN(n19326) );
  XNOR2_X1 U14058 ( .A(n19320), .B(n19321), .ZN(n6886) );
  NAND2_X1 U14059 ( .A1(n26168), .A2(n29610), .ZN(n6887) );
  NAND3_X1 U14060 ( .A1(n4751), .A2(n26914), .A3(n1872), .ZN(n6888) );
  NAND2_X1 U14061 ( .A1(n17518), .A2(n17106), .ZN(n6889) );
  XNOR2_X1 U14062 ( .A(n10303), .B(n1983), .ZN(n6891) );
  XNOR2_X1 U14064 ( .A(n13322), .B(n2025), .ZN(n6895) );
  NOR2_X1 U14065 ( .A1(n14310), .A2(n14309), .ZN(n14311) );
  NAND3_X2 U14066 ( .A1(n10979), .A2(n10978), .A3(n6896), .ZN(n12252) );
  INV_X1 U14067 ( .A(n12252), .ZN(n11933) );
  XNOR2_X1 U14068 ( .A(n12522), .B(n13434), .ZN(n12526) );
  XNOR2_X1 U14069 ( .A(n25178), .B(n25177), .ZN(n26374) );
  OR2_X1 U14070 ( .A1(n1030), .A2(n26380), .ZN(n26430) );
  AOI21_X1 U14071 ( .B1(n26991), .B2(n25770), .A(n25769), .ZN(n26537) );
  OR2_X1 U14072 ( .A1(n26254), .A2(n28053), .ZN(n26255) );
  BUF_X1 U14075 ( .A(n12762), .Z(n12735) );
  OAI211_X1 U14076 ( .C1(n28012), .C2(n443), .A(n28011), .B(n28010), .ZN(
        n28014) );
  OR2_X1 U14078 ( .A1(n29036), .A2(n28601), .ZN(n12796) );
  INV_X1 U14079 ( .A(n15738), .ZN(n16483) );
  XNOR2_X2 U14080 ( .A(n25085), .B(n25084), .ZN(n26917) );
  MUX2_X2 U14081 ( .A(n26916), .B(n26915), .S(n26914), .Z(n27531) );
  OR2_X1 U14082 ( .A1(n25957), .A2(n27357), .ZN(n25671) );
  OR2_X1 U14083 ( .A1(n25997), .A2(n28562), .ZN(n26002) );
  AOI22_X1 U14084 ( .A1(n27091), .A2(n27090), .B1(n27089), .B2(n27088), .ZN(
        n27271) );
  NAND2_X1 U14085 ( .A1(n23949), .A2(n23948), .ZN(n25922) );
  OAI22_X1 U14086 ( .A1(n28003), .A2(n28019), .B1(n28001), .B2(n28015), .ZN(
        n28022) );
  NOR2_X1 U14087 ( .A1(n17729), .A2(n18456), .ZN(n17731) );
  OR2_X1 U14088 ( .A1(n24556), .A2(n24551), .ZN(n24175) );
  AND3_X1 U14089 ( .A1(n27521), .A2(n27527), .A3(n27520), .ZN(n27522) );
  AND2_X1 U14091 ( .A1(n27843), .A2(n27101), .ZN(n27099) );
  NOR2_X1 U14092 ( .A1(n23906), .A2(n24373), .ZN(n24377) );
  AND2_X1 U14093 ( .A1(n13844), .A2(n15456), .ZN(n13845) );
  OR2_X1 U14094 ( .A1(n22451), .A2(n23387), .ZN(n23222) );
  OR2_X1 U14095 ( .A1(n21591), .A2(n21322), .ZN(n21323) );
  AND2_X1 U14096 ( .A1(n24427), .A2(n28531), .ZN(n24428) );
  AND2_X1 U14097 ( .A1(n25660), .A2(n26721), .ZN(n26217) );
  NOR2_X2 U14101 ( .A1(n23910), .A2(n23909), .ZN(n25375) );
  XNOR2_X1 U14102 ( .A(n25248), .B(n25830), .ZN(n26754) );
  OR2_X1 U14103 ( .A1(n14215), .A2(n13686), .ZN(n14419) );
  AND2_X1 U14104 ( .A1(n27562), .A2(n27551), .ZN(n27149) );
  OR2_X1 U14105 ( .A1(n27101), .A2(n27100), .ZN(n27248) );
  AOI21_X1 U14106 ( .B1(n27637), .B2(n26980), .A(n26672), .ZN(n26675) );
  OR2_X1 U14108 ( .A1(n339), .A2(n23776), .ZN(n23780) );
  XNOR2_X2 U14109 ( .A(n25326), .B(n25327), .ZN(n26204) );
  XNOR2_X2 U14110 ( .A(n7137), .B(Key[53]), .ZN(n8014) );
  INV_X1 U14112 ( .A(n27638), .ZN(n27637) );
  INV_X1 U14114 ( .A(n26933), .ZN(n24788) );
  AND2_X1 U14115 ( .A1(n24390), .A2(n24391), .ZN(n23900) );
  OAI21_X1 U14116 ( .B1(n24364), .B2(n28592), .A(n24363), .ZN(n26705) );
  NOR2_X1 U14117 ( .A1(n449), .A2(n29468), .ZN(n26605) );
  XNOR2_X1 U14118 ( .A(n22511), .B(n22510), .ZN(n22512) );
  OR2_X1 U14119 ( .A1(n20444), .A2(n415), .ZN(n19505) );
  XNOR2_X1 U14121 ( .A(n25507), .B(n25210), .ZN(n25212) );
  INV_X1 U14122 ( .A(n24858), .ZN(n25848) );
  XNOR2_X1 U14126 ( .A(n25351), .B(n25352), .ZN(n26077) );
  XNOR2_X2 U14127 ( .A(n16188), .B(n16187), .ZN(n17467) );
  OAI21_X1 U14128 ( .B1(n26159), .B2(n26457), .A(n25616), .ZN(n25633) );
  NOR2_X2 U14132 ( .A1(n17538), .A2(n17537), .ZN(n19555) );
  OAI211_X2 U14133 ( .C1(n18445), .C2(n18185), .A(n18184), .B(n18183), .ZN(
        n19397) );
  OR2_X1 U14134 ( .A1(n28524), .A2(n24716), .ZN(n24353) );
  AND2_X1 U14136 ( .A1(n9194), .A2(n329), .ZN(n6897) );
  XOR2_X1 U14137 ( .A(n10248), .B(n10247), .Z(n6898) );
  OR2_X1 U14138 ( .A1(n17561), .A2(n17560), .ZN(n6899) );
  OR3_X1 U14139 ( .A1(n17402), .A2(n29572), .A3(n17400), .ZN(n6900) );
  AND2_X1 U14140 ( .A1(n8381), .A2(n8384), .ZN(n6901) );
  OR2_X1 U14141 ( .A1(n29314), .A2(n1930), .ZN(n6904) );
  OR2_X1 U14142 ( .A1(n7626), .A2(n8217), .ZN(n6905) );
  AND2_X1 U14143 ( .A1(n2209), .A2(n29643), .ZN(n6906) );
  AND2_X1 U14144 ( .A1(n27859), .A2(n27847), .ZN(n6907) );
  OR2_X1 U14145 ( .A1(n8487), .A2(n8486), .ZN(n6908) );
  AOI21_X1 U14146 ( .B1(n25975), .B2(n26236), .A(n25974), .ZN(n28009) );
  AND2_X1 U14148 ( .A1(n8384), .A2(n8729), .ZN(n6909) );
  AND2_X1 U14149 ( .A1(n5425), .A2(n26880), .ZN(n6910) );
  AND2_X1 U14150 ( .A1(n21292), .A2(n20726), .ZN(n6911) );
  NAND2_X1 U14152 ( .A1(n26274), .A2(n26273), .ZN(n27582) );
  INV_X1 U14153 ( .A(n27582), .ZN(n26346) );
  INV_X1 U14154 ( .A(n2274), .ZN(n22755) );
  AND2_X1 U14155 ( .A1(n9033), .A2(n9032), .ZN(n6915) );
  AND2_X1 U14156 ( .A1(n11723), .A2(n11722), .ZN(n6917) );
  AND2_X1 U14157 ( .A1(n10761), .A2(n11119), .ZN(n6918) );
  OR2_X1 U14158 ( .A1(n12339), .A2(n12338), .ZN(n6919) );
  AND2_X1 U14159 ( .A1(n12049), .A2(n12050), .ZN(n6920) );
  OR2_X1 U14160 ( .A1(n14233), .A2(n14593), .ZN(n6921) );
  XOR2_X1 U14161 ( .A(n13099), .B(n13098), .Z(n6922) );
  XOR2_X1 U14162 ( .A(n12570), .B(n12569), .Z(n6923) );
  INV_X1 U14163 ( .A(n15420), .ZN(n15422) );
  OR2_X1 U14164 ( .A1(n17264), .A2(n16996), .ZN(n6926) );
  AND3_X2 U14165 ( .A1(n16998), .A2(n16997), .A3(n6926), .ZN(n6927) );
  AND2_X1 U14166 ( .A1(n16884), .A2(n16883), .ZN(n6928) );
  XOR2_X1 U14167 ( .A(n15563), .B(n15562), .Z(n6929) );
  AND2_X1 U14168 ( .A1(n17637), .A2(n17636), .ZN(n6930) );
  XNOR2_X1 U14170 ( .A(n18617), .B(n18616), .ZN(n20568) );
  OR2_X1 U14171 ( .A1(n20567), .A2(n20573), .ZN(n6932) );
  AND2_X1 U14172 ( .A1(n21412), .A2(n20663), .ZN(n6933) );
  AND2_X1 U14173 ( .A1(n20201), .A2(n20200), .ZN(n6935) );
  OR2_X1 U14174 ( .A1(n21500), .A2(n21192), .ZN(n6936) );
  AND2_X1 U14175 ( .A1(n20118), .A2(n21424), .ZN(n6937) );
  XOR2_X1 U14176 ( .A(n22591), .B(n22590), .Z(n6938) );
  XOR2_X1 U14177 ( .A(n22666), .B(n22665), .Z(n6939) );
  OR2_X1 U14178 ( .A1(n22402), .A2(n22401), .ZN(n6940) );
  AND2_X1 U14179 ( .A1(n23145), .A2(n23461), .ZN(n6941) );
  XNOR2_X1 U14180 ( .A(n17752), .B(n17751), .ZN(n20412) );
  OR2_X1 U14182 ( .A1(n1955), .A2(n28512), .ZN(n6943) );
  OR2_X1 U14183 ( .A1(n24672), .A2(n28635), .ZN(n6944) );
  OR3_X1 U14184 ( .A1(n24347), .A2(n24437), .A3(n24433), .ZN(n6945) );
  OR2_X1 U14185 ( .A1(n24806), .A2(n24261), .ZN(n6946) );
  XOR2_X1 U14186 ( .A(n25414), .B(n25413), .Z(n6947) );
  AND2_X1 U14187 ( .A1(n6768), .A2(n26940), .ZN(n6948) );
  AND2_X1 U14188 ( .A1(n27852), .A2(n27854), .ZN(n6949) );
  OR2_X1 U14189 ( .A1(n5505), .A2(n26933), .ZN(n6950) );
  OR2_X1 U14190 ( .A1(n27118), .A2(n26835), .ZN(n6951) );
  OR2_X1 U14191 ( .A1(n26146), .A2(n325), .ZN(n6952) );
  AND2_X1 U14192 ( .A1(n326), .A2(n26126), .ZN(n6953) );
  OR3_X1 U14193 ( .A1(n27855), .A2(n26641), .A3(n27847), .ZN(n6954) );
  AND2_X1 U14194 ( .A1(n28021), .A2(n28003), .ZN(n6955) );
  AND2_X1 U14195 ( .A1(n14230), .A2(n14101), .ZN(n6956) );
  OR2_X1 U14196 ( .A1(n7759), .A2(n8176), .ZN(n7345) );
  OR2_X1 U14197 ( .A1(n7958), .A2(n7589), .ZN(n7590) );
  INV_X1 U14198 ( .A(n8161), .ZN(n8166) );
  INV_X1 U14199 ( .A(Plaintext[159]), .ZN(n7049) );
  OR2_X1 U14200 ( .A1(n8270), .A2(n8267), .ZN(n7211) );
  OR2_X1 U14201 ( .A1(n8280), .A2(n8275), .ZN(n7407) );
  BUF_X1 U14202 ( .A(n7069), .Z(n7582) );
  XNOR2_X1 U14203 ( .A(Key[125]), .B(Plaintext[125]), .ZN(n8290) );
  OR2_X1 U14204 ( .A1(n8336), .A2(n8886), .ZN(n8007) );
  INV_X1 U14205 ( .A(n8462), .ZN(n7445) );
  OR2_X1 U14206 ( .A1(n7618), .A2(n8256), .ZN(n7389) );
  INV_X1 U14207 ( .A(Plaintext[167]), .ZN(n7058) );
  OR2_X1 U14208 ( .A1(n7763), .A2(n613), .ZN(n7764) );
  OR2_X1 U14209 ( .A1(n8300), .A2(n7400), .ZN(n7940) );
  INV_X1 U14210 ( .A(n29081), .ZN(n8002) );
  INV_X1 U14211 ( .A(n8397), .ZN(n8864) );
  INV_X1 U14212 ( .A(n8873), .ZN(n8876) );
  OR2_X1 U14213 ( .A1(n8917), .A2(n9108), .ZN(n8915) );
  OR2_X1 U14214 ( .A1(n8955), .A2(n8801), .ZN(n9162) );
  AOI22_X1 U14215 ( .A1(n7720), .A2(n8049), .B1(n7719), .B2(n7718), .ZN(n7726)
         );
  INV_X1 U14216 ( .A(n9060), .ZN(n8866) );
  INV_X1 U14217 ( .A(n9562), .ZN(n8765) );
  OR2_X1 U14218 ( .A1(n8549), .A2(n7410), .ZN(n7412) );
  OR2_X1 U14219 ( .A1(n9060), .A2(n8872), .ZN(n8395) );
  OR2_X1 U14220 ( .A1(n9582), .A2(n1196), .ZN(n9583) );
  OR2_X1 U14221 ( .A1(n8965), .A2(n8963), .ZN(n8640) );
  INV_X1 U14222 ( .A(n8763), .ZN(n8945) );
  INV_X1 U14223 ( .A(n8608), .ZN(n9529) );
  INV_X1 U14224 ( .A(n10956), .ZN(n9858) );
  XNOR2_X1 U14225 ( .A(n10271), .B(n10350), .ZN(n9849) );
  OAI211_X1 U14226 ( .C1(n9160), .C2(n8625), .A(n8624), .B(n8804), .ZN(n9306)
         );
  XNOR2_X1 U14227 ( .A(n9838), .B(n9495), .ZN(n9496) );
  INV_X1 U14228 ( .A(n9701), .ZN(n9666) );
  XNOR2_X1 U14229 ( .A(n10249), .B(n6898), .ZN(n10534) );
  XNOR2_X1 U14230 ( .A(n10175), .B(n10174), .ZN(n11067) );
  XNOR2_X1 U14231 ( .A(n7571), .B(n7570), .ZN(n7572) );
  OR2_X1 U14232 ( .A1(n11223), .A2(n29593), .ZN(n10660) );
  XNOR2_X1 U14233 ( .A(n9336), .B(n9780), .ZN(n9337) );
  NOR2_X1 U14234 ( .A1(n9860), .A2(n9859), .ZN(n9861) );
  AND2_X1 U14237 ( .A1(n11147), .A2(n10742), .ZN(n11148) );
  BUF_X1 U14238 ( .A(n10518), .Z(n11027) );
  XNOR2_X1 U14239 ( .A(n10299), .B(n10417), .ZN(n10301) );
  XNOR2_X1 U14240 ( .A(n10279), .B(n10278), .ZN(n11223) );
  XNOR2_X1 U14241 ( .A(n9337), .B(n9338), .ZN(n10912) );
  XNOR2_X1 U14242 ( .A(n8090), .B(n8089), .ZN(n10820) );
  AOI21_X1 U14243 ( .B1(n10807), .B2(n11149), .A(n11148), .ZN(n11419) );
  OR2_X1 U14244 ( .A1(n11039), .A2(n28612), .ZN(n11040) );
  OAI21_X1 U14245 ( .B1(n10894), .B2(n10893), .A(n10892), .ZN(n11660) );
  INV_X1 U14246 ( .A(n11739), .ZN(n11908) );
  NOR2_X1 U14247 ( .A1(n11940), .A2(n12517), .ZN(n12579) );
  INV_X1 U14248 ( .A(n12188), .ZN(n12192) );
  OR2_X1 U14249 ( .A1(n10908), .A2(n11927), .ZN(n10909) );
  AND2_X1 U14250 ( .A1(n12022), .A2(n12354), .ZN(n12429) );
  OR2_X1 U14251 ( .A1(n11395), .A2(n11951), .ZN(n11396) );
  AOI22_X1 U14252 ( .A1(n10782), .A2(n9858), .B1(n10781), .B2(n10780), .ZN(
        n10793) );
  OAI21_X1 U14253 ( .B1(n12100), .B2(n12099), .A(n12098), .ZN(n12101) );
  OAI21_X1 U14254 ( .B1(n12579), .B2(n12575), .A(n11591), .ZN(n11592) );
  AOI21_X1 U14255 ( .B1(n10645), .B2(n12219), .A(n10644), .ZN(n12608) );
  INV_X1 U14256 ( .A(n13012), .ZN(n13013) );
  OR2_X1 U14258 ( .A1(n11655), .A2(n11378), .ZN(n11379) );
  INV_X1 U14259 ( .A(n14830), .ZN(n14831) );
  AND2_X1 U14260 ( .A1(n14400), .A2(n14399), .ZN(n14403) );
  XNOR2_X1 U14261 ( .A(n12904), .B(n12298), .ZN(n11734) );
  OR2_X1 U14263 ( .A1(n14264), .A2(n14259), .ZN(n13762) );
  INV_X1 U14264 ( .A(n14287), .ZN(n14085) );
  XNOR2_X1 U14265 ( .A(n13520), .B(n12634), .ZN(n12635) );
  XNOR2_X1 U14266 ( .A(n13241), .B(n13242), .ZN(n14046) );
  XNOR2_X1 U14267 ( .A(n10444), .B(n10443), .ZN(n13606) );
  INV_X1 U14268 ( .A(n14314), .ZN(n13884) );
  XNOR2_X1 U14269 ( .A(n12386), .B(n12387), .ZN(n14407) );
  AND2_X1 U14270 ( .A1(n13629), .A2(n13628), .ZN(n13630) );
  OR2_X1 U14271 ( .A1(n14298), .A2(n13803), .ZN(n13658) );
  OR2_X1 U14272 ( .A1(n15127), .A2(n15001), .ZN(n14999) );
  INV_X1 U14273 ( .A(n15000), .ZN(n13632) );
  AND2_X1 U14275 ( .A1(n14563), .A2(n15083), .ZN(n14670) );
  INV_X1 U14277 ( .A(n14706), .ZN(n14431) );
  AND2_X1 U14279 ( .A1(n13632), .A2(n15123), .ZN(n14686) );
  OR2_X1 U14280 ( .A1(n14874), .A2(n15071), .ZN(n14876) );
  INV_X1 U14281 ( .A(n15015), .ZN(n15327) );
  AND2_X1 U14282 ( .A1(n17474), .A2(n17124), .ZN(n17480) );
  XNOR2_X1 U14283 ( .A(n16638), .B(n16637), .ZN(n16724) );
  BUF_X1 U14284 ( .A(n16477), .Z(n15777) );
  XNOR2_X1 U14286 ( .A(n15771), .B(n15770), .ZN(n15776) );
  XNOR2_X1 U14287 ( .A(n16218), .B(n16145), .ZN(n15820) );
  INV_X1 U14288 ( .A(n17350), .ZN(n17351) );
  INV_X1 U14289 ( .A(n18124), .ZN(n18125) );
  OR2_X1 U14290 ( .A1(n18513), .A2(n18516), .ZN(n18514) );
  INV_X1 U14291 ( .A(n18707), .ZN(n17980) );
  OR2_X1 U14292 ( .A1(n16726), .A2(n16725), .ZN(n16727) );
  XNOR2_X1 U14293 ( .A(n16350), .B(n16349), .ZN(n16712) );
  OAI211_X1 U14295 ( .C1(n17217), .C2(n16940), .A(n15809), .B(n15808), .ZN(
        n15810) );
  AND2_X1 U14296 ( .A1(n18042), .A2(n18422), .ZN(n17822) );
  INV_X1 U14297 ( .A(n18433), .ZN(n18149) );
  INV_X1 U14298 ( .A(n18314), .ZN(n16442) );
  INV_X1 U14299 ( .A(n18528), .ZN(n17699) );
  AND2_X1 U14300 ( .A1(n18261), .A2(n18262), .ZN(n17896) );
  INV_X1 U14301 ( .A(n17353), .ZN(n18706) );
  AND2_X1 U14302 ( .A1(n18190), .A2(n19562), .ZN(n17796) );
  NOR2_X1 U14304 ( .A1(n17775), .A2(n17774), .ZN(n17776) );
  NOR2_X1 U14305 ( .A1(n17703), .A2(n17702), .ZN(n17704) );
  XNOR2_X1 U14307 ( .A(n19718), .B(n3423), .ZN(n19180) );
  XNOR2_X1 U14308 ( .A(n19413), .B(n19412), .ZN(n19624) );
  OR2_X1 U14309 ( .A1(n20480), .A2(n20475), .ZN(n20355) );
  XNOR2_X1 U14310 ( .A(n17630), .B(n17631), .ZN(n17687) );
  XNOR2_X1 U14311 ( .A(n19074), .B(n19073), .ZN(n19093) );
  AND2_X1 U14312 ( .A1(n28140), .A2(n20413), .ZN(n20583) );
  XNOR2_X1 U14313 ( .A(n19444), .B(n19443), .ZN(n19795) );
  AND2_X1 U14314 ( .A1(n20157), .A2(n20159), .ZN(n19983) );
  INV_X1 U14315 ( .A(n21653), .ZN(n21012) );
  XNOR2_X1 U14317 ( .A(n18905), .B(n18904), .ZN(n19766) );
  XNOR2_X1 U14318 ( .A(n19239), .B(n19238), .ZN(n20013) );
  XNOR2_X1 U14319 ( .A(n18686), .B(n18685), .ZN(n18699) );
  NAND2_X1 U14320 ( .A1(n19950), .A2(n20314), .ZN(n19951) );
  INV_X1 U14321 ( .A(n21429), .ZN(n22397) );
  OR2_X1 U14323 ( .A1(n21435), .A2(n20339), .ZN(n20011) );
  OAI21_X1 U14324 ( .B1(n20392), .B2(n20545), .A(n20391), .ZN(n20393) );
  OR2_X1 U14325 ( .A1(n21401), .A2(n20658), .ZN(n21043) );
  AND2_X1 U14326 ( .A1(n20857), .A2(n21156), .ZN(n20527) );
  OAI22_X1 U14327 ( .A1(n20622), .A2(n20621), .B1(n20620), .B2(n20619), .ZN(
        n20722) );
  AND2_X1 U14328 ( .A1(n20241), .A2(n29527), .ZN(n19792) );
  INV_X1 U14329 ( .A(n21014), .ZN(n21664) );
  OAI211_X1 U14330 ( .C1(n20205), .C2(n20307), .A(n20204), .B(n20203), .ZN(
        n20207) );
  OR2_X1 U14331 ( .A1(n21347), .A2(n28440), .ZN(n21344) );
  XNOR2_X1 U14332 ( .A(n22677), .B(n5513), .ZN(n22680) );
  AND2_X1 U14333 ( .A1(n20951), .A2(n20184), .ZN(n20185) );
  INV_X1 U14334 ( .A(n21286), .ZN(n21297) );
  AOI21_X1 U14335 ( .B1(n3763), .B2(n21307), .A(n20772), .ZN(n20773) );
  AND2_X1 U14336 ( .A1(n21194), .A2(n21500), .ZN(n21195) );
  OR2_X1 U14337 ( .A1(n22404), .A2(n22398), .ZN(n20276) );
  INV_X1 U14338 ( .A(n28327), .ZN(n22534) );
  INV_X1 U14339 ( .A(n22677), .ZN(n22556) );
  OR2_X1 U14341 ( .A1(n23245), .A2(n23246), .ZN(n22984) );
  XNOR2_X1 U14342 ( .A(n22697), .B(n22879), .ZN(n22468) );
  XNOR2_X1 U14343 ( .A(n22615), .B(n22656), .ZN(n22350) );
  OR2_X1 U14344 ( .A1(n23456), .A2(n23148), .ZN(n23149) );
  AND2_X1 U14345 ( .A1(n23416), .A2(n23419), .ZN(n23098) );
  XNOR2_X1 U14346 ( .A(n22157), .B(n20470), .ZN(n20471) );
  XNOR2_X1 U14347 ( .A(n21937), .B(n22500), .ZN(n22205) );
  XNOR2_X1 U14348 ( .A(n22468), .B(n22467), .ZN(n22471) );
  XNOR2_X1 U14349 ( .A(n22478), .B(n22477), .ZN(n22494) );
  XNOR2_X1 U14350 ( .A(n22654), .B(n22653), .ZN(n23102) );
  XNOR2_X1 U14351 ( .A(n21546), .B(n21545), .ZN(n21559) );
  OR2_X1 U14352 ( .A1(n23427), .A2(n1873), .ZN(n23341) );
  XNOR2_X1 U14353 ( .A(n21852), .B(n21851), .ZN(n23156) );
  INV_X1 U14354 ( .A(n24502), .ZN(n24503) );
  XNOR2_X1 U14355 ( .A(n21341), .B(n21340), .ZN(n23422) );
  BUF_X1 U14357 ( .A(n22284), .Z(n23558) );
  AND2_X1 U14358 ( .A1(n23727), .A2(n23726), .ZN(n23728) );
  XNOR2_X1 U14359 ( .A(n22512), .B(n22513), .ZN(n23077) );
  OR2_X1 U14360 ( .A1(n24682), .A2(n24688), .ZN(n24311) );
  OR2_X1 U14363 ( .A1(n24891), .A2(n24631), .ZN(n24297) );
  NOR2_X1 U14364 ( .A1(n23036), .A2(n23482), .ZN(n23486) );
  OR2_X1 U14365 ( .A1(n21898), .A2(n23662), .ZN(n21724) );
  INV_X1 U14366 ( .A(n24600), .ZN(n24607) );
  NOR2_X1 U14367 ( .A1(n23729), .A2(n23728), .ZN(n23730) );
  AND2_X1 U14368 ( .A1(n404), .A2(n24678), .ZN(n24067) );
  AND2_X1 U14369 ( .A1(n29050), .A2(n24603), .ZN(n24285) );
  OR2_X1 U14371 ( .A1(n1883), .A2(n23378), .ZN(n23379) );
  AND2_X1 U14372 ( .A1(n24772), .A2(n24766), .ZN(n24774) );
  AND2_X1 U14373 ( .A1(n26240), .A2(n26761), .ZN(n25602) );
  AND2_X1 U14374 ( .A1(n26450), .A2(n26449), .ZN(n26451) );
  AOI21_X1 U14375 ( .B1(n26427), .B2(n26426), .A(n26425), .ZN(n26428) );
  XNOR2_X1 U14376 ( .A(n25138), .B(n25137), .ZN(n26436) );
  XNOR2_X1 U14377 ( .A(n26008), .B(n24955), .ZN(n24958) );
  INV_X1 U14378 ( .A(n25270), .ZN(n25056) );
  XNOR2_X1 U14379 ( .A(n25886), .B(n1225), .ZN(n25557) );
  OR2_X1 U14380 ( .A1(n28660), .A2(n27069), .ZN(n25963) );
  INV_X1 U14382 ( .A(n26240), .ZN(n25603) );
  OR2_X1 U14383 ( .A1(n26194), .A2(n26191), .ZN(n25240) );
  AND2_X1 U14384 ( .A1(n26949), .A2(n26266), .ZN(n26267) );
  XNOR2_X1 U14385 ( .A(n24882), .B(n24881), .ZN(n26263) );
  XNOR2_X1 U14386 ( .A(n26007), .B(n26008), .ZN(n26009) );
  XNOR2_X1 U14387 ( .A(n26077), .B(n26076), .ZN(n26078) );
  NOR2_X1 U14389 ( .A1(n26748), .A2(n25453), .ZN(n25461) );
  XNOR2_X1 U14390 ( .A(n25229), .B(n25228), .ZN(n26729) );
  OR2_X1 U14392 ( .A1(n28561), .A2(n28525), .ZN(n24200) );
  XNOR2_X1 U14393 ( .A(n25917), .B(n25918), .ZN(n26850) );
  AOI21_X1 U14394 ( .B1(n29482), .B2(n26998), .A(n26995), .ZN(n25972) );
  OR2_X1 U14395 ( .A1(n27388), .A2(n27402), .ZN(n25627) );
  AND3_X1 U14396 ( .A1(n24202), .A2(n24201), .A3(n24200), .ZN(n24203) );
  INV_X1 U14397 ( .A(n27282), .ZN(n27278) );
  NAND2_X1 U14398 ( .A1(n26434), .A2(n26433), .ZN(n26880) );
  AND2_X1 U14399 ( .A1(n26846), .A2(n27827), .ZN(n26902) );
  INV_X1 U14400 ( .A(n27852), .ZN(n27847) );
  AND2_X1 U14401 ( .A1(n27872), .A2(n27865), .ZN(n25897) );
  OR2_X1 U14402 ( .A1(n26984), .A2(n28001), .ZN(n28002) );
  BUF_X1 U14403 ( .A(n28009), .Z(n28003) );
  OR2_X1 U14404 ( .A1(n25957), .A2(n27328), .ZN(n25958) );
  OR2_X1 U14405 ( .A1(n26816), .A2(n24826), .ZN(n24827) );
  AOI22_X1 U14407 ( .A1(n26809), .A2(n25997), .B1(n25995), .B2(n27363), .ZN(
        n25996) );
  AND3_X1 U14408 ( .A1(n27615), .A2(n26973), .A3(n3154), .ZN(n27624) );
  INV_X1 U14409 ( .A(n25991), .ZN(n25992) );
  INV_X1 U14410 ( .A(Plaintext[113]), .ZN(n6957) );
  XNOR2_X1 U14411 ( .A(n6957), .B(Key[113]), .ZN(n6958) );
  XNOR2_X1 U14413 ( .A(Key[109]), .B(Plaintext[109]), .ZN(n7924) );
  NAND2_X1 U14414 ( .A1(n8214), .A2(n626), .ZN(n6963) );
  INV_X1 U14415 ( .A(n8216), .ZN(n7437) );
  OAI21_X1 U14416 ( .B1(n7437), .B2(n7626), .A(n7924), .ZN(n6962) );
  OAI21_X1 U14419 ( .B1(n8216), .B2(n8213), .A(n7625), .ZN(n6960) );
  INV_X1 U14420 ( .A(Plaintext[114]), .ZN(n6964) );
  XNOR2_X1 U14421 ( .A(n6964), .B(Key[114]), .ZN(n7613) );
  INV_X1 U14422 ( .A(n7614), .ZN(n7932) );
  INV_X1 U14424 ( .A(n7933), .ZN(n8308) );
  NAND2_X1 U14425 ( .A1(n8308), .A2(n7935), .ZN(n6965) );
  MUX2_X1 U14426 ( .A(n8310), .B(n6965), .S(n29135), .Z(n6967) );
  XNOR2_X1 U14427 ( .A(Key[115]), .B(Plaintext[115]), .ZN(n7393) );
  OAI211_X1 U14428 ( .C1(n7613), .C2(n7393), .A(n8310), .B(n7934), .ZN(n6966)
         );
  AND2_X1 U14429 ( .A1(n6967), .A2(n6966), .ZN(n9230) );
  INV_X1 U14430 ( .A(n9230), .ZN(n9047) );
  INV_X1 U14431 ( .A(Plaintext[103]), .ZN(n6968) );
  INV_X1 U14432 ( .A(n7619), .ZN(n8235) );
  INV_X1 U14433 ( .A(Plaintext[104]), .ZN(n6969) );
  INV_X1 U14434 ( .A(Plaintext[107]), .ZN(n6970) );
  INV_X1 U14435 ( .A(Plaintext[106]), .ZN(n6971) );
  NAND2_X1 U14437 ( .A1(n7358), .A2(n8237), .ZN(n7431) );
  INV_X1 U14438 ( .A(Plaintext[102]), .ZN(n6972) );
  NAND2_X1 U14439 ( .A1(n8232), .A2(n8231), .ZN(n6974) );
  XNOR2_X1 U14440 ( .A(Key[100]), .B(Plaintext[100]), .ZN(n7362) );
  INV_X1 U14441 ( .A(Plaintext[101]), .ZN(n6977) );
  AND2_X1 U14442 ( .A1(n8205), .A2(n7362), .ZN(n6983) );
  INV_X1 U14443 ( .A(Plaintext[97]), .ZN(n6978) );
  INV_X1 U14445 ( .A(n7634), .ZN(n8199) );
  INV_X1 U14446 ( .A(Plaintext[99]), .ZN(n6979) );
  INV_X1 U14447 ( .A(n7635), .ZN(n8201) );
  NAND2_X1 U14448 ( .A1(n8199), .A2(n8201), .ZN(n6982) );
  INV_X1 U14449 ( .A(Plaintext[96]), .ZN(n6980) );
  INV_X1 U14451 ( .A(n7363), .ZN(n8207) );
  MUX2_X1 U14452 ( .A(n7832), .B(n8207), .S(n28605), .Z(n6981) );
  INV_X1 U14454 ( .A(Plaintext[93]), .ZN(n6984) );
  XNOR2_X1 U14455 ( .A(n6984), .B(Key[93]), .ZN(n6988) );
  INV_X1 U14456 ( .A(Plaintext[94]), .ZN(n6985) );
  XNOR2_X1 U14457 ( .A(n6985), .B(Key[94]), .ZN(n7825) );
  INV_X1 U14458 ( .A(n7825), .ZN(n7695) );
  INV_X1 U14459 ( .A(Plaintext[90]), .ZN(n6986) );
  OAI21_X1 U14460 ( .B1(n7821), .B2(n7695), .A(n6987), .ZN(n6994) );
  INV_X1 U14461 ( .A(Plaintext[91]), .ZN(n6989) );
  INV_X1 U14463 ( .A(Plaintext[92]), .ZN(n6990) );
  XNOR2_X1 U14464 ( .A(n6990), .B(Key[92]), .ZN(n7371) );
  XNOR2_X1 U14465 ( .A(Key[95]), .B(Plaintext[95]), .ZN(n8221) );
  INV_X1 U14466 ( .A(n8221), .ZN(n8223) );
  NAND2_X1 U14467 ( .A1(n6991), .A2(n8223), .ZN(n6992) );
  INV_X1 U14468 ( .A(Plaintext[120]), .ZN(n6995) );
  INV_X1 U14470 ( .A(Plaintext[121]), .ZN(n6996) );
  INV_X1 U14471 ( .A(n8290), .ZN(n7910) );
  INV_X1 U14472 ( .A(Plaintext[122]), .ZN(n6997) );
  INV_X1 U14474 ( .A(n7909), .ZN(n7914) );
  XNOR2_X1 U14475 ( .A(Key[124]), .B(Plaintext[124]), .ZN(n8287) );
  INV_X1 U14476 ( .A(Plaintext[123]), .ZN(n6998) );
  XNOR2_X1 U14477 ( .A(n6998), .B(Key[123]), .ZN(n7911) );
  XNOR2_X1 U14478 ( .A(Key[73]), .B(Plaintext[73]), .ZN(n7498) );
  INV_X1 U14479 ( .A(n7498), .ZN(n7708) );
  XNOR2_X1 U14480 ( .A(Key[75]), .B(Plaintext[75]), .ZN(n7382) );
  AND2_X1 U14481 ( .A1(n7498), .A2(n7382), .ZN(n7855) );
  INV_X1 U14482 ( .A(n7855), .ZN(n7002) );
  XNOR2_X1 U14483 ( .A(Key[74]), .B(Plaintext[74]), .ZN(n7852) );
  NAND3_X1 U14484 ( .A1(n7856), .A2(n7002), .A3(n3594), .ZN(n7006) );
  XNOR2_X1 U14485 ( .A(Key[76]), .B(Plaintext[76]), .ZN(n7384) );
  INV_X1 U14486 ( .A(n7384), .ZN(n7494) );
  INV_X1 U14487 ( .A(n7852), .ZN(n7496) );
  INV_X1 U14488 ( .A(Plaintext[72]), .ZN(n7003) );
  NAND2_X1 U14489 ( .A1(n617), .A2(n7382), .ZN(n7707) );
  NAND2_X1 U14490 ( .A1(n7707), .A2(n371), .ZN(n7004) );
  XNOR2_X1 U14491 ( .A(Key[67]), .B(Plaintext[67]), .ZN(n7850) );
  INV_X1 U14492 ( .A(Plaintext[69]), .ZN(n7007) );
  INV_X1 U14493 ( .A(Plaintext[71]), .ZN(n7008) );
  INV_X1 U14494 ( .A(Plaintext[66]), .ZN(n7009) );
  INV_X1 U14495 ( .A(n7846), .ZN(n7843) );
  NAND2_X1 U14497 ( .A1(n7846), .A2(n8023), .ZN(n7520) );
  INV_X1 U14498 ( .A(n7011), .ZN(n7685) );
  INV_X1 U14500 ( .A(n7844), .ZN(n7517) );
  INV_X1 U14501 ( .A(n8023), .ZN(n7684) );
  INV_X1 U14505 ( .A(Plaintext[86]), .ZN(n7015) );
  XNOR2_X1 U14506 ( .A(n7015), .B(Key[86]), .ZN(n7838) );
  INV_X1 U14507 ( .A(n7838), .ZN(n7835) );
  XNOR2_X1 U14508 ( .A(Key[85]), .B(Plaintext[85]), .ZN(n7836) );
  INV_X1 U14509 ( .A(Plaintext[88]), .ZN(n7016) );
  INV_X1 U14512 ( .A(n7690), .ZN(n8244) );
  XNOR2_X1 U14513 ( .A(Key[79]), .B(Plaintext[79]), .ZN(n7377) );
  INV_X1 U14514 ( .A(n7377), .ZN(n8246) );
  XNOR2_X1 U14515 ( .A(Key[81]), .B(Plaintext[81]), .ZN(n7017) );
  NAND2_X1 U14516 ( .A1(n7017), .A2(n7690), .ZN(n7816) );
  INV_X1 U14517 ( .A(n7017), .ZN(n7691) );
  NAND2_X1 U14518 ( .A1(n7691), .A2(n7692), .ZN(n7018) );
  NAND3_X1 U14519 ( .A1(n7816), .A2(n7817), .A3(n7018), .ZN(n7021) );
  XNOR2_X1 U14520 ( .A(Key[82]), .B(Plaintext[82]), .ZN(n7376) );
  INV_X1 U14521 ( .A(n7376), .ZN(n8247) );
  NAND3_X1 U14523 ( .A1(n8247), .A2(n7690), .A3(n7692), .ZN(n7020) );
  OAI211_X1 U14524 ( .C1(n7501), .C2(n8246), .A(n7021), .B(n7020), .ZN(n8877)
         );
  INV_X1 U14525 ( .A(n8881), .ZN(n8709) );
  INV_X1 U14526 ( .A(Plaintext[56]), .ZN(n7022) );
  XNOR2_X1 U14527 ( .A(Key[58]), .B(Plaintext[58]), .ZN(n7508) );
  NAND2_X1 U14528 ( .A1(n7257), .A2(n7508), .ZN(n7258) );
  INV_X1 U14530 ( .A(n7508), .ZN(n7729) );
  OAI21_X1 U14532 ( .B1(n7729), .B2(n7507), .A(n7506), .ZN(n7023) );
  NAND2_X1 U14533 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  OAI21_X1 U14534 ( .B1(n7258), .B2(n29629), .A(n7025), .ZN(n8404) );
  INV_X1 U14535 ( .A(n8404), .ZN(n8875) );
  INV_X1 U14536 ( .A(Plaintext[62]), .ZN(n7026) );
  INV_X1 U14538 ( .A(n7265), .ZN(n8030) );
  INV_X1 U14539 ( .A(Plaintext[65]), .ZN(n7027) );
  NAND2_X1 U14540 ( .A1(n8030), .A2(n7268), .ZN(n7735) );
  INV_X1 U14541 ( .A(Plaintext[64]), .ZN(n7028) );
  INV_X1 U14543 ( .A(Plaintext[61]), .ZN(n7029) );
  INV_X1 U14545 ( .A(n8032), .ZN(n7267) );
  INV_X1 U14546 ( .A(Plaintext[63]), .ZN(n7030) );
  NAND3_X1 U14547 ( .A1(n7521), .A2(n7267), .A3(n7709), .ZN(n7031) );
  XNOR2_X1 U14548 ( .A(Key[60]), .B(Plaintext[60]), .ZN(n7737) );
  INV_X1 U14549 ( .A(n7737), .ZN(n8028) );
  NAND3_X1 U14550 ( .A1(n7268), .A2(n7267), .A3(n7709), .ZN(n7032) );
  OAI21_X1 U14551 ( .B1(n8875), .B2(n8699), .A(n8710), .ZN(n7033) );
  NOR2_X1 U14552 ( .A1(n7033), .A2(n8876), .ZN(n7034) );
  XNOR2_X1 U14553 ( .A(n9732), .B(n10297), .ZN(n10343) );
  INV_X1 U14554 ( .A(Plaintext[153]), .ZN(n7036) );
  XNOR2_X1 U14555 ( .A(n7036), .B(Key[153]), .ZN(n7040) );
  INV_X1 U14556 ( .A(Plaintext[150]), .ZN(n7037) );
  NAND2_X1 U14557 ( .A1(n7982), .A2(n7456), .ZN(n7194) );
  INV_X1 U14558 ( .A(Plaintext[154]), .ZN(n7038) );
  INV_X1 U14559 ( .A(Plaintext[155]), .ZN(n7039) );
  XNOR2_X1 U14560 ( .A(n7039), .B(Key[155]), .ZN(n7192) );
  NAND2_X1 U14561 ( .A1(n7641), .A2(n7985), .ZN(n7041) );
  INV_X1 U14562 ( .A(n7040), .ZN(n7643) );
  AOI21_X1 U14563 ( .B1(n7194), .B2(n7041), .A(n7643), .ZN(n7044) );
  INV_X1 U14564 ( .A(Plaintext[152]), .ZN(n7042) );
  XNOR2_X1 U14565 ( .A(n7042), .B(Key[152]), .ZN(n7191) );
  INV_X1 U14566 ( .A(Plaintext[151]), .ZN(n7043) );
  INV_X1 U14567 ( .A(Plaintext[157]), .ZN(n7045) );
  NAND2_X1 U14569 ( .A1(n7965), .A2(n7675), .ZN(n7188) );
  INV_X1 U14570 ( .A(Plaintext[161]), .ZN(n7047) );
  INV_X1 U14571 ( .A(Plaintext[160]), .ZN(n7048) );
  XNOR2_X1 U14572 ( .A(n7048), .B(Key[160]), .ZN(n7966) );
  INV_X1 U14573 ( .A(n7965), .ZN(n7968) );
  INV_X1 U14574 ( .A(n8809), .ZN(n8523) );
  XNOR2_X1 U14575 ( .A(Key[170]), .B(Plaintext[170]), .ZN(n7589) );
  INV_X1 U14576 ( .A(Plaintext[173]), .ZN(n7050) );
  XNOR2_X1 U14577 ( .A(n7050), .B(Key[173]), .ZN(n7233) );
  INV_X1 U14578 ( .A(Plaintext[172]), .ZN(n7051) );
  XNOR2_X1 U14579 ( .A(n7051), .B(Key[172]), .ZN(n7958) );
  INV_X1 U14580 ( .A(n7958), .ZN(n7872) );
  NAND2_X1 U14582 ( .A1(n7869), .A2(n441), .ZN(n7053) );
  INV_X1 U14583 ( .A(Plaintext[171]), .ZN(n7052) );
  INV_X1 U14584 ( .A(n7592), .ZN(n7873) );
  OAI211_X2 U14585 ( .C1(n7875), .C2(n7872), .A(n7055), .B(n7054), .ZN(n8810)
         );
  MUX2_X1 U14586 ( .A(n8808), .B(n8523), .S(n8810), .Z(n7081) );
  INV_X1 U14587 ( .A(Plaintext[165]), .ZN(n7056) );
  INV_X1 U14588 ( .A(n7241), .ZN(n7060) );
  INV_X1 U14589 ( .A(Plaintext[166]), .ZN(n7057) );
  INV_X1 U14591 ( .A(n7999), .ZN(n7649) );
  OAI21_X1 U14592 ( .B1(n7060), .B2(n7059), .A(n8002), .ZN(n7066) );
  INV_X1 U14593 ( .A(Plaintext[163]), .ZN(n7061) );
  NAND2_X1 U14595 ( .A1(n7995), .A2(n7993), .ZN(n7652) );
  INV_X1 U14596 ( .A(n7652), .ZN(n7064) );
  INV_X1 U14597 ( .A(Plaintext[162]), .ZN(n7062) );
  INV_X1 U14599 ( .A(n7992), .ZN(n7994) );
  NOR2_X1 U14600 ( .A1(n7993), .A2(n7994), .ZN(n7063) );
  OAI21_X1 U14601 ( .B1(n7064), .B2(n7063), .A(n29081), .ZN(n7065) );
  INV_X1 U14602 ( .A(Plaintext[176]), .ZN(n7067) );
  XNOR2_X1 U14603 ( .A(n7067), .B(Key[176]), .ZN(n7069) );
  NAND2_X1 U14604 ( .A1(n7582), .A2(n7071), .ZN(n7237) );
  INV_X1 U14605 ( .A(Plaintext[175]), .ZN(n7068) );
  INV_X1 U14606 ( .A(n7069), .ZN(n7583) );
  INV_X1 U14607 ( .A(Plaintext[177]), .ZN(n7070) );
  XNOR2_X1 U14608 ( .A(n7070), .B(Key[177]), .ZN(n7072) );
  INV_X1 U14610 ( .A(n7071), .ZN(n7884) );
  INV_X1 U14611 ( .A(Plaintext[179]), .ZN(n7073) );
  XNOR2_X1 U14612 ( .A(Key[178]), .B(Plaintext[178]), .ZN(n7082) );
  INV_X1 U14613 ( .A(n7082), .ZN(n7581) );
  NAND3_X1 U14614 ( .A1(n7581), .A2(n7585), .A3(n7583), .ZN(n7075) );
  OAI211_X1 U14615 ( .C1(n7237), .C2(n7584), .A(n7076), .B(n7075), .ZN(n8811)
         );
  INV_X1 U14616 ( .A(n8811), .ZN(n8680) );
  OAI21_X1 U14617 ( .B1(n29241), .B2(n8810), .A(n8679), .ZN(n7080) );
  INV_X1 U14618 ( .A(n7172), .ZN(n7310) );
  XNOR2_X1 U14619 ( .A(Key[181]), .B(Plaintext[181]), .ZN(n7308) );
  INV_X1 U14620 ( .A(n7308), .ZN(n7862) );
  XNOR2_X1 U14621 ( .A(Key[180]), .B(Plaintext[180]), .ZN(n7865) );
  AOI21_X1 U14622 ( .B1(n7310), .B2(n7862), .A(n7865), .ZN(n7079) );
  INV_X1 U14623 ( .A(Plaintext[185]), .ZN(n7077) );
  XNOR2_X1 U14626 ( .A(Key[184]), .B(Plaintext[184]), .ZN(n7867) );
  NAND2_X1 U14627 ( .A1(n7095), .A2(n5149), .ZN(n7078) );
  OAI21_X1 U14628 ( .B1(n7883), .B2(n7585), .A(n7083), .ZN(n7084) );
  INV_X1 U14629 ( .A(Plaintext[4]), .ZN(n7085) );
  INV_X1 U14630 ( .A(Plaintext[3]), .ZN(n7086) );
  INV_X1 U14631 ( .A(n7315), .ZN(n7774) );
  INV_X1 U14632 ( .A(Plaintext[5]), .ZN(n7087) );
  NAND2_X1 U14634 ( .A1(n7090), .A2(n1350), .ZN(n7091) );
  INV_X1 U14635 ( .A(n7092), .ZN(n7601) );
  INV_X1 U14636 ( .A(n7093), .ZN(n7864) );
  NAND2_X1 U14637 ( .A1(n7864), .A2(n7867), .ZN(n7094) );
  NAND2_X1 U14638 ( .A1(n8586), .A2(n8192), .ZN(n7102) );
  XNOR2_X1 U14639 ( .A(Key[12]), .B(Plaintext[12]), .ZN(n7100) );
  INV_X1 U14640 ( .A(n7100), .ZN(n7289) );
  INV_X1 U14641 ( .A(Plaintext[13]), .ZN(n7096) );
  XNOR2_X1 U14642 ( .A(n7096), .B(Key[13]), .ZN(n8173) );
  INV_X1 U14643 ( .A(Plaintext[14]), .ZN(n7097) );
  XNOR2_X1 U14644 ( .A(n7097), .B(Key[14]), .ZN(n7101) );
  INV_X1 U14645 ( .A(n7101), .ZN(n7758) );
  INV_X1 U14646 ( .A(Plaintext[17]), .ZN(n7098) );
  NAND2_X1 U14647 ( .A1(n7758), .A2(n7759), .ZN(n7763) );
  INV_X1 U14648 ( .A(Plaintext[16]), .ZN(n7099) );
  XNOR2_X1 U14649 ( .A(n7099), .B(Key[16]), .ZN(n8176) );
  NAND2_X1 U14650 ( .A1(n7102), .A2(n8824), .ZN(n7120) );
  INV_X1 U14651 ( .A(Plaintext[187]), .ZN(n7103) );
  INV_X1 U14653 ( .A(Plaintext[189]), .ZN(n7104) );
  XNOR2_X1 U14654 ( .A(n7104), .B(Key[189]), .ZN(n7106) );
  NAND2_X1 U14655 ( .A1(n7801), .A2(n7895), .ZN(n7597) );
  INV_X1 U14656 ( .A(Plaintext[186]), .ZN(n7105) );
  INV_X1 U14657 ( .A(n7106), .ZN(n7800) );
  NAND2_X1 U14658 ( .A1(n7312), .A2(n7800), .ZN(n7107) );
  XNOR2_X1 U14659 ( .A(Key[191]), .B(Plaintext[191]), .ZN(n7110) );
  AOI21_X1 U14660 ( .B1(n7597), .B2(n7107), .A(n7898), .ZN(n7113) );
  INV_X1 U14661 ( .A(Plaintext[188]), .ZN(n7108) );
  INV_X1 U14662 ( .A(Plaintext[190]), .ZN(n7109) );
  NAND2_X1 U14663 ( .A1(n7900), .A2(n7897), .ZN(n7313) );
  INV_X1 U14664 ( .A(n7900), .ZN(n7896) );
  INV_X1 U14665 ( .A(n7110), .ZN(n7176) );
  INV_X1 U14668 ( .A(n8826), .ZN(n8830) );
  INV_X1 U14669 ( .A(Plaintext[6]), .ZN(n7115) );
  XNOR2_X1 U14671 ( .A(Key[7]), .B(Plaintext[7]), .ZN(n7162) );
  INV_X1 U14672 ( .A(Plaintext[8]), .ZN(n7117) );
  OAI21_X1 U14674 ( .B1(n7164), .B2(n7342), .A(n7770), .ZN(n7118) );
  NAND2_X1 U14675 ( .A1(n7447), .A2(n8826), .ZN(n7119) );
  INV_X1 U14676 ( .A(n9799), .ZN(n7121) );
  XNOR2_X1 U14677 ( .A(n7121), .B(n10037), .ZN(n8953) );
  XNOR2_X1 U14678 ( .A(n8953), .B(n10343), .ZN(n7230) );
  XNOR2_X1 U14679 ( .A(Key[37]), .B(Plaintext[37]), .ZN(n7722) );
  INV_X1 U14680 ( .A(n7722), .ZN(n8139) );
  XNOR2_X1 U14681 ( .A(Key[36]), .B(Plaintext[36]), .ZN(n8138) );
  INV_X1 U14682 ( .A(n8138), .ZN(n8041) );
  XNOR2_X1 U14683 ( .A(Key[39]), .B(Plaintext[39]), .ZN(n7560) );
  INV_X1 U14685 ( .A(Plaintext[38]), .ZN(n7122) );
  INV_X1 U14686 ( .A(Plaintext[40]), .ZN(n7123) );
  NAND2_X1 U14688 ( .A1(n8141), .A2(n8143), .ZN(n7562) );
  INV_X1 U14690 ( .A(n8141), .ZN(n8142) );
  MUX2_X2 U14691 ( .A(n7125), .B(n7124), .S(n7336), .Z(n9245) );
  INV_X1 U14693 ( .A(n8048), .ZN(n8134) );
  XNOR2_X1 U14694 ( .A(Key[45]), .B(Plaintext[45]), .ZN(n8047) );
  INV_X1 U14695 ( .A(n8047), .ZN(n8135) );
  INV_X1 U14696 ( .A(Plaintext[42]), .ZN(n7126) );
  XNOR2_X1 U14697 ( .A(n7126), .B(Key[42]), .ZN(n7554) );
  INV_X1 U14698 ( .A(Plaintext[46]), .ZN(n7128) );
  NAND2_X1 U14700 ( .A1(n7127), .A2(n8131), .ZN(n7717) );
  NAND2_X1 U14701 ( .A1(n8134), .A2(n29119), .ZN(n7130) );
  AOI21_X1 U14702 ( .B1(n7717), .B2(n7130), .A(n8049), .ZN(n7131) );
  INV_X1 U14703 ( .A(n9041), .ZN(n9248) );
  NAND2_X1 U14704 ( .A1(n7257), .A2(n7514), .ZN(n7733) );
  OAI21_X1 U14705 ( .B1(n8039), .B2(n7257), .A(n7733), .ZN(n7135) );
  INV_X1 U14706 ( .A(n7514), .ZN(n7728) );
  AOI21_X1 U14707 ( .B1(n7133), .B2(n7132), .A(n7507), .ZN(n7134) );
  INV_X1 U14708 ( .A(Plaintext[51]), .ZN(n7136) );
  AND2_X1 U14709 ( .A1(n7744), .A2(n28161), .ZN(n7146) );
  INV_X1 U14710 ( .A(Plaintext[53]), .ZN(n7137) );
  INV_X1 U14711 ( .A(Plaintext[48]), .ZN(n7138) );
  OAI21_X1 U14712 ( .B1(n8014), .B2(n7744), .A(n8013), .ZN(n7145) );
  INV_X1 U14713 ( .A(Plaintext[52]), .ZN(n7139) );
  INV_X1 U14715 ( .A(n8014), .ZN(n7746) );
  INV_X1 U14716 ( .A(Plaintext[49]), .ZN(n7140) );
  INV_X1 U14717 ( .A(n7743), .ZN(n7745) );
  INV_X1 U14718 ( .A(n8013), .ZN(n7747) );
  NAND2_X1 U14719 ( .A1(n7745), .A2(n7747), .ZN(n7142) );
  INV_X1 U14720 ( .A(n7141), .ZN(n7523) );
  INV_X1 U14722 ( .A(n8693), .ZN(n9039) );
  NOR2_X1 U14723 ( .A1(n9410), .A2(n9039), .ZN(n7160) );
  XNOR2_X1 U14724 ( .A(Key[27]), .B(Plaintext[27]), .ZN(n7150) );
  INV_X1 U14725 ( .A(Plaintext[26]), .ZN(n7147) );
  XNOR2_X1 U14726 ( .A(n7147), .B(Key[26]), .ZN(n7283) );
  MUX2_X1 U14727 ( .A(n7541), .B(n8150), .S(n8151), .Z(n7152) );
  INV_X1 U14728 ( .A(Plaintext[29]), .ZN(n7148) );
  XNOR2_X1 U14729 ( .A(n7148), .B(Key[29]), .ZN(n7285) );
  INV_X1 U14730 ( .A(n7285), .ZN(n8148) );
  INV_X1 U14731 ( .A(Plaintext[24]), .ZN(n7149) );
  INV_X1 U14732 ( .A(n7150), .ZN(n8147) );
  INV_X1 U14733 ( .A(Plaintext[31]), .ZN(n7153) );
  INV_X1 U14735 ( .A(Plaintext[30]), .ZN(n7154) );
  NAND2_X1 U14736 ( .A1(n8165), .A2(n7348), .ZN(n7297) );
  INV_X1 U14737 ( .A(n8161), .ZN(n8159) );
  INV_X1 U14738 ( .A(Plaintext[34]), .ZN(n7155) );
  XNOR2_X1 U14739 ( .A(n7155), .B(Key[34]), .ZN(n8158) );
  INV_X1 U14740 ( .A(n8158), .ZN(n7750) );
  INV_X1 U14742 ( .A(Plaintext[33]), .ZN(n7156) );
  XNOR2_X1 U14743 ( .A(n7156), .B(Key[33]), .ZN(n7298) );
  INV_X1 U14744 ( .A(n8165), .ZN(n8167) );
  NAND3_X1 U14745 ( .A1(n7157), .A2(n8162), .A3(n8167), .ZN(n7158) );
  NAND2_X1 U14746 ( .A1(n8166), .A2(n7349), .ZN(n7296) );
  NAND2_X1 U14748 ( .A1(n9041), .A2(n9243), .ZN(n8110) );
  INV_X1 U14749 ( .A(n7890), .ZN(n7778) );
  INV_X1 U14750 ( .A(n7889), .ZN(n7777) );
  INV_X1 U14751 ( .A(n7162), .ZN(n7321) );
  INV_X1 U14752 ( .A(n7342), .ZN(n7163) );
  INV_X1 U14753 ( .A(Plaintext[20]), .ZN(n7166) );
  INV_X1 U14754 ( .A(n7291), .ZN(n7781) );
  NAND2_X1 U14755 ( .A1(n7781), .A2(n7330), .ZN(n7168) );
  XNOR2_X1 U14756 ( .A(Key[19]), .B(Plaintext[19]), .ZN(n7787) );
  XNOR2_X1 U14757 ( .A(Key[18]), .B(Plaintext[18]), .ZN(n7786) );
  XNOR2_X1 U14758 ( .A(Key[22]), .B(Plaintext[22]), .ZN(n7550) );
  INV_X1 U14759 ( .A(n7550), .ZN(n7785) );
  XNOR2_X1 U14760 ( .A(Key[21]), .B(Plaintext[21]), .ZN(n7292) );
  INV_X1 U14761 ( .A(n7292), .ZN(n7782) );
  INV_X1 U14762 ( .A(n7787), .ZN(n7331) );
  AOI21_X1 U14763 ( .B1(n7782), .B2(n7331), .A(n7786), .ZN(n7169) );
  OR2_X1 U14764 ( .A1(n7169), .A2(n7781), .ZN(n7170) );
  NAND2_X2 U14765 ( .A1(n7171), .A2(n7170), .ZN(n8381) );
  INV_X1 U14766 ( .A(n8381), .ZN(n8536) );
  NAND2_X1 U14767 ( .A1(n7862), .A2(n7172), .ZN(n7173) );
  INV_X1 U14768 ( .A(n7865), .ZN(n7174) );
  NAND2_X1 U14769 ( .A1(n7310), .A2(n7174), .ZN(n7604) );
  NAND2_X1 U14770 ( .A1(n7801), .A2(n7312), .ZN(n7595) );
  INV_X1 U14771 ( .A(n7595), .ZN(n7177) );
  OAI21_X1 U14772 ( .B1(n7177), .B2(n7176), .A(n7803), .ZN(n7179) );
  INV_X1 U14773 ( .A(n7801), .ZN(n7902) );
  OAI211_X1 U14774 ( .C1(n7897), .C2(n7176), .A(n7800), .B(n7902), .ZN(n7178)
         );
  AND2_X1 U14775 ( .A1(n7179), .A2(n7178), .ZN(n8729) );
  NAND3_X1 U14776 ( .A1(n8537), .A2(n8729), .A3(n8381), .ZN(n7185) );
  NAND2_X1 U14777 ( .A1(n7289), .A2(n8177), .ZN(n8175) );
  NAND3_X1 U14778 ( .A1(n8175), .A2(n8179), .A3(n7289), .ZN(n7183) );
  NAND3_X1 U14779 ( .A1(n8175), .A2(n8179), .A3(n613), .ZN(n7181) );
  NOR2_X1 U14780 ( .A1(n8381), .A2(n8733), .ZN(n8538) );
  NAND2_X1 U14781 ( .A1(n8538), .A2(n8739), .ZN(n7184) );
  XNOR2_X1 U14782 ( .A(n10346), .B(n9542), .ZN(n10169) );
  AOI21_X1 U14783 ( .B1(n7188), .B2(n7962), .A(n4696), .ZN(n7190) );
  NAND2_X1 U14784 ( .A1(n7965), .A2(n1938), .ZN(n7236) );
  AOI21_X1 U14785 ( .B1(n7236), .B2(n7675), .A(n29302), .ZN(n7189) );
  INV_X1 U14787 ( .A(n7191), .ZN(n7980) );
  INV_X1 U14789 ( .A(n7981), .ZN(n7243) );
  OAI211_X1 U14790 ( .C1(n7456), .C2(n7243), .A(n7194), .B(n7642), .ZN(n7195)
         );
  INV_X1 U14791 ( .A(n8685), .ZN(n8688) );
  XNOR2_X1 U14792 ( .A(Key[139]), .B(Plaintext[139]), .ZN(n7480) );
  INV_X1 U14793 ( .A(n7480), .ZN(n8284) );
  INV_X1 U14794 ( .A(Plaintext[141]), .ZN(n7196) );
  XNOR2_X1 U14795 ( .A(n7196), .B(Key[141]), .ZN(n7405) );
  INV_X1 U14796 ( .A(n7405), .ZN(n7975) );
  OAI21_X1 U14799 ( .B1(n8284), .B2(n7975), .A(n7477), .ZN(n7217) );
  INV_X1 U14800 ( .A(Plaintext[140]), .ZN(n7197) );
  XNOR2_X1 U14801 ( .A(n7197), .B(Key[140]), .ZN(n7198) );
  NAND2_X1 U14803 ( .A1(n8281), .A2(n7975), .ZN(n8279) );
  NAND2_X1 U14804 ( .A1(n7199), .A2(n8279), .ZN(n7214) );
  INV_X1 U14805 ( .A(Plaintext[143]), .ZN(n7200) );
  XNOR2_X1 U14806 ( .A(n7200), .B(Key[143]), .ZN(n7404) );
  INV_X1 U14807 ( .A(Plaintext[132]), .ZN(n7201) );
  XNOR2_X1 U14808 ( .A(n7201), .B(Key[132]), .ZN(n7942) );
  INV_X1 U14809 ( .A(Plaintext[133]), .ZN(n7202) );
  NAND2_X1 U14811 ( .A1(n7942), .A2(n7657), .ZN(n7941) );
  NAND2_X1 U14812 ( .A1(n7941), .A2(n29317), .ZN(n7209) );
  INV_X1 U14813 ( .A(Plaintext[134]), .ZN(n7203) );
  NAND2_X1 U14815 ( .A1(n8305), .A2(n8297), .ZN(n7208) );
  INV_X1 U14816 ( .A(Plaintext[135]), .ZN(n7204) );
  XNOR2_X1 U14817 ( .A(n7204), .B(Key[135]), .ZN(n7399) );
  INV_X1 U14818 ( .A(n7399), .ZN(n8301) );
  INV_X1 U14819 ( .A(n7657), .ZN(n8303) );
  INV_X1 U14820 ( .A(Plaintext[136]), .ZN(n7205) );
  INV_X1 U14821 ( .A(n7655), .ZN(n7939) );
  NAND2_X1 U14822 ( .A1(n7939), .A2(n29317), .ZN(n7206) );
  INV_X1 U14823 ( .A(n8525), .ZN(n9222) );
  XNOR2_X1 U14824 ( .A(Key[148]), .B(Plaintext[148]), .ZN(n8267) );
  XNOR2_X1 U14825 ( .A(Key[145]), .B(Plaintext[145]), .ZN(n7485) );
  INV_X1 U14826 ( .A(n7485), .ZN(n8271) );
  XNOR2_X1 U14827 ( .A(Key[149]), .B(Plaintext[149]), .ZN(n7488) );
  INV_X1 U14828 ( .A(Plaintext[144]), .ZN(n7212) );
  XNOR2_X1 U14829 ( .A(n7212), .B(Key[144]), .ZN(n7665) );
  INV_X1 U14830 ( .A(n7665), .ZN(n8268) );
  INV_X1 U14831 ( .A(n9221), .ZN(n8686) );
  NAND2_X1 U14832 ( .A1(n8098), .A2(n8687), .ZN(n7227) );
  INV_X1 U14833 ( .A(n7214), .ZN(n7215) );
  INV_X1 U14834 ( .A(Plaintext[130]), .ZN(n7218) );
  INV_X1 U14836 ( .A(Plaintext[128]), .ZN(n7219) );
  NAND2_X1 U14837 ( .A1(n29590), .A2(n8256), .ZN(n8259) );
  INV_X1 U14838 ( .A(Plaintext[129]), .ZN(n7220) );
  NAND2_X1 U14839 ( .A1(n6782), .A2(n28617), .ZN(n7221) );
  NAND2_X1 U14840 ( .A1(n8259), .A2(n7221), .ZN(n7224) );
  XNOR2_X2 U14841 ( .A(Key[131]), .B(Plaintext[131]), .ZN(n8258) );
  INV_X1 U14842 ( .A(n8258), .ZN(n7465) );
  INV_X1 U14844 ( .A(n8263), .ZN(n7463) );
  OAI21_X1 U14845 ( .B1(n6782), .B2(n7618), .A(n7463), .ZN(n7223) );
  XNOR2_X1 U14846 ( .A(Key[126]), .B(Plaintext[126]), .ZN(n7466) );
  NAND2_X1 U14847 ( .A1(n28618), .A2(n7946), .ZN(n7222) );
  OAI21_X1 U14849 ( .B1(n9220), .B2(n8686), .A(n8687), .ZN(n7225) );
  XNOR2_X1 U14850 ( .A(n9971), .B(n26214), .ZN(n7228) );
  XNOR2_X1 U14851 ( .A(n10169), .B(n7228), .ZN(n7229) );
  NOR2_X1 U14852 ( .A1(n7591), .A2(n7870), .ZN(n7232) );
  OAI21_X1 U14853 ( .B1(n7592), .B2(n7872), .A(n7960), .ZN(n7235) );
  INV_X1 U14854 ( .A(n7594), .ZN(n7234) );
  NAND2_X1 U14855 ( .A1(n7887), .A2(n7583), .ZN(n7305) );
  NAND2_X1 U14856 ( .A1(n7581), .A2(n7884), .ZN(n7238) );
  NAND2_X1 U14857 ( .A1(n7999), .A2(n7876), .ZN(n7877) );
  INV_X1 U14858 ( .A(n7877), .ZN(n7240) );
  INV_X1 U14859 ( .A(n7995), .ZN(n7879) );
  AOI21_X1 U14860 ( .B1(n7998), .B2(n7879), .A(n6615), .ZN(n7239) );
  OAI21_X1 U14861 ( .B1(n7240), .B2(n7998), .A(n7239), .ZN(n7242) );
  NAND2_X1 U14863 ( .A1(n7644), .A2(n7457), .ZN(n7244) );
  NAND2_X1 U14865 ( .A1(n7485), .A2(n8269), .ZN(n7990) );
  INV_X1 U14866 ( .A(n7488), .ZN(n7986) );
  NOR2_X1 U14867 ( .A1(n29639), .A2(n8264), .ZN(n7245) );
  NAND2_X1 U14868 ( .A1(n8270), .A2(n8267), .ZN(n8266) );
  OAI21_X1 U14869 ( .B1(n7662), .B2(n7245), .A(n8266), .ZN(n7246) );
  NAND2_X1 U14871 ( .A1(n8134), .A2(n8047), .ZN(n7248) );
  OAI21_X1 U14872 ( .B1(n8049), .B2(n615), .A(n8133), .ZN(n7249) );
  NAND2_X1 U14873 ( .A1(n7251), .A2(n3594), .ZN(n7253) );
  NAND2_X1 U14874 ( .A1(n7251), .A2(n3639), .ZN(n7252) );
  NAND3_X1 U14875 ( .A1(n7253), .A2(n7252), .A3(n7708), .ZN(n7256) );
  INV_X1 U14876 ( .A(n7851), .ZN(n7853) );
  NAND2_X1 U14877 ( .A1(n7256), .A2(n7255), .ZN(n8763) );
  INV_X1 U14878 ( .A(n7257), .ZN(n8038) );
  INV_X1 U14879 ( .A(n29629), .ZN(n7511) );
  NAND2_X1 U14880 ( .A1(n8763), .A2(n9562), .ZN(n9565) );
  NAND2_X1 U14883 ( .A1(n7260), .A2(n29106), .ZN(n7264) );
  INV_X1 U14884 ( .A(n8024), .ZN(n7515) );
  NAND3_X1 U14885 ( .A1(n7847), .A2(n7684), .A3(n7261), .ZN(n7263) );
  NAND3_X1 U14886 ( .A1(n7517), .A2(n7685), .A3(n29130), .ZN(n7262) );
  INV_X1 U14888 ( .A(n8944), .ZN(n10401) );
  NAND3_X1 U14889 ( .A1(n7268), .A2(n8032), .A3(n8030), .ZN(n7272) );
  NAND3_X1 U14890 ( .A1(n7268), .A2(n7265), .A3(n7521), .ZN(n7271) );
  NAND3_X1 U14891 ( .A1(n7266), .A2(n7267), .A3(n8030), .ZN(n7270) );
  NAND3_X1 U14892 ( .A1(n618), .A2(n7709), .A3(n7737), .ZN(n7269) );
  AOI21_X2 U14893 ( .B1(n8947), .B2(n10401), .A(n7274), .ZN(n10191) );
  INV_X1 U14894 ( .A(n7891), .ZN(n7773) );
  MUX2_X1 U14895 ( .A(n7275), .B(n7889), .S(n7315), .Z(n7276) );
  NAND2_X1 U14896 ( .A1(n7770), .A2(n7342), .ZN(n7278) );
  NAND2_X1 U14897 ( .A1(n7279), .A2(n7278), .ZN(n7280) );
  NAND2_X1 U14898 ( .A1(n8334), .A2(n8889), .ZN(n8079) );
  NAND2_X1 U14899 ( .A1(n8147), .A2(n7793), .ZN(n7282) );
  INV_X1 U14900 ( .A(n8151), .ZN(n7284) );
  AOI21_X1 U14901 ( .B1(n7284), .B2(n8148), .A(n7542), .ZN(n7287) );
  NAND2_X1 U14903 ( .A1(n8177), .A2(n7758), .ZN(n7288) );
  INV_X1 U14904 ( .A(n8177), .ZN(n7760) );
  NAND2_X1 U14905 ( .A1(n7330), .A2(n7291), .ZN(n8154) );
  NAND2_X1 U14906 ( .A1(n1899), .A2(n7787), .ZN(n8156) );
  INV_X1 U14908 ( .A(n7330), .ZN(n8153) );
  NAND3_X1 U14909 ( .A1(n1899), .A2(n8153), .A3(n7786), .ZN(n7294) );
  AOI21_X1 U14910 ( .B1(n7297), .B2(n7296), .A(n7750), .ZN(n7300) );
  NAND2_X1 U14911 ( .A1(n8165), .A2(n7298), .ZN(n7535) );
  AOI21_X1 U14912 ( .B1(n7535), .B2(n7348), .A(n7349), .ZN(n7299) );
  OR2_X2 U14913 ( .A1(n7300), .A2(n7299), .ZN(n8009) );
  NAND3_X1 U14914 ( .A1(n8891), .A2(n8009), .A3(n8335), .ZN(n7301) );
  OAI211_X1 U14915 ( .C1(n8079), .C2(n8887), .A(n7302), .B(n7301), .ZN(n9795)
         );
  INV_X1 U14916 ( .A(n9795), .ZN(n9266) );
  NAND2_X1 U14917 ( .A1(n7172), .A2(n7865), .ZN(n7306) );
  NAND3_X1 U14918 ( .A1(n7310), .A2(n7309), .A3(n7308), .ZN(n7311) );
  NAND2_X1 U14920 ( .A1(n7315), .A2(n7777), .ZN(n7317) );
  NAND2_X1 U14921 ( .A1(n29112), .A2(n7089), .ZN(n7316) );
  OAI21_X1 U14922 ( .B1(n7594), .B2(n7872), .A(n7318), .ZN(n7319) );
  AOI22_X1 U14923 ( .A1(n9425), .A2(n7569), .B1(n8574), .B2(n8327), .ZN(n7328)
         );
  AOI21_X1 U14924 ( .B1(n7323), .B2(n7322), .A(n7342), .ZN(n7324) );
  NAND2_X1 U14925 ( .A1(n8327), .A2(n9425), .ZN(n7326) );
  NAND2_X1 U14926 ( .A1(n8580), .A2(n7326), .ZN(n7327) );
  XNOR2_X1 U14927 ( .A(n9266), .B(n10007), .ZN(n9003) );
  OAI211_X1 U14928 ( .C1(n7781), .C2(n7550), .A(n7332), .B(n8153), .ZN(n7334)
         );
  OAI21_X1 U14929 ( .B1(n7782), .B2(n7786), .A(n7330), .ZN(n7333) );
  NAND2_X1 U14930 ( .A1(n8041), .A2(n8139), .ZN(n7725) );
  INV_X1 U14931 ( .A(n7336), .ZN(n8043) );
  INV_X1 U14932 ( .A(n8143), .ZN(n7721) );
  NAND2_X1 U14933 ( .A1(n29751), .A2(n8139), .ZN(n7337) );
  AOI21_X1 U14934 ( .B1(n7337), .B2(n8041), .A(n8142), .ZN(n7338) );
  NAND2_X1 U14936 ( .A1(n614), .A2(n7342), .ZN(n7341) );
  NAND2_X1 U14937 ( .A1(n7341), .A2(n7767), .ZN(n7344) );
  NOR2_X1 U14938 ( .A1(n5242), .A2(n7342), .ZN(n7343) );
  NAND3_X1 U14939 ( .A1(n7345), .A2(n613), .A3(n7760), .ZN(n7346) );
  NAND2_X1 U14940 ( .A1(n8563), .A2(n8185), .ZN(n8939) );
  INV_X1 U14941 ( .A(n7348), .ZN(n8160) );
  OAI21_X1 U14942 ( .B1(n8162), .B2(n8160), .A(n8159), .ZN(n7351) );
  OAI21_X1 U14943 ( .B1(n8168), .B2(n7750), .A(n8161), .ZN(n7350) );
  NAND2_X1 U14944 ( .A1(n8167), .A2(n8160), .ZN(n7352) );
  AOI21_X1 U14945 ( .B1(n8937), .B2(n8939), .A(n9140), .ZN(n7356) );
  OAI21_X1 U14946 ( .B1(n8148), .B2(n28149), .A(n7542), .ZN(n7353) );
  NAND2_X1 U14947 ( .A1(n9139), .A2(n8185), .ZN(n8330) );
  AOI21_X1 U14948 ( .B1(n8330), .B2(n8563), .A(n8562), .ZN(n7355) );
  MUX2_X1 U14949 ( .A(n7357), .B(n8232), .S(n29110), .Z(n7361) );
  INV_X1 U14950 ( .A(n8237), .ZN(n7919) );
  INV_X1 U14951 ( .A(n8232), .ZN(n8236) );
  INV_X1 U14952 ( .A(n7358), .ZN(n7920) );
  NAND2_X1 U14955 ( .A1(n7635), .A2(n7828), .ZN(n7366) );
  INV_X1 U14956 ( .A(n7828), .ZN(n8202) );
  NAND3_X1 U14957 ( .A1(n3431), .A2(n8205), .A3(n7363), .ZN(n7364) );
  OAI211_X1 U14958 ( .C1(n7366), .C2(n8205), .A(n7365), .B(n7364), .ZN(n9149)
         );
  INV_X1 U14959 ( .A(n7837), .ZN(n8208) );
  NAND2_X1 U14960 ( .A1(n7371), .A2(n7825), .ZN(n8225) );
  INV_X1 U14961 ( .A(n7371), .ZN(n7824) );
  NAND2_X1 U14962 ( .A1(n7822), .A2(n7824), .ZN(n7372) );
  AOI21_X1 U14963 ( .B1(n8225), .B2(n7372), .A(n8221), .ZN(n7375) );
  NAND3_X1 U14964 ( .A1(n7821), .A2(n7824), .A3(n3821), .ZN(n7373) );
  NAND2_X1 U14965 ( .A1(n7376), .A2(n7692), .ZN(n7378) );
  NAND3_X1 U14966 ( .A1(n7378), .A2(n8245), .A3(n7818), .ZN(n7381) );
  NAND2_X1 U14967 ( .A1(n8243), .A2(n7690), .ZN(n7380) );
  NAND3_X1 U14968 ( .A1(n8246), .A2(n7817), .A3(n7692), .ZN(n7379) );
  INV_X1 U14969 ( .A(n7382), .ZN(n7705) );
  NAND3_X1 U14970 ( .A1(n9374), .A2(n9149), .A3(n5958), .ZN(n7386) );
  XNOR2_X1 U14971 ( .A(n10364), .B(n10193), .ZN(n9094) );
  NAND2_X1 U14972 ( .A1(n8263), .A2(n7618), .ZN(n8260) );
  NAND3_X1 U14973 ( .A1(n7463), .A2(n8258), .A3(n7946), .ZN(n7388) );
  NAND2_X1 U14974 ( .A1(n6782), .A2(n28615), .ZN(n7390) );
  AOI21_X1 U14975 ( .B1(n7390), .B2(n7389), .A(n8258), .ZN(n7391) );
  INV_X1 U14977 ( .A(n7393), .ZN(n8311) );
  NAND2_X1 U14978 ( .A1(n7613), .A2(n8311), .ZN(n7427) );
  AND2_X1 U14979 ( .A1(n7393), .A2(n7614), .ZN(n7610) );
  NAND2_X1 U14980 ( .A1(n7933), .A2(n29135), .ZN(n7394) );
  NAND2_X1 U14981 ( .A1(n7610), .A2(n7394), .ZN(n7395) );
  OAI211_X2 U14982 ( .C1(n28810), .C2(n7427), .A(n7395), .B(n7609), .ZN(n9340)
         );
  NAND2_X1 U14983 ( .A1(n9132), .A2(n9340), .ZN(n8340) );
  INV_X1 U14984 ( .A(n8340), .ZN(n7397) );
  INV_X1 U14985 ( .A(n7911), .ZN(n7916) );
  AOI21_X1 U14986 ( .B1(n7628), .B2(n7916), .A(n8290), .ZN(n7396) );
  NAND2_X1 U14987 ( .A1(n7924), .A2(n7626), .ZN(n7926) );
  NAND2_X1 U14988 ( .A1(n8216), .A2(n8213), .ZN(n7398) );
  INV_X1 U14989 ( .A(n8213), .ZN(n7438) );
  INV_X1 U14990 ( .A(n7942), .ZN(n8302) );
  INV_X1 U14991 ( .A(n7400), .ZN(n8296) );
  NAND3_X1 U14992 ( .A1(n7655), .A2(n8296), .A3(n29317), .ZN(n7401) );
  NAND2_X1 U14993 ( .A1(n7403), .A2(n9134), .ZN(n7413) );
  NAND2_X1 U14994 ( .A1(n8342), .A2(n9134), .ZN(n8549) );
  NAND2_X1 U14995 ( .A1(n7976), .A2(n8281), .ZN(n7671) );
  NAND2_X1 U14996 ( .A1(n7406), .A2(n8275), .ZN(n8285) );
  OAI21_X1 U14997 ( .B1(n7671), .B2(n8280), .A(n8285), .ZN(n7409) );
  NAND2_X1 U14998 ( .A1(n7406), .A2(n8276), .ZN(n7408) );
  INV_X1 U14999 ( .A(n9133), .ZN(n7410) );
  INV_X1 U15000 ( .A(n29247), .ZN(n27952) );
  NOR2_X1 U15001 ( .A1(n8608), .A2(n9533), .ZN(n7416) );
  NAND3_X1 U15002 ( .A1(n29662), .A2(n8749), .A3(n9533), .ZN(n7417) );
  OAI21_X1 U15003 ( .B1(n370), .B2(n8208), .A(n7839), .ZN(n7421) );
  NAND3_X1 U15004 ( .A1(n619), .A2(n7840), .A3(n8208), .ZN(n7422) );
  INV_X1 U15005 ( .A(n8741), .ZN(n9074) );
  AND2_X1 U15006 ( .A1(n7827), .A2(n7695), .ZN(n7425) );
  INV_X1 U15007 ( .A(n8740), .ZN(n8378) );
  AOI21_X1 U15008 ( .B1(n7427), .B2(n7609), .A(n7933), .ZN(n7429) );
  AOI21_X1 U15009 ( .B1(n7930), .B2(n7613), .A(n7935), .ZN(n7428) );
  NOR2_X1 U15012 ( .A1(n9073), .A2(n8740), .ZN(n8855) );
  NAND2_X1 U15013 ( .A1(n7634), .A2(n7635), .ZN(n7829) );
  NAND2_X1 U15014 ( .A1(n7635), .A2(n7363), .ZN(n7433) );
  AOI21_X1 U15015 ( .B1(n8200), .B2(n7433), .A(n7830), .ZN(n7434) );
  INV_X1 U15016 ( .A(n9070), .ZN(n8856) );
  OAI21_X1 U15017 ( .B1(n8855), .B2(n8856), .A(n9075), .ZN(n7443) );
  NAND2_X1 U15018 ( .A1(n8217), .A2(n627), .ZN(n7441) );
  NAND3_X1 U15019 ( .A1(n7441), .A2(n7437), .A3(n7436), .ZN(n7440) );
  NAND3_X1 U15020 ( .A1(n7438), .A2(n8216), .A3(n7925), .ZN(n7439) );
  OAI211_X1 U15021 ( .C1(n7441), .C2(n7925), .A(n7440), .B(n7439), .ZN(n8857)
         );
  NAND2_X1 U15022 ( .A1(n8855), .A2(n8857), .ZN(n7442) );
  XNOR2_X1 U15023 ( .A(n9996), .B(n9754), .ZN(n7449) );
  NAND2_X1 U15024 ( .A1(n8824), .A2(n8826), .ZN(n7444) );
  OAI21_X1 U15025 ( .B1(n7445), .B2(n8824), .A(n7444), .ZN(n7446) );
  OAI21_X1 U15026 ( .B1(n7447), .B2(n8196), .A(n7446), .ZN(n9447) );
  XNOR2_X1 U15027 ( .A(n9447), .B(n3212), .ZN(n7448) );
  XNOR2_X1 U15028 ( .A(n7449), .B(n7448), .ZN(n7573) );
  NAND2_X1 U15029 ( .A1(n7399), .A2(n7657), .ZN(n7943) );
  NAND2_X1 U15030 ( .A1(n8305), .A2(n7655), .ZN(n7452) );
  NAND2_X1 U15031 ( .A1(n8296), .A2(n8304), .ZN(n7451) );
  NAND2_X1 U15034 ( .A1(n7456), .A2(n7981), .ZN(n7458) );
  AOI21_X1 U15035 ( .B1(n7459), .B2(n7458), .A(n7457), .ZN(n7460) );
  NAND2_X1 U15036 ( .A1(n29590), .A2(n8258), .ZN(n7464) );
  INV_X1 U15038 ( .A(n28614), .ZN(n7948) );
  INV_X1 U15039 ( .A(n7466), .ZN(n8257) );
  INV_X1 U15040 ( .A(n7618), .ZN(n7947) );
  INV_X1 U15042 ( .A(n8287), .ZN(n7631) );
  INV_X1 U15043 ( .A(n7912), .ZN(n7470) );
  OAI21_X1 U15044 ( .B1(n7631), .B2(n7470), .A(n7916), .ZN(n7472) );
  INV_X1 U15045 ( .A(n7628), .ZN(n7917) );
  NAND2_X1 U15046 ( .A1(n29568), .A2(n7917), .ZN(n7471) );
  AND2_X1 U15047 ( .A1(n7472), .A2(n7471), .ZN(n7476) );
  AOI21_X1 U15048 ( .B1(n7474), .B2(n7473), .A(n7915), .ZN(n7475) );
  OAI21_X1 U15050 ( .B1(n8280), .B2(n8281), .A(n7976), .ZN(n7478) );
  AND2_X1 U15052 ( .A1(n7480), .A2(n7975), .ZN(n7670) );
  INV_X1 U15053 ( .A(n7670), .ZN(n7481) );
  INV_X1 U15054 ( .A(n9080), .ZN(n7484) );
  NAND3_X1 U15055 ( .A1(n7484), .A2(n8605), .A3(n8603), .ZN(n7492) );
  OR2_X1 U15056 ( .A1(n9080), .A2(n8726), .ZN(n8851) );
  OAI21_X1 U15057 ( .B1(n341), .B2(n8268), .A(n7486), .ZN(n7487) );
  INV_X1 U15058 ( .A(n8270), .ZN(n7663) );
  NAND2_X1 U15059 ( .A1(n7487), .A2(n7663), .ZN(n9082) );
  INV_X1 U15061 ( .A(n9313), .ZN(n7530) );
  NAND2_X1 U15062 ( .A1(n7494), .A2(n7852), .ZN(n7495) );
  MUX2_X1 U15063 ( .A(n7497), .B(n7495), .S(n7851), .Z(n7500) );
  OAI21_X1 U15064 ( .B1(n8242), .B2(n8244), .A(n7501), .ZN(n7505) );
  NAND2_X1 U15065 ( .A1(n8247), .A2(n7817), .ZN(n7503) );
  AOI21_X1 U15067 ( .B1(n7503), .B2(n7502), .A(n7818), .ZN(n7504) );
  INV_X1 U15068 ( .A(n7507), .ZN(n7732) );
  NAND2_X1 U15069 ( .A1(n7732), .A2(n8034), .ZN(n8036) );
  NAND2_X1 U15070 ( .A1(n7507), .A2(n7506), .ZN(n8035) );
  NAND2_X1 U15071 ( .A1(n8034), .A2(n7508), .ZN(n7509) );
  NAND2_X1 U15072 ( .A1(n7510), .A2(n7509), .ZN(n7513) );
  NAND2_X1 U15075 ( .A1(n7850), .A2(n29130), .ZN(n7516) );
  OAI211_X1 U15076 ( .C1(n7517), .C2(n29130), .A(n7516), .B(n29106), .ZN(n7518) );
  NOR2_X1 U15077 ( .A1(n8817), .A2(n8592), .ZN(n8129) );
  INV_X1 U15078 ( .A(n8129), .ZN(n7529) );
  INV_X1 U15079 ( .A(n7521), .ZN(n7734) );
  NAND2_X1 U15081 ( .A1(n7266), .A2(n8032), .ZN(n7738) );
  OAI21_X1 U15082 ( .B1(n7266), .B2(n7737), .A(n7738), .ZN(n7522) );
  NAND2_X1 U15083 ( .A1(n7523), .A2(n8014), .ZN(n7748) );
  AOI21_X1 U15086 ( .B1(n7525), .B2(n7747), .A(n7744), .ZN(n7526) );
  NAND2_X1 U15087 ( .A1(n2024), .A2(n607), .ZN(n7528) );
  XNOR2_X1 U15088 ( .A(n7530), .B(n10395), .ZN(n10288) );
  INV_X1 U15089 ( .A(n10288), .ZN(n7571) );
  NAND2_X1 U15090 ( .A1(n7743), .A2(n7742), .ZN(n8015) );
  NAND2_X1 U15091 ( .A1(n8015), .A2(n8013), .ZN(n7532) );
  INV_X1 U15092 ( .A(n7533), .ZN(n7749) );
  INV_X1 U15093 ( .A(n9062), .ZN(n8393) );
  NAND3_X1 U15094 ( .A1(n7536), .A2(n8159), .A3(n7535), .ZN(n7539) );
  NAND2_X1 U15095 ( .A1(n7537), .A2(n8161), .ZN(n7538) );
  NAND2_X1 U15096 ( .A1(n8393), .A2(n9060), .ZN(n8871) );
  AND2_X1 U15097 ( .A1(n28149), .A2(n8148), .ZN(n7546) );
  INV_X1 U15098 ( .A(n7792), .ZN(n7540) );
  NAND2_X1 U15099 ( .A1(n7541), .A2(n7540), .ZN(n7545) );
  OAI21_X1 U15102 ( .B1(n7546), .B2(n7545), .A(n7544), .ZN(n8865) );
  OAI21_X1 U15103 ( .B1(n7785), .B2(n7787), .A(n1899), .ZN(n7548) );
  NAND2_X1 U15104 ( .A1(n7782), .A2(n7786), .ZN(n7547) );
  NAND2_X1 U15105 ( .A1(n7548), .A2(n7547), .ZN(n7553) );
  NAND2_X1 U15106 ( .A1(n7291), .A2(n7550), .ZN(n7549) );
  OAI21_X1 U15107 ( .B1(n7550), .B2(n1899), .A(n7549), .ZN(n7551) );
  NAND2_X1 U15108 ( .A1(n7551), .A2(n7330), .ZN(n7552) );
  NAND2_X1 U15109 ( .A1(n7553), .A2(n7552), .ZN(n8397) );
  NAND2_X1 U15110 ( .A1(n8865), .A2(n8397), .ZN(n8104) );
  NAND2_X1 U15111 ( .A1(n9062), .A2(n8104), .ZN(n7568) );
  MUX2_X1 U15112 ( .A(n29646), .B(n7127), .S(n8047), .Z(n7555) );
  NAND2_X1 U15113 ( .A1(n7555), .A2(n7554), .ZN(n7559) );
  NAND2_X1 U15115 ( .A1(n8044), .A2(n8138), .ZN(n7561) );
  NAND2_X1 U15116 ( .A1(n7561), .A2(n7336), .ZN(n7564) );
  NAND2_X1 U15117 ( .A1(n8043), .A2(n7562), .ZN(n7563) );
  NAND2_X1 U15118 ( .A1(n7564), .A2(n7563), .ZN(n7567) );
  MUX2_X1 U15119 ( .A(n7723), .B(n7565), .S(n7722), .Z(n7566) );
  INV_X1 U15120 ( .A(n8865), .ZN(n9059) );
  NAND2_X1 U15121 ( .A1(n8581), .A2(n606), .ZN(n9581) );
  NOR2_X1 U15122 ( .A1(n7569), .A2(n9421), .ZN(n8770) );
  XNOR2_X1 U15123 ( .A(n9779), .B(n10201), .ZN(n7570) );
  INV_X1 U15124 ( .A(n11146), .ZN(n7813) );
  INV_X1 U15125 ( .A(n8729), .ZN(n8734) );
  AND2_X1 U15126 ( .A1(n8381), .A2(n8733), .ZN(n8369) );
  NAND2_X1 U15127 ( .A1(n6909), .A2(n8537), .ZN(n7574) );
  AOI21_X1 U15129 ( .B1(n4696), .B2(n29301), .A(n1568), .ZN(n7577) );
  NAND2_X1 U15130 ( .A1(n7966), .A2(n7964), .ZN(n7576) );
  NAND2_X1 U15133 ( .A1(n7995), .A2(n7992), .ZN(n7651) );
  NAND2_X1 U15134 ( .A1(n8002), .A2(n7649), .ZN(n7579) );
  NAND2_X1 U15135 ( .A1(n7582), .A2(n7581), .ZN(n7587) );
  NAND2_X1 U15136 ( .A1(n7584), .A2(n7583), .ZN(n7586) );
  AOI21_X1 U15137 ( .B1(n7587), .B2(n7586), .A(n7585), .ZN(n7588) );
  INV_X1 U15139 ( .A(n8718), .ZN(n8785) );
  INV_X1 U15140 ( .A(n7897), .ZN(n7805) );
  AOI21_X1 U15141 ( .B1(n7596), .B2(n7595), .A(n7805), .ZN(n7599) );
  AOI21_X1 U15142 ( .B1(n7597), .B2(n7312), .A(n7896), .ZN(n7598) );
  NAND2_X1 U15143 ( .A1(n7862), .A2(n7865), .ZN(n7600) );
  NAND3_X1 U15144 ( .A1(n7604), .A2(n7601), .A3(n7600), .ZN(n7603) );
  NOR2_X1 U15145 ( .A1(n8788), .A2(n8718), .ZN(n7605) );
  AOI22_X1 U15146 ( .A1(n7606), .A2(n8787), .B1(n7605), .B2(n8717), .ZN(n7608)
         );
  OAI211_X2 U15147 ( .C1(n8438), .C2(n8442), .A(n7608), .B(n7607), .ZN(n10019)
         );
  OAI21_X1 U15148 ( .B1(n8311), .B2(n7934), .A(n7609), .ZN(n7612) );
  INV_X1 U15149 ( .A(n7610), .ZN(n7611) );
  INV_X1 U15151 ( .A(n7613), .ZN(n7931) );
  NAND2_X1 U15152 ( .A1(n7931), .A2(n7614), .ZN(n7615) );
  INV_X1 U15153 ( .A(n9196), .ZN(n8779) );
  INV_X1 U15154 ( .A(n329), .ZN(n9201) );
  NAND2_X1 U15155 ( .A1(n2089), .A2(n7920), .ZN(n7621) );
  NAND3_X1 U15156 ( .A1(n7621), .A2(n8231), .A3(n8235), .ZN(n7622) );
  NAND2_X1 U15158 ( .A1(n7925), .A2(n8213), .ZN(n7927) );
  NAND2_X1 U15159 ( .A1(n8217), .A2(n7626), .ZN(n7624) );
  NAND3_X1 U15160 ( .A1(n7626), .A2(n8216), .A3(n7925), .ZN(n7627) );
  INV_X1 U15161 ( .A(n9200), .ZN(n9194) );
  NAND2_X1 U15162 ( .A1(n29568), .A2(n7628), .ZN(n7633) );
  NAND2_X1 U15163 ( .A1(n7631), .A2(n7915), .ZN(n7632) );
  MUX2_X1 U15164 ( .A(n7636), .B(n8202), .S(n7635), .Z(n7637) );
  INV_X1 U15165 ( .A(n9197), .ZN(n9195) );
  NAND3_X1 U15166 ( .A1(n9195), .A2(n8779), .A3(n9201), .ZN(n7638) );
  INV_X1 U15168 ( .A(n9211), .ZN(n9435) );
  AOI21_X1 U15170 ( .B1(n7652), .B2(n7992), .A(n7998), .ZN(n7653) );
  NAND2_X1 U15172 ( .A1(n8304), .A2(n7655), .ZN(n7656) );
  AOI21_X1 U15173 ( .B1(n8298), .B2(n7656), .A(n29317), .ZN(n7661) );
  NAND2_X1 U15177 ( .A1(n7664), .A2(n7663), .ZN(n7668) );
  NAND3_X1 U15178 ( .A1(n631), .A2(n8270), .A3(n8264), .ZN(n7667) );
  NAND3_X1 U15179 ( .A1(n8265), .A2(n7986), .A3(n341), .ZN(n7666) );
  INV_X1 U15180 ( .A(n8777), .ZN(n9436) );
  INV_X1 U15181 ( .A(n8996), .ZN(n9209) );
  INV_X1 U15182 ( .A(n29301), .ZN(n7674) );
  OAI21_X1 U15183 ( .B1(n7675), .B2(n7968), .A(n7674), .ZN(n7677) );
  NAND2_X1 U15184 ( .A1(n7966), .A2(n29302), .ZN(n7676) );
  NAND3_X1 U15185 ( .A1(n9434), .A2(n8777), .A3(n9210), .ZN(n7681) );
  XNOR2_X1 U15186 ( .A(n9772), .B(n10322), .ZN(n9675) );
  XNOR2_X1 U15187 ( .A(n8883), .B(n9675), .ZN(n7812) );
  NAND2_X1 U15188 ( .A1(n8022), .A2(n7685), .ZN(n7689) );
  NAND2_X1 U15189 ( .A1(n7684), .A2(n29106), .ZN(n7688) );
  AND2_X1 U15190 ( .A1(n7850), .A2(n7843), .ZN(n7687) );
  NAND2_X1 U15192 ( .A1(n7821), .A2(n7822), .ZN(n7697) );
  NAND2_X1 U15193 ( .A1(n439), .A2(n7367), .ZN(n7704) );
  NAND2_X1 U15194 ( .A1(n619), .A2(n7839), .ZN(n7701) );
  OAI211_X1 U15195 ( .C1(n7840), .C2(n7839), .A(n7701), .B(n7700), .ZN(n7703)
         );
  NAND3_X1 U15196 ( .A1(n7837), .A2(n7835), .A3(n370), .ZN(n7702) );
  NAND2_X1 U15197 ( .A1(n9034), .A2(n8792), .ZN(n8360) );
  AOI21_X1 U15198 ( .B1(n7711), .B2(n7710), .A(n618), .ZN(n7712) );
  XNOR2_X1 U15199 ( .A(n10384), .B(n2511), .ZN(n7810) );
  AOI21_X1 U15200 ( .B1(n8135), .B2(n8048), .A(n8049), .ZN(n7719) );
  NAND2_X1 U15201 ( .A1(n9188), .A2(n9007), .ZN(n7741) );
  INV_X1 U15202 ( .A(n7726), .ZN(n8445) );
  NAND3_X1 U15203 ( .A1(n7729), .A2(n8038), .A3(n29629), .ZN(n7730) );
  NAND2_X1 U15205 ( .A1(n8445), .A2(n9186), .ZN(n7740) );
  NAND2_X1 U15206 ( .A1(n7265), .A2(n7737), .ZN(n8033) );
  OAI21_X1 U15207 ( .B1(n7738), .B2(n8030), .A(n8033), .ZN(n7739) );
  INV_X1 U15208 ( .A(n8782), .ZN(n9187) );
  AOI21_X1 U15209 ( .B1(n7741), .B2(n7740), .A(n9187), .ZN(n7757) );
  MUX2_X1 U15210 ( .A(n8160), .B(n8167), .S(n8162), .Z(n7754) );
  NAND2_X1 U15211 ( .A1(n7751), .A2(n8159), .ZN(n7753) );
  AND2_X1 U15212 ( .A1(n8162), .A2(n8158), .ZN(n7752) );
  AOI21_X2 U15213 ( .B1(n7754), .B2(n7753), .A(n7752), .ZN(n9009) );
  INV_X1 U15214 ( .A(n9007), .ZN(n9185) );
  NAND2_X1 U15215 ( .A1(n613), .A2(n7758), .ZN(n7762) );
  AND2_X1 U15217 ( .A1(n7775), .A2(n7089), .ZN(n7893) );
  INV_X1 U15218 ( .A(n7893), .ZN(n7780) );
  NAND3_X1 U15219 ( .A1(n7778), .A2(n7777), .A3(n438), .ZN(n7779) );
  INV_X1 U15221 ( .A(n7786), .ZN(n7783) );
  NAND2_X1 U15222 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  MUX2_X1 U15223 ( .A(n7789), .B(n7788), .S(n7291), .Z(n7790) );
  AOI21_X1 U15224 ( .B1(n7794), .B2(n7793), .A(n8150), .ZN(n7799) );
  NAND2_X1 U15225 ( .A1(n7796), .A2(n8150), .ZN(n7797) );
  OAI211_X1 U15226 ( .C1(n8353), .C2(n8351), .A(n7809), .B(n8077), .ZN(n7808)
         );
  XNOR2_X1 U15229 ( .A(n7810), .B(n10179), .ZN(n7811) );
  NAND2_X1 U15230 ( .A1(n8244), .A2(n7376), .ZN(n7815) );
  AND2_X1 U15231 ( .A1(n7815), .A2(n7816), .ZN(n7820) );
  NAND2_X1 U15232 ( .A1(n608), .A2(n9012), .ZN(n9019) );
  AOI21_X1 U15233 ( .B1(n7829), .B2(n7828), .A(n7363), .ZN(n7834) );
  AOI21_X1 U15234 ( .B1(n7832), .B2(n7831), .A(n7362), .ZN(n7833) );
  INV_X1 U15235 ( .A(n8910), .ZN(n9018) );
  NAND2_X1 U15236 ( .A1(n9019), .A2(n5674), .ZN(n7860) );
  AND2_X1 U15237 ( .A1(n7836), .A2(n7840), .ZN(n8209) );
  NAND2_X1 U15239 ( .A1(n7844), .A2(n8023), .ZN(n7845) );
  OAI211_X1 U15240 ( .C1(n7846), .C2(n7844), .A(n7845), .B(n29106), .ZN(n7848)
         );
  NAND2_X1 U15241 ( .A1(n8908), .A2(n9014), .ZN(n8906) );
  NAND2_X1 U15242 ( .A1(n8906), .A2(n8910), .ZN(n7859) );
  NAND2_X1 U15243 ( .A1(n7851), .A2(n7384), .ZN(n7854) );
  AOI22_X1 U15244 ( .A1(n7855), .A2(n7854), .B1(n7853), .B2(n7852), .ZN(n7858)
         );
  INV_X1 U15245 ( .A(n9015), .ZN(n9013) );
  NAND3_X1 U15246 ( .A1(n7865), .A2(n7172), .A3(n7864), .ZN(n7866) );
  NAND2_X1 U15247 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  INV_X1 U15248 ( .A(n8116), .ZN(n8655) );
  NAND2_X1 U15249 ( .A1(n29082), .A2(n7997), .ZN(n7881) );
  NAND3_X1 U15250 ( .A1(n7877), .A2(n7993), .A3(n7994), .ZN(n7880) );
  INV_X1 U15251 ( .A(n7993), .ZN(n7878) );
  INV_X1 U15252 ( .A(n8502), .ZN(n8651) );
  NOR2_X1 U15253 ( .A1(n7890), .A2(n7889), .ZN(n7892) );
  OAI21_X1 U15254 ( .B1(n7893), .B2(n7892), .A(n29112), .ZN(n7894) );
  NOR2_X1 U15255 ( .A1(n8658), .A2(n8502), .ZN(n7905) );
  NAND2_X1 U15256 ( .A1(n7895), .A2(n7312), .ZN(n7901) );
  MUX2_X1 U15257 ( .A(n7901), .B(n7899), .S(n7898), .Z(n7904) );
  OAI211_X1 U15258 ( .C1(n7312), .C2(n7902), .A(n7901), .B(n7900), .ZN(n7903)
         );
  AOI22_X1 U15259 ( .A1(n7906), .A2(n8658), .B1(n7905), .B2(n8653), .ZN(n7907)
         );
  NAND2_X1 U15260 ( .A1(n7910), .A2(n7909), .ZN(n8292) );
  INV_X1 U15261 ( .A(n9116), .ZN(n8917) );
  MUX2_X1 U15262 ( .A(n8231), .B(n7919), .S(n7920), .Z(n7923) );
  MUX2_X1 U15263 ( .A(n7921), .B(n8236), .S(n5946), .Z(n7922) );
  NAND2_X1 U15264 ( .A1(n8917), .A2(n9108), .ZN(n8671) );
  INV_X1 U15265 ( .A(n9108), .ZN(n9106) );
  NAND2_X1 U15266 ( .A1(n8212), .A2(n7925), .ZN(n7929) );
  INV_X1 U15267 ( .A(n7926), .ZN(n7928) );
  NAND2_X1 U15268 ( .A1(n9106), .A2(n8669), .ZN(n7938) );
  OAI21_X1 U15269 ( .B1(n7932), .B2(n7931), .A(n7930), .ZN(n9109) );
  INV_X1 U15270 ( .A(n7935), .ZN(n7934) );
  NAND2_X1 U15271 ( .A1(n7934), .A2(n7933), .ZN(n7937) );
  NAND2_X1 U15272 ( .A1(n7935), .A2(n7614), .ZN(n7936) );
  AND2_X1 U15273 ( .A1(n7937), .A2(n7936), .ZN(n9112) );
  MUX2_X2 U15274 ( .A(n9109), .B(n9112), .S(n29135), .Z(n8670) );
  AOI21_X1 U15275 ( .B1(n8671), .B2(n7938), .A(n8511), .ZN(n7956) );
  AOI21_X1 U15276 ( .B1(n7941), .B2(n7940), .A(n7939), .ZN(n7945) );
  AOI21_X1 U15277 ( .B1(n7943), .B2(n7942), .A(n8296), .ZN(n7944) );
  INV_X1 U15278 ( .A(n8914), .ZN(n8513) );
  NAND2_X1 U15279 ( .A1(n28618), .A2(n8257), .ZN(n7952) );
  NAND3_X1 U15280 ( .A1(n6782), .A2(n7948), .A3(n8258), .ZN(n7950) );
  NAND2_X1 U15281 ( .A1(n8513), .A2(n9107), .ZN(n7954) );
  NAND3_X1 U15282 ( .A1(n9108), .A2(n9116), .A3(n8914), .ZN(n7953) );
  INV_X1 U15284 ( .A(n8666), .ZN(n8492) );
  NAND2_X1 U15285 ( .A1(n7967), .A2(n7966), .ZN(n7971) );
  MUX2_X1 U15287 ( .A(n7971), .B(n7970), .S(n29302), .Z(n7972) );
  NAND2_X1 U15288 ( .A1(n8284), .A2(n8280), .ZN(n7974) );
  MUX2_X1 U15289 ( .A(n7974), .B(n8275), .S(n8276), .Z(n7979) );
  NOR2_X1 U15290 ( .A1(n7975), .A2(n8280), .ZN(n7977) );
  NAND2_X1 U15291 ( .A1(n8665), .A2(n8073), .ZN(n8006) );
  NAND2_X1 U15292 ( .A1(n7982), .A2(n7981), .ZN(n7983) );
  AND2_X1 U15293 ( .A1(n8267), .A2(n8264), .ZN(n7989) );
  NAND2_X1 U15294 ( .A1(n7986), .A2(n8270), .ZN(n7988) );
  NAND3_X1 U15295 ( .A1(n8271), .A2(n8265), .A3(n8264), .ZN(n7987) );
  NAND2_X1 U15296 ( .A1(n7993), .A2(n7992), .ZN(n8003) );
  NAND2_X1 U15297 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  NAND3_X1 U15298 ( .A1(n8003), .A2(n7997), .A3(n7996), .ZN(n8001) );
  NAND3_X1 U15299 ( .A1(n7999), .A2(n8002), .A3(n7998), .ZN(n8000) );
  OAI211_X1 U15300 ( .C1(n8003), .C2(n8002), .A(n8001), .B(n8000), .ZN(n9095)
         );
  OAI211_X1 U15301 ( .C1(n8492), .C2(n8006), .A(n8005), .B(n8004), .ZN(n10310)
         );
  XNOR2_X1 U15302 ( .A(n10310), .B(n10357), .ZN(n9672) );
  XNOR2_X1 U15303 ( .A(n10433), .B(n9672), .ZN(n8063) );
  OAI21_X1 U15304 ( .B1(n8334), .B2(n8889), .A(n8007), .ZN(n8008) );
  INV_X1 U15306 ( .A(n8009), .ZN(n8507) );
  NAND3_X1 U15307 ( .A1(n8507), .A2(n8891), .A3(n8335), .ZN(n8011) );
  NAND2_X1 U15308 ( .A1(n8009), .A2(n8336), .ZN(n8888) );
  NAND3_X1 U15310 ( .A1(n8016), .A2(n8015), .A3(n8014), .ZN(n8017) );
  NAND2_X1 U15311 ( .A1(n8019), .A2(n28161), .ZN(n8020) );
  NAND2_X1 U15312 ( .A1(n29106), .A2(n29130), .ZN(n8021) );
  AOI21_X1 U15313 ( .B1(n8022), .B2(n8021), .A(n7844), .ZN(n8026) );
  INV_X1 U15314 ( .A(n8899), .ZN(n8898) );
  NAND2_X1 U15316 ( .A1(n8898), .A2(n9124), .ZN(n9364) );
  NAND3_X1 U15317 ( .A1(n8036), .A2(n8035), .A3(n8038), .ZN(n8037) );
  AND2_X1 U15318 ( .A1(n29304), .A2(n8899), .ZN(n8663) );
  NAND2_X1 U15319 ( .A1(n8041), .A2(n29751), .ZN(n8146) );
  NAND2_X1 U15320 ( .A1(n8043), .A2(n8143), .ZN(n8042) );
  AOI21_X1 U15321 ( .B1(n8146), .B2(n8042), .A(n8044), .ZN(n8487) );
  NAND2_X1 U15322 ( .A1(n8043), .A2(n8141), .ZN(n8046) );
  AOI21_X1 U15324 ( .B1(n8046), .B2(n8045), .A(n8143), .ZN(n8486) );
  NAND2_X1 U15325 ( .A1(n8663), .A2(n9125), .ZN(n9365) );
  AND2_X1 U15326 ( .A1(n8048), .A2(n8047), .ZN(n8051) );
  NAND2_X1 U15327 ( .A1(n9125), .A2(n29304), .ZN(n8053) );
  OAI211_X1 U15328 ( .C1(n284), .C2(n9125), .A(n8053), .B(n3274), .ZN(n8054)
         );
  OAI211_X1 U15329 ( .C1(n3274), .C2(n9364), .A(n9365), .B(n8054), .ZN(n8055)
         );
  XNOR2_X1 U15330 ( .A(n9504), .B(n8055), .ZN(n10209) );
  NAND3_X1 U15331 ( .A1(n8431), .A2(n8351), .A3(n8353), .ZN(n8057) );
  INV_X1 U15332 ( .A(n8351), .ZN(n8428) );
  NAND3_X1 U15333 ( .A1(n8426), .A2(n8427), .A3(n8428), .ZN(n8056) );
  AND2_X1 U15334 ( .A1(n8056), .A2(n8057), .ZN(n8060) );
  NAND3_X1 U15335 ( .A1(n8430), .A2(n8428), .A3(n8058), .ZN(n8059) );
  XNOR2_X1 U15336 ( .A(n10071), .B(n1172), .ZN(n8061) );
  XNOR2_X1 U15337 ( .A(n10209), .B(n8061), .ZN(n8062) );
  INV_X1 U15338 ( .A(n284), .ZN(n8488) );
  NAND3_X1 U15339 ( .A1(n8898), .A2(n9125), .A3(n8488), .ZN(n8068) );
  NAND3_X1 U15340 ( .A1(n610), .A2(n284), .A3(n8899), .ZN(n8067) );
  NAND3_X1 U15341 ( .A1(n610), .A2(n284), .A3(n9124), .ZN(n8066) );
  NAND2_X1 U15342 ( .A1(n8899), .A2(n1793), .ZN(n8065) );
  NAND2_X1 U15343 ( .A1(n8656), .A2(n8116), .ZN(n8498) );
  NAND2_X1 U15344 ( .A1(n8498), .A2(n8502), .ZN(n8070) );
  OAI21_X1 U15345 ( .B1(n8498), .B2(n8635), .A(n8115), .ZN(n8069) );
  XNOR2_X1 U15346 ( .A(n10144), .B(n10219), .ZN(n9892) );
  INV_X1 U15347 ( .A(n9892), .ZN(n9336) );
  INV_X1 U15348 ( .A(n8669), .ZN(n9118) );
  AND2_X1 U15349 ( .A1(n8073), .A2(n8664), .ZN(n9096) );
  NAND2_X1 U15350 ( .A1(n9096), .A2(n8492), .ZN(n8076) );
  INV_X1 U15351 ( .A(n8665), .ZN(n8630) );
  INV_X1 U15352 ( .A(n8664), .ZN(n8491) );
  NAND3_X1 U15353 ( .A1(n8630), .A2(n8491), .A3(n9095), .ZN(n8075) );
  NAND3_X1 U15354 ( .A1(n8630), .A2(n8491), .A3(n8666), .ZN(n8074) );
  XNOR2_X1 U15355 ( .A(n28634), .B(n10028), .ZN(n9782) );
  XNOR2_X1 U15356 ( .A(n9336), .B(n9782), .ZN(n8090) );
  NAND2_X1 U15357 ( .A1(n8079), .A2(n8507), .ZN(n8080) );
  NAND2_X1 U15358 ( .A1(n8080), .A2(n8892), .ZN(n8083) );
  INV_X1 U15359 ( .A(n8889), .ZN(n8081) );
  INV_X1 U15360 ( .A(n8336), .ZN(n8890) );
  OAI211_X1 U15361 ( .C1(n8891), .C2(n8009), .A(n8081), .B(n8890), .ZN(n8082)
         );
  INV_X1 U15362 ( .A(n10289), .ZN(n9757) );
  XNOR2_X1 U15363 ( .A(n9992), .B(n9757), .ZN(n8088) );
  INV_X1 U15364 ( .A(n8481), .ZN(n8086) );
  NAND3_X1 U15365 ( .A1(n5674), .A2(n9013), .A3(n9014), .ZN(n8084) );
  AND3_X1 U15366 ( .A1(n8086), .A2(n8085), .A3(n8084), .ZN(n10143) );
  XNOR2_X1 U15367 ( .A(n10143), .B(n3087), .ZN(n8087) );
  XNOR2_X1 U15368 ( .A(n8088), .B(n8087), .ZN(n8089) );
  INV_X1 U15369 ( .A(n10820), .ZN(n11169) );
  NAND2_X1 U15370 ( .A1(n9238), .A2(n8544), .ZN(n8092) );
  INV_X1 U15371 ( .A(n9229), .ZN(n9237) );
  OAI21_X1 U15372 ( .B1(n9237), .B2(n9233), .A(n9232), .ZN(n8091) );
  AOI21_X1 U15374 ( .B1(n8433), .B2(n28210), .A(n9027), .ZN(n8094) );
  INV_X1 U15375 ( .A(n8526), .ZN(n8097) );
  NAND2_X1 U15376 ( .A1(n8097), .A2(n8688), .ZN(n8101) );
  NAND2_X1 U15377 ( .A1(n597), .A2(n9220), .ZN(n8100) );
  NAND2_X1 U15378 ( .A1(n8098), .A2(n597), .ZN(n8099) );
  NAND4_X2 U15379 ( .A1(n8102), .A2(n8101), .A3(n8099), .A4(n8100), .ZN(n9929)
         );
  INV_X1 U15382 ( .A(n8104), .ZN(n8105) );
  NAND2_X1 U15383 ( .A1(n8105), .A2(n9061), .ZN(n8106) );
  OAI211_X1 U15384 ( .C1(n8395), .C2(n9062), .A(n8107), .B(n8106), .ZN(n9963)
         );
  XNOR2_X1 U15385 ( .A(n9963), .B(n9929), .ZN(n8108) );
  XNOR2_X1 U15386 ( .A(n10123), .B(n8108), .ZN(n8126) );
  AND2_X1 U15387 ( .A1(n8109), .A2(n8693), .ZN(n9246) );
  INV_X1 U15388 ( .A(n9246), .ZN(n8114) );
  NAND2_X1 U15389 ( .A1(n8110), .A2(n9247), .ZN(n8111) );
  NAND2_X1 U15390 ( .A1(n8111), .A2(n9245), .ZN(n8113) );
  AND2_X1 U15391 ( .A1(n9247), .A2(n9243), .ZN(n9412) );
  NAND2_X1 U15392 ( .A1(n9412), .A2(n8693), .ZN(n8112) );
  OAI211_X2 U15393 ( .C1(n8114), .C2(n9245), .A(n8113), .B(n8112), .ZN(n10304)
         );
  XNOR2_X1 U15394 ( .A(n10009), .B(n10304), .ZN(n8124) );
  INV_X1 U15395 ( .A(n8427), .ZN(n8119) );
  AOI21_X1 U15396 ( .B1(n8119), .B2(n1910), .A(n8426), .ZN(n8122) );
  NAND2_X1 U15397 ( .A1(n8120), .A2(n8353), .ZN(n8121) );
  XNOR2_X1 U15398 ( .A(n10088), .B(n2602), .ZN(n8123) );
  XNOR2_X1 U15399 ( .A(n8124), .B(n8123), .ZN(n8125) );
  INV_X1 U15400 ( .A(n11330), .ZN(n11331) );
  INV_X1 U15402 ( .A(n8817), .ZN(n8976) );
  INV_X1 U15403 ( .A(n8593), .ZN(n8974) );
  INV_X1 U15404 ( .A(n8592), .ZN(n8591) );
  NAND3_X1 U15405 ( .A1(n8974), .A2(n607), .A3(n8591), .ZN(n8128) );
  NAND3_X1 U15406 ( .A1(n8977), .A2(n8819), .A3(n8594), .ZN(n8127) );
  AOI21_X1 U15407 ( .B1(n8135), .B2(n8134), .A(n8133), .ZN(n8137) );
  NAND2_X1 U15408 ( .A1(n8139), .A2(n8138), .ZN(n8140) );
  NAND3_X1 U15409 ( .A1(n8146), .A2(n8141), .A3(n8140), .ZN(n8145) );
  NAND3_X1 U15410 ( .A1(n8143), .A2(n7336), .A3(n8142), .ZN(n8144) );
  OAI211_X1 U15411 ( .C1(n8146), .C2(n7336), .A(n8145), .B(n8144), .ZN(n9396)
         );
  NAND2_X1 U15412 ( .A1(n8981), .A2(n9396), .ZN(n9398) );
  NAND2_X1 U15413 ( .A1(n8147), .A2(n8150), .ZN(n8149) );
  OAI211_X1 U15414 ( .C1(n28149), .C2(n1607), .A(n8149), .B(n8148), .ZN(n8152)
         );
  AND2_X1 U15415 ( .A1(n8153), .A2(n7550), .ZN(n8157) );
  NAND3_X1 U15416 ( .A1(n8162), .A2(n8161), .A3(n8160), .ZN(n8163) );
  NAND2_X1 U15418 ( .A1(n8166), .A2(n8165), .ZN(n8170) );
  AOI21_X1 U15420 ( .B1(n8170), .B2(n8169), .A(n8168), .ZN(n8171) );
  INV_X1 U15421 ( .A(n8176), .ZN(n8178) );
  NAND3_X1 U15422 ( .A1(n8173), .A2(n7760), .A3(n8178), .ZN(n8174) );
  NAND2_X1 U15423 ( .A1(n8175), .A2(n8174), .ZN(n8183) );
  NAND2_X1 U15424 ( .A1(n8177), .A2(n8176), .ZN(n8181) );
  INV_X1 U15425 ( .A(n8980), .ZN(n8644) );
  NAND3_X1 U15426 ( .A1(n8644), .A2(n596), .A3(n8982), .ZN(n8184) );
  INV_X1 U15427 ( .A(n9144), .ZN(n8561) );
  NAND2_X1 U15428 ( .A1(n8561), .A2(n8185), .ZN(n8186) );
  INV_X1 U15429 ( .A(n8563), .ZN(n9142) );
  NAND3_X1 U15430 ( .A1(n8561), .A2(n598), .A3(n9142), .ZN(n8188) );
  XNOR2_X1 U15431 ( .A(n9295), .B(n3770), .ZN(n8191) );
  XNOR2_X1 U15432 ( .A(n9770), .B(n8191), .ZN(n8319) );
  NAND2_X1 U15433 ( .A1(n8829), .A2(n8827), .ZN(n8198) );
  NAND2_X1 U15434 ( .A1(n8829), .A2(n8192), .ZN(n8195) );
  OAI21_X1 U15435 ( .B1(n8829), .B2(n8193), .A(n8826), .ZN(n8194) );
  OAI211_X1 U15436 ( .C1(n8196), .C2(n8826), .A(n8195), .B(n8194), .ZN(n8197)
         );
  NAND2_X1 U15437 ( .A1(n8203), .A2(n8205), .ZN(n8204) );
  NOR2_X1 U15438 ( .A1(n8836), .A2(n8838), .ZN(n9169) );
  INV_X1 U15439 ( .A(n8838), .ZN(n8229) );
  AOI21_X1 U15441 ( .B1(n8218), .B2(n8217), .A(n8216), .ZN(n8219) );
  OR2_X2 U15442 ( .A1(n8220), .A2(n8219), .ZN(n9171) );
  MUX2_X1 U15443 ( .A(n3821), .B(n8222), .S(n8221), .Z(n8228) );
  INV_X1 U15444 ( .A(n8230), .ZN(n8964) );
  OAI21_X1 U15445 ( .B1(n8229), .B2(n9171), .A(n8964), .ZN(n8250) );
  NAND2_X1 U15446 ( .A1(n8233), .A2(n8232), .ZN(n8241) );
  NAND2_X1 U15448 ( .A1(n8236), .A2(n8235), .ZN(n8238) );
  MUX2_X1 U15449 ( .A(n8239), .B(n8238), .S(n29110), .Z(n8240) );
  NAND3_X1 U15450 ( .A1(n8961), .A2(n9171), .A3(n9170), .ZN(n8249) );
  INV_X1 U15451 ( .A(n8836), .ZN(n8962) );
  NAND3_X1 U15452 ( .A1(n8962), .A2(n605), .A3(n8837), .ZN(n8248) );
  XNOR2_X1 U15453 ( .A(n10060), .B(n10178), .ZN(n9845) );
  NAND2_X1 U15454 ( .A1(n8521), .A2(n8811), .ZN(n8251) );
  AND2_X1 U15455 ( .A1(n8253), .A2(n8252), .ZN(n8254) );
  MUX2_X1 U15456 ( .A(n8257), .B(n28615), .S(n8258), .Z(n8262) );
  MUX2_X1 U15457 ( .A(n8260), .B(n8259), .S(n8258), .Z(n8261) );
  INV_X1 U15459 ( .A(n8954), .ZN(n8471) );
  INV_X1 U15460 ( .A(n8266), .ZN(n8274) );
  NAND2_X1 U15461 ( .A1(n8272), .A2(n8271), .ZN(n8273) );
  NAND2_X1 U15462 ( .A1(n8471), .A2(n8958), .ZN(n9167) );
  INV_X1 U15463 ( .A(n8275), .ZN(n8278) );
  INV_X1 U15464 ( .A(n8280), .ZN(n8282) );
  INV_X1 U15465 ( .A(n8956), .ZN(n9163) );
  INV_X1 U15466 ( .A(n8286), .ZN(n8289) );
  NAND2_X1 U15467 ( .A1(n7915), .A2(n8287), .ZN(n8288) );
  NAND2_X1 U15469 ( .A1(n8291), .A2(n7915), .ZN(n8293) );
  NAND3_X1 U15472 ( .A1(n8302), .A2(n8301), .A3(n29317), .ZN(n8307) );
  OAI211_X1 U15473 ( .C1(n9160), .C2(n8958), .A(n9162), .B(n29096), .ZN(n8317)
         );
  INV_X1 U15474 ( .A(n8958), .ZN(n9164) );
  NAND2_X1 U15475 ( .A1(n8308), .A2(n28810), .ZN(n8309) );
  AOI21_X1 U15476 ( .B1(n8310), .B2(n8309), .A(n7614), .ZN(n8315) );
  NAND3_X1 U15477 ( .A1(n7934), .A2(n28810), .A3(n7933), .ZN(n8313) );
  NAND3_X1 U15478 ( .A1(n8311), .A2(n7614), .A3(n7933), .ZN(n8312) );
  NAND2_X1 U15479 ( .A1(n8313), .A2(n8312), .ZN(n8314) );
  INV_X1 U15480 ( .A(n8802), .ZN(n9161) );
  INV_X1 U15481 ( .A(n8955), .ZN(n8800) );
  XNOR2_X1 U15482 ( .A(n28488), .B(n10059), .ZN(n9549) );
  XNOR2_X1 U15483 ( .A(n9845), .B(n9549), .ZN(n8318) );
  NOR2_X1 U15485 ( .A1(n9531), .A2(n9532), .ZN(n8322) );
  OAI21_X1 U15486 ( .B1(n9532), .B2(n8749), .A(n8747), .ZN(n8321) );
  NOR2_X1 U15488 ( .A1(n8610), .A2(n9530), .ZN(n8323) );
  NAND2_X1 U15489 ( .A1(n8323), .A2(n9531), .ZN(n9537) );
  NAND2_X1 U15491 ( .A1(n7569), .A2(n8579), .ZN(n8575) );
  INV_X1 U15494 ( .A(n9323), .ZN(n9870) );
  XNOR2_X1 U15495 ( .A(n10033), .B(n9870), .ZN(n10055) );
  NAND2_X1 U15496 ( .A1(n598), .A2(n8563), .ZN(n8560) );
  OAI21_X1 U15497 ( .B1(n8762), .B2(n8941), .A(n8764), .ZN(n8331) );
  XNOR2_X1 U15498 ( .A(n10055), .B(n9736), .ZN(n8348) );
  NAND3_X1 U15499 ( .A1(n8760), .A2(n9148), .A3(n9146), .ZN(n8333) );
  OAI21_X1 U15500 ( .B1(n8334), .B2(n8336), .A(n8009), .ZN(n8339) );
  NAND3_X1 U15501 ( .A1(n8507), .A2(n8336), .A3(n8335), .ZN(n8338) );
  NAND3_X1 U15502 ( .A1(n8507), .A2(n8504), .A3(n8891), .ZN(n8337) );
  XNOR2_X1 U15503 ( .A(n10171), .B(n9698), .ZN(n8346) );
  AOI21_X1 U15504 ( .B1(n8341), .B2(n8340), .A(n7410), .ZN(n8344) );
  XNOR2_X1 U15505 ( .A(n10138), .B(n5059), .ZN(n8345) );
  XNOR2_X1 U15506 ( .A(n8346), .B(n8345), .ZN(n8347) );
  XNOR2_X1 U15507 ( .A(n8348), .B(n8347), .ZN(n10467) );
  INV_X1 U15509 ( .A(n9186), .ZN(n9004) );
  OAI21_X1 U15510 ( .B1(n8445), .B2(n9186), .A(n8782), .ZN(n8350) );
  NOR2_X1 U15512 ( .A1(n8353), .A2(n1909), .ZN(n8355) );
  INV_X1 U15513 ( .A(n9202), .ZN(n8448) );
  NOR2_X1 U15514 ( .A1(n9196), .A2(n28862), .ZN(n8357) );
  OAI21_X1 U15515 ( .B1(n6897), .B2(n8357), .A(n8448), .ZN(n8359) );
  OAI21_X1 U15517 ( .B1(n9028), .B2(n8792), .A(n9030), .ZN(n8361) );
  XNOR2_X1 U15518 ( .A(n10183), .B(n9948), .ZN(n10157) );
  XNOR2_X1 U15519 ( .A(n9748), .B(n10157), .ZN(n8377) );
  NAND2_X1 U15521 ( .A1(n9435), .A2(n9434), .ZN(n8364) );
  OAI211_X1 U15522 ( .C1(n9434), .C2(n9208), .A(n8364), .B(n9210), .ZN(n8365)
         );
  NAND2_X1 U15523 ( .A1(n9437), .A2(n8365), .ZN(n8368) );
  NAND2_X1 U15524 ( .A1(n8718), .A2(n8787), .ZN(n8366) );
  INV_X1 U15525 ( .A(n8787), .ZN(n8439) );
  XNOR2_X1 U15526 ( .A(n9823), .B(n8368), .ZN(n10068) );
  INV_X1 U15527 ( .A(n8369), .ZN(n8738) );
  INV_X1 U15529 ( .A(n8733), .ZN(n8370) );
  NAND3_X1 U15530 ( .A1(n8730), .A2(n8370), .A3(n8734), .ZN(n8372) );
  NAND3_X1 U15531 ( .A1(n8739), .A2(n8370), .A3(n8381), .ZN(n8371) );
  XNOR2_X1 U15532 ( .A(n1895), .B(n3607), .ZN(n8375) );
  XNOR2_X1 U15533 ( .A(n8375), .B(n10068), .ZN(n8376) );
  NAND3_X1 U15534 ( .A1(n11331), .A2(n11166), .A3(n11168), .ZN(n8424) );
  OAI21_X1 U15536 ( .B1(n8378), .B2(n8741), .A(n9070), .ZN(n8379) );
  NAND2_X1 U15537 ( .A1(n8537), .A2(n8381), .ZN(n8382) );
  OAI21_X1 U15538 ( .B1(n8384), .B2(n8537), .A(n8382), .ZN(n8383) );
  NAND2_X1 U15539 ( .A1(n8383), .A2(n8735), .ZN(n8387) );
  NAND3_X1 U15540 ( .A1(n8384), .A2(n8536), .A3(n8733), .ZN(n8386) );
  NAND3_X1 U15541 ( .A1(n8731), .A2(n8739), .A3(n8729), .ZN(n8385) );
  XNOR2_X1 U15542 ( .A(n10074), .B(n10207), .ZN(n9850) );
  NAND2_X1 U15543 ( .A1(n29311), .A2(n2320), .ZN(n8391) );
  NAND2_X1 U15544 ( .A1(n9080), .A2(n8605), .ZN(n10240) );
  OAI211_X1 U15545 ( .C1(n29311), .C2(n28500), .A(n10240), .B(n8848), .ZN(
        n8389) );
  INV_X1 U15546 ( .A(n8848), .ZN(n9079) );
  OAI21_X1 U15547 ( .B1(n29311), .B2(n8726), .A(n9079), .ZN(n8388) );
  NAND2_X1 U15548 ( .A1(n8389), .A2(n8388), .ZN(n8390) );
  OAI21_X1 U15549 ( .B1(n8724), .B2(n8391), .A(n8390), .ZN(n9509) );
  INV_X1 U15550 ( .A(n9509), .ZN(n9368) );
  INV_X1 U15551 ( .A(n9064), .ZN(n8392) );
  NAND2_X1 U15552 ( .A1(n8392), .A2(n8397), .ZN(n8598) );
  NAND2_X1 U15555 ( .A1(n8396), .A2(n9062), .ZN(n8401) );
  NAND3_X1 U15556 ( .A1(n9060), .A2(n8864), .A3(n9059), .ZN(n8400) );
  NAND2_X1 U15557 ( .A1(n9064), .A2(n8397), .ZN(n9063) );
  INV_X1 U15558 ( .A(n9063), .ZN(n8398) );
  NAND2_X1 U15559 ( .A1(n8398), .A2(n9060), .ZN(n8399) );
  NAND4_X1 U15560 ( .A1(n8402), .A2(n8401), .A3(n8400), .A4(n8399), .ZN(n9592)
         );
  XNOR2_X1 U15561 ( .A(n9592), .B(n9368), .ZN(n9943) );
  XNOR2_X1 U15562 ( .A(n9850), .B(n9943), .ZN(n8421) );
  NAND2_X1 U15563 ( .A1(n8709), .A2(n8877), .ZN(n8708) );
  OR2_X1 U15564 ( .A1(n8708), .A2(n8873), .ZN(n8406) );
  NAND2_X1 U15565 ( .A1(n8875), .A2(n8881), .ZN(n8712) );
  OR2_X1 U15566 ( .A1(n8712), .A2(n8874), .ZN(n8405) );
  XNOR2_X1 U15567 ( .A(n10128), .B(n3493), .ZN(n8419) );
  MUX2_X1 U15568 ( .A(n8642), .B(n8984), .S(n8980), .Z(n8411) );
  OR2_X1 U15569 ( .A1(n9396), .A2(n8981), .ZN(n9177) );
  OAI21_X1 U15570 ( .B1(n8644), .B2(n8982), .A(n8981), .ZN(n8409) );
  NAND2_X1 U15573 ( .A1(n8413), .A2(n4321), .ZN(n8417) );
  INV_X1 U15574 ( .A(n8788), .ZN(n8440) );
  NAND3_X1 U15575 ( .A1(n8440), .A2(n8720), .A3(n8787), .ZN(n8416) );
  INV_X1 U15576 ( .A(n8719), .ZN(n8786) );
  NAND3_X1 U15577 ( .A1(n8717), .A2(n8786), .A3(n8414), .ZN(n8415) );
  XNOR2_X1 U15578 ( .A(n8419), .B(n8418), .ZN(n8420) );
  XNOR2_X1 U15579 ( .A(n8421), .B(n8420), .ZN(n10821) );
  INV_X1 U15580 ( .A(n9392), .ZN(n9614) );
  MUX2_X1 U15581 ( .A(n9027), .B(n9028), .S(n8433), .Z(n8434) );
  INV_X1 U15582 ( .A(n10295), .ZN(n10034) );
  XNOR2_X1 U15583 ( .A(n10034), .B(n9614), .ZN(n8444) );
  MUX2_X1 U15584 ( .A(n9211), .B(n9434), .S(n8777), .Z(n8437) );
  XNOR2_X1 U15586 ( .A(n9735), .B(n1920), .ZN(n8443) );
  XNOR2_X1 U15587 ( .A(n8444), .B(n8443), .ZN(n8455) );
  MUX2_X1 U15588 ( .A(n9009), .B(n9007), .S(n9184), .Z(n8447) );
  MUX2_X1 U15589 ( .A(n9184), .B(n9186), .S(n8445), .Z(n8446) );
  NOR2_X1 U15591 ( .A1(n329), .A2(n9200), .ZN(n8451) );
  NAND2_X1 U15592 ( .A1(n9199), .A2(n28862), .ZN(n8450) );
  XNOR2_X1 U15593 ( .A(n10298), .B(n10038), .ZN(n8453) );
  XNOR2_X1 U15594 ( .A(n1902), .B(n1184), .ZN(n8452) );
  XNOR2_X1 U15595 ( .A(n8453), .B(n8452), .ZN(n8454) );
  INV_X1 U15596 ( .A(n10748), .ZN(n11198) );
  AOI21_X1 U15597 ( .B1(n8456), .B2(n8980), .A(n8983), .ZN(n9399) );
  INV_X1 U15598 ( .A(n9399), .ZN(n8458) );
  NAND2_X1 U15599 ( .A1(n8642), .A2(n8980), .ZN(n9397) );
  OAI21_X1 U15600 ( .B1(n436), .B2(n596), .A(n9397), .ZN(n9179) );
  NAND2_X1 U15601 ( .A1(n9179), .A2(n9396), .ZN(n8457) );
  NAND2_X1 U15602 ( .A1(n8458), .A2(n8457), .ZN(n9656) );
  NAND2_X1 U15603 ( .A1(n8681), .A2(n8809), .ZN(n8459) );
  NAND2_X1 U15604 ( .A1(n8810), .A2(n8809), .ZN(n8460) );
  XNOR2_X1 U15605 ( .A(n9930), .B(n9656), .ZN(n8469) );
  INV_X1 U15606 ( .A(n8827), .ZN(n8825) );
  XNOR2_X1 U15607 ( .A(n9964), .B(n3386), .ZN(n8468) );
  XNOR2_X1 U15608 ( .A(n8469), .B(n8468), .ZN(n8480) );
  AOI22_X1 U15609 ( .A1(n8964), .A2(n9171), .B1(n8838), .B2(n8966), .ZN(n9174)
         );
  AND2_X1 U15610 ( .A1(n8836), .A2(n8838), .ZN(n8967) );
  OAI21_X1 U15611 ( .B1(n8967), .B2(n8837), .A(n8961), .ZN(n8470) );
  NAND2_X1 U15612 ( .A1(n8954), .A2(n8956), .ZN(n8805) );
  OAI21_X1 U15613 ( .B1(n8472), .B2(n9161), .A(n8471), .ZN(n8474) );
  NAND3_X1 U15614 ( .A1(n8801), .A2(n8802), .A3(n8956), .ZN(n8473) );
  OAI211_X1 U15615 ( .C1(n9164), .C2(n8805), .A(n8474), .B(n8473), .ZN(n10008)
         );
  XNOR2_X1 U15616 ( .A(n28616), .B(n10263), .ZN(n10306) );
  INV_X1 U15618 ( .A(n10193), .ZN(n8476) );
  XNOR2_X1 U15619 ( .A(n8476), .B(n10302), .ZN(n8477) );
  NAND2_X1 U15621 ( .A1(n11198), .A2(n28157), .ZN(n8623) );
  AOI22_X1 U15622 ( .A1(n8481), .A2(n9013), .B1(n9018), .B2(n8662), .ZN(n8484)
         );
  NAND2_X1 U15623 ( .A1(n284), .A2(n29304), .ZN(n8485) );
  OAI21_X1 U15624 ( .B1(n8664), .B2(n8665), .A(n8490), .ZN(n8496) );
  OR2_X1 U15626 ( .A1(n8500), .A2(n8499), .ZN(n8654) );
  NAND2_X1 U15627 ( .A1(n8634), .A2(n8653), .ZN(n8503) );
  INV_X1 U15628 ( .A(n9430), .ZN(n9976) );
  XNOR2_X1 U15629 ( .A(n9976), .B(n9771), .ZN(n9924) );
  NAND2_X1 U15630 ( .A1(n8009), .A2(n8889), .ZN(n8505) );
  AOI21_X1 U15631 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8510) );
  OAI21_X1 U15632 ( .B1(n8892), .B2(n8887), .A(n8508), .ZN(n8509) );
  NAND3_X1 U15634 ( .A1(n8916), .A2(n8512), .A3(n8511), .ZN(n8516) );
  NAND3_X1 U15635 ( .A1(n9106), .A2(n8513), .A3(n8917), .ZN(n8515) );
  NAND3_X2 U15636 ( .A1(n8515), .A2(n8516), .A3(n8514), .ZN(n10021) );
  XNOR2_X1 U15637 ( .A(n9678), .B(n10021), .ZN(n8518) );
  XNOR2_X1 U15638 ( .A(n9550), .B(n3211), .ZN(n8517) );
  XNOR2_X1 U15639 ( .A(n8518), .B(n8517), .ZN(n8519) );
  INV_X1 U15641 ( .A(n28638), .ZN(n10751) );
  NAND2_X1 U15642 ( .A1(n9224), .A2(n8687), .ZN(n8527) );
  NAND2_X1 U15643 ( .A1(n9228), .A2(n8687), .ZN(n8528) );
  XNOR2_X1 U15644 ( .A(n9991), .B(n9755), .ZN(n9936) );
  INV_X1 U15645 ( .A(n9412), .ZN(n8530) );
  INV_X1 U15646 ( .A(n9244), .ZN(n8529) );
  OAI21_X1 U15647 ( .B1(n8693), .B2(n8109), .A(n8529), .ZN(n9414) );
  NAND2_X1 U15648 ( .A1(n9410), .A2(n8109), .ZN(n9409) );
  OAI211_X1 U15649 ( .C1(n8530), .C2(n8109), .A(n9414), .B(n9409), .ZN(n8535)
         );
  AOI21_X1 U15650 ( .B1(n8404), .B2(n8874), .A(n8873), .ZN(n8534) );
  AND2_X1 U15651 ( .A1(n8873), .A2(n8881), .ZN(n8878) );
  INV_X1 U15652 ( .A(n8874), .ZN(n8531) );
  NAND3_X1 U15653 ( .A1(n8532), .A2(n8403), .A3(n8531), .ZN(n8533) );
  OAI21_X1 U15654 ( .B1(n8534), .B2(n8878), .A(n8533), .ZN(n9717) );
  XNOR2_X1 U15655 ( .A(n8535), .B(n9717), .ZN(n10291) );
  XNOR2_X1 U15656 ( .A(n9936), .B(n10291), .ZN(n8548) );
  NOR2_X1 U15657 ( .A1(n8537), .A2(n8734), .ZN(n8540) );
  OAI211_X1 U15659 ( .C1(n9045), .C2(n9047), .A(n9237), .B(n9233), .ZN(n8543)
         );
  OAI211_X1 U15660 ( .C1(n8544), .C2(n9045), .A(n8543), .B(n9238), .ZN(n10029)
         );
  XNOR2_X1 U15661 ( .A(n9626), .B(n10029), .ZN(n8546) );
  XNOR2_X1 U15662 ( .A(n9447), .B(n3336), .ZN(n8545) );
  XNOR2_X1 U15663 ( .A(n8546), .B(n8545), .ZN(n8547) );
  XNOR2_X1 U15664 ( .A(n8548), .B(n8547), .ZN(n10747) );
  INV_X1 U15665 ( .A(n10747), .ZN(n11197) );
  INV_X1 U15666 ( .A(n8550), .ZN(n9137) );
  INV_X1 U15667 ( .A(n9340), .ZN(n8924) );
  MUX2_X1 U15668 ( .A(n8550), .B(n8549), .S(n7410), .Z(n8551) );
  XNOR2_X1 U15669 ( .A(n9851), .B(n9504), .ZN(n8559) );
  NAND2_X1 U15670 ( .A1(n8553), .A2(n8941), .ZN(n8554) );
  NAND3_X1 U15671 ( .A1(n8557), .A2(n8765), .A3(n8554), .ZN(n8556) );
  NAND3_X1 U15672 ( .A1(n8945), .A2(n9562), .A3(n10401), .ZN(n8555) );
  OAI211_X1 U15673 ( .C1(n8557), .C2(n8945), .A(n8556), .B(n8555), .ZN(n10434)
         );
  XNOR2_X1 U15674 ( .A(n10434), .B(n3457), .ZN(n8558) );
  XNOR2_X1 U15675 ( .A(n8559), .B(n8558), .ZN(n8573) );
  NAND3_X1 U15676 ( .A1(n9144), .A2(n8563), .A3(n9139), .ZN(n8566) );
  INV_X1 U15677 ( .A(n8185), .ZN(n8564) );
  INV_X1 U15678 ( .A(n10436), .ZN(n8572) );
  INV_X1 U15679 ( .A(n9149), .ZN(n8931) );
  NAND2_X1 U15680 ( .A1(n8760), .A2(n8931), .ZN(n9152) );
  OAI211_X1 U15681 ( .C1(n8570), .C2(n8760), .A(n8930), .B(n9152), .ZN(n9378)
         );
  XNOR2_X1 U15682 ( .A(n8572), .B(n10311), .ZN(n9668) );
  AND2_X1 U15683 ( .A1(n8574), .A2(n603), .ZN(n9419) );
  INV_X1 U15684 ( .A(n9531), .ZN(n8751) );
  XNOR2_X1 U15685 ( .A(n9763), .B(n10359), .ZN(n9940) );
  NAND2_X1 U15686 ( .A1(n8580), .A2(n8579), .ZN(n8583) );
  OAI21_X1 U15687 ( .B1(n8828), .B2(n8826), .A(n8824), .ZN(n8585) );
  AOI22_X1 U15688 ( .A1(n8585), .A2(n8584), .B1(n1839), .B2(n8828), .ZN(n8588)
         );
  OR2_X1 U15689 ( .A1(n8588), .A2(n8587), .ZN(n9645) );
  XNOR2_X1 U15690 ( .A(n9645), .B(n1878), .ZN(n8602) );
  NAND2_X1 U15691 ( .A1(n8977), .A2(n8589), .ZN(n8973) );
  NAND2_X1 U15692 ( .A1(n8594), .A2(n8978), .ZN(n8590) );
  NAND2_X1 U15694 ( .A1(n8591), .A2(n8817), .ZN(n8595) );
  NAND2_X1 U15695 ( .A1(n8593), .A2(n8592), .ZN(n8818) );
  OAI21_X1 U15696 ( .B1(n8595), .B2(n8594), .A(n8818), .ZN(n8596) );
  NAND3_X1 U15697 ( .A1(n9064), .A2(n8872), .A3(n8865), .ZN(n8599) );
  AND2_X1 U15698 ( .A1(n8599), .A2(n8598), .ZN(n8600) );
  XNOR2_X1 U15699 ( .A(n10285), .B(n8602), .ZN(n8621) );
  NOR2_X1 U15700 ( .A1(n9080), .A2(n8603), .ZN(n10234) );
  NAND2_X1 U15701 ( .A1(n10234), .A2(n8724), .ZN(n8604) );
  OAI21_X1 U15702 ( .B1(n8724), .B2(n10240), .A(n8604), .ZN(n10245) );
  NAND2_X1 U15703 ( .A1(n8848), .A2(n28500), .ZN(n10237) );
  INV_X1 U15704 ( .A(n10237), .ZN(n8607) );
  OR3_X2 U15705 ( .A1(n10245), .A2(n8607), .A3(n8606), .ZN(n9749) );
  NAND2_X1 U15706 ( .A1(n8610), .A2(n9530), .ZN(n8752) );
  NAND3_X1 U15707 ( .A1(n9531), .A2(n8609), .A3(n9530), .ZN(n8613) );
  INV_X1 U15709 ( .A(n8857), .ZN(n8742) );
  NAND2_X1 U15710 ( .A1(n9075), .A2(n9070), .ZN(n8616) );
  NAND2_X1 U15711 ( .A1(n9075), .A2(n8857), .ZN(n8615) );
  NAND2_X1 U15712 ( .A1(n9071), .A2(n8740), .ZN(n8614) );
  NAND4_X1 U15713 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8614), .ZN(n8618)
         );
  XNOR2_X1 U15714 ( .A(n10043), .B(n3662), .ZN(n8619) );
  XNOR2_X1 U15715 ( .A(n9946), .B(n8619), .ZN(n8620) );
  NAND3_X1 U15716 ( .A1(n3585), .A2(n10563), .A3(n28207), .ZN(n8622) );
  NAND2_X1 U15718 ( .A1(n8802), .A2(n8955), .ZN(n8804) );
  XNOR2_X1 U15719 ( .A(n9306), .B(n1246), .ZN(n8626) );
  XNOR2_X1 U15720 ( .A(n8626), .B(n1877), .ZN(n8639) );
  INV_X1 U15721 ( .A(n9095), .ZN(n8627) );
  NAND3_X1 U15723 ( .A1(n9099), .A2(n8627), .A3(n8666), .ZN(n8628) );
  NAND2_X1 U15724 ( .A1(n8629), .A2(n8628), .ZN(n8633) );
  AOI21_X1 U15725 ( .B1(n8631), .B2(n9100), .A(n8630), .ZN(n8632) );
  NAND2_X1 U15726 ( .A1(n8634), .A2(n8635), .ZN(n8638) );
  NAND3_X1 U15727 ( .A1(n8635), .A2(n8656), .A3(n8655), .ZN(n8637) );
  NAND3_X1 U15728 ( .A1(n8653), .A2(n8652), .A3(n8658), .ZN(n8636) );
  XNOR2_X1 U15729 ( .A(n9986), .B(n10160), .ZN(n8904) );
  XNOR2_X1 U15730 ( .A(n8904), .B(n8639), .ZN(n8649) );
  NAND2_X1 U15731 ( .A1(n8836), .A2(n8966), .ZN(n8842) );
  NAND3_X1 U15732 ( .A1(n8963), .A2(n8962), .A3(n8838), .ZN(n8641) );
  NAND2_X1 U15733 ( .A1(n8836), .A2(n9171), .ZN(n8965) );
  NAND2_X1 U15734 ( .A1(n8982), .A2(n8642), .ZN(n8643) );
  AOI21_X1 U15735 ( .B1(n9398), .B2(n8644), .A(n8982), .ZN(n8645) );
  XNOR2_X1 U15736 ( .A(n9746), .B(n10184), .ZN(n8648) );
  OAI21_X1 U15737 ( .B1(n9566), .B2(n9561), .A(n8943), .ZN(n10403) );
  NAND2_X1 U15738 ( .A1(n10403), .A2(n8944), .ZN(n10407) );
  INV_X1 U15741 ( .A(n10283), .ZN(n8647) );
  OAI211_X1 U15742 ( .C1(n1966), .C2(n12202), .A(n11438), .B(n8650), .ZN(n9259) );
  OAI21_X1 U15743 ( .B1(n8656), .B2(n8655), .A(n8654), .ZN(n8657) );
  INV_X1 U15744 ( .A(n8657), .ZN(n8659) );
  XNOR2_X1 U15745 ( .A(n9614), .B(n9915), .ZN(n9660) );
  XNOR2_X1 U15746 ( .A(n10134), .B(n9696), .ZN(n10255) );
  XNOR2_X1 U15747 ( .A(n9660), .B(n10255), .ZN(n8677) );
  NAND2_X1 U15748 ( .A1(n8665), .A2(n8664), .ZN(n9098) );
  OAI21_X1 U15749 ( .B1(n9100), .B2(n8665), .A(n9098), .ZN(n8667) );
  MUX2_X1 U15750 ( .A(n8670), .B(n8669), .S(n8914), .Z(n8674) );
  MUX2_X1 U15751 ( .A(n8672), .B(n8671), .S(n8914), .Z(n8673) );
  XNOR2_X1 U15752 ( .A(n10133), .B(n10257), .ZN(n9831) );
  XNOR2_X1 U15753 ( .A(n9698), .B(n3191), .ZN(n8675) );
  XNOR2_X1 U15754 ( .A(n9831), .B(n8675), .ZN(n8676) );
  XNOR2_X1 U15755 ( .A(n8676), .B(n8677), .ZN(n10558) );
  NAND2_X1 U15756 ( .A1(n8810), .A2(n8811), .ZN(n8678) );
  AOI21_X1 U15757 ( .B1(n8679), .B2(n8678), .A(n8812), .ZN(n8684) );
  NAND2_X1 U15758 ( .A1(n8680), .A2(n8809), .ZN(n8682) );
  OAI21_X1 U15760 ( .B1(n8682), .B2(n8810), .A(n8814), .ZN(n8683) );
  XNOR2_X1 U15761 ( .A(n9645), .B(n9949), .ZN(n8692) );
  NAND3_X1 U15762 ( .A1(n8685), .A2(n9221), .A3(n9222), .ZN(n8690) );
  NAND3_X1 U15763 ( .A1(n8688), .A2(n8687), .A3(n8686), .ZN(n8689) );
  NAND3_X1 U15764 ( .A1(n9230), .A2(n9233), .A3(n9229), .ZN(n8691) );
  XNOR2_X1 U15765 ( .A(n8692), .B(n9603), .ZN(n8707) );
  NAND2_X1 U15766 ( .A1(n9042), .A2(n8693), .ZN(n8696) );
  NAND2_X1 U15767 ( .A1(n9041), .A2(n9247), .ZN(n8695) );
  XNOR2_X1 U15768 ( .A(n10330), .B(n10232), .ZN(n9304) );
  INV_X1 U15769 ( .A(n9304), .ZN(n8705) );
  INV_X1 U15770 ( .A(n8877), .ZN(n8698) );
  NAND2_X1 U15771 ( .A1(n8878), .A2(n8698), .ZN(n8703) );
  NAND2_X1 U15772 ( .A1(n8404), .A2(n8699), .ZN(n8702) );
  NAND3_X1 U15773 ( .A1(n8403), .A2(n8698), .A3(n8874), .ZN(n8701) );
  NAND3_X1 U15774 ( .A1(n8873), .A2(n8699), .A3(n8877), .ZN(n8700) );
  XNOR2_X1 U15775 ( .A(n10231), .B(n3180), .ZN(n8704) );
  XNOR2_X1 U15776 ( .A(n8705), .B(n8704), .ZN(n8706) );
  NAND3_X1 U15777 ( .A1(n8404), .A2(n8874), .A3(n8877), .ZN(n8711) );
  NAND2_X1 U15778 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  XNOR2_X1 U15780 ( .A(n9963), .B(n8715), .ZN(n9705) );
  NAND2_X1 U15781 ( .A1(n8719), .A2(n8718), .ZN(n8722) );
  AOI21_X1 U15782 ( .B1(n8722), .B2(n4321), .A(n8720), .ZN(n8723) );
  NAND2_X1 U15783 ( .A1(n8848), .A2(n8726), .ZN(n8725) );
  AOI21_X1 U15784 ( .B1(n8850), .B2(n8725), .A(n8724), .ZN(n8728) );
  NAND2_X1 U15785 ( .A1(n28500), .A2(n8726), .ZN(n9078) );
  AOI21_X1 U15786 ( .B1(n9078), .B2(n8848), .A(n29311), .ZN(n8727) );
  XNOR2_X1 U15787 ( .A(n10264), .B(n9877), .ZN(n9817) );
  XNOR2_X1 U15788 ( .A(n9705), .B(n9817), .ZN(n8746) );
  NOR2_X1 U15789 ( .A1(n8730), .A2(n8729), .ZN(n8732) );
  OAI21_X1 U15790 ( .B1(n8732), .B2(n8731), .A(n8739), .ZN(n8737) );
  AOI22_X1 U15791 ( .A1(n8856), .A2(n9075), .B1(n8740), .B2(n8741), .ZN(n8743)
         );
  XNOR2_X1 U15792 ( .A(n9931), .B(n10265), .ZN(n9742) );
  XNOR2_X1 U15793 ( .A(n9656), .B(n3323), .ZN(n8744) );
  XNOR2_X1 U15794 ( .A(n9742), .B(n8744), .ZN(n8745) );
  MUX2_X1 U15795 ( .A(n11345), .B(n1898), .S(n11334), .Z(n8846) );
  NAND3_X1 U15796 ( .A1(n9529), .A2(n29395), .A3(n29662), .ZN(n8750) );
  NAND2_X1 U15797 ( .A1(n9133), .A2(n9340), .ZN(n8754) );
  NOR2_X1 U15798 ( .A1(n9341), .A2(n8756), .ZN(n8757) );
  XNOR2_X1 U15799 ( .A(n10149), .B(n8757), .ZN(n9842) );
  NAND3_X1 U15800 ( .A1(n9148), .A2(n6747), .A3(n11), .ZN(n8758) );
  MUX2_X1 U15801 ( .A(n8762), .B(n8945), .S(n8941), .Z(n8766) );
  XNOR2_X1 U15802 ( .A(n9710), .B(n10151), .ZN(n10252) );
  XNOR2_X1 U15803 ( .A(n10252), .B(n9842), .ZN(n8775) );
  XNOR2_X1 U15805 ( .A(n9678), .B(n9908), .ZN(n8773) );
  INV_X1 U15806 ( .A(n1123), .ZN(n26656) );
  XNOR2_X1 U15808 ( .A(n8773), .B(n8772), .ZN(n8774) );
  INV_X1 U15809 ( .A(n11337), .ZN(n11174) );
  NOR2_X1 U15810 ( .A1(n8995), .A2(n9210), .ZN(n8776) );
  XNOR2_X1 U15814 ( .A(n9446), .B(n10218), .ZN(n9836) );
  NAND2_X1 U15815 ( .A1(n9188), .A2(n8782), .ZN(n9006) );
  NAND3_X1 U15816 ( .A1(n9187), .A2(n9009), .A3(n9007), .ZN(n8783) );
  XNOR2_X1 U15817 ( .A(n9992), .B(n9716), .ZN(n9310) );
  XNOR2_X1 U15818 ( .A(n9310), .B(n9836), .ZN(n8799) );
  OAI211_X1 U15819 ( .C1(n8788), .C2(n8787), .A(n8786), .B(n8785), .ZN(n8789)
         );
  XNOR2_X1 U15820 ( .A(n9626), .B(n9934), .ZN(n8797) );
  INV_X1 U15821 ( .A(n2353), .ZN(n25378) );
  XNOR2_X1 U15822 ( .A(n301), .B(n25378), .ZN(n8796) );
  XNOR2_X1 U15823 ( .A(n8797), .B(n8796), .ZN(n8798) );
  XNOR2_X1 U15824 ( .A(n8799), .B(n8798), .ZN(n10830) );
  AND2_X1 U15825 ( .A1(n8957), .A2(n8803), .ZN(n8807) );
  MUX2_X1 U15826 ( .A(n8805), .B(n8804), .S(n8958), .Z(n8806) );
  OAI21_X2 U15827 ( .B1(n8807), .B2(n29096), .A(n8806), .ZN(n10275) );
  XNOR2_X1 U15829 ( .A(n9852), .B(n10275), .ZN(n9591) );
  INV_X1 U15830 ( .A(n8818), .ZN(n8820) );
  NAND2_X1 U15831 ( .A1(n8820), .A2(n8819), .ZN(n8821) );
  NAND3_X1 U15832 ( .A1(n1839), .A2(n8826), .A3(n8825), .ZN(n8833) );
  NAND3_X1 U15833 ( .A1(n8830), .A2(n8829), .A3(n8828), .ZN(n8831) );
  XNOR2_X1 U15834 ( .A(n9591), .B(n8835), .ZN(n8845) );
  NOR2_X1 U15835 ( .A1(n8837), .A2(n8836), .ZN(n8840) );
  NOR2_X1 U15836 ( .A1(n8966), .A2(n8838), .ZN(n8839) );
  NAND3_X1 U15837 ( .A1(n8964), .A2(n605), .A3(n9170), .ZN(n8841) );
  INV_X1 U15838 ( .A(n2889), .ZN(n27778) );
  XNOR2_X1 U15839 ( .A(n10436), .B(n27778), .ZN(n8843) );
  INV_X1 U15840 ( .A(n8847), .ZN(n11702) );
  NAND2_X1 U15841 ( .A1(n11702), .A2(n12202), .ZN(n9058) );
  OAI21_X1 U15842 ( .B1(n28500), .B2(n8848), .A(n2320), .ZN(n8849) );
  NAND3_X1 U15843 ( .A1(n8852), .A2(n29311), .A3(n8851), .ZN(n8853) );
  OAI21_X2 U15846 ( .B1(n8862), .B2(n8861), .A(n8860), .ZN(n10385) );
  XNOR2_X1 U15847 ( .A(n10385), .B(n9619), .ZN(n10177) );
  XNOR2_X1 U15848 ( .A(n10321), .B(n2350), .ZN(n8863) );
  NAND3_X1 U15849 ( .A1(n9062), .A2(n8864), .A3(n9064), .ZN(n8870) );
  NAND2_X1 U15850 ( .A1(n9062), .A2(n8865), .ZN(n8867) );
  NAND3_X1 U15851 ( .A1(n8868), .A2(n8867), .A3(n8866), .ZN(n8869) );
  MUX2_X1 U15852 ( .A(n8403), .B(n8876), .S(n8874), .Z(n8882) );
  NAND3_X1 U15853 ( .A1(n8403), .A2(n8876), .A3(n8875), .ZN(n8880) );
  NAND2_X1 U15854 ( .A1(n8878), .A2(n8877), .ZN(n8879) );
  XNOR2_X1 U15855 ( .A(n8884), .B(n8885), .ZN(n10473) );
  INV_X1 U15856 ( .A(n10473), .ZN(n11323) );
  OAI22_X1 U15857 ( .A1(n8888), .A2(n8887), .B1(n8886), .B2(n8890), .ZN(n8895)
         );
  NAND2_X1 U15858 ( .A1(n8890), .A2(n8889), .ZN(n8893) );
  INV_X1 U15859 ( .A(n9824), .ZN(n8896) );
  XNOR2_X1 U15860 ( .A(n10282), .B(n8896), .ZN(n8903) );
  INV_X1 U15861 ( .A(n9125), .ZN(n8897) );
  NAND2_X1 U15862 ( .A1(n8900), .A2(n8899), .ZN(n8901) );
  XNOR2_X1 U15863 ( .A(n8902), .B(n8903), .ZN(n8923) );
  INV_X1 U15864 ( .A(n8904), .ZN(n8921) );
  INV_X1 U15865 ( .A(n9012), .ZN(n8905) );
  AND2_X1 U15866 ( .A1(n8907), .A2(n8906), .ZN(n8913) );
  NAND2_X1 U15867 ( .A1(n8908), .A2(n9012), .ZN(n8909) );
  OAI21_X1 U15868 ( .B1(n608), .B2(n9012), .A(n8909), .ZN(n8911) );
  NAND2_X1 U15869 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  NAND2_X1 U15870 ( .A1(n8913), .A2(n8912), .ZN(n10411) );
  NAND2_X1 U15871 ( .A1(n8916), .A2(n8915), .ZN(n8919) );
  AND2_X1 U15872 ( .A1(n8917), .A2(n9107), .ZN(n8918) );
  XNOR2_X1 U15873 ( .A(n10411), .B(n9647), .ZN(n9903) );
  XNOR2_X1 U15874 ( .A(n8921), .B(n9903), .ZN(n8922) );
  NAND2_X1 U15876 ( .A1(n11323), .A2(n10810), .ZN(n10859) );
  OAI21_X1 U15877 ( .B1(n9133), .B2(n9134), .A(n8924), .ZN(n8927) );
  XNOR2_X1 U15879 ( .A(n10202), .B(n3650), .ZN(n8928) );
  XNOR2_X1 U15880 ( .A(n9779), .B(n8928), .ZN(n8940) );
  NAND2_X1 U15881 ( .A1(n6747), .A2(n8929), .ZN(n9147) );
  NAND2_X1 U15882 ( .A1(n8931), .A2(n9148), .ZN(n8934) );
  NAND2_X1 U15883 ( .A1(n9374), .A2(n5958), .ZN(n8932) );
  AOI21_X2 U15884 ( .B1(n8935), .B2(n8934), .A(n8933), .ZN(n10396) );
  XNOR2_X1 U15885 ( .A(n10396), .B(n1868), .ZN(n9523) );
  XNOR2_X1 U15886 ( .A(n9996), .B(n10289), .ZN(n8951) );
  NOR2_X1 U15887 ( .A1(n8941), .A2(n9561), .ZN(n8942) );
  AOI21_X1 U15888 ( .B1(n8947), .B2(n8943), .A(n8942), .ZN(n8949) );
  NAND2_X1 U15889 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  NOR2_X1 U15890 ( .A1(n8947), .A2(n8946), .ZN(n8948) );
  INV_X1 U15891 ( .A(n10371), .ZN(n8950) );
  XNOR2_X1 U15892 ( .A(n8951), .B(n8950), .ZN(n8952) );
  INV_X1 U15893 ( .A(n10472), .ZN(n11184) );
  INV_X1 U15894 ( .A(n8953), .ZN(n8972) );
  MUX2_X1 U15895 ( .A(n8956), .B(n8955), .S(n29096), .Z(n8960) );
  NOR2_X1 U15896 ( .A1(n8962), .A2(n8961), .ZN(n8971) );
  OAI21_X1 U15897 ( .B1(n8964), .B2(n8963), .A(n605), .ZN(n8970) );
  OAI21_X1 U15898 ( .B1(n605), .B2(n8966), .A(n8965), .ZN(n8969) );
  INV_X1 U15899 ( .A(n8967), .ZN(n8968) );
  INV_X1 U15900 ( .A(n9540), .ZN(n10419) );
  XNOR2_X1 U15901 ( .A(n10419), .B(n9613), .ZN(n9872) );
  XNOR2_X1 U15902 ( .A(n9872), .B(n8972), .ZN(n8991) );
  XNOR2_X1 U15903 ( .A(n10294), .B(n2982), .ZN(n8989) );
  INV_X1 U15904 ( .A(n8973), .ZN(n8975) );
  NAND2_X1 U15905 ( .A1(n607), .A2(n8978), .ZN(n8979) );
  NAND3_X1 U15906 ( .A1(n8982), .A2(n8981), .A3(n8980), .ZN(n8986) );
  INV_X1 U15908 ( .A(n10258), .ZN(n9528) );
  XNOR2_X1 U15909 ( .A(n9528), .B(n10345), .ZN(n9833) );
  XNOR2_X1 U15910 ( .A(n8989), .B(n9833), .ZN(n8990) );
  NAND3_X1 U15911 ( .A1(n10859), .A2(n8992), .A3(n11322), .ZN(n9056) );
  NAND3_X1 U15912 ( .A1(n9434), .A2(n8996), .A3(n4305), .ZN(n8997) );
  NAND2_X1 U15913 ( .A1(n9196), .A2(n9206), .ZN(n8999) );
  AND2_X1 U15914 ( .A1(n8999), .A2(n9197), .ZN(n9002) );
  XNOR2_X1 U15915 ( .A(n10189), .B(n9003), .ZN(n9022) );
  NAND2_X1 U15916 ( .A1(n9009), .A2(n9007), .ZN(n9005) );
  AOI21_X1 U15917 ( .B1(n9006), .B2(n9005), .A(n9004), .ZN(n9011) );
  NAND2_X1 U15918 ( .A1(n9184), .A2(n9007), .ZN(n9008) );
  AOI21_X1 U15919 ( .B1(n9009), .B2(n9008), .A(n9188), .ZN(n9010) );
  NAND3_X1 U15920 ( .A1(n9013), .A2(n9012), .A3(n9014), .ZN(n9017) );
  XNOR2_X1 U15921 ( .A(n9512), .B(n10362), .ZN(n9820) );
  XNOR2_X1 U15922 ( .A(n10304), .B(n2598), .ZN(n9020) );
  XNOR2_X1 U15923 ( .A(n9820), .B(n9020), .ZN(n9021) );
  NAND2_X1 U15924 ( .A1(n9222), .A2(n9220), .ZN(n9023) );
  NAND2_X1 U15925 ( .A1(n597), .A2(n9023), .ZN(n9025) );
  NOR2_X1 U15927 ( .A1(n9035), .A2(n9034), .ZN(n9036) );
  NAND2_X1 U15928 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  NOR2_X1 U15929 ( .A1(n9039), .A2(n8109), .ZN(n9040) );
  INV_X1 U15931 ( .A(n9849), .ZN(n9044) );
  XNOR2_X1 U15932 ( .A(n9044), .B(n9631), .ZN(n9053) );
  XNOR2_X1 U15933 ( .A(n9592), .B(n10071), .ZN(n9051) );
  XNOR2_X1 U15934 ( .A(n10435), .B(n3321), .ZN(n9050) );
  XNOR2_X1 U15935 ( .A(n9051), .B(n9050), .ZN(n9052) );
  NAND3_X1 U15936 ( .A1(n11187), .A2(n11181), .A3(n11321), .ZN(n9054) );
  NAND2_X1 U15937 ( .A1(n12205), .A2(n12200), .ZN(n9057) );
  MUX2_X1 U15939 ( .A(n9059), .B(n9060), .S(n9062), .Z(n9065) );
  XNOR2_X1 U15940 ( .A(n10258), .B(n2509), .ZN(n9066) );
  XNOR2_X1 U15941 ( .A(n9066), .B(n1891), .ZN(n9068) );
  XNOR2_X1 U15942 ( .A(n10297), .B(n1902), .ZN(n9067) );
  XNOR2_X1 U15943 ( .A(n9068), .B(n9067), .ZN(n9093) );
  OAI21_X1 U15944 ( .B1(n9071), .B2(n9070), .A(n9069), .ZN(n9077) );
  OAI21_X1 U15945 ( .B1(n9074), .B2(n9073), .A(n9072), .ZN(n9076) );
  OAI21_X1 U15946 ( .B1(n9079), .B2(n28500), .A(n9078), .ZN(n9091) );
  NAND2_X1 U15947 ( .A1(n28500), .A2(n29310), .ZN(n9089) );
  INV_X1 U15948 ( .A(n9082), .ZN(n9086) );
  INV_X1 U15949 ( .A(n9083), .ZN(n9085) );
  OAI21_X1 U15950 ( .B1(n9086), .B2(n9085), .A(n9084), .ZN(n9087) );
  NAND2_X1 U15951 ( .A1(n9089), .A2(n9088), .ZN(n9090) );
  XNOR2_X1 U15952 ( .A(n9695), .B(n10344), .ZN(n10057) );
  XNOR2_X1 U15953 ( .A(n1920), .B(n10057), .ZN(n9092) );
  INV_X1 U15954 ( .A(n9094), .ZN(n9462) );
  OAI21_X1 U15955 ( .B1(n9097), .B2(n9096), .A(n9095), .ZN(n9103) );
  INV_X1 U15956 ( .A(n9098), .ZN(n9101) );
  OAI21_X1 U15957 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9102) );
  NAND2_X1 U15958 ( .A1(n9103), .A2(n9102), .ZN(n10363) );
  INV_X1 U15959 ( .A(n9107), .ZN(n9104) );
  NAND3_X1 U15960 ( .A1(n9108), .A2(n9118), .A3(n9107), .ZN(n9120) );
  INV_X1 U15961 ( .A(n9109), .ZN(n9111) );
  NAND2_X1 U15962 ( .A1(n9111), .A2(n28810), .ZN(n9117) );
  INV_X1 U15963 ( .A(n9112), .ZN(n9114) );
  NAND2_X1 U15964 ( .A1(n9114), .A2(n29135), .ZN(n9115) );
  NAND4_X1 U15965 ( .A1(n9118), .A2(n9117), .A3(n9116), .A4(n9115), .ZN(n9119)
         );
  XNOR2_X1 U15966 ( .A(n9462), .B(n10086), .ZN(n9130) );
  AOI22_X1 U15967 ( .A1(n9125), .A2(n9124), .B1(n29304), .B2(n9122), .ZN(n9126) );
  INV_X1 U15968 ( .A(n9512), .ZN(n9881) );
  XNOR2_X1 U15969 ( .A(n9794), .B(n9881), .ZN(n9128) );
  XNOR2_X1 U15970 ( .A(n9964), .B(n3232), .ZN(n9127) );
  XNOR2_X1 U15971 ( .A(n9128), .B(n9127), .ZN(n9129) );
  AND2_X1 U15972 ( .A1(n9132), .A2(n9133), .ZN(n9135) );
  XNOR2_X1 U15973 ( .A(n1877), .B(n10283), .ZN(n9138) );
  XNOR2_X1 U15974 ( .A(n10332), .B(n9138), .ZN(n9159) );
  OAI21_X1 U15975 ( .B1(n598), .B2(n9142), .A(n9141), .ZN(n9143) );
  XNOR2_X1 U15976 ( .A(n10159), .B(n9824), .ZN(n9157) );
  INV_X1 U15977 ( .A(n9147), .ZN(n9154) );
  AOI21_X1 U15978 ( .B1(n6747), .B2(n9149), .A(n9148), .ZN(n9151) );
  NAND2_X1 U15979 ( .A1(n9152), .A2(n9151), .ZN(n9153) );
  XNOR2_X1 U15980 ( .A(n1918), .B(n27452), .ZN(n9156) );
  XNOR2_X1 U15981 ( .A(n9157), .B(n9156), .ZN(n9158) );
  OAI21_X1 U15982 ( .B1(n9161), .B2(n9160), .A(n9164), .ZN(n9168) );
  INV_X1 U15983 ( .A(n9162), .ZN(n9166) );
  NAND2_X1 U15984 ( .A1(n9164), .A2(n9163), .ZN(n9165) );
  INV_X1 U15985 ( .A(n9357), .ZN(n9175) );
  XNOR2_X1 U15986 ( .A(n9175), .B(n10373), .ZN(n9182) );
  INV_X1 U15987 ( .A(n9176), .ZN(n9178) );
  XNOR2_X1 U15988 ( .A(n9684), .B(n10395), .ZN(n9450) );
  XNOR2_X1 U15989 ( .A(n1868), .B(n3035), .ZN(n9180) );
  XNOR2_X1 U15990 ( .A(n9450), .B(n9180), .ZN(n9181) );
  NAND2_X1 U15991 ( .A1(n10847), .A2(n11347), .ZN(n9219) );
  XNOR2_X1 U15992 ( .A(n9504), .B(n26909), .ZN(n9183) );
  XNOR2_X1 U15993 ( .A(n9183), .B(n10271), .ZN(n9193) );
  MUX2_X1 U15994 ( .A(n9188), .B(n9187), .S(n9184), .Z(n9192) );
  XNOR2_X1 U15997 ( .A(n10072), .B(n10353), .ZN(n9811) );
  XNOR2_X1 U15998 ( .A(n9811), .B(n9193), .ZN(n9217) );
  NAND2_X1 U15999 ( .A1(n9195), .A2(n9194), .ZN(n9205) );
  NOR2_X1 U16000 ( .A1(n9196), .A2(n9200), .ZN(n9198) );
  OAI21_X1 U16001 ( .B1(n9199), .B2(n9198), .A(n9197), .ZN(n9204) );
  NAND3_X1 U16002 ( .A1(n9202), .A2(n9201), .A3(n9200), .ZN(n9203) );
  OAI211_X1 U16003 ( .C1(n9206), .C2(n9205), .A(n9204), .B(n9203), .ZN(n9629)
         );
  INV_X1 U16004 ( .A(n9207), .ZN(n9215) );
  OAI21_X1 U16005 ( .B1(n9209), .B2(n4305), .A(n9208), .ZN(n9214) );
  NAND3_X1 U16006 ( .A1(n9211), .A2(n9210), .A3(n4305), .ZN(n9213) );
  NAND3_X1 U16007 ( .A1(n9434), .A2(n9436), .A3(n9438), .ZN(n9212) );
  XNOR2_X1 U16009 ( .A(n10356), .B(n9629), .ZN(n10432) );
  XNOR2_X1 U16010 ( .A(n10432), .B(n10359), .ZN(n9216) );
  INV_X1 U16012 ( .A(n11349), .ZN(n9218) );
  NAND3_X1 U16013 ( .A1(n9224), .A2(n9223), .A3(n9228), .ZN(n9225) );
  NOR2_X1 U16014 ( .A1(n9229), .A2(n9233), .ZN(n9231) );
  INV_X1 U16015 ( .A(n9232), .ZN(n9234) );
  OAI21_X1 U16016 ( .B1(n9238), .B2(n9237), .A(n9236), .ZN(n9239) );
  XNOR2_X1 U16018 ( .A(n10251), .B(n10384), .ZN(n9241) );
  NAND2_X1 U16019 ( .A1(n9246), .A2(n9245), .ZN(n9250) );
  XNOR2_X1 U16020 ( .A(n9677), .B(n9976), .ZN(n9253) );
  XNOR2_X1 U16021 ( .A(n9550), .B(n3625), .ZN(n9252) );
  XNOR2_X1 U16022 ( .A(n9253), .B(n9252), .ZN(n9254) );
  NAND2_X1 U16023 ( .A1(n10476), .A2(n11347), .ZN(n10477) );
  AOI21_X1 U16024 ( .B1(n10477), .B2(n10847), .A(n11192), .ZN(n9256) );
  MUX2_X2 U16025 ( .A(n9259), .B(n9258), .S(n5825), .Z(n12738) );
  XNOR2_X1 U16026 ( .A(n12738), .B(n3015), .ZN(n9478) );
  XNOR2_X1 U16027 ( .A(n9763), .B(n9629), .ZN(n9260) );
  XNOR2_X1 U16028 ( .A(n9849), .B(n9260), .ZN(n9264) );
  XNOR2_X1 U16029 ( .A(n9509), .B(n9852), .ZN(n10127) );
  INV_X1 U16030 ( .A(n10127), .ZN(n9262) );
  XNOR2_X1 U16031 ( .A(n10071), .B(n3722), .ZN(n9261) );
  XNOR2_X1 U16032 ( .A(n9262), .B(n9261), .ZN(n9263) );
  INV_X1 U16034 ( .A(n9820), .ZN(n9265) );
  XNOR2_X1 U16035 ( .A(n9929), .B(n9877), .ZN(n10119) );
  XNOR2_X1 U16036 ( .A(n9265), .B(n10119), .ZN(n9270) );
  XNOR2_X1 U16037 ( .A(n9930), .B(n1923), .ZN(n9267) );
  XNOR2_X1 U16038 ( .A(n9268), .B(n9267), .ZN(n9269) );
  INV_X1 U16040 ( .A(n10941), .ZN(n10110) );
  XNOR2_X1 U16041 ( .A(n10371), .B(n10391), .ZN(n10079) );
  XNOR2_X1 U16042 ( .A(n9755), .B(n9894), .ZN(n10220) );
  XNOR2_X1 U16043 ( .A(n10145), .B(n3196), .ZN(n9271) );
  XNOR2_X1 U16044 ( .A(n10220), .B(n9271), .ZN(n9272) );
  INV_X1 U16045 ( .A(n10940), .ZN(n10446) );
  XNOR2_X1 U16046 ( .A(n9824), .B(n9948), .ZN(n9520) );
  XNOR2_X1 U16047 ( .A(n10328), .B(n10412), .ZN(n10065) );
  INV_X1 U16048 ( .A(n10065), .ZN(n9646) );
  XNOR2_X1 U16049 ( .A(n9646), .B(n9520), .ZN(n9276) );
  XNOR2_X1 U16050 ( .A(n9749), .B(n9899), .ZN(n9274) );
  XNOR2_X1 U16051 ( .A(n10160), .B(n27956), .ZN(n9273) );
  XNOR2_X1 U16052 ( .A(n9274), .B(n9273), .ZN(n9275) );
  NAND2_X1 U16053 ( .A1(n10446), .A2(n10703), .ZN(n9281) );
  XNOR2_X1 U16054 ( .A(n9918), .B(n9833), .ZN(n9280) );
  XNOR2_X1 U16055 ( .A(n9695), .B(n10133), .ZN(n9278) );
  XNOR2_X1 U16056 ( .A(n9799), .B(n3369), .ZN(n9277) );
  XNOR2_X1 U16057 ( .A(n9278), .B(n9277), .ZN(n9279) );
  XNOR2_X1 U16059 ( .A(n10251), .B(n1884), .ZN(n9283) );
  INV_X1 U16060 ( .A(n9352), .ZN(n9711) );
  XNOR2_X1 U16061 ( .A(n10149), .B(n9711), .ZN(n9282) );
  XNOR2_X1 U16062 ( .A(n9282), .B(n9283), .ZN(n9288) );
  XNOR2_X1 U16063 ( .A(n1852), .B(n27231), .ZN(n9286) );
  XNOR2_X1 U16064 ( .A(n28488), .B(n9771), .ZN(n9285) );
  XNOR2_X1 U16065 ( .A(n9286), .B(n9285), .ZN(n9287) );
  NOR2_X1 U16067 ( .A1(n10705), .A2(n10942), .ZN(n10704) );
  INV_X1 U16068 ( .A(n10704), .ZN(n9290) );
  AOI21_X1 U16069 ( .B1(n10942), .B2(n10110), .A(n10703), .ZN(n9289) );
  NAND2_X1 U16070 ( .A1(n9290), .A2(n9289), .ZN(n9291) );
  XNOR2_X1 U16072 ( .A(n9710), .B(n10335), .ZN(n9293) );
  XNOR2_X1 U16073 ( .A(n10319), .B(n9293), .ZN(n9297) );
  INV_X1 U16074 ( .A(n3164), .ZN(n9294) );
  XNOR2_X1 U16075 ( .A(n10178), .B(n9294), .ZN(n9296) );
  XNOR2_X1 U16076 ( .A(n10356), .B(n2527), .ZN(n9298) );
  XNOR2_X1 U16077 ( .A(n9956), .B(n9298), .ZN(n9300) );
  XNOR2_X1 U16078 ( .A(n9851), .B(n9941), .ZN(n10315) );
  XNOR2_X1 U16079 ( .A(n10315), .B(n9590), .ZN(n9299) );
  XNOR2_X1 U16080 ( .A(n10038), .B(n9971), .ZN(n9302) );
  XNOR2_X1 U16081 ( .A(n10183), .B(n3422), .ZN(n9303) );
  XNOR2_X1 U16082 ( .A(n9303), .B(n10064), .ZN(n9305) );
  XNOR2_X1 U16083 ( .A(n9305), .B(n9304), .ZN(n9308) );
  XNOR2_X1 U16084 ( .A(n9949), .B(n10043), .ZN(n9307) );
  XNOR2_X1 U16086 ( .A(n9307), .B(n9725), .ZN(n10286) );
  XNOR2_X1 U16087 ( .A(n9308), .B(n10286), .ZN(n10973) );
  XNOR2_X1 U16089 ( .A(n9818), .B(n9705), .ZN(n9309) );
  XNOR2_X1 U16090 ( .A(n9311), .B(n9310), .ZN(n9317) );
  XNOR2_X1 U16091 ( .A(n10143), .B(n857), .ZN(n9315) );
  XNOR2_X1 U16092 ( .A(n5412), .B(n9997), .ZN(n9314) );
  XNOR2_X1 U16093 ( .A(n9315), .B(n9314), .ZN(n9316) );
  XNOR2_X1 U16095 ( .A(n10088), .B(n9930), .ZN(n10268) );
  INV_X1 U16096 ( .A(n10268), .ZN(n9319) );
  INV_X1 U16097 ( .A(n10264), .ZN(n9318) );
  XNOR2_X1 U16098 ( .A(n9319), .B(n9962), .ZN(n9322) );
  XNOR2_X1 U16099 ( .A(n9878), .B(n10304), .ZN(n9741) );
  XNOR2_X1 U16100 ( .A(n10426), .B(n1161), .ZN(n9320) );
  XNOR2_X1 U16101 ( .A(n9741), .B(n9320), .ZN(n9321) );
  XNOR2_X1 U16102 ( .A(n9322), .B(n9321), .ZN(n9344) );
  INV_X1 U16103 ( .A(n9344), .ZN(n10605) );
  XNOR2_X1 U16104 ( .A(n9735), .B(n9323), .ZN(n10256) );
  INV_X1 U16105 ( .A(n10256), .ZN(n9324) );
  XNOR2_X1 U16106 ( .A(n9324), .B(n9736), .ZN(n9328) );
  XNOR2_X1 U16107 ( .A(n10257), .B(n9971), .ZN(n9326) );
  XNOR2_X1 U16108 ( .A(n10419), .B(n2981), .ZN(n9325) );
  XNOR2_X1 U16109 ( .A(n9325), .B(n9326), .ZN(n9327) );
  NAND2_X1 U16110 ( .A1(n10605), .A2(n10913), .ZN(n10732) );
  INV_X1 U16111 ( .A(n10732), .ZN(n9333) );
  XNOR2_X1 U16112 ( .A(n10128), .B(n9592), .ZN(n9767) );
  XNOR2_X1 U16113 ( .A(n10277), .B(n9767), .ZN(n9332) );
  XNOR2_X1 U16114 ( .A(n10275), .B(n10310), .ZN(n9330) );
  XNOR2_X1 U16115 ( .A(n10435), .B(n3752), .ZN(n9329) );
  XNOR2_X1 U16116 ( .A(n9330), .B(n9329), .ZN(n9331) );
  XNOR2_X1 U16117 ( .A(n9332), .B(n9331), .ZN(n10735) );
  INV_X1 U16118 ( .A(n10735), .ZN(n10914) );
  NAND2_X1 U16119 ( .A1(n9333), .A2(n10914), .ZN(n11526) );
  XNOR2_X1 U16120 ( .A(n9997), .B(n9755), .ZN(n9335) );
  XNOR2_X1 U16121 ( .A(n10289), .B(n2274), .ZN(n9334) );
  XNOR2_X1 U16122 ( .A(n9335), .B(n9334), .ZN(n9338) );
  XNOR2_X1 U16123 ( .A(n10396), .B(n10218), .ZN(n9780) );
  INV_X1 U16124 ( .A(n10912), .ZN(n10689) );
  XNOR2_X1 U16125 ( .A(n10322), .B(n28693), .ZN(n9339) );
  XNOR2_X1 U16126 ( .A(n9771), .B(n9979), .ZN(n9342) );
  XNOR2_X1 U16127 ( .A(n9342), .B(n10060), .ZN(n10253) );
  XNOR2_X2 U16128 ( .A(n9343), .B(n10253), .ZN(n10911) );
  NAND2_X1 U16129 ( .A1(n10689), .A2(n10911), .ZN(n10733) );
  INV_X1 U16130 ( .A(n10913), .ZN(n10609) );
  OAI211_X1 U16131 ( .C1(n10605), .C2(n10689), .A(n10733), .B(n10609), .ZN(
        n11525) );
  XNOR2_X1 U16132 ( .A(n9749), .B(n9823), .ZN(n9491) );
  XNOR2_X1 U16133 ( .A(n9748), .B(n9491), .ZN(n9347) );
  XNOR2_X1 U16134 ( .A(n10411), .B(n3451), .ZN(n9345) );
  XNOR2_X1 U16135 ( .A(n9306), .B(n10227), .ZN(n9984) );
  XNOR2_X1 U16136 ( .A(n9345), .B(n9984), .ZN(n9346) );
  NAND3_X1 U16137 ( .A1(n10911), .A2(n10916), .A3(n9348), .ZN(n11523) );
  NAND2_X1 U16138 ( .A1(n13087), .A2(n11982), .ZN(n9349) );
  OAI21_X1 U16139 ( .B1(n11810), .B2(n13087), .A(n9349), .ZN(n9477) );
  XNOR2_X1 U16140 ( .A(n1917), .B(n1247), .ZN(n9350) );
  XNOR2_X1 U16141 ( .A(n9986), .B(n9948), .ZN(n9351) );
  XNOR2_X1 U16142 ( .A(n9647), .B(n9517), .ZN(n10188) );
  XNOR2_X1 U16143 ( .A(n10019), .B(n9352), .ZN(n10383) );
  INV_X1 U16144 ( .A(n10383), .ZN(n9620) );
  XNOR2_X1 U16145 ( .A(n10250), .B(n28488), .ZN(n9353) );
  XNOR2_X1 U16146 ( .A(n9620), .B(n9353), .ZN(n9356) );
  INV_X1 U16147 ( .A(n2973), .ZN(n24959) );
  XNOR2_X1 U16148 ( .A(n9619), .B(n24959), .ZN(n9354) );
  XNOR2_X1 U16149 ( .A(n10179), .B(n9354), .ZN(n9355) );
  XNOR2_X1 U16150 ( .A(n9356), .B(n9355), .ZN(n9863) );
  INV_X1 U16151 ( .A(n9863), .ZN(n9362) );
  XNOR2_X1 U16152 ( .A(n10372), .B(n9717), .ZN(n10027) );
  XNOR2_X1 U16153 ( .A(n9357), .B(n10027), .ZN(n9361) );
  XNOR2_X1 U16154 ( .A(n9996), .B(n28634), .ZN(n9359) );
  XNOR2_X1 U16155 ( .A(n10202), .B(n3015), .ZN(n9358) );
  XNOR2_X1 U16156 ( .A(n9358), .B(n9359), .ZN(n9360) );
  NAND2_X1 U16157 ( .A1(n9362), .A2(n10962), .ZN(n10602) );
  OAI21_X1 U16158 ( .B1(n10958), .B2(n28173), .A(n10602), .ZN(n9391) );
  XNOR2_X1 U16160 ( .A(n9368), .B(n10352), .ZN(n9369) );
  XNOR2_X1 U16161 ( .A(n9631), .B(n9369), .ZN(n9382) );
  INV_X1 U16162 ( .A(n9370), .ZN(n9372) );
  NAND2_X1 U16163 ( .A1(n9372), .A2(n11), .ZN(n9377) );
  INV_X1 U16164 ( .A(n9373), .ZN(n9375) );
  NAND2_X1 U16165 ( .A1(n9375), .A2(n9374), .ZN(n9376) );
  NAND3_X1 U16166 ( .A1(n9378), .A2(n9377), .A3(n9376), .ZN(n9379) );
  XNOR2_X1 U16167 ( .A(n9504), .B(n1911), .ZN(n9380) );
  XNOR2_X1 U16168 ( .A(n9721), .B(n9380), .ZN(n9381) );
  XNOR2_X1 U16169 ( .A(n9382), .B(n9381), .ZN(n10956) );
  INV_X1 U16170 ( .A(n9695), .ZN(n9383) );
  XNOR2_X1 U16171 ( .A(n10138), .B(n27462), .ZN(n9384) );
  XNOR2_X1 U16172 ( .A(n10169), .B(n9384), .ZN(n9385) );
  XNOR2_X1 U16173 ( .A(n9386), .B(n9385), .ZN(n10963) );
  XNOR2_X1 U16174 ( .A(n10191), .B(n10263), .ZN(n10005) );
  XNOR2_X1 U16175 ( .A(n10005), .B(n10424), .ZN(n9389) );
  XNOR2_X1 U16176 ( .A(n9639), .B(n9929), .ZN(n9388) );
  XNOR2_X1 U16177 ( .A(n10193), .B(n2446), .ZN(n9387) );
  OAI21_X1 U16178 ( .B1(n9858), .B2(n10780), .A(n10687), .ZN(n9390) );
  AOI22_X1 U16179 ( .A1(n9391), .A2(n9390), .B1(n28173), .B2(n9858), .ZN(
        n12226) );
  XNOR2_X1 U16180 ( .A(n10298), .B(n10134), .ZN(n9969) );
  XNOR2_X1 U16181 ( .A(n9732), .B(n9613), .ZN(n9453) );
  XNOR2_X1 U16182 ( .A(n9969), .B(n9453), .ZN(n9395) );
  XNOR2_X1 U16183 ( .A(n10344), .B(n9392), .ZN(n10418) );
  XNOR2_X1 U16184 ( .A(n1920), .B(n3378), .ZN(n9393) );
  XNOR2_X1 U16185 ( .A(n10418), .B(n9393), .ZN(n9394) );
  OAI22_X1 U16186 ( .A1(n436), .A2(n9398), .B1(n9397), .B2(n609), .ZN(n9400)
         );
  NOR2_X1 U16187 ( .A1(n9400), .A2(n9399), .ZN(n9401) );
  XNOR2_X1 U16188 ( .A(n9961), .B(n10425), .ZN(n9405) );
  XNOR2_X1 U16189 ( .A(n9964), .B(n1887), .ZN(n9402) );
  XNOR2_X1 U16190 ( .A(n9403), .B(n9402), .ZN(n9404) );
  XNOR2_X1 U16191 ( .A(n9985), .B(n10332), .ZN(n9408) );
  XNOR2_X1 U16192 ( .A(n9647), .B(n3483), .ZN(n9406) );
  XNOR2_X1 U16193 ( .A(n9687), .B(n9406), .ZN(n9407) );
  INV_X1 U16194 ( .A(n9409), .ZN(n9413) );
  OAI22_X1 U16195 ( .A1(n9413), .A2(n9412), .B1(n28211), .B2(n9410), .ZN(n9415) );
  XNOR2_X1 U16196 ( .A(n10202), .B(n3256), .ZN(n9416) );
  OAI21_X1 U16197 ( .B1(n11004), .B2(n6779), .A(n9417), .ZN(n9694) );
  OAI21_X1 U16198 ( .B1(n10997), .B2(n6779), .A(n9694), .ZN(n11528) );
  XNOR2_X1 U16199 ( .A(n10208), .B(n10356), .ZN(n9418) );
  XNOR2_X1 U16200 ( .A(n10272), .B(n10434), .ZN(n9958) );
  XNOR2_X1 U16201 ( .A(n9418), .B(n9958), .ZN(n9429) );
  INV_X1 U16202 ( .A(n9419), .ZN(n9424) );
  INV_X1 U16203 ( .A(n9420), .ZN(n9423) );
  OAI211_X1 U16204 ( .C1(n9425), .C2(n9424), .A(n9423), .B(n9422), .ZN(n9426)
         );
  XNOR2_X1 U16205 ( .A(n10436), .B(n3686), .ZN(n9427) );
  XNOR2_X1 U16206 ( .A(n9722), .B(n9427), .ZN(n9428) );
  XNOR2_X1 U16207 ( .A(n9428), .B(n9429), .ZN(n11000) );
  XNOR2_X1 U16208 ( .A(n9772), .B(n9430), .ZN(n10337) );
  INV_X1 U16209 ( .A(n10337), .ZN(n9712) );
  XNOR2_X1 U16210 ( .A(n10151), .B(n10386), .ZN(n9981) );
  XNOR2_X1 U16211 ( .A(n9712), .B(n9981), .ZN(n9432) );
  XNOR2_X1 U16212 ( .A(n9431), .B(n10335), .ZN(n10382) );
  OAI211_X1 U16213 ( .C1(n5573), .C2(n592), .A(n10936), .B(n10999), .ZN(n11524) );
  NAND2_X1 U16214 ( .A1(n11528), .A2(n11524), .ZN(n11980) );
  NAND2_X1 U16215 ( .A1(n9433), .A2(n12227), .ZN(n13082) );
  INV_X1 U16218 ( .A(n10045), .ZN(n9440) );
  XNOR2_X1 U16219 ( .A(n10283), .B(n9440), .ZN(n9442) );
  XNOR2_X1 U16220 ( .A(n9899), .B(n3219), .ZN(n9441) );
  XNOR2_X1 U16221 ( .A(n9442), .B(n9441), .ZN(n9445) );
  XNOR2_X1 U16222 ( .A(n10159), .B(n9746), .ZN(n9443) );
  XNOR2_X1 U16223 ( .A(n9443), .B(n10188), .ZN(n9444) );
  INV_X1 U16224 ( .A(n1879), .ZN(n10458) );
  XNOR2_X1 U16225 ( .A(n9446), .B(n10202), .ZN(n9893) );
  INV_X1 U16226 ( .A(n9893), .ZN(n9448) );
  XNOR2_X1 U16227 ( .A(n9447), .B(n10028), .ZN(n10199) );
  XNOR2_X1 U16228 ( .A(n10199), .B(n9448), .ZN(n9452) );
  XNOR2_X1 U16229 ( .A(n9754), .B(n2411), .ZN(n9449) );
  XNOR2_X1 U16230 ( .A(n9450), .B(n9449), .ZN(n9451) );
  XNOR2_X1 U16231 ( .A(n9452), .B(n9451), .ZN(n10924) );
  INV_X1 U16232 ( .A(n10924), .ZN(n9475) );
  NAND2_X1 U16233 ( .A1(n10458), .A2(n9475), .ZN(n10108) );
  INV_X1 U16234 ( .A(n9453), .ZN(n9455) );
  XNOR2_X1 U16235 ( .A(n10133), .B(n1892), .ZN(n9454) );
  XNOR2_X1 U16236 ( .A(n9455), .B(n9454), .ZN(n9459) );
  XNOR2_X1 U16237 ( .A(n10033), .B(n10297), .ZN(n9457) );
  XNOR2_X1 U16238 ( .A(n1902), .B(n25992), .ZN(n9456) );
  XNOR2_X1 U16239 ( .A(n9457), .B(n9456), .ZN(n9458) );
  XNOR2_X1 U16240 ( .A(n9639), .B(n9877), .ZN(n9461) );
  XNOR2_X1 U16241 ( .A(n10009), .B(n891), .ZN(n9460) );
  XNOR2_X1 U16242 ( .A(n9461), .B(n9460), .ZN(n9464) );
  XNOR2_X1 U16243 ( .A(n9462), .B(n9658), .ZN(n9463) );
  XNOR2_X1 U16246 ( .A(n9852), .B(n10208), .ZN(n9887) );
  XNOR2_X1 U16247 ( .A(n10357), .B(n9504), .ZN(n9466) );
  XNOR2_X1 U16248 ( .A(n10073), .B(n3633), .ZN(n9465) );
  XNOR2_X1 U16249 ( .A(n9772), .B(n10384), .ZN(n9470) );
  INV_X1 U16252 ( .A(n9906), .ZN(n9469) );
  XNOR2_X1 U16253 ( .A(n9469), .B(n9470), .ZN(n9474) );
  XNOR2_X1 U16254 ( .A(n9677), .B(n10059), .ZN(n9472) );
  XNOR2_X1 U16255 ( .A(n9550), .B(n5490), .ZN(n9471) );
  XNOR2_X1 U16256 ( .A(n9472), .B(n9471), .ZN(n9473) );
  AOI21_X1 U16257 ( .B1(n10459), .B2(n10458), .A(n590), .ZN(n9476) );
  XNOR2_X1 U16258 ( .A(n9478), .B(n13051), .ZN(n9869) );
  INV_X1 U16259 ( .A(n9771), .ZN(n9479) );
  XNOR2_X1 U16260 ( .A(n9479), .B(n10060), .ZN(n9480) );
  XNOR2_X1 U16261 ( .A(n9981), .B(n9480), .ZN(n9483) );
  XNOR2_X1 U16262 ( .A(n10021), .B(n3751), .ZN(n9481) );
  XNOR2_X1 U16263 ( .A(n10338), .B(n9481), .ZN(n9482) );
  XNOR2_X1 U16264 ( .A(n9851), .B(n10352), .ZN(n10018) );
  XNOR2_X1 U16265 ( .A(n10277), .B(n10018), .ZN(n9486) );
  XNOR2_X1 U16266 ( .A(n9958), .B(n9484), .ZN(n9485) );
  INV_X1 U16267 ( .A(n11318), .ZN(n11254) );
  XNOR2_X1 U16268 ( .A(n9969), .B(n10256), .ZN(n9490) );
  XNOR2_X1 U16269 ( .A(n28643), .B(n10038), .ZN(n9488) );
  XNOR2_X1 U16270 ( .A(n9698), .B(n2385), .ZN(n9487) );
  XNOR2_X1 U16271 ( .A(n9488), .B(n9487), .ZN(n9489) );
  XNOR2_X1 U16272 ( .A(n10043), .B(n27225), .ZN(n9492) );
  XNOR2_X1 U16273 ( .A(n10201), .B(n10392), .ZN(n9494) );
  INV_X1 U16274 ( .A(n3462), .ZN(n27656) );
  XNOR2_X1 U16275 ( .A(n301), .B(n27656), .ZN(n9493) );
  XNOR2_X1 U16276 ( .A(n9494), .B(n9493), .ZN(n9497) );
  XNOR2_X1 U16277 ( .A(n10029), .B(n10219), .ZN(n9838) );
  XNOR2_X1 U16278 ( .A(n9992), .B(n9755), .ZN(n9495) );
  XNOR2_X1 U16279 ( .A(n10191), .B(n9963), .ZN(n10367) );
  INV_X1 U16280 ( .A(n9743), .ZN(n9498) );
  XNOR2_X1 U16281 ( .A(n9498), .B(n10367), .ZN(n9501) );
  XNOR2_X1 U16282 ( .A(n10088), .B(n2402), .ZN(n9499) );
  XNOR2_X1 U16283 ( .A(n9961), .B(n9499), .ZN(n9500) );
  XNOR2_X1 U16284 ( .A(n9501), .B(n9500), .ZN(n10482) );
  MUX2_X2 U16285 ( .A(n9503), .B(n9502), .S(n4296), .Z(n12211) );
  XNOR2_X1 U16286 ( .A(n9505), .B(n9504), .ZN(n9506) );
  XNOR2_X1 U16287 ( .A(n9506), .B(n10271), .ZN(n9508) );
  XNOR2_X1 U16288 ( .A(n10128), .B(n3482), .ZN(n9507) );
  XNOR2_X1 U16289 ( .A(n9508), .B(n9507), .ZN(n9510) );
  XNOR2_X1 U16290 ( .A(n10435), .B(n10073), .ZN(n10212) );
  XNOR2_X1 U16291 ( .A(n10212), .B(n9509), .ZN(n9812) );
  XNOR2_X1 U16292 ( .A(n10193), .B(n1119), .ZN(n9511) );
  XNOR2_X1 U16293 ( .A(n9511), .B(n9878), .ZN(n9513) );
  XNOR2_X1 U16294 ( .A(n9513), .B(n1985), .ZN(n9516) );
  INV_X1 U16295 ( .A(n9929), .ZN(n9514) );
  XNOR2_X1 U16296 ( .A(n9515), .B(n9516), .ZN(n10522) );
  INV_X1 U16297 ( .A(n10522), .ZN(n11274) );
  NAND2_X1 U16298 ( .A1(n11038), .A2(n11274), .ZN(n9548) );
  XNOR2_X1 U16299 ( .A(n9900), .B(n1878), .ZN(n9518) );
  XNOR2_X1 U16300 ( .A(n10232), .B(n3223), .ZN(n9519) );
  XNOR2_X1 U16301 ( .A(n9520), .B(n9519), .ZN(n9521) );
  XNOR2_X1 U16302 ( .A(n9522), .B(n9521), .ZN(n11269) );
  INV_X1 U16303 ( .A(n11269), .ZN(n11034) );
  XNOR2_X1 U16304 ( .A(n9523), .B(n10199), .ZN(n9527) );
  XNOR2_X1 U16305 ( .A(n28634), .B(n10144), .ZN(n9525) );
  XNOR2_X1 U16306 ( .A(n9716), .B(n5633), .ZN(n9524) );
  XNOR2_X1 U16307 ( .A(n9525), .B(n9524), .ZN(n9526) );
  XNOR2_X1 U16308 ( .A(n9527), .B(n9526), .ZN(n11272) );
  NAND2_X1 U16309 ( .A1(n11034), .A2(n28612), .ZN(n9547) );
  XNOR2_X1 U16310 ( .A(n10137), .B(n9528), .ZN(n9873) );
  INV_X1 U16311 ( .A(n9873), .ZN(n9541) );
  OAI21_X1 U16312 ( .B1(n29662), .B2(n9533), .A(n9532), .ZN(n9535) );
  NAND2_X1 U16313 ( .A1(n9536), .A2(n9535), .ZN(n9538) );
  NAND2_X1 U16314 ( .A1(n9538), .A2(n9537), .ZN(n9539) );
  XNOR2_X1 U16315 ( .A(n9540), .B(n9539), .ZN(n10173) );
  XNOR2_X1 U16316 ( .A(n9541), .B(n10173), .ZN(n9546) );
  XNOR2_X1 U16317 ( .A(n9542), .B(n9696), .ZN(n9544) );
  XNOR2_X1 U16318 ( .A(n10138), .B(n2523), .ZN(n9543) );
  XNOR2_X1 U16319 ( .A(n9544), .B(n9543), .ZN(n9545) );
  MUX2_X1 U16320 ( .A(n9548), .B(n9547), .S(n279), .Z(n9557) );
  XNOR2_X1 U16321 ( .A(n9907), .B(n9549), .ZN(n9554) );
  XNOR2_X1 U16322 ( .A(n9710), .B(n10385), .ZN(n9552) );
  XNOR2_X1 U16323 ( .A(n9550), .B(n3660), .ZN(n9551) );
  XNOR2_X1 U16324 ( .A(n9552), .B(n9551), .ZN(n9553) );
  NAND2_X1 U16325 ( .A1(n9555), .A2(n11269), .ZN(n9556) );
  XNOR2_X1 U16326 ( .A(n10386), .B(n2984), .ZN(n9559) );
  INV_X1 U16327 ( .A(n9786), .ZN(n9558) );
  XNOR2_X1 U16328 ( .A(n9559), .B(n9558), .ZN(n9560) );
  XNOR2_X1 U16329 ( .A(n9560), .B(n9842), .ZN(n9571) );
  XNOR2_X1 U16330 ( .A(n10321), .B(n10178), .ZN(n9570) );
  NAND3_X1 U16331 ( .A1(n9566), .A2(n9562), .A3(n9561), .ZN(n9563) );
  OAI211_X1 U16332 ( .C1(n9566), .C2(n9565), .A(n9564), .B(n9563), .ZN(n9568)
         );
  NOR2_X1 U16333 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  XNOR2_X1 U16334 ( .A(n9570), .B(n9569), .ZN(n9926) );
  INV_X1 U16335 ( .A(n9817), .ZN(n9574) );
  XNOR2_X1 U16336 ( .A(n9795), .B(n3635), .ZN(n9572) );
  XNOR2_X1 U16337 ( .A(n9572), .B(n10302), .ZN(n9573) );
  XNOR2_X1 U16338 ( .A(n9574), .B(n9573), .ZN(n9578) );
  XNOR2_X1 U16339 ( .A(n9575), .B(n10304), .ZN(n9576) );
  NAND2_X1 U16342 ( .A1(n9579), .A2(n24906), .ZN(n9585) );
  NAND4_X1 U16343 ( .A1(n9581), .A2(n9582), .A3(n1196), .A4(n9580), .ZN(n9584)
         );
  NAND3_X1 U16344 ( .A1(n9585), .A2(n9584), .A3(n9583), .ZN(n9586) );
  XNOR2_X1 U16345 ( .A(n9586), .B(n10392), .ZN(n9587) );
  XNOR2_X1 U16346 ( .A(n9587), .B(n9836), .ZN(n9589) );
  XNOR2_X1 U16347 ( .A(n10143), .B(n9716), .ZN(n9588) );
  XNOR2_X1 U16348 ( .A(n9757), .B(n9588), .ZN(n9938) );
  XNOR2_X1 U16349 ( .A(n9589), .B(n9938), .ZN(n11252) );
  XNOR2_X1 U16350 ( .A(n9592), .B(n10434), .ZN(n10314) );
  XNOR2_X1 U16351 ( .A(n10071), .B(n3643), .ZN(n9593) );
  XNOR2_X1 U16352 ( .A(n9593), .B(n10314), .ZN(n9594) );
  XNOR2_X1 U16353 ( .A(n9595), .B(n9594), .ZN(n10524) );
  INV_X1 U16354 ( .A(n10524), .ZN(n10833) );
  XNOR2_X1 U16355 ( .A(n9596), .B(n10294), .ZN(n9919) );
  INV_X1 U16356 ( .A(n9919), .ZN(n9600) );
  XNOR2_X1 U16357 ( .A(n9799), .B(n3414), .ZN(n9597) );
  XNOR2_X1 U16358 ( .A(n10298), .B(n9597), .ZN(n9598) );
  XNOR2_X1 U16359 ( .A(n9598), .B(n9831), .ZN(n9599) );
  XNOR2_X1 U16361 ( .A(n10160), .B(n3317), .ZN(n9602) );
  INV_X1 U16362 ( .A(n9601), .ZN(n10409) );
  XNOR2_X1 U16363 ( .A(n9602), .B(n10409), .ZN(n9604) );
  XNOR2_X1 U16364 ( .A(n9604), .B(n9603), .ZN(n9607) );
  INV_X1 U16365 ( .A(n10282), .ZN(n9605) );
  XNOR2_X1 U16366 ( .A(n9606), .B(n9605), .ZN(n9947) );
  XNOR2_X1 U16367 ( .A(n9607), .B(n9947), .ZN(n10834) );
  MUX2_X1 U16369 ( .A(n11355), .B(n10476), .S(n11349), .Z(n9611) );
  INV_X1 U16370 ( .A(n9608), .ZN(n11351) );
  NAND2_X1 U16371 ( .A1(n11351), .A2(n11347), .ZN(n9609) );
  INV_X1 U16372 ( .A(n10847), .ZN(n11352) );
  OAI22_X1 U16373 ( .A1(n9609), .A2(n11349), .B1(n11352), .B2(n11351), .ZN(
        n9610) );
  AOI21_X2 U16374 ( .B1(n9611), .B2(n3161), .A(n9610), .ZN(n12110) );
  XNOR2_X1 U16376 ( .A(n9612), .B(n9613), .ZN(n10170) );
  INV_X1 U16377 ( .A(n10170), .ZN(n9616) );
  XNOR2_X1 U16378 ( .A(n9614), .B(n1892), .ZN(n9615) );
  XNOR2_X1 U16379 ( .A(n9616), .B(n9615), .ZN(n9618) );
  XNOR2_X1 U16381 ( .A(n9677), .B(n1853), .ZN(n9622) );
  INV_X1 U16382 ( .A(Key[122]), .ZN(n15576) );
  XNOR2_X1 U16383 ( .A(n9622), .B(n9621), .ZN(n9623) );
  NAND2_X1 U16384 ( .A1(n28204), .A2(n11045), .ZN(n9644) );
  XNOR2_X1 U16385 ( .A(n9684), .B(n10202), .ZN(n9625) );
  XNOR2_X1 U16386 ( .A(n10144), .B(n26531), .ZN(n9624) );
  XNOR2_X1 U16387 ( .A(n9625), .B(n9624), .ZN(n9628) );
  XNOR2_X1 U16388 ( .A(n9626), .B(n9996), .ZN(n10393) );
  INV_X1 U16389 ( .A(n10393), .ZN(n9627) );
  XNOR2_X1 U16390 ( .A(n10072), .B(n9629), .ZN(n9630) );
  XNOR2_X1 U16391 ( .A(n9631), .B(n9630), .ZN(n9635) );
  XNOR2_X1 U16392 ( .A(n10128), .B(n10436), .ZN(n9633) );
  INV_X1 U16393 ( .A(n3276), .ZN(n28013) );
  XNOR2_X1 U16394 ( .A(n10350), .B(n28013), .ZN(n9632) );
  XNOR2_X1 U16395 ( .A(n9633), .B(n9632), .ZN(n9634) );
  XNOR2_X1 U16396 ( .A(n10362), .B(n9878), .ZN(n9638) );
  INV_X1 U16397 ( .A(n2996), .ZN(n9636) );
  XNOR2_X1 U16398 ( .A(n9656), .B(n9636), .ZN(n9637) );
  XNOR2_X1 U16399 ( .A(n9638), .B(n9637), .ZN(n9643) );
  INV_X1 U16400 ( .A(n9639), .ZN(n9640) );
  XNOR2_X1 U16401 ( .A(n9794), .B(n9640), .ZN(n9641) );
  XNOR2_X1 U16402 ( .A(n10424), .B(n9641), .ZN(n9642) );
  XNOR2_X1 U16403 ( .A(n9642), .B(n9643), .ZN(n10528) );
  OAI22_X1 U16404 ( .A1(n9644), .A2(n11044), .B1(n11264), .B2(n28204), .ZN(
        n9654) );
  XNOR2_X1 U16405 ( .A(n9645), .B(n9986), .ZN(n10048) );
  XNOR2_X1 U16406 ( .A(n9646), .B(n10048), .ZN(n9652) );
  XNOR2_X1 U16407 ( .A(n9647), .B(n10159), .ZN(n9650) );
  XNOR2_X1 U16408 ( .A(n9648), .B(n1919), .ZN(n9649) );
  XNOR2_X1 U16409 ( .A(n9650), .B(n9649), .ZN(n9651) );
  NAND2_X1 U16410 ( .A1(n28204), .A2(n11267), .ZN(n11043) );
  XNOR2_X1 U16411 ( .A(n9656), .B(n1046), .ZN(n9657) );
  XNOR2_X1 U16412 ( .A(n10303), .B(n9657), .ZN(n9659) );
  INV_X1 U16413 ( .A(n9660), .ZN(n9664) );
  XNOR2_X1 U16416 ( .A(n9664), .B(n9663), .ZN(n9667) );
  XNOR2_X1 U16417 ( .A(n10295), .B(n9971), .ZN(n9665) );
  XNOR2_X1 U16418 ( .A(n9665), .B(n9732), .ZN(n9701) );
  XNOR2_X1 U16419 ( .A(n10072), .B(n10352), .ZN(n9670) );
  INV_X1 U16420 ( .A(n9668), .ZN(n9669) );
  XNOR2_X1 U16421 ( .A(n9669), .B(n9670), .ZN(n9673) );
  XNOR2_X1 U16422 ( .A(n9941), .B(n3537), .ZN(n9671) );
  INV_X1 U16423 ( .A(n9908), .ZN(n9922) );
  XNOR2_X1 U16424 ( .A(n9922), .B(n9674), .ZN(n9676) );
  XNOR2_X1 U16425 ( .A(n9676), .B(n9675), .ZN(n9682) );
  XNOR2_X1 U16426 ( .A(n9677), .B(n9678), .ZN(n9680) );
  XNOR2_X1 U16427 ( .A(n10022), .B(n2577), .ZN(n9679) );
  XNOR2_X1 U16428 ( .A(n9680), .B(n9679), .ZN(n9681) );
  XNOR2_X1 U16429 ( .A(n9681), .B(n9682), .ZN(n10855) );
  XNOR2_X1 U16430 ( .A(n9997), .B(n2522), .ZN(n9685) );
  XNOR2_X1 U16431 ( .A(n10046), .B(n9687), .ZN(n9691) );
  XNOR2_X1 U16432 ( .A(n10159), .B(n9949), .ZN(n9689) );
  XNOR2_X1 U16433 ( .A(n9725), .B(n2946), .ZN(n9688) );
  XNOR2_X1 U16434 ( .A(n9689), .B(n9688), .ZN(n9690) );
  XNOR2_X1 U16438 ( .A(n9695), .B(n1175), .ZN(n9697) );
  XNOR2_X1 U16439 ( .A(n9697), .B(n9696), .ZN(n9699) );
  XNOR2_X1 U16440 ( .A(n10342), .B(n9699), .ZN(n9700) );
  XNOR2_X1 U16441 ( .A(n9700), .B(n9701), .ZN(n10622) );
  INV_X1 U16442 ( .A(n10622), .ZN(n9709) );
  INV_X1 U16443 ( .A(n9964), .ZN(n9702) );
  XNOR2_X1 U16446 ( .A(n9705), .B(n9706), .ZN(n9707) );
  XNOR2_X2 U16447 ( .A(n9708), .B(n9707), .ZN(n10797) );
  NAND2_X1 U16448 ( .A1(n9709), .A2(n10797), .ZN(n10569) );
  XNOR2_X1 U16449 ( .A(n9710), .B(n9711), .ZN(n9713) );
  XNOR2_X1 U16450 ( .A(n9712), .B(n9713), .ZN(n9714) );
  XNOR2_X1 U16451 ( .A(n10391), .B(n9991), .ZN(n9715) );
  XNOR2_X1 U16452 ( .A(n10376), .B(n9715), .ZN(n9720) );
  XNOR2_X1 U16453 ( .A(n9313), .B(n2381), .ZN(n9718) );
  XNOR2_X1 U16454 ( .A(n9716), .B(n9717), .ZN(n10223) );
  XNOR2_X1 U16455 ( .A(n9718), .B(n10223), .ZN(n9719) );
  INV_X1 U16456 ( .A(n11227), .ZN(n10795) );
  XNOR2_X1 U16457 ( .A(n10330), .B(n9746), .ZN(n9723) );
  XNOR2_X1 U16458 ( .A(n9723), .B(n9724), .ZN(n9729) );
  XNOR2_X1 U16459 ( .A(n1917), .B(n9725), .ZN(n9727) );
  INV_X1 U16460 ( .A(n21865), .ZN(n27737) );
  XNOR2_X1 U16461 ( .A(n10232), .B(n27737), .ZN(n9726) );
  XNOR2_X1 U16462 ( .A(n9727), .B(n9726), .ZN(n9728) );
  XNOR2_X1 U16463 ( .A(n9729), .B(n9728), .ZN(n11225) );
  NAND2_X1 U16464 ( .A1(n28568), .A2(n11225), .ZN(n11231) );
  NAND2_X1 U16465 ( .A1(n10797), .A2(n11227), .ZN(n11898) );
  AOI21_X1 U16466 ( .B1(n11231), .B2(n11898), .A(n11099), .ZN(n9730) );
  INV_X1 U16467 ( .A(n12198), .ZN(n11818) );
  XNOR2_X1 U16468 ( .A(n10134), .B(n9732), .ZN(n9734) );
  XNOR2_X1 U16469 ( .A(n10038), .B(n2441), .ZN(n9733) );
  XNOR2_X1 U16470 ( .A(n9733), .B(n9734), .ZN(n9739) );
  XNOR2_X1 U16471 ( .A(n9915), .B(n9735), .ZN(n9737) );
  XNOR2_X1 U16472 ( .A(n9737), .B(n9736), .ZN(n9738) );
  INV_X1 U16473 ( .A(n11237), .ZN(n10628) );
  XNOR2_X1 U16474 ( .A(n9741), .B(n9740), .ZN(n9745) );
  XNOR2_X1 U16475 ( .A(n9742), .B(n9743), .ZN(n9744) );
  XNOR2_X1 U16476 ( .A(n9949), .B(n9746), .ZN(n9747) );
  XNOR2_X1 U16477 ( .A(n9748), .B(n9747), .ZN(n9753) );
  INV_X1 U16478 ( .A(n10231), .ZN(n10158) );
  XNOR2_X1 U16479 ( .A(n9749), .B(n10158), .ZN(n9751) );
  XNOR2_X1 U16481 ( .A(n9751), .B(n9750), .ZN(n9752) );
  XNOR2_X1 U16482 ( .A(n9753), .B(n9752), .ZN(n11013) );
  XNOR2_X1 U16483 ( .A(n9754), .B(n9755), .ZN(n9756) );
  XNOR2_X1 U16484 ( .A(n10287), .B(n9756), .ZN(n9761) );
  XNOR2_X1 U16485 ( .A(n9757), .B(n301), .ZN(n9759) );
  XNOR2_X1 U16486 ( .A(n10144), .B(n2541), .ZN(n9758) );
  XNOR2_X1 U16487 ( .A(n9759), .B(n9758), .ZN(n9760) );
  XNOR2_X1 U16488 ( .A(n9761), .B(n9760), .ZN(n11236) );
  NAND2_X1 U16489 ( .A1(n11013), .A2(n11236), .ZN(n11233) );
  INV_X1 U16490 ( .A(n11233), .ZN(n9762) );
  NAND2_X1 U16491 ( .A1(n9762), .A2(n5710), .ZN(n9778) );
  XNOR2_X1 U16492 ( .A(n9763), .B(n10272), .ZN(n9765) );
  INV_X1 U16493 ( .A(n10315), .ZN(n9764) );
  XNOR2_X1 U16494 ( .A(n9765), .B(n9764), .ZN(n9769) );
  XNOR2_X1 U16495 ( .A(n10357), .B(n2476), .ZN(n9766) );
  XNOR2_X1 U16496 ( .A(n9767), .B(n9766), .ZN(n9768) );
  XNOR2_X1 U16497 ( .A(n10319), .B(n9770), .ZN(n9776) );
  XNOR2_X1 U16498 ( .A(n9772), .B(n9771), .ZN(n9774) );
  INV_X1 U16499 ( .A(n22489), .ZN(n28007) );
  XNOR2_X1 U16500 ( .A(n10151), .B(n28007), .ZN(n9773) );
  XNOR2_X1 U16501 ( .A(n9774), .B(n9773), .ZN(n9775) );
  INV_X1 U16502 ( .A(n11235), .ZN(n11014) );
  INV_X1 U16503 ( .A(n11236), .ZN(n10776) );
  OAI211_X1 U16504 ( .C1(n3441), .C2(n1381), .A(n11014), .B(n10776), .ZN(n9777) );
  XNOR2_X1 U16505 ( .A(n10080), .B(n9780), .ZN(n9784) );
  XNOR2_X1 U16506 ( .A(n10395), .B(n28327), .ZN(n9781) );
  XNOR2_X1 U16507 ( .A(n9782), .B(n9781), .ZN(n9783) );
  XNOR2_X1 U16508 ( .A(n9784), .B(n9783), .ZN(n10990) );
  XNOR2_X1 U16509 ( .A(n28488), .B(n10385), .ZN(n9787) );
  INV_X1 U16510 ( .A(n10059), .ZN(n9788) );
  XNOR2_X1 U16511 ( .A(n9788), .B(n10384), .ZN(n9790) );
  XNOR2_X1 U16512 ( .A(n9979), .B(n3644), .ZN(n9789) );
  XNOR2_X1 U16513 ( .A(n9790), .B(n9789), .ZN(n9791) );
  INV_X1 U16514 ( .A(n10990), .ZN(n10785) );
  XNOR2_X1 U16515 ( .A(n9794), .B(n9795), .ZN(n10120) );
  INV_X1 U16516 ( .A(n10120), .ZN(n10085) );
  XNOR2_X1 U16517 ( .A(n10264), .B(n28294), .ZN(n9796) );
  XNOR2_X1 U16518 ( .A(n9796), .B(n10364), .ZN(n9797) );
  XNOR2_X1 U16519 ( .A(n10085), .B(n9797), .ZN(n9798) );
  XNOR2_X1 U16520 ( .A(n9799), .B(n9661), .ZN(n10135) );
  INV_X1 U16521 ( .A(n10135), .ZN(n9801) );
  XNOR2_X1 U16522 ( .A(n10257), .B(n10297), .ZN(n9800) );
  XNOR2_X1 U16523 ( .A(n9801), .B(n9800), .ZN(n9804) );
  XNOR2_X1 U16524 ( .A(n10138), .B(n27105), .ZN(n9802) );
  XNOR2_X1 U16525 ( .A(n10173), .B(n9802), .ZN(n9803) );
  INV_X1 U16526 ( .A(n10992), .ZN(n10791) );
  NAND3_X1 U16527 ( .A1(n10693), .A2(n10691), .A3(n10791), .ZN(n9816) );
  XNOR2_X1 U16528 ( .A(n10283), .B(n10159), .ZN(n9805) );
  XNOR2_X1 U16529 ( .A(n10227), .B(n9948), .ZN(n9807) );
  XNOR2_X1 U16530 ( .A(n10160), .B(n3742), .ZN(n9806) );
  XNOR2_X1 U16531 ( .A(n9807), .B(n9806), .ZN(n9808) );
  NAND3_X1 U16532 ( .A1(n10995), .A2(n10993), .A3(n4538), .ZN(n9815) );
  XNOR2_X1 U16533 ( .A(n10275), .B(n3565), .ZN(n9810) );
  MUX2_X1 U16537 ( .A(n11818), .B(n12189), .S(n12190), .Z(n9868) );
  XNOR2_X1 U16538 ( .A(n9818), .B(n9817), .ZN(n9822) );
  XNOR2_X1 U16539 ( .A(n10088), .B(n26032), .ZN(n9819) );
  XNOR2_X1 U16540 ( .A(n9820), .B(n9819), .ZN(n9821) );
  XNOR2_X1 U16541 ( .A(n9822), .B(n9821), .ZN(n10982) );
  XNOR2_X1 U16542 ( .A(n10229), .B(n9825), .ZN(n9829) );
  XNOR2_X1 U16543 ( .A(n10328), .B(n10043), .ZN(n9827) );
  XNOR2_X1 U16544 ( .A(n10183), .B(n72), .ZN(n9826) );
  XNOR2_X1 U16545 ( .A(n9827), .B(n9826), .ZN(n9828) );
  XNOR2_X1 U16546 ( .A(n9829), .B(n9828), .ZN(n10984) );
  NAND2_X1 U16547 ( .A1(n10982), .A2(n10984), .ZN(n10631) );
  XNOR2_X1 U16548 ( .A(n9870), .B(n10038), .ZN(n9830) );
  XNOR2_X1 U16549 ( .A(n9831), .B(n9830), .ZN(n9835) );
  XNOR2_X1 U16550 ( .A(n10171), .B(n2404), .ZN(n9832) );
  XNOR2_X1 U16551 ( .A(n9833), .B(n9832), .ZN(n9834) );
  NOR2_X1 U16552 ( .A1(n10989), .A2(n10982), .ZN(n10630) );
  XNOR2_X1 U16553 ( .A(n10371), .B(n10143), .ZN(n10200) );
  XNOR2_X1 U16554 ( .A(n10200), .B(n9836), .ZN(n9840) );
  XNOR2_X1 U16555 ( .A(n1868), .B(n26665), .ZN(n9837) );
  XNOR2_X1 U16556 ( .A(n9838), .B(n9837), .ZN(n9839) );
  XNOR2_X1 U16557 ( .A(n9840), .B(n9839), .ZN(n10981) );
  AND2_X1 U16558 ( .A1(n10985), .A2(n10982), .ZN(n9841) );
  NOR2_X1 U16559 ( .A1(n10630), .A2(n9841), .ZN(n9848) );
  XNOR2_X1 U16560 ( .A(n9843), .B(n9842), .ZN(n9847) );
  XNOR2_X1 U16561 ( .A(n10021), .B(n3654), .ZN(n9844) );
  XNOR2_X1 U16562 ( .A(n9845), .B(n9844), .ZN(n9846) );
  XNOR2_X1 U16563 ( .A(n9847), .B(n9846), .ZN(n10980) );
  XNOR2_X1 U16564 ( .A(n9849), .B(n9850), .ZN(n9856) );
  XNOR2_X1 U16565 ( .A(n9851), .B(n10275), .ZN(n9854) );
  XNOR2_X1 U16566 ( .A(n9852), .B(n3380), .ZN(n9853) );
  XNOR2_X1 U16567 ( .A(n9854), .B(n9853), .ZN(n9855) );
  INV_X1 U16568 ( .A(n10958), .ZN(n10686) );
  NAND2_X1 U16569 ( .A1(n10686), .A2(n10962), .ZN(n9857) );
  NAND2_X1 U16570 ( .A1(n9857), .A2(n10780), .ZN(n9862) );
  INV_X1 U16571 ( .A(n10966), .ZN(n9860) );
  NAND2_X1 U16572 ( .A1(n9862), .A2(n9861), .ZN(n12188) );
  MUX2_X1 U16573 ( .A(n10780), .B(n10687), .S(n10957), .Z(n9864) );
  NAND2_X1 U16574 ( .A1(n9864), .A2(n10958), .ZN(n12187) );
  NAND2_X1 U16575 ( .A1(n11816), .A2(n12128), .ZN(n12129) );
  NAND3_X1 U16576 ( .A1(n9865), .A2(n12194), .A3(n12190), .ZN(n9866) );
  NAND3_X1 U16577 ( .A1(n12129), .A2(n12186), .A3(n9866), .ZN(n9867) );
  XNOR2_X1 U16578 ( .A(n9869), .B(n12454), .ZN(n10444) );
  XNOR2_X1 U16579 ( .A(n9870), .B(n9915), .ZN(n9871) );
  XNOR2_X1 U16580 ( .A(n9872), .B(n9871), .ZN(n9876) );
  XNOR2_X1 U16581 ( .A(n10133), .B(n26825), .ZN(n9874) );
  XNOR2_X1 U16582 ( .A(n9873), .B(n9874), .ZN(n9875) );
  XNOR2_X1 U16583 ( .A(n9876), .B(n9875), .ZN(n9913) );
  INV_X1 U16584 ( .A(n9877), .ZN(n9879) );
  XNOR2_X1 U16585 ( .A(n9879), .B(n9878), .ZN(n9880) );
  XNOR2_X1 U16586 ( .A(n10189), .B(n9880), .ZN(n9885) );
  XNOR2_X1 U16587 ( .A(n9931), .B(n9881), .ZN(n9883) );
  XNOR2_X1 U16588 ( .A(n10088), .B(n730), .ZN(n9882) );
  XNOR2_X1 U16589 ( .A(n9883), .B(n9882), .ZN(n9884) );
  NAND2_X1 U16590 ( .A1(n11127), .A2(n11123), .ZN(n10507) );
  XNOR2_X1 U16591 ( .A(n10074), .B(n10271), .ZN(n9886) );
  XNOR2_X1 U16592 ( .A(n9887), .B(n9886), .ZN(n9891) );
  INV_X1 U16593 ( .A(n3606), .ZN(n25044) );
  XNOR2_X1 U16594 ( .A(n10128), .B(n25044), .ZN(n9889) );
  XNOR2_X1 U16595 ( .A(n9941), .B(n10435), .ZN(n9888) );
  XNOR2_X1 U16596 ( .A(n9888), .B(n9889), .ZN(n9890) );
  XNOR2_X1 U16597 ( .A(n9890), .B(n9891), .ZN(n11119) );
  INV_X1 U16598 ( .A(n11119), .ZN(n10504) );
  XNOR2_X1 U16599 ( .A(n9892), .B(n9893), .ZN(n9898) );
  XNOR2_X1 U16600 ( .A(n10396), .B(n9934), .ZN(n9896) );
  XNOR2_X1 U16601 ( .A(n1868), .B(n2987), .ZN(n9895) );
  XNOR2_X1 U16602 ( .A(n9896), .B(n9895), .ZN(n9897) );
  XNOR2_X1 U16603 ( .A(n9949), .B(n24897), .ZN(n9902) );
  INV_X1 U16605 ( .A(n10156), .ZN(n9901) );
  XNOR2_X1 U16606 ( .A(n9901), .B(n9902), .ZN(n9905) );
  XNOR2_X1 U16607 ( .A(n10229), .B(n9903), .ZN(n9904) );
  XNOR2_X1 U16608 ( .A(n9905), .B(n9904), .ZN(n10114) );
  XNOR2_X1 U16609 ( .A(n9906), .B(n9907), .ZN(n9912) );
  XNOR2_X1 U16610 ( .A(n9908), .B(n10385), .ZN(n9910) );
  XNOR2_X1 U16611 ( .A(n10060), .B(n3586), .ZN(n9909) );
  XNOR2_X1 U16612 ( .A(n9910), .B(n9909), .ZN(n9911) );
  INV_X1 U16613 ( .A(n11124), .ZN(n11126) );
  INV_X1 U16614 ( .A(n11390), .ZN(n11922) );
  XNOR2_X1 U16615 ( .A(n9915), .B(n3154), .ZN(n9917) );
  XNOR2_X1 U16616 ( .A(n9920), .B(n9919), .ZN(n10096) );
  XNOR2_X1 U16617 ( .A(n9921), .B(n3527), .ZN(n9923) );
  XNOR2_X1 U16618 ( .A(n9922), .B(n9923), .ZN(n9925) );
  XNOR2_X1 U16619 ( .A(n9924), .B(n9925), .ZN(n9927) );
  INV_X1 U16620 ( .A(n135), .ZN(n26176) );
  XNOR2_X1 U16621 ( .A(n9964), .B(n26176), .ZN(n9928) );
  XNOR2_X1 U16622 ( .A(n9931), .B(n9930), .ZN(n9932) );
  XNOR2_X1 U16623 ( .A(n9935), .B(n9934), .ZN(n9937) );
  XNOR2_X1 U16624 ( .A(n9936), .B(n9937), .ZN(n9939) );
  XNOR2_X1 U16625 ( .A(n9939), .B(n9938), .ZN(n10490) );
  INV_X1 U16626 ( .A(n10490), .ZN(n10492) );
  XNOR2_X1 U16627 ( .A(n9941), .B(n1927), .ZN(n9942) );
  XNOR2_X1 U16628 ( .A(n9943), .B(n9942), .ZN(n9944) );
  XNOR2_X1 U16629 ( .A(n9947), .B(n9946), .ZN(n9952) );
  XNOR2_X1 U16630 ( .A(n9948), .B(n3491), .ZN(n9950) );
  XNOR2_X1 U16631 ( .A(n9950), .B(n9949), .ZN(n9951) );
  INV_X1 U16632 ( .A(n10275), .ZN(n9954) );
  XNOR2_X1 U16633 ( .A(n9955), .B(n9954), .ZN(n9957) );
  XNOR2_X1 U16634 ( .A(n9956), .B(n9957), .ZN(n9960) );
  XNOR2_X1 U16635 ( .A(n10359), .B(n9958), .ZN(n9959) );
  XNOR2_X1 U16636 ( .A(n9962), .B(n9961), .ZN(n9968) );
  XNOR2_X1 U16637 ( .A(n10007), .B(n9963), .ZN(n9966) );
  XNOR2_X1 U16638 ( .A(n9964), .B(n2960), .ZN(n9965) );
  XNOR2_X1 U16639 ( .A(n9966), .B(n9965), .ZN(n9967) );
  INV_X1 U16640 ( .A(n9969), .ZN(n9970) );
  XNOR2_X1 U16641 ( .A(n9970), .B(n10342), .ZN(n9975) );
  XNOR2_X1 U16642 ( .A(n10037), .B(n10257), .ZN(n9973) );
  XNOR2_X1 U16643 ( .A(n9971), .B(n2505), .ZN(n9972) );
  XNOR2_X1 U16644 ( .A(n9973), .B(n9972), .ZN(n9974) );
  NAND2_X1 U16645 ( .A1(n5672), .A2(n10713), .ZN(n10457) );
  XNOR2_X1 U16647 ( .A(n9976), .B(n26713), .ZN(n9978) );
  XNOR2_X1 U16648 ( .A(n9978), .B(n9977), .ZN(n9983) );
  XNOR2_X1 U16649 ( .A(n10019), .B(n9979), .ZN(n9980) );
  XNOR2_X1 U16650 ( .A(n9981), .B(n9980), .ZN(n9982) );
  INV_X1 U16651 ( .A(n10498), .ZN(n11132) );
  XNOR2_X1 U16652 ( .A(n9985), .B(n9984), .ZN(n9990) );
  XNOR2_X1 U16653 ( .A(n9986), .B(n2477), .ZN(n9987) );
  XNOR2_X1 U16654 ( .A(n9988), .B(n9987), .ZN(n9989) );
  XNOR2_X1 U16655 ( .A(n9989), .B(n9990), .ZN(n10715) );
  INV_X1 U16656 ( .A(n10715), .ZN(n10500) );
  OAI21_X1 U16657 ( .B1(n10498), .B2(n10500), .A(n10502), .ZN(n10003) );
  XNOR2_X1 U16658 ( .A(n10392), .B(n9991), .ZN(n9995) );
  INV_X1 U16659 ( .A(n9992), .ZN(n9993) );
  XNOR2_X1 U16660 ( .A(n9993), .B(n10218), .ZN(n9994) );
  XNOR2_X1 U16661 ( .A(n9995), .B(n9994), .ZN(n10001) );
  XNOR2_X1 U16662 ( .A(n9996), .B(n301), .ZN(n9999) );
  XNOR2_X1 U16663 ( .A(n9997), .B(n3374), .ZN(n9998) );
  XNOR2_X1 U16664 ( .A(n9998), .B(n9999), .ZN(n10000) );
  XNOR2_X1 U16665 ( .A(n10000), .B(n10001), .ZN(n10711) );
  NAND2_X1 U16666 ( .A1(n10711), .A2(n1834), .ZN(n10714) );
  INV_X1 U16667 ( .A(n10714), .ZN(n10002) );
  INV_X1 U16668 ( .A(n10005), .ZN(n10006) );
  XNOR2_X1 U16669 ( .A(n10006), .B(n10425), .ZN(n10013) );
  XNOR2_X1 U16670 ( .A(n10007), .B(n28616), .ZN(n10011) );
  XNOR2_X1 U16671 ( .A(n10009), .B(n3516), .ZN(n10010) );
  XNOR2_X1 U16672 ( .A(n10010), .B(n10011), .ZN(n10012) );
  XNOR2_X2 U16673 ( .A(n10013), .B(n10012), .ZN(n11136) );
  INV_X1 U16674 ( .A(n11136), .ZN(n10718) );
  XNOR2_X1 U16675 ( .A(n10436), .B(n3372), .ZN(n10014) );
  XNOR2_X1 U16676 ( .A(n10015), .B(n10014), .ZN(n10017) );
  XNOR2_X1 U16677 ( .A(n10311), .B(n10073), .ZN(n10016) );
  INV_X1 U16678 ( .A(n11142), .ZN(n10920) );
  XNOR2_X1 U16679 ( .A(n10019), .B(n10250), .ZN(n10020) );
  XNOR2_X1 U16680 ( .A(n10382), .B(n10020), .ZN(n10026) );
  XNOR2_X1 U16681 ( .A(n10059), .B(n10021), .ZN(n10024) );
  XNOR2_X1 U16682 ( .A(n10022), .B(n26680), .ZN(n10023) );
  XNOR2_X1 U16683 ( .A(n10024), .B(n10023), .ZN(n10025) );
  XNOR2_X1 U16684 ( .A(n10026), .B(n10025), .ZN(n11140) );
  XNOR2_X1 U16685 ( .A(n5412), .B(n10028), .ZN(n10081) );
  XNOR2_X1 U16686 ( .A(n10029), .B(n1179), .ZN(n10030) );
  INV_X1 U16687 ( .A(n11135), .ZN(n10031) );
  XNOR2_X1 U16690 ( .A(n10034), .B(n10033), .ZN(n10036) );
  INV_X1 U16691 ( .A(n10418), .ZN(n10035) );
  XNOR2_X1 U16692 ( .A(n10036), .B(n10035), .ZN(n10042) );
  XNOR2_X1 U16693 ( .A(n28643), .B(n10037), .ZN(n10040) );
  XNOR2_X1 U16694 ( .A(n10038), .B(n1062), .ZN(n10039) );
  XNOR2_X1 U16695 ( .A(n10040), .B(n10039), .ZN(n10041) );
  XNOR2_X1 U16696 ( .A(n10043), .B(n3695), .ZN(n10044) );
  XNOR2_X1 U16697 ( .A(n10045), .B(n10044), .ZN(n10047) );
  XNOR2_X1 U16698 ( .A(n10047), .B(n10046), .ZN(n10049) );
  XNOR2_X1 U16699 ( .A(n10048), .B(n10064), .ZN(n10415) );
  OAI21_X1 U16700 ( .B1(n10458), .B2(n10726), .A(n10051), .ZN(n10054) );
  OAI21_X1 U16701 ( .B1(n10932), .B2(n10930), .A(n10927), .ZN(n10053) );
  NOR2_X1 U16702 ( .A1(n588), .A2(n10928), .ZN(n10052) );
  INV_X1 U16704 ( .A(n11853), .ZN(n11924) );
  XNOR2_X1 U16705 ( .A(n10345), .B(n1248), .ZN(n10056) );
  XNOR2_X1 U16706 ( .A(n10057), .B(n10056), .ZN(n10058) );
  XNOR2_X1 U16707 ( .A(n10059), .B(n1852), .ZN(n10176) );
  XNOR2_X1 U16708 ( .A(n10060), .B(n27894), .ZN(n10061) );
  XNOR2_X1 U16709 ( .A(n10176), .B(n10061), .ZN(n10062) );
  XNOR2_X1 U16710 ( .A(n10159), .B(n10064), .ZN(n10066) );
  XNOR2_X1 U16711 ( .A(n10065), .B(n10066), .ZN(n10070) );
  XNOR2_X1 U16712 ( .A(n10160), .B(n3622), .ZN(n10067) );
  XNOR2_X1 U16713 ( .A(n10068), .B(n10067), .ZN(n10069) );
  XNOR2_X1 U16714 ( .A(n10072), .B(n10071), .ZN(n10126) );
  XNOR2_X1 U16715 ( .A(n10432), .B(n10126), .ZN(n10078) );
  XNOR2_X1 U16716 ( .A(n10074), .B(n10073), .ZN(n10076) );
  XNOR2_X1 U16717 ( .A(n10350), .B(n22072), .ZN(n10075) );
  XNOR2_X1 U16718 ( .A(n10076), .B(n10075), .ZN(n10077) );
  INV_X1 U16719 ( .A(n10556), .ZN(n11153) );
  XNOR2_X1 U16720 ( .A(n10080), .B(n10079), .ZN(n10084) );
  XNOR2_X1 U16721 ( .A(n10219), .B(n3423), .ZN(n10082) );
  XNOR2_X1 U16722 ( .A(n10082), .B(n10081), .ZN(n10083) );
  XNOR2_X1 U16723 ( .A(n10087), .B(n10362), .ZN(n10190) );
  INV_X1 U16724 ( .A(n10190), .ZN(n10090) );
  XNOR2_X1 U16725 ( .A(n10088), .B(n2544), .ZN(n10089) );
  MUX2_X1 U16726 ( .A(n4788), .B(n593), .S(n11154), .Z(n10092) );
  INV_X1 U16727 ( .A(n10096), .ZN(n11115) );
  INV_X1 U16728 ( .A(n10097), .ZN(n10549) );
  MUX2_X1 U16729 ( .A(n10099), .B(n10098), .S(n29150), .Z(n10100) );
  NOR2_X1 U16730 ( .A1(n10502), .A2(n10715), .ZN(n10101) );
  NOR2_X1 U16731 ( .A1(n3862), .A2(n11136), .ZN(n10103) );
  NAND3_X1 U16732 ( .A1(n3862), .A2(n10919), .A3(n11136), .ZN(n10104) );
  MUX2_X1 U16733 ( .A(n10108), .B(n10932), .S(n10927), .Z(n10109) );
  INV_X1 U16734 ( .A(n10705), .ZN(n10946) );
  INV_X1 U16735 ( .A(n10592), .ZN(n10593) );
  NAND2_X1 U16736 ( .A1(n10593), .A2(n28495), .ZN(n10113) );
  NAND2_X1 U16737 ( .A1(n10110), .A2(n10703), .ZN(n10943) );
  OAI211_X1 U16738 ( .C1(n28176), .C2(n10592), .A(n10943), .B(n10942), .ZN(
        n10112) );
  INV_X1 U16739 ( .A(n10942), .ZN(n10445) );
  NAND3_X1 U16740 ( .A1(n1865), .A2(n10593), .A3(n10445), .ZN(n10111) );
  INV_X1 U16741 ( .A(n10114), .ZN(n11122) );
  AOI21_X1 U16742 ( .B1(n11120), .B2(n11126), .A(n11122), .ZN(n10116) );
  NAND2_X1 U16743 ( .A1(n10540), .A2(n11119), .ZN(n10115) );
  XNOR2_X1 U16744 ( .A(n13219), .B(n13167), .ZN(n10442) );
  XNOR2_X1 U16745 ( .A(n10120), .B(n10119), .ZN(n10125) );
  INV_X1 U16746 ( .A(n2916), .ZN(n10121) );
  XNOR2_X1 U16747 ( .A(n10265), .B(n10121), .ZN(n10122) );
  XNOR2_X1 U16748 ( .A(n10123), .B(n10122), .ZN(n10124) );
  XNOR2_X1 U16749 ( .A(n10126), .B(n10127), .ZN(n10132) );
  XNOR2_X1 U16750 ( .A(n10207), .B(n10272), .ZN(n10130) );
  XNOR2_X1 U16751 ( .A(n10128), .B(n3081), .ZN(n10129) );
  XNOR2_X1 U16752 ( .A(n10130), .B(n10129), .ZN(n10131) );
  XNOR2_X1 U16753 ( .A(n10132), .B(n10131), .ZN(n10882) );
  AND2_X1 U16754 ( .A1(n10882), .A2(n11210), .ZN(n10572) );
  XNOR2_X1 U16755 ( .A(n10134), .B(n10133), .ZN(n10136) );
  XNOR2_X1 U16756 ( .A(n10135), .B(n10136), .ZN(n10142) );
  XNOR2_X1 U16757 ( .A(n10137), .B(n10171), .ZN(n10140) );
  XNOR2_X1 U16758 ( .A(n10138), .B(n3134), .ZN(n10139) );
  XNOR2_X1 U16759 ( .A(n10140), .B(n10139), .ZN(n10141) );
  XNOR2_X1 U16760 ( .A(n10146), .B(n28634), .ZN(n10147) );
  XNOR2_X1 U16761 ( .A(n10149), .B(n28488), .ZN(n10150) );
  XNOR2_X1 U16762 ( .A(n10178), .B(n3666), .ZN(n10153) );
  XNOR2_X1 U16763 ( .A(n10152), .B(n10153), .ZN(n10154) );
  NAND3_X1 U16764 ( .A1(n11084), .A2(n11209), .A3(n11086), .ZN(n10166) );
  XNOR2_X1 U16765 ( .A(n10156), .B(n10157), .ZN(n10164) );
  XNOR2_X1 U16766 ( .A(n10159), .B(n10158), .ZN(n10162) );
  XNOR2_X1 U16767 ( .A(n10160), .B(n2961), .ZN(n10161) );
  XNOR2_X1 U16768 ( .A(n10162), .B(n10161), .ZN(n10163) );
  XNOR2_X1 U16769 ( .A(n10163), .B(n10164), .ZN(n11085) );
  NAND2_X1 U16770 ( .A1(n11084), .A2(n28624), .ZN(n11216) );
  NOR2_X1 U16771 ( .A1(n11216), .A2(n11209), .ZN(n10167) );
  XNOR2_X1 U16772 ( .A(n10169), .B(n10170), .ZN(n10175) );
  XNOR2_X1 U16773 ( .A(n10171), .B(n2389), .ZN(n10172) );
  XNOR2_X1 U16774 ( .A(n10173), .B(n10172), .ZN(n10174) );
  XNOR2_X1 U16775 ( .A(n10176), .B(n10177), .ZN(n10182) );
  XNOR2_X1 U16776 ( .A(n10178), .B(n3109), .ZN(n10180) );
  XNOR2_X1 U16777 ( .A(n10179), .B(n10180), .ZN(n10181) );
  XNOR2_X1 U16778 ( .A(n10183), .B(n27298), .ZN(n10186) );
  XNOR2_X1 U16779 ( .A(n10185), .B(n10186), .ZN(n10187) );
  INV_X1 U16780 ( .A(n11243), .ZN(n10640) );
  XNOR2_X1 U16781 ( .A(n10190), .B(n10189), .ZN(n10197) );
  XNOR2_X1 U16782 ( .A(n10191), .B(n10192), .ZN(n10195) );
  XNOR2_X1 U16783 ( .A(n10193), .B(n2510), .ZN(n10194) );
  XNOR2_X1 U16784 ( .A(n10195), .B(n10194), .ZN(n10196) );
  OAI211_X1 U16786 ( .C1(n1900), .C2(n11242), .A(n10640), .B(n10198), .ZN(
        n10217) );
  XNOR2_X1 U16787 ( .A(n10200), .B(n10199), .ZN(n10206) );
  XNOR2_X1 U16788 ( .A(n10201), .B(n10396), .ZN(n10204) );
  XNOR2_X1 U16789 ( .A(n10202), .B(n4029), .ZN(n10203) );
  XNOR2_X1 U16790 ( .A(n10204), .B(n10203), .ZN(n10205) );
  NAND3_X1 U16791 ( .A1(n1900), .A2(n11240), .A3(n11243), .ZN(n10216) );
  XNOR2_X1 U16792 ( .A(n10208), .B(n10207), .ZN(n10210) );
  XNOR2_X1 U16793 ( .A(n10210), .B(n10209), .ZN(n10214) );
  INV_X1 U16794 ( .A(n21537), .ZN(n27669) );
  XNOR2_X1 U16795 ( .A(n10350), .B(n27669), .ZN(n10211) );
  XNOR2_X1 U16796 ( .A(n10212), .B(n10211), .ZN(n10213) );
  NAND3_X1 U16797 ( .A1(n10880), .A2(n11069), .A3(n11066), .ZN(n10215) );
  XNOR2_X1 U16798 ( .A(n10219), .B(n10218), .ZN(n10221) );
  XNOR2_X1 U16799 ( .A(n10220), .B(n10221), .ZN(n10226) );
  INV_X1 U16800 ( .A(n2306), .ZN(n27850) );
  XNOR2_X1 U16801 ( .A(n10222), .B(n27850), .ZN(n10224) );
  XNOR2_X1 U16802 ( .A(n10223), .B(n10224), .ZN(n10225) );
  XNOR2_X1 U16803 ( .A(n10225), .B(n10226), .ZN(n11218) );
  XNOR2_X1 U16804 ( .A(n10227), .B(n10228), .ZN(n10230) );
  XNOR2_X1 U16805 ( .A(n10229), .B(n10230), .ZN(n10249) );
  XNOR2_X1 U16806 ( .A(n10232), .B(n10231), .ZN(n10248) );
  INV_X1 U16807 ( .A(n10233), .ZN(n10236) );
  INV_X1 U16808 ( .A(n10234), .ZN(n10235) );
  NAND3_X1 U16809 ( .A1(n10237), .A2(n10236), .A3(n10235), .ZN(n10239) );
  INV_X1 U16810 ( .A(n3116), .ZN(n27605) );
  NAND2_X1 U16811 ( .A1(n10237), .A2(n10241), .ZN(n10238) );
  NAND3_X1 U16812 ( .A1(n10239), .A2(n27605), .A3(n10238), .ZN(n10244) );
  INV_X1 U16813 ( .A(n10240), .ZN(n10242) );
  NAND3_X1 U16814 ( .A1(n10242), .A2(n10241), .A3(n27605), .ZN(n10243) );
  OAI211_X1 U16815 ( .C1(n10246), .C2(n10245), .A(n10244), .B(n10243), .ZN(
        n10247) );
  XNOR2_X1 U16816 ( .A(n10254), .B(n10253), .ZN(n10657) );
  XNOR2_X1 U16817 ( .A(n10256), .B(n10255), .ZN(n10262) );
  XNOR2_X1 U16818 ( .A(n10295), .B(n10257), .ZN(n10260) );
  XNOR2_X1 U16819 ( .A(n10258), .B(n1928), .ZN(n10259) );
  XNOR2_X1 U16820 ( .A(n10260), .B(n10259), .ZN(n10261) );
  NOR2_X1 U16821 ( .A1(n11222), .A2(n10876), .ZN(n10269) );
  XNOR2_X1 U16822 ( .A(n10264), .B(n10263), .ZN(n10267) );
  XNOR2_X1 U16823 ( .A(n10265), .B(n3036), .ZN(n10266) );
  XNOR2_X1 U16825 ( .A(n10272), .B(n3334), .ZN(n10273) );
  XNOR2_X1 U16826 ( .A(n10274), .B(n10273), .ZN(n10279) );
  XNOR2_X1 U16827 ( .A(n10311), .B(n10275), .ZN(n10276) );
  XNOR2_X1 U16828 ( .A(n10277), .B(n10276), .ZN(n10278) );
  INV_X1 U16830 ( .A(n10876), .ZN(n10871) );
  XNOR2_X1 U16833 ( .A(n10282), .B(n2465), .ZN(n10284) );
  XNOR2_X1 U16834 ( .A(n10288), .B(n10287), .ZN(n10293) );
  XNOR2_X1 U16835 ( .A(n10289), .B(n1215), .ZN(n10290) );
  XNOR2_X1 U16836 ( .A(n10291), .B(n10290), .ZN(n10292) );
  XNOR2_X1 U16837 ( .A(n10293), .B(n10292), .ZN(n11287) );
  XNOR2_X1 U16838 ( .A(n10294), .B(n1079), .ZN(n10296) );
  XNOR2_X1 U16839 ( .A(n10295), .B(n10296), .ZN(n10299) );
  XNOR2_X1 U16840 ( .A(n10298), .B(n10297), .ZN(n10417) );
  XNOR2_X1 U16841 ( .A(n10364), .B(n10302), .ZN(n10428) );
  XNOR2_X1 U16842 ( .A(n10303), .B(n10428), .ZN(n10308) );
  XNOR2_X1 U16843 ( .A(n10304), .B(n2995), .ZN(n10305) );
  XNOR2_X1 U16844 ( .A(n10306), .B(n10305), .ZN(n10307) );
  XNOR2_X1 U16845 ( .A(n10308), .B(n10307), .ZN(n10318) );
  OAI21_X1 U16846 ( .B1(n11290), .B2(n11287), .A(n10309), .ZN(n11292) );
  XNOR2_X1 U16847 ( .A(n10310), .B(n10311), .ZN(n10313) );
  XNOR2_X1 U16848 ( .A(n10353), .B(n1133), .ZN(n10312) );
  XNOR2_X1 U16849 ( .A(n10313), .B(n10312), .ZN(n10317) );
  XNOR2_X1 U16850 ( .A(n10315), .B(n10314), .ZN(n10316) );
  XNOR2_X1 U16851 ( .A(n10316), .B(n10317), .ZN(n11075) );
  INV_X1 U16852 ( .A(n10318), .ZN(n11072) );
  XNOR2_X1 U16853 ( .A(n10319), .B(n10320), .ZN(n10326) );
  XNOR2_X1 U16854 ( .A(n10321), .B(n10384), .ZN(n10324) );
  XNOR2_X1 U16855 ( .A(n10322), .B(n2894), .ZN(n10323) );
  XNOR2_X1 U16856 ( .A(n10324), .B(n10323), .ZN(n10325) );
  AND3_X1 U16857 ( .A1(n10891), .A2(n11287), .A3(n29116), .ZN(n10327) );
  XNOR2_X1 U16858 ( .A(n10328), .B(n3049), .ZN(n10329) );
  XNOR2_X1 U16859 ( .A(n10329), .B(n10330), .ZN(n10331) );
  XNOR2_X1 U16860 ( .A(n10331), .B(n10332), .ZN(n10333) );
  XNOR2_X1 U16861 ( .A(n10333), .B(n10334), .ZN(n10518) );
  XNOR2_X1 U16862 ( .A(n10335), .B(n10384), .ZN(n10336) );
  XNOR2_X1 U16863 ( .A(n10336), .B(n10337), .ZN(n10341) );
  XNOR2_X1 U16864 ( .A(n1852), .B(n3728), .ZN(n10339) );
  XNOR2_X1 U16865 ( .A(n10338), .B(n10339), .ZN(n10340) );
  NAND2_X1 U16866 ( .A1(n11027), .A2(n11282), .ZN(n11286) );
  XNOR2_X1 U16867 ( .A(n10342), .B(n10343), .ZN(n10349) );
  XNOR2_X1 U16868 ( .A(n10344), .B(n10345), .ZN(n10348) );
  XNOR2_X1 U16869 ( .A(n28643), .B(n900), .ZN(n10347) );
  INV_X1 U16870 ( .A(n2986), .ZN(n24060) );
  XNOR2_X1 U16871 ( .A(n10350), .B(n24060), .ZN(n10351) );
  XNOR2_X1 U16872 ( .A(n10351), .B(n10352), .ZN(n10355) );
  XNOR2_X1 U16873 ( .A(n10355), .B(n10354), .ZN(n10361) );
  XNOR2_X1 U16874 ( .A(n10357), .B(n10356), .ZN(n10358) );
  XNOR2_X1 U16875 ( .A(n10359), .B(n10358), .ZN(n10360) );
  XNOR2_X1 U16876 ( .A(n10361), .B(n10360), .ZN(n10517) );
  XNOR2_X1 U16877 ( .A(n10363), .B(n10362), .ZN(n10366) );
  XNOR2_X1 U16878 ( .A(n10364), .B(n3463), .ZN(n10365) );
  XNOR2_X1 U16879 ( .A(n10366), .B(n10365), .ZN(n10370) );
  XNOR2_X1 U16880 ( .A(n10368), .B(n10367), .ZN(n10369) );
  NAND3_X1 U16881 ( .A1(n585), .A2(n10517), .A3(n10884), .ZN(n10381) );
  INV_X1 U16882 ( .A(n10517), .ZN(n11283) );
  XNOR2_X1 U16884 ( .A(n10371), .B(n10372), .ZN(n10374) );
  XNOR2_X1 U16885 ( .A(n10373), .B(n10374), .ZN(n10378) );
  XNOR2_X1 U16886 ( .A(n10395), .B(n3673), .ZN(n10375) );
  XNOR2_X1 U16887 ( .A(n10376), .B(n10375), .ZN(n10377) );
  NAND3_X1 U16888 ( .A1(n10517), .A2(n584), .A3(n11281), .ZN(n10379) );
  XNOR2_X1 U16889 ( .A(n10383), .B(n10382), .ZN(n10390) );
  XNOR2_X1 U16890 ( .A(n10384), .B(n3710), .ZN(n10388) );
  XNOR2_X1 U16891 ( .A(n10386), .B(n10385), .ZN(n10387) );
  XNOR2_X1 U16892 ( .A(n10388), .B(n10387), .ZN(n10389) );
  XNOR2_X1 U16893 ( .A(n10391), .B(n10392), .ZN(n10394) );
  XNOR2_X1 U16894 ( .A(n10393), .B(n10394), .ZN(n10400) );
  XNOR2_X1 U16895 ( .A(n10396), .B(n10395), .ZN(n10398) );
  INV_X1 U16896 ( .A(n3508), .ZN(n26899) );
  XNOR2_X1 U16897 ( .A(n5412), .B(n26899), .ZN(n10397) );
  XNOR2_X1 U16898 ( .A(n10398), .B(n10397), .ZN(n10399) );
  NOR2_X1 U16899 ( .A1(n10401), .A2(n3787), .ZN(n10402) );
  NAND3_X1 U16900 ( .A1(n10407), .A2(n3787), .A3(n10406), .ZN(n10408) );
  XNOR2_X1 U16902 ( .A(n10411), .B(n1918), .ZN(n10413) );
  XNOR2_X1 U16903 ( .A(n10414), .B(n10413), .ZN(n10416) );
  XNOR2_X1 U16904 ( .A(n10417), .B(n10418), .ZN(n10423) );
  XNOR2_X1 U16905 ( .A(n10419), .B(n3062), .ZN(n10420) );
  XNOR2_X1 U16906 ( .A(n10421), .B(n10420), .ZN(n10422) );
  XNOR2_X1 U16907 ( .A(n10422), .B(n10423), .ZN(n11204) );
  INV_X1 U16908 ( .A(n11204), .ZN(n11090) );
  XNOR2_X1 U16909 ( .A(n10425), .B(n10424), .ZN(n10430) );
  XNOR2_X1 U16910 ( .A(n10426), .B(n3598), .ZN(n10427) );
  XNOR2_X1 U16911 ( .A(n10428), .B(n10427), .ZN(n10429) );
  NOR2_X1 U16913 ( .A1(n11204), .A2(n11206), .ZN(n10637) );
  XNOR2_X1 U16914 ( .A(n10432), .B(n10433), .ZN(n10440) );
  XNOR2_X1 U16915 ( .A(n10435), .B(n10434), .ZN(n10438) );
  XNOR2_X1 U16916 ( .A(n10436), .B(n3554), .ZN(n10437) );
  XNOR2_X1 U16917 ( .A(n10438), .B(n10437), .ZN(n10439) );
  XNOR2_X1 U16918 ( .A(n10440), .B(n10439), .ZN(n11093) );
  XNOR2_X1 U16919 ( .A(n13144), .B(n10442), .ZN(n10443) );
  INV_X1 U16920 ( .A(n13606), .ZN(n14102) );
  NAND2_X1 U16921 ( .A1(n10705), .A2(n28495), .ZN(n10448) );
  NOR2_X1 U16922 ( .A1(n10592), .A2(n28495), .ZN(n10706) );
  NAND2_X1 U16923 ( .A1(n10912), .A2(n10911), .ZN(n10449) );
  NAND2_X1 U16924 ( .A1(n10732), .A2(n10449), .ZN(n10450) );
  NAND2_X1 U16925 ( .A1(n10450), .A2(n10735), .ZN(n10451) );
  NOR2_X1 U16926 ( .A1(n10711), .A2(n10715), .ZN(n10454) );
  NAND2_X1 U16927 ( .A1(n10499), .A2(n10454), .ZN(n10456) );
  OAI211_X1 U16928 ( .C1(n10457), .C2(n2646), .A(n10456), .B(n10455), .ZN(
        n10868) );
  NAND2_X1 U16929 ( .A1(n10458), .A2(n10726), .ZN(n10926) );
  NAND2_X1 U16930 ( .A1(n10926), .A2(n10459), .ZN(n10460) );
  AND3_X1 U16931 ( .A1(n3862), .A2(n11138), .A3(n10718), .ZN(n10767) );
  INV_X1 U16932 ( .A(n11876), .ZN(n10464) );
  NAND2_X1 U16933 ( .A1(n10464), .A2(n287), .ZN(n10465) );
  NOR2_X1 U16934 ( .A1(n10745), .A2(n11168), .ZN(n10471) );
  INV_X1 U16935 ( .A(n11168), .ZN(n11170) );
  NAND2_X1 U16936 ( .A1(n11166), .A2(n11170), .ZN(n10466) );
  NAND2_X1 U16937 ( .A1(n10467), .A2(n11330), .ZN(n11332) );
  NOR2_X1 U16938 ( .A1(n10821), .A2(n11170), .ZN(n10468) );
  AOI21_X1 U16939 ( .B1(n10469), .B2(n11332), .A(n10468), .ZN(n10470) );
  NAND3_X1 U16941 ( .A1(n11184), .A2(n11181), .A3(n10810), .ZN(n10474) );
  OAI21_X1 U16943 ( .B1(n11349), .B2(n11192), .A(n10478), .ZN(n10479) );
  NAND2_X1 U16944 ( .A1(n11022), .A2(n11255), .ZN(n10484) );
  NOR2_X1 U16946 ( .A1(n10855), .A2(n11165), .ZN(n10487) );
  INV_X1 U16947 ( .A(n10855), .ZN(n11164) );
  NOR2_X1 U16948 ( .A1(n11164), .A2(n11053), .ZN(n10486) );
  INV_X1 U16949 ( .A(n12338), .ZN(n11913) );
  OAI21_X1 U16950 ( .B1(n12343), .B2(n11913), .A(n12339), .ZN(n10489) );
  XNOR2_X1 U16951 ( .A(n13097), .B(n13227), .ZN(n10539) );
  AOI21_X1 U16953 ( .B1(n10554), .B2(n10494), .A(n11154), .ZN(n10495) );
  MUX2_X1 U16954 ( .A(n10499), .B(n10498), .S(n10497), .Z(n10503) );
  MUX2_X1 U16955 ( .A(n10506), .B(n10505), .S(n4024), .Z(n10509) );
  OAI21_X1 U16956 ( .B1(n11461), .B2(n1836), .A(n11874), .ZN(n10516) );
  NAND2_X1 U16958 ( .A1(n11500), .A2(n11458), .ZN(n11870) );
  INV_X1 U16962 ( .A(n10518), .ZN(n11280) );
  MUX2_X1 U16963 ( .A(n10520), .B(n10519), .S(n11284), .Z(n10521) );
  INV_X1 U16964 ( .A(n11449), .ZN(n11888) );
  INV_X1 U16966 ( .A(n11037), .ZN(n11273) );
  INV_X1 U16967 ( .A(n12328), .ZN(n11884) );
  OAI21_X1 U16968 ( .B1(n11888), .B2(n11884), .A(n11747), .ZN(n10531) );
  INV_X1 U16969 ( .A(n10528), .ZN(n11266) );
  NOR2_X1 U16970 ( .A1(n11261), .A2(n11047), .ZN(n10530) );
  NAND2_X1 U16971 ( .A1(n10530), .A2(n28204), .ZN(n11886) );
  INV_X1 U16972 ( .A(n12327), .ZN(n12333) );
  NAND2_X1 U16973 ( .A1(n10665), .A2(n11076), .ZN(n10894) );
  INV_X1 U16974 ( .A(n11287), .ZN(n10893) );
  INV_X1 U16975 ( .A(n11075), .ZN(n11291) );
  NAND2_X1 U16976 ( .A1(n11291), .A2(n11072), .ZN(n10532) );
  INV_X1 U16977 ( .A(n11223), .ZN(n10878) );
  XNOR2_X1 U16978 ( .A(n10539), .B(n10538), .ZN(n10619) );
  NOR2_X1 U16979 ( .A1(n11119), .A2(n11118), .ZN(n10542) );
  INV_X1 U16980 ( .A(n11120), .ZN(n11125) );
  NAND2_X1 U16981 ( .A1(n11125), .A2(n11124), .ZN(n10541) );
  OAI21_X1 U16982 ( .B1(n10805), .B2(n11146), .A(n10543), .ZN(n10546) );
  NOR2_X2 U16983 ( .A1(n10546), .A2(n10545), .ZN(n11754) );
  OAI21_X1 U16984 ( .B1(n10548), .B2(n10461), .A(n10547), .ZN(n10552) );
  NAND2_X1 U16985 ( .A1(n29150), .A2(n11113), .ZN(n10551) );
  OAI21_X1 U16986 ( .B1(n11111), .B2(n11113), .A(n10549), .ZN(n10550) );
  NAND2_X1 U16987 ( .A1(n10555), .A2(n11158), .ZN(n10557) );
  AOI21_X1 U16988 ( .B1(n11338), .B2(n11337), .A(n10828), .ZN(n10561) );
  NOR2_X1 U16989 ( .A1(n10558), .A2(n11176), .ZN(n10827) );
  NOR2_X1 U16990 ( .A1(n10830), .A2(n1898), .ZN(n10559) );
  OAI21_X1 U16991 ( .B1(n10827), .B2(n10559), .A(n11341), .ZN(n10560) );
  OAI21_X1 U16992 ( .B1(n11345), .B2(n10561), .A(n10560), .ZN(n11755) );
  NOR2_X1 U16993 ( .A1(n10748), .A2(n10814), .ZN(n10815) );
  NOR2_X1 U16994 ( .A1(n11198), .A2(n10563), .ZN(n10564) );
  NOR3_X1 U16996 ( .A1(n5914), .A2(n5917), .A3(n28157), .ZN(n10566) );
  XNOR2_X1 U16997 ( .A(n13226), .B(n3752), .ZN(n10617) );
  INV_X1 U16998 ( .A(n10797), .ZN(n11232) );
  INV_X1 U16999 ( .A(n11225), .ZN(n10794) );
  NAND3_X1 U17000 ( .A1(n11099), .A2(n6814), .A3(n10794), .ZN(n11899) );
  OAI211_X1 U17001 ( .C1(n11066), .C2(n11244), .A(n11240), .B(n1851), .ZN(
        n10571) );
  INV_X1 U17002 ( .A(n11240), .ZN(n11063) );
  NAND3_X1 U17003 ( .A1(n10640), .A2(n11063), .A3(n11069), .ZN(n10570) );
  NAND2_X1 U17004 ( .A1(n12352), .A2(n11901), .ZN(n11468) );
  MUX2_X1 U17005 ( .A(n11212), .B(n11213), .S(n433), .Z(n10575) );
  NAND2_X1 U17006 ( .A1(n433), .A2(n11211), .ZN(n10573) );
  OAI21_X2 U17007 ( .B1(n10575), .B2(n10574), .A(n10573), .ZN(n12350) );
  INV_X1 U17008 ( .A(n12350), .ZN(n10586) );
  AND2_X1 U17009 ( .A1(n11205), .A2(n10576), .ZN(n10578) );
  NAND2_X1 U17010 ( .A1(n10579), .A2(n11013), .ZN(n10583) );
  NAND3_X1 U17011 ( .A1(n10628), .A2(n5710), .A3(n3441), .ZN(n10582) );
  NAND2_X1 U17013 ( .A1(n29648), .A2(n11237), .ZN(n11239) );
  INV_X1 U17014 ( .A(n11239), .ZN(n10580) );
  NAND2_X1 U17015 ( .A1(n10580), .A2(n10776), .ZN(n10581) );
  AOI22_X1 U17017 ( .A1(n10989), .A2(n3804), .B1(n10983), .B2(n10984), .ZN(
        n10585) );
  MUX2_X1 U17019 ( .A(n28405), .B(n10999), .S(n11003), .Z(n10589) );
  NOR2_X1 U17020 ( .A1(n10589), .A2(n10936), .ZN(n10590) );
  NAND2_X1 U17021 ( .A1(n10592), .A2(n28495), .ZN(n10944) );
  AOI21_X1 U17023 ( .B1(n10702), .B2(n28176), .A(n10946), .ZN(n10595) );
  INV_X1 U17024 ( .A(n10995), .ZN(n10787) );
  NAND2_X1 U17025 ( .A1(n10693), .A2(n10597), .ZN(n10601) );
  OAI21_X1 U17026 ( .B1(n10992), .B2(n10991), .A(n3454), .ZN(n10600) );
  INV_X1 U17027 ( .A(n10991), .ZN(n10598) );
  NOR2_X1 U17028 ( .A1(n10598), .A2(n10787), .ZN(n10599) );
  INV_X1 U17029 ( .A(n10602), .ZN(n10964) );
  OAI21_X1 U17030 ( .B1(n896), .B2(n9858), .A(n10964), .ZN(n10604) );
  INV_X1 U17031 ( .A(n10962), .ZN(n10778) );
  NAND2_X1 U17033 ( .A1(n11740), .A2(n12356), .ZN(n10898) );
  INV_X1 U17034 ( .A(n10911), .ZN(n10915) );
  INV_X1 U17037 ( .A(n12362), .ZN(n11741) );
  AOI21_X1 U17038 ( .B1(n10611), .B2(n10898), .A(n11741), .ZN(n10616) );
  NOR2_X1 U17041 ( .A1(n10616), .A2(n10615), .ZN(n12594) );
  INV_X1 U17042 ( .A(n12594), .ZN(n13381) );
  XNOR2_X1 U17043 ( .A(n13381), .B(n12593), .ZN(n12654) );
  XNOR2_X1 U17044 ( .A(n12654), .B(n10617), .ZN(n10618) );
  XNOR2_X2 U17045 ( .A(n10619), .B(n10618), .ZN(n14593) );
  NAND2_X1 U17046 ( .A1(n14102), .A2(n14593), .ZN(n11372) );
  MUX2_X1 U17048 ( .A(n10624), .B(n10623), .S(n10797), .Z(n10625) );
  NOR2_X2 U17049 ( .A1(n10626), .A2(n10625), .ZN(n12220) );
  NOR2_X1 U17050 ( .A1(n6108), .A2(n11013), .ZN(n10627) );
  INV_X1 U17052 ( .A(n10981), .ZN(n10985) );
  INV_X1 U17053 ( .A(n10631), .ZN(n10632) );
  NAND2_X1 U17054 ( .A1(n10632), .A2(n10783), .ZN(n10633) );
  MUX2_X1 U17055 ( .A(n12220), .B(n28726), .S(n12218), .Z(n10645) );
  NAND2_X1 U17056 ( .A1(n10785), .A2(n10786), .ZN(n10635) );
  NAND2_X1 U17057 ( .A1(n10995), .A2(n10786), .ZN(n10994) );
  OAI211_X1 U17058 ( .C1(n10785), .C2(n4538), .A(n10992), .B(n10994), .ZN(
        n11693) );
  INV_X1 U17059 ( .A(n12218), .ZN(n12041) );
  INV_X1 U17060 ( .A(n10637), .ZN(n10638) );
  NOR2_X1 U17061 ( .A1(n11069), .A2(n11066), .ZN(n10639) );
  NAND3_X1 U17062 ( .A1(n11066), .A2(n11242), .A3(n11244), .ZN(n10642) );
  INV_X1 U17063 ( .A(n11066), .ZN(n10641) );
  OAI22_X1 U17064 ( .A1(n10643), .A2(n12224), .B1(n12042), .B2(n11962), .ZN(
        n10644) );
  XNOR2_X1 U17065 ( .A(n13359), .B(n3114), .ZN(n10677) );
  NAND2_X1 U17066 ( .A1(n431), .A2(n12337), .ZN(n12027) );
  NAND2_X1 U17067 ( .A1(n12343), .A2(n12338), .ZN(n10646) );
  NAND2_X1 U17069 ( .A1(n10647), .A2(n1291), .ZN(n10651) );
  AOI22_X1 U17071 ( .A1(n10649), .A2(n12026), .B1(n10648), .B2(n12339), .ZN(
        n10650) );
  NOR2_X1 U17073 ( .A1(n11280), .A2(n11282), .ZN(n10652) );
  INV_X1 U17074 ( .A(n11281), .ZN(n11029) );
  AOI22_X1 U17075 ( .A1(n10883), .A2(n11086), .B1(n11211), .B2(n11212), .ZN(
        n10656) );
  NAND2_X1 U17076 ( .A1(n1986), .A2(n375), .ZN(n11682) );
  MUX2_X1 U17077 ( .A(n11218), .B(n10872), .S(n10659), .Z(n10658) );
  NAND2_X1 U17078 ( .A1(n10659), .A2(n29593), .ZN(n10661) );
  OAI22_X1 U17079 ( .A1(n10872), .A2(n10661), .B1(n10660), .B2(n10876), .ZN(
        n10662) );
  OAI21_X1 U17080 ( .B1(n10893), .B2(n10665), .A(n10664), .ZN(n10667) );
  NAND3_X1 U17081 ( .A1(n11290), .A2(n11072), .A3(n29116), .ZN(n10666) );
  NAND2_X1 U17082 ( .A1(n11048), .A2(n11261), .ZN(n10670) );
  INV_X1 U17083 ( .A(n11047), .ZN(n10888) );
  NAND3_X1 U17084 ( .A1(n11979), .A2(n12232), .A3(n12233), .ZN(n10675) );
  OAI21_X2 U17085 ( .B1(n10673), .B2(n11274), .A(n10672), .ZN(n12234) );
  NAND4_X2 U17086 ( .A1(n11977), .A2(n10676), .A3(n10674), .A4(n10675), .ZN(
        n13337) );
  XNOR2_X1 U17087 ( .A(n12560), .B(n13337), .ZN(n13549) );
  XNOR2_X1 U17088 ( .A(n13549), .B(n10677), .ZN(n10773) );
  NAND2_X1 U17089 ( .A1(n10973), .A2(n29577), .ZN(n10679) );
  MUX2_X1 U17090 ( .A(n10679), .B(n10678), .S(n10681), .Z(n11495) );
  MUX2_X1 U17091 ( .A(n10936), .B(n6779), .S(n10937), .Z(n10685) );
  INV_X1 U17092 ( .A(n12304), .ZN(n10701) );
  OAI21_X1 U17093 ( .B1(n10913), .B2(n10916), .A(n10688), .ZN(n10737) );
  NAND2_X1 U17094 ( .A1(n10690), .A2(n10913), .ZN(n11494) );
  NAND2_X1 U17095 ( .A1(n10791), .A2(n3454), .ZN(n10692) );
  NAND2_X1 U17096 ( .A1(n12304), .A2(n12303), .ZN(n10700) );
  INV_X1 U17097 ( .A(n10983), .ZN(n10694) );
  MUX2_X1 U17099 ( .A(n10695), .B(n589), .S(n10783), .Z(n10699) );
  INV_X1 U17101 ( .A(n10982), .ZN(n10988) );
  NAND2_X1 U17102 ( .A1(n10701), .A2(n11491), .ZN(n11363) );
  NAND2_X1 U17104 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  OAI211_X1 U17105 ( .C1(n10710), .C2(n10110), .A(n10708), .B(n10707), .ZN(
        n11794) );
  NAND2_X1 U17106 ( .A1(n10711), .A2(n10715), .ZN(n10712) );
  AOI21_X1 U17107 ( .B1(n10715), .B2(n10714), .A(n10713), .ZN(n10716) );
  OAI21_X1 U17108 ( .B1(n3862), .B2(n2968), .A(n10919), .ZN(n10720) );
  OAI21_X1 U17109 ( .B1(n10721), .B2(n10720), .A(n10719), .ZN(n10722) );
  NAND2_X1 U17110 ( .A1(n6482), .A2(n11486), .ZN(n11718) );
  OAI21_X1 U17111 ( .B1(n10976), .B2(n29577), .A(n10970), .ZN(n10724) );
  NAND2_X1 U17112 ( .A1(n11718), .A2(n11430), .ZN(n10731) );
  OAI21_X1 U17113 ( .B1(n10924), .B2(n10927), .A(n590), .ZN(n10729) );
  NAND2_X1 U17115 ( .A1(n10731), .A2(n28436), .ZN(n10739) );
  NAND2_X1 U17116 ( .A1(n10737), .A2(n10732), .ZN(n10734) );
  NAND2_X1 U17117 ( .A1(n10734), .A2(n10733), .ZN(n11428) );
  NAND2_X1 U17118 ( .A1(n10735), .A2(n10916), .ZN(n10736) );
  INV_X1 U17120 ( .A(n11486), .ZN(n11431) );
  NAND3_X1 U17121 ( .A1(n11487), .A2(n11431), .A3(n2194), .ZN(n10738) );
  XNOR2_X1 U17122 ( .A(n13036), .B(n12919), .ZN(n12065) );
  INV_X1 U17123 ( .A(n11166), .ZN(n10819) );
  MUX2_X1 U17124 ( .A(n28638), .B(n28157), .S(n10563), .Z(n10750) );
  OAI21_X1 U17125 ( .B1(n11152), .B2(n10752), .A(n28175), .ZN(n10753) );
  NAND2_X1 U17126 ( .A1(n10753), .A2(n10803), .ZN(n10756) );
  NOR2_X1 U17128 ( .A1(n11401), .A2(n11672), .ZN(n10758) );
  INV_X1 U17129 ( .A(n10828), .ZN(n11336) );
  NAND2_X1 U17130 ( .A1(n11341), .A2(n11176), .ZN(n10757) );
  OR2_X1 U17131 ( .A1(n11340), .A2(n1898), .ZN(n11634) );
  INV_X1 U17132 ( .A(n11515), .ZN(n11845) );
  OAI21_X1 U17133 ( .B1(n11677), .B2(n10758), .A(n11845), .ZN(n10765) );
  NOR2_X1 U17134 ( .A1(n11640), .A2(n29139), .ZN(n10763) );
  NAND2_X1 U17135 ( .A1(n11120), .A2(n11124), .ZN(n10759) );
  AOI21_X1 U17136 ( .B1(n10760), .B2(n10759), .A(n11119), .ZN(n10762) );
  NOR2_X1 U17137 ( .A1(n11124), .A2(n11123), .ZN(n10761) );
  INV_X1 U17138 ( .A(n11848), .ZN(n11641) );
  AOI22_X1 U17139 ( .A1(n10763), .A2(n11515), .B1(n11641), .B2(n11401), .ZN(
        n10764) );
  INV_X1 U17140 ( .A(n10868), .ZN(n11583) );
  NAND2_X1 U17141 ( .A1(n11877), .A2(n11583), .ZN(n10771) );
  INV_X1 U17142 ( .A(n11881), .ZN(n11582) );
  INV_X1 U17143 ( .A(n10766), .ZN(n10769) );
  INV_X1 U17144 ( .A(n10767), .ZN(n10768) );
  NAND4_X1 U17145 ( .A1(n10769), .A2(n11583), .A3(n10768), .A4(n10453), .ZN(
        n10770) );
  XNOR2_X1 U17146 ( .A(n13109), .B(n13547), .ZN(n13237) );
  XNOR2_X1 U17147 ( .A(n13237), .B(n12065), .ZN(n10772) );
  NOR2_X1 U17148 ( .A1(n29648), .A2(n11235), .ZN(n10775) );
  NOR2_X1 U17149 ( .A1(n11012), .A2(n10776), .ZN(n10777) );
  OAI21_X1 U17151 ( .B1(n9362), .B2(n10962), .A(n10958), .ZN(n10781) );
  AND3_X1 U17154 ( .A1(n10980), .A2(n10988), .A3(n589), .ZN(n10784) );
  INV_X1 U17155 ( .A(n10784), .ZN(n12094) );
  MUX2_X1 U17156 ( .A(n10785), .B(n10787), .S(n10786), .Z(n10792) );
  NAND2_X1 U17157 ( .A1(n10791), .A2(n10991), .ZN(n10789) );
  NAND2_X1 U17158 ( .A1(n10787), .A2(n10786), .ZN(n10788) );
  MUX2_X1 U17159 ( .A(n10789), .B(n10788), .S(n3454), .Z(n10790) );
  OAI21_X1 U17160 ( .B1(n10792), .B2(n10791), .A(n10790), .ZN(n11385) );
  INV_X1 U17161 ( .A(n11385), .ZN(n12100) );
  AND2_X1 U17162 ( .A1(n11099), .A2(n333), .ZN(n11893) );
  NAND2_X1 U17163 ( .A1(n6814), .A2(n10795), .ZN(n10796) );
  NAND2_X1 U17164 ( .A1(n11896), .A2(n10797), .ZN(n10798) );
  AOI21_X1 U17165 ( .B1(n12100), .B2(n12155), .A(n12088), .ZN(n10801) );
  NOR2_X1 U17166 ( .A1(n10431), .A2(n11093), .ZN(n10800) );
  OAI21_X1 U17167 ( .B1(n11206), .B2(n587), .A(n11207), .ZN(n10799) );
  MUX2_X1 U17168 ( .A(n10800), .B(n10799), .S(n11094), .Z(n12091) );
  NOR2_X1 U17169 ( .A1(n11205), .A2(n29517), .ZN(n12092) );
  OAI21_X1 U17170 ( .B1(n11146), .B2(n10806), .A(n10805), .ZN(n10807) );
  OAI211_X1 U17171 ( .C1(n10808), .C2(n11149), .A(n11146), .B(n28627), .ZN(
        n10809) );
  AOI22_X1 U17172 ( .A1(n11322), .A2(n11323), .B1(n11321), .B2(n10810), .ZN(
        n10811) );
  NOR2_X1 U17173 ( .A1(n10811), .A2(n11183), .ZN(n10812) );
  NOR3_X1 U17174 ( .A1(n581), .A2(n11198), .A3(n28157), .ZN(n10817) );
  INV_X1 U17175 ( .A(n11646), .ZN(n11645) );
  NAND2_X1 U17176 ( .A1(n11645), .A2(n11715), .ZN(n11414) );
  INV_X1 U17177 ( .A(n10821), .ZN(n11329) );
  OR2_X1 U17178 ( .A1(n10823), .A2(n11331), .ZN(n10824) );
  NOR2_X1 U17179 ( .A1(n11335), .A2(n11176), .ZN(n10826) );
  NOR2_X1 U17180 ( .A1(n11338), .A2(n434), .ZN(n10825) );
  MUX2_X1 U17181 ( .A(n10826), .B(n10825), .S(n11345), .Z(n10832) );
  INV_X1 U17182 ( .A(n10827), .ZN(n11179) );
  NAND3_X1 U17183 ( .A1(n11176), .A2(n11174), .A3(n1898), .ZN(n10829) );
  OAI21_X1 U17184 ( .B1(n11179), .B2(n10830), .A(n10829), .ZN(n10831) );
  XNOR2_X1 U17185 ( .A(n12723), .B(n13386), .ZN(n10867) );
  NAND2_X1 U17186 ( .A1(n586), .A2(n10833), .ZN(n10837) );
  AND2_X1 U17187 ( .A1(n10834), .A2(n11252), .ZN(n11250) );
  INV_X1 U17188 ( .A(n11250), .ZN(n10835) );
  MUX2_X1 U17189 ( .A(n10837), .B(n10836), .S(n29148), .Z(n10841) );
  INV_X1 U17190 ( .A(n10838), .ZN(n10839) );
  NAND2_X1 U17191 ( .A1(n10839), .A2(n11033), .ZN(n10840) );
  NAND2_X1 U17192 ( .A1(n11034), .A2(n279), .ZN(n10843) );
  NAND3_X1 U17193 ( .A1(n10847), .A2(n11350), .A3(n11347), .ZN(n10848) );
  INV_X1 U17194 ( .A(n11347), .ZN(n11191) );
  OAI21_X1 U17195 ( .B1(n11349), .B2(n11348), .A(n10849), .ZN(n10850) );
  NOR2_X1 U17196 ( .A1(n11308), .A2(n10851), .ZN(n10854) );
  INV_X1 U17197 ( .A(n11053), .ZN(n11312) );
  AOI22_X1 U17198 ( .A1(n10854), .A2(n1933), .B1(n10852), .B2(n10851), .ZN(
        n10857) );
  INV_X1 U17199 ( .A(n11321), .ZN(n10858) );
  NAND3_X1 U17200 ( .A1(n11184), .A2(n10858), .A3(n10473), .ZN(n10860) );
  OAI21_X1 U17201 ( .B1(n12037), .B2(n12241), .A(n10861), .ZN(n12239) );
  OAI211_X1 U17203 ( .C1(n3653), .C2(n12507), .A(n12512), .B(n11990), .ZN(
        n10865) );
  XNOR2_X1 U17204 ( .A(n11684), .B(n10867), .ZN(n10904) );
  NAND2_X1 U17205 ( .A1(n11878), .A2(n11877), .ZN(n10870) );
  INV_X1 U17206 ( .A(n13195), .ZN(n12914) );
  NAND2_X1 U17207 ( .A1(n10871), .A2(n435), .ZN(n10874) );
  MUX2_X1 U17209 ( .A(n10874), .B(n28329), .S(n11220), .Z(n11658) );
  INV_X1 U17210 ( .A(n11217), .ZN(n10879) );
  NOR2_X1 U17211 ( .A1(n10876), .A2(n435), .ZN(n10877) );
  AOI22_X1 U17212 ( .A1(n10879), .A2(n10878), .B1(n10877), .B2(n11222), .ZN(
        n11657) );
  AOI21_X1 U17213 ( .B1(n11063), .B2(n11242), .A(n11243), .ZN(n10881) );
  INV_X1 U17214 ( .A(n10882), .ZN(n11083) );
  NAND2_X1 U17215 ( .A1(n1854), .A2(n10884), .ZN(n11028) );
  NAND3_X1 U17216 ( .A1(n11027), .A2(n11284), .A3(n11281), .ZN(n10886) );
  OAI211_X1 U17217 ( .C1(n11283), .C2(n10884), .A(n11029), .B(n584), .ZN(
        n10885) );
  INV_X1 U17218 ( .A(n12164), .ZN(n10887) );
  OAI21_X1 U17219 ( .B1(n1931), .B2(n12163), .A(n10887), .ZN(n10897) );
  AND2_X1 U17220 ( .A1(n11264), .A2(n11267), .ZN(n10890) );
  OAI21_X1 U17221 ( .B1(n10890), .B2(n29510), .A(n10889), .ZN(n11656) );
  MUX2_X1 U17223 ( .A(n11294), .B(n11290), .S(n10318), .Z(n11659) );
  AND2_X1 U17224 ( .A1(n11659), .A2(n29116), .ZN(n10895) );
  XNOR2_X1 U17225 ( .A(n12914), .B(n13556), .ZN(n10902) );
  NOR2_X1 U17226 ( .A1(n12359), .A2(n12362), .ZN(n10900) );
  INV_X1 U17227 ( .A(n12356), .ZN(n11907) );
  XNOR2_X1 U17228 ( .A(n13101), .B(n3742), .ZN(n10901) );
  XNOR2_X1 U17229 ( .A(n10902), .B(n10901), .ZN(n10903) );
  XNOR2_X1 U17230 ( .A(n10904), .B(n10903), .ZN(n14105) );
  NAND2_X1 U17231 ( .A1(n11547), .A2(n11855), .ZN(n10907) );
  MUX2_X1 U17232 ( .A(n10907), .B(n10906), .S(n11549), .Z(n10910) );
  NAND3_X1 U17233 ( .A1(n11137), .A2(n10918), .A3(n10919), .ZN(n10922) );
  NAND2_X1 U17234 ( .A1(n1879), .A2(n10924), .ZN(n10925) );
  AOI21_X1 U17235 ( .B1(n10926), .B2(n10925), .A(n590), .ZN(n10935) );
  NAND2_X1 U17236 ( .A1(n10930), .A2(n10929), .ZN(n10931) );
  NAND2_X1 U17237 ( .A1(n11951), .A2(n11861), .ZN(n10955) );
  NOR2_X1 U17238 ( .A1(n11002), .A2(n592), .ZN(n10938) );
  INV_X1 U17239 ( .A(n11944), .ZN(n11857) );
  OAI22_X1 U17240 ( .A1(n10944), .A2(n10946), .B1(n10943), .B2(n10942), .ZN(
        n10945) );
  NAND2_X1 U17241 ( .A1(n10949), .A2(n28608), .ZN(n10951) );
  NAND3_X1 U17242 ( .A1(n11862), .A2(n11945), .A3(n11943), .ZN(n10953) );
  INV_X1 U17243 ( .A(n11859), .ZN(n11948) );
  NOR2_X1 U17244 ( .A1(n10956), .A2(n10963), .ZN(n10961) );
  NAND2_X1 U17245 ( .A1(n10963), .A2(n10962), .ZN(n10965) );
  NOR2_X1 U17246 ( .A1(n29577), .A2(n10970), .ZN(n10974) );
  OAI21_X1 U17247 ( .B1(n10974), .B2(n10973), .A(n10972), .ZN(n10979) );
  OAI211_X1 U17248 ( .C1(n10983), .C2(n10982), .A(n10981), .B(n10980), .ZN(
        n10987) );
  NAND3_X1 U17249 ( .A1(n10985), .A2(n10988), .A3(n10984), .ZN(n10986) );
  AOI21_X1 U17251 ( .B1(n10999), .B2(n10998), .A(n10997), .ZN(n11009) );
  NOR2_X1 U17252 ( .A1(n5573), .A2(n11000), .ZN(n11001) );
  NOR2_X1 U17253 ( .A1(n11001), .A2(n28405), .ZN(n11008) );
  NAND2_X1 U17254 ( .A1(n11005), .A2(n28405), .ZN(n11006) );
  NOR2_X1 U17255 ( .A1(n3441), .A2(n11010), .ZN(n11011) );
  NAND2_X1 U17256 ( .A1(n11237), .A2(n11011), .ZN(n11018) );
  NAND3_X1 U17257 ( .A1(n5709), .A2(n11236), .A3(n11014), .ZN(n11015) );
  NOR2_X1 U17258 ( .A1(n12252), .A2(n12253), .ZN(n11019) );
  AOI22_X1 U17259 ( .A1(n11020), .A2(n12070), .B1(n11019), .B2(n349), .ZN(
        n11021) );
  AND2_X1 U17260 ( .A1(n11022), .A2(n11315), .ZN(n11319) );
  NAND2_X1 U17261 ( .A1(n11319), .A2(n11258), .ZN(n11025) );
  NAND4_X1 U17262 ( .A1(n11317), .A2(n11025), .A3(n11024), .A4(n11023), .ZN(
        n12263) );
  INV_X1 U17263 ( .A(n12263), .ZN(n12133) );
  NAND2_X1 U17264 ( .A1(n11282), .A2(n11281), .ZN(n11026) );
  INV_X1 U17266 ( .A(n11028), .ZN(n11031) );
  NOR2_X1 U17267 ( .A1(n11280), .A2(n11029), .ZN(n11030) );
  OAI21_X1 U17268 ( .B1(n12133), .B2(n11435), .A(n12132), .ZN(n11062) );
  NAND2_X1 U17269 ( .A1(n11273), .A2(n28612), .ZN(n11036) );
  MUX2_X1 U17271 ( .A(n11036), .B(n11035), .S(n28147), .Z(n11042) );
  NAND2_X1 U17272 ( .A1(n12133), .A2(n11574), .ZN(n11928) );
  INV_X1 U17273 ( .A(n11928), .ZN(n11061) );
  AOI21_X1 U17274 ( .B1(n11045), .B2(n11266), .A(n11267), .ZN(n11046) );
  NAND2_X1 U17275 ( .A1(n11262), .A2(n11046), .ZN(n11050) );
  NAND3_X1 U17276 ( .A1(n11048), .A2(n11047), .A3(n11266), .ZN(n11049) );
  NAND2_X1 U17277 ( .A1(n10855), .A2(n11165), .ZN(n11052) );
  NAND2_X1 U17278 ( .A1(n11164), .A2(n11053), .ZN(n11054) );
  OAI211_X1 U17279 ( .C1(n11057), .C2(n29637), .A(n11055), .B(n11054), .ZN(
        n12264) );
  NAND3_X1 U17280 ( .A1(n12134), .A2(n11574), .A3(n12267), .ZN(n11059) );
  XNOR2_X1 U17281 ( .A(n12827), .B(n13371), .ZN(n12466) );
  XNOR2_X1 U17282 ( .A(n12087), .B(n12466), .ZN(n11203) );
  NOR2_X1 U17283 ( .A1(n1900), .A2(n11063), .ZN(n11065) );
  NAND2_X1 U17284 ( .A1(n1900), .A2(n11066), .ZN(n11241) );
  OAI22_X1 U17285 ( .A1(n11069), .A2(n11241), .B1(n11068), .B2(n11240), .ZN(
        n11070) );
  INV_X1 U17286 ( .A(n11290), .ZN(n11071) );
  NAND2_X1 U17287 ( .A1(n11071), .A2(n10665), .ZN(n11080) );
  OAI21_X1 U17288 ( .B1(n11075), .B2(n11072), .A(n10665), .ZN(n11074) );
  OAI21_X1 U17289 ( .B1(n11291), .B2(n11287), .A(n29116), .ZN(n11073) );
  NAND2_X1 U17290 ( .A1(n11074), .A2(n11073), .ZN(n11079) );
  NAND3_X1 U17291 ( .A1(n11077), .A2(n11076), .A3(n11075), .ZN(n11078) );
  INV_X1 U17292 ( .A(n12270), .ZN(n12576) );
  NAND2_X1 U17293 ( .A1(n11213), .A2(n28624), .ZN(n11081) );
  NOR2_X1 U17294 ( .A1(n11084), .A2(n11083), .ZN(n11088) );
  NOR2_X1 U17295 ( .A1(n11086), .A2(n11085), .ZN(n11087) );
  MUX2_X1 U17296 ( .A(n11088), .B(n11087), .S(n11210), .Z(n11089) );
  NAND2_X1 U17297 ( .A1(n11207), .A2(n10431), .ZN(n11091) );
  AOI21_X1 U17298 ( .B1(n11092), .B2(n11091), .A(n11090), .ZN(n11098) );
  NAND2_X1 U17299 ( .A1(n29517), .A2(n11093), .ZN(n11096) );
  OAI21_X1 U17300 ( .B1(n5277), .B2(n11096), .A(n11095), .ZN(n11097) );
  NOR2_X1 U17301 ( .A1(n12578), .A2(n12517), .ZN(n12273) );
  OAI21_X1 U17302 ( .B1(n11099), .B2(n333), .A(n11225), .ZN(n11100) );
  NAND2_X1 U17303 ( .A1(n11100), .A2(n9709), .ZN(n11102) );
  INV_X1 U17304 ( .A(n11898), .ZN(n11101) );
  INV_X1 U17305 ( .A(n12516), .ZN(n11940) );
  MUX2_X1 U17306 ( .A(n11103), .B(n12273), .S(n11940), .Z(n11110) );
  NOR2_X1 U17307 ( .A1(n11222), .A2(n435), .ZN(n11107) );
  NAND2_X1 U17308 ( .A1(n11104), .A2(n11220), .ZN(n11105) );
  OAI21_X1 U17309 ( .B1(n5974), .B2(n28202), .A(n12578), .ZN(n11108) );
  NOR2_X1 U17310 ( .A1(n11121), .A2(n11120), .ZN(n11130) );
  NAND3_X1 U17311 ( .A1(n11124), .A2(n11123), .A3(n11122), .ZN(n11129) );
  NAND3_X1 U17312 ( .A1(n11127), .A2(n11126), .A3(n11125), .ZN(n11128) );
  NAND2_X1 U17313 ( .A1(n11774), .A2(n11131), .ZN(n11134) );
  NAND3_X1 U17314 ( .A1(n11133), .A2(n11132), .A3(n4555), .ZN(n11775) );
  INV_X1 U17315 ( .A(n11551), .ZN(n11422) );
  NAND2_X1 U17316 ( .A1(n11422), .A2(n11782), .ZN(n11151) );
  AOI22_X1 U17317 ( .A1(n11137), .A2(n11136), .B1(n11135), .B2(n3862), .ZN(
        n11143) );
  NAND2_X1 U17319 ( .A1(n11421), .A2(n11553), .ZN(n11150) );
  OAI21_X1 U17320 ( .B1(n11146), .B2(n28627), .A(n11144), .ZN(n11147) );
  MUX2_X1 U17321 ( .A(n11151), .B(n11150), .S(n11785), .Z(n11161) );
  NAND2_X1 U17322 ( .A1(n28175), .A2(n11153), .ZN(n11156) );
  INV_X1 U17323 ( .A(n11154), .ZN(n11155) );
  XNOR2_X1 U17324 ( .A(n13249), .B(n1905), .ZN(n13532) );
  NAND2_X1 U17325 ( .A1(n11166), .A2(n11168), .ZN(n11167) );
  OAI211_X1 U17326 ( .C1(n11169), .C2(n11168), .A(n11167), .B(n11330), .ZN(
        n11172) );
  NAND3_X1 U17327 ( .A1(n28208), .A2(n11331), .A3(n11170), .ZN(n11171) );
  NAND3_X1 U17331 ( .A1(n11349), .A2(n11192), .A3(n11350), .ZN(n11193) );
  XNOR2_X1 U17332 ( .A(n13118), .B(n3378), .ZN(n11201) );
  XNOR2_X1 U17333 ( .A(n13532), .B(n11201), .ZN(n11202) );
  OAI211_X1 U17334 ( .C1(n11211), .C2(n28624), .A(n433), .B(n11209), .ZN(
        n11215) );
  OAI21_X1 U17335 ( .B1(n11222), .B2(n11218), .A(n11217), .ZN(n11224) );
  OAI21_X1 U17336 ( .B1(n11223), .B2(n11220), .A(n11219), .ZN(n11221) );
  OAI21_X1 U17337 ( .B1(n333), .B2(n11225), .A(n11231), .ZN(n11229) );
  NAND2_X1 U17338 ( .A1(n11232), .A2(n28270), .ZN(n11228) );
  AND2_X1 U17342 ( .A1(n12315), .A2(n12321), .ZN(n11246) );
  NOR2_X1 U17343 ( .A1(n11243), .A2(n11242), .ZN(n11245) );
  NAND2_X1 U17344 ( .A1(n11254), .A2(n11315), .ZN(n11256) );
  MUX2_X1 U17345 ( .A(n11256), .B(n11314), .S(n11255), .Z(n11257) );
  OAI21_X1 U17346 ( .B1(n11259), .B2(n11258), .A(n11257), .ZN(n12081) );
  NOR2_X1 U17347 ( .A1(n12080), .A2(n12081), .ZN(n11297) );
  NAND2_X1 U17348 ( .A1(n11264), .A2(n28204), .ZN(n11265) );
  NAND3_X1 U17349 ( .A1(n28174), .A2(n11267), .A3(n11266), .ZN(n12290) );
  NAND2_X1 U17350 ( .A1(n12289), .A2(n12081), .ZN(n12062) );
  OAI21_X1 U17351 ( .B1(n11271), .B2(n10523), .A(n11270), .ZN(n11279) );
  NAND2_X1 U17352 ( .A1(n10523), .A2(n11272), .ZN(n11277) );
  AOI21_X1 U17353 ( .B1(n11277), .B2(n11276), .A(n11275), .ZN(n11278) );
  NOR2_X1 U17354 ( .A1(n11288), .A2(n11287), .ZN(n11289) );
  MUX2_X1 U17355 ( .A(n12062), .B(n11295), .S(n29324), .Z(n11296) );
  XNOR2_X1 U17356 ( .A(n13539), .B(n12841), .ZN(n11307) );
  NAND2_X1 U17357 ( .A1(n11782), .A2(n11785), .ZN(n11301) );
  OR2_X1 U17358 ( .A1(n11552), .A2(n11785), .ZN(n11300) );
  INV_X1 U17359 ( .A(n11782), .ZN(n11298) );
  OAI211_X1 U17360 ( .C1(n11551), .C2(n29137), .A(n11552), .B(n11298), .ZN(
        n11299) );
  OAI211_X1 U17361 ( .C1(n11550), .C2(n11301), .A(n11300), .B(n11299), .ZN(
        n12931) );
  NAND2_X1 U17362 ( .A1(n11789), .A2(n28436), .ZN(n11305) );
  NAND3_X1 U17363 ( .A1(n10717), .A2(n2194), .A3(n2748), .ZN(n11304) );
  NAND2_X1 U17364 ( .A1(n10717), .A2(n11302), .ZN(n11303) );
  XNOR2_X1 U17365 ( .A(n12931), .B(n13075), .ZN(n12136) );
  XNOR2_X1 U17366 ( .A(n11307), .B(n12136), .ZN(n11370) );
  NOR2_X1 U17367 ( .A1(n11315), .A2(n11314), .ZN(n11320) );
  NOR2_X1 U17370 ( .A1(n11330), .A2(n11329), .ZN(n11333) );
  INV_X1 U17371 ( .A(n12402), .ZN(n11346) );
  NAND2_X1 U17372 ( .A1(n11335), .A2(n11334), .ZN(n11344) );
  NOR2_X1 U17373 ( .A1(n11341), .A2(n11337), .ZN(n11339) );
  AOI22_X1 U17374 ( .A1(n11339), .A2(n11338), .B1(n11337), .B2(n11336), .ZN(
        n11343) );
  OAI21_X1 U17375 ( .B1(n11346), .B2(n12281), .A(n12286), .ZN(n11357) );
  NAND3_X1 U17377 ( .A1(n11352), .A2(n11351), .A3(n11350), .ZN(n11353) );
  OAI211_X2 U17378 ( .C1(n11356), .C2(n11355), .A(n11354), .B(n11353), .ZN(
        n12407) );
  OAI211_X1 U17381 ( .C1(n11868), .C2(n11500), .A(n11457), .B(n578), .ZN(
        n11361) );
  INV_X1 U17382 ( .A(n12303), .ZN(n11769) );
  OAI21_X1 U17385 ( .B1(n569), .B2(n12300), .A(n12305), .ZN(n11365) );
  INV_X1 U17386 ( .A(n11363), .ZN(n11364) );
  AOI22_X2 U17387 ( .A1(n11366), .A2(n11365), .B1(n11364), .B2(n12300), .ZN(
        n13404) );
  XNOR2_X1 U17388 ( .A(n13404), .B(n3164), .ZN(n11367) );
  XNOR2_X1 U17389 ( .A(n11368), .B(n11367), .ZN(n11369) );
  NOR2_X1 U17390 ( .A1(n12111), .A2(n12110), .ZN(n11831) );
  OAI21_X1 U17391 ( .B1(n12207), .B2(n12208), .A(n28203), .ZN(n11375) );
  NOR2_X1 U17392 ( .A1(n12110), .A2(n9692), .ZN(n11374) );
  INV_X1 U17394 ( .A(n12171), .ZN(n11382) );
  INV_X1 U17395 ( .A(n11656), .ZN(n12103) );
  NAND2_X1 U17396 ( .A1(n12103), .A2(n12164), .ZN(n11376) );
  INV_X1 U17397 ( .A(n12163), .ZN(n11378) );
  XNOR2_X1 U17398 ( .A(n13297), .B(n13401), .ZN(n12490) );
  NOR2_X1 U17399 ( .A1(n12151), .A2(n579), .ZN(n11384) );
  NOR2_X1 U17400 ( .A1(n11856), .A2(n12088), .ZN(n11383) );
  NOR3_X1 U17401 ( .A1(n11384), .A2(n12150), .A3(n11383), .ZN(n11388) );
  AND2_X1 U17402 ( .A1(n12151), .A2(n11856), .ZN(n12152) );
  NAND2_X1 U17403 ( .A1(n12152), .A2(n12990), .ZN(n11386) );
  NAND2_X1 U17404 ( .A1(n11927), .A2(n11851), .ZN(n11394) );
  OAI21_X1 U17405 ( .B1(n11853), .B2(n11855), .A(n11852), .ZN(n11392) );
  NAND3_X1 U17407 ( .A1(n11944), .A2(n11858), .A3(n11945), .ZN(n11397) );
  NAND2_X1 U17408 ( .A1(n11952), .A2(n11947), .ZN(n11395) );
  NAND2_X1 U17409 ( .A1(n11397), .A2(n11396), .ZN(n11400) );
  NAND2_X1 U17410 ( .A1(n11857), .A2(n11948), .ZN(n11398) );
  AOI21_X1 U17411 ( .B1(n11665), .B2(n11398), .A(n11862), .ZN(n11399) );
  NOR2_X2 U17412 ( .A1(n11400), .A2(n11399), .ZN(n13208) );
  XNOR2_X1 U17413 ( .A(n13025), .B(n13208), .ZN(n12930) );
  NOR2_X1 U17414 ( .A1(n11402), .A2(n11848), .ZN(n11407) );
  INV_X1 U17415 ( .A(n11672), .ZN(n11404) );
  NOR3_X1 U17416 ( .A1(n11405), .A2(n11404), .A3(n11403), .ZN(n11406) );
  XNOR2_X1 U17417 ( .A(n12747), .B(n13405), .ZN(n11409) );
  XNOR2_X1 U17418 ( .A(n12930), .B(n11409), .ZN(n11410) );
  INV_X1 U17419 ( .A(n12176), .ZN(n12124) );
  INV_X1 U17420 ( .A(n11824), .ZN(n12180) );
  AOI22_X1 U17421 ( .A1(n11730), .A2(n12125), .B1(n12124), .B2(n12180), .ZN(
        n11413) );
  MUX2_X1 U17422 ( .A(n11411), .B(n12124), .S(n11730), .Z(n11412) );
  XNOR2_X1 U17423 ( .A(n12788), .B(n12595), .ZN(n11432) );
  INV_X1 U17424 ( .A(n11419), .ZN(n11502) );
  AOI21_X1 U17425 ( .B1(n11422), .B2(n11778), .A(n11421), .ZN(n11423) );
  INV_X1 U17426 ( .A(n11426), .ZN(n11427) );
  NOR2_X1 U17427 ( .A1(n11427), .A2(n11430), .ZN(n11429) );
  NAND3_X1 U17429 ( .A1(n12128), .A2(n12189), .A3(n11818), .ZN(n11434) );
  INV_X1 U17430 ( .A(n12189), .ZN(n11724) );
  OAI211_X2 U17431 ( .C1(n11727), .C2(n11816), .A(n11434), .B(n11433), .ZN(
        n13230) );
  AOI22_X1 U17432 ( .A1(n12132), .A2(n11058), .B1(n12264), .B2(n12263), .ZN(
        n11930) );
  NAND2_X1 U17433 ( .A1(n575), .A2(n12263), .ZN(n11436) );
  NAND2_X1 U17434 ( .A1(n11436), .A2(n12264), .ZN(n11437) );
  XNOR2_X1 U17435 ( .A(n13230), .B(n13380), .ZN(n11443) );
  NAND2_X1 U17436 ( .A1(n12200), .A2(n12203), .ZN(n11441) );
  OAI211_X1 U17437 ( .C1(n12204), .C2(n11441), .A(n11440), .B(n11439), .ZN(
        n12948) );
  XNOR2_X1 U17438 ( .A(n12948), .B(n3334), .ZN(n11442) );
  XNOR2_X1 U17439 ( .A(n11443), .B(n11442), .ZN(n11444) );
  XNOR2_X2 U17440 ( .A(n11445), .B(n11444), .ZN(n15194) );
  INV_X1 U17441 ( .A(n11740), .ZN(n12357) );
  OAI21_X1 U17442 ( .B1(n12363), .B2(n12362), .A(n11446), .ZN(n11447) );
  NAND3_X1 U17443 ( .A1(n12327), .A2(n12018), .A3(n11449), .ZN(n11452) );
  INV_X1 U17444 ( .A(n11747), .ZN(n12329) );
  OAI211_X1 U17445 ( .C1(n11888), .C2(n12328), .A(n11450), .B(n12332), .ZN(
        n11451) );
  XNOR2_X1 U17447 ( .A(n13166), .B(n13278), .ZN(n11466) );
  NAND2_X1 U17448 ( .A1(n11875), .A2(n11877), .ZN(n11454) );
  AOI22_X1 U17449 ( .A1(n130), .A2(n11454), .B1(n287), .B2(n11453), .ZN(n11456) );
  NAND3_X1 U17450 ( .A1(n11881), .A2(n11877), .A3(n11876), .ZN(n11455) );
  NOR2_X1 U17452 ( .A1(n4712), .A2(n11458), .ZN(n11459) );
  OAI211_X1 U17453 ( .C1(n1836), .C2(n11869), .A(n11462), .B(n11500), .ZN(
        n11464) );
  XNOR2_X1 U17454 ( .A(n12894), .B(n12817), .ZN(n11465) );
  XNOR2_X1 U17455 ( .A(n11465), .B(n11466), .ZN(n11481) );
  INV_X1 U17456 ( .A(n12352), .ZN(n11467) );
  NAND3_X1 U17458 ( .A1(n29209), .A2(n12353), .A3(n29735), .ZN(n11470) );
  NAND2_X1 U17459 ( .A1(n12339), .A2(n12337), .ZN(n11474) );
  XNOR2_X1 U17460 ( .A(n13018), .B(n12514), .ZN(n12681) );
  INV_X1 U17461 ( .A(n11755), .ZN(n11996) );
  AND2_X1 U17462 ( .A1(n11754), .A2(n12000), .ZN(n11995) );
  NAND3_X1 U17463 ( .A1(n11998), .A2(n11754), .A3(n11755), .ZN(n11476) );
  OAI211_X1 U17464 ( .C1(n11995), .C2(n11755), .A(n11477), .B(n11476), .ZN(
        n11478) );
  XNOR2_X1 U17466 ( .A(n12763), .B(n26531), .ZN(n11479) );
  XNOR2_X1 U17467 ( .A(n12681), .B(n11479), .ZN(n11480) );
  INV_X1 U17468 ( .A(n12081), .ZN(n12291) );
  NAND2_X1 U17469 ( .A1(n29498), .A2(n11795), .ZN(n12296) );
  NOR2_X1 U17470 ( .A1(n12058), .A2(n29499), .ZN(n11796) );
  INV_X1 U17471 ( .A(n12289), .ZN(n11482) );
  NOR2_X1 U17473 ( .A1(n12053), .A2(n12313), .ZN(n12312) );
  INV_X1 U17474 ( .A(n12312), .ZN(n11485) );
  NOR2_X1 U17475 ( .A1(n12315), .A2(n12049), .ZN(n11484) );
  INV_X1 U17476 ( .A(n12320), .ZN(n12054) );
  NAND2_X1 U17477 ( .A1(n12054), .A2(n12313), .ZN(n11613) );
  OR2_X1 U17478 ( .A1(n11613), .A2(n12049), .ZN(n11483) );
  NAND3_X1 U17480 ( .A1(n11793), .A2(n2194), .A3(n4046), .ZN(n11488) );
  INV_X1 U17481 ( .A(n13263), .ZN(n11498) );
  AND3_X1 U17482 ( .A1(n11769), .A2(n12304), .A3(n11768), .ZN(n11496) );
  NOR2_X2 U17483 ( .A1(n11497), .A2(n11496), .ZN(n13104) );
  XNOR2_X1 U17484 ( .A(n11498), .B(n13104), .ZN(n12912) );
  INV_X1 U17485 ( .A(n12912), .ZN(n11499) );
  XNOR2_X1 U17486 ( .A(n11499), .B(n12966), .ZN(n11511) );
  OAI211_X1 U17487 ( .C1(n3900), .C2(n11502), .A(n11551), .B(n11553), .ZN(
        n11503) );
  INV_X1 U17488 ( .A(n12722), .ZN(n11937) );
  XNOR2_X1 U17489 ( .A(n11937), .B(n12965), .ZN(n11509) );
  OR2_X1 U17490 ( .A1(n12402), .A2(n12407), .ZN(n11507) );
  NAND2_X1 U17491 ( .A1(n11801), .A2(n12400), .ZN(n12283) );
  NAND3_X1 U17492 ( .A1(n12280), .A2(n12402), .A3(n12281), .ZN(n11506) );
  XNOR2_X1 U17493 ( .A(n13150), .B(n3223), .ZN(n11508) );
  XNOR2_X1 U17494 ( .A(n11509), .B(n11508), .ZN(n11510) );
  INV_X1 U17495 ( .A(n14241), .ZN(n14243) );
  NAND3_X1 U17496 ( .A1(n11970), .A2(n12159), .A3(n12037), .ZN(n11513) );
  INV_X1 U17497 ( .A(n11673), .ZN(n11639) );
  NAND3_X1 U17499 ( .A1(n11848), .A2(n29139), .A3(n11640), .ZN(n11516) );
  XNOR2_X1 U17500 ( .A(n12780), .B(n13137), .ZN(n13375) );
  NOR2_X1 U17501 ( .A1(n3653), .A2(n12508), .ZN(n11836) );
  NAND3_X1 U17502 ( .A1(n12512), .A2(n6374), .A3(n10863), .ZN(n11520) );
  INV_X1 U17503 ( .A(n13081), .ZN(n13084) );
  INV_X1 U17504 ( .A(n303), .ZN(n11522) );
  NAND3_X1 U17505 ( .A1(n13083), .A2(n13084), .A3(n11522), .ZN(n11531) );
  AND2_X1 U17506 ( .A1(n11524), .A2(n11523), .ZN(n11527) );
  NAND4_X1 U17507 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11529) );
  XNOR2_X1 U17508 ( .A(n13270), .B(n13533), .ZN(n12905) );
  XNOR2_X1 U17509 ( .A(n13375), .B(n12905), .ZN(n11546) );
  INV_X1 U17510 ( .A(n12220), .ZN(n11963) );
  INV_X1 U17511 ( .A(n12219), .ZN(n11965) );
  NAND2_X1 U17512 ( .A1(n12043), .A2(n11965), .ZN(n11534) );
  NAND2_X1 U17513 ( .A1(n12044), .A2(n11963), .ZN(n11533) );
  NAND3_X1 U17514 ( .A1(n12220), .A2(n12219), .A3(n12218), .ZN(n11532) );
  NAND4_X2 U17515 ( .A1(n11535), .A2(n11533), .A3(n11534), .A4(n11532), .ZN(
        n13420) );
  OAI21_X1 U17516 ( .B1(n11754), .B2(n11536), .A(n12000), .ZN(n11537) );
  INV_X1 U17517 ( .A(n11998), .ZN(n12001) );
  NAND3_X1 U17518 ( .A1(n12001), .A2(n11754), .A3(n11996), .ZN(n11539) );
  XNOR2_X1 U17519 ( .A(n12830), .B(n13420), .ZN(n11544) );
  NAND3_X1 U17520 ( .A1(n1986), .A2(n12236), .A3(n375), .ZN(n11542) );
  XNOR2_X1 U17521 ( .A(n11544), .B(n11543), .ZN(n11545) );
  INV_X1 U17522 ( .A(n14171), .ZN(n14239) );
  INV_X1 U17524 ( .A(n11861), .ZN(n11558) );
  NOR2_X1 U17525 ( .A1(n11952), .A2(n11947), .ZN(n11555) );
  AOI22_X1 U17526 ( .A1(n11951), .A2(n11555), .B1(n11944), .B2(n11858), .ZN(
        n11557) );
  INV_X1 U17527 ( .A(n11947), .ZN(n11556) );
  AOI21_X1 U17528 ( .B1(n349), .B2(n12249), .A(n12070), .ZN(n11559) );
  NAND2_X1 U17529 ( .A1(n11559), .A2(n11934), .ZN(n11562) );
  NAND2_X1 U17530 ( .A1(n11594), .A2(n12070), .ZN(n11561) );
  INV_X1 U17531 ( .A(n12253), .ZN(n11932) );
  NOR2_X1 U17532 ( .A1(n349), .A2(n11932), .ZN(n11560) );
  XNOR2_X1 U17533 ( .A(n13364), .B(n13190), .ZN(n12920) );
  XNOR2_X1 U17534 ( .A(n11563), .B(n12920), .ZN(n11578) );
  NOR2_X1 U17535 ( .A1(n12271), .A2(n12270), .ZN(n12583) );
  INV_X1 U17536 ( .A(n12583), .ZN(n11565) );
  INV_X1 U17537 ( .A(n28202), .ZN(n11564) );
  NAND3_X1 U17538 ( .A1(n12271), .A2(n12517), .A3(n11564), .ZN(n12519) );
  AND2_X1 U17539 ( .A1(n11565), .A2(n12519), .ZN(n11566) );
  INV_X1 U17540 ( .A(n11622), .ZN(n11953) );
  OAI21_X1 U17541 ( .B1(n571), .B2(n11953), .A(n6706), .ZN(n11569) );
  AOI21_X1 U17543 ( .B1(n11574), .B2(n12266), .A(n12267), .ZN(n11571) );
  OAI21_X1 U17544 ( .B1(n12265), .B2(n12266), .A(n11571), .ZN(n11573) );
  NAND3_X1 U17545 ( .A1(n11574), .A2(n568), .A3(n12263), .ZN(n11572) );
  INV_X1 U17546 ( .A(n2402), .ZN(n27678) );
  XNOR2_X1 U17547 ( .A(n13291), .B(n27678), .ZN(n11575) );
  XNOR2_X1 U17548 ( .A(n11578), .B(n11577), .ZN(n14238) );
  NAND3_X1 U17549 ( .A1(n28172), .A2(n14239), .A3(n563), .ZN(n11579) );
  NAND2_X1 U17550 ( .A1(n14893), .A2(n15415), .ZN(n15412) );
  INV_X1 U17551 ( .A(n15412), .ZN(n12012) );
  XNOR2_X1 U17552 ( .A(n12881), .B(n12841), .ZN(n13540) );
  NOR2_X1 U17553 ( .A1(n11881), .A2(n11877), .ZN(n11589) );
  OAI21_X1 U17554 ( .B1(n11878), .B2(n11582), .A(n11876), .ZN(n11588) );
  NOR2_X1 U17555 ( .A1(n11877), .A2(n11583), .ZN(n11584) );
  NOR2_X1 U17556 ( .A1(n10453), .A2(n11876), .ZN(n11585) );
  NAND2_X1 U17557 ( .A1(n287), .A2(n11585), .ZN(n11586) );
  XNOR2_X1 U17559 ( .A(n13540), .B(n12349), .ZN(n11606) );
  NAND2_X1 U17560 ( .A1(n12583), .A2(n11940), .ZN(n12581) );
  NAND2_X1 U17561 ( .A1(n28202), .A2(n12270), .ZN(n11590) );
  NAND2_X1 U17562 ( .A1(n12575), .A2(n11590), .ZN(n11591) );
  INV_X1 U17563 ( .A(n12251), .ZN(n12256) );
  NOR2_X1 U17564 ( .A1(n12253), .A2(n12249), .ZN(n11593) );
  AOI21_X1 U17565 ( .B1(n349), .B2(n12253), .A(n11593), .ZN(n11598) );
  NAND2_X1 U17566 ( .A1(n11595), .A2(n12256), .ZN(n11596) );
  XNOR2_X1 U17567 ( .A(n13504), .B(n13458), .ZN(n12933) );
  NAND2_X1 U17568 ( .A1(n12204), .A2(n4844), .ZN(n11600) );
  AOI21_X1 U17569 ( .B1(n11601), .B2(n11600), .A(n11702), .ZN(n11603) );
  NOR2_X1 U17570 ( .A1(n12205), .A2(n11807), .ZN(n11602) );
  XNOR2_X1 U17571 ( .A(n12933), .B(n11604), .ZN(n11605) );
  XNOR2_X1 U17572 ( .A(n11606), .B(n11605), .ZN(n14157) );
  INV_X1 U17573 ( .A(n14157), .ZN(n13935) );
  NOR2_X1 U17574 ( .A1(n12303), .A2(n12302), .ZN(n11607) );
  NOR2_X1 U17575 ( .A1(n12305), .A2(n11607), .ZN(n11611) );
  INV_X1 U17576 ( .A(n11608), .ZN(n11609) );
  INV_X1 U17577 ( .A(n12548), .ZN(n13473) );
  NAND2_X1 U17578 ( .A1(n285), .A2(n12313), .ZN(n11614) );
  AOI21_X1 U17579 ( .B1(n11614), .B2(n12054), .A(n12316), .ZN(n11615) );
  XNOR2_X1 U17580 ( .A(n13473), .B(n13450), .ZN(n12899) );
  OAI21_X1 U17581 ( .B1(n11617), .B2(n11616), .A(n3653), .ZN(n11620) );
  NOR2_X1 U17582 ( .A1(n12512), .A2(n12508), .ZN(n11618) );
  XNOR2_X1 U17583 ( .A(n13563), .B(n13055), .ZN(n11621) );
  XNOR2_X1 U17584 ( .A(n12899), .B(n11621), .ZN(n11631) );
  INV_X1 U17585 ( .A(n11800), .ZN(n11623) );
  NAND2_X1 U17586 ( .A1(n11623), .A2(n12286), .ZN(n11624) );
  XNOR2_X1 U17587 ( .A(n13567), .B(n3372), .ZN(n11628) );
  XNOR2_X1 U17588 ( .A(n11629), .B(n11628), .ZN(n11630) );
  XNOR2_X2 U17589 ( .A(n11631), .B(n11630), .ZN(n14480) );
  INV_X1 U17590 ( .A(n11632), .ZN(n11638) );
  INV_X1 U17591 ( .A(n11633), .ZN(n11635) );
  NAND2_X1 U17592 ( .A1(n11635), .A2(n11634), .ZN(n11637) );
  NOR3_X1 U17593 ( .A1(n11638), .A2(n11637), .A3(n11636), .ZN(n11675) );
  MUX2_X1 U17594 ( .A(n11675), .B(n11640), .S(n11671), .Z(n11644) );
  NOR2_X1 U17595 ( .A1(n11640), .A2(n11672), .ZN(n11849) );
  NOR2_X1 U17596 ( .A1(n11849), .A2(n29139), .ZN(n11643) );
  NAND3_X1 U17597 ( .A1(n11641), .A2(n11640), .A3(n11639), .ZN(n11642) );
  XNOR2_X1 U17599 ( .A(n29140), .B(n13219), .ZN(n11652) );
  XNOR2_X1 U17600 ( .A(n12867), .B(n13523), .ZN(n13168) );
  XNOR2_X1 U17601 ( .A(n11652), .B(n13168), .ZN(n11670) );
  NOR2_X1 U17602 ( .A1(n12150), .A2(n12100), .ZN(n11653) );
  NAND2_X1 U17603 ( .A1(n1931), .A2(n12164), .ZN(n11654) );
  AOI21_X1 U17605 ( .B1(n11655), .B2(n11654), .A(n28828), .ZN(n11664) );
  INV_X1 U17607 ( .A(n11660), .ZN(n11661) );
  MUX2_X1 U17608 ( .A(n11844), .B(n11662), .S(n12102), .Z(n11663) );
  MUX2_X1 U17609 ( .A(n11951), .B(n11948), .S(n11945), .Z(n11666) );
  XNOR2_X1 U17610 ( .A(n13048), .B(n2274), .ZN(n11669) );
  NOR2_X1 U17612 ( .A1(n11676), .A2(n11675), .ZN(n11679) );
  INV_X1 U17613 ( .A(n11680), .ZN(n11683) );
  OAI21_X2 U17614 ( .B1(n11682), .B2(n11683), .A(n11681), .ZN(n13245) );
  XNOR2_X1 U17615 ( .A(n13553), .B(n13245), .ZN(n12911) );
  XNOR2_X1 U17616 ( .A(n11684), .B(n12911), .ZN(n11701) );
  NOR2_X1 U17617 ( .A1(n12000), .A2(n6661), .ZN(n11757) );
  AND2_X1 U17619 ( .A1(n13081), .A2(n12231), .ZN(n11811) );
  INV_X1 U17620 ( .A(n11811), .ZN(n11689) );
  AND2_X1 U17621 ( .A1(n11980), .A2(n12226), .ZN(n12228) );
  OAI211_X1 U17622 ( .C1(n13081), .C2(n13086), .A(n13083), .B(n11809), .ZN(
        n11690) );
  INV_X1 U17623 ( .A(n13043), .ZN(n11692) );
  XNOR2_X1 U17624 ( .A(n12686), .B(n11692), .ZN(n11699) );
  OAI211_X1 U17625 ( .C1(n12219), .C2(n12218), .A(n12224), .B(n12042), .ZN(
        n11696) );
  NAND4_X1 U17626 ( .A1(n2846), .A2(n12221), .A3(n11694), .A4(n11693), .ZN(
        n11695) );
  XNOR2_X1 U17627 ( .A(n13484), .B(n3422), .ZN(n11698) );
  XNOR2_X1 U17628 ( .A(n11699), .B(n11698), .ZN(n11700) );
  XNOR2_X1 U17629 ( .A(n11701), .B(n11700), .ZN(n13755) );
  INV_X1 U17630 ( .A(n13755), .ZN(n13934) );
  NOR2_X1 U17631 ( .A1(n12202), .A2(n12201), .ZN(n11706) );
  NAND2_X1 U17632 ( .A1(n12204), .A2(n11706), .ZN(n11707) );
  XNOR2_X1 U17633 ( .A(n12495), .B(n12827), .ZN(n13535) );
  INV_X1 U17634 ( .A(n13535), .ZN(n11717) );
  OAI211_X1 U17635 ( .C1(n11712), .C2(n11711), .A(n11710), .B(n11709), .ZN(
        n11713) );
  XNOR2_X1 U17636 ( .A(n1857), .B(n3369), .ZN(n11716) );
  XNOR2_X1 U17637 ( .A(n11717), .B(n11716), .ZN(n11735) );
  INV_X1 U17638 ( .A(n11718), .ZN(n11720) );
  NOR2_X1 U17639 ( .A1(n11787), .A2(n2748), .ZN(n11719) );
  XNOR2_X1 U17640 ( .A(n13249), .B(n13067), .ZN(n12298) );
  NAND3_X1 U17641 ( .A1(n11819), .A2(n12198), .A3(n12186), .ZN(n11722) );
  NOR2_X1 U17642 ( .A1(n12186), .A2(n11724), .ZN(n11725) );
  NAND2_X1 U17643 ( .A1(n2483), .A2(n11725), .ZN(n11726) );
  OAI211_X1 U17644 ( .C1(n11727), .C2(n2483), .A(n6917), .B(n11726), .ZN(
        n12554) );
  INV_X1 U17645 ( .A(n12554), .ZN(n12826) );
  INV_X1 U17646 ( .A(n11730), .ZN(n12179) );
  NOR2_X1 U17647 ( .A1(n12179), .A2(n11824), .ZN(n11729) );
  NOR2_X1 U17648 ( .A1(n12125), .A2(n12124), .ZN(n11728) );
  MUX2_X1 U17649 ( .A(n11729), .B(n11728), .S(n570), .Z(n11733) );
  NAND2_X1 U17650 ( .A1(n1890), .A2(n12177), .ZN(n12183) );
  NOR2_X1 U17651 ( .A1(n13206), .A2(n11731), .ZN(n11732) );
  NOR2_X2 U17652 ( .A1(n11733), .A2(n11732), .ZN(n13418) );
  XNOR2_X1 U17653 ( .A(n13418), .B(n12826), .ZN(n12904) );
  NAND2_X1 U17654 ( .A1(n13934), .A2(n14158), .ZN(n14163) );
  OAI21_X1 U17655 ( .B1(n29735), .B2(n12022), .A(n12354), .ZN(n11738) );
  MUX2_X1 U17656 ( .A(n580), .B(n12350), .S(n12352), .Z(n11737) );
  NOR2_X1 U17657 ( .A1(n12353), .A2(n12352), .ZN(n11736) );
  INV_X1 U17658 ( .A(n13511), .ZN(n11746) );
  INV_X1 U17659 ( .A(n12363), .ZN(n12358) );
  NAND3_X1 U17660 ( .A1(n12358), .A2(n11741), .A3(n12359), .ZN(n11745) );
  NAND3_X1 U17661 ( .A1(n11741), .A2(n11908), .A3(n12356), .ZN(n11744) );
  NAND3_X1 U17662 ( .A1(n12362), .A2(n11742), .A3(n12359), .ZN(n11743) );
  XNOR2_X1 U17663 ( .A(n11746), .B(n13039), .ZN(n12809) );
  NAND2_X1 U17665 ( .A1(n11449), .A2(n11747), .ZN(n12330) );
  XNOR2_X1 U17666 ( .A(n13432), .B(n13547), .ZN(n11749) );
  XNOR2_X1 U17667 ( .A(n12809), .B(n11749), .ZN(n11764) );
  NOR2_X1 U17668 ( .A1(n11751), .A2(n390), .ZN(n11753) );
  NAND2_X1 U17669 ( .A1(n4712), .A2(n11868), .ZN(n11752) );
  XNOR2_X1 U17670 ( .A(n12560), .B(n12699), .ZN(n11762) );
  NAND2_X1 U17672 ( .A1(n11998), .A2(n1831), .ZN(n11758) );
  XNOR2_X1 U17673 ( .A(n13191), .B(n2446), .ZN(n11761) );
  XNOR2_X1 U17674 ( .A(n11762), .B(n11761), .ZN(n11763) );
  XNOR2_X1 U17675 ( .A(n11764), .B(n11763), .ZN(n13936) );
  INV_X1 U17676 ( .A(n13936), .ZN(n13754) );
  NAND2_X1 U17677 ( .A1(n14163), .A2(n13754), .ZN(n11765) );
  NAND2_X1 U17678 ( .A1(n14473), .A2(n13935), .ZN(n11766) );
  INV_X1 U17679 ( .A(n11770), .ZN(n11773) );
  OAI211_X2 U17680 ( .C1(n11773), .C2(n285), .A(n11772), .B(n11771), .ZN(
        n13170) );
  XNOR2_X1 U17681 ( .A(n13170), .B(n13014), .ZN(n13277) );
  INV_X1 U17682 ( .A(n11774), .ZN(n11777) );
  INV_X1 U17683 ( .A(n11131), .ZN(n11776) );
  OAI21_X1 U17684 ( .B1(n11777), .B2(n11776), .A(n11775), .ZN(n11779) );
  MUX2_X1 U17685 ( .A(n11780), .B(n11779), .S(n11778), .Z(n11781) );
  INV_X1 U17686 ( .A(n11781), .ZN(n11786) );
  INV_X1 U17687 ( .A(n12542), .ZN(n12866) );
  NAND2_X1 U17688 ( .A1(n11789), .A2(n2194), .ZN(n11790) );
  XNOR2_X1 U17690 ( .A(n13020), .B(n12866), .ZN(n12634) );
  XNOR2_X1 U17691 ( .A(n12634), .B(n13277), .ZN(n11805) );
  NAND3_X1 U17692 ( .A1(n12289), .A2(n12080), .A3(n29499), .ZN(n11798) );
  NAND2_X1 U17693 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  XNOR2_X1 U17694 ( .A(n12734), .B(n12817), .ZN(n11803) );
  INV_X1 U17695 ( .A(n12407), .ZN(n12278) );
  INV_X1 U17696 ( .A(n3087), .ZN(n27560) );
  XNOR2_X1 U17697 ( .A(n12760), .B(n27560), .ZN(n11802) );
  XNOR2_X1 U17698 ( .A(n11803), .B(n11802), .ZN(n11804) );
  NAND3_X1 U17699 ( .A1(n12201), .A2(n12202), .A3(n12200), .ZN(n11806) );
  NAND3_X1 U17700 ( .A1(n8847), .A2(n11807), .A3(n12201), .ZN(n11808) );
  XNOR2_X1 U17701 ( .A(n12776), .B(n29247), .ZN(n11815) );
  OAI21_X1 U17702 ( .B1(n11812), .B2(n303), .A(n11982), .ZN(n11813) );
  XNOR2_X1 U17703 ( .A(n11815), .B(n12985), .ZN(n11829) );
  INV_X1 U17704 ( .A(n12128), .ZN(n11820) );
  NOR2_X1 U17705 ( .A1(n11819), .A2(n12186), .ZN(n11817) );
  NAND2_X1 U17706 ( .A1(n12128), .A2(n11817), .ZN(n11822) );
  NAND3_X1 U17707 ( .A1(n11820), .A2(n11819), .A3(n12189), .ZN(n11821) );
  NAND4_X1 U17708 ( .A1(n11823), .A2(n11822), .A3(n12127), .A4(n11821), .ZN(
        n13436) );
  AOI21_X1 U17709 ( .B1(n12179), .B2(n11824), .A(n570), .ZN(n11828) );
  NAND2_X1 U17710 ( .A1(n12125), .A2(n12176), .ZN(n11825) );
  AND2_X1 U17711 ( .A1(n12183), .A2(n11825), .ZN(n11827) );
  NAND2_X1 U17712 ( .A1(n1890), .A2(n12180), .ZN(n11826) );
  XNOR2_X1 U17713 ( .A(n13360), .B(n13436), .ZN(n13290) );
  XNOR2_X1 U17714 ( .A(n11829), .B(n13290), .ZN(n11839) );
  OAI21_X2 U17717 ( .B1(n11833), .B2(n12109), .A(n11832), .ZN(n13035) );
  INV_X1 U17718 ( .A(n12512), .ZN(n12510) );
  OAI21_X1 U17719 ( .B1(n12512), .B2(n10863), .A(n6374), .ZN(n11834) );
  XNOR2_X1 U17720 ( .A(n11839), .B(n11838), .ZN(n13778) );
  INV_X1 U17721 ( .A(n13778), .ZN(n14249) );
  NAND3_X1 U17722 ( .A1(n12210), .A2(n12206), .A3(n12211), .ZN(n11841) );
  OAI21_X1 U17723 ( .B1(n11849), .B2(n11848), .A(n5079), .ZN(n11850) );
  AOI21_X1 U17724 ( .B1(n11858), .B2(n11943), .A(n11857), .ZN(n11863) );
  XNOR2_X1 U17725 ( .A(n13566), .B(n13175), .ZN(n12792) );
  XNOR2_X1 U17726 ( .A(n12595), .B(n3537), .ZN(n11864) );
  XNOR2_X1 U17727 ( .A(n12792), .B(n11864), .ZN(n11865) );
  MUX2_X1 U17728 ( .A(n13744), .B(n14249), .S(n29312), .Z(n12010) );
  OAI21_X1 U17729 ( .B1(n578), .B2(n11869), .A(n390), .ZN(n11871) );
  OAI211_X1 U17730 ( .C1(n390), .C2(n4712), .A(n11871), .B(n11870), .ZN(n11873) );
  OAI21_X1 U17731 ( .B1(n11875), .B2(n11877), .A(n567), .ZN(n11882) );
  NOR2_X1 U17732 ( .A1(n11877), .A2(n11876), .ZN(n11880) );
  XNOR2_X1 U17733 ( .A(n12849), .B(n13478), .ZN(n12638) );
  OAI21_X1 U17734 ( .B1(n11884), .B2(n12332), .A(n12327), .ZN(n11891) );
  NAND3_X1 U17735 ( .A1(n11888), .A2(n12018), .A3(n12329), .ZN(n11889) );
  OAI211_X2 U17736 ( .C1(n12014), .C2(n11891), .A(n11890), .B(n11889), .ZN(
        n13136) );
  XNOR2_X1 U17737 ( .A(n12830), .B(n13136), .ZN(n11892) );
  XNOR2_X1 U17738 ( .A(n12638), .B(n11892), .ZN(n11920) );
  INV_X1 U17740 ( .A(n11893), .ZN(n11895) );
  NAND2_X1 U17741 ( .A1(n11895), .A2(n11894), .ZN(n11897) );
  NAND2_X1 U17742 ( .A1(n11900), .A2(n11899), .ZN(n11903) );
  NOR2_X1 U17743 ( .A1(n11903), .A2(n11901), .ZN(n12427) );
  INV_X1 U17744 ( .A(n12427), .ZN(n11902) );
  INV_X1 U17745 ( .A(n11903), .ZN(n11904) );
  NAND3_X1 U17746 ( .A1(n11904), .A2(n29209), .A3(n12350), .ZN(n12430) );
  NAND2_X1 U17748 ( .A1(n12362), .A2(n12359), .ZN(n11911) );
  NAND3_X1 U17749 ( .A1(n12361), .A2(n11908), .A3(n12357), .ZN(n11909) );
  INV_X1 U17752 ( .A(n431), .ZN(n12340) );
  NAND2_X1 U17753 ( .A1(n11915), .A2(n12338), .ZN(n11914) );
  INV_X1 U17754 ( .A(n12339), .ZN(n12344) );
  NAND3_X1 U17755 ( .A1(n12344), .A2(n12343), .A3(n11915), .ZN(n11916) );
  XNOR2_X1 U17756 ( .A(n13482), .B(n2982), .ZN(n11918) );
  XNOR2_X1 U17757 ( .A(n13274), .B(n11918), .ZN(n11919) );
  XNOR2_X1 U17758 ( .A(n11919), .B(n11920), .ZN(n13775) );
  AOI21_X1 U17759 ( .B1(n11922), .B2(n11927), .A(n11921), .ZN(n11926) );
  NOR2_X1 U17760 ( .A1(n11924), .A2(n10905), .ZN(n11925) );
  NOR2_X1 U17761 ( .A1(n12132), .A2(n12267), .ZN(n11929) );
  OAI21_X1 U17762 ( .B1(n11930), .B2(n11929), .A(n11928), .ZN(n11931) );
  INV_X1 U17763 ( .A(n12249), .ZN(n12072) );
  OAI22_X1 U17764 ( .A1(n12251), .A2(n11933), .B1(n11932), .B2(n12072), .ZN(
        n12071) );
  NAND2_X1 U17765 ( .A1(n12071), .A2(n11934), .ZN(n11936) );
  OAI211_X1 U17766 ( .C1(n12070), .C2(n12252), .A(n349), .B(n12072), .ZN(
        n11935) );
  XNOR2_X1 U17767 ( .A(n13265), .B(n11937), .ZN(n11938) );
  XNOR2_X1 U17768 ( .A(n11939), .B(n11938), .ZN(n11961) );
  XNOR2_X1 U17769 ( .A(n13008), .B(n13262), .ZN(n11959) );
  NAND3_X1 U17770 ( .A1(n571), .A2(n6706), .A3(n11953), .ZN(n11957) );
  XNOR2_X1 U17771 ( .A(n13488), .B(n3180), .ZN(n11958) );
  XNOR2_X1 U17772 ( .A(n11958), .B(n11959), .ZN(n11960) );
  XNOR2_X1 U17773 ( .A(n11961), .B(n11960), .ZN(n14078) );
  NAND2_X1 U17774 ( .A1(n12224), .A2(n11962), .ZN(n11968) );
  AOI21_X1 U17775 ( .B1(n11963), .B2(n12042), .A(n11962), .ZN(n11964) );
  NAND3_X1 U17777 ( .A1(n11963), .A2(n11965), .A3(n12218), .ZN(n11966) );
  XNOR2_X1 U17778 ( .A(n13209), .B(n3625), .ZN(n11975) );
  NAND3_X1 U17779 ( .A1(n5839), .A2(n12035), .A3(n12037), .ZN(n11974) );
  INV_X1 U17780 ( .A(n11969), .ZN(n11970) );
  NAND3_X1 U17781 ( .A1(n11970), .A2(n12157), .A3(n12241), .ZN(n11972) );
  NAND3_X1 U17782 ( .A1(n11969), .A2(n12159), .A3(n12241), .ZN(n11971) );
  NOR2_X1 U17783 ( .A1(n776), .A2(n12234), .ZN(n11976) );
  NOR2_X1 U17784 ( .A1(n11976), .A2(n5009), .ZN(n11978) );
  NAND3_X1 U17785 ( .A1(n13081), .A2(n11982), .A3(n303), .ZN(n11986) );
  NAND4_X1 U17786 ( .A1(n11984), .A2(n13086), .A3(n13084), .A4(n11983), .ZN(
        n11985) );
  XNOR2_X1 U17787 ( .A(n13133), .B(n13543), .ZN(n12492) );
  XNOR2_X1 U17788 ( .A(n11988), .B(n12492), .ZN(n12007) );
  INV_X1 U17789 ( .A(n12747), .ZN(n12005) );
  NAND2_X1 U17791 ( .A1(n11990), .A2(n11989), .ZN(n11991) );
  NAND2_X1 U17792 ( .A1(n12000), .A2(n11996), .ZN(n12003) );
  INV_X1 U17793 ( .A(n11995), .ZN(n11999) );
  NAND2_X1 U17794 ( .A1(n11996), .A2(n1831), .ZN(n11997) );
  NAND3_X1 U17795 ( .A1(n6658), .A2(n572), .A3(n12001), .ZN(n12002) );
  XNOR2_X1 U17796 ( .A(n13028), .B(n12879), .ZN(n12648) );
  XNOR2_X1 U17797 ( .A(n12005), .B(n12648), .ZN(n12006) );
  XNOR2_X1 U17798 ( .A(n12007), .B(n12006), .ZN(n13776) );
  NAND2_X1 U17799 ( .A1(n13776), .A2(n14252), .ZN(n13745) );
  INV_X1 U17800 ( .A(n13745), .ZN(n12008) );
  NAND2_X1 U17801 ( .A1(n12008), .A2(n14254), .ZN(n12009) );
  AOI22_X1 U17803 ( .A1(n12012), .A2(n15406), .B1(n12011), .B2(n3362), .ZN(
        n12372) );
  AND2_X1 U17804 ( .A1(n12013), .A2(n12018), .ZN(n12021) );
  INV_X1 U17805 ( .A(n12014), .ZN(n12020) );
  OAI21_X1 U17806 ( .B1(n12021), .B2(n12020), .A(n12019), .ZN(n12388) );
  XNOR2_X1 U17807 ( .A(n12684), .B(n3787), .ZN(n12025) );
  OAI211_X1 U17808 ( .C1(n12022), .C2(n12354), .A(n11467), .B(n580), .ZN(
        n12023) );
  OAI211_X1 U17809 ( .C1(n29735), .C2(n29209), .A(n12024), .B(n12023), .ZN(
        n13348) );
  XNOR2_X1 U17810 ( .A(n13246), .B(n12025), .ZN(n12033) );
  XNOR2_X1 U17811 ( .A(n13195), .B(n12965), .ZN(n12797) );
  NOR2_X1 U17812 ( .A1(n12026), .A2(n12337), .ZN(n12031) );
  OAI21_X1 U17813 ( .B1(n12028), .B2(n12337), .A(n12027), .ZN(n12029) );
  XNOR2_X1 U17814 ( .A(n12913), .B(n12686), .ZN(n13425) );
  XNOR2_X1 U17815 ( .A(n13425), .B(n12797), .ZN(n12032) );
  XNOR2_X1 U17816 ( .A(n12033), .B(n12032), .ZN(n14481) );
  XNOR2_X1 U17817 ( .A(n12954), .B(n2381), .ZN(n12034) );
  XNOR2_X1 U17818 ( .A(n12396), .B(n13012), .ZN(n13441) );
  MUX2_X1 U17819 ( .A(n12042), .B(n12041), .S(n12220), .Z(n12046) );
  XNOR2_X1 U17820 ( .A(n13525), .B(n13171), .ZN(n13015) );
  XNOR2_X1 U17821 ( .A(n13051), .B(n13015), .ZN(n12047) );
  NOR2_X1 U17822 ( .A1(n12053), .A2(n12051), .ZN(n12052) );
  OAI21_X1 U17823 ( .B1(n6920), .B2(n12052), .A(n566), .ZN(n12056) );
  NAND2_X1 U17824 ( .A1(n12054), .A2(n285), .ZN(n12055) );
  OAI211_X1 U17825 ( .C1(n566), .C2(n12057), .A(n12056), .B(n12055), .ZN(
        n13341) );
  INV_X1 U17826 ( .A(n12058), .ZN(n12297) );
  NAND2_X1 U17827 ( .A1(n12288), .A2(n12297), .ZN(n12063) );
  XNOR2_X1 U17828 ( .A(n13341), .B(n12697), .ZN(n12410) );
  NAND2_X1 U17829 ( .A1(n12279), .A2(n12401), .ZN(n12068) );
  NAND3_X1 U17830 ( .A1(n12408), .A2(n12278), .A3(n12402), .ZN(n12066) );
  NAND4_X1 U17831 ( .A1(n12068), .A2(n12067), .A3(n12404), .A4(n12066), .ZN(
        n12069) );
  NAND2_X1 U17832 ( .A1(n29306), .A2(n12120), .ZN(n13766) );
  OAI21_X1 U17833 ( .B1(n349), .B2(n12072), .A(n12253), .ZN(n12073) );
  NAND2_X1 U17834 ( .A1(n12073), .A2(n12251), .ZN(n12074) );
  OAI21_X1 U17835 ( .B1(n12271), .B2(n28202), .A(n12576), .ZN(n12076) );
  XNOR2_X1 U17836 ( .A(n12677), .B(n3565), .ZN(n12078) );
  XNOR2_X1 U17837 ( .A(n13229), .B(n12078), .ZN(n12086) );
  XNOR2_X1 U17838 ( .A(n12948), .B(n565), .ZN(n12789) );
  NOR2_X1 U17839 ( .A1(n12080), .A2(n3558), .ZN(n12083) );
  XNOR2_X1 U17842 ( .A(n13451), .B(n13447), .ZN(n13283) );
  XNOR2_X1 U17843 ( .A(n13283), .B(n12789), .ZN(n12085) );
  NAND2_X1 U17845 ( .A1(n12990), .A2(n12088), .ZN(n12089) );
  INV_X1 U17847 ( .A(n12091), .ZN(n12095) );
  INV_X1 U17848 ( .A(n12092), .ZN(n12093) );
  NAND3_X1 U17849 ( .A1(n12095), .A2(n12094), .A3(n12093), .ZN(n12096) );
  NOR2_X1 U17850 ( .A1(n12097), .A2(n12096), .ZN(n12992) );
  NAND2_X1 U17851 ( .A1(n12155), .A2(n12992), .ZN(n12098) );
  MUX2_X1 U17852 ( .A(n28828), .B(n12102), .S(n12164), .Z(n12107) );
  OAI21_X2 U17854 ( .B1(n12107), .B2(n12167), .A(n12106), .ZN(n13370) );
  XNOR2_X1 U17855 ( .A(n13331), .B(n13370), .ZN(n12383) );
  OAI21_X1 U17857 ( .B1(n12211), .B2(n12206), .A(n12210), .ZN(n12114) );
  NAND3_X1 U17858 ( .A1(n12111), .A2(n12110), .A3(n12109), .ZN(n12112) );
  XNOR2_X1 U17859 ( .A(n1857), .B(n2441), .ZN(n12116) );
  XNOR2_X1 U17860 ( .A(n12117), .B(n12116), .ZN(n12118) );
  INV_X1 U17861 ( .A(n29306), .ZN(n14485) );
  NAND2_X1 U17862 ( .A1(n570), .A2(n12180), .ZN(n13205) );
  MUX2_X1 U17863 ( .A(n1890), .B(n12177), .S(n12176), .Z(n13202) );
  INV_X1 U17864 ( .A(n13202), .ZN(n12123) );
  MUX2_X1 U17865 ( .A(n13205), .B(n12123), .S(n13206), .Z(n12126) );
  NAND3_X1 U17866 ( .A1(n12181), .A2(n12125), .A3(n12124), .ZN(n13203) );
  NAND3_X1 U17868 ( .A1(n12129), .A2(n12186), .A3(n12128), .ZN(n12130) );
  INV_X1 U17869 ( .A(n13027), .ZN(n12135) );
  XNOR2_X1 U17870 ( .A(n12135), .B(n13296), .ZN(n12139) );
  XNOR2_X1 U17871 ( .A(n13405), .B(n3654), .ZN(n12137) );
  XNOR2_X1 U17872 ( .A(n12136), .B(n12137), .ZN(n12138) );
  NAND3_X1 U17873 ( .A1(n14485), .A2(n14484), .A3(n13947), .ZN(n12140) );
  INV_X1 U17874 ( .A(n12142), .ZN(n12143) );
  NOR2_X1 U17875 ( .A1(n12146), .A2(n12145), .ZN(n12147) );
  NOR3_X1 U17876 ( .A1(n12151), .A2(n3961), .A3(n12991), .ZN(n12153) );
  NOR2_X1 U17877 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  XNOR2_X1 U17878 ( .A(n13433), .B(n12559), .ZN(n12717) );
  INV_X1 U17879 ( .A(n12717), .ZN(n12160) );
  XNOR2_X1 U17880 ( .A(n13236), .B(n13039), .ZN(n12609) );
  XNOR2_X1 U17881 ( .A(n12160), .B(n12609), .ZN(n12175) );
  XNOR2_X1 U17882 ( .A(n13547), .B(n13338), .ZN(n12173) );
  AND2_X1 U17883 ( .A1(n12163), .A2(n1931), .ZN(n12161) );
  NAND2_X1 U17884 ( .A1(n12162), .A2(n12161), .ZN(n12170) );
  NAND3_X1 U17885 ( .A1(n28828), .A2(n11378), .A3(n12164), .ZN(n12169) );
  NAND3_X1 U17886 ( .A1(n12167), .A2(n11378), .A3(n1931), .ZN(n12168) );
  XNOR2_X1 U17887 ( .A(n13113), .B(n1923), .ZN(n12172) );
  XNOR2_X1 U17888 ( .A(n12173), .B(n12172), .ZN(n12174) );
  NOR2_X1 U17889 ( .A1(n12177), .A2(n12176), .ZN(n12178) );
  MUX2_X1 U17890 ( .A(n12179), .B(n12178), .S(n570), .Z(n12185) );
  NOR2_X1 U17891 ( .A1(n12181), .A2(n12180), .ZN(n12182) );
  NOR2_X1 U17892 ( .A1(n12183), .A2(n12182), .ZN(n12184) );
  NAND2_X1 U17894 ( .A1(n12186), .A2(n12189), .ZN(n12197) );
  NAND2_X1 U17895 ( .A1(n12187), .A2(n12186), .ZN(n12193) );
  NOR2_X1 U17896 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  OAI21_X1 U17897 ( .B1(n12193), .B2(n12192), .A(n12191), .ZN(n12196) );
  OAI211_X1 U17898 ( .C1(n12198), .C2(n12197), .A(n12196), .B(n12195), .ZN(
        n13428) );
  XNOR2_X1 U17899 ( .A(n13261), .B(n13428), .ZN(n12721) );
  XNOR2_X1 U17900 ( .A(n13552), .B(n12854), .ZN(n12199) );
  XNOR2_X1 U17901 ( .A(n12721), .B(n12199), .ZN(n12216) );
  OAI21_X1 U17902 ( .B1(n12206), .B2(n12210), .A(n12207), .ZN(n12213) );
  AOI22_X1 U17903 ( .A1(n12211), .A2(n12210), .B1(n12209), .B2(n12208), .ZN(
        n12212) );
  OAI21_X1 U17904 ( .B1(n6281), .B2(n12213), .A(n12212), .ZN(n12658) );
  XNOR2_X1 U17905 ( .A(n12658), .B(n12799), .ZN(n12484) );
  XNOR2_X1 U17906 ( .A(n13043), .B(n3695), .ZN(n12214) );
  XNOR2_X1 U17907 ( .A(n12484), .B(n12214), .ZN(n12215) );
  XNOR2_X1 U17908 ( .A(n12216), .B(n12215), .ZN(n14268) );
  AOI22_X1 U17909 ( .A1(n28726), .A2(n12220), .B1(n12221), .B2(n12218), .ZN(
        n12225) );
  MUX2_X1 U17910 ( .A(n12222), .B(n12221), .S(n12220), .Z(n12223) );
  XNOR2_X1 U17911 ( .A(n12872), .B(n13285), .ZN(n12238) );
  NAND2_X1 U17912 ( .A1(n12228), .A2(n13086), .ZN(n12229) );
  XNOR2_X1 U17913 ( .A(n13448), .B(n12472), .ZN(n12423) );
  INV_X1 U17914 ( .A(n12423), .ZN(n12237) );
  XNOR2_X1 U17915 ( .A(n12237), .B(n12238), .ZN(n12248) );
  XNOR2_X1 U17916 ( .A(n13055), .B(n13226), .ZN(n12246) );
  NAND2_X1 U17917 ( .A1(n12242), .A2(n12241), .ZN(n12243) );
  INV_X1 U17918 ( .A(n22072), .ZN(n25361) );
  XNOR2_X1 U17919 ( .A(n12790), .B(n25361), .ZN(n12245) );
  XNOR2_X1 U17920 ( .A(n12245), .B(n12246), .ZN(n12247) );
  NAND2_X1 U17921 ( .A1(n12252), .A2(n12249), .ZN(n12250) );
  OAI21_X1 U17922 ( .B1(n12251), .B2(n12252), .A(n12250), .ZN(n12255) );
  XNOR2_X1 U17923 ( .A(n12262), .B(n12735), .ZN(n12269) );
  XNOR2_X1 U17924 ( .A(n12866), .B(n12632), .ZN(n12268) );
  XNOR2_X1 U17925 ( .A(n12269), .B(n12268), .ZN(n12277) );
  MUX2_X1 U17926 ( .A(n28202), .B(n12270), .S(n12271), .Z(n12274) );
  INV_X1 U17927 ( .A(n12271), .ZN(n12272) );
  XNOR2_X1 U17928 ( .A(n13080), .B(n13048), .ZN(n12275) );
  XNOR2_X1 U17929 ( .A(n13219), .B(n12275), .ZN(n12276) );
  XNOR2_X1 U17930 ( .A(n12277), .B(n12276), .ZN(n13749) );
  INV_X1 U17931 ( .A(n13749), .ZN(n14099) );
  MUX2_X1 U17932 ( .A(n12278), .B(n12280), .S(n12402), .Z(n12287) );
  OAI21_X1 U17933 ( .B1(n12407), .B2(n12281), .A(n12280), .ZN(n12282) );
  NAND3_X1 U17934 ( .A1(n12284), .A2(n12283), .A3(n12282), .ZN(n12285) );
  OAI21_X1 U17935 ( .B1(n12287), .B2(n12286), .A(n12285), .ZN(n12752) );
  NAND4_X1 U17936 ( .A1(n12061), .A2(n29324), .A3(n12291), .A4(n12290), .ZN(
        n12294) );
  XNOR2_X1 U17937 ( .A(n12783), .B(n13121), .ZN(n12465) );
  XNOR2_X1 U17938 ( .A(n12465), .B(n12298), .ZN(n12326) );
  OAI21_X1 U17940 ( .B1(n12305), .B2(n28807), .A(n12300), .ZN(n12310) );
  AND2_X1 U17941 ( .A1(n12302), .A2(n12304), .ZN(n12308) );
  NOR2_X1 U17942 ( .A1(n12304), .A2(n12303), .ZN(n12306) );
  AOI22_X1 U17943 ( .A1(n12308), .A2(n4197), .B1(n12306), .B2(n12305), .ZN(
        n12309) );
  NAND2_X1 U17945 ( .A1(n12312), .A2(n12316), .ZN(n12319) );
  NAND2_X1 U17946 ( .A1(n12321), .A2(n12313), .ZN(n12314) );
  OAI21_X1 U17947 ( .B1(n12316), .B2(n12315), .A(n12314), .ZN(n12317) );
  INV_X1 U17948 ( .A(n12317), .ZN(n12318) );
  NAND3_X1 U17949 ( .A1(n12322), .A2(n12321), .A3(n12320), .ZN(n12323) );
  XNOR2_X1 U17950 ( .A(n13419), .B(n13272), .ZN(n13140) );
  XNOR2_X1 U17951 ( .A(n12849), .B(n3154), .ZN(n12324) );
  XNOR2_X1 U17952 ( .A(n13140), .B(n12324), .ZN(n12325) );
  XNOR2_X2 U17953 ( .A(n12326), .B(n12325), .ZN(n14262) );
  NOR2_X1 U17954 ( .A1(n14262), .A2(n1743), .ZN(n12367) );
  AOI21_X1 U17955 ( .B1(n12329), .B2(n12328), .A(n12327), .ZN(n12331) );
  MUX2_X1 U17956 ( .A(n12332), .B(n12331), .S(n12330), .Z(n12336) );
  NOR2_X1 U17957 ( .A1(n12334), .A2(n12333), .ZN(n12335) );
  OAI22_X1 U17958 ( .A1(n1291), .A2(n12341), .B1(n6919), .B2(n12340), .ZN(
        n12348) );
  AOI21_X1 U17960 ( .B1(n12346), .B2(n12345), .A(n12344), .ZN(n12347) );
  NOR2_X1 U17961 ( .A1(n12348), .A2(n12347), .ZN(n12572) );
  INV_X1 U17962 ( .A(n12572), .ZN(n12768) );
  XNOR2_X1 U17963 ( .A(n12768), .B(n12644), .ZN(n12460) );
  XNOR2_X1 U17964 ( .A(n12460), .B(n12349), .ZN(n12366) );
  MUX2_X1 U17965 ( .A(n11467), .B(n580), .S(n12350), .Z(n12351) );
  NAND2_X1 U17966 ( .A1(n12351), .A2(n29735), .ZN(n12355) );
  XNOR2_X1 U17967 ( .A(n13298), .B(n13461), .ZN(n12749) );
  XNOR2_X1 U17968 ( .A(n12879), .B(n3586), .ZN(n12364) );
  XNOR2_X1 U17969 ( .A(n12749), .B(n12364), .ZN(n12365) );
  XNOR2_X1 U17970 ( .A(n12365), .B(n12366), .ZN(n14264) );
  OAI21_X1 U17971 ( .B1(n13613), .B2(n12367), .A(n13762), .ZN(n12368) );
  XNOR2_X1 U17972 ( .A(n16310), .B(n27105), .ZN(n12631) );
  XNOR2_X1 U17973 ( .A(n13297), .B(n29064), .ZN(n12374) );
  XNOR2_X1 U17974 ( .A(n13459), .B(n2511), .ZN(n12373) );
  XNOR2_X1 U17975 ( .A(n12374), .B(n12373), .ZN(n12376) );
  XNOR2_X1 U17976 ( .A(n13027), .B(n13542), .ZN(n12375) );
  XNOR2_X1 U17977 ( .A(n12677), .B(n3457), .ZN(n12378) );
  XNOR2_X1 U17978 ( .A(n12379), .B(n12378), .ZN(n12382) );
  XNOR2_X1 U17979 ( .A(n13179), .B(n13226), .ZN(n13565) );
  INV_X1 U17982 ( .A(n14331), .ZN(n14336) );
  XNOR2_X1 U17983 ( .A(n13249), .B(n13533), .ZN(n12691) );
  XNOR2_X1 U17984 ( .A(n12383), .B(n12691), .ZN(n12387) );
  XNOR2_X1 U17985 ( .A(n12385), .B(n12384), .ZN(n12386) );
  INV_X1 U17986 ( .A(n12388), .ZN(n13005) );
  XNOR2_X1 U17987 ( .A(n12913), .B(n12723), .ZN(n12391) );
  XNOR2_X1 U17988 ( .A(n13348), .B(n3491), .ZN(n12390) );
  XNOR2_X1 U17989 ( .A(n12391), .B(n12390), .ZN(n12392) );
  INV_X1 U17991 ( .A(n14406), .ZN(n13878) );
  NAND2_X1 U17992 ( .A1(n14332), .A2(n13878), .ZN(n12399) );
  INV_X1 U17993 ( .A(n13015), .ZN(n12395) );
  XNOR2_X1 U17994 ( .A(n13278), .B(n2987), .ZN(n12394) );
  XNOR2_X1 U17995 ( .A(n12395), .B(n12394), .ZN(n12398) );
  XNOR2_X1 U17996 ( .A(n12738), .B(n12868), .ZN(n12815) );
  XNOR2_X1 U17997 ( .A(n13522), .B(n12815), .ZN(n12397) );
  INV_X1 U17998 ( .A(n14407), .ZN(n13879) );
  NAND2_X1 U17999 ( .A1(n12402), .A2(n12278), .ZN(n12403) );
  NAND3_X1 U18000 ( .A1(n12405), .A2(n12404), .A3(n12403), .ZN(n12406) );
  OAI21_X1 U18001 ( .B1(n12408), .B2(n12407), .A(n12406), .ZN(n12860) );
  XNOR2_X1 U18002 ( .A(n13109), .B(n12860), .ZN(n12807) );
  XNOR2_X1 U18003 ( .A(n13547), .B(n13190), .ZN(n12698) );
  XNOR2_X1 U18004 ( .A(n12698), .B(n12807), .ZN(n12412) );
  XNOR2_X1 U18005 ( .A(n13291), .B(n3516), .ZN(n12409) );
  XNOR2_X1 U18006 ( .A(n12410), .B(n12409), .ZN(n12411) );
  XNOR2_X1 U18007 ( .A(n12411), .B(n12412), .ZN(n14330) );
  INV_X1 U18008 ( .A(n14330), .ZN(n14405) );
  NAND3_X1 U18009 ( .A1(n13879), .A2(n14405), .A3(n29607), .ZN(n12415) );
  NOR2_X1 U18010 ( .A1(n29607), .A2(n13878), .ZN(n12413) );
  NAND2_X1 U18011 ( .A1(n14411), .A2(n12413), .ZN(n12414) );
  NAND2_X1 U18012 ( .A1(n14904), .A2(n14906), .ZN(n14903) );
  INV_X1 U18013 ( .A(n14903), .ZN(n13993) );
  XNOR2_X1 U18014 ( .A(n13402), .B(n12588), .ZN(n12419) );
  XNOR2_X1 U18015 ( .A(n13461), .B(n22489), .ZN(n12416) );
  XNOR2_X1 U18016 ( .A(n12417), .B(n12416), .ZN(n12418) );
  INV_X1 U18017 ( .A(n13287), .ZN(n13378) );
  XNOR2_X1 U18018 ( .A(n12421), .B(n13378), .ZN(n12425) );
  XNOR2_X1 U18019 ( .A(n13451), .B(n3380), .ZN(n12422) );
  XNOR2_X1 U18020 ( .A(n12423), .B(n12422), .ZN(n12424) );
  NOR2_X1 U18021 ( .A1(n30), .A2(n29628), .ZN(n12452) );
  XNOR2_X1 U18022 ( .A(n13121), .B(n13482), .ZN(n12616) );
  INV_X1 U18023 ( .A(n12616), .ZN(n12426) );
  XNOR2_X1 U18024 ( .A(n13419), .B(n13270), .ZN(n13374) );
  XNOR2_X1 U18025 ( .A(n12426), .B(n13374), .ZN(n12434) );
  XNOR2_X1 U18026 ( .A(n13269), .B(n13136), .ZN(n12433) );
  AND2_X1 U18027 ( .A1(n12427), .A2(n12428), .ZN(n12431) );
  XNOR2_X1 U18028 ( .A(n13369), .B(n1175), .ZN(n12432) );
  XNOR2_X1 U18029 ( .A(n12658), .B(n13488), .ZN(n12620) );
  XNOR2_X1 U18030 ( .A(n12620), .B(n12435), .ZN(n12439) );
  XNOR2_X1 U18031 ( .A(n13262), .B(n12686), .ZN(n12437) );
  XNOR2_X1 U18032 ( .A(n13428), .B(n27298), .ZN(n12436) );
  XNOR2_X1 U18033 ( .A(n12437), .B(n12436), .ZN(n12438) );
  NAND2_X1 U18034 ( .A1(n13877), .A2(n14399), .ZN(n12451) );
  XNOR2_X1 U18035 ( .A(n12776), .B(n3036), .ZN(n12440) );
  XNOR2_X1 U18036 ( .A(n13433), .B(n12440), .ZN(n12443) );
  INV_X1 U18037 ( .A(n13360), .ZN(n12441) );
  XNOR2_X1 U18038 ( .A(n13236), .B(n12441), .ZN(n12442) );
  XNOR2_X1 U18039 ( .A(n12443), .B(n12442), .ZN(n12446) );
  INV_X1 U18040 ( .A(n13035), .ZN(n12444) );
  XNOR2_X1 U18041 ( .A(n13364), .B(n12699), .ZN(n12987) );
  XNOR2_X1 U18042 ( .A(n12444), .B(n12987), .ZN(n12445) );
  NOR2_X1 U18043 ( .A1(n14402), .A2(n14399), .ZN(n13963) );
  XNOR2_X1 U18044 ( .A(n12894), .B(n12632), .ZN(n12449) );
  XNOR2_X1 U18045 ( .A(n12760), .B(n3508), .ZN(n12447) );
  XNOR2_X1 U18046 ( .A(n12447), .B(n13445), .ZN(n12448) );
  XNOR2_X1 U18047 ( .A(n13170), .B(n12734), .ZN(n12450) );
  INV_X1 U18048 ( .A(n15097), .ZN(n14901) );
  XNOR2_X1 U18049 ( .A(n13020), .B(n12453), .ZN(n13147) );
  INV_X1 U18050 ( .A(n13147), .ZN(n13497) );
  XNOR2_X1 U18051 ( .A(n13497), .B(n12454), .ZN(n12458) );
  XNOR2_X1 U18052 ( .A(n12763), .B(n12632), .ZN(n12456) );
  XNOR2_X1 U18053 ( .A(n12735), .B(n5633), .ZN(n12455) );
  XOR2_X1 U18054 ( .A(n12455), .B(n12456), .Z(n12457) );
  XNOR2_X1 U18055 ( .A(n12841), .B(n13405), .ZN(n12459) );
  XNOR2_X1 U18056 ( .A(n12460), .B(n12459), .ZN(n12464) );
  XNOR2_X1 U18057 ( .A(n13404), .B(n3728), .ZN(n12462) );
  XNOR2_X1 U18058 ( .A(n13028), .B(n12461), .ZN(n13505) );
  XNOR2_X1 U18059 ( .A(n12462), .B(n13505), .ZN(n12463) );
  XNOR2_X1 U18061 ( .A(n13478), .B(n12780), .ZN(n13141) );
  XNOR2_X1 U18062 ( .A(n13141), .B(n12465), .ZN(n12469) );
  XNOR2_X1 U18063 ( .A(n13272), .B(n2912), .ZN(n12467) );
  XNOR2_X1 U18064 ( .A(n12467), .B(n12466), .ZN(n12468) );
  XNOR2_X1 U18065 ( .A(n12469), .B(n12468), .ZN(n13686) );
  INV_X1 U18066 ( .A(n13686), .ZN(n12481) );
  NAND2_X1 U18067 ( .A1(n14417), .A2(n12470), .ZN(n12475) );
  XNOR2_X1 U18068 ( .A(n13285), .B(n12978), .ZN(n13474) );
  XNOR2_X1 U18069 ( .A(n13054), .B(n13563), .ZN(n12471) );
  XNOR2_X1 U18070 ( .A(n12948), .B(n13231), .ZN(n12474) );
  INV_X1 U18071 ( .A(n1133), .ZN(n28073) );
  XNOR2_X1 U18072 ( .A(n13381), .B(n28073), .ZN(n12473) );
  NAND2_X1 U18073 ( .A1(n12475), .A2(n14414), .ZN(n12489) );
  XNOR2_X1 U18074 ( .A(n13236), .B(n13359), .ZN(n12477) );
  XNOR2_X1 U18076 ( .A(n13113), .B(n12985), .ZN(n13509) );
  XNOR2_X1 U18077 ( .A(n12560), .B(n1046), .ZN(n12478) );
  XNOR2_X1 U18078 ( .A(n13509), .B(n12478), .ZN(n12479) );
  XNOR2_X1 U18079 ( .A(n13261), .B(n13008), .ZN(n13487) );
  XNOR2_X1 U18080 ( .A(n12965), .B(n13386), .ZN(n12482) );
  XNOR2_X1 U18081 ( .A(n13487), .B(n12482), .ZN(n12486) );
  XNOR2_X1 U18082 ( .A(n12566), .B(n3317), .ZN(n12483) );
  XNOR2_X1 U18083 ( .A(n12484), .B(n12483), .ZN(n12485) );
  XNOR2_X1 U18084 ( .A(n12486), .B(n12485), .ZN(n14215) );
  INV_X1 U18085 ( .A(n14215), .ZN(n13891) );
  NAND3_X1 U18086 ( .A1(n13891), .A2(n14415), .A3(n14217), .ZN(n12487) );
  AND2_X1 U18087 ( .A1(n14413), .A2(n12487), .ZN(n12488) );
  NAND2_X1 U18088 ( .A1(n12489), .A2(n12488), .ZN(n14902) );
  INV_X1 U18089 ( .A(n14902), .ZN(n14578) );
  XNOR2_X1 U18091 ( .A(n13457), .B(n12490), .ZN(n12494) );
  XNOR2_X1 U18092 ( .A(n12881), .B(n27231), .ZN(n12491) );
  XNOR2_X1 U18093 ( .A(n12492), .B(n12491), .ZN(n12493) );
  XNOR2_X1 U18095 ( .A(n13414), .B(n13136), .ZN(n12498) );
  INV_X1 U18096 ( .A(n12495), .ZN(n12496) );
  XNOR2_X1 U18097 ( .A(n12496), .B(n13137), .ZN(n12847) );
  INV_X1 U18098 ( .A(n12847), .ZN(n12497) );
  XNOR2_X1 U18099 ( .A(n12497), .B(n12498), .ZN(n12502) );
  XNOR2_X1 U18100 ( .A(n13413), .B(n13420), .ZN(n12500) );
  XNOR2_X1 U18101 ( .A(n12500), .B(n12499), .ZN(n12501) );
  INV_X1 U18102 ( .A(n857), .ZN(n12503) );
  XNOR2_X1 U18103 ( .A(n12504), .B(n12503), .ZN(n12505) );
  XNOR2_X1 U18104 ( .A(n12505), .B(n13278), .ZN(n12506) );
  XNOR2_X1 U18105 ( .A(n13018), .B(n12734), .ZN(n13146) );
  XNOR2_X1 U18106 ( .A(n12506), .B(n13146), .ZN(n12515) );
  NOR2_X1 U18107 ( .A1(n12508), .A2(n12507), .ZN(n12509) );
  AOI22_X1 U18108 ( .A1(n12511), .A2(n12510), .B1(n12509), .B2(n3653), .ZN(
        n12513) );
  XNOR2_X1 U18109 ( .A(n12515), .B(n13442), .ZN(n13703) );
  XNOR2_X1 U18111 ( .A(n12696), .B(n13035), .ZN(n13155) );
  INV_X1 U18112 ( .A(n13155), .ZN(n12522) );
  AOI21_X1 U18113 ( .B1(n5947), .B2(n12578), .A(n12516), .ZN(n12518) );
  OAI22_X1 U18114 ( .A1(n12518), .A2(n12583), .B1(n5947), .B2(n12272), .ZN(
        n12520) );
  NAND2_X1 U18115 ( .A1(n12520), .A2(n12519), .ZN(n12521) );
  XNOR2_X1 U18117 ( .A(n13191), .B(n13436), .ZN(n12524) );
  XNOR2_X1 U18118 ( .A(n13291), .B(n28294), .ZN(n12523) );
  XNOR2_X1 U18119 ( .A(n12524), .B(n12523), .ZN(n12525) );
  INV_X1 U18121 ( .A(n3633), .ZN(n12527) );
  XNOR2_X1 U18122 ( .A(n13159), .B(n12527), .ZN(n12528) );
  XNOR2_X1 U18123 ( .A(n13380), .B(n13567), .ZN(n12876) );
  XNOR2_X1 U18124 ( .A(n12528), .B(n12876), .ZN(n12531) );
  XNOR2_X1 U18125 ( .A(n13566), .B(n12788), .ZN(n13284) );
  XNOR2_X1 U18126 ( .A(n13230), .B(n12529), .ZN(n13180) );
  NAND2_X1 U18128 ( .A1(n13872), .A2(n12534), .ZN(n14425) );
  INV_X1 U18129 ( .A(n14425), .ZN(n14306) );
  XNOR2_X1 U18130 ( .A(n13150), .B(n3483), .ZN(n12535) );
  XNOR2_X1 U18131 ( .A(n12535), .B(n13260), .ZN(n12537) );
  INV_X1 U18132 ( .A(n13265), .ZN(n12536) );
  XNOR2_X1 U18133 ( .A(n12914), .B(n12536), .ZN(n13426) );
  XNOR2_X1 U18134 ( .A(n13426), .B(n12537), .ZN(n12540) );
  INV_X1 U18135 ( .A(n13553), .ZN(n12657) );
  XNOR2_X1 U18136 ( .A(n12657), .B(n12538), .ZN(n12539) );
  NAND2_X1 U18137 ( .A1(n14306), .A2(n14426), .ZN(n14905) );
  INV_X1 U18140 ( .A(n15098), .ZN(n15095) );
  XNOR2_X1 U18141 ( .A(n12762), .B(n3035), .ZN(n12543) );
  XNOR2_X1 U18142 ( .A(n12543), .B(n13051), .ZN(n12544) );
  XNOR2_X1 U18143 ( .A(n12544), .B(n13315), .ZN(n12547) );
  XNOR2_X1 U18144 ( .A(n13171), .B(n12600), .ZN(n12545) );
  XNOR2_X1 U18145 ( .A(n12816), .B(n12545), .ZN(n12546) );
  XNOR2_X1 U18146 ( .A(n12547), .B(n12546), .ZN(n14319) );
  INV_X1 U18147 ( .A(n14319), .ZN(n14310) );
  XNOR2_X1 U18148 ( .A(n12548), .B(n12872), .ZN(n13095) );
  XNOR2_X1 U18149 ( .A(n13097), .B(n13563), .ZN(n12549) );
  XNOR2_X1 U18150 ( .A(n12549), .B(n13095), .ZN(n12553) );
  XNOR2_X1 U18151 ( .A(n12677), .B(n3643), .ZN(n12550) );
  XNOR2_X1 U18152 ( .A(n12550), .B(n12551), .ZN(n12552) );
  XNOR2_X1 U18153 ( .A(n13418), .B(n13069), .ZN(n12851) );
  XNOR2_X1 U18154 ( .A(n12851), .B(n13332), .ZN(n12558) );
  XNOR2_X1 U18155 ( .A(n13370), .B(n12783), .ZN(n12556) );
  XNOR2_X1 U18156 ( .A(n12827), .B(n3501), .ZN(n12555) );
  XNOR2_X1 U18157 ( .A(n12556), .B(n12555), .ZN(n12557) );
  XNOR2_X1 U18158 ( .A(n12558), .B(n12557), .ZN(n13257) );
  MUX2_X1 U18159 ( .A(n14310), .B(n14313), .S(n14320), .Z(n12587) );
  XNOR2_X1 U18160 ( .A(n13432), .B(n13034), .ZN(n12562) );
  XNOR2_X1 U18161 ( .A(n12560), .B(n12697), .ZN(n13192) );
  INV_X1 U18162 ( .A(n13192), .ZN(n12561) );
  XNOR2_X1 U18163 ( .A(n12561), .B(n12562), .ZN(n12565) );
  XNOR2_X1 U18164 ( .A(n13511), .B(n13036), .ZN(n13112) );
  XNOR2_X1 U18165 ( .A(n13338), .B(n3323), .ZN(n12563) );
  XNOR2_X1 U18166 ( .A(n13112), .B(n12563), .ZN(n12564) );
  INV_X1 U18168 ( .A(n14318), .ZN(n13711) );
  XNOR2_X1 U18169 ( .A(n13005), .B(n12566), .ZN(n13197) );
  INV_X1 U18170 ( .A(n13197), .ZN(n12567) );
  XNOR2_X1 U18171 ( .A(n12567), .B(n13347), .ZN(n12571) );
  XNOR2_X1 U18172 ( .A(n12568), .B(n13245), .ZN(n12570) );
  XNOR2_X1 U18173 ( .A(n13101), .B(n3528), .ZN(n12569) );
  NAND3_X1 U18175 ( .A1(n14319), .A2(n13711), .A3(n13884), .ZN(n12586) );
  XNOR2_X1 U18176 ( .A(n13406), .B(n12841), .ZN(n12574) );
  XNOR2_X1 U18177 ( .A(n12572), .B(n13075), .ZN(n12573) );
  XNOR2_X1 U18178 ( .A(n12574), .B(n12573), .ZN(n12584) );
  OAI21_X1 U18179 ( .B1(n28202), .B2(n12576), .A(n12575), .ZN(n12582) );
  NAND2_X1 U18180 ( .A1(n12579), .A2(n12578), .ZN(n12580) );
  OAI211_X1 U18181 ( .C1(n12583), .C2(n12582), .A(n12581), .B(n12580), .ZN(
        n12883) );
  XNOR2_X1 U18182 ( .A(n13504), .B(n12879), .ZN(n13322) );
  XNOR2_X1 U18183 ( .A(n12747), .B(n13404), .ZN(n13503) );
  XNOR2_X1 U18184 ( .A(n12588), .B(n13503), .ZN(n12592) );
  XNOR2_X1 U18185 ( .A(n13458), .B(n3666), .ZN(n12590) );
  XNOR2_X1 U18186 ( .A(n13061), .B(n12589), .ZN(n13324) );
  XNOR2_X1 U18187 ( .A(n12590), .B(n13324), .ZN(n12591) );
  INV_X1 U18188 ( .A(n13803), .ZN(n14297) );
  XNOR2_X1 U18189 ( .A(n12594), .B(n12595), .ZN(n13471) );
  XNOR2_X1 U18190 ( .A(n12833), .B(n13471), .ZN(n12599) );
  XNOR2_X1 U18191 ( .A(n12787), .B(n13231), .ZN(n12597) );
  XNOR2_X1 U18192 ( .A(n13450), .B(n21537), .ZN(n12596) );
  XNOR2_X1 U18193 ( .A(n12597), .B(n12596), .ZN(n12598) );
  XNOR2_X1 U18194 ( .A(n12599), .B(n12598), .ZN(n12607) );
  XNOR2_X1 U18195 ( .A(n12760), .B(n1215), .ZN(n12601) );
  XNOR2_X1 U18196 ( .A(n12601), .B(n12600), .ZN(n12602) );
  XNOR2_X1 U18197 ( .A(n12817), .B(n13396), .ZN(n13494) );
  XNOR2_X1 U18198 ( .A(n12602), .B(n13494), .ZN(n12606) );
  XNOR2_X1 U18199 ( .A(n12603), .B(n13048), .ZN(n12604) );
  XNOR2_X1 U18200 ( .A(n12604), .B(n12813), .ZN(n12605) );
  XNOR2_X1 U18201 ( .A(n13038), .B(n12609), .ZN(n12613) );
  XNOR2_X1 U18202 ( .A(n13432), .B(n13337), .ZN(n12611) );
  XNOR2_X1 U18203 ( .A(n12776), .B(n1119), .ZN(n12610) );
  XNOR2_X1 U18204 ( .A(n12611), .B(n12610), .ZN(n12612) );
  XNOR2_X1 U18205 ( .A(n12613), .B(n12612), .ZN(n14293) );
  AOI22_X1 U18206 ( .A1(n12614), .A2(n14298), .B1(n14292), .B2(n14293), .ZN(
        n12625) );
  XNOR2_X1 U18207 ( .A(n13418), .B(n1928), .ZN(n12615) );
  XNOR2_X1 U18208 ( .A(n13067), .B(n1906), .ZN(n13329) );
  XNOR2_X1 U18209 ( .A(n13329), .B(n12615), .ZN(n12618) );
  XNOR2_X1 U18210 ( .A(n13479), .B(n12616), .ZN(n12617) );
  INV_X1 U18212 ( .A(n14292), .ZN(n13697) );
  OAI22_X1 U18213 ( .A1(n14297), .A2(n14293), .B1(n14295), .B2(n13697), .ZN(
        n12623) );
  XNOR2_X1 U18214 ( .A(n12722), .B(n13386), .ZN(n13490) );
  XNOR2_X1 U18215 ( .A(n13556), .B(n13043), .ZN(n13350) );
  XNOR2_X1 U18216 ( .A(n13490), .B(n13350), .ZN(n12622) );
  XNOR2_X1 U18217 ( .A(n13245), .B(n3049), .ZN(n12619) );
  XNOR2_X1 U18218 ( .A(n12620), .B(n12619), .ZN(n12621) );
  XNOR2_X1 U18219 ( .A(n12622), .B(n12621), .ZN(n13306) );
  NAND2_X1 U18220 ( .A1(n12623), .A2(n14291), .ZN(n12624) );
  AND2_X1 U18221 ( .A1(n3315), .A2(n15094), .ZN(n12627) );
  NOR2_X1 U18222 ( .A1(n14578), .A2(n3315), .ZN(n12626) );
  AOI22_X1 U18223 ( .A1(n15095), .A2(n12627), .B1(n12626), .B2(n14903), .ZN(
        n12628) );
  NAND2_X1 U18224 ( .A1(n12629), .A2(n12628), .ZN(n16527) );
  INV_X1 U18225 ( .A(n16527), .ZN(n12630) );
  XNOR2_X1 U18226 ( .A(n12631), .B(n12630), .ZN(n13130) );
  XNOR2_X1 U18227 ( .A(n1885), .B(n3423), .ZN(n12633) );
  XNOR2_X1 U18228 ( .A(n13220), .B(n12633), .ZN(n12636) );
  XNOR2_X1 U18229 ( .A(n12637), .B(n13121), .ZN(n13247) );
  XNOR2_X1 U18230 ( .A(n13247), .B(n12638), .ZN(n12643) );
  INV_X1 U18231 ( .A(n13371), .ZN(n12639) );
  XNOR2_X1 U18232 ( .A(n1905), .B(n12639), .ZN(n12641) );
  XNOR2_X1 U18233 ( .A(n12495), .B(n26214), .ZN(n12640) );
  XNOR2_X1 U18234 ( .A(n12641), .B(n12640), .ZN(n12642) );
  XNOR2_X1 U18235 ( .A(n12746), .B(n12644), .ZN(n13224) );
  INV_X1 U18236 ( .A(n13224), .ZN(n12647) );
  INV_X1 U18237 ( .A(n12881), .ZN(n12645) );
  XNOR2_X1 U18238 ( .A(n13539), .B(n12645), .ZN(n12646) );
  XNOR2_X1 U18239 ( .A(n12647), .B(n12646), .ZN(n12651) );
  XNOR2_X1 U18240 ( .A(n13404), .B(n3211), .ZN(n12649) );
  XNOR2_X1 U18241 ( .A(n12649), .B(n12648), .ZN(n12650) );
  XNOR2_X1 U18242 ( .A(n12651), .B(n12650), .ZN(n13851) );
  INV_X1 U18243 ( .A(n13851), .ZN(n14176) );
  MUX2_X1 U18244 ( .A(n14177), .B(n14181), .S(n14176), .Z(n12673) );
  INV_X1 U18245 ( .A(n13227), .ZN(n12729) );
  XNOR2_X1 U18246 ( .A(n12729), .B(n13231), .ZN(n13096) );
  XNOR2_X1 U18247 ( .A(n12652), .B(n13096), .ZN(n12656) );
  XNOR2_X1 U18248 ( .A(n13567), .B(n2889), .ZN(n12653) );
  XNOR2_X1 U18249 ( .A(n12654), .B(n12653), .ZN(n12655) );
  XNOR2_X1 U18250 ( .A(n12657), .B(n12854), .ZN(n12659) );
  XNOR2_X1 U18251 ( .A(n12659), .B(n13243), .ZN(n12663) );
  XNOR2_X1 U18252 ( .A(n13386), .B(n13556), .ZN(n12661) );
  XNOR2_X1 U18253 ( .A(n4670), .B(n24897), .ZN(n12660) );
  XNOR2_X1 U18254 ( .A(n12661), .B(n12660), .ZN(n12662) );
  XNOR2_X1 U18255 ( .A(n12663), .B(n12662), .ZN(n13753) );
  NAND2_X1 U18256 ( .A1(n5693), .A2(n14451), .ZN(n12671) );
  INV_X1 U18257 ( .A(n12985), .ZN(n12664) );
  XNOR2_X1 U18258 ( .A(n13236), .B(n12664), .ZN(n12666) );
  XNOR2_X1 U18259 ( .A(n13338), .B(n13109), .ZN(n12665) );
  XNOR2_X1 U18260 ( .A(n12665), .B(n12666), .ZN(n12670) );
  XNOR2_X1 U18261 ( .A(n13359), .B(n13337), .ZN(n12668) );
  XNOR2_X1 U18262 ( .A(n13191), .B(n2960), .ZN(n12667) );
  XNOR2_X1 U18263 ( .A(n12668), .B(n12667), .ZN(n12669) );
  XNOR2_X1 U18264 ( .A(n12670), .B(n12669), .ZN(n14178) );
  OAI21_X1 U18265 ( .B1(n12671), .B2(n14176), .A(n13932), .ZN(n12672) );
  XNOR2_X1 U18266 ( .A(n13230), .B(n2527), .ZN(n12675) );
  INV_X1 U18267 ( .A(n12787), .ZN(n12674) );
  XNOR2_X1 U18268 ( .A(n12675), .B(n12674), .ZN(n12676) );
  XNOR2_X1 U18269 ( .A(n12676), .B(n13565), .ZN(n12679) );
  XNOR2_X1 U18270 ( .A(n13451), .B(n12677), .ZN(n12678) );
  XNOR2_X1 U18271 ( .A(n12678), .B(n13380), .ZN(n12983) );
  XNOR2_X1 U18272 ( .A(n12679), .B(n12983), .ZN(n12711) );
  XNOR2_X1 U18273 ( .A(n12760), .B(n28327), .ZN(n12680) );
  XNOR2_X1 U18274 ( .A(n29140), .B(n12681), .ZN(n12682) );
  XNOR2_X1 U18275 ( .A(n12683), .B(n12682), .ZN(n12712) );
  XNOR2_X1 U18276 ( .A(n13150), .B(n12684), .ZN(n13388) );
  XNOR2_X1 U18277 ( .A(n12685), .B(n13388), .ZN(n12690) );
  XNOR2_X1 U18278 ( .A(n13488), .B(n72), .ZN(n12687) );
  XNOR2_X1 U18279 ( .A(n12688), .B(n12687), .ZN(n12689) );
  XNOR2_X1 U18280 ( .A(n12690), .B(n12689), .ZN(n13967) );
  XNOR2_X1 U18282 ( .A(n13370), .B(n13137), .ZN(n13000) );
  XNOR2_X1 U18283 ( .A(n13000), .B(n12691), .ZN(n12695) );
  XNOR2_X1 U18284 ( .A(n1857), .B(n13420), .ZN(n12693) );
  XNOR2_X1 U18285 ( .A(n13482), .B(n27462), .ZN(n12692) );
  XNOR2_X1 U18286 ( .A(n12693), .B(n12692), .ZN(n12694) );
  XNOR2_X1 U18287 ( .A(n12696), .B(n12697), .ZN(n13363) );
  XNOR2_X1 U18288 ( .A(n12698), .B(n13363), .ZN(n12703) );
  XNOR2_X1 U18289 ( .A(n12776), .B(n2325), .ZN(n12700) );
  XNOR2_X1 U18290 ( .A(n12701), .B(n12700), .ZN(n12702) );
  OAI21_X1 U18291 ( .B1(n14463), .B2(n13967), .A(n12704), .ZN(n12715) );
  INV_X1 U18292 ( .A(n13967), .ZN(n14456) );
  NOR2_X1 U18293 ( .A1(n14455), .A2(n14456), .ZN(n12714) );
  XNOR2_X1 U18294 ( .A(n13406), .B(n13401), .ZN(n12706) );
  XNOR2_X1 U18295 ( .A(n12705), .B(n12706), .ZN(n12710) );
  XNOR2_X1 U18296 ( .A(n13208), .B(n3697), .ZN(n12708) );
  XNOR2_X1 U18297 ( .A(n12707), .B(n12708), .ZN(n12709) );
  NOR2_X1 U18298 ( .A1(n12711), .A2(n427), .ZN(n12713) );
  XNOR2_X1 U18299 ( .A(n13035), .B(n13109), .ZN(n12716) );
  XNOR2_X1 U18300 ( .A(n12717), .B(n12716), .ZN(n12720) );
  XNOR2_X1 U18301 ( .A(n13113), .B(n13364), .ZN(n13293) );
  XNOR2_X1 U18302 ( .A(n12808), .B(n2602), .ZN(n12718) );
  XNOR2_X1 U18303 ( .A(n12718), .B(n13293), .ZN(n12719) );
  INV_X1 U18304 ( .A(n13933), .ZN(n14465) );
  XNOR2_X1 U18305 ( .A(n13346), .B(n12721), .ZN(n12726) );
  XNOR2_X1 U18306 ( .A(n12722), .B(n12723), .ZN(n12822) );
  XNOR2_X1 U18307 ( .A(n13263), .B(n27452), .ZN(n12724) );
  XNOR2_X1 U18308 ( .A(n12822), .B(n12724), .ZN(n12725) );
  INV_X1 U18309 ( .A(n14469), .ZN(n14185) );
  XNOR2_X1 U18310 ( .A(n12595), .B(n13159), .ZN(n12728) );
  XNOR2_X1 U18311 ( .A(n12980), .B(n13285), .ZN(n12727) );
  XNOR2_X1 U18312 ( .A(n12727), .B(n12728), .ZN(n12733) );
  XNOR2_X1 U18313 ( .A(n12790), .B(n12729), .ZN(n12731) );
  XNOR2_X1 U18314 ( .A(n13448), .B(n3482), .ZN(n12730) );
  XNOR2_X1 U18315 ( .A(n12731), .B(n12730), .ZN(n12732) );
  XNOR2_X1 U18316 ( .A(n12732), .B(n12733), .ZN(n12743) );
  NAND2_X1 U18317 ( .A1(n14185), .A2(n12743), .ZN(n12744) );
  XNOR2_X1 U18318 ( .A(n12894), .B(n13080), .ZN(n13280) );
  INV_X1 U18319 ( .A(n13280), .ZN(n12737) );
  INV_X1 U18320 ( .A(n12734), .ZN(n12736) );
  XNOR2_X1 U18321 ( .A(n12736), .B(n12762), .ZN(n13318) );
  XNOR2_X1 U18322 ( .A(n12737), .B(n13318), .ZN(n12742) );
  XNOR2_X1 U18323 ( .A(n12738), .B(n2522), .ZN(n12740) );
  XNOR2_X1 U18324 ( .A(n13445), .B(n12817), .ZN(n12739) );
  XNOR2_X1 U18325 ( .A(n12740), .B(n12739), .ZN(n12741) );
  XNOR2_X1 U18326 ( .A(n12742), .B(n12741), .ZN(n13677) );
  INV_X1 U18327 ( .A(n13677), .ZN(n14184) );
  XNOR2_X1 U18330 ( .A(n13025), .B(n2984), .ZN(n12748) );
  XNOR2_X1 U18331 ( .A(n12747), .B(n29064), .ZN(n12839) );
  XNOR2_X1 U18332 ( .A(n12839), .B(n12748), .ZN(n12751) );
  XNOR2_X1 U18333 ( .A(n13325), .B(n12749), .ZN(n12750) );
  XNOR2_X1 U18334 ( .A(n12750), .B(n12751), .ZN(n13678) );
  INV_X1 U18335 ( .A(n12752), .ZN(n12753) );
  XNOR2_X1 U18336 ( .A(n13374), .B(n13328), .ZN(n12757) );
  XNOR2_X1 U18337 ( .A(n12830), .B(n13272), .ZN(n12755) );
  XNOR2_X1 U18338 ( .A(n13118), .B(n2385), .ZN(n12754) );
  XNOR2_X1 U18339 ( .A(n12755), .B(n12754), .ZN(n12756) );
  NAND3_X1 U18340 ( .A1(n14182), .A2(n14469), .A3(n14464), .ZN(n12758) );
  XNOR2_X1 U18341 ( .A(n12760), .B(n13278), .ZN(n13496) );
  INV_X1 U18342 ( .A(n13496), .ZN(n12761) );
  XNOR2_X1 U18343 ( .A(n12761), .B(n13277), .ZN(n12767) );
  XNOR2_X1 U18344 ( .A(n12762), .B(n2306), .ZN(n12764) );
  XNOR2_X1 U18345 ( .A(n12764), .B(n12763), .ZN(n12765) );
  XNOR2_X1 U18346 ( .A(n12765), .B(n13167), .ZN(n12766) );
  XNOR2_X1 U18348 ( .A(n12768), .B(n13405), .ZN(n12769) );
  XNOR2_X1 U18349 ( .A(n13501), .B(n12769), .ZN(n12773) );
  XNOR2_X1 U18350 ( .A(n13543), .B(n12931), .ZN(n12771) );
  XNOR2_X1 U18351 ( .A(n13209), .B(n3109), .ZN(n12770) );
  XNOR2_X1 U18352 ( .A(n12771), .B(n12770), .ZN(n12772) );
  XNOR2_X1 U18353 ( .A(n12773), .B(n12772), .ZN(n14497) );
  XNOR2_X1 U18355 ( .A(n13290), .B(n12775), .ZN(n12779) );
  XNOR2_X1 U18356 ( .A(n12919), .B(n2996), .ZN(n12777) );
  XNOR2_X1 U18357 ( .A(n12777), .B(n13513), .ZN(n12778) );
  XNOR2_X1 U18358 ( .A(n12780), .B(n13414), .ZN(n12782) );
  INV_X1 U18359 ( .A(n12944), .ZN(n12781) );
  XNOR2_X1 U18360 ( .A(n12781), .B(n12782), .ZN(n12786) );
  INV_X1 U18361 ( .A(n3134), .ZN(n27643) );
  XNOR2_X1 U18362 ( .A(n12783), .B(n27643), .ZN(n12784) );
  XNOR2_X1 U18363 ( .A(n12784), .B(n13274), .ZN(n12785) );
  XNOR2_X1 U18364 ( .A(n12786), .B(n12785), .ZN(n13672) );
  INV_X1 U18365 ( .A(n13672), .ZN(n14491) );
  NAND2_X1 U18366 ( .A1(n14154), .A2(n14491), .ZN(n12795) );
  INV_X1 U18367 ( .A(n12949), .ZN(n13472) );
  XNOR2_X1 U18368 ( .A(n13472), .B(n12789), .ZN(n12794) );
  XNOR2_X1 U18369 ( .A(n12790), .B(n3554), .ZN(n12791) );
  XNOR2_X1 U18370 ( .A(n12791), .B(n12792), .ZN(n12793) );
  MUX2_X1 U18371 ( .A(n12796), .B(n12795), .S(n14492), .Z(n12805) );
  XNOR2_X1 U18372 ( .A(n13265), .B(n13485), .ZN(n12798) );
  XNOR2_X1 U18373 ( .A(n12798), .B(n12797), .ZN(n12803) );
  XNOR2_X1 U18374 ( .A(n12799), .B(n13262), .ZN(n12801) );
  XNOR2_X1 U18375 ( .A(n13488), .B(n2465), .ZN(n12800) );
  XNOR2_X1 U18376 ( .A(n12801), .B(n12800), .ZN(n12802) );
  XNOR2_X1 U18377 ( .A(n12803), .B(n12802), .ZN(n13855) );
  INV_X1 U18378 ( .A(n13855), .ZN(n14493) );
  OAI21_X1 U18379 ( .B1(n4549), .B2(n15101), .A(n549), .ZN(n12891) );
  INV_X1 U18380 ( .A(n13549), .ZN(n12806) );
  XNOR2_X1 U18381 ( .A(n12806), .B(n12807), .ZN(n12812) );
  XNOR2_X1 U18382 ( .A(n12808), .B(n2544), .ZN(n12810) );
  INV_X1 U18383 ( .A(n12809), .ZN(n13342) );
  XNOR2_X1 U18384 ( .A(n13342), .B(n12810), .ZN(n12811) );
  INV_X1 U18385 ( .A(n13048), .ZN(n12814) );
  XNOR2_X1 U18386 ( .A(n12814), .B(n12813), .ZN(n13314) );
  XNOR2_X1 U18387 ( .A(n13314), .B(n12815), .ZN(n12821) );
  XNOR2_X1 U18388 ( .A(n12816), .B(n13493), .ZN(n12819) );
  XNOR2_X1 U18389 ( .A(n12817), .B(n2353), .ZN(n12818) );
  XNOR2_X1 U18390 ( .A(n12819), .B(n12818), .ZN(n12820) );
  XNOR2_X1 U18391 ( .A(n13557), .B(n12913), .ZN(n12824) );
  XNOR2_X1 U18392 ( .A(n13484), .B(n3662), .ZN(n12823) );
  XNOR2_X1 U18393 ( .A(n12824), .B(n12823), .ZN(n12825) );
  XNOR2_X1 U18394 ( .A(n12827), .B(n5059), .ZN(n12828) );
  XNOR2_X1 U18395 ( .A(n13118), .B(n12830), .ZN(n12831) );
  INV_X1 U18396 ( .A(n13329), .ZN(n12832) );
  XNOR2_X1 U18397 ( .A(n13563), .B(n12595), .ZN(n12836) );
  XNOR2_X1 U18398 ( .A(n13473), .B(n26909), .ZN(n12835) );
  XNOR2_X1 U18399 ( .A(n12836), .B(n12835), .ZN(n12837) );
  INV_X1 U18400 ( .A(n12839), .ZN(n12840) );
  XNOR2_X1 U18401 ( .A(n12840), .B(n13324), .ZN(n12845) );
  XNOR2_X1 U18402 ( .A(n12841), .B(n13459), .ZN(n12843) );
  XNOR2_X1 U18403 ( .A(n13504), .B(n2350), .ZN(n12842) );
  XNOR2_X1 U18404 ( .A(n12843), .B(n12842), .ZN(n12844) );
  NAND3_X1 U18405 ( .A1(n4549), .A2(n15422), .A3(n14575), .ZN(n12890) );
  XNOR2_X1 U18406 ( .A(n13331), .B(n12849), .ZN(n12850) );
  INV_X1 U18407 ( .A(n12851), .ZN(n13248) );
  XNOR2_X1 U18408 ( .A(n13150), .B(n3219), .ZN(n12852) );
  XNOR2_X1 U18409 ( .A(n13553), .B(n12852), .ZN(n12853) );
  XNOR2_X1 U18410 ( .A(n13246), .B(n12853), .ZN(n12857) );
  XNOR2_X1 U18411 ( .A(n12913), .B(n13245), .ZN(n12855) );
  XNOR2_X1 U18412 ( .A(n12855), .B(n12854), .ZN(n12856) );
  XNOR2_X1 U18413 ( .A(n12857), .B(n12856), .ZN(n14207) );
  INV_X1 U18414 ( .A(n13036), .ZN(n12858) );
  XNOR2_X1 U18415 ( .A(n13341), .B(n12858), .ZN(n13240) );
  XNOR2_X1 U18416 ( .A(n13338), .B(n13432), .ZN(n12859) );
  XNOR2_X1 U18417 ( .A(n13240), .B(n12859), .ZN(n12864) );
  XNOR2_X1 U18418 ( .A(n12860), .B(n13191), .ZN(n12924) );
  INV_X1 U18419 ( .A(n1161), .ZN(n27730) );
  XNOR2_X1 U18420 ( .A(n12861), .B(n27730), .ZN(n12862) );
  XNOR2_X1 U18421 ( .A(n12924), .B(n12862), .ZN(n12863) );
  XNOR2_X1 U18422 ( .A(n12864), .B(n12863), .ZN(n14433) );
  MUX2_X1 U18423 ( .A(n1841), .B(n14207), .S(n14433), .Z(n12888) );
  XNOR2_X1 U18424 ( .A(n13018), .B(n1179), .ZN(n12865) );
  XNOR2_X1 U18425 ( .A(n12868), .B(n12867), .ZN(n12892) );
  XNOR2_X1 U18426 ( .A(n13444), .B(n13525), .ZN(n12869) );
  XNOR2_X1 U18427 ( .A(n12869), .B(n13051), .ZN(n13221) );
  INV_X1 U18428 ( .A(n13221), .ZN(n12870) );
  XNOR2_X2 U18429 ( .A(n12871), .B(n12870), .ZN(n14438) );
  XNOR2_X1 U18430 ( .A(n12872), .B(n13447), .ZN(n12874) );
  INV_X1 U18431 ( .A(n13229), .ZN(n12873) );
  XNOR2_X1 U18432 ( .A(n13450), .B(n25044), .ZN(n12875) );
  XNOR2_X1 U18433 ( .A(n12876), .B(n12875), .ZN(n12877) );
  XNOR2_X1 U18434 ( .A(n12879), .B(n3527), .ZN(n12880) );
  XNOR2_X1 U18435 ( .A(n12880), .B(n29494), .ZN(n12882) );
  XNOR2_X1 U18436 ( .A(n12881), .B(n13459), .ZN(n12929) );
  XNOR2_X1 U18437 ( .A(n12883), .B(n13075), .ZN(n12884) );
  INV_X1 U18439 ( .A(n15423), .ZN(n14577) );
  NAND3_X1 U18440 ( .A1(n15102), .A2(n15105), .A3(n14577), .ZN(n12889) );
  XNOR2_X1 U18441 ( .A(n13167), .B(n13493), .ZN(n12893) );
  XNOR2_X1 U18442 ( .A(n12892), .B(n12893), .ZN(n12898) );
  XNOR2_X1 U18443 ( .A(n13166), .B(n1225), .ZN(n12896) );
  XNOR2_X1 U18444 ( .A(n12894), .B(n13444), .ZN(n12895) );
  XNOR2_X1 U18445 ( .A(n12895), .B(n12896), .ZN(n12897) );
  XNOR2_X1 U18446 ( .A(n13179), .B(n13447), .ZN(n12900) );
  XNOR2_X1 U18447 ( .A(n12899), .B(n12900), .ZN(n12903) );
  XNOR2_X1 U18448 ( .A(n13567), .B(n3083), .ZN(n12901) );
  XNOR2_X1 U18449 ( .A(n12904), .B(n12905), .ZN(n12910) );
  XNOR2_X1 U18450 ( .A(n12495), .B(n2389), .ZN(n12907) );
  XNOR2_X1 U18451 ( .A(n12908), .B(n12907), .ZN(n12909) );
  MUX2_X1 U18452 ( .A(n14082), .B(n14084), .S(n14287), .Z(n12928) );
  INV_X1 U18453 ( .A(n12913), .ZN(n12915) );
  XNOR2_X1 U18454 ( .A(n12914), .B(n12915), .ZN(n12917) );
  XNOR2_X1 U18455 ( .A(n13484), .B(n3116), .ZN(n12916) );
  XNOR2_X1 U18456 ( .A(n12917), .B(n12916), .ZN(n12918) );
  NOR2_X1 U18457 ( .A1(n28625), .A2(n14282), .ZN(n12927) );
  XNOR2_X1 U18459 ( .A(n12921), .B(n12920), .ZN(n12926) );
  INV_X1 U18460 ( .A(n3463), .ZN(n12922) );
  XNOR2_X1 U18461 ( .A(n13511), .B(n12922), .ZN(n12923) );
  XNOR2_X1 U18462 ( .A(n12924), .B(n12923), .ZN(n12925) );
  XNOR2_X1 U18463 ( .A(n12926), .B(n12925), .ZN(n14083) );
  XNOR2_X1 U18464 ( .A(n12929), .B(n12930), .ZN(n12935) );
  XNOR2_X1 U18465 ( .A(n12931), .B(n3710), .ZN(n12932) );
  XNOR2_X1 U18466 ( .A(n12933), .B(n12932), .ZN(n12934) );
  XNOR2_X1 U18467 ( .A(n12935), .B(n12934), .ZN(n14286) );
  INV_X1 U18468 ( .A(n14084), .ZN(n14281) );
  AND2_X1 U18471 ( .A1(n14106), .A2(n14105), .ZN(n14234) );
  NAND2_X1 U18472 ( .A1(n14234), .A2(n14102), .ZN(n12941) );
  BUF_X2 U18473 ( .A(n13606), .Z(n14230) );
  NAND2_X1 U18474 ( .A1(n12938), .A2(n14230), .ZN(n12940) );
  NAND2_X1 U18475 ( .A1(n14102), .A2(n14107), .ZN(n12939) );
  XNOR2_X1 U18478 ( .A(n13141), .B(n12943), .ZN(n12947) );
  XNOR2_X1 U18479 ( .A(n13419), .B(n1184), .ZN(n12945) );
  XNOR2_X1 U18480 ( .A(n12944), .B(n12945), .ZN(n12946) );
  XNOR2_X1 U18481 ( .A(n13448), .B(n12948), .ZN(n13379) );
  XNOR2_X1 U18482 ( .A(n12949), .B(n13379), .ZN(n12953) );
  XNOR2_X1 U18483 ( .A(n13230), .B(n3493), .ZN(n12951) );
  XNOR2_X1 U18484 ( .A(n12978), .B(n13055), .ZN(n12950) );
  XNOR2_X1 U18485 ( .A(n12951), .B(n12950), .ZN(n12952) );
  XNOR2_X1 U18486 ( .A(n12954), .B(n13445), .ZN(n13394) );
  XNOR2_X1 U18487 ( .A(n13394), .B(n13496), .ZN(n12959) );
  XNOR2_X1 U18488 ( .A(n13020), .B(n13048), .ZN(n12957) );
  XNOR2_X1 U18489 ( .A(n12955), .B(n3212), .ZN(n12956) );
  XNOR2_X1 U18490 ( .A(n12956), .B(n12957), .ZN(n12958) );
  INV_X1 U18491 ( .A(n13061), .ZN(n12960) );
  XNOR2_X1 U18492 ( .A(n13028), .B(n1123), .ZN(n12961) );
  XNOR2_X1 U18493 ( .A(n12962), .B(n12961), .ZN(n12964) );
  XNOR2_X1 U18494 ( .A(n13428), .B(n12965), .ZN(n13389) );
  XNOR2_X1 U18495 ( .A(n12966), .B(n13389), .ZN(n12970) );
  XNOR2_X1 U18496 ( .A(n13008), .B(n13043), .ZN(n12968) );
  XNOR2_X1 U18497 ( .A(n13488), .B(n3622), .ZN(n12967) );
  XNOR2_X1 U18498 ( .A(n12968), .B(n12967), .ZN(n12969) );
  XNOR2_X1 U18499 ( .A(n13039), .B(n135), .ZN(n12971) );
  XNOR2_X1 U18500 ( .A(n12985), .B(n12971), .ZN(n12973) );
  XNOR2_X1 U18501 ( .A(n12973), .B(n12972), .ZN(n12975) );
  XNOR2_X1 U18502 ( .A(n13513), .B(n13433), .ZN(n12974) );
  NAND2_X1 U18503 ( .A1(n12976), .A2(n14365), .ZN(n14370) );
  XNOR2_X1 U18504 ( .A(n12978), .B(n3276), .ZN(n12979) );
  XNOR2_X1 U18505 ( .A(n12979), .B(n28587), .ZN(n12982) );
  XNOR2_X1 U18506 ( .A(n12980), .B(n13562), .ZN(n12981) );
  XNOR2_X1 U18507 ( .A(n12982), .B(n12981), .ZN(n12984) );
  XNOR2_X1 U18508 ( .A(n12985), .B(n2598), .ZN(n12986) );
  XNOR2_X1 U18509 ( .A(n13341), .B(n13436), .ZN(n13545) );
  XNOR2_X1 U18510 ( .A(n12986), .B(n13545), .ZN(n12989) );
  XNOR2_X1 U18511 ( .A(n13363), .B(n12987), .ZN(n12988) );
  XNOR2_X1 U18512 ( .A(n12989), .B(n12988), .ZN(n13832) );
  MUX2_X1 U18513 ( .A(n12992), .B(n12991), .S(n12990), .Z(n12993) );
  NAND2_X1 U18514 ( .A1(n12994), .A2(n12993), .ZN(n12997) );
  INV_X1 U18515 ( .A(n12995), .ZN(n12996) );
  NAND2_X1 U18516 ( .A1(n12997), .A2(n12996), .ZN(n12999) );
  INV_X1 U18517 ( .A(n13413), .ZN(n12998) );
  XNOR2_X1 U18518 ( .A(n12998), .B(n12999), .ZN(n13530) );
  XNOR2_X1 U18519 ( .A(n13000), .B(n13530), .ZN(n13004) );
  XNOR2_X1 U18520 ( .A(n1857), .B(n13478), .ZN(n13002) );
  XNOR2_X1 U18521 ( .A(n13270), .B(n3414), .ZN(n13001) );
  XNOR2_X1 U18522 ( .A(n13002), .B(n13001), .ZN(n13003) );
  NAND3_X1 U18523 ( .A1(n13829), .A2(n13832), .A3(n14278), .ZN(n13024) );
  XNOR2_X1 U18524 ( .A(n13005), .B(n13263), .ZN(n13007) );
  INV_X1 U18525 ( .A(n13348), .ZN(n13006) );
  XNOR2_X1 U18526 ( .A(n13006), .B(n13265), .ZN(n13554) );
  XNOR2_X1 U18527 ( .A(n13150), .B(n2946), .ZN(n13009) );
  XNOR2_X1 U18528 ( .A(n13010), .B(n13009), .ZN(n13011) );
  XNOR2_X1 U18529 ( .A(n13013), .B(n13014), .ZN(n13016) );
  XNOR2_X1 U18530 ( .A(n13016), .B(n13015), .ZN(n13023) );
  INV_X1 U18531 ( .A(n13017), .ZN(n13019) );
  XNOR2_X1 U18532 ( .A(n13018), .B(n13019), .ZN(n13393) );
  XNOR2_X1 U18533 ( .A(n13020), .B(n3462), .ZN(n13021) );
  XNOR2_X1 U18534 ( .A(n13393), .B(n13021), .ZN(n13022) );
  NAND2_X1 U18535 ( .A1(n14362), .A2(n14358), .ZN(n14275) );
  XNOR2_X1 U18536 ( .A(n13025), .B(n29495), .ZN(n13026) );
  XNOR2_X1 U18537 ( .A(n13027), .B(n13026), .ZN(n13031) );
  XNOR2_X1 U18538 ( .A(n13028), .B(n3660), .ZN(n13029) );
  XNOR2_X1 U18539 ( .A(n13456), .B(n13029), .ZN(n13030) );
  XNOR2_X1 U18540 ( .A(n13031), .B(n13030), .ZN(n14360) );
  OAI21_X1 U18541 ( .B1(n14275), .B2(n14360), .A(n13032), .ZN(n13033) );
  XNOR2_X1 U18542 ( .A(n13035), .B(n13034), .ZN(n13340) );
  XNOR2_X1 U18543 ( .A(n13036), .B(n13360), .ZN(n13037) );
  XNOR2_X1 U18544 ( .A(n13340), .B(n13037), .ZN(n13041) );
  XNOR2_X1 U18545 ( .A(n13039), .B(n1887), .ZN(n13040) );
  INV_X1 U18546 ( .A(n13490), .ZN(n13042) );
  XNOR2_X1 U18547 ( .A(n13346), .B(n13042), .ZN(n13047) );
  XNOR2_X1 U18548 ( .A(n13043), .B(n13262), .ZN(n13045) );
  XNOR2_X1 U18549 ( .A(n13101), .B(n3451), .ZN(n13044) );
  XNOR2_X1 U18550 ( .A(n13045), .B(n13044), .ZN(n13046) );
  XNOR2_X1 U18551 ( .A(n13170), .B(n3196), .ZN(n13049) );
  XNOR2_X1 U18552 ( .A(n13049), .B(n13048), .ZN(n13050) );
  XNOR2_X1 U18553 ( .A(n13050), .B(n13318), .ZN(n13053) );
  XNOR2_X1 U18554 ( .A(n13494), .B(n13051), .ZN(n13052) );
  XNOR2_X1 U18555 ( .A(n13353), .B(n13471), .ZN(n13059) );
  XNOR2_X1 U18556 ( .A(n13097), .B(n13175), .ZN(n13057) );
  XNOR2_X1 U18557 ( .A(n13055), .B(n3385), .ZN(n13056) );
  XNOR2_X1 U18558 ( .A(n13057), .B(n13056), .ZN(n13058) );
  XNOR2_X1 U18559 ( .A(n13059), .B(n13058), .ZN(n13824) );
  XNOR2_X1 U18560 ( .A(n13325), .B(n13503), .ZN(n13065) );
  XNOR2_X1 U18561 ( .A(n13061), .B(n13075), .ZN(n13063) );
  XNOR2_X1 U18562 ( .A(n13209), .B(n26680), .ZN(n13062) );
  XNOR2_X1 U18563 ( .A(n13063), .B(n13062), .ZN(n13064) );
  INV_X1 U18564 ( .A(n13369), .ZN(n13066) );
  XNOR2_X1 U18565 ( .A(n13066), .B(n13067), .ZN(n13068) );
  XNOR2_X1 U18566 ( .A(n13328), .B(n13068), .ZN(n13072) );
  XNOR2_X1 U18567 ( .A(n429), .B(n25992), .ZN(n13070) );
  XNOR2_X1 U18568 ( .A(n13479), .B(n13070), .ZN(n13071) );
  OAI211_X1 U18569 ( .C1(n14351), .C2(n13826), .A(n4893), .B(n14354), .ZN(
        n13073) );
  INV_X1 U18570 ( .A(n13073), .ZN(n13074) );
  AOI21_X2 U18571 ( .B1(n14015), .B2(n14350), .A(n13074), .ZN(n15077) );
  XNOR2_X1 U18572 ( .A(n13298), .B(n13075), .ZN(n13077) );
  XNOR2_X1 U18573 ( .A(n13208), .B(n3644), .ZN(n13076) );
  XNOR2_X1 U18574 ( .A(n13077), .B(n13076), .ZN(n13079) );
  XNOR2_X1 U18575 ( .A(n13224), .B(n13322), .ZN(n13078) );
  XNOR2_X1 U18576 ( .A(n13078), .B(n13079), .ZN(n14342) );
  XNOR2_X1 U18577 ( .A(n13166), .B(n13080), .ZN(n13092) );
  NAND2_X1 U18578 ( .A1(n13082), .A2(n13081), .ZN(n13089) );
  NAND2_X1 U18579 ( .A1(n13087), .A2(n13083), .ZN(n13085) );
  OAI211_X1 U18580 ( .C1(n13087), .C2(n13086), .A(n13085), .B(n13084), .ZN(
        n13088) );
  NAND2_X1 U18581 ( .A1(n13089), .A2(n13088), .ZN(n13090) );
  XNOR2_X1 U18582 ( .A(n13090), .B(n2541), .ZN(n13091) );
  XNOR2_X1 U18583 ( .A(n13092), .B(n13091), .ZN(n13093) );
  INV_X1 U18584 ( .A(n13095), .ZN(n13354) );
  XNOR2_X1 U18585 ( .A(n13354), .B(n13096), .ZN(n13100) );
  XNOR2_X1 U18586 ( .A(n13179), .B(n13285), .ZN(n13099) );
  XNOR2_X1 U18587 ( .A(n13097), .B(n1911), .ZN(n13098) );
  INV_X1 U18589 ( .A(n13101), .ZN(n13102) );
  XNOR2_X1 U18590 ( .A(n28603), .B(n13102), .ZN(n13103) );
  XNOR2_X1 U18591 ( .A(n13103), .B(n13347), .ZN(n13107) );
  XNOR2_X1 U18592 ( .A(n13104), .B(n21865), .ZN(n13105) );
  XNOR2_X1 U18593 ( .A(n13243), .B(n13105), .ZN(n13106) );
  XNOR2_X1 U18594 ( .A(n13107), .B(n13106), .ZN(n13842) );
  XNOR2_X1 U18595 ( .A(n13338), .B(n13236), .ZN(n13111) );
  INV_X1 U18596 ( .A(n13190), .ZN(n13108) );
  XNOR2_X1 U18597 ( .A(n13108), .B(n13109), .ZN(n13110) );
  XNOR2_X1 U18598 ( .A(n13111), .B(n13110), .ZN(n13117) );
  INV_X1 U18599 ( .A(n13112), .ZN(n13115) );
  XNOR2_X1 U18600 ( .A(n13113), .B(n2510), .ZN(n13114) );
  XNOR2_X1 U18601 ( .A(n13115), .B(n13114), .ZN(n13116) );
  XNOR2_X1 U18602 ( .A(n13116), .B(n13117), .ZN(n14010) );
  XNOR2_X1 U18603 ( .A(n429), .B(n13533), .ZN(n13120) );
  XNOR2_X1 U18604 ( .A(n13118), .B(n2404), .ZN(n13119) );
  XNOR2_X1 U18605 ( .A(n13120), .B(n13119), .ZN(n13124) );
  XNOR2_X1 U18606 ( .A(n13272), .B(n13121), .ZN(n13122) );
  XNOR2_X1 U18607 ( .A(n13122), .B(n13332), .ZN(n13123) );
  INV_X1 U18608 ( .A(n14342), .ZN(n14135) );
  INV_X1 U18609 ( .A(n14131), .ZN(n14343) );
  NAND2_X1 U18610 ( .A1(n14135), .A2(n14343), .ZN(n13125) );
  MUX2_X1 U18611 ( .A(n14948), .B(n15077), .S(n15073), .Z(n13126) );
  INV_X1 U18612 ( .A(n14874), .ZN(n14572) );
  NAND2_X1 U18613 ( .A1(n13126), .A2(n14572), .ZN(n13127) );
  INV_X1 U18614 ( .A(n14948), .ZN(n15072) );
  XNOR2_X1 U18615 ( .A(n16606), .B(n16476), .ZN(n13129) );
  XNOR2_X1 U18616 ( .A(n13130), .B(n13129), .ZN(n13605) );
  XNOR2_X1 U18617 ( .A(n13539), .B(n29494), .ZN(n13132) );
  XNOR2_X1 U18618 ( .A(n13131), .B(n13132), .ZN(n13135) );
  XNOR2_X1 U18619 ( .A(n13133), .B(n2973), .ZN(n13134) );
  XNOR2_X1 U18620 ( .A(n1906), .B(n13136), .ZN(n13139) );
  XNOR2_X1 U18621 ( .A(n13137), .B(n27105), .ZN(n13138) );
  XNOR2_X1 U18622 ( .A(n13139), .B(n13138), .ZN(n13143) );
  XNOR2_X1 U18623 ( .A(n13140), .B(n13141), .ZN(n13142) );
  XNOR2_X1 U18624 ( .A(n13143), .B(n13142), .ZN(n14061) );
  XNOR2_X1 U18625 ( .A(n13144), .B(n26665), .ZN(n13145) );
  XNOR2_X1 U18626 ( .A(n13145), .B(n13394), .ZN(n13149) );
  XNOR2_X1 U18627 ( .A(n13147), .B(n13146), .ZN(n13148) );
  MUX2_X1 U18628 ( .A(n14325), .B(n14064), .S(n14327), .Z(n13165) );
  XNOR2_X1 U18629 ( .A(n13487), .B(n13389), .ZN(n13154) );
  XNOR2_X1 U18630 ( .A(n13150), .B(n27422), .ZN(n13151) );
  XNOR2_X1 U18631 ( .A(n13152), .B(n13151), .ZN(n13153) );
  XNOR2_X1 U18632 ( .A(n13154), .B(n13153), .ZN(n13653) );
  XNOR2_X1 U18633 ( .A(n13362), .B(n13155), .ZN(n13158) );
  XNOR2_X1 U18634 ( .A(n13337), .B(n3598), .ZN(n13156) );
  XNOR2_X1 U18635 ( .A(n13509), .B(n13156), .ZN(n13157) );
  XNOR2_X1 U18636 ( .A(n13157), .B(n13158), .ZN(n13652) );
  XNOR2_X1 U18637 ( .A(n13474), .B(n13379), .ZN(n13163) );
  XNOR2_X1 U18638 ( .A(n13159), .B(n13380), .ZN(n13161) );
  XNOR2_X1 U18639 ( .A(n12593), .B(n3686), .ZN(n13160) );
  XNOR2_X1 U18640 ( .A(n13161), .B(n13160), .ZN(n13162) );
  XNOR2_X2 U18641 ( .A(n13163), .B(n13162), .ZN(n14328) );
  INV_X1 U18642 ( .A(n15692), .ZN(n15084) );
  XNOR2_X1 U18643 ( .A(n13166), .B(n13167), .ZN(n13169) );
  XNOR2_X1 U18644 ( .A(n13169), .B(n13168), .ZN(n13174) );
  XNOR2_X1 U18645 ( .A(n13170), .B(n13171), .ZN(n13398) );
  XNOR2_X1 U18646 ( .A(n13218), .B(n3336), .ZN(n13172) );
  XNOR2_X1 U18647 ( .A(n13172), .B(n13398), .ZN(n13173) );
  XNOR2_X1 U18648 ( .A(n13174), .B(n13173), .ZN(n14029) );
  XNOR2_X1 U18649 ( .A(n13567), .B(n3321), .ZN(n13176) );
  XNOR2_X1 U18650 ( .A(n13177), .B(n13176), .ZN(n13183) );
  XNOR2_X1 U18651 ( .A(n13178), .B(n13179), .ZN(n13181) );
  XNOR2_X1 U18652 ( .A(n13181), .B(n13180), .ZN(n13182) );
  XNOR2_X1 U18653 ( .A(n13370), .B(n13414), .ZN(n13184) );
  XNOR2_X1 U18654 ( .A(n13535), .B(n13184), .ZN(n13188) );
  XNOR2_X1 U18655 ( .A(n13369), .B(n13420), .ZN(n13186) );
  XNOR2_X1 U18656 ( .A(n13533), .B(n3191), .ZN(n13185) );
  XNOR2_X1 U18657 ( .A(n13186), .B(n13185), .ZN(n13187) );
  MUX2_X1 U18659 ( .A(n14029), .B(n29107), .S(n14031), .Z(n13217) );
  XNOR2_X1 U18660 ( .A(n13360), .B(n730), .ZN(n13189) );
  XNOR2_X1 U18661 ( .A(n13189), .B(n13434), .ZN(n13194) );
  XNOR2_X1 U18662 ( .A(n13190), .B(n13191), .ZN(n13546) );
  XNOR2_X1 U18663 ( .A(n13192), .B(n13546), .ZN(n13193) );
  XNOR2_X1 U18664 ( .A(n13553), .B(n13195), .ZN(n13196) );
  XNOR2_X1 U18665 ( .A(n13197), .B(n13196), .ZN(n13201) );
  XNOR2_X1 U18666 ( .A(n13104), .B(n1246), .ZN(n13199) );
  XNOR2_X1 U18667 ( .A(n13244), .B(n13262), .ZN(n13198) );
  XNOR2_X1 U18668 ( .A(n13199), .B(n13198), .ZN(n13200) );
  XNOR2_X1 U18669 ( .A(n13201), .B(n13200), .ZN(n13917) );
  NAND2_X1 U18670 ( .A1(n13917), .A2(n13793), .ZN(n13215) );
  XNOR2_X1 U18671 ( .A(n13540), .B(n13457), .ZN(n13213) );
  NAND2_X1 U18672 ( .A1(n13206), .A2(n13202), .ZN(n13204) );
  OAI211_X1 U18673 ( .C1(n13206), .C2(n13205), .A(n13204), .B(n13203), .ZN(
        n13207) );
  XNOR2_X1 U18674 ( .A(n13208), .B(n13207), .ZN(n13211) );
  XNOR2_X1 U18675 ( .A(n13209), .B(n3770), .ZN(n13210) );
  XNOR2_X1 U18676 ( .A(n13211), .B(n13210), .ZN(n13212) );
  XNOR2_X2 U18677 ( .A(n13213), .B(n13212), .ZN(n14030) );
  NAND2_X1 U18678 ( .A1(n14030), .A2(n29107), .ZN(n13214) );
  MUX2_X1 U18679 ( .A(n13215), .B(n13214), .S(n14029), .Z(n13216) );
  XNOR2_X1 U18680 ( .A(n13223), .B(n13224), .ZN(n13225) );
  NAND2_X1 U18681 ( .A1(n14045), .A2(n14043), .ZN(n13578) );
  INV_X1 U18682 ( .A(n13578), .ZN(n13256) );
  XNOR2_X1 U18683 ( .A(n13227), .B(n13226), .ZN(n13228) );
  XNOR2_X1 U18684 ( .A(n13229), .B(n13228), .ZN(n13235) );
  XNOR2_X1 U18685 ( .A(n13230), .B(n13231), .ZN(n13233) );
  XNOR2_X1 U18686 ( .A(n13450), .B(n2986), .ZN(n13232) );
  XNOR2_X1 U18687 ( .A(n13233), .B(n13232), .ZN(n13234) );
  XNOR2_X2 U18688 ( .A(n13235), .B(n13234), .ZN(n14051) );
  NAND2_X1 U18689 ( .A1(n14045), .A2(n14051), .ZN(n13909) );
  XNOR2_X1 U18690 ( .A(n13432), .B(n13236), .ZN(n13238) );
  XNOR2_X1 U18691 ( .A(n13238), .B(n13237), .ZN(n13242) );
  XNOR2_X1 U18692 ( .A(n13240), .B(n13239), .ZN(n13241) );
  XNOR2_X1 U18693 ( .A(n13244), .B(n13245), .ZN(n13430) );
  NOR2_X1 U18694 ( .A1(n14046), .A2(n14044), .ZN(n13255) );
  XNOR2_X1 U18695 ( .A(n13248), .B(n13247), .ZN(n13253) );
  XNOR2_X1 U18696 ( .A(n13249), .B(n13331), .ZN(n13251) );
  XNOR2_X1 U18697 ( .A(n13420), .B(n2523), .ZN(n13250) );
  XNOR2_X1 U18698 ( .A(n13251), .B(n13250), .ZN(n13252) );
  NAND2_X1 U18699 ( .A1(n1896), .A2(n14043), .ZN(n13254) );
  AOI21_X1 U18700 ( .B1(n14309), .B2(n14317), .A(n14318), .ZN(n13259) );
  NOR2_X1 U18701 ( .A1(n14320), .A2(n13884), .ZN(n13258) );
  XNOR2_X1 U18702 ( .A(n28603), .B(n13260), .ZN(n13264) );
  XNOR2_X1 U18703 ( .A(n13263), .B(n13262), .ZN(n13390) );
  XNOR2_X1 U18704 ( .A(n13390), .B(n13264), .ZN(n13268) );
  XNOR2_X1 U18705 ( .A(n13265), .B(n27956), .ZN(n13266) );
  XNOR2_X1 U18706 ( .A(n13425), .B(n13266), .ZN(n13267) );
  XNOR2_X1 U18707 ( .A(n13270), .B(n1062), .ZN(n13271) );
  XNOR2_X1 U18708 ( .A(n13412), .B(n13271), .ZN(n13276) );
  XNOR2_X1 U18709 ( .A(n13272), .B(n13273), .ZN(n13481) );
  XNOR2_X1 U18710 ( .A(n13481), .B(n13274), .ZN(n13275) );
  XNOR2_X1 U18711 ( .A(n13441), .B(n13277), .ZN(n13282) );
  XNOR2_X1 U18712 ( .A(n13278), .B(n2411), .ZN(n13279) );
  XNOR2_X1 U18713 ( .A(n13280), .B(n13279), .ZN(n13281) );
  XNOR2_X1 U18714 ( .A(n13283), .B(n13284), .ZN(n13289) );
  XNOR2_X1 U18715 ( .A(n13285), .B(n1927), .ZN(n13286) );
  XNOR2_X1 U18716 ( .A(n13287), .B(n13286), .ZN(n13288) );
  XNOR2_X1 U18718 ( .A(n13438), .B(n13290), .ZN(n13295) );
  XNOR2_X1 U18719 ( .A(n13291), .B(n3244), .ZN(n13292) );
  XNOR2_X1 U18720 ( .A(n13293), .B(n13292), .ZN(n13294) );
  XNOR2_X1 U18721 ( .A(n13294), .B(n13295), .ZN(n13646) );
  INV_X1 U18722 ( .A(n14053), .ZN(n14303) );
  NAND3_X1 U18723 ( .A1(n29611), .A2(n13646), .A3(n14303), .ZN(n13304) );
  INV_X1 U18724 ( .A(n14301), .ZN(n14054) );
  XNOR2_X1 U18725 ( .A(n13402), .B(n13296), .ZN(n13302) );
  XNOR2_X1 U18726 ( .A(n13297), .B(n13298), .ZN(n13300) );
  XNOR2_X1 U18727 ( .A(n13543), .B(n1193), .ZN(n13299) );
  XNOR2_X1 U18728 ( .A(n13300), .B(n13299), .ZN(n13301) );
  XNOR2_X1 U18729 ( .A(n13302), .B(n13301), .ZN(n14302) );
  NAND3_X1 U18730 ( .A1(n14054), .A2(n14302), .A3(n14304), .ZN(n13303) );
  NAND3_X1 U18731 ( .A1(n14563), .A2(n15690), .A3(n15691), .ZN(n13305) );
  INV_X1 U18732 ( .A(n15690), .ZN(n15087) );
  INV_X1 U18733 ( .A(n14563), .ZN(n15088) );
  NOR2_X1 U18734 ( .A1(n13803), .A2(n13699), .ZN(n13310) );
  OAI21_X1 U18736 ( .B1(n14293), .B2(n13306), .A(n14294), .ZN(n13307) );
  NAND2_X1 U18737 ( .A1(n14298), .A2(n13307), .ZN(n13308) );
  INV_X1 U18738 ( .A(n15083), .ZN(n15689) );
  NAND2_X1 U18739 ( .A1(n15088), .A2(n15689), .ZN(n13311) );
  AOI21_X1 U18740 ( .B1(n14878), .B2(n13311), .A(n15692), .ZN(n13312) );
  INV_X1 U18741 ( .A(n13314), .ZN(n13317) );
  INV_X1 U18742 ( .A(n13315), .ZN(n13316) );
  XNOR2_X1 U18743 ( .A(n13317), .B(n13316), .ZN(n13321) );
  XNOR2_X1 U18744 ( .A(n13525), .B(n4029), .ZN(n13319) );
  XNOR2_X1 U18745 ( .A(n13319), .B(n13318), .ZN(n13320) );
  XNOR2_X1 U18746 ( .A(n13538), .B(n3003), .ZN(n13323) );
  XNOR2_X1 U18747 ( .A(n13322), .B(n13323), .ZN(n13327) );
  XNOR2_X1 U18748 ( .A(n13325), .B(n13324), .ZN(n13326) );
  INV_X1 U18750 ( .A(n13328), .ZN(n13330) );
  XNOR2_X1 U18751 ( .A(n13329), .B(n13330), .ZN(n13335) );
  XNOR2_X1 U18752 ( .A(n13331), .B(n3062), .ZN(n13333) );
  XNOR2_X1 U18753 ( .A(n13332), .B(n13333), .ZN(n13334) );
  XNOR2_X1 U18754 ( .A(n13335), .B(n13334), .ZN(n13913) );
  INV_X1 U18755 ( .A(n13913), .ZN(n13729) );
  NOR2_X1 U18756 ( .A1(n6351), .A2(n13729), .ZN(n13336) );
  XNOR2_X1 U18757 ( .A(n13338), .B(n13337), .ZN(n13339) );
  XNOR2_X1 U18758 ( .A(n13340), .B(n13339), .ZN(n13345) );
  XNOR2_X1 U18759 ( .A(n13341), .B(n2995), .ZN(n13343) );
  XNOR2_X1 U18760 ( .A(n13343), .B(n13342), .ZN(n13344) );
  XNOR2_X1 U18762 ( .A(n13346), .B(n13347), .ZN(n13352) );
  XNOR2_X1 U18763 ( .A(n13348), .B(n2961), .ZN(n13349) );
  XNOR2_X1 U18764 ( .A(n13350), .B(n13349), .ZN(n13351) );
  XNOR2_X1 U18765 ( .A(n13352), .B(n13351), .ZN(n13583) );
  MUX2_X1 U18766 ( .A(n13912), .B(n13583), .S(n13729), .Z(n13358) );
  XNOR2_X1 U18767 ( .A(n13354), .B(n13353), .ZN(n13357) );
  XNOR2_X1 U18768 ( .A(n13562), .B(n2476), .ZN(n13355) );
  XNOR2_X1 U18769 ( .A(n13360), .B(n13359), .ZN(n13361) );
  XNOR2_X1 U18770 ( .A(n13362), .B(n13361), .ZN(n13368) );
  INV_X1 U18771 ( .A(n13363), .ZN(n13366) );
  XNOR2_X1 U18772 ( .A(n13364), .B(n891), .ZN(n13365) );
  XNOR2_X1 U18773 ( .A(n13366), .B(n13365), .ZN(n13367) );
  XNOR2_X1 U18774 ( .A(n13369), .B(n13370), .ZN(n13373) );
  XNOR2_X1 U18775 ( .A(n13371), .B(n26825), .ZN(n13372) );
  XNOR2_X1 U18776 ( .A(n13373), .B(n13372), .ZN(n13377) );
  XNOR2_X1 U18777 ( .A(n13374), .B(n13375), .ZN(n13376) );
  NAND2_X1 U18778 ( .A1(n13716), .A2(n14016), .ZN(n14142) );
  XNOR2_X1 U18779 ( .A(n13378), .B(n13379), .ZN(n13385) );
  XNOR2_X1 U18780 ( .A(n13381), .B(n1172), .ZN(n13382) );
  XNOR2_X1 U18781 ( .A(n13383), .B(n13382), .ZN(n13384) );
  XNOR2_X2 U18782 ( .A(n13385), .B(n13384), .ZN(n14144) );
  INV_X1 U18783 ( .A(n14144), .ZN(n13900) );
  XNOR2_X1 U18784 ( .A(n13386), .B(n2477), .ZN(n13387) );
  XNOR2_X1 U18785 ( .A(n13388), .B(n13387), .ZN(n13392) );
  XNOR2_X1 U18786 ( .A(n13390), .B(n13389), .ZN(n13391) );
  XNOR2_X1 U18787 ( .A(n13391), .B(n13392), .ZN(n13902) );
  INV_X1 U18788 ( .A(n13393), .ZN(n13395) );
  XNOR2_X1 U18789 ( .A(n13395), .B(n13394), .ZN(n13399) );
  XNOR2_X1 U18790 ( .A(n13396), .B(n2403), .ZN(n13397) );
  XNOR2_X1 U18791 ( .A(n13461), .B(n27894), .ZN(n13400) );
  XNOR2_X1 U18792 ( .A(n13400), .B(n29495), .ZN(n13403) );
  XNOR2_X1 U18793 ( .A(n13403), .B(n13402), .ZN(n13409) );
  XNOR2_X1 U18794 ( .A(n13405), .B(n13404), .ZN(n13407) );
  XNOR2_X1 U18795 ( .A(n13406), .B(n13407), .ZN(n13408) );
  INV_X1 U18796 ( .A(n13412), .ZN(n13417) );
  XNOR2_X1 U18797 ( .A(n13413), .B(n2509), .ZN(n13415) );
  XNOR2_X1 U18798 ( .A(n13415), .B(n13414), .ZN(n13416) );
  XNOR2_X1 U18799 ( .A(n13417), .B(n13416), .ZN(n13424) );
  INV_X1 U18800 ( .A(n13418), .ZN(n13422) );
  XNOR2_X1 U18801 ( .A(n13419), .B(n13420), .ZN(n13421) );
  XNOR2_X1 U18802 ( .A(n13422), .B(n13421), .ZN(n13423) );
  INV_X1 U18803 ( .A(n13425), .ZN(n13427) );
  XNOR2_X1 U18804 ( .A(n13428), .B(n3607), .ZN(n13429) );
  XNOR2_X1 U18805 ( .A(n13430), .B(n13429), .ZN(n13431) );
  XNOR2_X1 U18806 ( .A(n13432), .B(n13433), .ZN(n13435) );
  XNOR2_X1 U18807 ( .A(n13434), .B(n13435), .ZN(n13439) );
  INV_X1 U18808 ( .A(n3386), .ZN(n19658) );
  XNOR2_X1 U18809 ( .A(n13436), .B(n19658), .ZN(n13437) );
  NOR2_X1 U18810 ( .A1(n13440), .A2(n13726), .ZN(n13464) );
  INV_X1 U18811 ( .A(n13441), .ZN(n13443) );
  XNOR2_X1 U18812 ( .A(n13444), .B(n3650), .ZN(n13446) );
  XNOR2_X1 U18813 ( .A(n13448), .B(n13447), .ZN(n13449) );
  XNOR2_X1 U18814 ( .A(n28587), .B(n13450), .ZN(n13453) );
  INV_X1 U18815 ( .A(n1187), .ZN(n27534) );
  XNOR2_X1 U18816 ( .A(n13451), .B(n27534), .ZN(n13452) );
  XNOR2_X1 U18817 ( .A(n13453), .B(n13452), .ZN(n13454) );
  XNOR2_X1 U18818 ( .A(n13455), .B(n13454), .ZN(n13595) );
  XNOR2_X1 U18819 ( .A(n13461), .B(n2577), .ZN(n13462) );
  NAND2_X1 U18821 ( .A1(n14881), .A2(n388), .ZN(n13519) );
  NAND2_X1 U18822 ( .A1(n14030), .A2(n14031), .ZN(n13465) );
  OAI21_X1 U18823 ( .B1(n14029), .B2(n14030), .A(n13465), .ZN(n13467) );
  INV_X1 U18824 ( .A(n14030), .ZN(n13796) );
  INV_X1 U18825 ( .A(n14031), .ZN(n13916) );
  INV_X1 U18826 ( .A(n13793), .ZN(n14032) );
  NAND2_X1 U18827 ( .A1(n14031), .A2(n14032), .ZN(n13466) );
  INV_X1 U18828 ( .A(n14046), .ZN(n13662) );
  NAND3_X1 U18829 ( .A1(n13662), .A2(n14051), .A3(n13661), .ZN(n13468) );
  NAND3_X1 U18830 ( .A1(n14043), .A2(n14044), .A3(n14051), .ZN(n13469) );
  INV_X1 U18831 ( .A(n14045), .ZN(n13907) );
  XNOR2_X1 U18832 ( .A(n13472), .B(n13471), .ZN(n13477) );
  XNOR2_X1 U18833 ( .A(n13473), .B(n3722), .ZN(n13475) );
  XNOR2_X1 U18834 ( .A(n13474), .B(n13475), .ZN(n13476) );
  XNOR2_X1 U18836 ( .A(n29640), .B(n13478), .ZN(n13480) );
  XNOR2_X1 U18837 ( .A(n13479), .B(n13480), .ZN(n13483) );
  INV_X1 U18838 ( .A(n3067), .ZN(n27515) );
  XNOR2_X1 U18839 ( .A(n13485), .B(n13484), .ZN(n13486) );
  XNOR2_X1 U18840 ( .A(n13487), .B(n13486), .ZN(n13492) );
  XNOR2_X1 U18841 ( .A(n13488), .B(n1247), .ZN(n13489) );
  XNOR2_X1 U18842 ( .A(n13490), .B(n13489), .ZN(n13491) );
  XNOR2_X1 U18843 ( .A(n13493), .B(n3256), .ZN(n13495) );
  XNOR2_X1 U18844 ( .A(n13495), .B(n13494), .ZN(n13499) );
  XNOR2_X1 U18845 ( .A(n13496), .B(n13497), .ZN(n13498) );
  NAND2_X1 U18846 ( .A1(n13589), .A2(n13719), .ZN(n14000) );
  INV_X1 U18847 ( .A(n13501), .ZN(n13502) );
  XNOR2_X1 U18848 ( .A(n13502), .B(n13503), .ZN(n13508) );
  XNOR2_X1 U18849 ( .A(n13504), .B(n28693), .ZN(n13506) );
  XNOR2_X1 U18850 ( .A(n13505), .B(n13506), .ZN(n13507) );
  XNOR2_X1 U18851 ( .A(n13509), .B(n13510), .ZN(n13515) );
  XNOR2_X1 U18852 ( .A(n13511), .B(n26032), .ZN(n13512) );
  XNOR2_X1 U18853 ( .A(n13513), .B(n13512), .ZN(n13514) );
  INV_X1 U18855 ( .A(n14974), .ZN(n13517) );
  NAND2_X1 U18856 ( .A1(n13517), .A2(n14972), .ZN(n13518) );
  XNOR2_X1 U18857 ( .A(n16346), .B(n16312), .ZN(n13603) );
  XNOR2_X1 U18858 ( .A(n13522), .B(n13521), .ZN(n13529) );
  XNOR2_X1 U18859 ( .A(n13524), .B(n13523), .ZN(n13527) );
  XNOR2_X1 U18860 ( .A(n13525), .B(n3673), .ZN(n13526) );
  XNOR2_X1 U18861 ( .A(n13527), .B(n13526), .ZN(n13528) );
  INV_X1 U18862 ( .A(n14007), .ZN(n14386) );
  INV_X1 U18863 ( .A(n13530), .ZN(n13531) );
  XNOR2_X1 U18864 ( .A(n13531), .B(n13532), .ZN(n13537) );
  XNOR2_X1 U18865 ( .A(n13533), .B(n1079), .ZN(n13534) );
  XNOR2_X1 U18866 ( .A(n13535), .B(n13534), .ZN(n13536) );
  XNOR2_X1 U18867 ( .A(n13537), .B(n13536), .ZN(n13837) );
  XNOR2_X1 U18868 ( .A(n13538), .B(n13539), .ZN(n13541) );
  XNOR2_X1 U18869 ( .A(n13540), .B(n13541), .ZN(n13544) );
  XNOR2_X1 U18870 ( .A(n13546), .B(n13545), .ZN(n13551) );
  XNOR2_X1 U18871 ( .A(n13547), .B(n3635), .ZN(n13548) );
  XNOR2_X1 U18872 ( .A(n13549), .B(n13548), .ZN(n13550) );
  XNOR2_X1 U18873 ( .A(n13551), .B(n13550), .ZN(n14381) );
  AOI22_X1 U18874 ( .A1(n14386), .A2(n14150), .B1(n13572), .B2(n14381), .ZN(
        n13575) );
  XNOR2_X1 U18875 ( .A(n13552), .B(n13553), .ZN(n13555) );
  XNOR2_X1 U18876 ( .A(n13554), .B(n13555), .ZN(n13561) );
  XNOR2_X1 U18877 ( .A(n13104), .B(n1919), .ZN(n13559) );
  XNOR2_X1 U18878 ( .A(n13557), .B(n13556), .ZN(n13558) );
  XNOR2_X1 U18879 ( .A(n13559), .B(n13558), .ZN(n13560) );
  XNOR2_X1 U18880 ( .A(n13563), .B(n13562), .ZN(n13564) );
  XNOR2_X1 U18881 ( .A(n13565), .B(n13564), .ZN(n13571) );
  XNOR2_X1 U18882 ( .A(n13567), .B(n3081), .ZN(n13568) );
  XNOR2_X1 U18883 ( .A(n13569), .B(n13568), .ZN(n13570) );
  NOR2_X1 U18884 ( .A1(n14007), .A2(n14381), .ZN(n13734) );
  NOR2_X1 U18885 ( .A1(n13573), .A2(n13734), .ZN(n13574) );
  NAND2_X1 U18886 ( .A1(n14043), .A2(n13661), .ZN(n13576) );
  INV_X1 U18887 ( .A(n14043), .ZN(n13906) );
  NAND2_X1 U18888 ( .A1(n14047), .A2(n13906), .ZN(n13577) );
  NAND3_X1 U18889 ( .A1(n13578), .A2(n5731), .A3(n13577), .ZN(n13579) );
  NOR2_X1 U18890 ( .A1(n13716), .A2(n29589), .ZN(n13581) );
  NAND2_X1 U18891 ( .A1(n13912), .A2(n13583), .ZN(n13582) );
  NAND2_X1 U18892 ( .A1(n6351), .A2(n13914), .ZN(n13585) );
  INV_X1 U18893 ( .A(n13583), .ZN(n13910) );
  OAI211_X1 U18894 ( .C1(n13730), .C2(n13914), .A(n5847), .B(n13910), .ZN(
        n13584) );
  MUX2_X1 U18895 ( .A(n13589), .B(n13587), .S(n13719), .Z(n13588) );
  NOR2_X1 U18896 ( .A1(n13588), .A2(n14039), .ZN(n13590) );
  NAND2_X1 U18897 ( .A1(n13719), .A2(n28569), .ZN(n13999) );
  NAND2_X1 U18898 ( .A1(n13592), .A2(n28196), .ZN(n13600) );
  NOR2_X1 U18899 ( .A1(n13593), .A2(n13726), .ZN(n13597) );
  NOR2_X1 U18900 ( .A1(n28518), .A2(n13638), .ZN(n14895) );
  INV_X1 U18901 ( .A(n14895), .ZN(n13598) );
  NAND2_X1 U18902 ( .A1(n13598), .A2(n15400), .ZN(n13599) );
  NAND2_X1 U18903 ( .A1(n13600), .A2(n13599), .ZN(n13601) );
  XNOR2_X1 U18904 ( .A(n13603), .B(n15777), .ZN(n13604) );
  NOR2_X1 U18905 ( .A1(n14231), .A2(n14107), .ZN(n13607) );
  MUX2_X1 U18906 ( .A(n6956), .B(n13607), .S(n14593), .Z(n13610) );
  AOI21_X1 U18907 ( .B1(n14235), .B2(n13608), .A(n14230), .ZN(n13609) );
  NOR2_X2 U18908 ( .A1(n13610), .A2(n13609), .ZN(n15004) );
  NAND2_X1 U18909 ( .A1(n1743), .A2(n14262), .ZN(n13763) );
  INV_X1 U18910 ( .A(n13763), .ZN(n13612) );
  NAND2_X1 U18912 ( .A1(n14362), .A2(n28507), .ZN(n13617) );
  INV_X1 U18913 ( .A(n13832), .ZN(n14271) );
  NAND3_X1 U18914 ( .A1(n14272), .A2(n14271), .A3(n14278), .ZN(n13616) );
  NAND2_X1 U18916 ( .A1(n15001), .A2(n15127), .ZN(n14688) );
  INV_X1 U18917 ( .A(n13770), .ZN(n13620) );
  INV_X1 U18920 ( .A(n14091), .ZN(n14369) );
  NAND2_X1 U18921 ( .A1(n14091), .A2(n14365), .ZN(n14118) );
  NOR2_X1 U18922 ( .A1(n14118), .A2(n14366), .ZN(n13624) );
  AOI21_X2 U18923 ( .B1(n13625), .B2(n1960), .A(n13624), .ZN(n15000) );
  NAND2_X1 U18924 ( .A1(n14351), .A2(n4893), .ZN(n13626) );
  NAND3_X1 U18925 ( .A1(n13627), .A2(n13626), .A3(n13826), .ZN(n13631) );
  INV_X1 U18926 ( .A(n14354), .ZN(n14353) );
  NAND3_X1 U18927 ( .A1(n13825), .A2(n4893), .A3(n14353), .ZN(n13629) );
  NAND2_X1 U18928 ( .A1(n14126), .A2(n14355), .ZN(n13628) );
  NAND2_X1 U18929 ( .A1(n13631), .A2(n13630), .ZN(n15123) );
  INV_X1 U18930 ( .A(n15004), .ZN(n15125) );
  NOR2_X1 U18931 ( .A1(n15127), .A2(n15123), .ZN(n13633) );
  AOI21_X1 U18932 ( .B1(n14686), .B2(n15125), .A(n13633), .ZN(n13634) );
  OAI21_X1 U18933 ( .B1(n14944), .B2(n13637), .A(n13636), .ZN(n14945) );
  INV_X1 U18934 ( .A(n13638), .ZN(n15401) );
  NAND2_X1 U18935 ( .A1(n14945), .A2(n15401), .ZN(n13642) );
  OAI21_X1 U18936 ( .B1(n14944), .B2(n14943), .A(n13639), .ZN(n13640) );
  NAND2_X1 U18937 ( .A1(n13640), .A2(n28196), .ZN(n13641) );
  NAND2_X1 U18938 ( .A1(n5887), .A2(n13583), .ZN(n13643) );
  AOI21_X2 U18939 ( .B1(n13645), .B2(n13730), .A(n13644), .ZN(n15115) );
  NAND2_X1 U18940 ( .A1(n14301), .A2(n14304), .ZN(n13651) );
  INV_X1 U18941 ( .A(n13647), .ZN(n13648) );
  NAND2_X1 U18942 ( .A1(n13648), .A2(n14054), .ZN(n13649) );
  INV_X1 U18943 ( .A(n13652), .ZN(n14324) );
  INV_X1 U18944 ( .A(n13653), .ZN(n14065) );
  INV_X1 U18945 ( .A(n14328), .ZN(n13654) );
  NOR2_X1 U18946 ( .A1(n14327), .A2(n13654), .ZN(n13656) );
  OAI211_X1 U18947 ( .C1(n29626), .C2(n14328), .A(n13653), .B(n14064), .ZN(
        n13655) );
  NAND2_X1 U18948 ( .A1(n13808), .A2(n13803), .ZN(n13659) );
  INV_X1 U18949 ( .A(n14295), .ZN(n13806) );
  NAND3_X1 U18950 ( .A1(n14295), .A2(n14291), .A3(n14297), .ZN(n13657) );
  OAI21_X1 U18951 ( .B1(n15115), .B2(n1001), .A(n13660), .ZN(n14114) );
  NOR2_X1 U18952 ( .A1(n14045), .A2(n13661), .ZN(n13664) );
  NOR2_X1 U18953 ( .A1(n1896), .A2(n14051), .ZN(n13663) );
  MUX2_X1 U18954 ( .A(n13664), .B(n13663), .S(n13662), .Z(n13665) );
  INV_X1 U18955 ( .A(n14514), .ZN(n15116) );
  INV_X1 U18956 ( .A(n14029), .ZN(n13921) );
  NAND2_X1 U18957 ( .A1(n13916), .A2(n29107), .ZN(n13666) );
  OR2_X1 U18958 ( .A1(n13666), .A2(n14032), .ZN(n13667) );
  XNOR2_X1 U18960 ( .A(n29319), .B(n28557), .ZN(n13669) );
  XNOR2_X1 U18961 ( .A(n13669), .B(n13670), .ZN(n13760) );
  INV_X1 U18962 ( .A(n14207), .ZN(n14439) );
  NOR2_X1 U18963 ( .A1(n14207), .A2(n1876), .ZN(n13671) );
  INV_X1 U18964 ( .A(n13672), .ZN(n13673) );
  OAI21_X1 U18965 ( .B1(n14492), .B2(n14497), .A(n13856), .ZN(n13676) );
  NAND2_X1 U18967 ( .A1(n14492), .A2(n29036), .ZN(n13675) );
  NAND2_X1 U18968 ( .A1(n15389), .A2(n15388), .ZN(n14723) );
  INV_X1 U18969 ( .A(n14464), .ZN(n13852) );
  INV_X1 U18970 ( .A(n13678), .ZN(n14467) );
  NAND3_X1 U18971 ( .A1(n14467), .A2(n13852), .A3(n4840), .ZN(n13681) );
  NAND3_X1 U18972 ( .A1(n14185), .A2(n13678), .A3(n14464), .ZN(n13679) );
  NOR2_X1 U18973 ( .A1(n12711), .A2(n14456), .ZN(n13682) );
  NAND2_X1 U18977 ( .A1(n14416), .A2(n14414), .ZN(n13893) );
  INV_X1 U18978 ( .A(n14193), .ZN(n13867) );
  NAND3_X1 U18979 ( .A1(n28805), .A2(n14192), .A3(n13867), .ZN(n13688) );
  INV_X1 U18982 ( .A(n14992), .ZN(n15391) );
  MUX2_X1 U18985 ( .A(n29133), .B(n14406), .S(n14407), .Z(n13693) );
  INV_X1 U18986 ( .A(n14333), .ZN(n13692) );
  OAI21_X1 U18987 ( .B1(n13653), .B2(n14061), .A(n14324), .ZN(n13694) );
  AOI21_X1 U18989 ( .B1(n14291), .B2(n14293), .A(n13697), .ZN(n13698) );
  NAND2_X1 U18990 ( .A1(n13698), .A2(n13702), .ZN(n13701) );
  NOR2_X1 U18991 ( .A1(n14292), .A2(n13699), .ZN(n13807) );
  NAND2_X1 U18992 ( .A1(n13807), .A2(n13803), .ZN(n13700) );
  OAI211_X1 U18993 ( .C1(n13702), .C2(n14294), .A(n13701), .B(n13700), .ZN(
        n15137) );
  NAND2_X1 U18994 ( .A1(n15248), .A2(n15137), .ZN(n15247) );
  NOR2_X1 U18995 ( .A1(n13872), .A2(n14429), .ZN(n13706) );
  INV_X1 U18996 ( .A(n14426), .ZN(n13873) );
  NAND2_X1 U18998 ( .A1(n15250), .A2(n15137), .ZN(n13710) );
  OAI21_X1 U19000 ( .B1(n14398), .B2(n28804), .A(n14402), .ZN(n13707) );
  MUX2_X1 U19001 ( .A(n13710), .B(n14733), .S(n15246), .Z(n13715) );
  NAND3_X1 U19002 ( .A1(n14312), .A2(n13711), .A3(n14313), .ZN(n13713) );
  NAND3_X1 U19003 ( .A1(n15249), .A2(n15135), .A3(n15250), .ZN(n13714) );
  XNOR2_X1 U19004 ( .A(n16160), .B(n16126), .ZN(n16418) );
  INV_X1 U19005 ( .A(n15372), .ZN(n15374) );
  NAND3_X1 U19006 ( .A1(n13726), .A2(n5404), .A3(n14146), .ZN(n13727) );
  INV_X1 U19008 ( .A(n14010), .ZN(n14344) );
  NAND2_X1 U19009 ( .A1(n14346), .A2(n14132), .ZN(n14134) );
  NOR2_X1 U19011 ( .A1(n14344), .A2(n14345), .ZN(n13728) );
  INV_X1 U19012 ( .A(n14380), .ZN(n14385) );
  MUX2_X1 U19013 ( .A(n14007), .B(n14385), .S(n14150), .Z(n13736) );
  INV_X1 U19014 ( .A(n13572), .ZN(n13836) );
  NOR2_X1 U19015 ( .A1(n13836), .A2(n14380), .ZN(n13733) );
  AOI22_X1 U19016 ( .A1(n13734), .A2(n14004), .B1(n13733), .B2(n14007), .ZN(
        n13735) );
  NAND2_X1 U19017 ( .A1(n28172), .A2(n14241), .ZN(n13769) );
  NOR2_X1 U19018 ( .A1(n15194), .A2(n14241), .ZN(n15192) );
  NAND2_X1 U19019 ( .A1(n15192), .A2(n29097), .ZN(n13741) );
  OAI211_X1 U19020 ( .C1(n29097), .C2(n14238), .A(n15194), .B(n13739), .ZN(
        n13740) );
  INV_X1 U19021 ( .A(n15379), .ZN(n15152) );
  NOR2_X1 U19022 ( .A1(n14166), .A2(n14484), .ZN(n13742) );
  INV_X1 U19023 ( .A(n14481), .ZN(n14164) );
  INV_X1 U19024 ( .A(n15382), .ZN(n13752) );
  OAI22_X1 U19025 ( .A1(n13744), .A2(n14252), .B1(n14078), .B2(n13778), .ZN(
        n14076) );
  INV_X1 U19026 ( .A(n14078), .ZN(n14251) );
  NOR2_X1 U19027 ( .A1(n14251), .A2(n14250), .ZN(n13746) );
  INV_X1 U19028 ( .A(n15383), .ZN(n15150) );
  NOR2_X1 U19029 ( .A1(n14268), .A2(n14262), .ZN(n13748) );
  MUX2_X1 U19030 ( .A(n13748), .B(n13747), .S(n14264), .Z(n13751) );
  NAND2_X1 U19031 ( .A1(n14261), .A2(n14259), .ZN(n14266) );
  OAI21_X1 U19032 ( .B1(n14264), .B2(n14266), .A(n14098), .ZN(n13750) );
  AOI21_X1 U19033 ( .B1(n13752), .B2(n15150), .A(n15151), .ZN(n13758) );
  OAI22_X1 U19034 ( .A1(n14177), .A2(n14452), .B1(n13753), .B2(n14178), .ZN(
        n13850) );
  OAI22_X1 U19035 ( .A1(n15155), .A2(n15379), .B1(n15151), .B2(n15383), .ZN(
        n15381) );
  NAND2_X1 U19036 ( .A1(n14475), .A2(n13936), .ZN(n13756) );
  NOR2_X1 U19037 ( .A1(n14480), .A2(n13936), .ZN(n13757) );
  INV_X1 U19038 ( .A(n14986), .ZN(n15384) );
  XNOR2_X1 U19039 ( .A(n16456), .B(n16318), .ZN(n16162) );
  XNOR2_X1 U19040 ( .A(n16162), .B(n16418), .ZN(n13759) );
  XNOR2_X1 U19041 ( .A(n13760), .B(n13759), .ZN(n17716) );
  INV_X1 U19042 ( .A(n17716), .ZN(n17720) );
  MUX2_X1 U19043 ( .A(n13762), .B(n13761), .S(n14099), .Z(n13764) );
  NAND3_X1 U19045 ( .A1(n29306), .A2(n14481), .A3(n14486), .ZN(n13765) );
  NAND2_X1 U19046 ( .A1(n15201), .A2(n15207), .ZN(n14968) );
  MUX2_X1 U19047 ( .A(n15195), .B(n13943), .S(n28172), .Z(n13768) );
  AND3_X1 U19048 ( .A1(n13767), .A2(n14174), .A3(n14241), .ZN(n15193) );
  MUX2_X1 U19049 ( .A(n14285), .B(n14083), .S(n14287), .Z(n13774) );
  NAND2_X1 U19050 ( .A1(n14082), .A2(n14084), .ZN(n13771) );
  AND2_X1 U19051 ( .A1(n13771), .A2(n13770), .ZN(n13773) );
  INV_X1 U19052 ( .A(n14286), .ZN(n14081) );
  NOR2_X1 U19053 ( .A1(n14287), .A2(n14081), .ZN(n13772) );
  INV_X1 U19054 ( .A(n14963), .ZN(n15209) );
  INV_X1 U19055 ( .A(n13775), .ZN(n14077) );
  MUX2_X1 U19056 ( .A(n14252), .B(n14077), .S(n14078), .Z(n13781) );
  INV_X1 U19057 ( .A(n13776), .ZN(n14253) );
  NAND3_X1 U19058 ( .A1(n13778), .A2(n14252), .A3(n14077), .ZN(n13779) );
  INV_X1 U19060 ( .A(n15208), .ZN(n13782) );
  INV_X1 U19061 ( .A(n15207), .ZN(n15204) );
  NAND3_X1 U19062 ( .A1(n15209), .A2(n13782), .A3(n15204), .ZN(n13787) );
  NAND2_X1 U19063 ( .A1(n14230), .A2(n14593), .ZN(n13784) );
  OAI211_X1 U19064 ( .C1(n14960), .C2(n15207), .A(n13785), .B(n15202), .ZN(
        n13786) );
  INV_X1 U19066 ( .A(n14881), .ZN(n14976) );
  NAND2_X1 U19067 ( .A1(n14882), .A2(n13789), .ZN(n14970) );
  OAI21_X1 U19068 ( .B1(n14976), .B2(n14970), .A(n13788), .ZN(n13792) );
  NOR2_X1 U19069 ( .A1(n13789), .A2(n14972), .ZN(n13790) );
  XNOR2_X1 U19070 ( .A(n15070), .B(n16284), .ZN(n16171) );
  NAND2_X1 U19071 ( .A1(n6066), .A2(n14032), .ZN(n13797) );
  AOI21_X1 U19072 ( .B1(n6066), .B2(n14031), .A(n13793), .ZN(n13795) );
  NOR2_X1 U19074 ( .A1(n14324), .A2(n14328), .ZN(n13798) );
  NAND2_X1 U19075 ( .A1(n14314), .A2(n14318), .ZN(n13886) );
  NAND2_X1 U19076 ( .A1(n13886), .A2(n14313), .ZN(n13801) );
  AOI21_X1 U19077 ( .B1(n14313), .B2(n560), .A(n14314), .ZN(n13800) );
  MUX2_X1 U19078 ( .A(n13805), .B(n13804), .S(n14294), .Z(n13810) );
  AOI22_X1 U19079 ( .A1(n13808), .A2(n14291), .B1(n13807), .B2(n13806), .ZN(
        n13809) );
  NAND2_X1 U19080 ( .A1(n14332), .A2(n14405), .ZN(n13812) );
  OAI21_X1 U19081 ( .B1(n14408), .B2(n13878), .A(n13879), .ZN(n13811) );
  OAI21_X1 U19082 ( .B1(n13813), .B2(n13812), .A(n13811), .ZN(n13814) );
  NOR2_X1 U19083 ( .A1(n15184), .A2(n14784), .ZN(n15187) );
  NAND2_X1 U19084 ( .A1(n28625), .A2(n14084), .ZN(n14284) );
  OAI21_X1 U19085 ( .B1(n14085), .B2(n14285), .A(n561), .ZN(n13821) );
  NAND2_X1 U19086 ( .A1(n13821), .A2(n14082), .ZN(n13823) );
  NAND3_X1 U19087 ( .A1(n14286), .A2(n561), .A3(n14282), .ZN(n13822) );
  NAND2_X1 U19088 ( .A1(n14362), .A2(n13832), .ZN(n14363) );
  INV_X1 U19089 ( .A(n14363), .ZN(n13828) );
  NAND2_X1 U19090 ( .A1(n13828), .A2(n13827), .ZN(n13831) );
  INV_X1 U19091 ( .A(n14360), .ZN(n14273) );
  NAND3_X1 U19092 ( .A1(n14359), .A2(n14273), .A3(n28507), .ZN(n13830) );
  NOR2_X1 U19093 ( .A1(n308), .A2(n14091), .ZN(n13834) );
  NAND2_X1 U19095 ( .A1(n13836), .A2(n14380), .ZN(n13840) );
  NAND3_X1 U19096 ( .A1(n14006), .A2(n557), .A3(n14150), .ZN(n13839) );
  OAI21_X1 U19097 ( .B1(n13572), .B2(n14004), .A(n556), .ZN(n13838) );
  OAI21_X1 U19098 ( .B1(n14797), .B2(n15460), .A(n13841), .ZN(n13846) );
  OAI21_X1 U19099 ( .B1(n14135), .B2(n14346), .A(n14343), .ZN(n13843) );
  MUX2_X1 U19100 ( .A(n28803), .B(n15180), .S(n15175), .Z(n13844) );
  XNOR2_X1 U19101 ( .A(n15738), .B(n16366), .ZN(n16044) );
  XNOR2_X1 U19102 ( .A(n16171), .B(n16044), .ZN(n13927) );
  AOI21_X1 U19103 ( .B1(n14435), .B2(n14439), .A(n14433), .ZN(n13849) );
  OAI22_X1 U19104 ( .A1(n14438), .A2(n14434), .B1(n14207), .B2(n14433), .ZN(
        n14206) );
  NAND2_X1 U19105 ( .A1(n14206), .A2(n14432), .ZN(n13848) );
  NOR2_X1 U19106 ( .A1(n15476), .A2(n15168), .ZN(n13861) );
  NAND2_X1 U19107 ( .A1(n13851), .A2(n14452), .ZN(n14453) );
  NAND3_X1 U19108 ( .A1(n14453), .A2(n13753), .A3(n14451), .ZN(n14548) );
  OAI21_X1 U19109 ( .B1(n14466), .B2(n4840), .A(n14182), .ZN(n14183) );
  NAND2_X1 U19110 ( .A1(n13933), .A2(n14464), .ZN(n13854) );
  NAND2_X1 U19111 ( .A1(n14492), .A2(n14497), .ZN(n14155) );
  NAND2_X1 U19112 ( .A1(n14493), .A2(n13674), .ZN(n13858) );
  NAND3_X1 U19114 ( .A1(n14498), .A2(n14491), .A3(n14494), .ZN(n13859) );
  OAI211_X1 U19115 ( .C1(n29037), .C2(n14155), .A(n13860), .B(n13859), .ZN(
        n15167) );
  INV_X1 U19116 ( .A(n15168), .ZN(n14551) );
  NAND2_X1 U19117 ( .A1(n13967), .A2(n14459), .ZN(n13862) );
  INV_X1 U19119 ( .A(n15166), .ZN(n15471) );
  NAND3_X1 U19120 ( .A1(n14193), .A2(n14393), .A3(n14194), .ZN(n13869) );
  OAI211_X1 U19121 ( .C1(n13873), .C2(n13872), .A(n13871), .B(n28199), .ZN(
        n13876) );
  NOR2_X1 U19122 ( .A1(n15466), .A2(n4515), .ZN(n13890) );
  MUX2_X1 U19123 ( .A(n13879), .B(n13878), .S(n14405), .Z(n13880) );
  NAND3_X1 U19124 ( .A1(n14332), .A2(n1830), .A3(n29133), .ZN(n13881) );
  OAI21_X1 U19125 ( .B1(n13884), .B2(n14312), .A(n14318), .ZN(n13885) );
  OR2_X1 U19126 ( .A1(n560), .A2(n13886), .ZN(n13887) );
  NAND3_X1 U19129 ( .A1(n13891), .A2(n14216), .A3(n28647), .ZN(n13892) );
  XNOR2_X1 U19130 ( .A(n16192), .B(n16634), .ZN(n16397) );
  INV_X1 U19132 ( .A(n14773), .ZN(n14808) );
  NAND2_X1 U19133 ( .A1(n14020), .A2(n13901), .ZN(n13905) );
  NOR2_X1 U19134 ( .A1(n14808), .A2(n14807), .ZN(n14712) );
  OAI211_X1 U19135 ( .C1(n14030), .C2(n14033), .A(n13917), .B(n13916), .ZN(
        n13919) );
  NAND3_X1 U19136 ( .A1(n6066), .A2(n14032), .A3(n29107), .ZN(n13918) );
  OAI211_X1 U19137 ( .C1(n13921), .C2(n29107), .A(n13919), .B(n13918), .ZN(
        n14806) );
  INV_X1 U19138 ( .A(n14806), .ZN(n14767) );
  NAND2_X1 U19139 ( .A1(n14807), .A2(n28493), .ZN(n13923) );
  INV_X1 U19140 ( .A(n14302), .ZN(n14059) );
  AOI21_X1 U19141 ( .B1(n14059), .B2(n5956), .A(n29611), .ZN(n14771) );
  MUX2_X1 U19142 ( .A(n14300), .B(n14299), .S(n28478), .Z(n14770) );
  NAND2_X1 U19143 ( .A1(n14302), .A2(n14303), .ZN(n14769) );
  NAND3_X1 U19144 ( .A1(n14810), .A2(n14807), .A3(n14713), .ZN(n13925) );
  NAND2_X1 U19145 ( .A1(n14176), .A2(n14452), .ZN(n13928) );
  NAND2_X1 U19146 ( .A1(n1320), .A2(n13928), .ZN(n13929) );
  OAI21_X1 U19147 ( .B1(n13930), .B2(n1320), .A(n13929), .ZN(n13931) );
  NAND2_X1 U19149 ( .A1(n14249), .A2(n14250), .ZN(n14237) );
  NAND2_X1 U19150 ( .A1(n14251), .A2(n14077), .ZN(n13938) );
  NAND2_X1 U19151 ( .A1(n15438), .A2(n15300), .ZN(n13941) );
  INV_X1 U19152 ( .A(n15438), .ZN(n15302) );
  INV_X1 U19153 ( .A(n15018), .ZN(n15437) );
  NOR2_X1 U19154 ( .A1(n15444), .A2(n15437), .ZN(n14667) );
  NAND2_X1 U19155 ( .A1(n15303), .A2(n15302), .ZN(n13949) );
  NOR2_X1 U19156 ( .A1(n14193), .A2(n14192), .ZN(n13952) );
  NAND2_X1 U19158 ( .A1(n13956), .A2(n13955), .ZN(n15015) );
  INV_X1 U19159 ( .A(n13957), .ZN(n13958) );
  AOI21_X1 U19160 ( .B1(n14438), .B2(n14432), .A(n14437), .ZN(n13960) );
  OAI21_X1 U19161 ( .B1(n13963), .B2(n13962), .A(n30), .ZN(n13964) );
  OAI21_X2 U19162 ( .B1(n13965), .B2(n14400), .A(n13964), .ZN(n15014) );
  INV_X1 U19163 ( .A(n14459), .ZN(n13966) );
  NAND3_X1 U19164 ( .A1(n14204), .A2(n14456), .A3(n13966), .ZN(n13971) );
  AND2_X1 U19165 ( .A1(n14455), .A2(n13967), .ZN(n13968) );
  NAND2_X1 U19166 ( .A1(n13968), .A2(n14200), .ZN(n13970) );
  NAND4_X1 U19167 ( .A1(n14463), .A2(n13971), .A3(n13970), .A4(n13969), .ZN(
        n15013) );
  AOI21_X1 U19168 ( .B1(n14155), .B2(n14494), .A(n14491), .ZN(n13975) );
  NAND2_X1 U19169 ( .A1(n14493), .A2(n14491), .ZN(n13972) );
  AOI21_X1 U19170 ( .B1(n13973), .B2(n13972), .A(n14497), .ZN(n13974) );
  NAND2_X1 U19171 ( .A1(n15447), .A2(n15321), .ZN(n13976) );
  XNOR2_X1 U19172 ( .A(n16564), .B(n16146), .ZN(n16424) );
  NOR2_X1 U19173 ( .A1(n15115), .A2(n15117), .ZN(n14112) );
  INV_X1 U19174 ( .A(n14112), .ZN(n13982) );
  INV_X1 U19175 ( .A(n14743), .ZN(n15114) );
  OAI21_X1 U19176 ( .B1(n15113), .B2(n1904), .A(n14744), .ZN(n13981) );
  NOR2_X1 U19177 ( .A1(n14514), .A2(n14740), .ZN(n13980) );
  AOI21_X1 U19178 ( .B1(n13982), .B2(n13981), .A(n13980), .ZN(n13984) );
  NOR2_X1 U19179 ( .A1(n15115), .A2(n15113), .ZN(n15120) );
  AND2_X1 U19180 ( .A1(n15120), .A2(n15116), .ZN(n13983) );
  NOR2_X1 U19181 ( .A1(n15125), .A2(n15000), .ZN(n13987) );
  AOI22_X1 U19182 ( .A1(n15132), .A2(n13987), .B1(n15004), .B2(n13986), .ZN(
        n13988) );
  XNOR2_X1 U19183 ( .A(n28579), .B(n15788), .ZN(n16183) );
  XNOR2_X1 U19184 ( .A(n16183), .B(n16424), .ZN(n14028) );
  INV_X1 U19185 ( .A(n15085), .ZN(n13989) );
  NAND2_X1 U19186 ( .A1(n13989), .A2(n15691), .ZN(n13992) );
  NAND2_X1 U19187 ( .A1(n15691), .A2(n323), .ZN(n14566) );
  OAI21_X1 U19188 ( .B1(n1886), .B2(n14563), .A(n15690), .ZN(n13991) );
  OAI21_X1 U19190 ( .B1(n15098), .B2(n15094), .A(n15099), .ZN(n13996) );
  OAI21_X1 U19191 ( .B1(n13993), .B2(n14902), .A(n14679), .ZN(n13995) );
  AND2_X1 U19192 ( .A1(n13993), .A2(n15094), .ZN(n13994) );
  XNOR2_X1 U19193 ( .A(n16062), .B(n16295), .ZN(n14026) );
  MUX2_X1 U19194 ( .A(n13999), .B(n13998), .S(n14036), .Z(n14003) );
  INV_X1 U19195 ( .A(n14000), .ZN(n14001) );
  AOI22_X1 U19196 ( .A1(n14001), .A2(n14036), .B1(n13587), .B2(n28569), .ZN(
        n14002) );
  NAND2_X1 U19197 ( .A1(n14003), .A2(n14002), .ZN(n14824) );
  INV_X1 U19198 ( .A(n14004), .ZN(n14382) );
  AND2_X1 U19199 ( .A1(n14824), .A2(n15431), .ZN(n14823) );
  INV_X1 U19200 ( .A(n14823), .ZN(n14024) );
  NAND3_X1 U19202 ( .A1(n14341), .A2(n14344), .A3(n14345), .ZN(n14012) );
  NAND3_X1 U19203 ( .A1(n14132), .A2(n14135), .A3(n14136), .ZN(n14011) );
  INV_X1 U19204 ( .A(n14821), .ZN(n15432) );
  NAND2_X1 U19205 ( .A1(n2974), .A2(n14144), .ZN(n14019) );
  NOR2_X1 U19206 ( .A1(n29589), .A2(n4425), .ZN(n14017) );
  AOI22_X1 U19207 ( .A1(n14020), .A2(n14019), .B1(n14018), .B2(n14017), .ZN(
        n14825) );
  INV_X1 U19208 ( .A(n14825), .ZN(n15027) );
  NAND3_X1 U19209 ( .A1(n15031), .A2(n14821), .A3(n15027), .ZN(n14021) );
  XNOR2_X1 U19210 ( .A(n16059), .B(n3380), .ZN(n14025) );
  XNOR2_X1 U19211 ( .A(n14026), .B(n14025), .ZN(n14027) );
  INV_X1 U19213 ( .A(n17428), .ZN(n17005) );
  MUX2_X1 U19215 ( .A(n14030), .B(n14031), .S(n14029), .Z(n14035) );
  MUX2_X1 U19216 ( .A(n14032), .B(n6066), .S(n14031), .Z(n14034) );
  NAND2_X1 U19218 ( .A1(n14046), .A2(n14051), .ZN(n14048) );
  MUX2_X1 U19219 ( .A(n14049), .B(n14048), .S(n14047), .Z(n14050) );
  NOR2_X1 U19220 ( .A1(n14300), .A2(n28478), .ZN(n14055) );
  INV_X1 U19221 ( .A(n14055), .ZN(n14058) );
  OAI21_X1 U19222 ( .B1(n14055), .B2(n5956), .A(n14054), .ZN(n14057) );
  NAND3_X1 U19223 ( .A1(n29611), .A2(n14300), .A3(n14299), .ZN(n14056) );
  OAI211_X2 U19224 ( .C1(n14058), .C2(n14059), .A(n14057), .B(n14056), .ZN(
        n14842) );
  NOR2_X1 U19225 ( .A1(n28842), .A2(n14060), .ZN(n14074) );
  INV_X1 U19226 ( .A(n14061), .ZN(n14063) );
  MUX2_X1 U19227 ( .A(n14323), .B(n14063), .S(n29626), .Z(n14067) );
  NAND2_X1 U19228 ( .A1(n15286), .A2(n14601), .ZN(n14073) );
  NAND2_X1 U19229 ( .A1(n14068), .A2(n13583), .ZN(n14069) );
  NOR2_X1 U19230 ( .A1(n14696), .A2(n14071), .ZN(n14072) );
  AOI21_X2 U19231 ( .B1(n14074), .B2(n14073), .A(n14072), .ZN(n15801) );
  INV_X1 U19232 ( .A(n15292), .ZN(n15289) );
  OAI21_X1 U19233 ( .B1(n14078), .B2(n14077), .A(n14249), .ZN(n14079) );
  NOR2_X1 U19234 ( .A1(n14080), .A2(n14082), .ZN(n14090) );
  NAND3_X1 U19236 ( .A1(n14085), .A2(n14083), .A3(n14084), .ZN(n14087) );
  INV_X1 U19237 ( .A(n14365), .ZN(n14368) );
  OAI21_X1 U19238 ( .B1(n14094), .B2(n564), .A(n14368), .ZN(n14095) );
  MUX2_X1 U19239 ( .A(n1743), .B(n14262), .S(n14260), .Z(n14100) );
  INV_X1 U19240 ( .A(n14101), .ZN(n14232) );
  NOR2_X1 U19241 ( .A1(n14106), .A2(n14593), .ZN(n14108) );
  INV_X1 U19242 ( .A(n14517), .ZN(n15293) );
  XNOR2_X1 U19243 ( .A(n15801), .B(n29516), .ZN(n16179) );
  NAND2_X1 U19244 ( .A1(n15115), .A2(n14514), .ZN(n14111) );
  NAND2_X1 U19245 ( .A1(n14112), .A2(n14744), .ZN(n14113) );
  NAND2_X1 U19246 ( .A1(n15138), .A2(n15250), .ZN(n14730) );
  INV_X1 U19247 ( .A(n15137), .ZN(n15251) );
  XNOR2_X1 U19248 ( .A(n16329), .B(n16377), .ZN(n14117) );
  XNOR2_X1 U19249 ( .A(n16179), .B(n14117), .ZN(n14225) );
  NAND2_X1 U19250 ( .A1(n14119), .A2(n14118), .ZN(n14124) );
  NAND2_X1 U19251 ( .A1(n14120), .A2(n14365), .ZN(n14121) );
  INV_X1 U19253 ( .A(n14153), .ZN(n15355) );
  OAI211_X1 U19255 ( .C1(n14127), .C2(n14355), .A(n14126), .B(n14125), .ZN(
        n14130) );
  INV_X1 U19256 ( .A(n14752), .ZN(n15243) );
  NAND2_X1 U19257 ( .A1(n14132), .A2(n14131), .ZN(n14133) );
  MUX2_X1 U19258 ( .A(n14134), .B(n14133), .S(n14345), .Z(n14140) );
  NAND2_X1 U19259 ( .A1(n14135), .A2(n14341), .ZN(n14138) );
  NAND2_X1 U19260 ( .A1(n14344), .A2(n14343), .ZN(n14137) );
  MUX2_X1 U19261 ( .A(n14138), .B(n14137), .S(n14136), .Z(n14139) );
  AOI21_X2 U19262 ( .B1(n14144), .B2(n14145), .A(n14143), .ZN(n15060) );
  NOR2_X1 U19263 ( .A1(n15060), .A2(n15355), .ZN(n14149) );
  NAND2_X1 U19264 ( .A1(n13594), .A2(n2849), .ZN(n14147) );
  MUX2_X1 U19265 ( .A(n14150), .B(n13572), .S(n14386), .Z(n14152) );
  NOR2_X1 U19266 ( .A1(n15359), .A2(n14153), .ZN(n14751) );
  XNOR2_X1 U19267 ( .A(n16467), .B(n3516), .ZN(n14223) );
  OAI22_X1 U19268 ( .A1(n29036), .A2(n14491), .B1(n28601), .B2(n14494), .ZN(
        n14156) );
  NAND2_X1 U19269 ( .A1(n14156), .A2(n14493), .ZN(n15344) );
  NAND2_X1 U19270 ( .A1(n14157), .A2(n14480), .ZN(n14476) );
  OAI21_X1 U19271 ( .B1(n293), .B2(n14161), .A(n14476), .ZN(n14160) );
  AND2_X1 U19272 ( .A1(n15222), .A2(n15343), .ZN(n15228) );
  NAND2_X1 U19273 ( .A1(n29565), .A2(n14164), .ZN(n14168) );
  NOR2_X1 U19274 ( .A1(n14757), .A2(n15222), .ZN(n14191) );
  INV_X1 U19275 ( .A(n15342), .ZN(n15225) );
  NAND2_X1 U19276 ( .A1(n14178), .A2(n14451), .ZN(n14179) );
  NAND2_X1 U19277 ( .A1(n14183), .A2(n14182), .ZN(n14190) );
  AOI21_X1 U19278 ( .B1(n14465), .B2(n14185), .A(n14184), .ZN(n14186) );
  NAND2_X1 U19279 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  AOI21_X1 U19280 ( .B1(n12534), .B2(n14426), .A(n29558), .ZN(n14197) );
  NAND2_X1 U19281 ( .A1(n14199), .A2(n14198), .ZN(n15238) );
  NAND2_X1 U19282 ( .A1(n427), .A2(n14456), .ZN(n14202) );
  MUX2_X1 U19283 ( .A(n14202), .B(n14459), .S(n28806), .Z(n14203) );
  INV_X1 U19285 ( .A(n15238), .ZN(n15233) );
  INV_X1 U19286 ( .A(n14206), .ZN(n14209) );
  OAI211_X1 U19287 ( .C1(n14432), .C2(n14437), .A(n1841), .B(n14207), .ZN(
        n14208) );
  NAND3_X1 U19288 ( .A1(n15338), .A2(n15233), .A3(n15334), .ZN(n14222) );
  NAND2_X1 U19289 ( .A1(n14402), .A2(n14399), .ZN(n14211) );
  MUX2_X1 U19290 ( .A(n14211), .B(n14210), .S(n14400), .Z(n14212) );
  INV_X1 U19292 ( .A(n15334), .ZN(n15339) );
  OAI211_X1 U19293 ( .C1(n14216), .C2(n14215), .A(n14214), .B(n29638), .ZN(
        n14219) );
  NAND3_X1 U19294 ( .A1(n14220), .A2(n15339), .A3(n15333), .ZN(n14221) );
  XNOR2_X1 U19295 ( .A(n14225), .B(n14224), .ZN(n17426) );
  MUX2_X1 U19296 ( .A(n14227), .B(n14226), .S(n17426), .Z(n14507) );
  MUX2_X1 U19297 ( .A(n14767), .B(n14713), .S(n14810), .Z(n14228) );
  INV_X1 U19298 ( .A(n14595), .ZN(n14233) );
  INV_X1 U19299 ( .A(n14234), .ZN(n14236) );
  AND2_X1 U19300 ( .A1(n14235), .A2(n14236), .ZN(n14594) );
  OR2_X1 U19301 ( .A1(n14237), .A2(n14252), .ZN(n14596) );
  INV_X1 U19302 ( .A(n14596), .ZN(n14248) );
  OAI21_X1 U19303 ( .B1(n14240), .B2(n14239), .A(n14238), .ZN(n14242) );
  NAND2_X1 U19304 ( .A1(n14242), .A2(n14241), .ZN(n14247) );
  NAND3_X1 U19305 ( .A1(n13943), .A2(n14243), .A3(n15194), .ZN(n14246) );
  MUX2_X1 U19306 ( .A(n14251), .B(n14250), .S(n14249), .Z(n14257) );
  NAND2_X1 U19307 ( .A1(n14253), .A2(n14252), .ZN(n14256) );
  INV_X1 U19308 ( .A(n14254), .ZN(n14255) );
  NOR2_X1 U19309 ( .A1(n14260), .A2(n14259), .ZN(n14263) );
  INV_X1 U19310 ( .A(n14264), .ZN(n14265) );
  OAI22_X1 U19311 ( .A1(n14268), .A2(n14267), .B1(n14266), .B2(n14265), .ZN(
        n14269) );
  NAND2_X1 U19313 ( .A1(n14275), .A2(n14274), .ZN(n14276) );
  NAND2_X1 U19314 ( .A1(n14276), .A2(n14360), .ZN(n14277) );
  NAND2_X1 U19315 ( .A1(n14286), .A2(n14285), .ZN(n14288) );
  INV_X1 U19316 ( .A(n15054), .ZN(n15259) );
  OAI21_X1 U19318 ( .B1(n14298), .B2(n14297), .A(n14296), .ZN(n14606) );
  NAND2_X1 U19319 ( .A1(n15309), .A2(n14851), .ZN(n14340) );
  AND2_X1 U19320 ( .A1(n12534), .A2(n4522), .ZN(n14607) );
  NOR2_X2 U19321 ( .A1(n14610), .A2(n14607), .ZN(n15319) );
  INV_X1 U19322 ( .A(n15319), .ZN(n14854) );
  NAND2_X1 U19323 ( .A1(n14311), .A2(n14313), .ZN(n14316) );
  NOR2_X1 U19324 ( .A1(n14314), .A2(n14313), .ZN(n14315) );
  MUX2_X1 U19325 ( .A(n14319), .B(n14318), .S(n14317), .Z(n14321) );
  NOR2_X1 U19326 ( .A1(n14325), .A2(n14328), .ZN(n14326) );
  NAND2_X1 U19327 ( .A1(n14327), .A2(n14326), .ZN(n14329) );
  AND2_X1 U19328 ( .A1(n14406), .A2(n29133), .ZN(n14409) );
  INV_X1 U19329 ( .A(n14409), .ZN(n14337) );
  NOR2_X1 U19330 ( .A1(n14332), .A2(n14406), .ZN(n14334) );
  OAI21_X1 U19331 ( .B1(n14337), .B2(n1830), .A(n14335), .ZN(n15307) );
  OAI21_X1 U19332 ( .B1(n15309), .B2(n15307), .A(n14851), .ZN(n14338) );
  OAI21_X1 U19333 ( .B1(n14340), .B2(n14854), .A(n14339), .ZN(n16339) );
  INV_X1 U19334 ( .A(n16339), .ZN(n16130) );
  MUX2_X1 U19335 ( .A(n14343), .B(n14342), .S(n14341), .Z(n14348) );
  MUX2_X1 U19336 ( .A(n14345), .B(n14344), .S(n14343), .Z(n14347) );
  MUX2_X2 U19337 ( .A(n14348), .B(n14347), .S(n14346), .Z(n15514) );
  NOR2_X1 U19339 ( .A1(n15274), .A2(n15515), .ZN(n14364) );
  NAND2_X1 U19340 ( .A1(n15510), .A2(n15276), .ZN(n14388) );
  AOI22_X1 U19341 ( .A1(n13725), .A2(n14373), .B1(n14376), .B2(n14372), .ZN(
        n14375) );
  INV_X1 U19342 ( .A(n15511), .ZN(n14918) );
  OAI211_X1 U19344 ( .C1(n14918), .C2(n15274), .A(n14920), .B(n15515), .ZN(
        n14387) );
  XNOR2_X1 U19345 ( .A(n16130), .B(n16443), .ZN(n16028) );
  XNOR2_X1 U19346 ( .A(n16028), .B(n16154), .ZN(n14506) );
  NOR2_X1 U19347 ( .A1(n15285), .A2(n14695), .ZN(n14844) );
  INV_X1 U19348 ( .A(n14844), .ZN(n14390) );
  OAI21_X1 U19349 ( .B1(n6048), .B2(n14842), .A(n14695), .ZN(n14392) );
  XNOR2_X1 U19350 ( .A(n15452), .B(n3528), .ZN(n14504) );
  AOI21_X1 U19352 ( .B1(n14332), .B2(n14406), .A(n14405), .ZN(n14412) );
  INV_X1 U19354 ( .A(n14413), .ZN(n14423) );
  NAND2_X1 U19355 ( .A1(n28648), .A2(n14414), .ZN(n14422) );
  AOI21_X1 U19356 ( .B1(n29638), .B2(n14415), .A(n14414), .ZN(n14418) );
  INV_X1 U19357 ( .A(n14621), .ZN(n14705) );
  NAND2_X1 U19358 ( .A1(n14436), .A2(n14435), .ZN(n14443) );
  NAND3_X1 U19359 ( .A1(n14438), .A2(n14440), .A3(n14437), .ZN(n14442) );
  NAND3_X1 U19360 ( .A1(n1841), .A2(n14440), .A3(n14439), .ZN(n14441) );
  INV_X1 U19361 ( .A(n28647), .ZN(n14445) );
  OR2_X1 U19362 ( .A1(n14446), .A2(n14445), .ZN(n14447) );
  NOR2_X1 U19363 ( .A1(n427), .A2(n14459), .ZN(n14457) );
  OAI21_X1 U19364 ( .B1(n14458), .B2(n14457), .A(n14456), .ZN(n14462) );
  NAND2_X1 U19365 ( .A1(n14460), .A2(n14459), .ZN(n14461) );
  OAI211_X1 U19366 ( .C1(n427), .C2(n14463), .A(n14462), .B(n14461), .ZN(
        n15490) );
  INV_X1 U19367 ( .A(n15490), .ZN(n14702) );
  NAND2_X1 U19368 ( .A1(n14465), .A2(n14464), .ZN(n14468) );
  MUX2_X1 U19369 ( .A(n14471), .B(n14470), .S(n14469), .Z(n14472) );
  NAND2_X1 U19370 ( .A1(n14473), .A2(n14480), .ZN(n14478) );
  NAND3_X1 U19371 ( .A1(n14476), .A2(n14475), .A3(n14474), .ZN(n14477) );
  NAND2_X1 U19373 ( .A1(n15491), .A2(n15485), .ZN(n14917) );
  NAND2_X1 U19374 ( .A1(n29565), .A2(n14481), .ZN(n14482) );
  MUX2_X1 U19375 ( .A(n14483), .B(n14482), .S(n14166), .Z(n14490) );
  NOR2_X1 U19376 ( .A1(n14485), .A2(n14484), .ZN(n14488) );
  AOI22_X1 U19377 ( .A1(n14488), .A2(n14166), .B1(n14487), .B2(n14486), .ZN(
        n14489) );
  NOR2_X1 U19378 ( .A1(n29037), .A2(n14493), .ZN(n14495) );
  AND3_X1 U19379 ( .A1(n29036), .A2(n14498), .A3(n14497), .ZN(n14616) );
  NOR2_X1 U19380 ( .A1(n15490), .A2(n14616), .ZN(n14500) );
  XNOR2_X1 U19381 ( .A(n16653), .B(n16558), .ZN(n16406) );
  XNOR2_X1 U19382 ( .A(n16406), .B(n14504), .ZN(n14505) );
  XNOR2_X1 U19383 ( .A(n14505), .B(n14506), .ZN(n17424) );
  OAI21_X1 U19385 ( .B1(n15138), .B2(n15246), .A(n15252), .ZN(n14511) );
  INV_X1 U19387 ( .A(n15250), .ZN(n15136) );
  NAND3_X1 U19388 ( .A1(n15135), .A2(n15136), .A3(n15248), .ZN(n14509) );
  NOR2_X1 U19390 ( .A1(n14514), .A2(n15117), .ZN(n14742) );
  NAND2_X1 U19391 ( .A1(n14742), .A2(n15115), .ZN(n14515) );
  OR2_X1 U19392 ( .A1(n15215), .A2(n15292), .ZN(n14522) );
  NAND3_X1 U19393 ( .A1(n15036), .A2(n15290), .A3(n14517), .ZN(n14519) );
  NAND4_X2 U19394 ( .A1(n14522), .A2(n14521), .A3(n14520), .A4(n14519), .ZN(
        n16262) );
  XNOR2_X1 U19395 ( .A(n16262), .B(n72), .ZN(n14523) );
  INV_X1 U19396 ( .A(n15224), .ZN(n15348) );
  MUX2_X1 U19397 ( .A(n15225), .B(n15348), .S(n15046), .Z(n14525) );
  NAND2_X1 U19399 ( .A1(n15338), .A2(n15333), .ZN(n14526) );
  AND3_X1 U19400 ( .A1(n15238), .A2(n14526), .A3(n14781), .ZN(n14527) );
  INV_X1 U19401 ( .A(n16024), .ZN(n14529) );
  XNOR2_X1 U19402 ( .A(n14529), .B(n16405), .ZN(n15893) );
  NAND3_X1 U19403 ( .A1(n15183), .A2(n552), .A3(n14785), .ZN(n14530) );
  NAND3_X1 U19404 ( .A1(n553), .A2(n15457), .A3(n15174), .ZN(n14538) );
  NOR2_X1 U19405 ( .A1(n15456), .A2(n15174), .ZN(n15458) );
  NAND3_X1 U19406 ( .A1(n15180), .A2(n15174), .A3(n28803), .ZN(n14536) );
  NAND3_X1 U19407 ( .A1(n14534), .A2(n5635), .A3(n15456), .ZN(n14535) );
  XNOR2_X1 U19408 ( .A(n16052), .B(n15927), .ZN(n16311) );
  NAND3_X1 U19409 ( .A1(n15202), .A2(n15204), .A3(n14967), .ZN(n14543) );
  NOR2_X1 U19410 ( .A1(n15202), .A2(n15208), .ZN(n14539) );
  AND2_X1 U19411 ( .A1(n15207), .A2(n15208), .ZN(n14964) );
  NAND2_X1 U19412 ( .A1(n15209), .A2(n14960), .ZN(n14540) );
  NAND3_X2 U19413 ( .A1(n14542), .A2(n14543), .A3(n14541), .ZN(n16247) );
  XNOR2_X1 U19414 ( .A(n16247), .B(n5059), .ZN(n14544) );
  XNOR2_X1 U19415 ( .A(n16311), .B(n14544), .ZN(n14562) );
  INV_X1 U19416 ( .A(n15466), .ZN(n15159) );
  NAND2_X1 U19417 ( .A1(n15159), .A2(n15463), .ZN(n14546) );
  NOR3_X1 U19418 ( .A1(n15462), .A2(n14652), .A3(n29153), .ZN(n14545) );
  NAND2_X1 U19420 ( .A1(n15168), .A2(n15474), .ZN(n15170) );
  INV_X1 U19421 ( .A(n15167), .ZN(n14958) );
  NAND3_X1 U19422 ( .A1(n15166), .A2(n14551), .A3(n1848), .ZN(n14552) );
  OAI211_X1 U19423 ( .C1(n1809), .C2(n15170), .A(n14553), .B(n14552), .ZN(
        n16435) );
  INV_X1 U19424 ( .A(n16435), .ZN(n14554) );
  XNOR2_X1 U19425 ( .A(n14554), .B(n16603), .ZN(n16343) );
  NOR2_X1 U19426 ( .A1(n14810), .A2(n14713), .ZN(n14559) );
  INV_X1 U19427 ( .A(n14713), .ZN(n14766) );
  OAI21_X1 U19428 ( .B1(n14767), .B2(n14766), .A(n13922), .ZN(n14558) );
  NAND2_X1 U19429 ( .A1(n14559), .A2(n14715), .ZN(n14557) );
  NAND2_X1 U19430 ( .A1(n14775), .A2(n14555), .ZN(n14556) );
  XNOR2_X1 U19431 ( .A(n16618), .B(n16312), .ZN(n14560) );
  XNOR2_X1 U19432 ( .A(n16343), .B(n14560), .ZN(n14561) );
  NAND2_X1 U19433 ( .A1(n15690), .A2(n15083), .ZN(n14877) );
  AND2_X1 U19434 ( .A1(n14877), .A2(n14563), .ZN(n14565) );
  NAND2_X1 U19435 ( .A1(n14670), .A2(n323), .ZN(n14564) );
  OAI21_X1 U19436 ( .B1(n15692), .B2(n14565), .A(n14564), .ZN(n14568) );
  NOR2_X1 U19437 ( .A1(n15084), .A2(n14566), .ZN(n14567) );
  NOR2_X1 U19438 ( .A1(n14568), .A2(n14567), .ZN(n14921) );
  INV_X1 U19439 ( .A(n15082), .ZN(n14574) );
  INV_X1 U19441 ( .A(n15077), .ZN(n15075) );
  OR2_X1 U19442 ( .A1(n14948), .A2(n15077), .ZN(n14872) );
  NAND2_X1 U19443 ( .A1(n14872), .A2(n14571), .ZN(n14573) );
  INV_X1 U19445 ( .A(n16320), .ZN(n14581) );
  OAI21_X1 U19446 ( .B1(n15420), .B2(n15101), .A(n4549), .ZN(n14576) );
  AOI21_X1 U19447 ( .B1(n14903), .B2(n15097), .A(n14578), .ZN(n14580) );
  XNOR2_X1 U19448 ( .A(n14581), .B(n15903), .ZN(n14592) );
  NAND2_X1 U19449 ( .A1(n14881), .A2(n13789), .ZN(n14585) );
  XNOR2_X1 U19450 ( .A(n29319), .B(n16256), .ZN(n14590) );
  NAND2_X1 U19451 ( .A1(n15406), .A2(n14894), .ZN(n14939) );
  INV_X1 U19452 ( .A(n15407), .ZN(n15416) );
  AOI21_X1 U19453 ( .B1(n14940), .B2(n14939), .A(n15416), .ZN(n14588) );
  NAND2_X1 U19454 ( .A1(n15415), .A2(n15409), .ZN(n14586) );
  AOI21_X1 U19455 ( .B1(n14586), .B2(n14893), .A(n14894), .ZN(n14587) );
  XNOR2_X1 U19456 ( .A(n16257), .B(n3728), .ZN(n14589) );
  XNOR2_X1 U19457 ( .A(n14590), .B(n14589), .ZN(n14591) );
  INV_X1 U19459 ( .A(n29297), .ZN(n16996) );
  INV_X1 U19460 ( .A(n14762), .ZN(n15056) );
  NAND2_X1 U19461 ( .A1(n14597), .A2(n14596), .ZN(n15053) );
  NAND2_X1 U19462 ( .A1(n15053), .A2(n14761), .ZN(n14598) );
  NAND3_X1 U19463 ( .A1(n15055), .A2(n15261), .A3(n14763), .ZN(n14599) );
  INV_X1 U19464 ( .A(n15366), .ZN(n14603) );
  NOR2_X1 U19466 ( .A1(n15274), .A2(n15511), .ZN(n14605) );
  NOR2_X1 U19467 ( .A1(n15514), .A2(n14697), .ZN(n14604) );
  INV_X1 U19468 ( .A(n15307), .ZN(n15308) );
  INV_X1 U19469 ( .A(n15306), .ZN(n15312) );
  OAI21_X1 U19470 ( .B1(n15312), .B2(n15310), .A(n14851), .ZN(n14613) );
  INV_X1 U19471 ( .A(n14606), .ZN(n14609) );
  INV_X1 U19472 ( .A(n14607), .ZN(n14608) );
  NAND3_X1 U19473 ( .A1(n1096), .A2(n14609), .A3(n14608), .ZN(n14611) );
  OAI21_X1 U19474 ( .B1(n14611), .B2(n14610), .A(n15311), .ZN(n14612) );
  NAND2_X1 U19476 ( .A1(n14702), .A2(n15485), .ZN(n14617) );
  INV_X1 U19478 ( .A(n15489), .ZN(n15486) );
  NAND3_X1 U19479 ( .A1(n15486), .A2(n14702), .A3(n14703), .ZN(n14619) );
  NOR2_X1 U19480 ( .A1(n15503), .A2(n15265), .ZN(n14623) );
  AOI22_X1 U19481 ( .A1(n14623), .A2(n15502), .B1(n14622), .B2(n15500), .ZN(
        n14627) );
  INV_X1 U19482 ( .A(n15506), .ZN(n14625) );
  INV_X1 U19483 ( .A(n14623), .ZN(n14624) );
  OAI211_X1 U19484 ( .C1(n14625), .C2(n15497), .A(n14624), .B(n14922), .ZN(
        n14626) );
  XNOR2_X1 U19485 ( .A(n16399), .B(n16043), .ZN(n16367) );
  XNOR2_X1 U19486 ( .A(n16278), .B(n16367), .ZN(n14628) );
  NOR2_X1 U19487 ( .A1(n14992), .A2(n15394), .ZN(n14632) );
  AOI22_X1 U19488 ( .A1(n15395), .A2(n14632), .B1(n15391), .B2(n14631), .ZN(
        n14635) );
  MUX2_X1 U19491 ( .A(n15382), .B(n15152), .S(n14986), .Z(n14638) );
  OR2_X1 U19492 ( .A1(n15382), .A2(n15151), .ZN(n15154) );
  NAND3_X1 U19493 ( .A1(n15382), .A2(n14986), .A3(n15150), .ZN(n14636) );
  AND2_X1 U19494 ( .A1(n15154), .A2(n14636), .ZN(n14637) );
  OAI21_X1 U19495 ( .B1(n14638), .B2(n15155), .A(n14637), .ZN(n16426) );
  XNOR2_X1 U19496 ( .A(n16426), .B(n16567), .ZN(n16362) );
  INV_X1 U19497 ( .A(n16362), .ZN(n14643) );
  OAI21_X1 U19498 ( .B1(n15077), .B2(n15072), .A(n15081), .ZN(n14640) );
  XNOR2_X1 U19499 ( .A(n16272), .B(n16295), .ZN(n15426) );
  INV_X1 U19500 ( .A(n15426), .ZN(n14642) );
  XNOR2_X1 U19501 ( .A(n14643), .B(n14642), .ZN(n14656) );
  NAND3_X1 U19502 ( .A1(n15184), .A2(n15183), .A3(n15190), .ZN(n14648) );
  INV_X1 U19503 ( .A(n15183), .ZN(n14644) );
  NAND3_X1 U19504 ( .A1(n15186), .A2(n14644), .A3(n15185), .ZN(n14647) );
  NAND2_X1 U19505 ( .A1(n14645), .A2(n14644), .ZN(n14646) );
  NAND3_X1 U19507 ( .A1(n3784), .A2(n6879), .A3(n15370), .ZN(n14651) );
  NOR2_X1 U19508 ( .A1(n15372), .A2(n14863), .ZN(n14650) );
  XNOR2_X1 U19509 ( .A(n15817), .B(n16294), .ZN(n14654) );
  XNOR2_X1 U19510 ( .A(n321), .B(n2889), .ZN(n14653) );
  XNOR2_X1 U19511 ( .A(n14654), .B(n14653), .ZN(n14655) );
  OAI21_X1 U19512 ( .B1(n16863), .B2(n16996), .A(n16991), .ZN(n14694) );
  NOR2_X1 U19513 ( .A1(n16992), .A2(n17269), .ZN(n14693) );
  NOR2_X1 U19514 ( .A1(n15438), .A2(n15436), .ZN(n15020) );
  INV_X1 U19515 ( .A(n14658), .ZN(n14663) );
  INV_X1 U19516 ( .A(n14659), .ZN(n14662) );
  NAND2_X1 U19518 ( .A1(n14670), .A2(n28666), .ZN(n14672) );
  OAI211_X1 U19519 ( .C1(n323), .C2(n15691), .A(n15087), .B(n15689), .ZN(
        n14671) );
  XNOR2_X1 U19520 ( .A(n28597), .B(n16641), .ZN(n14676) );
  NAND2_X1 U19521 ( .A1(n15321), .A2(n15013), .ZN(n15326) );
  INV_X1 U19522 ( .A(n15013), .ZN(n15445) );
  OAI211_X1 U19523 ( .C1(n15014), .C2(n15015), .A(n15322), .B(n15445), .ZN(
        n14674) );
  NAND2_X1 U19524 ( .A1(n1926), .A2(n15014), .ZN(n14673) );
  XNOR2_X1 U19525 ( .A(n14676), .B(n14675), .ZN(n14692) );
  INV_X1 U19526 ( .A(n15094), .ZN(n14680) );
  AOI21_X1 U19527 ( .B1(n3315), .B2(n14680), .A(n14679), .ZN(n14681) );
  INV_X1 U19528 ( .A(n14824), .ZN(n15032) );
  INV_X1 U19529 ( .A(n15029), .ZN(n14684) );
  XNOR2_X1 U19530 ( .A(n15909), .B(n15802), .ZN(n16331) );
  NAND2_X1 U19531 ( .A1(n14685), .A2(n15000), .ZN(n14690) );
  INV_X1 U19532 ( .A(n15132), .ZN(n14689) );
  XNOR2_X1 U19533 ( .A(n16329), .B(n16238), .ZN(n16082) );
  XNOR2_X1 U19534 ( .A(n16082), .B(n16331), .ZN(n14691) );
  XNOR2_X1 U19535 ( .A(n14692), .B(n14691), .ZN(n16995) );
  XNOR2_X1 U19536 ( .A(n16563), .B(n1911), .ZN(n14701) );
  NAND2_X1 U19537 ( .A1(n14698), .A2(n15512), .ZN(n14699) );
  NAND3_X1 U19538 ( .A1(n15309), .A2(n15312), .A3(n15307), .ZN(n14700) );
  XNOR2_X1 U19539 ( .A(n16216), .B(n16421), .ZN(n16536) );
  XNOR2_X1 U19540 ( .A(n16536), .B(n14701), .ZN(n14721) );
  INV_X1 U19541 ( .A(n15494), .ZN(n15269) );
  AND2_X1 U19542 ( .A1(n14922), .A2(n15503), .ZN(n14707) );
  INV_X1 U19544 ( .A(n16185), .ZN(n14709) );
  INV_X1 U19545 ( .A(n16270), .ZN(n15878) );
  INV_X1 U19546 ( .A(n15053), .ZN(n15262) );
  NOR2_X1 U19547 ( .A1(n15262), .A2(n15260), .ZN(n14710) );
  INV_X1 U19549 ( .A(n16568), .ZN(n14719) );
  INV_X1 U19550 ( .A(n14712), .ZN(n14714) );
  AOI21_X1 U19551 ( .B1(n14714), .B2(n14713), .A(n14810), .ZN(n14718) );
  NAND2_X1 U19552 ( .A1(n14810), .A2(n28493), .ZN(n14716) );
  AOI21_X1 U19553 ( .B1(n14811), .B2(n14716), .A(n14773), .ZN(n14717) );
  XNOR2_X1 U19554 ( .A(n15878), .B(n16145), .ZN(n14720) );
  NAND2_X1 U19555 ( .A1(n15387), .A2(n15388), .ZN(n14728) );
  NAND2_X1 U19556 ( .A1(n15395), .A2(n14722), .ZN(n14727) );
  NAND2_X1 U19557 ( .A1(n15389), .A2(n3210), .ZN(n14725) );
  INV_X1 U19558 ( .A(n15389), .ZN(n15145) );
  OAI21_X1 U19559 ( .B1(n15387), .B2(n15144), .A(n15145), .ZN(n14724) );
  OAI211_X1 U19560 ( .C1(n14990), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        n14726) );
  NAND3_X1 U19561 ( .A1(n15252), .A2(n15138), .A3(n15246), .ZN(n14731) );
  XNOR2_X1 U19562 ( .A(n16280), .B(n543), .ZN(n15863) );
  INV_X1 U19563 ( .A(n15863), .ZN(n14736) );
  NAND2_X1 U19564 ( .A1(n28196), .A2(n28518), .ZN(n15399) );
  XNOR2_X1 U19565 ( .A(n16365), .B(n1225), .ZN(n14735) );
  XNOR2_X1 U19566 ( .A(n14736), .B(n14735), .ZN(n14749) );
  MUX2_X1 U19567 ( .A(n15155), .B(n15382), .S(n15383), .Z(n14739) );
  NOR2_X1 U19568 ( .A1(n14740), .A2(n1904), .ZN(n14741) );
  NAND2_X1 U19569 ( .A1(n15115), .A2(n14743), .ZN(n14745) );
  NAND2_X1 U19570 ( .A1(n15000), .A2(n15127), .ZN(n14747) );
  XNOR2_X1 U19571 ( .A(n16116), .B(n16506), .ZN(n14748) );
  OAI21_X1 U19573 ( .B1(n15060), .B2(n14753), .A(n15359), .ZN(n14754) );
  AND2_X1 U19575 ( .A1(n15343), .A2(n15342), .ZN(n14756) );
  NAND2_X1 U19576 ( .A1(n15226), .A2(n14756), .ZN(n14759) );
  AOI22_X1 U19577 ( .A1(n14757), .A2(n15223), .B1(n15348), .B2(n15343), .ZN(
        n14758) );
  INV_X1 U19578 ( .A(n16578), .ZN(n14760) );
  XNOR2_X1 U19579 ( .A(n14760), .B(n16495), .ZN(n16124) );
  OAI21_X1 U19580 ( .B1(n14810), .B2(n14767), .A(n14766), .ZN(n14768) );
  NAND2_X1 U19581 ( .A1(n14768), .A2(n13922), .ZN(n14777) );
  INV_X1 U19582 ( .A(n14772), .ZN(n14774) );
  XNOR2_X1 U19583 ( .A(n16416), .B(n16012), .ZN(n16497) );
  INV_X1 U19584 ( .A(n16497), .ZN(n14778) );
  XNOR2_X1 U19585 ( .A(n14778), .B(n16124), .ZN(n14791) );
  XNOR2_X1 U19586 ( .A(n16579), .B(n3586), .ZN(n14789) );
  INV_X1 U19587 ( .A(n15239), .ZN(n15235) );
  NAND3_X1 U19588 ( .A1(n15234), .A2(n15338), .A3(n15334), .ZN(n14782) );
  INV_X1 U19589 ( .A(n14784), .ZN(n14783) );
  AOI21_X1 U19590 ( .B1(n15184), .B2(n15185), .A(n14783), .ZN(n14788) );
  OAI21_X1 U19591 ( .B1(n14785), .B2(n15182), .A(n14799), .ZN(n14786) );
  NAND2_X1 U19592 ( .A1(n14786), .A2(n15183), .ZN(n14787) );
  XNOR2_X1 U19593 ( .A(n16321), .B(n16077), .ZN(n16253) );
  XNOR2_X1 U19594 ( .A(n14789), .B(n16253), .ZN(n14790) );
  XNOR2_X1 U19595 ( .A(n14791), .B(n14790), .ZN(n14871) );
  OAI211_X1 U19596 ( .C1(n14881), .C2(n13789), .A(n14793), .B(n5813), .ZN(
        n14794) );
  AOI22_X1 U19597 ( .A1(n15459), .A2(n15174), .B1(n15456), .B2(n28803), .ZN(
        n15461) );
  OAI211_X1 U19598 ( .C1(n14534), .C2(n28803), .A(n28462), .B(n15457), .ZN(
        n14798) );
  XNOR2_X1 U19599 ( .A(n28585), .B(n15760), .ZN(n16514) );
  XNOR2_X1 U19600 ( .A(n16119), .B(n16514), .ZN(n14815) );
  INV_X1 U19601 ( .A(n15171), .ZN(n15475) );
  NAND2_X1 U19602 ( .A1(n15475), .A2(n15476), .ZN(n15473) );
  OAI211_X1 U19603 ( .C1(n15166), .C2(n15168), .A(n15171), .B(n14958), .ZN(
        n14801) );
  NAND2_X1 U19604 ( .A1(n545), .A2(n15462), .ZN(n15164) );
  INV_X1 U19605 ( .A(n15164), .ZN(n14804) );
  NAND2_X1 U19606 ( .A1(n14802), .A2(n15161), .ZN(n14803) );
  AOI21_X1 U19607 ( .B1(n14808), .B2(n14807), .A(n28493), .ZN(n14809) );
  XNOR2_X1 U19608 ( .A(n16586), .B(n135), .ZN(n14813) );
  XNOR2_X1 U19609 ( .A(n16243), .B(n14813), .ZN(n14814) );
  XNOR2_X1 U19610 ( .A(n14815), .B(n14814), .ZN(n16999) );
  MUX2_X1 U19611 ( .A(n29572), .B(n14871), .S(n16999), .Z(n14915) );
  AND3_X1 U19612 ( .A1(n15437), .A2(n15438), .A3(n15300), .ZN(n14816) );
  AOI21_X1 U19613 ( .B1(n15444), .B2(n15302), .A(n14816), .ZN(n14820) );
  INV_X1 U19614 ( .A(n15300), .ZN(n15440) );
  OAI21_X1 U19615 ( .B1(n15444), .B2(n15436), .A(n15440), .ZN(n14819) );
  INV_X1 U19616 ( .A(n15303), .ZN(n14817) );
  NOR2_X1 U19617 ( .A1(n14817), .A2(n15022), .ZN(n14818) );
  NOR2_X1 U19618 ( .A1(n14821), .A2(n14826), .ZN(n14822) );
  NAND2_X1 U19619 ( .A1(n15032), .A2(n14825), .ZN(n14827) );
  AOI21_X1 U19620 ( .B1(n15433), .B2(n14827), .A(n15430), .ZN(n14828) );
  NOR2_X1 U19621 ( .A1(n14832), .A2(n14831), .ZN(n14835) );
  OAI21_X1 U19622 ( .B1(n14837), .B2(n15294), .A(n14836), .ZN(n14840) );
  INV_X1 U19623 ( .A(n15291), .ZN(n15037) );
  OAI21_X1 U19624 ( .B1(n15215), .B2(n15037), .A(n14838), .ZN(n14839) );
  INV_X1 U19625 ( .A(n15284), .ZN(n14841) );
  NOR2_X1 U19626 ( .A1(n28996), .A2(n14842), .ZN(n14843) );
  XNOR2_X1 U19627 ( .A(n16017), .B(n15887), .ZN(n16524) );
  INV_X1 U19628 ( .A(n16524), .ZN(n14850) );
  INV_X1 U19629 ( .A(n15309), .ZN(n14852) );
  NAND3_X1 U19630 ( .A1(n14854), .A2(n14851), .A3(n14852), .ZN(n14858) );
  NOR2_X1 U19631 ( .A1(n14852), .A2(n15310), .ZN(n14853) );
  NAND2_X1 U19632 ( .A1(n14854), .A2(n14853), .ZN(n14857) );
  NAND3_X1 U19633 ( .A1(n15310), .A2(n15311), .A3(n15306), .ZN(n14856) );
  NAND3_X1 U19634 ( .A1(n15322), .A2(n546), .A3(n15321), .ZN(n14862) );
  NAND3_X1 U19635 ( .A1(n15447), .A2(n15321), .A3(n15014), .ZN(n14861) );
  INV_X1 U19636 ( .A(n15321), .ZN(n15446) );
  NAND3_X1 U19637 ( .A1(n15446), .A2(n546), .A3(n15445), .ZN(n14860) );
  INV_X1 U19638 ( .A(n15014), .ZN(n15448) );
  NAND3_X1 U19639 ( .A1(n1926), .A2(n15448), .A3(n15015), .ZN(n14859) );
  XNOR2_X1 U19640 ( .A(n16165), .B(n16313), .ZN(n16249) );
  NOR2_X1 U19641 ( .A1(n15009), .A2(n14863), .ZN(n14864) );
  OAI21_X1 U19642 ( .B1(n14865), .B2(n14864), .A(n15373), .ZN(n14866) );
  XNOR2_X1 U19643 ( .A(n16249), .B(n14868), .ZN(n14869) );
  XNOR2_X1 U19644 ( .A(n14870), .B(n14869), .ZN(n17396) );
  OAI21_X1 U19645 ( .B1(n15073), .B2(n15072), .A(n14872), .ZN(n14873) );
  NAND2_X1 U19646 ( .A1(n14873), .A2(n15071), .ZN(n14875) );
  AND2_X1 U19647 ( .A1(n15072), .A2(n14874), .ZN(n15078) );
  MUX2_X1 U19648 ( .A(n323), .B(n15690), .S(n15692), .Z(n14880) );
  NAND2_X1 U19649 ( .A1(n14878), .A2(n14877), .ZN(n14879) );
  XNOR2_X1 U19650 ( .A(n15849), .B(n15982), .ZN(n16518) );
  INV_X1 U19651 ( .A(n16518), .ZN(n14892) );
  NAND2_X1 U19652 ( .A1(n14882), .A2(n14881), .ZN(n14883) );
  NAND2_X1 U19653 ( .A1(n14883), .A2(n388), .ZN(n14889) );
  NOR2_X1 U19654 ( .A1(n14884), .A2(n5813), .ZN(n14888) );
  NAND3_X1 U19655 ( .A1(n14886), .A2(n13789), .A3(n14885), .ZN(n14887) );
  XNOR2_X1 U19656 ( .A(n16131), .B(n14890), .ZN(n14891) );
  XNOR2_X1 U19657 ( .A(n14892), .B(n14891), .ZN(n14914) );
  NAND2_X1 U19658 ( .A1(n14895), .A2(n28196), .ZN(n14899) );
  NAND2_X1 U19659 ( .A1(n14944), .A2(n15402), .ZN(n14897) );
  OAI211_X1 U19660 ( .C1(n28196), .C2(n15398), .A(n14899), .B(n14898), .ZN(
        n16409) );
  XNOR2_X1 U19661 ( .A(n16409), .B(n16556), .ZN(n16134) );
  NAND2_X1 U19662 ( .A1(n14903), .A2(n14901), .ZN(n15096) );
  NAND3_X1 U19663 ( .A1(n15096), .A2(n15099), .A3(n15100), .ZN(n14911) );
  NAND2_X1 U19664 ( .A1(n14908), .A2(n14907), .ZN(n14909) );
  OAI211_X1 U19665 ( .C1(n15095), .C2(n15094), .A(n3315), .B(n14909), .ZN(
        n14910) );
  XNOR2_X1 U19666 ( .A(n16070), .B(n2946), .ZN(n14912) );
  XNOR2_X1 U19667 ( .A(n16134), .B(n14912), .ZN(n14913) );
  INV_X1 U19668 ( .A(n17397), .ZN(n17402) );
  INV_X1 U19669 ( .A(n16498), .ZN(n15855) );
  NAND2_X1 U19670 ( .A1(n15510), .A2(n14918), .ZN(n14919) );
  XNOR2_X1 U19673 ( .A(n16455), .B(n16038), .ZN(n14931) );
  NAND2_X1 U19674 ( .A1(n14927), .A2(n14967), .ZN(n14929) );
  XNOR2_X1 U19675 ( .A(n15654), .B(n3109), .ZN(n14930) );
  XNOR2_X1 U19676 ( .A(n14931), .B(n14930), .ZN(n14932) );
  INV_X1 U19677 ( .A(n15802), .ZN(n14933) );
  XNOR2_X1 U19678 ( .A(n14933), .B(n16509), .ZN(n14941) );
  INV_X1 U19679 ( .A(n15101), .ZN(n15417) );
  OAI211_X1 U19680 ( .C1(n15407), .C2(n15406), .A(n14937), .B(n15410), .ZN(
        n14938) );
  XNOR2_X1 U19681 ( .A(n15583), .B(n16241), .ZN(n15948) );
  XNOR2_X1 U19682 ( .A(n15948), .B(n14941), .ZN(n14955) );
  XNOR2_X1 U19683 ( .A(n16641), .B(n2916), .ZN(n14953) );
  NOR2_X1 U19684 ( .A1(n15401), .A2(n28518), .ZN(n14947) );
  NAND2_X1 U19685 ( .A1(n14945), .A2(n15399), .ZN(n14946) );
  AOI21_X1 U19686 ( .B1(n14949), .B2(n15071), .A(n15076), .ZN(n14951) );
  XNOR2_X1 U19688 ( .A(n15949), .B(n15999), .ZN(n16639) );
  XNOR2_X1 U19689 ( .A(n16639), .B(n14953), .ZN(n14954) );
  AOI22_X1 U19690 ( .A1(n15475), .A2(n14958), .B1(n1850), .B2(n15168), .ZN(
        n14956) );
  MUX2_X1 U19691 ( .A(n14956), .B(n15170), .S(n15166), .Z(n14957) );
  NOR2_X1 U19693 ( .A1(n15208), .A2(n14960), .ZN(n14962) );
  AOI22_X1 U19694 ( .A1(n14963), .A2(n15208), .B1(n14962), .B2(n14961), .ZN(
        n14966) );
  XNOR2_X1 U19696 ( .A(n16296), .B(n16534), .ZN(n15944) );
  XNOR2_X1 U19697 ( .A(n321), .B(n3537), .ZN(n14978) );
  NAND2_X1 U19698 ( .A1(n14972), .A2(n14971), .ZN(n14973) );
  AOI21_X2 U19700 ( .B1(n14977), .B2(n14976), .A(n14975), .ZN(n16211) );
  XNOR2_X1 U19701 ( .A(n14978), .B(n16211), .ZN(n14979) );
  XNOR2_X1 U19702 ( .A(n14979), .B(n15944), .ZN(n14985) );
  NAND2_X1 U19703 ( .A1(n15180), .A2(n15174), .ZN(n14982) );
  INV_X1 U19704 ( .A(n16422), .ZN(n14983) );
  MUX2_X1 U19705 ( .A(n15383), .B(n15151), .S(n15382), .Z(n14988) );
  MUX2_X1 U19706 ( .A(n15382), .B(n14986), .S(n15379), .Z(n14987) );
  NOR2_X1 U19707 ( .A1(n15394), .A2(n15388), .ZN(n14991) );
  XNOR2_X1 U19708 ( .A(n16023), .B(n3422), .ZN(n14996) );
  INV_X1 U19709 ( .A(n16409), .ZN(n14995) );
  XNOR2_X1 U19710 ( .A(n14996), .B(n14995), .ZN(n14997) );
  INV_X1 U19711 ( .A(n14999), .ZN(n15005) );
  NAND2_X1 U19712 ( .A1(n15001), .A2(n15000), .ZN(n15002) );
  NOR2_X1 U19713 ( .A1(n15002), .A2(n15132), .ZN(n15003) );
  AOI21_X1 U19714 ( .B1(n15005), .B2(n15004), .A(n15003), .ZN(n15006) );
  XNOR2_X1 U19715 ( .A(n15007), .B(n15772), .ZN(n15986) );
  XNOR2_X1 U19716 ( .A(n15986), .B(n2206), .ZN(n16658) );
  XNOR2_X1 U19717 ( .A(n16393), .B(n15011), .ZN(n15026) );
  AND2_X1 U19718 ( .A1(n15447), .A2(n15445), .ZN(n15012) );
  NAND2_X1 U19719 ( .A1(n15320), .A2(n546), .ZN(n15017) );
  NOR2_X1 U19720 ( .A1(n15022), .A2(n15301), .ZN(n15019) );
  NOR2_X1 U19721 ( .A1(n15020), .A2(n15019), .ZN(n15021) );
  NAND2_X1 U19722 ( .A1(n15021), .A2(n15444), .ZN(n15024) );
  NOR2_X1 U19723 ( .A1(n15438), .A2(n15022), .ZN(n15435) );
  NAND2_X1 U19724 ( .A1(n15435), .A2(n15440), .ZN(n15023) );
  XNOR2_X1 U19725 ( .A(n15026), .B(n15965), .ZN(n15044) );
  NAND3_X1 U19727 ( .A1(n15037), .A2(n15036), .A3(n15293), .ZN(n15038) );
  XNOR2_X1 U19729 ( .A(n15042), .B(n16232), .ZN(n16633) );
  INV_X1 U19730 ( .A(n16633), .ZN(n15043) );
  INV_X1 U19731 ( .A(n15338), .ZN(n15052) );
  XNOR2_X1 U19736 ( .A(n15780), .B(n16618), .ZN(n15057) );
  XNOR2_X1 U19737 ( .A(n15973), .B(n15057), .ZN(n15068) );
  INV_X1 U19738 ( .A(n15359), .ZN(n15245) );
  NOR3_X1 U19740 ( .A1(n15245), .A2(n15361), .A3(n28197), .ZN(n15059) );
  NOR3_X1 U19741 ( .A1(n15359), .A2(n14752), .A3(n15355), .ZN(n15058) );
  NOR2_X1 U19742 ( .A1(n15059), .A2(n15058), .ZN(n15064) );
  NOR2_X1 U19743 ( .A1(n15060), .A2(n15360), .ZN(n15061) );
  XNOR2_X1 U19745 ( .A(n16619), .B(n2385), .ZN(n15066) );
  XNOR2_X1 U19746 ( .A(n16526), .B(n16052), .ZN(n15065) );
  XNOR2_X1 U19747 ( .A(n15066), .B(n15065), .ZN(n15067) );
  NAND3_X1 U19748 ( .A1(n17435), .A2(n17438), .A3(n17440), .ZN(n15069) );
  INV_X1 U19749 ( .A(n18304), .ZN(n18475) );
  XNOR2_X1 U19750 ( .A(n15070), .B(n2403), .ZN(n15093) );
  NOR2_X1 U19751 ( .A1(n15072), .A2(n15071), .ZN(n15074) );
  NAND2_X1 U19752 ( .A1(n15078), .A2(n15077), .ZN(n15079) );
  NOR2_X1 U19753 ( .A1(n15084), .A2(n15083), .ZN(n15091) );
  OAI21_X1 U19754 ( .B1(n15692), .B2(n323), .A(n15691), .ZN(n15090) );
  XNOR2_X1 U19756 ( .A(n16598), .B(n15093), .ZN(n15112) );
  NAND2_X1 U19757 ( .A1(n15102), .A2(n15101), .ZN(n15104) );
  INV_X1 U19758 ( .A(n16191), .ZN(n15110) );
  NAND2_X1 U19759 ( .A1(n15410), .A2(n15107), .ZN(n15109) );
  XNOR2_X1 U19760 ( .A(n16365), .B(n16398), .ZN(n15741) );
  XNOR2_X1 U19761 ( .A(n15110), .B(n15741), .ZN(n15111) );
  INV_X1 U19762 ( .A(n17304), .ZN(n17305) );
  XNOR2_X1 U19763 ( .A(n16477), .B(n2509), .ZN(n15133) );
  AND2_X1 U19764 ( .A1(n15116), .A2(n15115), .ZN(n15118) );
  NOR2_X1 U19766 ( .A1(n13632), .A2(n15123), .ZN(n15124) );
  AOI22_X1 U19767 ( .A1(n15126), .A2(n15125), .B1(n15124), .B2(n1744), .ZN(
        n15130) );
  NOR2_X1 U19768 ( .A1(n551), .A2(n15127), .ZN(n15128) );
  NAND2_X1 U19769 ( .A1(n15132), .A2(n15128), .ZN(n15129) );
  XNOR2_X1 U19770 ( .A(n15133), .B(n16140), .ZN(n15158) );
  INV_X1 U19771 ( .A(n15246), .ZN(n15134) );
  OAI21_X1 U19772 ( .B1(n15249), .B2(n15135), .A(n15134), .ZN(n15143) );
  AND2_X1 U19773 ( .A1(n15135), .A2(n15138), .ZN(n15142) );
  NAND2_X1 U19774 ( .A1(n15246), .A2(n15136), .ZN(n15140) );
  NAND2_X1 U19775 ( .A1(n15138), .A2(n15137), .ZN(n15139) );
  MUX2_X1 U19776 ( .A(n15140), .B(n15139), .S(n14733), .Z(n15141) );
  OAI21_X1 U19777 ( .B1(n15143), .B2(n15142), .A(n15141), .ZN(n16620) );
  MUX2_X1 U19778 ( .A(n15388), .B(n15389), .S(n15144), .Z(n15146) );
  NOR3_X1 U19779 ( .A1(n15395), .A2(n15391), .A3(n15387), .ZN(n15148) );
  INV_X1 U19780 ( .A(n16196), .ZN(n15156) );
  NAND3_X1 U19781 ( .A1(n15155), .A2(n15152), .A3(n15384), .ZN(n15153) );
  XNOR2_X1 U19782 ( .A(n15156), .B(n16050), .ZN(n15157) );
  AND2_X1 U19783 ( .A1(n15161), .A2(n29153), .ZN(n15162) );
  NOR2_X1 U19784 ( .A1(n15171), .A2(n15170), .ZN(n15172) );
  XNOR2_X1 U19785 ( .A(n16449), .B(n1247), .ZN(n15173) );
  XNOR2_X1 U19786 ( .A(n16203), .B(n15173), .ZN(n15214) );
  NAND2_X1 U19787 ( .A1(n28462), .A2(n15180), .ZN(n15178) );
  MUX2_X1 U19788 ( .A(n15178), .B(n15177), .S(n5635), .Z(n15179) );
  MUX2_X1 U19789 ( .A(n15184), .B(n15183), .S(n15182), .Z(n15191) );
  NOR2_X1 U19790 ( .A1(n15186), .A2(n15185), .ZN(n15188) );
  OAI21_X1 U19791 ( .B1(n15188), .B2(n15187), .A(n15190), .ZN(n15189) );
  XNOR2_X1 U19793 ( .A(n15850), .B(n16407), .ZN(n16554) );
  INV_X1 U19794 ( .A(n15192), .ZN(n15198) );
  INV_X1 U19795 ( .A(n15193), .ZN(n15197) );
  NAND2_X1 U19796 ( .A1(n15195), .A2(n15194), .ZN(n15196) );
  OAI211_X1 U19797 ( .C1(n15199), .C2(n15198), .A(n15197), .B(n15196), .ZN(
        n15200) );
  NAND2_X1 U19798 ( .A1(n15201), .A2(n15200), .ZN(n15205) );
  NAND2_X1 U19799 ( .A1(n15202), .A2(n15208), .ZN(n15203) );
  OAI211_X1 U19801 ( .C1(n15209), .C2(n15208), .A(n15207), .B(n15206), .ZN(
        n15210) );
  INV_X1 U19802 ( .A(n16404), .ZN(n15212) );
  XNOR2_X1 U19803 ( .A(n16554), .B(n15745), .ZN(n15213) );
  XNOR2_X1 U19804 ( .A(n15213), .B(n15214), .ZN(n17012) );
  MUX2_X1 U19806 ( .A(n15216), .B(n15215), .S(n15217), .Z(n15221) );
  INV_X1 U19807 ( .A(n15217), .ZN(n15297) );
  NAND2_X1 U19808 ( .A1(n15291), .A2(n14517), .ZN(n15218) );
  AND2_X1 U19809 ( .A1(n15219), .A2(n15218), .ZN(n15220) );
  XNOR2_X1 U19810 ( .A(n16563), .B(n15642), .ZN(n16058) );
  NOR2_X1 U19811 ( .A1(n15222), .A2(n15224), .ZN(n15232) );
  OAI21_X1 U19813 ( .B1(n15229), .B2(n15228), .A(n15227), .ZN(n15230) );
  NOR2_X1 U19814 ( .A1(n15234), .A2(n15233), .ZN(n15237) );
  AND2_X1 U19815 ( .A1(n15334), .A2(n15333), .ZN(n15236) );
  AND2_X1 U19816 ( .A1(n15238), .A2(n15239), .ZN(n15335) );
  INV_X1 U19817 ( .A(n16105), .ZN(n15241) );
  XNOR2_X1 U19818 ( .A(n15241), .B(n16271), .ZN(n16218) );
  INV_X1 U19819 ( .A(n16218), .ZN(n15242) );
  XNOR2_X1 U19820 ( .A(n16058), .B(n15242), .ZN(n15258) );
  XNOR2_X1 U19821 ( .A(n15788), .B(n3321), .ZN(n15256) );
  NAND2_X1 U19822 ( .A1(n15355), .A2(n14752), .ZN(n15244) );
  AOI21_X1 U19823 ( .B1(n15247), .B2(n15246), .A(n15252), .ZN(n15255) );
  XNOR2_X1 U19824 ( .A(n15727), .B(n16360), .ZN(n16566) );
  INV_X1 U19825 ( .A(n16566), .ZN(n16147) );
  NOR2_X1 U19827 ( .A1(n15260), .A2(n15259), .ZN(n15263) );
  XNOR2_X1 U19828 ( .A(n16388), .B(n16586), .ZN(n16031) );
  XNOR2_X1 U19829 ( .A(n16084), .B(n16242), .ZN(n15834) );
  XNOR2_X1 U19830 ( .A(n16031), .B(n15834), .ZN(n15281) );
  NAND2_X1 U19831 ( .A1(n15312), .A2(n15311), .ZN(n15955) );
  NAND2_X1 U19832 ( .A1(n15956), .A2(n15955), .ZN(n15273) );
  OR2_X1 U19833 ( .A1(n15319), .A2(n15272), .ZN(n15954) );
  OR3_X1 U19834 ( .A1(n15276), .A2(n15275), .A3(n15274), .ZN(n15278) );
  XNOR2_X1 U19836 ( .A(n16387), .B(n15545), .ZN(n16588) );
  NAND2_X1 U19837 ( .A1(n17013), .A2(n16788), .ZN(n15331) );
  OAI21_X1 U19838 ( .B1(n15293), .B2(n15292), .A(n15291), .ZN(n15295) );
  NAND2_X1 U19839 ( .A1(n15295), .A2(n15294), .ZN(n15296) );
  INV_X1 U19841 ( .A(n16580), .ZN(n15299) );
  XNOR2_X1 U19842 ( .A(n15299), .B(n16575), .ZN(n16123) );
  OAI21_X1 U19843 ( .B1(n15302), .B2(n15301), .A(n15300), .ZN(n15305) );
  AOI22_X2 U19844 ( .A1(n15305), .A2(n548), .B1(n15304), .B2(n15303), .ZN(
        n16414) );
  XNOR2_X1 U19845 ( .A(n16414), .B(n16579), .ZN(n15762) );
  XNOR2_X1 U19846 ( .A(n16123), .B(n15762), .ZN(n15330) );
  NAND2_X1 U19847 ( .A1(n15307), .A2(n15306), .ZN(n15318) );
  OAI21_X1 U19848 ( .B1(n15309), .B2(n15308), .A(n15315), .ZN(n15314) );
  OAI21_X1 U19849 ( .B1(n15312), .B2(n15311), .A(n15310), .ZN(n15313) );
  NAND2_X1 U19850 ( .A1(n15314), .A2(n15313), .ZN(n15317) );
  OAI21_X1 U19851 ( .B1(n15322), .B2(n15445), .A(n15321), .ZN(n15324) );
  NAND2_X1 U19852 ( .A1(n15324), .A2(n546), .ZN(n15325) );
  XNOR2_X1 U19853 ( .A(n16625), .B(n16255), .ZN(n16223) );
  XNOR2_X1 U19854 ( .A(n16456), .B(n3029), .ZN(n15328) );
  XNOR2_X1 U19855 ( .A(n16223), .B(n15328), .ZN(n15329) );
  MUX2_X2 U19857 ( .A(n15332), .B(n15331), .S(n29152), .Z(n18011) );
  MUX2_X1 U19858 ( .A(n18476), .B(n18475), .S(n18011), .Z(n15523) );
  NOR2_X1 U19859 ( .A1(n15334), .A2(n15333), .ZN(n15336) );
  XNOR2_X1 U19860 ( .A(n16170), .B(n16366), .ZN(n16484) );
  AOI21_X1 U19861 ( .B1(n550), .B2(n15342), .A(n15343), .ZN(n15354) );
  AND2_X1 U19862 ( .A1(n15345), .A2(n15344), .ZN(n15347) );
  NAND4_X1 U19863 ( .A1(n15349), .A2(n15348), .A3(n15347), .A4(n15346), .ZN(
        n15350) );
  OAI21_X1 U19864 ( .B1(n15351), .B2(n425), .A(n15350), .ZN(n15352) );
  AOI21_X1 U19865 ( .B1(n15361), .B2(n15360), .A(n15359), .ZN(n15362) );
  XNOR2_X1 U19867 ( .A(n16279), .B(n16230), .ZN(n15994) );
  XNOR2_X1 U19868 ( .A(n16484), .B(n15994), .ZN(n15368) );
  XNOR2_X1 U19869 ( .A(n29084), .B(n3508), .ZN(n15365) );
  XNOR2_X1 U19870 ( .A(n15366), .B(n15365), .ZN(n15367) );
  NAND2_X1 U19872 ( .A1(n15373), .A2(n426), .ZN(n15375) );
  NAND2_X1 U19873 ( .A1(n15375), .A2(n15374), .ZN(n15377) );
  NAND2_X1 U19874 ( .A1(n15381), .A2(n15380), .ZN(n15386) );
  NAND2_X1 U19875 ( .A1(n15386), .A2(n15385), .ZN(n16373) );
  XNOR2_X1 U19876 ( .A(n16081), .B(n16373), .ZN(n15997) );
  XNOR2_X1 U19877 ( .A(n16082), .B(n15997), .ZN(n15397) );
  XNOR2_X1 U19878 ( .A(n15949), .B(n2544), .ZN(n15396) );
  OAI22_X1 U19879 ( .A1(n15389), .A2(n15388), .B1(n15387), .B2(n15390), .ZN(
        n15393) );
  NAND3_X1 U19880 ( .A1(n15391), .A2(n15394), .A3(n15390), .ZN(n15392) );
  XNOR2_X1 U19881 ( .A(n16589), .B(n16377), .ZN(n16468) );
  NAND2_X1 U19882 ( .A1(n17298), .A2(n29072), .ZN(n16831) );
  NAND2_X1 U19883 ( .A1(n15402), .A2(n15400), .ZN(n15403) );
  MUX2_X1 U19884 ( .A(n15403), .B(n15402), .S(n15401), .Z(n15405) );
  OAI21_X1 U19885 ( .B1(n3362), .B2(n15407), .A(n15406), .ZN(n15413) );
  NAND2_X1 U19886 ( .A1(n15410), .A2(n15409), .ZN(n15411) );
  NAND3_X1 U19887 ( .A1(n15413), .A2(n15412), .A3(n15411), .ZN(n15414) );
  XNOR2_X1 U19889 ( .A(n15914), .B(n16649), .ZN(n15789) );
  NAND3_X1 U19890 ( .A1(n15420), .A2(n15423), .A3(n15417), .ZN(n15418) );
  OAI211_X1 U19891 ( .C1(n15423), .C2(n15422), .A(n15421), .B(n14575), .ZN(
        n15424) );
  XNOR2_X1 U19892 ( .A(n16062), .B(n16569), .ZN(n16461) );
  INV_X1 U19893 ( .A(n16461), .ZN(n15425) );
  XNOR2_X1 U19894 ( .A(n15425), .B(n15789), .ZN(n15429) );
  XNOR2_X1 U19895 ( .A(n16211), .B(n2527), .ZN(n15427) );
  XNOR2_X1 U19896 ( .A(n15426), .B(n15427), .ZN(n15428) );
  NAND2_X1 U19898 ( .A1(n16831), .A2(n17411), .ZN(n15522) );
  NAND2_X1 U19899 ( .A1(n15444), .A2(n15435), .ZN(n15443) );
  NOR2_X1 U19900 ( .A1(n15438), .A2(n15437), .ZN(n15441) );
  NOR2_X1 U19901 ( .A1(n15437), .A2(n15436), .ZN(n15439) );
  AOI22_X1 U19902 ( .A1(n15441), .A2(n15440), .B1(n15439), .B2(n15438), .ZN(
        n15442) );
  XNOR2_X1 U19903 ( .A(n16071), .B(n16303), .ZN(n15769) );
  MUX2_X1 U19904 ( .A(n15446), .B(n15445), .S(n15447), .Z(n15450) );
  XNOR2_X1 U19905 ( .A(n16557), .B(n16339), .ZN(n16450) );
  INV_X1 U19906 ( .A(n16450), .ZN(n15451) );
  XNOR2_X1 U19907 ( .A(n15769), .B(n15451), .ZN(n15455) );
  XNOR2_X1 U19908 ( .A(n16262), .B(n3317), .ZN(n15453) );
  XNOR2_X1 U19909 ( .A(n15852), .B(n15453), .ZN(n15454) );
  XNOR2_X1 U19910 ( .A(n16252), .B(n29319), .ZN(n15470) );
  INV_X1 U19914 ( .A(n16453), .ZN(n15469) );
  XNOR2_X1 U19915 ( .A(n15469), .B(n15470), .ZN(n15483) );
  AOI21_X1 U19916 ( .B1(n15473), .B2(n15472), .A(n15471), .ZN(n15479) );
  NAND2_X1 U19917 ( .A1(n15475), .A2(n15474), .ZN(n15477) );
  AOI21_X1 U19918 ( .B1(n15477), .B2(n15476), .A(n1848), .ZN(n15478) );
  XNOR2_X1 U19919 ( .A(n16319), .B(n15977), .ZN(n15481) );
  XNOR2_X1 U19920 ( .A(n16257), .B(n2511), .ZN(n15480) );
  XNOR2_X1 U19921 ( .A(n15481), .B(n15480), .ZN(n15482) );
  XNOR2_X2 U19922 ( .A(n15483), .B(n15482), .ZN(n17413) );
  NAND2_X1 U19923 ( .A1(n17411), .A2(n29072), .ZN(n15484) );
  NAND2_X1 U19924 ( .A1(n15486), .A2(n15485), .ZN(n15488) );
  NAND2_X1 U19925 ( .A1(n15491), .A2(n15489), .ZN(n15487) );
  NAND3_X1 U19926 ( .A1(n15491), .A2(n3748), .A3(n15489), .ZN(n15492) );
  XNOR2_X1 U19928 ( .A(n16309), .B(n2981), .ZN(n15496) );
  XNOR2_X1 U19929 ( .A(n15496), .B(n16619), .ZN(n15508) );
  NAND2_X1 U19930 ( .A1(n15497), .A2(n15500), .ZN(n15507) );
  NAND3_X1 U19931 ( .A1(n15503), .A2(n15499), .A3(n15498), .ZN(n15505) );
  NAND2_X1 U19932 ( .A1(n15500), .A2(n15502), .ZN(n15501) );
  OAI211_X1 U19933 ( .C1(n15503), .C2(n15502), .A(n15501), .B(n14923), .ZN(
        n15504) );
  XNOR2_X1 U19934 ( .A(n16346), .B(n16607), .ZN(n16481) );
  INV_X1 U19935 ( .A(n16481), .ZN(n15648) );
  XNOR2_X1 U19936 ( .A(n15648), .B(n15508), .ZN(n15521) );
  XNOR2_X1 U19937 ( .A(n16312), .B(n16247), .ZN(n15520) );
  INV_X1 U19938 ( .A(n15509), .ZN(n15519) );
  OAI21_X1 U19939 ( .B1(n5049), .B2(n15511), .A(n15510), .ZN(n15518) );
  NAND2_X1 U19940 ( .A1(n15519), .A2(n15515), .ZN(n15516) );
  XNOR2_X1 U19941 ( .A(n15928), .B(n15520), .ZN(n16098) );
  XNOR2_X1 U19943 ( .A(n16229), .B(n16634), .ZN(n16503) );
  XNOR2_X1 U19944 ( .A(n29084), .B(n15992), .ZN(n16190) );
  INV_X1 U19945 ( .A(n16190), .ZN(n15525) );
  XNOR2_X1 U19946 ( .A(n15525), .B(n16503), .ZN(n15528) );
  XNOR2_X1 U19947 ( .A(n15865), .B(n16284), .ZN(n16369) );
  XNOR2_X1 U19948 ( .A(n16398), .B(n2274), .ZN(n15526) );
  XNOR2_X1 U19949 ( .A(n16369), .B(n15526), .ZN(n15527) );
  XNOR2_X1 U19950 ( .A(n15528), .B(n15527), .ZN(n15551) );
  XNOR2_X1 U19951 ( .A(n16619), .B(n16434), .ZN(n15530) );
  XNOR2_X1 U19952 ( .A(n16310), .B(n26214), .ZN(n15529) );
  XNOR2_X1 U19953 ( .A(n15530), .B(n15529), .ZN(n15534) );
  XNOR2_X1 U19954 ( .A(n16051), .B(n16527), .ZN(n15532) );
  XNOR2_X1 U19955 ( .A(n16017), .B(n3661), .ZN(n15531) );
  XNOR2_X1 U19956 ( .A(n15532), .B(n15531), .ZN(n15533) );
  XNOR2_X1 U19957 ( .A(n15533), .B(n15534), .ZN(n17349) );
  XNOR2_X1 U19958 ( .A(n16264), .B(n15535), .ZN(n16517) );
  INV_X1 U19959 ( .A(n16517), .ZN(n15536) );
  INV_X1 U19960 ( .A(n16305), .ZN(n15537) );
  XNOR2_X1 U19961 ( .A(n15537), .B(n15850), .ZN(n16340) );
  XNOR2_X1 U19962 ( .A(n16404), .B(n3787), .ZN(n15538) );
  XNOR2_X1 U19963 ( .A(n16340), .B(n15538), .ZN(n15539) );
  XNOR2_X1 U19964 ( .A(n16360), .B(n16211), .ZN(n15877) );
  XNOR2_X1 U19965 ( .A(n16271), .B(n16146), .ZN(n16532) );
  XNOR2_X1 U19966 ( .A(n16532), .B(n15877), .ZN(n15544) );
  XNOR2_X1 U19967 ( .A(n28579), .B(n15642), .ZN(n15542) );
  XNOR2_X1 U19968 ( .A(n16216), .B(n22072), .ZN(n15541) );
  XNOR2_X1 U19969 ( .A(n15542), .B(n15541), .ZN(n15543) );
  XNOR2_X1 U19970 ( .A(n15544), .B(n15543), .ZN(n17346) );
  INV_X1 U19971 ( .A(n17346), .ZN(n17029) );
  XNOR2_X1 U19972 ( .A(n16510), .B(n2402), .ZN(n15546) );
  XNOR2_X1 U19973 ( .A(n16376), .B(n15546), .ZN(n15550) );
  XNOR2_X1 U19974 ( .A(n15949), .B(n15760), .ZN(n16208) );
  INV_X1 U19975 ( .A(n16208), .ZN(n15548) );
  XNOR2_X1 U19976 ( .A(n16388), .B(n16242), .ZN(n15547) );
  XNOR2_X1 U19977 ( .A(n15548), .B(n15547), .ZN(n15549) );
  INV_X1 U19978 ( .A(n15551), .ZN(n17192) );
  MUX2_X1 U19979 ( .A(n17029), .B(n17347), .S(n17192), .Z(n15557) );
  INV_X1 U19980 ( .A(n16318), .ZN(n15552) );
  XNOR2_X1 U19981 ( .A(n16414), .B(n15552), .ZN(n15553) );
  XNOR2_X1 U19982 ( .A(n16224), .B(n15553), .ZN(n15556) );
  XNOR2_X1 U19984 ( .A(n29151), .B(n2984), .ZN(n15554) );
  XNOR2_X1 U19985 ( .A(n16499), .B(n15554), .ZN(n15555) );
  XNOR2_X1 U19986 ( .A(n16568), .B(n15790), .ZN(n16214) );
  XNOR2_X1 U19987 ( .A(n15944), .B(n16214), .ZN(n15560) );
  XNOR2_X1 U19988 ( .A(n16185), .B(n16295), .ZN(n16102) );
  XNOR2_X1 U19989 ( .A(n16102), .B(n15558), .ZN(n15559) );
  XNOR2_X1 U19990 ( .A(n15561), .B(n15965), .ZN(n15564) );
  XNOR2_X1 U19991 ( .A(n16090), .B(n15668), .ZN(n15563) );
  XNOR2_X1 U19992 ( .A(n29571), .B(n2411), .ZN(n15562) );
  NOR2_X1 U19993 ( .A1(n17338), .A2(n17340), .ZN(n15582) );
  XNOR2_X1 U19994 ( .A(n16444), .B(n15565), .ZN(n16300) );
  XNOR2_X1 U19995 ( .A(n15900), .B(n16519), .ZN(n15566) );
  XNOR2_X1 U19996 ( .A(n16300), .B(n15566), .ZN(n15570) );
  XNOR2_X1 U19997 ( .A(n15772), .B(n16070), .ZN(n15567) );
  XNOR2_X1 U19998 ( .A(n15568), .B(n15567), .ZN(n15569) );
  XNOR2_X1 U19999 ( .A(n16165), .B(n16312), .ZN(n15572) );
  XNOR2_X1 U20000 ( .A(n15927), .B(n3191), .ZN(n15571) );
  XNOR2_X1 U20001 ( .A(n15572), .B(n15571), .ZN(n15574) );
  XNOR2_X1 U20002 ( .A(n15780), .B(n16605), .ZN(n16197) );
  XNOR2_X1 U20003 ( .A(n15973), .B(n16197), .ZN(n15573) );
  INV_X1 U20004 ( .A(n17155), .ZN(n17200) );
  XNOR2_X1 U20005 ( .A(n16322), .B(n16077), .ZN(n15858) );
  XNOR2_X1 U20006 ( .A(n16578), .B(n15654), .ZN(n16221) );
  XNOR2_X1 U20007 ( .A(n15858), .B(n16221), .ZN(n15580) );
  XNOR2_X1 U20008 ( .A(n6454), .B(n16498), .ZN(n15578) );
  XNOR2_X1 U20009 ( .A(n15578), .B(n15577), .ZN(n15579) );
  INV_X1 U20010 ( .A(n17204), .ZN(n17339) );
  XNOR2_X1 U20012 ( .A(n16085), .B(n16329), .ZN(n15872) );
  XNOR2_X1 U20013 ( .A(n15999), .B(n16585), .ZN(n16207) );
  XNOR2_X1 U20014 ( .A(n15872), .B(n16207), .ZN(n15587) );
  XNOR2_X1 U20015 ( .A(n15583), .B(n15909), .ZN(n15585) );
  XNOR2_X1 U20016 ( .A(n16241), .B(n1119), .ZN(n15584) );
  XNOR2_X1 U20017 ( .A(n15585), .B(n15584), .ZN(n15586) );
  MUX2_X1 U20018 ( .A(n28564), .B(n17335), .S(n17338), .Z(n15588) );
  NOR2_X1 U20019 ( .A1(n17336), .A2(n15588), .ZN(n15589) );
  XNOR2_X1 U20020 ( .A(n16449), .B(n16023), .ZN(n15770) );
  XNOR2_X1 U20021 ( .A(n16557), .B(n16519), .ZN(n15591) );
  XNOR2_X1 U20022 ( .A(n15770), .B(n15591), .ZN(n15594) );
  XNOR2_X1 U20023 ( .A(n16303), .B(n3607), .ZN(n15592) );
  XNOR2_X1 U20024 ( .A(n15594), .B(n15593), .ZN(n17389) );
  XNOR2_X1 U20025 ( .A(n16456), .B(n16038), .ZN(n15782) );
  XNOR2_X1 U20026 ( .A(n16319), .B(n16498), .ZN(n15595) );
  XNOR2_X1 U20027 ( .A(n15782), .B(n15595), .ZN(n15599) );
  XNOR2_X1 U20028 ( .A(n16257), .B(n26680), .ZN(n15596) );
  XNOR2_X1 U20029 ( .A(n15597), .B(n15596), .ZN(n15598) );
  XNOR2_X1 U20030 ( .A(n15598), .B(n15599), .ZN(n16700) );
  NAND2_X1 U20031 ( .A1(n17389), .A2(n29045), .ZN(n17162) );
  XNOR2_X1 U20032 ( .A(n15802), .B(n16467), .ZN(n16032) );
  INV_X1 U20033 ( .A(n16238), .ZN(n15711) );
  XNOR2_X1 U20034 ( .A(n15801), .B(n15711), .ZN(n15600) );
  XNOR2_X1 U20035 ( .A(n15600), .B(n16032), .ZN(n15604) );
  XNOR2_X1 U20036 ( .A(n16373), .B(n16589), .ZN(n15602) );
  XNOR2_X1 U20037 ( .A(n16241), .B(n891), .ZN(n15601) );
  XNOR2_X1 U20038 ( .A(n15602), .B(n15601), .ZN(n15603) );
  XNOR2_X1 U20039 ( .A(n15788), .B(n16272), .ZN(n15606) );
  XNOR2_X1 U20040 ( .A(n16569), .B(n16534), .ZN(n15605) );
  XNOR2_X1 U20041 ( .A(n15605), .B(n15606), .ZN(n15610) );
  INV_X1 U20042 ( .A(n2476), .ZN(n24356) );
  XNOR2_X1 U20043 ( .A(n321), .B(n24356), .ZN(n15607) );
  XNOR2_X1 U20044 ( .A(n15608), .B(n15607), .ZN(n15609) );
  NAND2_X1 U20045 ( .A1(n17386), .A2(n17385), .ZN(n15611) );
  NAND2_X1 U20046 ( .A1(n17162), .A2(n15611), .ZN(n15616) );
  XNOR2_X1 U20047 ( .A(n16247), .B(n2404), .ZN(n15612) );
  XNOR2_X1 U20048 ( .A(n16309), .B(n16607), .ZN(n15613) );
  XNOR2_X1 U20049 ( .A(n15777), .B(n15613), .ZN(n15614) );
  XNOR2_X1 U20050 ( .A(n16483), .B(n16233), .ZN(n15698) );
  OAI21_X1 U20052 ( .B1(n17382), .B2(n28497), .A(n17385), .ZN(n15615) );
  OAI21_X1 U20054 ( .B1(n18493), .B2(n18292), .A(n28633), .ZN(n15737) );
  XNOR2_X1 U20057 ( .A(n16280), .B(n16636), .ZN(n15620) );
  XNOR2_X1 U20058 ( .A(n15620), .B(n15619), .ZN(n15624) );
  XNOR2_X1 U20059 ( .A(n16596), .B(n16230), .ZN(n15622) );
  XNOR2_X1 U20060 ( .A(n16398), .B(n5633), .ZN(n15621) );
  XNOR2_X1 U20061 ( .A(n15622), .B(n15621), .ZN(n15623) );
  XNOR2_X1 U20062 ( .A(n15624), .B(n15623), .ZN(n17355) );
  XNOR2_X1 U20064 ( .A(n16321), .B(n16416), .ZN(n15859) );
  XNOR2_X1 U20065 ( .A(n15625), .B(n15859), .ZN(n15628) );
  XNOR2_X1 U20066 ( .A(n16256), .B(n16625), .ZN(n15822) );
  XNOR2_X1 U20067 ( .A(n16578), .B(n27231), .ZN(n15626) );
  XNOR2_X1 U20068 ( .A(n15822), .B(n15626), .ZN(n15627) );
  XNOR2_X1 U20069 ( .A(n16081), .B(n16641), .ZN(n16240) );
  XNOR2_X1 U20070 ( .A(n28585), .B(n16471), .ZN(n15629) );
  XNOR2_X1 U20071 ( .A(n16240), .B(n15629), .ZN(n15633) );
  XNOR2_X1 U20072 ( .A(n15631), .B(n15630), .ZN(n15632) );
  XNOR2_X1 U20073 ( .A(n15633), .B(n15632), .ZN(n17357) );
  MUX2_X1 U20074 ( .A(n17355), .B(n17359), .S(n17357), .Z(n15647) );
  XNOR2_X1 U20075 ( .A(n16404), .B(n3662), .ZN(n15634) );
  INV_X1 U20076 ( .A(n15849), .ZN(n16408) );
  XNOR2_X1 U20077 ( .A(n16408), .B(n16556), .ZN(n15636) );
  XNOR2_X1 U20078 ( .A(n15636), .B(n16654), .ZN(n15637) );
  NOR2_X1 U20080 ( .A1(n17354), .A2(n17359), .ZN(n17198) );
  XNOR2_X1 U20081 ( .A(n16605), .B(n16434), .ZN(n15639) );
  XNOR2_X1 U20082 ( .A(n15928), .B(n16618), .ZN(n16246) );
  INV_X1 U20083 ( .A(n16620), .ZN(n16095) );
  XNOR2_X1 U20084 ( .A(n16436), .B(n16095), .ZN(n15975) );
  INV_X1 U20085 ( .A(n17356), .ZN(n17196) );
  NAND2_X1 U20086 ( .A1(n17198), .A2(n17196), .ZN(n15646) );
  XNOR2_X1 U20087 ( .A(n15914), .B(n15817), .ZN(n16269) );
  INV_X1 U20088 ( .A(n16269), .ZN(n15641) );
  XNOR2_X1 U20089 ( .A(n16291), .B(n16568), .ZN(n15640) );
  XNOR2_X1 U20090 ( .A(n16105), .B(n3554), .ZN(n15643) );
  XNOR2_X1 U20091 ( .A(n15644), .B(n15643), .ZN(n15645) );
  INV_X1 U20092 ( .A(n17030), .ZN(n16953) );
  INV_X1 U20093 ( .A(n18489), .ZN(n17674) );
  NOR2_X1 U20094 ( .A1(n18487), .A2(n17674), .ZN(n15736) );
  XNOR2_X1 U20095 ( .A(n15649), .B(n15648), .ZN(n15653) );
  XNOR2_X1 U20096 ( .A(n29525), .B(n15927), .ZN(n15651) );
  XNOR2_X1 U20097 ( .A(n16247), .B(n26825), .ZN(n15650) );
  XNOR2_X1 U20098 ( .A(n15651), .B(n15650), .ZN(n15652) );
  XNOR2_X1 U20099 ( .A(n28557), .B(n6449), .ZN(n15656) );
  XNOR2_X1 U20100 ( .A(n16574), .B(n15654), .ZN(n15655) );
  XNOR2_X1 U20101 ( .A(n15656), .B(n15655), .ZN(n15660) );
  INV_X1 U20102 ( .A(n2577), .ZN(n25902) );
  XNOR2_X1 U20103 ( .A(n16257), .B(n25902), .ZN(n15657) );
  XNOR2_X1 U20104 ( .A(n15658), .B(n15657), .ZN(n15659) );
  XNOR2_X1 U20105 ( .A(n16426), .B(n16272), .ZN(n16107) );
  INV_X1 U20106 ( .A(n16107), .ZN(n15661) );
  INV_X1 U20107 ( .A(n16062), .ZN(n16143) );
  XNOR2_X1 U20108 ( .A(n16143), .B(n16563), .ZN(n16359) );
  XNOR2_X1 U20109 ( .A(n16359), .B(n15661), .ZN(n15665) );
  XNOR2_X1 U20110 ( .A(n16294), .B(n15790), .ZN(n15663) );
  XNOR2_X1 U20111 ( .A(n16569), .B(n1927), .ZN(n15662) );
  XNOR2_X1 U20112 ( .A(n15663), .B(n15662), .ZN(n15664) );
  XNOR2_X1 U20113 ( .A(n15665), .B(n15664), .ZN(n16762) );
  INV_X1 U20115 ( .A(n16484), .ZN(n15667) );
  XNOR2_X1 U20116 ( .A(n16233), .B(n16365), .ZN(n15666) );
  XNOR2_X1 U20117 ( .A(n15667), .B(n15666), .ZN(n15672) );
  XNOR2_X1 U20118 ( .A(n16399), .B(n15668), .ZN(n15670) );
  XNOR2_X1 U20119 ( .A(n15989), .B(n3256), .ZN(n15669) );
  XNOR2_X1 U20120 ( .A(n15670), .B(n15669), .ZN(n15671) );
  INV_X1 U20121 ( .A(n15772), .ZN(n16199) );
  XNOR2_X1 U20122 ( .A(n15900), .B(n15673), .ZN(n15677) );
  XNOR2_X1 U20123 ( .A(n16262), .B(n2961), .ZN(n15674) );
  XNOR2_X1 U20124 ( .A(n15674), .B(n16405), .ZN(n15675) );
  XNOR2_X1 U20125 ( .A(n15675), .B(n16450), .ZN(n15676) );
  XNOR2_X1 U20126 ( .A(n15676), .B(n15677), .ZN(n16943) );
  NAND2_X1 U20128 ( .A1(n17549), .A2(n16944), .ZN(n16947) );
  INV_X1 U20129 ( .A(n16947), .ZN(n15686) );
  XNOR2_X1 U20130 ( .A(n16238), .B(n28597), .ZN(n15680) );
  INV_X1 U20131 ( .A(n15999), .ZN(n15678) );
  XNOR2_X1 U20132 ( .A(n15678), .B(n16586), .ZN(n15679) );
  XNOR2_X1 U20133 ( .A(n15679), .B(n15680), .ZN(n15684) );
  XNOR2_X1 U20134 ( .A(n16589), .B(n3232), .ZN(n15681) );
  XNOR2_X1 U20135 ( .A(n15682), .B(n15681), .ZN(n15683) );
  INV_X1 U20136 ( .A(n17548), .ZN(n17239) );
  OAI21_X1 U20137 ( .B1(n15686), .B2(n15685), .A(n17552), .ZN(n15687) );
  INV_X1 U20138 ( .A(n18490), .ZN(n18015) );
  XNOR2_X1 U20141 ( .A(n16395), .B(n1849), .ZN(n15696) );
  XNOR2_X1 U20142 ( .A(n16043), .B(n16393), .ZN(n16504) );
  XNOR2_X1 U20143 ( .A(n15696), .B(n16504), .ZN(n15700) );
  XNOR2_X1 U20144 ( .A(n16284), .B(n3462), .ZN(n15697) );
  XNOR2_X1 U20145 ( .A(n15698), .B(n15697), .ZN(n15699) );
  INV_X1 U20147 ( .A(n17368), .ZN(n17366) );
  XNOR2_X1 U20148 ( .A(n16495), .B(n15701), .ZN(n16415) );
  XNOR2_X1 U20149 ( .A(n16160), .B(n16494), .ZN(n16577) );
  XNOR2_X1 U20150 ( .A(n16577), .B(n16415), .ZN(n15705) );
  XNOR2_X1 U20151 ( .A(n16257), .B(n3164), .ZN(n15702) );
  XNOR2_X1 U20152 ( .A(n15703), .B(n15702), .ZN(n15704) );
  XNOR2_X1 U20153 ( .A(n15705), .B(n15704), .ZN(n17361) );
  XNOR2_X1 U20154 ( .A(n15706), .B(n15971), .ZN(n16433) );
  INV_X1 U20155 ( .A(n16433), .ZN(n15707) );
  XNOR2_X1 U20156 ( .A(n15707), .B(n259), .ZN(n15710) );
  XNOR2_X1 U20157 ( .A(n16606), .B(n16310), .ZN(n16166) );
  XNOR2_X1 U20158 ( .A(n16247), .B(n2389), .ZN(n15708) );
  XNOR2_X1 U20159 ( .A(n16166), .B(n15708), .ZN(n15709) );
  INV_X1 U20160 ( .A(n17365), .ZN(n17369) );
  XNOR2_X1 U20161 ( .A(n15711), .B(n16509), .ZN(n15712) );
  XNOR2_X1 U20162 ( .A(n15712), .B(n16591), .ZN(n15716) );
  XNOR2_X1 U20163 ( .A(n16387), .B(n16467), .ZN(n15714) );
  XNOR2_X1 U20164 ( .A(n16332), .B(n1887), .ZN(n15713) );
  XNOR2_X1 U20165 ( .A(n15714), .B(n15713), .ZN(n15715) );
  XNOR2_X1 U20166 ( .A(n15716), .B(n15715), .ZN(n15731) );
  XNOR2_X1 U20167 ( .A(n16558), .B(n16407), .ZN(n15718) );
  XNOR2_X1 U20168 ( .A(n16024), .B(n16409), .ZN(n16521) );
  XNOR2_X1 U20169 ( .A(n15718), .B(n16521), .ZN(n15722) );
  XNOR2_X1 U20170 ( .A(n16305), .B(n3622), .ZN(n15719) );
  XNOR2_X1 U20171 ( .A(n15720), .B(n15719), .ZN(n15721) );
  XNOR2_X1 U20173 ( .A(n16422), .B(n15723), .ZN(n16533) );
  INV_X1 U20174 ( .A(n16533), .ZN(n15726) );
  XNOR2_X1 U20175 ( .A(n16059), .B(n3081), .ZN(n15724) );
  XNOR2_X1 U20176 ( .A(n15724), .B(n16272), .ZN(n15725) );
  XNOR2_X1 U20177 ( .A(n15725), .B(n15726), .ZN(n15730) );
  XNOR2_X1 U20178 ( .A(n28579), .B(n16427), .ZN(n15728) );
  INV_X1 U20179 ( .A(n16564), .ZN(n16213) );
  XNOR2_X1 U20180 ( .A(n16213), .B(n15728), .ZN(n15729) );
  XNOR2_X1 U20181 ( .A(n15730), .B(n15729), .ZN(n17234) );
  INV_X1 U20182 ( .A(n28632), .ZN(n18486) );
  OAI211_X1 U20183 ( .C1(n18015), .C2(n18489), .A(n15734), .B(n18486), .ZN(
        n15735) );
  XNOR2_X1 U20184 ( .A(n19495), .B(n19103), .ZN(n19650) );
  XNOR2_X1 U20185 ( .A(n15668), .B(n2541), .ZN(n15740) );
  XNOR2_X1 U20186 ( .A(n15738), .B(n15992), .ZN(n15739) );
  XNOR2_X1 U20187 ( .A(n15740), .B(n15739), .ZN(n15743) );
  XNOR2_X1 U20188 ( .A(n16397), .B(n15741), .ZN(n15742) );
  XNOR2_X1 U20189 ( .A(n16443), .B(n1919), .ZN(n15744) );
  XNOR2_X1 U20190 ( .A(n15744), .B(n15982), .ZN(n15747) );
  INV_X1 U20191 ( .A(n15745), .ZN(n15746) );
  XNOR2_X1 U20192 ( .A(n15747), .B(n15746), .ZN(n15749) );
  XNOR2_X1 U20193 ( .A(n16406), .B(n15900), .ZN(n15748) );
  XNOR2_X1 U20194 ( .A(n16527), .B(n16606), .ZN(n16432) );
  XNOR2_X1 U20195 ( .A(n16432), .B(n16050), .ZN(n15753) );
  XNOR2_X1 U20196 ( .A(n16017), .B(n16476), .ZN(n15751) );
  XNOR2_X1 U20197 ( .A(n15927), .B(n25992), .ZN(n15750) );
  XNOR2_X1 U20198 ( .A(n15751), .B(n15750), .ZN(n15752) );
  XNOR2_X1 U20199 ( .A(n15753), .B(n15752), .ZN(n16918) );
  NOR2_X1 U20200 ( .A1(n17317), .A2(n16918), .ZN(n15754) );
  AOI21_X1 U20201 ( .B1(n17316), .B2(n17317), .A(n15754), .ZN(n15768) );
  INV_X1 U20202 ( .A(n16058), .ZN(n15755) );
  XNOR2_X1 U20203 ( .A(n15755), .B(n16424), .ZN(n15759) );
  XNOR2_X1 U20204 ( .A(n16294), .B(n16216), .ZN(n15757) );
  XNOR2_X1 U20205 ( .A(n16059), .B(n3722), .ZN(n15756) );
  XNOR2_X1 U20206 ( .A(n15757), .B(n15756), .ZN(n15758) );
  XNOR2_X1 U20207 ( .A(n16467), .B(n3386), .ZN(n15761) );
  INV_X1 U20208 ( .A(n15760), .ZN(n16000) );
  XNOR2_X1 U20210 ( .A(n16418), .B(n15762), .ZN(n15766) );
  XNOR2_X1 U20211 ( .A(n15764), .B(n15763), .ZN(n15765) );
  XNOR2_X1 U20212 ( .A(n15766), .B(n15765), .ZN(n17312) );
  INV_X1 U20213 ( .A(n17312), .ZN(n17560) );
  INV_X1 U20214 ( .A(n15769), .ZN(n15771) );
  XNOR2_X1 U20215 ( .A(n16408), .B(n15772), .ZN(n15774) );
  XNOR2_X1 U20216 ( .A(n16444), .B(n3491), .ZN(n15773) );
  XNOR2_X1 U20217 ( .A(n15774), .B(n15773), .ZN(n15775) );
  XNOR2_X1 U20218 ( .A(n15928), .B(n16052), .ZN(n15778) );
  XNOR2_X1 U20219 ( .A(n16309), .B(n15780), .ZN(n16617) );
  XNOR2_X1 U20220 ( .A(n15781), .B(n16319), .ZN(n16629) );
  INV_X1 U20221 ( .A(n16629), .ZN(n16011) );
  XNOR2_X1 U20222 ( .A(n16011), .B(n15782), .ZN(n15786) );
  XNOR2_X1 U20223 ( .A(n16416), .B(n16252), .ZN(n15784) );
  XNOR2_X1 U20224 ( .A(n16323), .B(n2973), .ZN(n15783) );
  XNOR2_X1 U20225 ( .A(n15784), .B(n15783), .ZN(n15785) );
  INV_X1 U20227 ( .A(n17541), .ZN(n15787) );
  XNOR2_X1 U20228 ( .A(n16296), .B(n15788), .ZN(n16462) );
  XNOR2_X1 U20229 ( .A(n15789), .B(n16462), .ZN(n15794) );
  XNOR2_X1 U20230 ( .A(n16421), .B(n15790), .ZN(n15792) );
  XNOR2_X1 U20231 ( .A(n321), .B(n1133), .ZN(n15791) );
  XNOR2_X1 U20232 ( .A(n15792), .B(n15791), .ZN(n15793) );
  INV_X1 U20233 ( .A(n15994), .ZN(n15795) );
  XNOR2_X1 U20234 ( .A(n15795), .B(n15796), .ZN(n15800) );
  XNOR2_X1 U20235 ( .A(n16400), .B(n16283), .ZN(n15798) );
  XNOR2_X1 U20236 ( .A(n15989), .B(n3035), .ZN(n15797) );
  XNOR2_X1 U20237 ( .A(n15798), .B(n15797), .ZN(n15799) );
  OAI22_X1 U20238 ( .A1(n17542), .A2(n17545), .B1(n17543), .B2(n17540), .ZN(
        n15807) );
  XNOR2_X1 U20239 ( .A(n15801), .B(n16328), .ZN(n16472) );
  XNOR2_X1 U20240 ( .A(n16472), .B(n15997), .ZN(n15806) );
  INV_X1 U20241 ( .A(n28585), .ZN(n16386) );
  XNOR2_X1 U20242 ( .A(n15802), .B(n16386), .ZN(n15804) );
  XNOR2_X1 U20243 ( .A(n15999), .B(n28294), .ZN(n15803) );
  XNOR2_X1 U20244 ( .A(n15804), .B(n15803), .ZN(n15805) );
  XNOR2_X1 U20245 ( .A(n15806), .B(n15805), .ZN(n17539) );
  INV_X1 U20246 ( .A(n17539), .ZN(n17213) );
  NAND2_X1 U20247 ( .A1(n15807), .A2(n17213), .ZN(n15809) );
  NAND2_X1 U20248 ( .A1(n17217), .A2(n17545), .ZN(n15808) );
  INV_X1 U20250 ( .A(n17413), .ZN(n17297) );
  INV_X1 U20251 ( .A(n17414), .ZN(n17300) );
  NAND2_X1 U20252 ( .A1(n15812), .A2(n17300), .ZN(n15816) );
  NAND3_X1 U20253 ( .A1(n17298), .A2(n17297), .A3(n17414), .ZN(n15814) );
  NAND2_X1 U20254 ( .A1(n17298), .A2(n17411), .ZN(n15813) );
  AND2_X1 U20255 ( .A1(n15814), .A2(n15813), .ZN(n15815) );
  NAND2_X1 U20256 ( .A1(n15816), .A2(n15815), .ZN(n17926) );
  INV_X1 U20257 ( .A(n17926), .ZN(n18059) );
  XNOR2_X1 U20258 ( .A(n16360), .B(n15817), .ZN(n15819) );
  XNOR2_X1 U20259 ( .A(n16059), .B(n3276), .ZN(n15818) );
  XNOR2_X1 U20260 ( .A(n15819), .B(n15818), .ZN(n15821) );
  XNOR2_X1 U20262 ( .A(n15822), .B(n29630), .ZN(n15827) );
  XNOR2_X1 U20263 ( .A(n29151), .B(n3654), .ZN(n15824) );
  XNOR2_X1 U20264 ( .A(n15825), .B(n15824), .ZN(n15826) );
  XNOR2_X1 U20265 ( .A(n16203), .B(n16134), .ZN(n15832) );
  XNOR2_X1 U20266 ( .A(n15828), .B(n15850), .ZN(n15830) );
  XNOR2_X1 U20267 ( .A(n16443), .B(n3695), .ZN(n15829) );
  XNOR2_X1 U20268 ( .A(n15830), .B(n15829), .ZN(n15831) );
  INV_X1 U20269 ( .A(n16119), .ZN(n15833) );
  XNOR2_X1 U20270 ( .A(n15833), .B(n15834), .ZN(n15838) );
  XNOR2_X1 U20271 ( .A(n16641), .B(n3114), .ZN(n15835) );
  XNOR2_X1 U20272 ( .A(n15836), .B(n15835), .ZN(n15837) );
  XNOR2_X1 U20273 ( .A(n16191), .B(n16116), .ZN(n15842) );
  XNOR2_X1 U20274 ( .A(n16483), .B(n16232), .ZN(n15840) );
  XNOR2_X1 U20275 ( .A(n15865), .B(n3087), .ZN(n15839) );
  XNOR2_X1 U20276 ( .A(n15840), .B(n15839), .ZN(n15841) );
  INV_X1 U20277 ( .A(n17554), .ZN(n16911) );
  XNOR2_X1 U20278 ( .A(n16196), .B(n16138), .ZN(n15846) );
  XNOR2_X1 U20279 ( .A(n16618), .B(n3661), .ZN(n15844) );
  XNOR2_X1 U20280 ( .A(n16476), .B(n900), .ZN(n15843) );
  XNOR2_X1 U20281 ( .A(n15844), .B(n15843), .ZN(n15845) );
  INV_X1 U20282 ( .A(n16908), .ZN(n17221) );
  OAI21_X1 U20283 ( .B1(n18298), .B2(n18059), .A(n29561), .ZN(n15938) );
  XNOR2_X1 U20285 ( .A(n15851), .B(n15850), .ZN(n15853) );
  XNOR2_X1 U20286 ( .A(n16519), .B(n16070), .ZN(n15854) );
  XNOR2_X1 U20287 ( .A(n15855), .B(n15977), .ZN(n15857) );
  XNOR2_X1 U20288 ( .A(n29151), .B(n2350), .ZN(n15856) );
  XNOR2_X1 U20289 ( .A(n15857), .B(n15856), .ZN(n15861) );
  XNOR2_X1 U20290 ( .A(n15859), .B(n15858), .ZN(n15860) );
  XNOR2_X1 U20291 ( .A(n15863), .B(n15862), .ZN(n16237) );
  XNOR2_X1 U20292 ( .A(n15966), .B(n28327), .ZN(n15864) );
  XNOR2_X1 U20293 ( .A(n15864), .B(n16090), .ZN(n15867) );
  XNOR2_X1 U20294 ( .A(n15865), .B(n16400), .ZN(n15866) );
  XNOR2_X1 U20295 ( .A(n15867), .B(n15866), .ZN(n15868) );
  INV_X1 U20296 ( .A(n15949), .ZN(n15870) );
  XNOR2_X1 U20298 ( .A(n15872), .B(n15871), .ZN(n15876) );
  XNOR2_X1 U20299 ( .A(n16241), .B(n2602), .ZN(n15873) );
  XNOR2_X1 U20300 ( .A(n15874), .B(n15873), .ZN(n15875) );
  NAND2_X1 U20301 ( .A1(n1166), .A2(n4118), .ZN(n15884) );
  INV_X1 U20302 ( .A(n15877), .ZN(n15879) );
  XNOR2_X1 U20303 ( .A(n15878), .B(n15879), .ZN(n15883) );
  XNOR2_X1 U20304 ( .A(n16295), .B(n16421), .ZN(n15881) );
  XNOR2_X1 U20305 ( .A(n16534), .B(n3372), .ZN(n15880) );
  XNOR2_X1 U20306 ( .A(n15881), .B(n15880), .ZN(n15882) );
  INV_X1 U20307 ( .A(n29098), .ZN(n17037) );
  XNOR2_X1 U20308 ( .A(n1967), .B(n3661), .ZN(n15886) );
  XNOR2_X1 U20309 ( .A(n16619), .B(n16165), .ZN(n15885) );
  XNOR2_X1 U20310 ( .A(n15886), .B(n15885), .ZN(n15891) );
  XNOR2_X1 U20311 ( .A(n15887), .B(n16312), .ZN(n15889) );
  XNOR2_X1 U20312 ( .A(n16313), .B(n2505), .ZN(n15888) );
  XNOR2_X1 U20313 ( .A(n15889), .B(n15888), .ZN(n15890) );
  XNOR2_X1 U20314 ( .A(n15891), .B(n15890), .ZN(n17566) );
  INV_X1 U20315 ( .A(n17566), .ZN(n17038) );
  XNOR2_X1 U20317 ( .A(n16154), .B(n15893), .ZN(n15902) );
  XNOR2_X1 U20318 ( .A(n15894), .B(n27956), .ZN(n15897) );
  XNOR2_X1 U20319 ( .A(n15895), .B(n27956), .ZN(n15896) );
  XNOR2_X1 U20320 ( .A(n15898), .B(n16407), .ZN(n15899) );
  XNOR2_X1 U20321 ( .A(n15899), .B(n15900), .ZN(n15901) );
  XNOR2_X1 U20322 ( .A(n15902), .B(n15901), .ZN(n17571) );
  XNOR2_X1 U20323 ( .A(n16162), .B(n15903), .ZN(n15907) );
  XNOR2_X1 U20324 ( .A(n16575), .B(n16252), .ZN(n15905) );
  XNOR2_X1 U20325 ( .A(n15905), .B(n15904), .ZN(n15906) );
  XNOR2_X1 U20326 ( .A(n15906), .B(n15907), .ZN(n16904) );
  NAND2_X1 U20327 ( .A1(n17571), .A2(n16904), .ZN(n17404) );
  INV_X1 U20328 ( .A(n16179), .ZN(n15908) );
  XNOR2_X1 U20329 ( .A(n15908), .B(n16375), .ZN(n15913) );
  XNOR2_X1 U20330 ( .A(n16387), .B(n16081), .ZN(n15911) );
  XNOR2_X1 U20331 ( .A(n15909), .B(n3598), .ZN(n15910) );
  XNOR2_X1 U20332 ( .A(n15911), .B(n15910), .ZN(n15912) );
  XNOR2_X1 U20333 ( .A(n15914), .B(n16294), .ZN(n15915) );
  XNOR2_X1 U20334 ( .A(n16183), .B(n15915), .ZN(n15918) );
  XNOR2_X1 U20335 ( .A(n16427), .B(n3643), .ZN(n15916) );
  XNOR2_X1 U20336 ( .A(n16362), .B(n15916), .ZN(n15917) );
  XNOR2_X1 U20337 ( .A(n15917), .B(n15918), .ZN(n17405) );
  NAND2_X1 U20338 ( .A1(n17572), .A2(n17405), .ZN(n17403) );
  XNOR2_X1 U20343 ( .A(n16395), .B(n15668), .ZN(n15920) );
  XNOR2_X1 U20345 ( .A(n16230), .B(n3336), .ZN(n15922) );
  XNOR2_X1 U20346 ( .A(n16367), .B(n15922), .ZN(n15923) );
  XNOR2_X1 U20347 ( .A(n15924), .B(n15923), .ZN(n16822) );
  XNOR2_X1 U20348 ( .A(n16310), .B(n2523), .ZN(n15926) );
  INV_X1 U20349 ( .A(n15971), .ZN(n15925) );
  XNOR2_X1 U20350 ( .A(n15928), .B(n15927), .ZN(n15929) );
  XNOR2_X1 U20351 ( .A(n15929), .B(n15777), .ZN(n15930) );
  INV_X1 U20352 ( .A(n17572), .ZN(n17320) );
  NAND3_X1 U20353 ( .A1(n17707), .A2(n17570), .A3(n17320), .ZN(n15933) );
  NAND3_X1 U20354 ( .A1(n17707), .A2(n16904), .A3(n17320), .ZN(n15932) );
  NOR2_X1 U20355 ( .A1(n18298), .A2(n1861), .ZN(n15935) );
  INV_X1 U20356 ( .A(n18060), .ZN(n17928) );
  NAND2_X1 U20357 ( .A1(n15935), .A2(n17928), .ZN(n15936) );
  XNOR2_X1 U20359 ( .A(n15940), .B(n21865), .ZN(n15941) );
  XNOR2_X1 U20360 ( .A(n16654), .B(n16407), .ZN(n15942) );
  XNOR2_X1 U20361 ( .A(n16105), .B(n16211), .ZN(n16648) );
  INV_X1 U20362 ( .A(n16648), .ZN(n15943) );
  XNOR2_X1 U20363 ( .A(n15943), .B(n15944), .ZN(n15946) );
  INV_X1 U20364 ( .A(n16514), .ZN(n15947) );
  XNOR2_X1 U20365 ( .A(n15947), .B(n15948), .ZN(n15963) );
  XNOR2_X1 U20366 ( .A(n15949), .B(n16084), .ZN(n15961) );
  INV_X1 U20367 ( .A(n15955), .ZN(n15950) );
  NAND2_X1 U20368 ( .A1(n15950), .A2(n3635), .ZN(n15952) );
  INV_X1 U20369 ( .A(n15954), .ZN(n15951) );
  MUX2_X1 U20370 ( .A(n15952), .B(n3635), .S(n15951), .Z(n15959) );
  INV_X1 U20371 ( .A(n15956), .ZN(n15953) );
  NAND3_X1 U20372 ( .A1(n15954), .A2(n15953), .A3(n3635), .ZN(n15958) );
  INV_X1 U20373 ( .A(n3635), .ZN(n27384) );
  NAND3_X1 U20374 ( .A1(n15956), .A2(n27384), .A3(n15955), .ZN(n15957) );
  NAND3_X1 U20375 ( .A1(n15959), .A2(n15958), .A3(n15957), .ZN(n15960) );
  XNOR2_X1 U20376 ( .A(n15961), .B(n15960), .ZN(n15962) );
  XNOR2_X1 U20377 ( .A(n15963), .B(n15962), .ZN(n16764) );
  INV_X1 U20378 ( .A(n16764), .ZN(n17278) );
  XNOR2_X1 U20379 ( .A(n15965), .B(n16636), .ZN(n15970) );
  XNOR2_X1 U20380 ( .A(n29084), .B(n3196), .ZN(n15967) );
  XNOR2_X1 U20381 ( .A(n16395), .B(n15967), .ZN(n15968) );
  XNOR2_X1 U20382 ( .A(n15968), .B(n16506), .ZN(n15969) );
  XNOR2_X1 U20383 ( .A(n15971), .B(n1184), .ZN(n15972) );
  INV_X1 U20384 ( .A(n16017), .ZN(n15974) );
  XNOR2_X1 U20385 ( .A(n15974), .B(n16619), .ZN(n16198) );
  XNOR2_X1 U20386 ( .A(n16575), .B(n16498), .ZN(n15976) );
  XNOR2_X1 U20387 ( .A(n16497), .B(n15976), .ZN(n15979) );
  XNOR2_X1 U20388 ( .A(n15977), .B(n3660), .ZN(n15978) );
  XNOR2_X1 U20389 ( .A(n16071), .B(n15982), .ZN(n15984) );
  INV_X1 U20390 ( .A(n16557), .ZN(n15983) );
  XNOR2_X1 U20391 ( .A(n15983), .B(n16070), .ZN(n16156) );
  XNOR2_X1 U20392 ( .A(n16156), .B(n15984), .ZN(n15988) );
  XNOR2_X1 U20393 ( .A(n16303), .B(n3180), .ZN(n15985) );
  XNOR2_X1 U20394 ( .A(n15986), .B(n15985), .ZN(n15987) );
  XNOR2_X1 U20395 ( .A(n15987), .B(n15988), .ZN(n17255) );
  XNOR2_X1 U20396 ( .A(n15989), .B(n26531), .ZN(n15990) );
  XNOR2_X1 U20397 ( .A(n15991), .B(n15990), .ZN(n15996) );
  XNOR2_X1 U20398 ( .A(n16170), .B(n15992), .ZN(n15993) );
  XNOR2_X1 U20399 ( .A(n15994), .B(n15993), .ZN(n15995) );
  INV_X1 U20401 ( .A(n17248), .ZN(n17016) );
  XNOR2_X1 U20402 ( .A(n15998), .B(n15997), .ZN(n16004) );
  XNOR2_X1 U20403 ( .A(n16641), .B(n1923), .ZN(n16002) );
  XNOR2_X1 U20404 ( .A(n15999), .B(n16000), .ZN(n16001) );
  XNOR2_X1 U20405 ( .A(n16002), .B(n16001), .ZN(n16003) );
  XNOR2_X1 U20406 ( .A(n16004), .B(n16003), .ZN(n17250) );
  INV_X1 U20407 ( .A(n17250), .ZN(n17017) );
  XNOR2_X1 U20408 ( .A(n16569), .B(n16216), .ZN(n16006) );
  XNOR2_X1 U20409 ( .A(n15914), .B(n16006), .ZN(n16007) );
  OAI21_X1 U20410 ( .B1(n17016), .B2(n17017), .A(n16977), .ZN(n16008) );
  XNOR2_X1 U20411 ( .A(n16009), .B(n16077), .ZN(n16159) );
  INV_X1 U20412 ( .A(n16159), .ZN(n16010) );
  XNOR2_X1 U20413 ( .A(n16010), .B(n16011), .ZN(n16016) );
  XNOR2_X1 U20414 ( .A(n16252), .B(n16012), .ZN(n16014) );
  XNOR2_X1 U20415 ( .A(n16256), .B(n5490), .ZN(n16013) );
  XNOR2_X1 U20416 ( .A(n16014), .B(n16013), .ZN(n16015) );
  AOI22_X1 U20417 ( .A1(n17251), .A2(n17249), .B1(n16977), .B2(n29503), .ZN(
        n17015) );
  XNOR2_X1 U20418 ( .A(n16246), .B(n16617), .ZN(n16021) );
  XNOR2_X1 U20419 ( .A(n16017), .B(n16165), .ZN(n16019) );
  XNOR2_X1 U20420 ( .A(n16607), .B(n2441), .ZN(n16018) );
  XNOR2_X1 U20421 ( .A(n16019), .B(n16018), .ZN(n16020) );
  OR2_X1 U20422 ( .A1(n17015), .A2(n6539), .ZN(n16022) );
  XNOR2_X1 U20424 ( .A(n16264), .B(n16023), .ZN(n16026) );
  XNOR2_X1 U20427 ( .A(n16404), .B(n27298), .ZN(n16027) );
  XNOR2_X1 U20428 ( .A(n16028), .B(n16027), .ZN(n16029) );
  INV_X1 U20430 ( .A(n16031), .ZN(n16033) );
  XNOR2_X1 U20431 ( .A(n16033), .B(n16032), .ZN(n16037) );
  XNOR2_X1 U20432 ( .A(n16377), .B(n16242), .ZN(n16035) );
  XNOR2_X1 U20433 ( .A(n16035), .B(n16034), .ZN(n16036) );
  XNOR2_X1 U20434 ( .A(n16037), .B(n16036), .ZN(n17098) );
  INV_X1 U20435 ( .A(n17098), .ZN(n16814) );
  XNOR2_X1 U20436 ( .A(n16038), .B(n16414), .ZN(n16040) );
  XNOR2_X1 U20437 ( .A(n16351), .B(n16040), .ZN(n16042) );
  XNOR2_X1 U20438 ( .A(n16255), .B(n3751), .ZN(n16041) );
  XNOR2_X1 U20439 ( .A(n16043), .B(n16365), .ZN(n16594) );
  INV_X1 U20440 ( .A(n16044), .ZN(n16045) );
  XNOR2_X1 U20441 ( .A(n16594), .B(n16045), .ZN(n16049) );
  XNOR2_X1 U20442 ( .A(n16229), .B(n16398), .ZN(n16047) );
  XNOR2_X1 U20443 ( .A(n16047), .B(n16046), .ZN(n16048) );
  XNOR2_X1 U20445 ( .A(n16051), .B(n16052), .ZN(n16054) );
  XNOR2_X1 U20446 ( .A(n16346), .B(n1248), .ZN(n16053) );
  XNOR2_X1 U20447 ( .A(n16054), .B(n16053), .ZN(n16055) );
  XNOR2_X1 U20448 ( .A(n320), .B(n3606), .ZN(n16056) );
  XNOR2_X1 U20449 ( .A(n16056), .B(n16567), .ZN(n16057) );
  XNOR2_X1 U20450 ( .A(n16058), .B(n16057), .ZN(n16064) );
  INV_X1 U20451 ( .A(n16059), .ZN(n16060) );
  XNOR2_X1 U20452 ( .A(n16271), .B(n16060), .ZN(n16061) );
  XNOR2_X1 U20453 ( .A(n16062), .B(n16061), .ZN(n16063) );
  NAND2_X1 U20454 ( .A1(n16860), .A2(n17097), .ZN(n16065) );
  MUX2_X1 U20455 ( .A(n16066), .B(n16065), .S(n17282), .Z(n16067) );
  XNOR2_X1 U20456 ( .A(n16262), .B(n3116), .ZN(n16068) );
  XNOR2_X1 U20457 ( .A(n16068), .B(n16405), .ZN(n16069) );
  XNOR2_X1 U20458 ( .A(n16300), .B(n16069), .ZN(n16074) );
  XNOR2_X1 U20459 ( .A(n16071), .B(n16070), .ZN(n16072) );
  XNOR2_X1 U20460 ( .A(n16654), .B(n16072), .ZN(n16073) );
  XNOR2_X1 U20461 ( .A(n16252), .B(n16625), .ZN(n16076) );
  XNOR2_X1 U20462 ( .A(n16323), .B(n16077), .ZN(n16079) );
  INV_X1 U20463 ( .A(n3625), .ZN(n28097) );
  XNOR2_X1 U20464 ( .A(n16257), .B(n28097), .ZN(n16078) );
  XNOR2_X1 U20465 ( .A(n16078), .B(n16079), .ZN(n16080) );
  XNOR2_X1 U20466 ( .A(n16081), .B(n16470), .ZN(n16083) );
  XNOR2_X1 U20467 ( .A(n16082), .B(n16083), .ZN(n16089) );
  XNOR2_X1 U20468 ( .A(n16328), .B(n16084), .ZN(n16087) );
  XNOR2_X1 U20469 ( .A(n16085), .B(n2598), .ZN(n16086) );
  XNOR2_X1 U20470 ( .A(n16087), .B(n16086), .ZN(n16088) );
  XNOR2_X1 U20471 ( .A(n16486), .B(n3015), .ZN(n16091) );
  XNOR2_X1 U20472 ( .A(n29571), .B(n16399), .ZN(n16092) );
  XNOR2_X1 U20473 ( .A(n16092), .B(n16636), .ZN(n16093) );
  AND2_X1 U20474 ( .A1(n17120), .A2(n16811), .ZN(n16100) );
  XNOR2_X1 U20475 ( .A(n29525), .B(n3154), .ZN(n16094) );
  XNOR2_X1 U20476 ( .A(n16094), .B(n16480), .ZN(n16097) );
  XNOR2_X1 U20477 ( .A(n16165), .B(n16095), .ZN(n16096) );
  XNOR2_X1 U20478 ( .A(n16097), .B(n16096), .ZN(n16099) );
  XNOR2_X1 U20479 ( .A(n16099), .B(n16098), .ZN(n17459) );
  INV_X1 U20480 ( .A(n17459), .ZN(n16676) );
  OAI21_X1 U20481 ( .B1(n16101), .B2(n16100), .A(n16676), .ZN(n16111) );
  AND2_X1 U20482 ( .A1(n17459), .A2(n16812), .ZN(n17113) );
  XNOR2_X1 U20483 ( .A(n16103), .B(n16102), .ZN(n16109) );
  INV_X1 U20484 ( .A(n3385), .ZN(n16104) );
  XNOR2_X1 U20485 ( .A(n16105), .B(n16104), .ZN(n16106) );
  XNOR2_X1 U20486 ( .A(n16107), .B(n16106), .ZN(n16108) );
  XNOR2_X1 U20487 ( .A(n16108), .B(n16109), .ZN(n16810) );
  INV_X1 U20488 ( .A(n29083), .ZN(n17457) );
  OAI21_X1 U20489 ( .B1(n17113), .B2(n16810), .A(n17457), .ZN(n16110) );
  NAND2_X1 U20490 ( .A1(n16111), .A2(n16110), .ZN(n17601) );
  INV_X1 U20491 ( .A(n16598), .ZN(n16113) );
  XNOR2_X1 U20492 ( .A(n16280), .B(n1196), .ZN(n16112) );
  XNOR2_X1 U20493 ( .A(n16113), .B(n16112), .ZN(n16118) );
  INV_X1 U20494 ( .A(n16366), .ZN(n16114) );
  XNOR2_X1 U20495 ( .A(n16634), .B(n16114), .ZN(n16115) );
  XNOR2_X1 U20496 ( .A(n16116), .B(n16115), .ZN(n16117) );
  XNOR2_X1 U20497 ( .A(n16510), .B(n3244), .ZN(n16120) );
  XNOR2_X1 U20498 ( .A(n16121), .B(n16120), .ZN(n16122) );
  INV_X1 U20499 ( .A(n16123), .ZN(n16125) );
  XNOR2_X1 U20500 ( .A(n16124), .B(n16125), .ZN(n16129) );
  XNOR2_X1 U20501 ( .A(n28557), .B(n28693), .ZN(n16127) );
  XNOR2_X1 U20502 ( .A(n16321), .B(n16126), .ZN(n16628) );
  XNOR2_X1 U20503 ( .A(n16127), .B(n16628), .ZN(n16128) );
  XNOR2_X1 U20504 ( .A(n16129), .B(n16128), .ZN(n16137) );
  XNOR2_X1 U20505 ( .A(n16130), .B(n16131), .ZN(n16132) );
  XNOR2_X1 U20506 ( .A(n16554), .B(n16132), .ZN(n16136) );
  XNOR2_X1 U20507 ( .A(n16653), .B(n1246), .ZN(n16133) );
  XNOR2_X1 U20508 ( .A(n16134), .B(n16133), .ZN(n16135) );
  XNOR2_X1 U20509 ( .A(n16136), .B(n16135), .ZN(n16668) );
  INV_X1 U20510 ( .A(n16137), .ZN(n16806) );
  XNOR2_X1 U20511 ( .A(n16527), .B(n16313), .ZN(n16616) );
  XNOR2_X1 U20512 ( .A(n16346), .B(n3062), .ZN(n16141) );
  XNOR2_X1 U20513 ( .A(n16143), .B(n21537), .ZN(n16144) );
  XNOR2_X1 U20514 ( .A(n16145), .B(n16144), .ZN(n16149) );
  XNOR2_X1 U20515 ( .A(n16291), .B(n16146), .ZN(n16647) );
  XNOR2_X1 U20516 ( .A(n16147), .B(n16647), .ZN(n16148) );
  XNOR2_X1 U20517 ( .A(n16148), .B(n16149), .ZN(n17260) );
  NAND2_X1 U20518 ( .A1(n17762), .A2(n17941), .ZN(n16152) );
  XNOR2_X1 U20519 ( .A(n16154), .B(n16302), .ZN(n16158) );
  XNOR2_X1 U20520 ( .A(n16558), .B(n24897), .ZN(n16155) );
  XNOR2_X1 U20521 ( .A(n16156), .B(n16155), .ZN(n16157) );
  XNOR2_X1 U20522 ( .A(n16320), .B(n16159), .ZN(n16164) );
  XNOR2_X1 U20523 ( .A(n16160), .B(n3697), .ZN(n16161) );
  XNOR2_X1 U20524 ( .A(n16162), .B(n16161), .ZN(n16163) );
  XNOR2_X1 U20525 ( .A(n16477), .B(n16165), .ZN(n16167) );
  XNOR2_X1 U20526 ( .A(n16607), .B(n3134), .ZN(n16168) );
  XNOR2_X1 U20527 ( .A(n16311), .B(n16168), .ZN(n16169) );
  XNOR2_X1 U20528 ( .A(n16192), .B(n16170), .ZN(n16595) );
  XNOR2_X1 U20529 ( .A(n16171), .B(n16595), .ZN(n16175) );
  XNOR2_X1 U20530 ( .A(n29571), .B(n2522), .ZN(n16173) );
  XNOR2_X1 U20531 ( .A(n16278), .B(n16173), .ZN(n16174) );
  INV_X1 U20532 ( .A(n16176), .ZN(n16204) );
  XNOR2_X1 U20533 ( .A(n16204), .B(n2446), .ZN(n16178) );
  XNOR2_X1 U20534 ( .A(n16178), .B(n16177), .ZN(n16181) );
  XNOR2_X1 U20535 ( .A(n16179), .B(n16331), .ZN(n16180) );
  XNOR2_X1 U20536 ( .A(n321), .B(n3334), .ZN(n16182) );
  XNOR2_X1 U20537 ( .A(n16182), .B(n16294), .ZN(n16184) );
  XNOR2_X1 U20538 ( .A(n16183), .B(n16184), .ZN(n16188) );
  XNOR2_X1 U20539 ( .A(n16569), .B(n16185), .ZN(n16186) );
  XNOR2_X1 U20540 ( .A(n16564), .B(n16186), .ZN(n16187) );
  XNOR2_X1 U20541 ( .A(n19650), .B(n19607), .ZN(n16698) );
  XNOR2_X1 U20542 ( .A(n16191), .B(n16190), .ZN(n16195) );
  XNOR2_X1 U20543 ( .A(n16192), .B(n2987), .ZN(n16193) );
  INV_X1 U20545 ( .A(n16888), .ZN(n17140) );
  XNOR2_X1 U20546 ( .A(n16199), .B(n16556), .ZN(n16202) );
  XNOR2_X1 U20547 ( .A(n16558), .B(n3483), .ZN(n16200) );
  XNOR2_X1 U20548 ( .A(n16206), .B(n16205), .ZN(n16210) );
  XNOR2_X1 U20549 ( .A(n16207), .B(n16208), .ZN(n16209) );
  NAND2_X1 U20550 ( .A1(n17140), .A2(n16887), .ZN(n16702) );
  INV_X1 U20551 ( .A(n16211), .ZN(n16212) );
  XNOR2_X1 U20552 ( .A(n16213), .B(n16212), .ZN(n16215) );
  XNOR2_X1 U20553 ( .A(n16215), .B(n16214), .ZN(n16220) );
  XNOR2_X1 U20554 ( .A(n16216), .B(n26909), .ZN(n16217) );
  XNOR2_X1 U20555 ( .A(n16218), .B(n16217), .ZN(n16219) );
  NAND2_X1 U20556 ( .A1(n16888), .A2(n17139), .ZN(n17136) );
  NAND2_X1 U20557 ( .A1(n16702), .A2(n17136), .ZN(n16227) );
  XNOR2_X1 U20558 ( .A(n16160), .B(n3666), .ZN(n16222) );
  XNOR2_X1 U20559 ( .A(n16221), .B(n16222), .ZN(n16226) );
  XNOR2_X1 U20560 ( .A(n16223), .B(n16224), .ZN(n16225) );
  XNOR2_X1 U20561 ( .A(n16231), .B(n16230), .ZN(n16235) );
  XNOR2_X1 U20562 ( .A(n16233), .B(n16232), .ZN(n16234) );
  XNOR2_X1 U20563 ( .A(n16235), .B(n16234), .ZN(n16236) );
  XNOR2_X1 U20564 ( .A(n16236), .B(n16237), .ZN(n16736) );
  XNOR2_X1 U20565 ( .A(n16238), .B(n730), .ZN(n16239) );
  XNOR2_X1 U20566 ( .A(n16240), .B(n16239), .ZN(n16245) );
  XNOR2_X1 U20567 ( .A(n16242), .B(n16241), .ZN(n16513) );
  XNOR2_X1 U20568 ( .A(n16513), .B(n16243), .ZN(n16244) );
  XNOR2_X1 U20569 ( .A(n16244), .B(n16245), .ZN(n17147) );
  NAND2_X1 U20570 ( .A1(n16736), .A2(n17147), .ZN(n17485) );
  XNOR2_X1 U20571 ( .A(n16525), .B(n16246), .ZN(n16251) );
  XNOR2_X1 U20572 ( .A(n16247), .B(n3067), .ZN(n16248) );
  XNOR2_X1 U20573 ( .A(n16249), .B(n16248), .ZN(n16250) );
  XNOR2_X1 U20574 ( .A(n16251), .B(n16250), .ZN(n17076) );
  XNOR2_X1 U20575 ( .A(n16252), .B(n16498), .ZN(n16254) );
  XNOR2_X1 U20576 ( .A(n16254), .B(n16253), .ZN(n16261) );
  XNOR2_X1 U20577 ( .A(n16256), .B(n16255), .ZN(n16259) );
  XNOR2_X1 U20578 ( .A(n16257), .B(n27894), .ZN(n16258) );
  XNOR2_X1 U20579 ( .A(n16258), .B(n16259), .ZN(n16260) );
  XNOR2_X2 U20580 ( .A(n16261), .B(n16260), .ZN(n17489) );
  OR2_X1 U20581 ( .A1(n17076), .A2(n17489), .ZN(n16735) );
  XNOR2_X1 U20582 ( .A(n16262), .B(n27225), .ZN(n16263) );
  XNOR2_X1 U20583 ( .A(n16263), .B(n28406), .ZN(n16265) );
  XNOR2_X1 U20584 ( .A(n16266), .B(n16265), .ZN(n16268) );
  MUX2_X1 U20585 ( .A(n17485), .B(n16735), .S(n17487), .Z(n16277) );
  INV_X1 U20586 ( .A(n16736), .ZN(n17078) );
  XNOR2_X1 U20587 ( .A(n16269), .B(n16270), .ZN(n16276) );
  XNOR2_X1 U20588 ( .A(n16271), .B(n16272), .ZN(n16274) );
  XNOR2_X1 U20589 ( .A(n16534), .B(n3686), .ZN(n16273) );
  XNOR2_X1 U20590 ( .A(n16274), .B(n16273), .ZN(n16275) );
  INV_X1 U20592 ( .A(n17487), .ZN(n17153) );
  INV_X1 U20593 ( .A(n17147), .ZN(n17146) );
  XNOR2_X1 U20594 ( .A(n16280), .B(n16279), .ZN(n16632) );
  XNOR2_X1 U20595 ( .A(n16281), .B(n16632), .ZN(n16288) );
  XNOR2_X1 U20596 ( .A(n16282), .B(n16283), .ZN(n16286) );
  XNOR2_X1 U20597 ( .A(n16284), .B(n3212), .ZN(n16285) );
  XNOR2_X1 U20598 ( .A(n16286), .B(n16285), .ZN(n16287) );
  XNOR2_X1 U20599 ( .A(n16288), .B(n16287), .ZN(n16612) );
  XNOR2_X1 U20600 ( .A(n320), .B(n1187), .ZN(n16290) );
  XNOR2_X1 U20601 ( .A(n16290), .B(n16291), .ZN(n16293) );
  XNOR2_X1 U20602 ( .A(n28579), .B(n16649), .ZN(n16358) );
  XNOR2_X1 U20603 ( .A(n16358), .B(n16293), .ZN(n16299) );
  XNOR2_X1 U20604 ( .A(n16295), .B(n16294), .ZN(n16297) );
  XNOR2_X1 U20605 ( .A(n16296), .B(n16297), .ZN(n16298) );
  XNOR2_X1 U20606 ( .A(n16299), .B(n16298), .ZN(n16730) );
  NOR2_X1 U20607 ( .A1(n16612), .A2(n17497), .ZN(n16337) );
  INV_X1 U20608 ( .A(n16300), .ZN(n16301) );
  XNOR2_X1 U20609 ( .A(n16301), .B(n16302), .ZN(n16308) );
  XNOR2_X1 U20610 ( .A(n16304), .B(n16303), .ZN(n16656) );
  XNOR2_X1 U20611 ( .A(n16305), .B(n3451), .ZN(n16306) );
  XNOR2_X1 U20612 ( .A(n16656), .B(n16306), .ZN(n16307) );
  XNOR2_X1 U20613 ( .A(n16310), .B(n16309), .ZN(n16344) );
  XNOR2_X1 U20614 ( .A(n16344), .B(n16311), .ZN(n16317) );
  XNOR2_X1 U20615 ( .A(n16480), .B(n16312), .ZN(n16315) );
  XNOR2_X1 U20616 ( .A(n16313), .B(n3414), .ZN(n16314) );
  XNOR2_X1 U20617 ( .A(n16315), .B(n16314), .ZN(n16316) );
  XNOR2_X1 U20618 ( .A(n16319), .B(n16318), .ZN(n16352) );
  XNOR2_X1 U20619 ( .A(n16320), .B(n16352), .ZN(n16327) );
  XNOR2_X1 U20620 ( .A(n16321), .B(n16322), .ZN(n16325) );
  XNOR2_X1 U20621 ( .A(n16323), .B(n3710), .ZN(n16324) );
  XNOR2_X1 U20622 ( .A(n16325), .B(n16324), .ZN(n16326) );
  XNOR2_X1 U20623 ( .A(n16327), .B(n16326), .ZN(n17498) );
  XNOR2_X1 U20624 ( .A(n16328), .B(n16329), .ZN(n16330) );
  XNOR2_X1 U20625 ( .A(n16331), .B(n16330), .ZN(n16336) );
  INV_X1 U20626 ( .A(n16640), .ZN(n16334) );
  XNOR2_X1 U20627 ( .A(n29516), .B(n2510), .ZN(n16333) );
  XNOR2_X1 U20628 ( .A(n16334), .B(n16333), .ZN(n16335) );
  NOR2_X1 U20629 ( .A1(n6079), .A2(n18465), .ZN(n16338) );
  XNOR2_X1 U20630 ( .A(n16303), .B(n3742), .ZN(n16341) );
  XNOR2_X1 U20631 ( .A(n16555), .B(n16341), .ZN(n16342) );
  INV_X1 U20632 ( .A(n16343), .ZN(n16345) );
  XNOR2_X1 U20633 ( .A(n16345), .B(n16344), .ZN(n16350) );
  XNOR2_X1 U20634 ( .A(n16346), .B(n2982), .ZN(n16348) );
  XNOR2_X1 U20635 ( .A(n16348), .B(n16347), .ZN(n16349) );
  INV_X1 U20636 ( .A(n16712), .ZN(n16381) );
  INV_X1 U20637 ( .A(n16351), .ZN(n16353) );
  XNOR2_X1 U20638 ( .A(n16353), .B(n16352), .ZN(n16357) );
  XNOR2_X1 U20639 ( .A(n6449), .B(n16579), .ZN(n16355) );
  INV_X1 U20640 ( .A(n2894), .ZN(n26877) );
  XNOR2_X1 U20641 ( .A(n29151), .B(n26877), .ZN(n16354) );
  XNOR2_X1 U20642 ( .A(n16355), .B(n16354), .ZN(n16356) );
  NAND2_X1 U20644 ( .A1(n16381), .A2(n28776), .ZN(n16383) );
  XNOR2_X1 U20646 ( .A(n16359), .B(n16358), .ZN(n16364) );
  XNOR2_X1 U20647 ( .A(n16360), .B(n3493), .ZN(n16361) );
  XNOR2_X1 U20648 ( .A(n16362), .B(n16361), .ZN(n16363) );
  INV_X1 U20649 ( .A(n17374), .ZN(n17173) );
  XNOR2_X1 U20650 ( .A(n16366), .B(n16365), .ZN(n16368) );
  XNOR2_X1 U20651 ( .A(n16367), .B(n16368), .ZN(n16372) );
  XNOR2_X1 U20652 ( .A(n16369), .B(n16370), .ZN(n16371) );
  XNOR2_X1 U20653 ( .A(n16373), .B(n16586), .ZN(n16374) );
  XNOR2_X1 U20654 ( .A(n16375), .B(n16374), .ZN(n16380) );
  INV_X1 U20655 ( .A(n16376), .ZN(n16379) );
  XNOR2_X1 U20656 ( .A(n16377), .B(n3463), .ZN(n16378) );
  NAND3_X1 U20657 ( .A1(n29635), .A2(n16381), .A3(n17375), .ZN(n16382) );
  XNOR2_X1 U20658 ( .A(n16509), .B(n28597), .ZN(n16385) );
  XNOR2_X1 U20659 ( .A(n16384), .B(n16385), .ZN(n16392) );
  XNOR2_X1 U20660 ( .A(n16387), .B(n16386), .ZN(n16390) );
  XNOR2_X1 U20661 ( .A(n16388), .B(n2960), .ZN(n16389) );
  XNOR2_X1 U20662 ( .A(n16390), .B(n16389), .ZN(n16391) );
  XNOR2_X1 U20663 ( .A(n16392), .B(n16391), .ZN(n16884) );
  INV_X1 U20664 ( .A(n16393), .ZN(n16394) );
  XNOR2_X1 U20665 ( .A(n16395), .B(n16394), .ZN(n16396) );
  XNOR2_X1 U20666 ( .A(n16397), .B(n16396), .ZN(n16403) );
  XNOR2_X1 U20667 ( .A(n16400), .B(n2306), .ZN(n16401) );
  XNOR2_X1 U20668 ( .A(n16488), .B(n16401), .ZN(n16402) );
  XNOR2_X1 U20669 ( .A(n16404), .B(n16405), .ZN(n16447) );
  XNOR2_X1 U20670 ( .A(n16406), .B(n16447), .ZN(n16413) );
  XNOR2_X1 U20671 ( .A(n16408), .B(n16407), .ZN(n16411) );
  XNOR2_X1 U20672 ( .A(n16409), .B(n27452), .ZN(n16410) );
  XNOR2_X1 U20673 ( .A(n16411), .B(n16410), .ZN(n16412) );
  XNOR2_X1 U20674 ( .A(n16415), .B(n16454), .ZN(n16420) );
  XNOR2_X1 U20675 ( .A(n16416), .B(n3527), .ZN(n16417) );
  XNOR2_X1 U20676 ( .A(n16418), .B(n16417), .ZN(n16419) );
  NOR2_X1 U20677 ( .A1(n17181), .A2(n17528), .ZN(n17531) );
  INV_X1 U20678 ( .A(n17531), .ZN(n16431) );
  XNOR2_X1 U20679 ( .A(n16422), .B(n16421), .ZN(n16423) );
  XNOR2_X1 U20680 ( .A(n16424), .B(n16423), .ZN(n16429) );
  XNOR2_X1 U20681 ( .A(n16425), .B(n16426), .ZN(n16464) );
  XNOR2_X1 U20682 ( .A(n16429), .B(n16428), .ZN(n16706) );
  INV_X1 U20683 ( .A(n16884), .ZN(n17157) );
  OAI22_X1 U20684 ( .A1(n6928), .A2(n16431), .B1(n16430), .B2(n17158), .ZN(
        n16441) );
  XNOR2_X1 U20685 ( .A(n16433), .B(n16432), .ZN(n16439) );
  XNOR2_X1 U20686 ( .A(n16434), .B(n16435), .ZN(n16478) );
  XNOR2_X1 U20687 ( .A(n16436), .B(n27462), .ZN(n16437) );
  XNOR2_X1 U20688 ( .A(n16437), .B(n16478), .ZN(n16438) );
  XNOR2_X1 U20689 ( .A(n16438), .B(n16439), .ZN(n17524) );
  NAND2_X1 U20690 ( .A1(n6928), .A2(n4979), .ZN(n16440) );
  XNOR2_X1 U20691 ( .A(n16443), .B(n3223), .ZN(n16446) );
  INV_X1 U20692 ( .A(n16444), .ZN(n16445) );
  XNOR2_X1 U20693 ( .A(n16446), .B(n16445), .ZN(n16448) );
  XNOR2_X1 U20694 ( .A(n16448), .B(n16447), .ZN(n16452) );
  XNOR2_X1 U20695 ( .A(n29511), .B(n16450), .ZN(n16451) );
  XNOR2_X1 U20696 ( .A(n16453), .B(n16454), .ZN(n16460) );
  XNOR2_X1 U20697 ( .A(n16456), .B(n3211), .ZN(n16457) );
  XNOR2_X1 U20698 ( .A(n16458), .B(n16457), .ZN(n16459) );
  XNOR2_X1 U20699 ( .A(n16460), .B(n16459), .ZN(n16549) );
  INV_X1 U20700 ( .A(n16549), .ZN(n17508) );
  XNOR2_X1 U20701 ( .A(n16461), .B(n16462), .ZN(n16466) );
  XNOR2_X1 U20702 ( .A(n16059), .B(n3752), .ZN(n16463) );
  XNOR2_X1 U20703 ( .A(n16464), .B(n16463), .ZN(n16465) );
  XNOR2_X1 U20704 ( .A(n16467), .B(n29247), .ZN(n16469) );
  XNOR2_X1 U20705 ( .A(n16468), .B(n16469), .ZN(n16475) );
  XNOR2_X1 U20706 ( .A(n28597), .B(n16471), .ZN(n16473) );
  XNOR2_X1 U20707 ( .A(n16472), .B(n16473), .ZN(n16474) );
  XNOR2_X1 U20708 ( .A(n16477), .B(n16476), .ZN(n16479) );
  XNOR2_X1 U20709 ( .A(n16480), .B(n3369), .ZN(n16482) );
  XNOR2_X1 U20710 ( .A(n15070), .B(n16483), .ZN(n16485) );
  XNOR2_X1 U20711 ( .A(n16484), .B(n16485), .ZN(n16490) );
  XNOR2_X1 U20712 ( .A(n16486), .B(n2381), .ZN(n16487) );
  XNOR2_X1 U20713 ( .A(n16487), .B(n16488), .ZN(n16489) );
  OAI21_X1 U20714 ( .B1(n4271), .B2(n17505), .A(n17506), .ZN(n16491) );
  INV_X1 U20715 ( .A(n18471), .ZN(n18464) );
  XNOR2_X1 U20716 ( .A(n16494), .B(n16495), .ZN(n16496) );
  XNOR2_X1 U20717 ( .A(n16497), .B(n16496), .ZN(n16502) );
  XNOR2_X1 U20718 ( .A(n16498), .B(n3770), .ZN(n16500) );
  XNOR2_X1 U20719 ( .A(n16499), .B(n16500), .ZN(n16501) );
  XNOR2_X1 U20720 ( .A(n16503), .B(n16504), .ZN(n16508) );
  INV_X1 U20721 ( .A(n17452), .ZN(n17067) );
  XNOR2_X1 U20722 ( .A(n16510), .B(n16509), .ZN(n16512) );
  XNOR2_X1 U20723 ( .A(n16512), .B(n16511), .ZN(n16516) );
  XNOR2_X1 U20724 ( .A(n16513), .B(n16514), .ZN(n16515) );
  INV_X1 U20725 ( .A(n17450), .ZN(n17066) );
  MUX2_X1 U20726 ( .A(n6772), .B(n17067), .S(n17066), .Z(n16539) );
  XNOR2_X1 U20727 ( .A(n16517), .B(n16518), .ZN(n16523) );
  XNOR2_X1 U20728 ( .A(n16519), .B(n3049), .ZN(n16520) );
  XNOR2_X1 U20729 ( .A(n16521), .B(n16520), .ZN(n16522) );
  XNOR2_X1 U20730 ( .A(n16523), .B(n16522), .ZN(n17455) );
  XNOR2_X1 U20731 ( .A(n16524), .B(n16525), .ZN(n16531) );
  XNOR2_X1 U20732 ( .A(n16526), .B(n16603), .ZN(n16529) );
  XNOR2_X1 U20733 ( .A(n16527), .B(n1062), .ZN(n16528) );
  XNOR2_X1 U20734 ( .A(n16529), .B(n16528), .ZN(n16530) );
  XNOR2_X1 U20735 ( .A(n16531), .B(n16530), .ZN(n17129) );
  INV_X1 U20736 ( .A(n17129), .ZN(n17068) );
  NOR2_X1 U20737 ( .A1(n28193), .A2(n16797), .ZN(n16538) );
  XNOR2_X1 U20738 ( .A(n16534), .B(n3633), .ZN(n16535) );
  XNOR2_X1 U20739 ( .A(n16536), .B(n16535), .ZN(n16537) );
  INV_X1 U20740 ( .A(n17456), .ZN(n17120) );
  NAND2_X1 U20741 ( .A1(n17120), .A2(n16810), .ZN(n16540) );
  AOI21_X1 U20742 ( .B1(n17117), .B2(n16540), .A(n16676), .ZN(n16545) );
  NAND2_X1 U20746 ( .A1(n18353), .A2(n16611), .ZN(n17918) );
  INV_X1 U20747 ( .A(n16728), .ZN(n16546) );
  NAND2_X1 U20748 ( .A1(n16546), .A2(n4271), .ZN(n16553) );
  NAND3_X1 U20749 ( .A1(n4271), .A2(n4270), .A3(n17505), .ZN(n16548) );
  BUF_X2 U20750 ( .A(n16549), .Z(n17830) );
  XNOR2_X1 U20751 ( .A(n16555), .B(n16554), .ZN(n16562) );
  XNOR2_X1 U20752 ( .A(n16557), .B(n16556), .ZN(n16560) );
  XNOR2_X1 U20753 ( .A(n16558), .B(n3219), .ZN(n16559) );
  XNOR2_X1 U20754 ( .A(n16560), .B(n16559), .ZN(n16561) );
  XNOR2_X1 U20755 ( .A(n16563), .B(n16564), .ZN(n16565) );
  XNOR2_X1 U20756 ( .A(n16566), .B(n16565), .ZN(n16573) );
  XNOR2_X1 U20757 ( .A(n16568), .B(n16567), .ZN(n16571) );
  XNOR2_X1 U20758 ( .A(n16569), .B(n3482), .ZN(n16570) );
  XNOR2_X1 U20759 ( .A(n16570), .B(n16571), .ZN(n16572) );
  INV_X1 U20760 ( .A(n17516), .ZN(n17083) );
  XNOR2_X1 U20761 ( .A(n16574), .B(n16575), .ZN(n16576) );
  XNOR2_X1 U20762 ( .A(n16577), .B(n16576), .ZN(n16584) );
  XNOR2_X1 U20763 ( .A(n16578), .B(n16579), .ZN(n16582) );
  XNOR2_X1 U20764 ( .A(n16580), .B(n22489), .ZN(n16581) );
  XNOR2_X1 U20765 ( .A(n16582), .B(n16581), .ZN(n16583) );
  XNOR2_X1 U20767 ( .A(n16585), .B(n16586), .ZN(n16587) );
  XNOR2_X1 U20768 ( .A(n16588), .B(n16587), .ZN(n16593) );
  XNOR2_X1 U20769 ( .A(n16589), .B(n2325), .ZN(n16590) );
  XNOR2_X1 U20770 ( .A(n16591), .B(n16590), .ZN(n16592) );
  XNOR2_X1 U20771 ( .A(n16593), .B(n16592), .ZN(n17469) );
  NOR2_X1 U20772 ( .A1(n29406), .A2(n17469), .ZN(n16601) );
  XNOR2_X1 U20773 ( .A(n16596), .B(n2353), .ZN(n16597) );
  XNOR2_X1 U20774 ( .A(n16598), .B(n16597), .ZN(n16599) );
  INV_X1 U20775 ( .A(n17518), .ZN(n17109) );
  INV_X1 U20776 ( .A(n16603), .ZN(n16604) );
  XNOR2_X1 U20777 ( .A(n16607), .B(n2912), .ZN(n16608) );
  XNOR2_X1 U20778 ( .A(n16609), .B(n16608), .ZN(n16610) );
  NAND2_X1 U20779 ( .A1(n536), .A2(n538), .ZN(n16614) );
  NOR2_X1 U20780 ( .A1(n29373), .A2(n17062), .ZN(n16613) );
  AOI21_X1 U20781 ( .B1(n16611), .B2(n18312), .A(n18353), .ZN(n16615) );
  XNOR2_X1 U20782 ( .A(n16616), .B(n16617), .ZN(n16624) );
  XNOR2_X1 U20783 ( .A(n16619), .B(n16618), .ZN(n16622) );
  XNOR2_X1 U20784 ( .A(n16620), .B(n1079), .ZN(n16621) );
  XNOR2_X1 U20785 ( .A(n16622), .B(n16621), .ZN(n16623) );
  XNOR2_X1 U20786 ( .A(n16625), .B(n3644), .ZN(n16626) );
  XNOR2_X1 U20787 ( .A(n16627), .B(n16626), .ZN(n16631) );
  XNOR2_X1 U20788 ( .A(n16629), .B(n16628), .ZN(n16630) );
  XNOR2_X1 U20789 ( .A(n16630), .B(n16631), .ZN(n17478) );
  NOR2_X1 U20790 ( .A1(n534), .A2(n3883), .ZN(n16660) );
  XNOR2_X1 U20791 ( .A(n16633), .B(n16632), .ZN(n16638) );
  XNOR2_X1 U20792 ( .A(n16634), .B(n3650), .ZN(n16635) );
  XNOR2_X1 U20793 ( .A(n16636), .B(n16635), .ZN(n16637) );
  INV_X1 U20794 ( .A(n16724), .ZN(n17481) );
  XNOR2_X1 U20795 ( .A(n16639), .B(n16640), .ZN(n16646) );
  XNOR2_X1 U20796 ( .A(n16642), .B(n16641), .ZN(n16644) );
  XNOR2_X1 U20797 ( .A(n16644), .B(n16643), .ZN(n16645) );
  XNOR2_X1 U20798 ( .A(n16648), .B(n16647), .ZN(n16652) );
  XNOR2_X1 U20799 ( .A(n16649), .B(n2986), .ZN(n16650) );
  XNOR2_X1 U20800 ( .A(n16652), .B(n16651), .ZN(n16691) );
  INV_X1 U20801 ( .A(n16691), .ZN(n16723) );
  XNOR2_X1 U20802 ( .A(n16653), .B(n2477), .ZN(n16655) );
  XNOR2_X1 U20803 ( .A(n16655), .B(n16654), .ZN(n16657) );
  XNOR2_X1 U20804 ( .A(n16657), .B(n16656), .ZN(n16659) );
  XNOR2_X1 U20805 ( .A(n16659), .B(n16658), .ZN(n17474) );
  NOR2_X1 U20806 ( .A1(n16661), .A2(n17667), .ZN(n16662) );
  NAND4_X1 U20807 ( .A1(n2055), .A2(n16663), .A3(n518), .A4(n16662), .ZN(
        n16664) );
  NOR2_X1 U20808 ( .A1(n17276), .A2(n17278), .ZN(n16665) );
  INV_X1 U20811 ( .A(n16685), .ZN(n17663) );
  INV_X1 U20812 ( .A(n16668), .ZN(n16805) );
  OAI211_X1 U20813 ( .C1(n17259), .C2(n16805), .A(n17260), .B(n16669), .ZN(
        n16671) );
  INV_X1 U20814 ( .A(n17466), .ZN(n16673) );
  AOI22_X1 U20815 ( .A1(n17090), .A2(n16675), .B1(n6830), .B2(n16674), .ZN(
        n16693) );
  NAND2_X1 U20816 ( .A1(n16810), .A2(n421), .ZN(n16678) );
  NAND2_X1 U20817 ( .A1(n16813), .A2(n29083), .ZN(n16677) );
  NAND2_X1 U20818 ( .A1(n29559), .A2(n16679), .ZN(n17284) );
  INV_X1 U20819 ( .A(n17283), .ZN(n16857) );
  OAI21_X1 U20820 ( .B1(n17284), .B2(n16857), .A(n16680), .ZN(n16688) );
  NAND2_X1 U20821 ( .A1(n16688), .A2(n17117), .ZN(n16683) );
  MUX2_X1 U20823 ( .A(n29086), .B(n17282), .S(n17101), .Z(n16681) );
  INV_X1 U20824 ( .A(n17102), .ZN(n16815) );
  NAND3_X1 U20825 ( .A1(n16681), .A2(n16815), .A3(n17117), .ZN(n16682) );
  NAND2_X1 U20826 ( .A1(n16683), .A2(n16682), .ZN(n16684) );
  NAND3_X1 U20827 ( .A1(n514), .A2(n16932), .A3(n16684), .ZN(n16694) );
  OAI21_X1 U20828 ( .B1(n16814), .B2(n17282), .A(n16815), .ZN(n16686) );
  NOR2_X1 U20829 ( .A1(n16687), .A2(n16686), .ZN(n16689) );
  AOI22_X1 U20830 ( .A1(n17475), .A2(n3883), .B1(n17476), .B2(n17477), .ZN(
        n16692) );
  XNOR2_X1 U20832 ( .A(n29505), .B(n3244), .ZN(n16695) );
  XNOR2_X1 U20833 ( .A(n16696), .B(n16695), .ZN(n16697) );
  XNOR2_X1 U20834 ( .A(n16698), .B(n16697), .ZN(n20551) );
  INV_X1 U20835 ( .A(n17385), .ZN(n17188) );
  MUX2_X1 U20836 ( .A(n17188), .B(n28497), .S(n16879), .Z(n16701) );
  INV_X1 U20837 ( .A(n16700), .ZN(n18069) );
  AND2_X1 U20838 ( .A1(n16702), .A2(n17139), .ZN(n16705) );
  NAND2_X1 U20840 ( .A1(n17139), .A2(n16887), .ZN(n17500) );
  NOR2_X1 U20841 ( .A1(n17500), .A2(n17502), .ZN(n16703) );
  NOR2_X1 U20842 ( .A1(n17087), .A2(n16703), .ZN(n16704) );
  NOR2_X1 U20844 ( .A1(n16706), .A2(n16883), .ZN(n18221) );
  INV_X1 U20845 ( .A(n18221), .ZN(n17532) );
  MUX2_X1 U20846 ( .A(n16707), .B(n17532), .S(n17158), .Z(n16708) );
  AOI21_X1 U20847 ( .B1(n17200), .B2(n17339), .A(n28564), .ZN(n16710) );
  NOR2_X1 U20848 ( .A1(n17338), .A2(n17204), .ZN(n16709) );
  NAND2_X1 U20849 ( .A1(n17336), .A2(n17204), .ZN(n16711) );
  INV_X1 U20850 ( .A(n16711), .ZN(n16936) );
  INV_X1 U20852 ( .A(n17357), .ZN(n17195) );
  OAI21_X1 U20854 ( .B1(n17198), .B2(n16713), .A(n17356), .ZN(n16716) );
  OAI21_X1 U20858 ( .B1(n16717), .B2(n29502), .A(n18195), .ZN(n16720) );
  OAI211_X1 U20859 ( .C1(n18195), .C2(n17746), .A(n16720), .B(n16719), .ZN(
        n18737) );
  NOR2_X1 U20860 ( .A1(n17129), .A2(n16797), .ZN(n16721) );
  NOR2_X1 U20861 ( .A1(n16723), .A2(n17124), .ZN(n16722) );
  INV_X1 U20862 ( .A(n17804), .ZN(n16747) );
  NAND3_X1 U20863 ( .A1(n4271), .A2(n17506), .A3(n17508), .ZN(n16729) );
  NOR2_X1 U20864 ( .A1(n17492), .A2(n17498), .ZN(n17495) );
  INV_X1 U20865 ( .A(n16730), .ZN(n16882) );
  NAND2_X1 U20866 ( .A1(n16882), .A2(n17491), .ZN(n16880) );
  OAI21_X1 U20868 ( .B1(n538), .B2(n16880), .A(n17493), .ZN(n16733) );
  NAND3_X1 U20869 ( .A1(n16880), .A2(n4314), .A3(n536), .ZN(n16732) );
  MUX2_X1 U20870 ( .A(n16735), .B(n16734), .S(n17078), .Z(n16739) );
  INV_X1 U20871 ( .A(n17486), .ZN(n16737) );
  AOI22_X1 U20872 ( .A1(n16737), .A2(n4655), .B1(n17488), .B2(n5737), .ZN(
        n16738) );
  NAND3_X1 U20873 ( .A1(n3995), .A2(n18276), .A3(n18204), .ZN(n16746) );
  INV_X1 U20874 ( .A(n17110), .ZN(n17520) );
  INV_X1 U20875 ( .A(n17469), .ZN(n17517) );
  NAND3_X1 U20876 ( .A1(n17109), .A2(n17106), .A3(n17517), .ZN(n16742) );
  NAND3_X1 U20877 ( .A1(n17518), .A2(n29406), .A3(n17083), .ZN(n16741) );
  NAND3_X1 U20878 ( .A1(n17106), .A2(n17470), .A3(n17469), .ZN(n16740) );
  NOR2_X1 U20880 ( .A1(n18203), .A2(n18277), .ZN(n16744) );
  OAI21_X1 U20881 ( .B1(n16744), .B2(n3994), .A(n16898), .ZN(n16745) );
  OAI211_X1 U20882 ( .C1(n16747), .C2(n16898), .A(n16746), .B(n16745), .ZN(
        n18899) );
  XNOR2_X1 U20883 ( .A(n18899), .B(n18737), .ZN(n19646) );
  NOR2_X1 U20884 ( .A1(n17025), .A2(n17344), .ZN(n17350) );
  NOR2_X1 U20885 ( .A1(n17029), .A2(n17347), .ZN(n16748) );
  NOR2_X1 U20887 ( .A1(n17348), .A2(n17347), .ZN(n16749) );
  OAI21_X1 U20888 ( .B1(n16749), .B2(n17029), .A(n17025), .ZN(n18093) );
  NOR2_X1 U20889 ( .A1(n17546), .A2(n17539), .ZN(n18091) );
  AOI21_X1 U20890 ( .B1(n18090), .B2(n18093), .A(n18091), .ZN(n16758) );
  OR2_X1 U20891 ( .A1(n17542), .A2(n17543), .ZN(n17215) );
  NOR2_X1 U20892 ( .A1(n16939), .A2(n17545), .ZN(n16750) );
  INV_X1 U20893 ( .A(n18096), .ZN(n16757) );
  MUX2_X1 U20894 ( .A(n17555), .B(n17556), .S(n17554), .Z(n16754) );
  OAI21_X1 U20895 ( .B1(n16913), .B2(n17221), .A(n29142), .ZN(n16753) );
  NOR2_X1 U20896 ( .A1(n16911), .A2(n16908), .ZN(n16752) );
  AOI22_X1 U20897 ( .A1(n16758), .A2(n16757), .B1(n18179), .B2(n18178), .ZN(
        n18442) );
  INV_X1 U20898 ( .A(n17234), .ZN(n17043) );
  NAND2_X1 U20899 ( .A1(n17046), .A2(n17365), .ZN(n16759) );
  INV_X1 U20900 ( .A(n17364), .ZN(n16761) );
  NAND2_X1 U20901 ( .A1(n16761), .A2(n6180), .ZN(n17788) );
  NAND3_X1 U20902 ( .A1(n16844), .A2(n17002), .A3(n17275), .ZN(n16765) );
  OAI21_X1 U20903 ( .B1(n17001), .B2(n16766), .A(n16765), .ZN(n16769) );
  NOR2_X1 U20904 ( .A1(n16767), .A2(n17271), .ZN(n16768) );
  INV_X1 U20905 ( .A(n18109), .ZN(n17799) );
  NOR2_X1 U20906 ( .A1(n17265), .A2(n16995), .ZN(n16772) );
  INV_X1 U20907 ( .A(n29600), .ZN(n16970) );
  NAND2_X1 U20909 ( .A1(n16772), .A2(n29600), .ZN(n16770) );
  OAI211_X2 U20910 ( .C1(n16772), .C2(n16773), .A(n16771), .B(n16770), .ZN(
        n18111) );
  NAND2_X1 U20911 ( .A1(n17248), .A2(n17017), .ZN(n16775) );
  NAND3_X1 U20912 ( .A1(n16865), .A2(n16775), .A3(n17249), .ZN(n16778) );
  NOR2_X1 U20913 ( .A1(n17016), .A2(n17249), .ZN(n16776) );
  NAND2_X1 U20914 ( .A1(n16776), .A2(n17251), .ZN(n16777) );
  NAND3_X1 U20915 ( .A1(n17799), .A2(n18111), .A3(n17903), .ZN(n16796) );
  NOR2_X1 U20916 ( .A1(n17259), .A2(n16779), .ZN(n16780) );
  NAND2_X1 U20917 ( .A1(n17425), .A2(n29088), .ZN(n16787) );
  NAND2_X1 U20918 ( .A1(n17428), .A2(n28194), .ZN(n16783) );
  NAND2_X1 U20919 ( .A1(n16974), .A2(n16783), .ZN(n16784) );
  NAND2_X1 U20920 ( .A1(n16784), .A2(n2826), .ZN(n16786) );
  NAND3_X1 U20921 ( .A1(n28792), .A2(n17005), .A3(n17720), .ZN(n16785) );
  NAND3_X1 U20922 ( .A1(n17799), .A2(n17902), .A3(n18107), .ZN(n16795) );
  INV_X1 U20923 ( .A(n17902), .ZN(n18459) );
  NAND2_X1 U20924 ( .A1(n17903), .A2(n18459), .ZN(n16794) );
  NAND2_X1 U20925 ( .A1(n17012), .A2(n29152), .ZN(n16789) );
  XNOR2_X1 U20926 ( .A(n19252), .B(n19549), .ZN(n19582) );
  XNOR2_X1 U20927 ( .A(n19646), .B(n19582), .ZN(n16871) );
  NAND2_X1 U20928 ( .A1(n28193), .A2(n16797), .ZN(n16798) );
  NAND2_X1 U20929 ( .A1(n16798), .A2(n17068), .ZN(n16799) );
  OAI211_X1 U20930 ( .C1(n16803), .C2(n3883), .A(n17124), .B(n17481), .ZN(
        n16804) );
  NAND2_X1 U20931 ( .A1(n16805), .A2(n29574), .ZN(n16809) );
  NAND2_X1 U20932 ( .A1(n17283), .A2(n1466), .ZN(n16816) );
  MUX2_X1 U20933 ( .A(n16817), .B(n16816), .S(n16815), .Z(n16818) );
  NOR2_X1 U20934 ( .A1(n18174), .A2(n18168), .ZN(n17689) );
  NOR2_X1 U20935 ( .A1(n29605), .A2(n17405), .ZN(n16823) );
  INV_X1 U20937 ( .A(n17401), .ZN(n17394) );
  INV_X1 U20938 ( .A(n16999), .ZN(n17293) );
  NOR2_X1 U20939 ( .A1(n17394), .A2(n17293), .ZN(n16824) );
  OAI211_X1 U20941 ( .C1(n17435), .C2(n29566), .A(n17437), .B(n336), .ZN(
        n16828) );
  NAND2_X1 U20942 ( .A1(n17298), .A2(n17413), .ZN(n17412) );
  NAND2_X1 U20943 ( .A1(n15811), .A2(n17413), .ZN(n16830) );
  NAND3_X1 U20945 ( .A1(n5430), .A2(n17297), .A3(n17411), .ZN(n16829) );
  NAND2_X1 U20946 ( .A1(n16922), .A2(n15811), .ZN(n16832) );
  AOI21_X1 U20947 ( .B1(n16985), .B2(n18188), .A(n29044), .ZN(n16842) );
  NOR2_X1 U20948 ( .A1(n17553), .A2(n17554), .ZN(n16834) );
  NOR2_X1 U20949 ( .A1(n17555), .A2(n16908), .ZN(n16833) );
  NAND2_X1 U20951 ( .A1(n17312), .A2(n16918), .ZN(n17563) );
  INV_X1 U20952 ( .A(n17563), .ZN(n16839) );
  XNOR2_X1 U20953 ( .A(n19474), .B(n18395), .ZN(n16869) );
  NOR2_X1 U20954 ( .A1(n17277), .A2(n17002), .ZN(n17273) );
  NOR2_X1 U20955 ( .A1(n17428), .A2(n28194), .ZN(n16845) );
  OAI21_X1 U20956 ( .B1(n16846), .B2(n16845), .A(n17425), .ZN(n16849) );
  OAI21_X1 U20957 ( .B1(n16973), .B2(n17428), .A(n2826), .ZN(n16848) );
  NAND2_X1 U20960 ( .A1(n17101), .A2(n16860), .ZN(n16856) );
  NAND2_X1 U20961 ( .A1(n16856), .A2(n17284), .ZN(n16858) );
  NAND2_X1 U20962 ( .A1(n16858), .A2(n16857), .ZN(n16859) );
  NOR2_X1 U20963 ( .A1(n16863), .A2(n29298), .ZN(n16864) );
  NOR2_X1 U20965 ( .A1(n18172), .A2(n18170), .ZN(n17688) );
  NOR2_X1 U20966 ( .A1(n17688), .A2(n17780), .ZN(n16872) );
  NAND2_X1 U20967 ( .A1(n28649), .A2(n16872), .ZN(n16873) );
  NAND3_X1 U20969 ( .A1(n17375), .A2(n17374), .A3(n16874), .ZN(n16875) );
  NAND3_X1 U20970 ( .A1(n17382), .A2(n17386), .A3(n17388), .ZN(n18071) );
  NAND2_X1 U20971 ( .A1(n16879), .A2(n17385), .ZN(n18070) );
  INV_X1 U20972 ( .A(n16880), .ZN(n16881) );
  MUX2_X1 U20973 ( .A(n17524), .B(n17527), .S(n17181), .Z(n16886) );
  INV_X1 U20974 ( .A(n18516), .ZN(n18078) );
  OAI211_X1 U20975 ( .C1(n29127), .C2(n17138), .A(n28574), .B(n17501), .ZN(
        n18073) );
  NOR2_X1 U20976 ( .A1(n17139), .A2(n17138), .ZN(n16889) );
  NOR2_X1 U20977 ( .A1(n18508), .A2(n18507), .ZN(n16896) );
  NOR2_X1 U20978 ( .A1(n17153), .A2(n17148), .ZN(n16890) );
  NOR2_X1 U20979 ( .A1(n17148), .A2(n17489), .ZN(n16891) );
  NAND2_X1 U20980 ( .A1(n17488), .A2(n16891), .ZN(n16894) );
  INV_X1 U20981 ( .A(n17076), .ZN(n17149) );
  NAND3_X1 U20982 ( .A1(n17153), .A2(n17489), .A3(n17149), .ZN(n16893) );
  NAND3_X1 U20983 ( .A1(n17487), .A2(n17147), .A3(n17148), .ZN(n16892) );
  NAND2_X1 U20985 ( .A1(n18509), .A2(n29057), .ZN(n16895) );
  XNOR2_X1 U20986 ( .A(n18906), .B(n19686), .ZN(n16903) );
  AND2_X1 U20987 ( .A1(n18203), .A2(n18277), .ZN(n16899) );
  OAI21_X1 U20988 ( .B1(n3994), .B2(n18203), .A(n17803), .ZN(n16897) );
  OAI21_X1 U20989 ( .B1(n17803), .B2(n16899), .A(n16897), .ZN(n16901) );
  AOI22_X1 U20990 ( .A1(n16899), .A2(n18276), .B1(n18279), .B2(n17696), .ZN(
        n16900) );
  XNOR2_X1 U20991 ( .A(n19111), .B(n25044), .ZN(n16902) );
  XNOR2_X1 U20992 ( .A(n16903), .B(n16902), .ZN(n16983) );
  MUX2_X1 U20993 ( .A(n17707), .B(n17573), .S(n423), .Z(n16905) );
  NAND2_X1 U20994 ( .A1(n29605), .A2(n17572), .ZN(n17406) );
  NAND2_X1 U20995 ( .A1(n17707), .A2(n17405), .ZN(n17322) );
  AND2_X1 U20996 ( .A1(n17322), .A2(n17406), .ZN(n17706) );
  NAND2_X1 U20997 ( .A1(n17038), .A2(n17568), .ZN(n16907) );
  INV_X1 U20998 ( .A(n17557), .ZN(n17219) );
  NOR2_X1 U20999 ( .A1(n17555), .A2(n17219), .ZN(n16910) );
  NOR2_X1 U21000 ( .A1(n29142), .A2(n16908), .ZN(n16909) );
  AOI22_X1 U21001 ( .A1(n16910), .A2(n16911), .B1(n16909), .B2(n17553), .ZN(
        n16915) );
  NOR2_X1 U21002 ( .A1(n16911), .A2(n17555), .ZN(n16912) );
  NAND2_X1 U21003 ( .A1(n16913), .A2(n16912), .ZN(n16914) );
  NOR2_X1 U21004 ( .A1(n17562), .A2(n17315), .ZN(n16920) );
  NOR2_X1 U21005 ( .A1(n17316), .A2(n17560), .ZN(n16919) );
  NAND2_X1 U21006 ( .A1(n16921), .A2(n17301), .ZN(n16923) );
  NAND2_X1 U21007 ( .A1(n18263), .A2(n18324), .ZN(n17985) );
  MUX2_X1 U21008 ( .A(n17434), .B(n17309), .S(n17435), .Z(n16928) );
  INV_X1 U21009 ( .A(n17435), .ZN(n16924) );
  NAND3_X1 U21010 ( .A1(n16924), .A2(n529), .A3(n337), .ZN(n16925) );
  INV_X1 U21011 ( .A(n18324), .ZN(n17895) );
  OAI22_X1 U21012 ( .A1(n17713), .A2(n17985), .B1(n29603), .B2(n17986), .ZN(
        n16929) );
  NAND2_X1 U21013 ( .A1(n16932), .A2(n17117), .ZN(n18341) );
  NOR2_X1 U21014 ( .A1(n18341), .A2(n18342), .ZN(n17665) );
  OAI21_X1 U21015 ( .B1(n17043), .B2(n17368), .A(n17233), .ZN(n16934) );
  MUX2_X1 U21016 ( .A(n17368), .B(n17365), .S(n17362), .Z(n16933) );
  INV_X1 U21017 ( .A(n17335), .ZN(n17342) );
  NOR2_X1 U21018 ( .A1(n17338), .A2(n17342), .ZN(n16935) );
  INV_X1 U21019 ( .A(n17542), .ZN(n16941) );
  OAI21_X1 U21020 ( .B1(n16941), .B2(n17539), .A(n17540), .ZN(n16942) );
  INV_X1 U21021 ( .A(n16943), .ZN(n17242) );
  NAND2_X1 U21022 ( .A1(n17552), .A2(n5398), .ZN(n16945) );
  AOI22_X1 U21023 ( .A1(n1121), .A2(n16949), .B1(n16948), .B2(n17029), .ZN(
        n16950) );
  NOR2_X1 U21024 ( .A1(n18538), .A2(n18527), .ZN(n16956) );
  NOR2_X1 U21025 ( .A1(n17356), .A2(n2449), .ZN(n16952) );
  NOR2_X1 U21026 ( .A1(n16953), .A2(n17359), .ZN(n16954) );
  AND2_X1 U21027 ( .A1(n17358), .A2(n16954), .ZN(n18530) );
  MUX2_X1 U21028 ( .A(n17402), .B(n17400), .S(n17394), .Z(n16961) );
  NOR2_X1 U21029 ( .A1(n17400), .A2(n17396), .ZN(n16959) );
  MUX2_X1 U21030 ( .A(n16959), .B(n16958), .S(n17402), .Z(n16960) );
  NOR2_X1 U21032 ( .A1(n17305), .A2(n16964), .ZN(n16965) );
  INV_X1 U21034 ( .A(n16995), .ZN(n16969) );
  NAND2_X1 U21036 ( .A1(n6539), .A2(n29503), .ZN(n16976) );
  NAND2_X1 U21037 ( .A1(n17018), .A2(n17249), .ZN(n16975) );
  MUX2_X1 U21038 ( .A(n16976), .B(n16975), .S(n17248), .Z(n16979) );
  NAND2_X1 U21039 ( .A1(n17248), .A2(n16977), .ZN(n16978) );
  XNOR2_X1 U21040 ( .A(n19634), .B(n19598), .ZN(n16982) );
  INV_X1 U21041 ( .A(n18088), .ZN(n16987) );
  INV_X1 U21042 ( .A(n16985), .ZN(n16986) );
  OAI21_X1 U21043 ( .B1(n527), .B2(n16987), .A(n18186), .ZN(n16988) );
  NOR2_X1 U21044 ( .A1(n29600), .A2(n16991), .ZN(n16994) );
  NAND2_X1 U21045 ( .A1(n16994), .A2(n29298), .ZN(n16997) );
  NAND2_X1 U21046 ( .A1(n16992), .A2(n16995), .ZN(n17264) );
  NAND3_X1 U21047 ( .A1(n17277), .A2(n17002), .A3(n17271), .ZN(n17003) );
  NOR2_X1 U21049 ( .A1(n2825), .A2(n17426), .ZN(n17006) );
  OAI211_X1 U21050 ( .C1(n6927), .C2(n18600), .A(n17014), .B(n17990), .ZN(
        n17024) );
  NAND2_X1 U21052 ( .A1(n2656), .A2(n28142), .ZN(n17023) );
  OAI211_X1 U21053 ( .C1(n17018), .C2(n17249), .A(n17017), .B(n17016), .ZN(
        n17019) );
  INV_X1 U21054 ( .A(n17019), .ZN(n17020) );
  INV_X1 U21055 ( .A(n17854), .ZN(n18599) );
  AND3_X1 U21056 ( .A1(n29065), .A2(n28142), .A3(n18599), .ZN(n17022) );
  AOI21_X2 U21057 ( .B1(n17024), .B2(n17023), .A(n17022), .ZN(n19507) );
  NAND2_X1 U21058 ( .A1(n17349), .A2(n17344), .ZN(n17027) );
  NAND2_X1 U21059 ( .A1(n17029), .A2(n17347), .ZN(n17026) );
  INV_X1 U21060 ( .A(n18338), .ZN(n18370) );
  OR2_X1 U21061 ( .A1(n17199), .A2(n17356), .ZN(n17036) );
  NAND2_X1 U21062 ( .A1(n29546), .A2(n17195), .ZN(n17033) );
  NAND3_X1 U21063 ( .A1(n17358), .A2(n28793), .A3(n17033), .ZN(n17035) );
  NOR2_X1 U21064 ( .A1(n18370), .A2(n18332), .ZN(n18001) );
  NAND2_X1 U21065 ( .A1(n17569), .A2(n17568), .ZN(n17039) );
  AOI21_X1 U21066 ( .B1(n17040), .B2(n17039), .A(n17038), .ZN(n17041) );
  MUX2_X1 U21067 ( .A(n17045), .B(n17044), .S(n17366), .Z(n17049) );
  NOR2_X1 U21068 ( .A1(n18338), .A2(n18332), .ZN(n17060) );
  INV_X1 U21069 ( .A(n17241), .ZN(n17052) );
  NOR2_X1 U21070 ( .A1(n17052), .A2(n17051), .ZN(n17053) );
  MUX2_X2 U21071 ( .A(n17054), .B(n17053), .S(n5398), .Z(n18337) );
  NAND2_X1 U21072 ( .A1(n17540), .A2(n17539), .ZN(n17057) );
  INV_X1 U21073 ( .A(n17545), .ZN(n17055) );
  AOI21_X1 U21074 ( .B1(n17057), .B2(n5695), .A(n15787), .ZN(n17058) );
  XNOR2_X1 U21075 ( .A(n19507), .B(n19096), .ZN(n19628) );
  OAI21_X1 U21076 ( .B1(n17497), .B2(n29373), .A(n17063), .ZN(n17064) );
  INV_X1 U21077 ( .A(n17206), .ZN(n18591) );
  NOR2_X1 U21078 ( .A1(n18591), .A2(n18588), .ZN(n18596) );
  INV_X1 U21080 ( .A(n17506), .ZN(n17071) );
  AND2_X1 U21081 ( .A1(n17074), .A2(n17071), .ZN(n17831) );
  MUX2_X1 U21082 ( .A(n17072), .B(n17831), .S(n17830), .Z(n17075) );
  OR2_X2 U21083 ( .A1(n17075), .A2(n17828), .ZN(n18124) );
  NAND2_X1 U21084 ( .A1(n5737), .A2(n17489), .ZN(n17080) );
  NAND2_X1 U21085 ( .A1(n17076), .A2(n17489), .ZN(n17077) );
  NAND2_X1 U21086 ( .A1(n17078), .A2(n17077), .ZN(n17079) );
  MUX2_X1 U21087 ( .A(n17080), .B(n17079), .S(n17147), .Z(n17081) );
  NOR2_X1 U21088 ( .A1(n18124), .A2(n18128), .ZN(n17082) );
  INV_X1 U21089 ( .A(n17515), .ZN(n17085) );
  AOI22_X1 U21090 ( .A1(n17840), .A2(n18595), .B1(n17835), .B2(n18124), .ZN(
        n17089) );
  NAND2_X1 U21091 ( .A1(n17090), .A2(n28800), .ZN(n17096) );
  NOR2_X1 U21092 ( .A1(n17093), .A2(n387), .ZN(n17092) );
  AOI21_X1 U21093 ( .B1(n17094), .B2(n17093), .A(n17092), .ZN(n17095) );
  INV_X1 U21094 ( .A(n18144), .ZN(n17627) );
  OAI21_X1 U21095 ( .B1(n17102), .B2(n1466), .A(n17099), .ZN(n17285) );
  NAND2_X1 U21096 ( .A1(n17285), .A2(n17283), .ZN(n17105) );
  NAND2_X1 U21097 ( .A1(n17110), .A2(n17106), .ZN(n17107) );
  NOR2_X1 U21098 ( .A1(n17110), .A2(n17109), .ZN(n17111) );
  INV_X1 U21100 ( .A(n17117), .ZN(n17121) );
  INV_X1 U21101 ( .A(n17118), .ZN(n17119) );
  NAND3_X1 U21102 ( .A1(n17481), .A2(n3883), .A3(n17476), .ZN(n17123) );
  NOR2_X1 U21103 ( .A1(n28193), .A2(n17450), .ZN(n17130) );
  AND2_X1 U21104 ( .A1(n17130), .A2(n17454), .ZN(n17131) );
  XNOR2_X1 U21105 ( .A(n18695), .B(n19697), .ZN(n17170) );
  AOI21_X1 U21106 ( .B1(n17136), .B2(n17135), .A(n28574), .ZN(n17145) );
  NAND3_X1 U21107 ( .A1(n17140), .A2(n17139), .A3(n17138), .ZN(n17141) );
  OAI21_X1 U21108 ( .B1(n17143), .B2(n17142), .A(n17141), .ZN(n17144) );
  AOI21_X1 U21109 ( .B1(n17488), .B2(n17146), .A(n17148), .ZN(n17154) );
  NOR2_X1 U21110 ( .A1(n17148), .A2(n17147), .ZN(n17150) );
  OAI21_X1 U21111 ( .B1(n17151), .B2(n17150), .A(n17149), .ZN(n17152) );
  AOI21_X1 U21112 ( .B1(n17156), .B2(n17338), .A(n17340), .ZN(n17994) );
  INV_X1 U21113 ( .A(n17181), .ZN(n17183) );
  NAND2_X1 U21114 ( .A1(n17159), .A2(n17382), .ZN(n17161) );
  NAND2_X1 U21115 ( .A1(n18069), .A2(n17385), .ZN(n17160) );
  INV_X1 U21118 ( .A(n18376), .ZN(n18000) );
  AOI22_X1 U21120 ( .A1(n18383), .A2(n17166), .B1(n17165), .B2(n18382), .ZN(
        n17167) );
  XNOR2_X1 U21121 ( .A(n19412), .B(n28097), .ZN(n17169) );
  XNOR2_X1 U21122 ( .A(n17170), .B(n17169), .ZN(n17171) );
  INV_X1 U21123 ( .A(n20551), .ZN(n17172) );
  MUX2_X1 U21124 ( .A(n29294), .B(n17375), .S(n17173), .Z(n17180) );
  NAND2_X1 U21126 ( .A1(n29294), .A2(n17374), .ZN(n17176) );
  MUX2_X1 U21127 ( .A(n17177), .B(n17176), .S(n28776), .Z(n17178) );
  NAND2_X1 U21128 ( .A1(n17182), .A2(n17181), .ZN(n17187) );
  OAI21_X1 U21129 ( .B1(n17527), .B2(n16884), .A(n531), .ZN(n17184) );
  NAND2_X1 U21130 ( .A1(n17184), .A2(n17183), .ZN(n17186) );
  INV_X1 U21131 ( .A(n18122), .ZN(n18418) );
  NOR2_X1 U21132 ( .A1(n417), .A2(n18418), .ZN(n17205) );
  NAND2_X1 U21133 ( .A1(n17386), .A2(n29045), .ZN(n17190) );
  NAND3_X1 U21134 ( .A1(n17382), .A2(n17188), .A3(n18069), .ZN(n17189) );
  AOI21_X1 U21135 ( .B1(n1121), .B2(n5420), .A(n17344), .ZN(n17194) );
  NAND2_X1 U21136 ( .A1(n17348), .A2(n17349), .ZN(n17193) );
  INV_X1 U21137 ( .A(n18121), .ZN(n18028) );
  OAI211_X1 U21138 ( .C1(n2449), .C2(n17196), .A(n17355), .B(n17195), .ZN(
        n17197) );
  NAND2_X1 U21139 ( .A1(n17340), .A2(n17201), .ZN(n17202) );
  AOI21_X1 U21140 ( .B1(n18128), .B2(n18126), .A(n18591), .ZN(n17209) );
  NOR2_X1 U21141 ( .A1(n18126), .A2(n18124), .ZN(n17208) );
  XNOR2_X1 U21142 ( .A(n19243), .B(n18690), .ZN(n19665) );
  INV_X1 U21143 ( .A(n18426), .ZN(n17212) );
  OAI21_X1 U21144 ( .B1(n18042), .B2(n17802), .A(n17824), .ZN(n17211) );
  NAND2_X1 U21145 ( .A1(n18423), .A2(n18421), .ZN(n17210) );
  MUX2_X1 U21146 ( .A(n17540), .B(n15787), .S(n17213), .Z(n17218) );
  NAND2_X1 U21147 ( .A1(n17540), .A2(n17545), .ZN(n17214) );
  MUX2_X1 U21148 ( .A(n17215), .B(n17214), .S(n15787), .Z(n17216) );
  OAI21_X1 U21149 ( .B1(n29142), .B2(n17221), .A(n17554), .ZN(n17222) );
  MUX2_X1 U21150 ( .A(n17223), .B(n17222), .S(n17556), .Z(n17225) );
  OAI21_X1 U21151 ( .B1(n29550), .B2(n17314), .A(n17560), .ZN(n17226) );
  NAND2_X1 U21152 ( .A1(n17228), .A2(n17229), .ZN(n17231) );
  AOI21_X1 U21153 ( .B1(n17233), .B2(n17234), .A(n17232), .ZN(n17238) );
  AOI21_X1 U21154 ( .B1(n17236), .B2(n17235), .A(n17369), .ZN(n17237) );
  NAND2_X1 U21155 ( .A1(n17549), .A2(n16762), .ZN(n17551) );
  NAND2_X1 U21156 ( .A1(n17241), .A2(n17240), .ZN(n17244) );
  NAND3_X1 U21157 ( .A1(n17242), .A2(n4624), .A3(n5398), .ZN(n17243) );
  XNOR2_X1 U21160 ( .A(n19246), .B(n19617), .ZN(n18722) );
  XNOR2_X1 U21161 ( .A(n18722), .B(n19665), .ZN(n17334) );
  MUX2_X1 U21162 ( .A(n1880), .B(n17249), .S(n17248), .Z(n17253) );
  NOR2_X1 U21163 ( .A1(n17251), .A2(n29503), .ZN(n17252) );
  INV_X1 U21164 ( .A(n18241), .ZN(n17843) );
  NAND2_X1 U21165 ( .A1(n17264), .A2(n17263), .ZN(n17270) );
  NAND2_X1 U21166 ( .A1(n17843), .A2(n17842), .ZN(n17290) );
  NOR2_X1 U21167 ( .A1(n17271), .A2(n17275), .ZN(n17274) );
  NOR2_X1 U21168 ( .A1(n18242), .A2(n17842), .ZN(n17970) );
  NOR2_X1 U21169 ( .A1(n28800), .A2(n17280), .ZN(n17281) );
  NAND2_X1 U21170 ( .A1(n17970), .A2(n17969), .ZN(n17289) );
  NAND2_X1 U21171 ( .A1(n17285), .A2(n17284), .ZN(n17286) );
  NOR2_X1 U21172 ( .A1(n17969), .A2(n18236), .ZN(n17287) );
  OAI21_X1 U21173 ( .B1(n17607), .B2(n17287), .A(n18241), .ZN(n17288) );
  OAI211_X1 U21175 ( .C1(n17400), .C2(n17294), .A(n29572), .B(n17293), .ZN(
        n17295) );
  INV_X1 U21176 ( .A(n17411), .ZN(n17416) );
  INV_X1 U21178 ( .A(n17423), .ZN(n17615) );
  OAI21_X1 U21181 ( .B1(n17309), .B2(n17439), .A(n17308), .ZN(n17311) );
  MUX2_X1 U21182 ( .A(n17435), .B(n17309), .S(n17438), .Z(n17310) );
  INV_X1 U21183 ( .A(n18156), .ZN(n18153) );
  INV_X1 U21184 ( .A(n17826), .ZN(n18154) );
  INV_X1 U21185 ( .A(n17405), .ZN(n17575) );
  NOR2_X1 U21186 ( .A1(n17707), .A2(n17575), .ZN(n17319) );
  MUX2_X1 U21187 ( .A(n17319), .B(n17318), .S(n17710), .Z(n17324) );
  NAND2_X1 U21188 ( .A1(n17320), .A2(n17575), .ZN(n17321) );
  AOI21_X1 U21189 ( .B1(n17322), .B2(n17321), .A(n29513), .ZN(n17323) );
  NOR2_X2 U21190 ( .A1(n17324), .A2(n17323), .ZN(n18032) );
  INV_X1 U21191 ( .A(n18032), .ZN(n17745) );
  NAND3_X1 U21192 ( .A1(n17745), .A2(n18160), .A3(n18153), .ZN(n17325) );
  XNOR2_X1 U21193 ( .A(n29554), .B(n29038), .ZN(n17332) );
  XNOR2_X1 U21195 ( .A(n19136), .B(n26531), .ZN(n17331) );
  XNOR2_X1 U21196 ( .A(n17332), .B(n17331), .ZN(n17333) );
  NOR2_X1 U21197 ( .A1(n17340), .A2(n17335), .ZN(n17337) );
  NAND3_X1 U21199 ( .A1(n17346), .A2(n17345), .A3(n29632), .ZN(n17352) );
  OAI21_X1 U21200 ( .B1(n17365), .B2(n17362), .A(n17361), .ZN(n17363) );
  NAND2_X1 U21201 ( .A1(n17364), .A2(n17363), .ZN(n17372) );
  NAND2_X1 U21202 ( .A1(n17366), .A2(n17365), .ZN(n17371) );
  NOR2_X1 U21203 ( .A1(n17368), .A2(n15731), .ZN(n17370) );
  OAI21_X1 U21204 ( .B1(n29636), .B2(n530), .A(n17374), .ZN(n17380) );
  NAND2_X1 U21205 ( .A1(n17375), .A2(n17374), .ZN(n17376) );
  NAND2_X1 U21206 ( .A1(n17377), .A2(n17376), .ZN(n17378) );
  AND2_X1 U21207 ( .A1(n28558), .A2(n18404), .ZN(n17381) );
  NAND2_X1 U21208 ( .A1(n18707), .A2(n17381), .ZN(n18712) );
  OAI21_X1 U21209 ( .B1(n17382), .B2(n29045), .A(n17385), .ZN(n17383) );
  NOR2_X1 U21210 ( .A1(n17388), .A2(n29045), .ZN(n17390) );
  OAI211_X1 U21211 ( .C1(n18707), .C2(n17392), .A(n18712), .B(n17391), .ZN(
        n17446) );
  OAI21_X1 U21212 ( .B1(n17397), .B2(n17396), .A(n17395), .ZN(n17398) );
  NAND2_X1 U21213 ( .A1(n17406), .A2(n17405), .ZN(n17407) );
  NAND2_X1 U21214 ( .A1(n5430), .A2(n17415), .ZN(n17410) );
  NAND3_X1 U21215 ( .A1(n17412), .A2(n17411), .A3(n17410), .ZN(n17419) );
  NAND3_X1 U21216 ( .A1(n17415), .A2(n17414), .A3(n17413), .ZN(n17418) );
  NAND3_X1 U21217 ( .A1(n18232), .A2(n17977), .A3(n18231), .ZN(n17445) );
  INV_X1 U21218 ( .A(n17425), .ZN(n17427) );
  NAND2_X1 U21219 ( .A1(n17427), .A2(n17426), .ZN(n17429) );
  MUX2_X1 U21220 ( .A(n17429), .B(n17428), .S(n28792), .Z(n17430) );
  INV_X1 U21221 ( .A(n18398), .ZN(n17442) );
  NAND2_X1 U21222 ( .A1(n17438), .A2(n17437), .ZN(n17441) );
  NAND3_X1 U21223 ( .A1(n17442), .A2(n18399), .A3(n18234), .ZN(n17444) );
  NAND3_X1 U21224 ( .A1(n18232), .A2(n18400), .A3(n18233), .ZN(n17443) );
  XNOR2_X1 U21225 ( .A(n19468), .B(n17446), .ZN(n19639) );
  NAND3_X1 U21226 ( .A1(n17762), .A2(n519), .A3(n517), .ZN(n17448) );
  AOI21_X1 U21227 ( .B1(n17762), .B2(n17872), .A(n17941), .ZN(n17447) );
  XNOR2_X1 U21228 ( .A(n18942), .B(n27737), .ZN(n17449) );
  XNOR2_X1 U21229 ( .A(n19639), .B(n17449), .ZN(n17581) );
  NOR2_X1 U21230 ( .A1(n17451), .A2(n17450), .ZN(n17453) );
  NAND2_X1 U21231 ( .A1(n17466), .A2(n17463), .ZN(n17465) );
  MUX2_X1 U21232 ( .A(n17467), .B(n17465), .S(n17464), .Z(n17468) );
  NAND2_X1 U21233 ( .A1(n17516), .A2(n17469), .ZN(n17514) );
  OR2_X1 U21234 ( .A1(n17514), .A2(n17470), .ZN(n17471) );
  NOR2_X1 U21235 ( .A1(n17477), .A2(n17476), .ZN(n17479) );
  NOR2_X1 U21236 ( .A1(n17505), .A2(n4270), .ZN(n17482) );
  NAND2_X1 U21238 ( .A1(n17484), .A2(n17506), .ZN(n17507) );
  OAI21_X1 U21239 ( .B1(n16736), .B2(n17487), .A(n17486), .ZN(n17490) );
  NOR2_X1 U21240 ( .A1(n17492), .A2(n17491), .ZN(n17494) );
  OAI21_X1 U21241 ( .B1(n17495), .B2(n17494), .A(n17493), .ZN(n18226) );
  NAND2_X1 U21243 ( .A1(n18388), .A2(n18393), .ZN(n18229) );
  OAI211_X1 U21244 ( .C1(n17506), .C2(n17505), .A(n17507), .B(n17829), .ZN(
        n17511) );
  INV_X1 U21245 ( .A(n17507), .ZN(n17509) );
  NAND2_X1 U21246 ( .A1(n17509), .A2(n17508), .ZN(n17510) );
  NAND2_X1 U21247 ( .A1(n17515), .A2(n17514), .ZN(n17521) );
  OAI21_X1 U21248 ( .B1(n17518), .B2(n17517), .A(n17516), .ZN(n17519) );
  AOI21_X1 U21249 ( .B1(n5234), .B2(n18393), .A(n18227), .ZN(n17522) );
  INV_X1 U21250 ( .A(n17522), .ZN(n17523) );
  OAI21_X1 U21252 ( .B1(n17526), .B2(n16884), .A(n17524), .ZN(n17530) );
  OAI21_X1 U21253 ( .B1(n17528), .B2(n17527), .A(n4979), .ZN(n17529) );
  INV_X1 U21254 ( .A(n18387), .ZN(n18391) );
  NAND3_X1 U21255 ( .A1(n5233), .A2(n18227), .A3(n18391), .ZN(n17533) );
  XNOR2_X1 U21256 ( .A(n19122), .B(n19377), .ZN(n17579) );
  NOR2_X1 U21258 ( .A1(n17969), .A2(n18243), .ZN(n17536) );
  NOR2_X1 U21259 ( .A1(n18241), .A2(n18236), .ZN(n17535) );
  NAND2_X1 U21260 ( .A1(n18243), .A2(n18241), .ZN(n17966) );
  NOR2_X1 U21261 ( .A1(n17542), .A2(n28454), .ZN(n17544) );
  MUX2_X1 U21262 ( .A(n16908), .B(n17554), .S(n17553), .Z(n17559) );
  MUX2_X1 U21263 ( .A(n17556), .B(n17555), .S(n17554), .Z(n17558) );
  INV_X1 U21264 ( .A(n17564), .ZN(n18253) );
  NAND2_X1 U21265 ( .A1(n17573), .A2(n17572), .ZN(n17574) );
  XNOR2_X1 U21266 ( .A(n19373), .B(n19555), .ZN(n19574) );
  XNOR2_X1 U21267 ( .A(n19574), .B(n17579), .ZN(n17580) );
  XNOR2_X1 U21268 ( .A(n17581), .B(n17580), .ZN(n19855) );
  NAND2_X1 U21269 ( .A1(n18251), .A2(n18253), .ZN(n17582) );
  INV_X1 U21270 ( .A(n6912), .ZN(n17962) );
  AOI21_X1 U21271 ( .B1(n17583), .B2(n17772), .A(n18251), .ZN(n17584) );
  NAND2_X1 U21273 ( .A1(n18214), .A2(n18506), .ZN(n17588) );
  NOR2_X1 U21274 ( .A1(n18500), .A2(n520), .ZN(n17586) );
  NAND2_X1 U21275 ( .A1(n18215), .A2(n17586), .ZN(n17587) );
  NAND2_X1 U21276 ( .A1(n17588), .A2(n17587), .ZN(n17591) );
  NAND2_X1 U21277 ( .A1(n520), .A2(n2363), .ZN(n17589) );
  NAND2_X1 U21278 ( .A1(n18388), .A2(n18387), .ZN(n17596) );
  INV_X1 U21279 ( .A(n18389), .ZN(n17593) );
  NAND2_X1 U21280 ( .A1(n17593), .A2(n17592), .ZN(n17595) );
  MUX2_X1 U21281 ( .A(n18707), .B(n18706), .S(n18404), .Z(n17600) );
  NOR2_X1 U21282 ( .A1(n18707), .A2(n18404), .ZN(n17599) );
  XNOR2_X1 U21283 ( .A(n19615), .B(n29038), .ZN(n17604) );
  XNOR2_X1 U21284 ( .A(n19490), .B(n26665), .ZN(n17603) );
  XNOR2_X1 U21285 ( .A(n17604), .B(n17603), .ZN(n17605) );
  AOI21_X1 U21286 ( .B1(n17757), .B2(n17756), .A(n18240), .ZN(n17608) );
  XNOR2_X1 U21287 ( .A(n18799), .B(n19256), .ZN(n17623) );
  AOI21_X1 U21289 ( .B1(n17610), .B2(n18431), .A(n18148), .ZN(n17611) );
  NAND3_X1 U21291 ( .A1(n17615), .A2(n17614), .A3(n17613), .ZN(n17618) );
  INV_X1 U21292 ( .A(n17616), .ZN(n17617) );
  NAND2_X1 U21293 ( .A1(n17825), .A2(n18033), .ZN(n17619) );
  OAI21_X1 U21294 ( .B1(n18160), .B2(n18156), .A(n17619), .ZN(n18036) );
  AOI21_X1 U21295 ( .B1(n17621), .B2(n17620), .A(n18153), .ZN(n17622) );
  XNOR2_X1 U21296 ( .A(n18408), .B(n18738), .ZN(n19362) );
  XNOR2_X1 U21297 ( .A(n17623), .B(n19362), .ZN(n17631) );
  NAND2_X1 U21298 ( .A1(n18028), .A2(n18414), .ZN(n17624) );
  OAI21_X1 U21299 ( .B1(n18413), .B2(n18122), .A(n17624), .ZN(n17625) );
  NAND2_X1 U21300 ( .A1(n18137), .A2(n17847), .ZN(n17626) );
  XNOR2_X1 U21301 ( .A(n18735), .B(n19584), .ZN(n17629) );
  XNOR2_X1 U21302 ( .A(n18949), .B(n1079), .ZN(n17628) );
  XNOR2_X1 U21303 ( .A(n17628), .B(n17629), .ZN(n17630) );
  NAND2_X1 U21304 ( .A1(n20414), .A2(n20941), .ZN(n17686) );
  INV_X1 U21305 ( .A(n20414), .ZN(n20192) );
  NOR2_X1 U21306 ( .A1(n18124), .A2(n18589), .ZN(n18592) );
  NOR2_X1 U21309 ( .A1(n17846), .A2(n18137), .ZN(n17635) );
  NAND2_X1 U21310 ( .A1(n17635), .A2(n17845), .ZN(n17638) );
  NAND3_X1 U21311 ( .A1(n18137), .A2(n526), .A3(n17847), .ZN(n17637) );
  XNOR2_X1 U21312 ( .A(n19215), .B(n19305), .ZN(n17644) );
  NAND2_X1 U21313 ( .A1(n18087), .A2(n18188), .ZN(n17642) );
  NOR2_X1 U21314 ( .A1(n18190), .A2(n29125), .ZN(n17641) );
  OAI211_X1 U21315 ( .C1(n17642), .C2(n17641), .A(n17640), .B(n17797), .ZN(
        n19339) );
  XNOR2_X1 U21316 ( .A(n19339), .B(n1187), .ZN(n17643) );
  XNOR2_X1 U21317 ( .A(n17644), .B(n17643), .ZN(n17656) );
  INV_X1 U21319 ( .A(n18382), .ZN(n17645) );
  NAND2_X1 U21320 ( .A1(n17645), .A2(n18379), .ZN(n18349) );
  NAND3_X1 U21321 ( .A1(n17883), .A2(n17647), .A3(n18376), .ZN(n17646) );
  NAND2_X1 U21323 ( .A1(n17883), .A2(n18376), .ZN(n18348) );
  NAND3_X1 U21324 ( .A1(n18348), .A2(n17647), .A3(n18380), .ZN(n17648) );
  XNOR2_X1 U21325 ( .A(n19686), .B(n19108), .ZN(n17654) );
  INV_X1 U21326 ( .A(n6927), .ZN(n17890) );
  NOR2_X1 U21327 ( .A1(n18338), .A2(n18372), .ZN(n17653) );
  XNOR2_X1 U21328 ( .A(n18773), .B(n19632), .ZN(n19597) );
  XNOR2_X1 U21329 ( .A(n19597), .B(n17654), .ZN(n17655) );
  NOR2_X1 U21331 ( .A1(n18465), .A2(n18471), .ZN(n18008) );
  NAND2_X1 U21332 ( .A1(n18008), .A2(n18469), .ZN(n17658) );
  NAND2_X1 U21333 ( .A1(n18314), .A2(n6079), .ZN(n17657) );
  XNOR2_X1 U21335 ( .A(n18942), .B(n3219), .ZN(n17662) );
  XNOR2_X1 U21336 ( .A(n19123), .B(n17662), .ZN(n17670) );
  INV_X1 U21337 ( .A(n18341), .ZN(n17908) );
  OAI21_X1 U21338 ( .B1(n17908), .B2(n514), .A(n18343), .ZN(n17664) );
  INV_X1 U21339 ( .A(n17947), .ZN(n18346) );
  NOR2_X1 U21340 ( .A1(n16611), .A2(n18312), .ZN(n17666) );
  INV_X1 U21341 ( .A(n18311), .ZN(n18357) );
  XNOR2_X1 U21342 ( .A(n19465), .B(n19232), .ZN(n17669) );
  XNOR2_X1 U21343 ( .A(n17670), .B(n17669), .ZN(n17684) );
  NAND3_X1 U21344 ( .A1(n29561), .A2(n18298), .A3(n18059), .ZN(n17673) );
  INV_X1 U21345 ( .A(n18057), .ZN(n17671) );
  NAND2_X1 U21346 ( .A1(n18298), .A2(n1861), .ZN(n17672) );
  NOR2_X1 U21347 ( .A1(n18493), .A2(n28632), .ZN(n18297) );
  MUX2_X1 U21349 ( .A(n17674), .B(n28633), .S(n18488), .Z(n17676) );
  XNOR2_X1 U21350 ( .A(n29318), .B(n18520), .ZN(n17683) );
  NOR2_X1 U21351 ( .A1(n18476), .A2(n18305), .ZN(n17677) );
  NAND2_X1 U21352 ( .A1(n17677), .A2(n18478), .ZN(n17678) );
  OAI21_X1 U21353 ( .B1(n18477), .B2(n18012), .A(n17678), .ZN(n17682) );
  NOR2_X1 U21354 ( .A1(n18476), .A2(n18306), .ZN(n18310) );
  INV_X1 U21355 ( .A(n18306), .ZN(n18474) );
  INV_X1 U21356 ( .A(n17679), .ZN(n17934) );
  NOR3_X1 U21357 ( .A1(n18310), .A2(n18011), .A3(n17680), .ZN(n17681) );
  XNOR2_X1 U21358 ( .A(n17683), .B(n19637), .ZN(n19336) );
  INV_X1 U21359 ( .A(n17687), .ZN(n20193) );
  NOR2_X1 U21360 ( .A1(n20414), .A2(n20193), .ZN(n17753) );
  XNOR2_X1 U21361 ( .A(n19707), .B(n29247), .ZN(n17690) );
  NOR2_X1 U21362 ( .A1(n510), .A2(n18078), .ZN(n17692) );
  NOR2_X1 U21363 ( .A1(n18510), .A2(n18508), .ZN(n17691) );
  INV_X1 U21365 ( .A(n18277), .ZN(n18275) );
  XNOR2_X1 U21366 ( .A(n19194), .B(n18913), .ZN(n17697) );
  NAND2_X1 U21368 ( .A1(n17700), .A2(n17699), .ZN(n17705) );
  AND2_X1 U21369 ( .A1(n18529), .A2(n18537), .ZN(n17701) );
  NOR3_X1 U21370 ( .A1(n18260), .A2(n17864), .A3(n18529), .ZN(n17702) );
  INV_X1 U21371 ( .A(n17706), .ZN(n17711) );
  OAI21_X1 U21372 ( .B1(n423), .B2(n17707), .A(n17710), .ZN(n17708) );
  OAI22_X1 U21373 ( .A1(n17711), .A2(n17710), .B1(n17709), .B2(n17708), .ZN(
        n17712) );
  INV_X1 U21374 ( .A(n18325), .ZN(n18322) );
  OR2_X1 U21375 ( .A1(n17717), .A2(n17431), .ZN(n17718) );
  XNOR2_X1 U21377 ( .A(n18369), .B(n28623), .ZN(n17725) );
  XNOR2_X1 U21378 ( .A(n17725), .B(n19603), .ZN(n19357) );
  XNOR2_X1 U21379 ( .A(n17726), .B(n19357), .ZN(n19747) );
  BUF_X2 U21380 ( .A(n19747), .Z(n20577) );
  AOI21_X2 U21381 ( .B1(n17728), .B2(n18217), .A(n17727), .ZN(n19321) );
  INV_X1 U21382 ( .A(n18107), .ZN(n18455) );
  XNOR2_X1 U21383 ( .A(n19321), .B(n19626), .ZN(n17742) );
  INV_X1 U21385 ( .A(n17592), .ZN(n17732) );
  INV_X1 U21387 ( .A(n18227), .ZN(n17766) );
  AND2_X1 U21388 ( .A1(n18390), .A2(n17766), .ZN(n17735) );
  NAND2_X1 U21389 ( .A1(n5233), .A2(n17592), .ZN(n17734) );
  INV_X1 U21391 ( .A(n17965), .ZN(n18960) );
  NOR2_X1 U21392 ( .A1(n18441), .A2(n18179), .ZN(n17737) );
  OAI21_X1 U21393 ( .B1(n18444), .B2(n18181), .A(n17737), .ZN(n17740) );
  XNOR2_X1 U21396 ( .A(n19331), .B(n18960), .ZN(n17741) );
  XNOR2_X1 U21397 ( .A(n17741), .B(n17742), .ZN(n17752) );
  NAND2_X1 U21398 ( .A1(n18156), .A2(n18154), .ZN(n18035) );
  NOR2_X1 U21399 ( .A1(n18160), .A2(n18032), .ZN(n18157) );
  NAND2_X1 U21400 ( .A1(n18159), .A2(n18034), .ZN(n17744) );
  AND2_X1 U21401 ( .A1(n18032), .A2(n18033), .ZN(n17743) );
  NAND3_X1 U21402 ( .A1(n17746), .A2(n29502), .A3(n18193), .ZN(n17748) );
  INV_X1 U21403 ( .A(n18449), .ZN(n18450) );
  NOR2_X1 U21404 ( .A1(n18450), .A2(n18198), .ZN(n17747) );
  XNOR2_X1 U21405 ( .A(n19332), .B(n18856), .ZN(n17750) );
  XNOR2_X1 U21406 ( .A(n19697), .B(n3666), .ZN(n17749) );
  XNOR2_X1 U21407 ( .A(n17750), .B(n17749), .ZN(n17751) );
  AOI22_X1 U21408 ( .A1(n17753), .A2(n20577), .B1(n503), .B2(n20412), .ZN(
        n17754) );
  NOR2_X1 U21409 ( .A1(n18506), .A2(n18500), .ZN(n17755) );
  NOR2_X1 U21410 ( .A1(n4725), .A2(n18236), .ZN(n17759) );
  NAND2_X1 U21411 ( .A1(n18240), .A2(n17842), .ZN(n17758) );
  OAI211_X1 U21412 ( .C1(n17977), .C2(n18402), .A(n18399), .B(n18400), .ZN(
        n17760) );
  OAI211_X1 U21413 ( .C1(n18397), .C2(n17977), .A(n18396), .B(n17760), .ZN(
        n19535) );
  XNOR2_X1 U21414 ( .A(n19084), .B(n19045), .ZN(n17779) );
  INV_X1 U21415 ( .A(n17761), .ZN(n17765) );
  OAI22_X1 U21416 ( .A1(n17937), .A2(n517), .B1(n17941), .B2(n17762), .ZN(
        n17873) );
  NAND2_X1 U21417 ( .A1(n18393), .A2(n17592), .ZN(n17769) );
  NAND3_X1 U21418 ( .A1(n17767), .A2(n18387), .A3(n18227), .ZN(n17768) );
  OAI21_X1 U21420 ( .B1(n18019), .B2(n1888), .A(n17773), .ZN(n17775) );
  XNOR2_X1 U21421 ( .A(n19481), .B(n19685), .ZN(n18670) );
  XNOR2_X1 U21425 ( .A(n18675), .B(n19378), .ZN(n17801) );
  NOR2_X1 U21426 ( .A1(n16985), .A2(n29125), .ZN(n17794) );
  NAND2_X1 U21427 ( .A1(n18087), .A2(n17794), .ZN(n19564) );
  OAI21_X1 U21428 ( .B1(n18087), .B2(n19560), .A(n29044), .ZN(n17795) );
  OAI21_X1 U21429 ( .B1(n17796), .B2(n29044), .A(n17795), .ZN(n19559) );
  OAI211_X1 U21430 ( .C1(n18188), .C2(n17797), .A(n19564), .B(n19559), .ZN(
        n19299) );
  XNOR2_X1 U21432 ( .A(n19077), .B(n17801), .ZN(n17813) );
  XNOR2_X1 U21433 ( .A(n28530), .B(n3622), .ZN(n17811) );
  NAND3_X1 U21434 ( .A1(n18450), .A2(n29502), .A3(n6663), .ZN(n17808) );
  XNOR2_X1 U21436 ( .A(n29492), .B(n19679), .ZN(n19156) );
  XNOR2_X1 U21437 ( .A(n19156), .B(n17811), .ZN(n17812) );
  XNOR2_X1 U21438 ( .A(n17813), .B(n17812), .ZN(n20310) );
  INV_X1 U21439 ( .A(n20310), .ZN(n20584) );
  XNOR2_X1 U21442 ( .A(n19283), .B(n19278), .ZN(n19105) );
  XNOR2_X1 U21443 ( .A(n19105), .B(n19285), .ZN(n17853) );
  INV_X1 U21444 ( .A(n17828), .ZN(n17833) );
  OAI21_X1 U21445 ( .B1(n17835), .B2(n17838), .A(n17834), .ZN(n17836) );
  NAND2_X1 U21446 ( .A1(n17840), .A2(n18128), .ZN(n17841) );
  NAND2_X1 U21448 ( .A1(n18241), .A2(n17842), .ZN(n18239) );
  XNOR2_X1 U21449 ( .A(n19704), .B(n19354), .ZN(n17851) );
  XNOR2_X1 U21450 ( .A(n17851), .B(n17850), .ZN(n17852) );
  XNOR2_X2 U21451 ( .A(n17853), .B(n17852), .ZN(n20585) );
  AOI22_X1 U21452 ( .A1(n17890), .A2(n18366), .B1(n18367), .B2(n2656), .ZN(
        n17855) );
  OR2_X1 U21453 ( .A1(n17855), .A2(n17854), .ZN(n17857) );
  AND2_X2 U21454 ( .A1(n17857), .A2(n17856), .ZN(n19359) );
  OAI22_X1 U21455 ( .A1(n17858), .A2(n374), .B1(n18286), .B2(n18081), .ZN(
        n17860) );
  XNOR2_X1 U21456 ( .A(n19359), .B(n19251), .ZN(n17865) );
  AOI21_X1 U21457 ( .B1(n18508), .B2(n18507), .A(n18510), .ZN(n17862) );
  XNOR2_X1 U21458 ( .A(n19725), .B(n19475), .ZN(n18681) );
  XNOR2_X1 U21459 ( .A(n17865), .B(n18681), .ZN(n17879) );
  NOR2_X1 U21460 ( .A1(n18500), .A2(n18213), .ZN(n18503) );
  NOR2_X1 U21461 ( .A1(n515), .A2(n17868), .ZN(n17869) );
  AOI22_X1 U21464 ( .A1(n18063), .A2(n18064), .B1(n18057), .B2(n17926), .ZN(
        n18303) );
  AOI21_X1 U21465 ( .B1(n17928), .B2(n1861), .A(n18059), .ZN(n17871) );
  XNOR2_X1 U21466 ( .A(n18760), .B(n19727), .ZN(n17877) );
  AOI21_X1 U21467 ( .B1(n17939), .B2(n28656), .A(n517), .ZN(n17875) );
  INV_X1 U21468 ( .A(n17942), .ZN(n17938) );
  XNOR2_X1 U21469 ( .A(n19643), .B(n1175), .ZN(n17876) );
  XNOR2_X1 U21470 ( .A(n17877), .B(n17876), .ZN(n17878) );
  XNOR2_X1 U21471 ( .A(n17879), .B(n17878), .ZN(n17954) );
  INV_X1 U21472 ( .A(n18350), .ZN(n17882) );
  NOR2_X1 U21473 ( .A1(n18382), .A2(n18379), .ZN(n18378) );
  AOI22_X1 U21474 ( .A1(n17882), .A2(n18000), .B1(n18378), .B2(n5383), .ZN(
        n17886) );
  NAND3_X1 U21475 ( .A1(n18383), .A2(n18382), .A3(n17883), .ZN(n17885) );
  MUX2_X1 U21476 ( .A(n18337), .B(n18372), .S(n18333), .Z(n17887) );
  INV_X1 U21477 ( .A(n18334), .ZN(n18371) );
  NOR2_X1 U21479 ( .A1(n17890), .A2(n29065), .ZN(n17891) );
  NOR2_X1 U21480 ( .A1(n17892), .A2(n6927), .ZN(n17893) );
  MUX2_X1 U21481 ( .A(n18262), .B(n17895), .S(n18325), .Z(n17897) );
  XNOR2_X1 U21482 ( .A(n19315), .B(n19066), .ZN(n17913) );
  NOR2_X1 U21483 ( .A1(n18311), .A2(n16611), .ZN(n17899) );
  INV_X1 U21484 ( .A(n18354), .ZN(n17898) );
  INV_X1 U21485 ( .A(n18312), .ZN(n18355) );
  NOR2_X1 U21486 ( .A1(n17918), .A2(n18355), .ZN(n17900) );
  XNOR2_X1 U21488 ( .A(n18778), .B(n19346), .ZN(n17911) );
  NOR2_X1 U21489 ( .A1(n18343), .A2(n18344), .ZN(n17909) );
  NOR2_X1 U21490 ( .A1(n514), .A2(n17947), .ZN(n17907) );
  XNOR2_X1 U21491 ( .A(n18646), .B(n2274), .ZN(n17910) );
  XNOR2_X1 U21492 ( .A(n17911), .B(n17910), .ZN(n17912) );
  XNOR2_X1 U21493 ( .A(n17913), .B(n17912), .ZN(n19827) );
  NOR2_X1 U21494 ( .A1(n20585), .A2(n19827), .ZN(n17956) );
  OAI21_X1 U21496 ( .B1(n145), .B2(n17917), .A(n18472), .ZN(n19173) );
  XNOR2_X1 U21499 ( .A(n18628), .B(n19692), .ZN(n17932) );
  AOI21_X1 U21500 ( .B1(n18493), .B2(n18292), .A(n28633), .ZN(n17925) );
  NOR2_X1 U21501 ( .A1(n18489), .A2(n18488), .ZN(n18293) );
  AOI21_X1 U21502 ( .B1(n18015), .B2(n18489), .A(n18293), .ZN(n17924) );
  OR2_X1 U21503 ( .A1(n18292), .A2(n18489), .ZN(n17923) );
  OAI21_X1 U21504 ( .B1(n17925), .B2(n17924), .A(n17923), .ZN(n18806) );
  NAND2_X1 U21505 ( .A1(n17928), .A2(n18064), .ZN(n17931) );
  NOR2_X1 U21506 ( .A1(n29561), .A2(n17926), .ZN(n17927) );
  XNOR2_X1 U21507 ( .A(n19508), .B(n18806), .ZN(n19322) );
  XNOR2_X1 U21508 ( .A(n19322), .B(n17932), .ZN(n17953) );
  NAND2_X1 U21509 ( .A1(n18304), .A2(n17934), .ZN(n17935) );
  INV_X1 U21510 ( .A(n18305), .ZN(n18479) );
  OAI22_X1 U21511 ( .A1(n18477), .A2(n17935), .B1(n18480), .B2(n18479), .ZN(
        n17936) );
  NAND2_X1 U21512 ( .A1(n17944), .A2(n17943), .ZN(n17945) );
  XNOR2_X1 U21513 ( .A(n19267), .B(n19323), .ZN(n19095) );
  NAND3_X1 U21515 ( .A1(n17948), .A2(n17947), .A3(n514), .ZN(n17949) );
  XNOR2_X1 U21516 ( .A(n19622), .B(n3654), .ZN(n17951) );
  XNOR2_X1 U21517 ( .A(n19095), .B(n17951), .ZN(n17952) );
  XNOR2_X1 U21518 ( .A(n17953), .B(n17952), .ZN(n20196) );
  NOR2_X1 U21519 ( .A1(n20196), .A2(n29144), .ZN(n17955) );
  MUX2_X1 U21520 ( .A(n17956), .B(n17955), .S(n20311), .Z(n17957) );
  NOR2_X1 U21521 ( .A1(n17960), .A2(n17959), .ZN(n17964) );
  OAI22_X1 U21522 ( .A1(n17961), .A2(n18253), .B1(n18018), .B2(n524), .ZN(
        n17963) );
  AOI21_X2 U21523 ( .B1(n17964), .B2(n17963), .A(n17962), .ZN(n19691) );
  XNOR2_X1 U21524 ( .A(n17965), .B(n19691), .ZN(n19210) );
  INV_X1 U21525 ( .A(n17966), .ZN(n17968) );
  OAI21_X1 U21526 ( .B1(n17968), .B2(n17967), .A(n18240), .ZN(n17973) );
  AOI22_X1 U21527 ( .A1(n29034), .A2(n17970), .B1(n17969), .B2(n4725), .ZN(
        n17972) );
  XNOR2_X1 U21528 ( .A(n17974), .B(n19409), .ZN(n17975) );
  XNOR2_X1 U21529 ( .A(n17975), .B(n19210), .ZN(n17984) );
  NAND3_X1 U21530 ( .A1(n17977), .A2(n18233), .A3(n18402), .ZN(n17978) );
  XNOR2_X1 U21531 ( .A(n19321), .B(n17982), .ZN(n17983) );
  XNOR2_X1 U21532 ( .A(n17984), .B(n17983), .ZN(n20199) );
  NOR2_X1 U21533 ( .A1(n18262), .A2(n18261), .ZN(n17987) );
  XNOR2_X1 U21534 ( .A(n18812), .B(n19462), .ZN(n17991) );
  XNOR2_X1 U21535 ( .A(n18815), .B(n17991), .ZN(n18005) );
  OR3_X1 U21536 ( .A1(n18383), .A2(n18382), .A3(n18376), .ZN(n17999) );
  INV_X1 U21537 ( .A(n17992), .ZN(n17993) );
  NAND2_X1 U21538 ( .A1(n17993), .A2(n2048), .ZN(n17995) );
  NOR3_X1 U21539 ( .A1(n18379), .A2(n17995), .A3(n17994), .ZN(n17996) );
  XNOR2_X1 U21540 ( .A(n19428), .B(n19232), .ZN(n19557) );
  XNOR2_X1 U21541 ( .A(n19427), .B(n3483), .ZN(n18003) );
  XNOR2_X1 U21542 ( .A(n19557), .B(n18003), .ZN(n18004) );
  NAND2_X1 U21543 ( .A1(n20199), .A2(n20200), .ZN(n20121) );
  INV_X1 U21544 ( .A(n18466), .ZN(n18006) );
  NOR3_X1 U21545 ( .A1(n18465), .A2(n18467), .A3(n18006), .ZN(n18007) );
  AOI21_X1 U21546 ( .B1(n6079), .B2(n18008), .A(n18007), .ZN(n18009) );
  XNOR2_X1 U21547 ( .A(n18735), .B(n18762), .ZN(n19548) );
  NAND2_X1 U21548 ( .A1(n18011), .A2(n18306), .ZN(n18013) );
  XNOR2_X1 U21551 ( .A(n18802), .B(n19198), .ZN(n19723) );
  XNOR2_X1 U21552 ( .A(n19723), .B(n19548), .ZN(n18025) );
  OAI21_X1 U21553 ( .B1(n18018), .B2(n18017), .A(n17771), .ZN(n18022) );
  XNOR2_X1 U21555 ( .A(n19440), .B(n3414), .ZN(n18023) );
  XNOR2_X1 U21556 ( .A(n19473), .B(n18023), .ZN(n18024) );
  XNOR2_X2 U21557 ( .A(n18024), .B(n18025), .ZN(n20302) );
  INV_X1 U21558 ( .A(n20199), .ZN(n20202) );
  XNOR2_X1 U21559 ( .A(n19273), .B(n3493), .ZN(n18031) );
  AOI21_X1 U21560 ( .B1(n18413), .B2(n18027), .A(n18122), .ZN(n18030) );
  NAND2_X1 U21561 ( .A1(n18028), .A2(n18122), .ZN(n18029) );
  XNOR2_X1 U21562 ( .A(n19215), .B(n18981), .ZN(n18966) );
  XNOR2_X1 U21563 ( .A(n18966), .B(n18031), .ZN(n18051) );
  AND2_X1 U21564 ( .A1(n18032), .A2(n18160), .ZN(n18039) );
  INV_X1 U21566 ( .A(n18164), .ZN(n18038) );
  NAND2_X1 U21567 ( .A1(n18036), .A2(n18035), .ZN(n18037) );
  OAI21_X1 U21568 ( .B1(n18039), .B2(n18038), .A(n18037), .ZN(n18633) );
  XNOR2_X1 U21569 ( .A(n18633), .B(n19305), .ZN(n18824) );
  NOR2_X1 U21570 ( .A1(n4805), .A2(n29507), .ZN(n18043) );
  INV_X1 U21571 ( .A(n18430), .ZN(n18432) );
  INV_X1 U21572 ( .A(n18146), .ZN(n18046) );
  NAND2_X1 U21573 ( .A1(n18046), .A2(n18431), .ZN(n18048) );
  NAND2_X1 U21574 ( .A1(n1758), .A2(n3467), .ZN(n18047) );
  XNOR2_X1 U21576 ( .A(n19421), .B(n19389), .ZN(n18622) );
  XNOR2_X1 U21577 ( .A(n18622), .B(n18824), .ZN(n18050) );
  XNOR2_X1 U21578 ( .A(n18050), .B(n18051), .ZN(n20201) );
  NOR2_X1 U21579 ( .A1(n18260), .A2(n18536), .ZN(n18052) );
  MUX2_X1 U21580 ( .A(n18054), .B(n18052), .S(n18539), .Z(n18056) );
  OAI21_X1 U21581 ( .B1(n18535), .B2(n18537), .A(n18536), .ZN(n18053) );
  NOR2_X2 U21582 ( .A1(n18056), .A2(n18055), .ZN(n19229) );
  AOI21_X1 U21583 ( .B1(n18059), .B2(n1861), .A(n18063), .ZN(n18058) );
  INV_X1 U21584 ( .A(n18058), .ZN(n18068) );
  NOR2_X1 U21585 ( .A1(n29561), .A2(n18059), .ZN(n18067) );
  INV_X1 U21586 ( .A(n18061), .ZN(n18062) );
  NAND3_X1 U21587 ( .A1(n18063), .A2(n18298), .A3(n18062), .ZN(n18066) );
  NAND2_X1 U21588 ( .A1(n18067), .A2(n18064), .ZN(n18065) );
  NAND3_X1 U21589 ( .A1(n18071), .A2(n18070), .A3(n18069), .ZN(n18072) );
  XNOR2_X1 U21590 ( .A(n19448), .B(n18725), .ZN(n19519) );
  XNOR2_X1 U21592 ( .A(n19717), .B(n18085), .ZN(n18791) );
  XNOR2_X1 U21593 ( .A(n18791), .B(n19519), .ZN(n18086) );
  XNOR2_X1 U21594 ( .A(n19452), .B(n19278), .ZN(n18099) );
  INV_X1 U21595 ( .A(n18090), .ZN(n18095) );
  INV_X1 U21596 ( .A(n18091), .ZN(n18092) );
  NAND2_X1 U21597 ( .A1(n18093), .A2(n18092), .ZN(n18094) );
  NOR3_X1 U21598 ( .A1(n18096), .A2(n18095), .A3(n18094), .ZN(n18097) );
  XNOR2_X1 U21599 ( .A(n18099), .B(n19702), .ZN(n18105) );
  NAND2_X1 U21600 ( .A1(n18100), .A2(n18452), .ZN(n18104) );
  XNOR2_X1 U21601 ( .A(n19194), .B(n19004), .ZN(n19541) );
  XNOR2_X1 U21602 ( .A(n18105), .B(n19541), .ZN(n18116) );
  MUX2_X1 U21603 ( .A(n18107), .B(n18111), .S(n18106), .Z(n18108) );
  NAND2_X1 U21604 ( .A1(n18108), .A2(n18456), .ZN(n18112) );
  NAND2_X1 U21605 ( .A1(n18111), .A2(n18109), .ZN(n18110) );
  XNOR2_X1 U21606 ( .A(n19700), .B(n2960), .ZN(n18113) );
  XNOR2_X1 U21607 ( .A(n18114), .B(n18113), .ZN(n18115) );
  MUX2_X1 U21608 ( .A(n18118), .B(n18117), .S(n19947), .Z(n18119) );
  AND3_X1 U21609 ( .A1(n18410), .A2(n18122), .A3(n18121), .ZN(n18123) );
  NOR3_X1 U21611 ( .A1(n18129), .A2(n18588), .A3(n18128), .ZN(n18132) );
  NOR2_X1 U21612 ( .A1(n18591), .A2(n18130), .ZN(n18131) );
  NOR3_X1 U21613 ( .A1(n18133), .A2(n18132), .A3(n18131), .ZN(n18134) );
  NAND3_X1 U21614 ( .A1(n18137), .A2(n18136), .A3(n3264), .ZN(n18139) );
  XNOR2_X1 U21615 ( .A(n18852), .B(n3317), .ZN(n18145) );
  AND3_X1 U21616 ( .A1(n18147), .A2(n18148), .A3(n18146), .ZN(n18152) );
  NOR2_X1 U21617 ( .A1(n18431), .A2(n18430), .ZN(n18150) );
  XNOR2_X1 U21618 ( .A(n19555), .B(n19376), .ZN(n18165) );
  OAI21_X1 U21619 ( .B1(n18155), .B2(n18154), .A(n18153), .ZN(n18163) );
  NAND2_X1 U21620 ( .A1(n18157), .A2(n18156), .ZN(n18162) );
  XNOR2_X1 U21622 ( .A(n28530), .B(n19678), .ZN(n19125) );
  XNOR2_X1 U21623 ( .A(n19125), .B(n18165), .ZN(n18166) );
  NAND2_X1 U21624 ( .A1(n4884), .A2(n18168), .ZN(n18169) );
  NAND2_X1 U21625 ( .A1(n18171), .A2(n18170), .ZN(n18175) );
  NAND3_X1 U21626 ( .A1(n513), .A2(n18179), .A3(n18180), .ZN(n18184) );
  NOR2_X1 U21627 ( .A1(n18181), .A2(n18180), .ZN(n18182) );
  NAND2_X1 U21628 ( .A1(n18182), .A2(n17793), .ZN(n18183) );
  XNOR2_X1 U21629 ( .A(n18880), .B(n19397), .ZN(n19065) );
  NAND2_X1 U21631 ( .A1(n18190), .A2(n18189), .ZN(n18191) );
  XNOR2_X1 U21633 ( .A(n19141), .B(n19065), .ZN(n18212) );
  MUX2_X1 U21635 ( .A(n18449), .B(n18195), .S(n18194), .Z(n18196) );
  INV_X1 U21636 ( .A(n18196), .ZN(n18202) );
  NOR2_X1 U21637 ( .A1(n18451), .A2(n18197), .ZN(n18201) );
  NAND2_X1 U21638 ( .A1(n18199), .A2(n18198), .ZN(n18200) );
  MUX2_X1 U21639 ( .A(n18203), .B(n18277), .S(n18204), .Z(n18205) );
  AND2_X1 U21640 ( .A1(n18275), .A2(n18204), .ZN(n18278) );
  AOI22_X1 U21641 ( .A1(n18205), .A2(n16898), .B1(n18278), .B2(n18279), .ZN(
        n18208) );
  NAND2_X1 U21642 ( .A1(n18206), .A2(n18276), .ZN(n18207) );
  XNOR2_X1 U21644 ( .A(n19617), .B(n3336), .ZN(n18209) );
  XNOR2_X1 U21645 ( .A(n18210), .B(n18209), .ZN(n18211) );
  XNOR2_X1 U21646 ( .A(n18212), .B(n18211), .ZN(n20544) );
  NOR3_X1 U21647 ( .A1(n18223), .A2(n18222), .A3(n18221), .ZN(n18225) );
  NAND3_X1 U21648 ( .A1(n18226), .A2(n18225), .A3(n18224), .ZN(n18228) );
  AOI21_X1 U21649 ( .B1(n18229), .B2(n18228), .A(n18227), .ZN(n18230) );
  XNOR2_X1 U21650 ( .A(n19024), .B(n18877), .ZN(n18583) );
  OAI21_X1 U21652 ( .B1(n18242), .B2(n18236), .A(n18243), .ZN(n18237) );
  AOI21_X1 U21653 ( .B1(n18238), .B2(n18242), .A(n18237), .ZN(n18246) );
  NOR2_X1 U21654 ( .A1(n18240), .A2(n18239), .ZN(n18245) );
  NOR3_X1 U21655 ( .A1(n18243), .A2(n18242), .A3(n18241), .ZN(n18244) );
  NOR3_X1 U21656 ( .A1(n18246), .A2(n18245), .A3(n18244), .ZN(n18247) );
  XNOR2_X1 U21657 ( .A(n18667), .B(n18247), .ZN(n19130) );
  XNOR2_X1 U21658 ( .A(n19130), .B(n18583), .ZN(n18258) );
  XNOR2_X1 U21659 ( .A(n19402), .B(n18256), .ZN(n18257) );
  MUX2_X1 U21660 ( .A(n19820), .B(n20544), .S(n20547), .Z(n18365) );
  XNOR2_X1 U21661 ( .A(n19525), .B(n1193), .ZN(n18269) );
  INV_X1 U21662 ( .A(n18326), .ZN(n18330) );
  NAND2_X1 U21663 ( .A1(n18330), .A2(n18261), .ZN(n18267) );
  OAI21_X1 U21664 ( .B1(n18326), .B2(n18324), .A(n18263), .ZN(n18264) );
  NAND2_X1 U21665 ( .A1(n18265), .A2(n18264), .ZN(n18266) );
  OAI21_X1 U21666 ( .B1(n18268), .B2(n18267), .A(n18266), .ZN(n18975) );
  XNOR2_X1 U21667 ( .A(n18975), .B(n19511), .ZN(n19410) );
  XNOR2_X1 U21668 ( .A(n19410), .B(n18269), .ZN(n18290) );
  INV_X1 U21669 ( .A(n18510), .ZN(n18271) );
  NAND3_X1 U21670 ( .A1(n18276), .A2(n18279), .A3(n18275), .ZN(n18284) );
  INV_X1 U21671 ( .A(n18276), .ZN(n18280) );
  NAND3_X1 U21672 ( .A1(n3995), .A2(n18280), .A3(n18277), .ZN(n18283) );
  INV_X1 U21673 ( .A(n18278), .ZN(n18282) );
  NAND3_X1 U21674 ( .A1(n18280), .A2(n16898), .A3(n18279), .ZN(n18281) );
  NAND4_X1 U21675 ( .A1(n18284), .A2(n18283), .A3(n18282), .A4(n18281), .ZN(
        n18857) );
  XNOR2_X1 U21676 ( .A(n18857), .B(n19320), .ZN(n18578) );
  XNOR2_X1 U21677 ( .A(n19695), .B(n19622), .ZN(n19116) );
  XNOR2_X1 U21678 ( .A(n19116), .B(n18578), .ZN(n18289) );
  XNOR2_X1 U21679 ( .A(n18290), .B(n18289), .ZN(n20388) );
  AND2_X1 U21680 ( .A1(n18291), .A2(n28633), .ZN(n18296) );
  NAND2_X1 U21681 ( .A1(n18292), .A2(n28633), .ZN(n18294) );
  NAND2_X1 U21682 ( .A1(n18294), .A2(n18293), .ZN(n18295) );
  NAND2_X1 U21683 ( .A1(n18301), .A2(n18300), .ZN(n18302) );
  XNOR2_X1 U21684 ( .A(n19631), .B(n19482), .ZN(n19391) );
  NAND3_X1 U21685 ( .A1(n18306), .A2(n17679), .A3(n18305), .ZN(n18307) );
  OAI21_X1 U21686 ( .B1(n18011), .B2(n17679), .A(n18307), .ZN(n18308) );
  XNOR2_X1 U21687 ( .A(n18868), .B(n19391), .ZN(n18321) );
  AOI21_X1 U21688 ( .B1(n18471), .B2(n18466), .A(n18467), .ZN(n18313) );
  NAND2_X1 U21690 ( .A1(n18465), .A2(n18315), .ZN(n18316) );
  OAI21_X2 U21691 ( .B1(n18318), .B2(n18317), .A(n18316), .ZN(n19306) );
  XNOR2_X1 U21692 ( .A(n19087), .B(n19306), .ZN(n18620) );
  XNOR2_X1 U21693 ( .A(n19534), .B(n1911), .ZN(n18319) );
  XNOR2_X1 U21694 ( .A(n18620), .B(n18319), .ZN(n18320) );
  MUX2_X1 U21695 ( .A(n20388), .B(n20539), .S(n19820), .Z(n18364) );
  NAND2_X1 U21696 ( .A1(n18323), .A2(n18322), .ZN(n18328) );
  NOR2_X1 U21697 ( .A1(n29603), .A2(n18324), .ZN(n18327) );
  XNOR2_X1 U21698 ( .A(n19359), .B(n19726), .ZN(n18862) );
  OAI21_X1 U21699 ( .B1(n18337), .B2(n18332), .A(n18331), .ZN(n18339) );
  XNOR2_X1 U21701 ( .A(n19384), .B(n18680), .ZN(n19071) );
  XNOR2_X1 U21702 ( .A(n18862), .B(n19071), .ZN(n18363) );
  AOI21_X1 U21703 ( .B1(n18349), .B2(n18348), .A(n18380), .ZN(n18352) );
  NAND2_X1 U21704 ( .A1(n18382), .A2(n18376), .ZN(n18351) );
  NOR2_X1 U21705 ( .A1(n18355), .A2(n18353), .ZN(n18360) );
  OAI21_X1 U21706 ( .B1(n18355), .B2(n18354), .A(n18356), .ZN(n18359) );
  XNOR2_X1 U21707 ( .A(n18798), .B(n18900), .ZN(n19472) );
  XNOR2_X1 U21708 ( .A(n19549), .B(n25992), .ZN(n18361) );
  XNOR2_X1 U21709 ( .A(n19472), .B(n18361), .ZN(n18362) );
  MUX2_X1 U21710 ( .A(n18365), .B(n18364), .S(n20546), .Z(n21346) );
  MUX2_X1 U21711 ( .A(n6314), .B(n21692), .S(n21346), .Z(n18548) );
  XNOR2_X1 U21712 ( .A(n19277), .B(n18638), .ZN(n18766) );
  MUX2_X2 U21713 ( .A(n18374), .B(n18373), .S(n18372), .Z(n19191) );
  XNOR2_X1 U21714 ( .A(n19700), .B(n19191), .ZN(n18375) );
  XNOR2_X1 U21715 ( .A(n18766), .B(n18375), .ZN(n18386) );
  AND2_X1 U21716 ( .A1(n18376), .A2(n18379), .ZN(n18377) );
  NOR2_X1 U21717 ( .A1(n18380), .A2(n18379), .ZN(n18381) );
  XNOR2_X1 U21718 ( .A(n29505), .B(n26032), .ZN(n18384) );
  XNOR2_X1 U21719 ( .A(n19356), .B(n18384), .ZN(n18385) );
  AOI22_X1 U21721 ( .A1(n29024), .A2(n18388), .B1(n17592), .B2(n18387), .ZN(
        n18394) );
  XNOR2_X1 U21724 ( .A(n18863), .B(n18395), .ZN(n18987) );
  OAI21_X1 U21725 ( .B1(n18707), .B2(n18706), .A(n4757), .ZN(n18407) );
  XNOR2_X1 U21726 ( .A(n28798), .B(n18948), .ZN(n18409) );
  NAND2_X1 U21727 ( .A1(n20290), .A2(n20295), .ZN(n20128) );
  INV_X1 U21728 ( .A(n18410), .ZN(n18412) );
  MUX2_X1 U21729 ( .A(n18413), .B(n18412), .S(n18411), .Z(n18419) );
  NAND3_X1 U21730 ( .A1(n18410), .A2(n417), .A3(n18414), .ZN(n18415) );
  XNOR2_X1 U21731 ( .A(n19409), .B(n19332), .ZN(n18420) );
  XNOR2_X1 U21732 ( .A(n19330), .B(n18420), .ZN(n18440) );
  NAND2_X1 U21733 ( .A1(n29507), .A2(n18421), .ZN(n18424) );
  AOI21_X1 U21734 ( .B1(n1942), .B2(n18424), .A(n18423), .ZN(n18428) );
  XNOR2_X1 U21735 ( .A(n19697), .B(n19592), .ZN(n18438) );
  XNOR2_X1 U21736 ( .A(n19207), .B(n3211), .ZN(n18437) );
  XNOR2_X1 U21737 ( .A(n18438), .B(n18437), .ZN(n18439) );
  XNOR2_X1 U21738 ( .A(n18440), .B(n18439), .ZN(n20125) );
  NAND2_X1 U21739 ( .A1(n18441), .A2(n523), .ZN(n18447) );
  INV_X1 U21740 ( .A(n18442), .ZN(n18443) );
  OAI21_X1 U21741 ( .B1(n18445), .B2(n18444), .A(n18443), .ZN(n18446) );
  XNOR2_X1 U21742 ( .A(n19686), .B(n19219), .ZN(n18967) );
  NAND3_X1 U21743 ( .A1(n18452), .A2(n6663), .A3(n18451), .ZN(n18453) );
  XNOR2_X1 U21744 ( .A(n19338), .B(n18967), .ZN(n18462) );
  XNOR2_X1 U21745 ( .A(n19595), .B(n19339), .ZN(n18774) );
  XNOR2_X1 U21746 ( .A(n19389), .B(n3633), .ZN(n18460) );
  XNOR2_X1 U21747 ( .A(n18774), .B(n18460), .ZN(n18461) );
  XNOR2_X1 U21748 ( .A(n18462), .B(n18461), .ZN(n19815) );
  NAND2_X1 U21749 ( .A1(n20125), .A2(n19815), .ZN(n18463) );
  NAND2_X1 U21750 ( .A1(n20128), .A2(n18463), .ZN(n18547) );
  NOR2_X1 U21751 ( .A1(n18465), .A2(n18464), .ZN(n18470) );
  NOR2_X1 U21752 ( .A1(n18467), .A2(n18466), .ZN(n18468) );
  NOR2_X1 U21753 ( .A1(n18472), .A2(n18471), .ZN(n18473) );
  XNOR2_X1 U21754 ( .A(n19225), .B(n19136), .ZN(n18991) );
  AOI21_X1 U21755 ( .B1(n18474), .B2(n18479), .A(n18477), .ZN(n18485) );
  AOI21_X1 U21756 ( .B1(n18478), .B2(n18475), .A(n18011), .ZN(n18484) );
  NOR3_X1 U21757 ( .A1(n18477), .A2(n18479), .A3(n18476), .ZN(n18482) );
  NOR3_X1 U21758 ( .A1(n18480), .A2(n18479), .A3(n18478), .ZN(n18481) );
  NOR2_X1 U21759 ( .A1(n18482), .A2(n18481), .ZN(n18483) );
  OAI21_X1 U21760 ( .B1(n18485), .B2(n18484), .A(n18483), .ZN(n19611) );
  XNOR2_X1 U21761 ( .A(n19611), .B(n19245), .ZN(n18779) );
  INV_X1 U21762 ( .A(n18488), .ZN(n18491) );
  XNOR2_X1 U21763 ( .A(n19228), .B(n2522), .ZN(n18497) );
  XNOR2_X1 U21764 ( .A(n19717), .B(n18935), .ZN(n18496) );
  XNOR2_X1 U21765 ( .A(n18497), .B(n18496), .ZN(n18498) );
  XNOR2_X1 U21766 ( .A(n18499), .B(n18498), .ZN(n20123) );
  NOR2_X1 U21767 ( .A1(n18500), .A2(n2363), .ZN(n18501) );
  AND2_X1 U21768 ( .A1(n18503), .A2(n18506), .ZN(n18504) );
  XNOR2_X1 U21771 ( .A(n18517), .B(n18652), .ZN(n19333) );
  XNOR2_X1 U21772 ( .A(n18942), .B(n3116), .ZN(n18518) );
  XNOR2_X1 U21773 ( .A(n18518), .B(n18812), .ZN(n18519) );
  XNOR2_X1 U21774 ( .A(n19333), .B(n18519), .ZN(n18545) );
  XNOR2_X1 U21775 ( .A(n19262), .B(n19577), .ZN(n18755) );
  NOR2_X1 U21776 ( .A1(n18528), .A2(n18527), .ZN(n18534) );
  MUX2_X1 U21779 ( .A(n18534), .B(n29327), .S(n509), .Z(n18543) );
  NOR2_X1 U21780 ( .A1(n18538), .A2(n18537), .ZN(n18540) );
  XNOR2_X1 U21781 ( .A(n28144), .B(n18755), .ZN(n18544) );
  XNOR2_X1 U21782 ( .A(n18544), .B(n18545), .ZN(n20293) );
  INV_X1 U21783 ( .A(n20290), .ZN(n19967) );
  INV_X1 U21785 ( .A(n19370), .ZN(n18550) );
  XNOR2_X1 U21786 ( .A(n19123), .B(n18550), .ZN(n18894) );
  XNOR2_X1 U21787 ( .A(n19122), .B(n19376), .ZN(n18551) );
  XNOR2_X1 U21788 ( .A(n18894), .B(n18551), .ZN(n18555) );
  XNOR2_X1 U21789 ( .A(n19636), .B(n19232), .ZN(n18553) );
  XNOR2_X1 U21790 ( .A(n19468), .B(n24897), .ZN(n18552) );
  XNOR2_X1 U21791 ( .A(n18552), .B(n18553), .ZN(n18554) );
  XNOR2_X1 U21792 ( .A(n19346), .B(n19397), .ZN(n19666) );
  XNOR2_X1 U21793 ( .A(n18556), .B(n19666), .ZN(n18560) );
  XNOR2_X1 U21794 ( .A(n19487), .B(n29554), .ZN(n18558) );
  XNOR2_X1 U21795 ( .A(n19136), .B(n857), .ZN(n18557) );
  XNOR2_X1 U21796 ( .A(n18558), .B(n18557), .ZN(n18559) );
  INV_X1 U21798 ( .A(n19194), .ZN(n18744) );
  XNOR2_X1 U21799 ( .A(n18744), .B(n2598), .ZN(n18561) );
  XNOR2_X1 U21800 ( .A(n19402), .B(n18561), .ZN(n18564) );
  XNOR2_X1 U21801 ( .A(n19495), .B(n19655), .ZN(n18562) );
  XNOR2_X1 U21802 ( .A(n18562), .B(n19133), .ZN(n18563) );
  XNOR2_X1 U21804 ( .A(n18695), .B(n18856), .ZN(n19117) );
  XNOR2_X1 U21805 ( .A(n19410), .B(n19117), .ZN(n18568) );
  XNOR2_X1 U21806 ( .A(n19507), .B(n18960), .ZN(n18566) );
  XNOR2_X1 U21807 ( .A(n19622), .B(n22489), .ZN(n18565) );
  XNOR2_X1 U21808 ( .A(n18566), .B(n18565), .ZN(n18567) );
  NOR2_X1 U21809 ( .A1(n29315), .A2(n20077), .ZN(n18573) );
  INV_X1 U21810 ( .A(n19384), .ZN(n19291) );
  XNOR2_X1 U21811 ( .A(n19291), .B(n19474), .ZN(n18989) );
  XNOR2_X1 U21812 ( .A(n18989), .B(n19359), .ZN(n19649) );
  XNOR2_X1 U21813 ( .A(n18569), .B(n18395), .ZN(n18571) );
  XNOR2_X1 U21814 ( .A(n19162), .B(n19256), .ZN(n18570) );
  XNOR2_X1 U21815 ( .A(n18571), .B(n18570), .ZN(n18572) );
  XNOR2_X1 U21816 ( .A(n19691), .B(n18628), .ZN(n18576) );
  XNOR2_X1 U21818 ( .A(n18578), .B(n18577), .ZN(n18579) );
  BUF_X2 U21820 ( .A(n18834), .Z(n20381) );
  XNOR2_X1 U21821 ( .A(n18581), .B(n19702), .ZN(n18582) );
  XNOR2_X1 U21822 ( .A(n18582), .B(n18583), .ZN(n18586) );
  XNOR2_X1 U21823 ( .A(n19700), .B(n3114), .ZN(n18584) );
  INV_X1 U21824 ( .A(n19004), .ZN(n18769) );
  XNOR2_X1 U21825 ( .A(n18769), .B(n18584), .ZN(n18585) );
  XNOR2_X1 U21827 ( .A(n18852), .B(n2465), .ZN(n18587) );
  XNOR2_X1 U21828 ( .A(n18587), .B(n19378), .ZN(n18597) );
  XNOR2_X1 U21829 ( .A(n19428), .B(n19300), .ZN(n18754) );
  XNOR2_X1 U21830 ( .A(n18597), .B(n18754), .ZN(n18609) );
  OR2_X1 U21831 ( .A1(n6927), .A2(n18598), .ZN(n18606) );
  MUX2_X1 U21832 ( .A(n28142), .B(n18600), .S(n18599), .Z(n18602) );
  NAND2_X1 U21833 ( .A1(n18602), .A2(n6927), .ZN(n18605) );
  AOI21_X1 U21834 ( .B1(n18606), .B2(n18605), .A(n18604), .ZN(n18607) );
  XNOR2_X1 U21835 ( .A(n18607), .B(n19427), .ZN(n18608) );
  INV_X1 U21836 ( .A(n20573), .ZN(n19837) );
  XNOR2_X1 U21837 ( .A(n19198), .B(n18762), .ZN(n19439) );
  XNOR2_X1 U21838 ( .A(n19039), .B(n19439), .ZN(n18612) );
  XNOR2_X1 U21839 ( .A(n18680), .B(n26825), .ZN(n18610) );
  XNOR2_X1 U21840 ( .A(n19727), .B(n18798), .ZN(n19289) );
  XNOR2_X1 U21841 ( .A(n18610), .B(n19289), .ZN(n18611) );
  XNOR2_X1 U21842 ( .A(n18612), .B(n18611), .ZN(n18613) );
  INV_X1 U21843 ( .A(n18613), .ZN(n19838) );
  AOI21_X1 U21844 ( .B1(n28637), .B2(n19837), .A(n19833), .ZN(n18627) );
  XNOR2_X1 U21846 ( .A(n18928), .B(n19229), .ZN(n19715) );
  XNOR2_X1 U21847 ( .A(n19399), .B(n19715), .ZN(n18617) );
  INV_X1 U21848 ( .A(n19491), .ZN(n19313) );
  XNOR2_X1 U21849 ( .A(n6489), .B(n18880), .ZN(n18615) );
  XNOR2_X1 U21850 ( .A(n19448), .B(n3035), .ZN(n18614) );
  XNOR2_X1 U21851 ( .A(n18615), .B(n18614), .ZN(n18616) );
  NAND2_X1 U21852 ( .A1(n29143), .A2(n20568), .ZN(n18625) );
  XNOR2_X1 U21853 ( .A(n18981), .B(n3722), .ZN(n18619) );
  INV_X1 U21854 ( .A(n19045), .ZN(n18618) );
  XNOR2_X1 U21855 ( .A(n18619), .B(n18618), .ZN(n18621) );
  XNOR2_X1 U21856 ( .A(n18621), .B(n18620), .ZN(n18623) );
  XNOR2_X1 U21857 ( .A(n18622), .B(n19535), .ZN(n19690) );
  MUX2_X1 U21858 ( .A(n18625), .B(n18624), .S(n28637), .Z(n18626) );
  XNOR2_X1 U21859 ( .A(n19321), .B(n18628), .ZN(n18629) );
  XNOR2_X1 U21860 ( .A(n19206), .B(n19692), .ZN(n18730) );
  XNOR2_X1 U21861 ( .A(n18629), .B(n18730), .ZN(n18632) );
  XNOR2_X1 U21862 ( .A(n19592), .B(n3164), .ZN(n18630) );
  XNOR2_X1 U21863 ( .A(n19528), .B(n18630), .ZN(n18631) );
  XNOR2_X1 U21864 ( .A(n19045), .B(n19595), .ZN(n18634) );
  INV_X1 U21865 ( .A(n18633), .ZN(n19423) );
  XNOR2_X1 U21866 ( .A(n19423), .B(n19219), .ZN(n19532) );
  XNOR2_X1 U21867 ( .A(n19532), .B(n18634), .ZN(n18637) );
  XNOR2_X1 U21868 ( .A(n19220), .B(n19687), .ZN(n18720) );
  XNOR2_X1 U21869 ( .A(n19305), .B(n3554), .ZN(n18635) );
  XNOR2_X1 U21870 ( .A(n18720), .B(n18635), .ZN(n18636) );
  XNOR2_X1 U21871 ( .A(n18637), .B(n18636), .ZN(n19849) );
  NOR2_X1 U21872 ( .A1(n20401), .A2(n29041), .ZN(n18650) );
  INV_X1 U21873 ( .A(n18114), .ZN(n19166) );
  XNOR2_X1 U21874 ( .A(n19166), .B(n18638), .ZN(n18639) );
  XNOR2_X1 U21875 ( .A(n19192), .B(n19704), .ZN(n18743) );
  XNOR2_X1 U21876 ( .A(n18743), .B(n18640), .ZN(n18641) );
  XNOR2_X1 U21877 ( .A(n18760), .B(n18863), .ZN(n18643) );
  XNOR2_X1 U21878 ( .A(n19643), .B(n27462), .ZN(n18642) );
  XNOR2_X1 U21879 ( .A(n18643), .B(n18642), .ZN(n18645) );
  XNOR2_X1 U21880 ( .A(n18948), .B(n19440), .ZN(n19546) );
  XNOR2_X1 U21881 ( .A(n19290), .B(n19546), .ZN(n18644) );
  XNOR2_X1 U21882 ( .A(n18644), .B(n18645), .ZN(n19851) );
  NOR2_X1 U21883 ( .A1(n20209), .A2(n19851), .ZN(n20559) );
  XNOR2_X1 U21884 ( .A(n18646), .B(n3374), .ZN(n18647) );
  XNOR2_X1 U21885 ( .A(n19225), .B(n18647), .ZN(n18648) );
  XNOR2_X1 U21886 ( .A(n19518), .B(n18648), .ZN(n18649) );
  XNOR2_X1 U21887 ( .A(n19611), .B(n19490), .ZN(n19317) );
  XNOR2_X1 U21888 ( .A(n18778), .B(n19317), .ZN(n19183) );
  XNOR2_X1 U21890 ( .A(n19577), .B(n19465), .ZN(n19296) );
  XNOR2_X1 U21891 ( .A(n28144), .B(n19378), .ZN(n18651) );
  XNOR2_X1 U21892 ( .A(n19296), .B(n18651), .ZN(n18657) );
  INV_X1 U21893 ( .A(n18652), .ZN(n19235) );
  XNOR2_X1 U21894 ( .A(n19568), .B(n19235), .ZN(n18655) );
  XNOR2_X1 U21895 ( .A(n29492), .B(n3607), .ZN(n18654) );
  XNOR2_X1 U21896 ( .A(n18655), .B(n18654), .ZN(n18656) );
  XNOR2_X1 U21897 ( .A(n18656), .B(n18657), .ZN(n20208) );
  NOR2_X1 U21898 ( .A1(n20208), .A2(n29041), .ZN(n20398) );
  OAI21_X1 U21899 ( .B1(n20398), .B2(n20401), .A(n20209), .ZN(n18658) );
  NAND2_X1 U21901 ( .A1(n29315), .A2(n29551), .ZN(n20075) );
  INV_X1 U21902 ( .A(n19391), .ZN(n18661) );
  XNOR2_X1 U21903 ( .A(n19215), .B(n19108), .ZN(n18660) );
  XNOR2_X1 U21904 ( .A(n18661), .B(n18660), .ZN(n18665) );
  XNOR2_X1 U21905 ( .A(n19111), .B(n19483), .ZN(n18663) );
  XNOR2_X1 U21906 ( .A(n18663), .B(n18662), .ZN(n18664) );
  XNOR2_X1 U21907 ( .A(n18665), .B(n18664), .ZN(n18838) );
  NOR2_X1 U21908 ( .A1(n20075), .A2(n18838), .ZN(n18753) );
  INV_X1 U21909 ( .A(n18753), .ZN(n19914) );
  XNOR2_X1 U21911 ( .A(n19285), .B(n18666), .ZN(n18669) );
  XNOR2_X1 U21912 ( .A(n18912), .B(n18877), .ZN(n19102) );
  INV_X1 U21913 ( .A(n18667), .ZN(n19709) );
  XNOR2_X1 U21914 ( .A(n19709), .B(n19278), .ZN(n19502) );
  XNOR2_X1 U21915 ( .A(n19102), .B(n19502), .ZN(n18668) );
  XNOR2_X1 U21916 ( .A(n18668), .B(n18669), .ZN(n18843) );
  INV_X1 U21917 ( .A(n18843), .ZN(n20372) );
  XNOR2_X1 U21918 ( .A(n19688), .B(n19273), .ZN(n19480) );
  XNOR2_X1 U21919 ( .A(n19480), .B(n18670), .ZN(n18674) );
  XNOR2_X1 U21920 ( .A(n18906), .B(n19087), .ZN(n18672) );
  XNOR2_X1 U21922 ( .A(n18672), .B(n18671), .ZN(n18673) );
  INV_X1 U21924 ( .A(n20374), .ZN(n19739) );
  XNOR2_X1 U21925 ( .A(n29580), .B(n19679), .ZN(n19298) );
  XNOR2_X1 U21926 ( .A(n18852), .B(n19377), .ZN(n19078) );
  XNOR2_X1 U21927 ( .A(n19298), .B(n19078), .ZN(n18679) );
  XNOR2_X1 U21928 ( .A(n19122), .B(n19462), .ZN(n18677) );
  INV_X1 U21929 ( .A(n1247), .ZN(n26701) );
  XNOR2_X1 U21930 ( .A(n19464), .B(n26701), .ZN(n18676) );
  XNOR2_X1 U21931 ( .A(n18677), .B(n18676), .ZN(n18678) );
  NOR3_X1 U21932 ( .A1(n20372), .A2(n19739), .A3(n20375), .ZN(n18688) );
  INV_X1 U21933 ( .A(n18680), .ZN(n19250) );
  XNOR2_X1 U21934 ( .A(n19250), .B(n18395), .ZN(n18682) );
  XNOR2_X1 U21935 ( .A(n18681), .B(n18682), .ZN(n18686) );
  XNOR2_X1 U21936 ( .A(n19251), .B(n19726), .ZN(n18684) );
  XNOR2_X1 U21937 ( .A(n18899), .B(n2385), .ZN(n18683) );
  XNOR2_X1 U21938 ( .A(n18684), .B(n18683), .ZN(n18685) );
  NOR2_X1 U21939 ( .A1(n20071), .A2(n20374), .ZN(n18687) );
  XNOR2_X1 U21940 ( .A(n19136), .B(n1225), .ZN(n18689) );
  INV_X1 U21941 ( .A(n19486), .ZN(n19716) );
  XNOR2_X1 U21942 ( .A(n19716), .B(n18927), .ZN(n18692) );
  XNOR2_X1 U21943 ( .A(n18692), .B(n18691), .ZN(n18693) );
  NAND2_X1 U21944 ( .A1(n20373), .A2(n18699), .ZN(n18701) );
  XNOR2_X1 U21945 ( .A(n19267), .B(n19695), .ZN(n19513) );
  XNOR2_X1 U21946 ( .A(n19322), .B(n19513), .ZN(n18698) );
  XNOR2_X1 U21947 ( .A(n18695), .B(n3660), .ZN(n18696) );
  XNOR2_X1 U21948 ( .A(n18696), .B(n19097), .ZN(n18697) );
  XNOR2_X1 U21949 ( .A(n18698), .B(n18697), .ZN(n19841) );
  INV_X1 U21950 ( .A(n18699), .ZN(n19740) );
  NAND3_X1 U21951 ( .A1(n19841), .A2(n351), .A3(n19740), .ZN(n18700) );
  OAI21_X1 U21952 ( .B1(n18843), .B2(n18701), .A(n18700), .ZN(n18702) );
  NOR2_X2 U21953 ( .A1(n18703), .A2(n18702), .ZN(n20972) );
  INV_X1 U21954 ( .A(n20972), .ZN(n21216) );
  XNOR2_X1 U21955 ( .A(n18704), .B(n19637), .ZN(n18705) );
  XNOR2_X1 U21956 ( .A(n18705), .B(n19574), .ZN(n18717) );
  MUX2_X1 U21957 ( .A(n28558), .B(n18707), .S(n18706), .Z(n18711) );
  INV_X1 U21958 ( .A(n18712), .ZN(n18713) );
  XNOR2_X1 U21959 ( .A(n19235), .B(n19232), .ZN(n18715) );
  XNOR2_X1 U21960 ( .A(n19075), .B(n18715), .ZN(n18716) );
  XNOR2_X1 U21961 ( .A(n19215), .B(n3565), .ZN(n18719) );
  XNOR2_X1 U21962 ( .A(n19632), .B(n19085), .ZN(n18718) );
  XNOR2_X1 U21963 ( .A(n18719), .B(n18718), .ZN(n18721) );
  INV_X1 U21964 ( .A(n18749), .ZN(n18751) );
  XNOR2_X1 U21965 ( .A(n19243), .B(n3212), .ZN(n18724) );
  INV_X1 U21966 ( .A(n18722), .ZN(n18723) );
  XNOR2_X1 U21967 ( .A(n18724), .B(n18723), .ZN(n18728) );
  INV_X1 U21968 ( .A(n18725), .ZN(n19226) );
  XNOR2_X1 U21969 ( .A(n18726), .B(n19226), .ZN(n18727) );
  XNOR2_X1 U21970 ( .A(n19525), .B(n19626), .ZN(n18729) );
  XNOR2_X1 U21971 ( .A(n18729), .B(n18730), .ZN(n18734) );
  XNOR2_X1 U21972 ( .A(n18960), .B(n19408), .ZN(n18732) );
  XNOR2_X1 U21973 ( .A(n19096), .B(n26680), .ZN(n18731) );
  XNOR2_X1 U21974 ( .A(n18732), .B(n18731), .ZN(n18733) );
  INV_X1 U21975 ( .A(n19582), .ZN(n18736) );
  XNOR2_X1 U21976 ( .A(n18735), .B(n18863), .ZN(n19203) );
  XNOR2_X1 U21977 ( .A(n18736), .B(n19203), .ZN(n18742) );
  XNOR2_X1 U21978 ( .A(n18760), .B(n3369), .ZN(n18740) );
  INV_X1 U21979 ( .A(n18738), .ZN(n19644) );
  XNOR2_X1 U21980 ( .A(n18737), .B(n19644), .ZN(n18739) );
  XNOR2_X1 U21981 ( .A(n18740), .B(n18739), .ZN(n18741) );
  XNOR2_X1 U21982 ( .A(n19607), .B(n18743), .ZN(n18748) );
  XNOR2_X1 U21983 ( .A(n18744), .B(n3036), .ZN(n18745) );
  XNOR2_X1 U21984 ( .A(n18745), .B(n18746), .ZN(n18747) );
  XNOR2_X1 U21985 ( .A(n18755), .B(n18754), .ZN(n18759) );
  XNOR2_X1 U21986 ( .A(n29318), .B(n3787), .ZN(n18757) );
  XNOR2_X1 U21987 ( .A(n29492), .B(n18942), .ZN(n19681) );
  XNOR2_X1 U21988 ( .A(n18757), .B(n19681), .ZN(n18758) );
  XNOR2_X1 U21989 ( .A(n18759), .B(n18758), .ZN(n20064) );
  XNOR2_X1 U21990 ( .A(n18761), .B(n18760), .ZN(n19438) );
  XNOR2_X1 U21991 ( .A(n19585), .B(n18798), .ZN(n18764) );
  XNOR2_X1 U21992 ( .A(n28798), .B(n3191), .ZN(n18763) );
  INV_X1 U21993 ( .A(n18766), .ZN(n19165) );
  XNOR2_X1 U21995 ( .A(n19165), .B(n18768), .ZN(n18771) );
  XNOR2_X1 U21996 ( .A(n29506), .B(n19704), .ZN(n18770) );
  XNOR2_X1 U21997 ( .A(n18770), .B(n18769), .ZN(n19455) );
  NOR2_X1 U21998 ( .A1(n20063), .A2(n20049), .ZN(n18846) );
  XNOR2_X1 U21999 ( .A(n19306), .B(n19686), .ZN(n18772) );
  XNOR2_X1 U22000 ( .A(n18981), .B(n19687), .ZN(n19420) );
  XNOR2_X1 U22001 ( .A(n18772), .B(n19420), .ZN(n18775) );
  INV_X1 U22002 ( .A(n18773), .ZN(n19110) );
  NOR2_X1 U22003 ( .A1(n20064), .A2(n19761), .ZN(n18776) );
  XNOR2_X1 U22004 ( .A(n19448), .B(n19615), .ZN(n18995) );
  XNOR2_X1 U22005 ( .A(n19313), .B(n5633), .ZN(n18777) );
  XNOR2_X1 U22006 ( .A(n18777), .B(n18995), .ZN(n18781) );
  XNOR2_X1 U22007 ( .A(n18778), .B(n18935), .ZN(n19447) );
  XNOR2_X1 U22008 ( .A(n19447), .B(n18779), .ZN(n18780) );
  XNOR2_X1 U22009 ( .A(n18781), .B(n18780), .ZN(n18845) );
  XNOR2_X1 U22010 ( .A(n19320), .B(n2350), .ZN(n18783) );
  XNOR2_X1 U22011 ( .A(n19697), .B(n18959), .ZN(n18784) );
  XNOR2_X1 U22012 ( .A(n18784), .B(n19692), .ZN(n19436) );
  XNOR2_X1 U22013 ( .A(n18785), .B(n19436), .ZN(n20066) );
  NAND3_X1 U22014 ( .A1(n21221), .A2(n20972), .A3(n20966), .ZN(n18786) );
  INV_X1 U22016 ( .A(n20089), .ZN(n19778) );
  NOR2_X1 U22017 ( .A1(n18790), .A2(n20039), .ZN(n20877) );
  INV_X1 U22018 ( .A(n18791), .ZN(n18793) );
  XNOR2_X1 U22019 ( .A(n19349), .B(n18937), .ZN(n18792) );
  XNOR2_X1 U22020 ( .A(n18793), .B(n18792), .ZN(n18797) );
  XNOR2_X1 U22021 ( .A(n19491), .B(n19228), .ZN(n18795) );
  XNOR2_X1 U22022 ( .A(n18927), .B(n2541), .ZN(n18794) );
  XNOR2_X1 U22023 ( .A(n18795), .B(n18794), .ZN(n18796) );
  XNOR2_X1 U22024 ( .A(n18798), .B(n18799), .ZN(n18801) );
  XNOR2_X1 U22025 ( .A(n18899), .B(n900), .ZN(n18800) );
  XNOR2_X1 U22026 ( .A(n18801), .B(n18800), .ZN(n18805) );
  XNOR2_X1 U22027 ( .A(n18802), .B(n19725), .ZN(n18803) );
  XNOR2_X1 U22028 ( .A(n19546), .B(n18803), .ZN(n18804) );
  INV_X1 U22029 ( .A(n20098), .ZN(n20096) );
  INV_X1 U22030 ( .A(n18806), .ZN(n19696) );
  XNOR2_X1 U22031 ( .A(n19321), .B(n19696), .ZN(n18807) );
  XNOR2_X1 U22032 ( .A(n19528), .B(n18807), .ZN(n18811) );
  XNOR2_X1 U22033 ( .A(n19409), .B(n3029), .ZN(n18809) );
  XNOR2_X1 U22034 ( .A(n19320), .B(n19412), .ZN(n18808) );
  XNOR2_X1 U22035 ( .A(n18809), .B(n18808), .ZN(n18810) );
  XNOR2_X1 U22036 ( .A(n18811), .B(n18810), .ZN(n20150) );
  INV_X1 U22037 ( .A(n18812), .ZN(n19371) );
  XNOR2_X1 U22038 ( .A(n19371), .B(n19300), .ZN(n18814) );
  XNOR2_X1 U22039 ( .A(n19377), .B(n27956), .ZN(n18813) );
  XNOR2_X1 U22040 ( .A(n18814), .B(n18813), .ZN(n18819) );
  XNOR2_X1 U22041 ( .A(n28144), .B(n19679), .ZN(n18817) );
  INV_X1 U22042 ( .A(n18815), .ZN(n18816) );
  XNOR2_X1 U22043 ( .A(n18816), .B(n18817), .ZN(n18818) );
  XNOR2_X1 U22044 ( .A(n18912), .B(n19706), .ZN(n18821) );
  XNOR2_X1 U22045 ( .A(n19700), .B(n2544), .ZN(n18820) );
  XNOR2_X1 U22046 ( .A(n18821), .B(n18820), .ZN(n18823) );
  XNOR2_X1 U22047 ( .A(n18114), .B(n19024), .ZN(n19498) );
  XNOR2_X1 U22048 ( .A(n19498), .B(n19540), .ZN(n18822) );
  XNOR2_X1 U22049 ( .A(n18906), .B(n19219), .ZN(n18826) );
  INV_X1 U22050 ( .A(n18824), .ZN(n18825) );
  XNOR2_X1 U22051 ( .A(n18826), .B(n18825), .ZN(n18830) );
  XNOR2_X1 U22052 ( .A(n19389), .B(n19306), .ZN(n18828) );
  INV_X1 U22053 ( .A(n3537), .ZN(n27324) );
  XNOR2_X1 U22054 ( .A(n19685), .B(n27324), .ZN(n18827) );
  XNOR2_X1 U22055 ( .A(n18828), .B(n18827), .ZN(n18829) );
  XNOR2_X1 U22056 ( .A(n18830), .B(n18829), .ZN(n18887) );
  INV_X1 U22059 ( .A(n18834), .ZN(n20574) );
  NOR2_X1 U22061 ( .A1(n29145), .A2(n18838), .ZN(n18836) );
  NOR2_X1 U22062 ( .A1(n20077), .A2(n28526), .ZN(n18835) );
  INV_X1 U22063 ( .A(n18838), .ZN(n20083) );
  INV_X1 U22064 ( .A(n20375), .ZN(n20371) );
  INV_X1 U22065 ( .A(n19841), .ZN(n20377) );
  MUX2_X1 U22066 ( .A(n19739), .B(n20371), .S(n20377), .Z(n18844) );
  INV_X1 U22067 ( .A(n20373), .ZN(n20074) );
  NOR2_X1 U22068 ( .A1(n20379), .A2(n20074), .ZN(n18841) );
  NOR2_X1 U22069 ( .A1(n19740), .A2(n19841), .ZN(n18840) );
  AOI22_X1 U22070 ( .A1(n18843), .A2(n18841), .B1(n18840), .B2(n20371), .ZN(
        n18842) );
  NOR2_X1 U22071 ( .A1(n21266), .A2(n20816), .ZN(n18849) );
  INV_X1 U22072 ( .A(n18845), .ZN(n20065) );
  INV_X1 U22073 ( .A(n20066), .ZN(n20048) );
  INV_X1 U22074 ( .A(n20063), .ZN(n18892) );
  INV_X1 U22075 ( .A(n18846), .ZN(n19764) );
  NOR2_X1 U22076 ( .A1(n21268), .A2(n20875), .ZN(n21271) );
  AOI22_X1 U22077 ( .A1(n21269), .A2(n18849), .B1(n21271), .B2(n21266), .ZN(
        n18850) );
  XNOR2_X1 U22079 ( .A(n19123), .B(n18852), .ZN(n19575) );
  XNOR2_X1 U22081 ( .A(n19235), .B(n3049), .ZN(n18853) );
  XNOR2_X1 U22082 ( .A(n19125), .B(n18853), .ZN(n18854) );
  XNOR2_X1 U22083 ( .A(n18855), .B(n18854), .ZN(n20158) );
  XNOR2_X1 U22084 ( .A(n19206), .B(n27894), .ZN(n18858) );
  INV_X1 U22086 ( .A(n19096), .ZN(n18859) );
  XNOR2_X1 U22087 ( .A(n19508), .B(n18859), .ZN(n19033) );
  XNOR2_X1 U22088 ( .A(n19116), .B(n19033), .ZN(n18860) );
  XNOR2_X1 U22089 ( .A(n18861), .B(n18860), .ZN(n20159) );
  NAND2_X1 U22090 ( .A1(n20158), .A2(n20159), .ZN(n19874) );
  XNOR2_X1 U22091 ( .A(n19250), .B(n19256), .ZN(n19583) );
  XNOR2_X1 U22092 ( .A(n19583), .B(n18862), .ZN(n18866) );
  XNOR2_X1 U22094 ( .A(n18863), .B(n3154), .ZN(n18864) );
  XNOR2_X1 U22095 ( .A(n19040), .B(n18864), .ZN(n18865) );
  INV_X1 U22096 ( .A(n20161), .ZN(n19984) );
  NAND2_X1 U22097 ( .A1(n19874), .A2(n19984), .ZN(n18886) );
  INV_X1 U22098 ( .A(n18868), .ZN(n18869) );
  XNOR2_X1 U22099 ( .A(n18869), .B(n19599), .ZN(n18873) );
  XNOR2_X1 U22100 ( .A(n19085), .B(n19220), .ZN(n18871) );
  XNOR2_X1 U22101 ( .A(n19481), .B(n3752), .ZN(n18870) );
  XNOR2_X1 U22102 ( .A(n18871), .B(n18870), .ZN(n18872) );
  INV_X1 U22104 ( .A(n20157), .ZN(n20044) );
  XNOR2_X1 U22106 ( .A(n19192), .B(n19103), .ZN(n18876) );
  XNOR2_X1 U22107 ( .A(n19500), .B(n2325), .ZN(n18875) );
  INV_X1 U22108 ( .A(n19604), .ZN(n19281) );
  NAND3_X1 U22109 ( .A1(n19985), .A2(n20158), .A3(n29066), .ZN(n18885) );
  XNOR2_X1 U22110 ( .A(n19243), .B(n3650), .ZN(n18879) );
  XNOR2_X1 U22111 ( .A(n19484), .B(n19225), .ZN(n18878) );
  XNOR2_X1 U22112 ( .A(n18879), .B(n18878), .ZN(n18882) );
  XNOR2_X1 U22113 ( .A(n18880), .B(n19139), .ZN(n19613) );
  XNOR2_X1 U22114 ( .A(n19141), .B(n19613), .ZN(n18881) );
  XNOR2_X1 U22115 ( .A(n18881), .B(n18882), .ZN(n20162) );
  NAND2_X1 U22117 ( .A1(n28187), .A2(n20161), .ZN(n20045) );
  INV_X1 U22118 ( .A(n21288), .ZN(n20916) );
  INV_X1 U22119 ( .A(n18887), .ZN(n20151) );
  NOR2_X1 U22121 ( .A1(n18888), .A2(n28188), .ZN(n18889) );
  NAND2_X1 U22122 ( .A1(n20916), .A2(n20988), .ZN(n21286) );
  OAI21_X1 U22123 ( .B1(n18765), .B2(n19761), .A(n20066), .ZN(n18891) );
  XNOR2_X1 U22124 ( .A(n19462), .B(n19378), .ZN(n18893) );
  XNOR2_X1 U22125 ( .A(n18894), .B(n18893), .ZN(n18898) );
  XNOR2_X1 U22126 ( .A(n19299), .B(n19377), .ZN(n18896) );
  XNOR2_X1 U22127 ( .A(n19427), .B(n3180), .ZN(n18895) );
  XNOR2_X1 U22128 ( .A(n18896), .B(n18895), .ZN(n18897) );
  XNOR2_X2 U22129 ( .A(n18898), .B(n18897), .ZN(n18919) );
  XNOR2_X1 U22130 ( .A(n19251), .B(n19256), .ZN(n18901) );
  XNOR2_X1 U22131 ( .A(n18899), .B(n18900), .ZN(n19381) );
  XNOR2_X1 U22132 ( .A(n18901), .B(n19381), .ZN(n18905) );
  XNOR2_X1 U22133 ( .A(n19198), .B(n19727), .ZN(n18903) );
  XNOR2_X1 U22134 ( .A(n19643), .B(n27105), .ZN(n18902) );
  XNOR2_X1 U22135 ( .A(n18903), .B(n18902), .ZN(n18904) );
  XNOR2_X1 U22136 ( .A(n19086), .B(n19045), .ZN(n19635) );
  INV_X1 U22137 ( .A(n19635), .ZN(n18907) );
  XNOR2_X1 U22138 ( .A(n19421), .B(n19482), .ZN(n19153) );
  XNOR2_X1 U22139 ( .A(n18907), .B(n19153), .ZN(n18911) );
  INV_X1 U22140 ( .A(n19084), .ZN(n18909) );
  XNOR2_X1 U22141 ( .A(n19108), .B(n21537), .ZN(n18908) );
  XNOR2_X1 U22142 ( .A(n18909), .B(n18908), .ZN(n18910) );
  MUX2_X1 U22143 ( .A(n18919), .B(n21091), .S(n20144), .Z(n18918) );
  XNOR2_X1 U22144 ( .A(n18912), .B(n19025), .ZN(n19651) );
  XNOR2_X1 U22145 ( .A(n19496), .B(n19702), .ZN(n19164) );
  XNOR2_X1 U22146 ( .A(n19651), .B(n19164), .ZN(n18917) );
  INV_X1 U22147 ( .A(n19105), .ZN(n18915) );
  XNOR2_X1 U22148 ( .A(n18913), .B(n3635), .ZN(n18914) );
  XNOR2_X1 U22149 ( .A(n18915), .B(n18914), .ZN(n18916) );
  NOR2_X1 U22150 ( .A1(n18918), .A2(n20145), .ZN(n19011) );
  INV_X1 U22151 ( .A(n19011), .ZN(n18932) );
  XNOR2_X1 U22152 ( .A(n19691), .B(n19511), .ZN(n18921) );
  INV_X1 U22153 ( .A(n19095), .ZN(n18920) );
  XNOR2_X1 U22154 ( .A(n18920), .B(n18921), .ZN(n18926) );
  XNOR2_X1 U22155 ( .A(n19413), .B(n18922), .ZN(n18924) );
  XNOR2_X1 U22156 ( .A(n19412), .B(n3697), .ZN(n18923) );
  XNOR2_X1 U22157 ( .A(n18924), .B(n18923), .ZN(n18925) );
  INV_X1 U22158 ( .A(n18928), .ZN(n19520) );
  XNOR2_X1 U22159 ( .A(n19487), .B(n19229), .ZN(n19181) );
  NOR2_X1 U22160 ( .A1(n20102), .A2(n21091), .ZN(n18930) );
  AOI22_X1 U22161 ( .A1(n19010), .A2(n21091), .B1(n18930), .B2(n20145), .ZN(
        n18931) );
  NAND2_X1 U22162 ( .A1(n18932), .A2(n18931), .ZN(n18934) );
  INV_X1 U22163 ( .A(n18934), .ZN(n19014) );
  INV_X1 U22164 ( .A(n21291), .ZN(n21289) );
  XNOR2_X1 U22165 ( .A(n19669), .B(n29038), .ZN(n18936) );
  XNOR2_X1 U22166 ( .A(n19519), .B(n18936), .ZN(n18941) );
  XNOR2_X1 U22167 ( .A(n19228), .B(n18937), .ZN(n18939) );
  XNOR2_X1 U22168 ( .A(n19246), .B(n3256), .ZN(n18938) );
  XNOR2_X1 U22169 ( .A(n18939), .B(n18938), .ZN(n18940) );
  XNOR2_X1 U22170 ( .A(n18941), .B(n18940), .ZN(n20165) );
  XNOR2_X1 U22171 ( .A(n28143), .B(n19637), .ZN(n18945) );
  XNOR2_X1 U22172 ( .A(n18942), .B(n3491), .ZN(n18943) );
  XNOR2_X1 U22173 ( .A(n18943), .B(n19679), .ZN(n18944) );
  XNOR2_X1 U22174 ( .A(n18944), .B(n18945), .ZN(n18947) );
  XNOR2_X1 U22176 ( .A(n19557), .B(n29484), .ZN(n18946) );
  XNOR2_X1 U22177 ( .A(n18946), .B(n18947), .ZN(n18972) );
  XNOR2_X1 U22178 ( .A(n19144), .B(n19548), .ZN(n18953) );
  XNOR2_X1 U22179 ( .A(n19725), .B(n19644), .ZN(n18951) );
  XNOR2_X1 U22180 ( .A(n18949), .B(n2389), .ZN(n18950) );
  XNOR2_X1 U22181 ( .A(n18951), .B(n18950), .ZN(n18952) );
  AOI21_X1 U22182 ( .B1(n18972), .B2(n20165), .A(n20166), .ZN(n18974) );
  XNOR2_X1 U22183 ( .A(n29506), .B(n2602), .ZN(n18954) );
  XNOR2_X1 U22184 ( .A(n18955), .B(n18954), .ZN(n18957) );
  XNOR2_X1 U22185 ( .A(n19191), .B(n19403), .ZN(n19132) );
  XNOR2_X1 U22186 ( .A(n19132), .B(n19541), .ZN(n18956) );
  XNOR2_X1 U22187 ( .A(n18956), .B(n18957), .ZN(n19993) );
  INV_X1 U22189 ( .A(n19626), .ZN(n18958) );
  XNOR2_X1 U22190 ( .A(n18958), .B(n19408), .ZN(n18961) );
  XNOR2_X1 U22191 ( .A(n18960), .B(n18959), .ZN(n19526) );
  XNOR2_X1 U22192 ( .A(n19526), .B(n18961), .ZN(n18965) );
  XNOR2_X1 U22193 ( .A(n19696), .B(n19697), .ZN(n18963) );
  XNOR2_X1 U22194 ( .A(n19207), .B(n3003), .ZN(n18962) );
  XNOR2_X1 U22195 ( .A(n18963), .B(n18962), .ZN(n18964) );
  MUX2_X1 U22196 ( .A(n29587), .B(n297), .S(n19989), .Z(n18973) );
  INV_X1 U22197 ( .A(n18966), .ZN(n19533) );
  XNOR2_X1 U22198 ( .A(n19533), .B(n18967), .ZN(n18971) );
  XNOR2_X1 U22199 ( .A(n19272), .B(n19632), .ZN(n18969) );
  XNOR2_X1 U22200 ( .A(n19685), .B(n3276), .ZN(n18968) );
  XNOR2_X1 U22201 ( .A(n18969), .B(n18968), .ZN(n18970) );
  INV_X1 U22202 ( .A(n21290), .ZN(n20986) );
  INV_X1 U22203 ( .A(n19331), .ZN(n18976) );
  INV_X1 U22204 ( .A(n18975), .ZN(n19625) );
  XNOR2_X1 U22205 ( .A(n18976), .B(n19625), .ZN(n19094) );
  XNOR2_X1 U22206 ( .A(n19094), .B(n19330), .ZN(n18979) );
  XNOR2_X1 U22207 ( .A(n19525), .B(n19507), .ZN(n19212) );
  XNOR2_X1 U22208 ( .A(n19212), .B(n18977), .ZN(n18978) );
  XNOR2_X1 U22209 ( .A(n18979), .B(n18978), .ZN(n19054) );
  XNOR2_X1 U22210 ( .A(n18981), .B(n18980), .ZN(n18983) );
  XNOR2_X1 U22211 ( .A(n19483), .B(n3457), .ZN(n18982) );
  XNOR2_X1 U22212 ( .A(n18983), .B(n18982), .ZN(n18986) );
  XNOR2_X1 U22213 ( .A(n19631), .B(n19110), .ZN(n19082) );
  XNOR2_X1 U22214 ( .A(n19082), .B(n18984), .ZN(n18985) );
  XNOR2_X1 U22215 ( .A(n19549), .B(n3501), .ZN(n18990) );
  XNOR2_X1 U22217 ( .A(n29554), .B(n19397), .ZN(n18992) );
  XNOR2_X1 U22219 ( .A(n19617), .B(n2306), .ZN(n18994) );
  XNOR2_X1 U22220 ( .A(n18995), .B(n18994), .ZN(n18996) );
  XNOR2_X1 U22221 ( .A(n18997), .B(n18996), .ZN(n20053) );
  INV_X1 U22222 ( .A(n19333), .ZN(n18998) );
  XNOR2_X1 U22223 ( .A(n29318), .B(n19376), .ZN(n19079) );
  XNOR2_X1 U22224 ( .A(n19428), .B(n3742), .ZN(n18999) );
  XNOR2_X1 U22225 ( .A(n19079), .B(n18999), .ZN(n19000) );
  XNOR2_X1 U22226 ( .A(n19000), .B(n19001), .ZN(n20178) );
  OAI21_X1 U22229 ( .B1(n20174), .B2(n4886), .A(n19002), .ZN(n19008) );
  XNOR2_X1 U22230 ( .A(n28516), .B(n19603), .ZN(n19101) );
  XNOR2_X1 U22231 ( .A(n19495), .B(n19356), .ZN(n19005) );
  XNOR2_X1 U22232 ( .A(n19006), .B(n19005), .ZN(n20176) );
  INV_X1 U22233 ( .A(n19052), .ZN(n19007) );
  NOR2_X1 U22234 ( .A1(n21291), .A2(n21287), .ZN(n19013) );
  XNOR2_X1 U22235 ( .A(n22582), .B(n21884), .ZN(n19738) );
  XNOR2_X1 U22236 ( .A(n19371), .B(n19378), .ZN(n19015) );
  XNOR2_X1 U22237 ( .A(n19313), .B(n24906), .ZN(n19019) );
  XNOR2_X1 U22238 ( .A(n19020), .B(n19019), .ZN(n19023) );
  XNOR2_X1 U22239 ( .A(n19484), .B(n19487), .ZN(n19021) );
  XNOR2_X1 U22240 ( .A(n19399), .B(n19021), .ZN(n19022) );
  XNOR2_X1 U22241 ( .A(n19023), .B(n19022), .ZN(n20479) );
  XNOR2_X1 U22242 ( .A(n19496), .B(n19024), .ZN(n19027) );
  XNOR2_X1 U22243 ( .A(n19027), .B(n19026), .ZN(n19031) );
  XNOR2_X1 U22244 ( .A(n19700), .B(n2446), .ZN(n19029) );
  XNOR2_X1 U22245 ( .A(n19500), .B(n19452), .ZN(n19028) );
  XNOR2_X1 U22246 ( .A(n19029), .B(n19028), .ZN(n19030) );
  XNOR2_X1 U22247 ( .A(n19409), .B(n19511), .ZN(n19034) );
  XNOR2_X1 U22248 ( .A(n19033), .B(n19034), .ZN(n19038) );
  XNOR2_X1 U22249 ( .A(n19413), .B(n3770), .ZN(n19035) );
  XNOR2_X1 U22250 ( .A(n19036), .B(n19035), .ZN(n19037) );
  INV_X1 U22251 ( .A(n19039), .ZN(n19382) );
  XNOR2_X1 U22252 ( .A(n19382), .B(n19040), .ZN(n19044) );
  INV_X1 U22253 ( .A(n1184), .ZN(n19041) );
  XNOR2_X1 U22254 ( .A(n19440), .B(n19041), .ZN(n19042) );
  XNOR2_X1 U22255 ( .A(n19472), .B(n19042), .ZN(n19043) );
  XNOR2_X1 U22256 ( .A(n19044), .B(n19043), .ZN(n19995) );
  XNOR2_X1 U22257 ( .A(n19423), .B(n19085), .ZN(n19047) );
  XNOR2_X1 U22258 ( .A(n19045), .B(n19481), .ZN(n19046) );
  XNOR2_X1 U22259 ( .A(n19047), .B(n19046), .ZN(n19051) );
  XNOR2_X1 U22260 ( .A(n19482), .B(n19306), .ZN(n19049) );
  XNOR2_X1 U22261 ( .A(n19049), .B(n19048), .ZN(n19050) );
  INV_X1 U22262 ( .A(n19054), .ZN(n19976) );
  OAI21_X1 U22263 ( .B1(n19055), .B2(n19976), .A(n20171), .ZN(n19056) );
  INV_X1 U22264 ( .A(n21277), .ZN(n21278) );
  NOR2_X1 U22265 ( .A1(n297), .A2(n20219), .ZN(n19059) );
  NOR3_X1 U22266 ( .A1(n19860), .A2(n19059), .A3(n20222), .ZN(n19063) );
  NAND3_X1 U22267 ( .A1(n19989), .A2(n385), .A3(n296), .ZN(n19061) );
  NAND2_X1 U22268 ( .A1(n21278), .A2(n21703), .ZN(n21378) );
  XNOR2_X1 U22269 ( .A(n19615), .B(n2381), .ZN(n19064) );
  XNOR2_X1 U22270 ( .A(n19665), .B(n19064), .ZN(n19068) );
  XNOR2_X1 U22271 ( .A(n19066), .B(n19065), .ZN(n19067) );
  XNOR2_X1 U22272 ( .A(n19251), .B(n19727), .ZN(n19070) );
  XNOR2_X1 U22273 ( .A(n19584), .B(n2912), .ZN(n19069) );
  XNOR2_X1 U22274 ( .A(n19070), .B(n19069), .ZN(n19074) );
  INV_X1 U22275 ( .A(n19071), .ZN(n19072) );
  XNOR2_X1 U22276 ( .A(n19646), .B(n19072), .ZN(n19073) );
  INV_X1 U22277 ( .A(n19093), .ZN(n20486) );
  NOR2_X1 U22278 ( .A1(n20481), .A2(n20486), .ZN(n20238) );
  XNOR2_X1 U22279 ( .A(n19075), .B(n3451), .ZN(n19076) );
  XNOR2_X1 U22280 ( .A(n19077), .B(n19076), .ZN(n19081) );
  XNOR2_X1 U22281 ( .A(n19079), .B(n19078), .ZN(n19080) );
  INV_X1 U22282 ( .A(n19082), .ZN(n19083) );
  XNOR2_X1 U22283 ( .A(n19083), .B(n19084), .ZN(n19091) );
  XNOR2_X1 U22284 ( .A(n19086), .B(n19085), .ZN(n19089) );
  XNOR2_X1 U22285 ( .A(n19087), .B(n26909), .ZN(n19088) );
  XNOR2_X1 U22286 ( .A(n19089), .B(n19088), .ZN(n19090) );
  INV_X1 U22287 ( .A(n20483), .ZN(n20000) );
  XNOR2_X1 U22288 ( .A(n19094), .B(n19095), .ZN(n19100) );
  XNOR2_X1 U22289 ( .A(n19096), .B(n2894), .ZN(n19098) );
  XNOR2_X1 U22290 ( .A(n19098), .B(n19097), .ZN(n19099) );
  XNOR2_X1 U22291 ( .A(n19101), .B(n19102), .ZN(n19107) );
  XNOR2_X1 U22292 ( .A(n19103), .B(n730), .ZN(n19104) );
  XNOR2_X1 U22293 ( .A(n19105), .B(n19104), .ZN(n19106) );
  NOR2_X1 U22294 ( .A1(n20488), .A2(n20239), .ZN(n20482) );
  XNOR2_X1 U22295 ( .A(n19272), .B(n19688), .ZN(n19388) );
  XNOR2_X1 U22296 ( .A(n19219), .B(n19108), .ZN(n19109) );
  XNOR2_X1 U22297 ( .A(n19109), .B(n19388), .ZN(n19115) );
  XNOR2_X1 U22298 ( .A(n19110), .B(n3081), .ZN(n19113) );
  XNOR2_X1 U22299 ( .A(n19113), .B(n19112), .ZN(n19114) );
  XNOR2_X1 U22300 ( .A(n19115), .B(n19114), .ZN(n20499) );
  INV_X1 U22301 ( .A(n20499), .ZN(n20227) );
  XNOR2_X1 U22302 ( .A(n19116), .B(n19117), .ZN(n19121) );
  XNOR2_X1 U22303 ( .A(n19207), .B(n24959), .ZN(n19118) );
  XNOR2_X1 U22304 ( .A(n19119), .B(n19118), .ZN(n19120) );
  XNOR2_X1 U22306 ( .A(n28144), .B(n19373), .ZN(n19124) );
  XNOR2_X1 U22307 ( .A(n29318), .B(n3662), .ZN(n19126) );
  XNOR2_X1 U22308 ( .A(n19125), .B(n19126), .ZN(n19127) );
  MUX2_X1 U22310 ( .A(n20227), .B(n28621), .S(n20500), .Z(n19151) );
  INV_X1 U22311 ( .A(n19130), .ZN(n19131) );
  XNOR2_X1 U22312 ( .A(n19603), .B(n2402), .ZN(n19134) );
  XNOR2_X1 U22313 ( .A(n19133), .B(n19134), .ZN(n19135) );
  XNOR2_X1 U22314 ( .A(n19616), .B(n19228), .ZN(n19138) );
  XNOR2_X1 U22315 ( .A(n19136), .B(n2411), .ZN(n19137) );
  XNOR2_X1 U22316 ( .A(n19138), .B(n19137), .ZN(n19143) );
  XNOR2_X1 U22317 ( .A(n19139), .B(n19615), .ZN(n19140) );
  XNOR2_X1 U22318 ( .A(n19141), .B(n19140), .ZN(n19142) );
  XNOR2_X1 U22319 ( .A(n18395), .B(n19359), .ZN(n19145) );
  XNOR2_X1 U22320 ( .A(n19256), .B(n19726), .ZN(n19147) );
  XNOR2_X1 U22321 ( .A(n19584), .B(n2404), .ZN(n19146) );
  XNOR2_X1 U22322 ( .A(n19147), .B(n19146), .ZN(n19148) );
  NOR2_X1 U22323 ( .A1(n20500), .A2(n20339), .ZN(n19149) );
  AOI21_X2 U22324 ( .B1(n19151), .B2(n19150), .A(n19149), .ZN(n21704) );
  XNOR2_X1 U22325 ( .A(n19687), .B(n19305), .ZN(n19152) );
  INV_X1 U22326 ( .A(n3380), .ZN(n27811) );
  XNOR2_X1 U22327 ( .A(n19370), .B(n2946), .ZN(n19155) );
  XNOR2_X1 U22328 ( .A(n19155), .B(n19234), .ZN(n19158) );
  XNOR2_X1 U22329 ( .A(n19156), .B(n19296), .ZN(n19157) );
  INV_X1 U22330 ( .A(n20493), .ZN(n20179) );
  XNOR2_X1 U22331 ( .A(n18760), .B(n28798), .ZN(n19161) );
  XNOR2_X1 U22332 ( .A(n19198), .B(n2981), .ZN(n19160) );
  XNOR2_X1 U22333 ( .A(n19161), .B(n19160), .ZN(n19163) );
  XNOR2_X1 U22334 ( .A(n19164), .B(n19165), .ZN(n19169) );
  XNOR2_X1 U22335 ( .A(n19166), .B(n19706), .ZN(n19167) );
  XNOR2_X1 U22336 ( .A(n19691), .B(n19321), .ZN(n19171) );
  XNOR2_X1 U22337 ( .A(n19696), .B(n19511), .ZN(n19170) );
  XNOR2_X1 U22338 ( .A(n19171), .B(n19170), .ZN(n19178) );
  INV_X1 U22339 ( .A(n19173), .ZN(n19172) );
  NAND2_X1 U22340 ( .A1(n19172), .A2(n5490), .ZN(n19174) );
  INV_X1 U22341 ( .A(Key[26]), .ZN(n24166) );
  XNOR2_X1 U22342 ( .A(n19176), .B(n19175), .ZN(n19177) );
  INV_X1 U22343 ( .A(n20496), .ZN(n19863) );
  XNOR2_X1 U22344 ( .A(n19180), .B(n19348), .ZN(n19182) );
  XNOR2_X1 U22345 ( .A(n19182), .B(n19181), .ZN(n19184) );
  XNOR2_X1 U22346 ( .A(n19184), .B(n19183), .ZN(n20182) );
  MUX2_X1 U22348 ( .A(n19187), .B(n21374), .S(n21372), .Z(n19188) );
  XNOR2_X1 U22351 ( .A(n19191), .B(n19702), .ZN(n19193) );
  XNOR2_X1 U22352 ( .A(n19194), .B(n19277), .ZN(n19195) );
  XNOR2_X1 U22353 ( .A(n19495), .B(n19195), .ZN(n19196) );
  XNOR2_X1 U22354 ( .A(n19197), .B(n19196), .ZN(n20017) );
  XNOR2_X1 U22355 ( .A(n19199), .B(n19198), .ZN(n19201) );
  XNOR2_X1 U22356 ( .A(n19549), .B(n2505), .ZN(n19200) );
  XNOR2_X1 U22357 ( .A(n19201), .B(n19200), .ZN(n19205) );
  XNOR2_X1 U22358 ( .A(n28798), .B(n19474), .ZN(n19202) );
  XNOR2_X1 U22359 ( .A(n19202), .B(n19203), .ZN(n19204) );
  XNOR2_X1 U22360 ( .A(n19206), .B(n19332), .ZN(n19209) );
  XNOR2_X1 U22361 ( .A(n19207), .B(n3586), .ZN(n19208) );
  XNOR2_X1 U22362 ( .A(n19209), .B(n19208), .ZN(n19214) );
  INV_X1 U22365 ( .A(n19215), .ZN(n19216) );
  XNOR2_X1 U22366 ( .A(n19216), .B(n19483), .ZN(n19218) );
  XNOR2_X1 U22367 ( .A(n19339), .B(n2527), .ZN(n19217) );
  XNOR2_X1 U22368 ( .A(n19218), .B(n19217), .ZN(n19224) );
  XNOR2_X1 U22369 ( .A(n19534), .B(n19219), .ZN(n19222) );
  XNOR2_X1 U22370 ( .A(n19421), .B(n19220), .ZN(n19221) );
  XNOR2_X1 U22371 ( .A(n19222), .B(n19221), .ZN(n19223) );
  XNOR2_X1 U22373 ( .A(n19348), .B(n19226), .ZN(n19227) );
  XNOR2_X1 U22374 ( .A(n19670), .B(n19228), .ZN(n19230) );
  XNOR2_X1 U22375 ( .A(n19230), .B(n19229), .ZN(n19231) );
  INV_X1 U22376 ( .A(n20342), .ZN(n20509) );
  XNOR2_X1 U22377 ( .A(n19232), .B(n1919), .ZN(n19233) );
  XNOR2_X1 U22378 ( .A(n19234), .B(n19233), .ZN(n19239) );
  XNOR2_X1 U22379 ( .A(n28143), .B(n19235), .ZN(n19237) );
  XNOR2_X1 U22380 ( .A(n19236), .B(n19237), .ZN(n19238) );
  OAI21_X1 U22381 ( .B1(n20509), .B2(n20510), .A(n20343), .ZN(n19240) );
  XNOR2_X1 U22383 ( .A(n19670), .B(n3462), .ZN(n19242) );
  XNOR2_X1 U22384 ( .A(n19242), .B(n19243), .ZN(n19244) );
  XNOR2_X1 U22385 ( .A(n19244), .B(n19613), .ZN(n19249) );
  XNOR2_X1 U22386 ( .A(n19245), .B(n19246), .ZN(n19247) );
  XNOR2_X1 U22387 ( .A(n19249), .B(n19248), .ZN(n20458) );
  INV_X1 U22388 ( .A(n20458), .ZN(n20028) );
  XNOR2_X1 U22389 ( .A(n19250), .B(n19251), .ZN(n19254) );
  XNOR2_X1 U22391 ( .A(n19256), .B(n28798), .ZN(n19258) );
  XNOR2_X1 U22392 ( .A(n19474), .B(n26214), .ZN(n19257) );
  XNOR2_X1 U22393 ( .A(n19258), .B(n19257), .ZN(n19259) );
  XNOR2_X1 U22394 ( .A(n19462), .B(n29484), .ZN(n19261) );
  XNOR2_X1 U22395 ( .A(n19575), .B(n19261), .ZN(n19264) );
  XNOR2_X1 U22396 ( .A(n19262), .B(n2961), .ZN(n19263) );
  INV_X1 U22397 ( .A(n19628), .ZN(n19266) );
  XNOR2_X1 U22398 ( .A(n19408), .B(n19332), .ZN(n19265) );
  XNOR2_X1 U22400 ( .A(n19267), .B(n1123), .ZN(n19268) );
  XNOR2_X1 U22401 ( .A(n19269), .B(n19268), .ZN(n19270) );
  XNOR2_X1 U22402 ( .A(n19272), .B(n19273), .ZN(n19275) );
  XNOR2_X1 U22403 ( .A(n19339), .B(n3372), .ZN(n19274) );
  XNOR2_X1 U22404 ( .A(n19275), .B(n19274), .ZN(n19276) );
  XNOR2_X1 U22405 ( .A(n19277), .B(n28294), .ZN(n19280) );
  XNOR2_X1 U22406 ( .A(n19278), .B(n19403), .ZN(n19279) );
  INV_X1 U22407 ( .A(n19283), .ZN(n19701) );
  XNOR2_X1 U22408 ( .A(n19701), .B(n3323), .ZN(n19284) );
  XNOR2_X1 U22409 ( .A(n19284), .B(n19285), .ZN(n19288) );
  XNOR2_X1 U22410 ( .A(n28516), .B(n18638), .ZN(n19286) );
  XNOR2_X1 U22411 ( .A(n19498), .B(n19286), .ZN(n19287) );
  XNOR2_X1 U22414 ( .A(n19291), .B(n28571), .ZN(n19293) );
  XNOR2_X1 U22415 ( .A(n19475), .B(n3134), .ZN(n19292) );
  XNOR2_X1 U22416 ( .A(n19293), .B(n19292), .ZN(n19294) );
  XNOR2_X2 U22417 ( .A(n19295), .B(n19294), .ZN(n20334) );
  INV_X1 U22418 ( .A(n19296), .ZN(n19297) );
  XNOR2_X1 U22419 ( .A(n19297), .B(n19298), .ZN(n19304) );
  XNOR2_X1 U22420 ( .A(n19299), .B(n19300), .ZN(n19302) );
  XNOR2_X1 U22421 ( .A(n19376), .B(n2477), .ZN(n19301) );
  XNOR2_X1 U22422 ( .A(n19302), .B(n19301), .ZN(n19303) );
  XNOR2_X2 U22423 ( .A(n19304), .B(n19303), .ZN(n20623) );
  XNOR2_X1 U22424 ( .A(n19631), .B(n19481), .ZN(n19307) );
  XNOR2_X1 U22425 ( .A(n19308), .B(n19307), .ZN(n19312) );
  XNOR2_X1 U22426 ( .A(n19595), .B(n19535), .ZN(n19310) );
  XNOR2_X1 U22427 ( .A(n19685), .B(n3482), .ZN(n19309) );
  XNOR2_X1 U22428 ( .A(n19310), .B(n19309), .ZN(n19311) );
  XNOR2_X1 U22430 ( .A(n6489), .B(n19397), .ZN(n19314) );
  XNOR2_X1 U22431 ( .A(n19520), .B(n3015), .ZN(n19316) );
  XNOR2_X1 U22432 ( .A(n19317), .B(n19316), .ZN(n19318) );
  INV_X1 U22433 ( .A(n20630), .ZN(n20335) );
  XNOR2_X1 U22434 ( .A(n19592), .B(n19323), .ZN(n19529) );
  XNOR2_X1 U22435 ( .A(n19625), .B(n3710), .ZN(n19324) );
  XNOR2_X1 U22436 ( .A(n19529), .B(n19324), .ZN(n19325) );
  NAND2_X1 U22438 ( .A1(n20625), .A2(n20623), .ZN(n19327) );
  MUX2_X1 U22439 ( .A(n19328), .B(n19327), .S(n20005), .Z(n19329) );
  OAI21_X1 U22440 ( .B1(n21364), .B2(n21713), .A(n21714), .ZN(n19461) );
  INV_X1 U22441 ( .A(n21364), .ZN(n21258) );
  XNOR2_X1 U22442 ( .A(n19331), .B(n19626), .ZN(n19591) );
  XNOR2_X1 U22443 ( .A(n19333), .B(n28530), .ZN(n19335) );
  XNOR2_X1 U22444 ( .A(n19568), .B(n3422), .ZN(n19334) );
  XNOR2_X1 U22445 ( .A(n19335), .B(n19334), .ZN(n19337) );
  XNOR2_X2 U22446 ( .A(n19337), .B(n19336), .ZN(n20617) );
  INV_X1 U22447 ( .A(n19339), .ZN(n19340) );
  XNOR2_X1 U22448 ( .A(n19423), .B(n19340), .ZN(n19342) );
  XNOR2_X1 U22449 ( .A(n19342), .B(n19341), .ZN(n19343) );
  XNOR2_X1 U22450 ( .A(n19343), .B(n19344), .ZN(n20431) );
  NOR2_X1 U22451 ( .A1(n20617), .A2(n29040), .ZN(n19345) );
  XNOR2_X1 U22452 ( .A(n19346), .B(n19669), .ZN(n19347) );
  XNOR2_X1 U22453 ( .A(n19348), .B(n19615), .ZN(n19351) );
  XNOR2_X1 U22454 ( .A(n19349), .B(n3508), .ZN(n19350) );
  XNOR2_X1 U22455 ( .A(n19350), .B(n19351), .ZN(n19352) );
  XNOR2_X1 U22456 ( .A(n19452), .B(n135), .ZN(n19355) );
  INV_X1 U22458 ( .A(n20616), .ZN(n20433) );
  XNOR2_X1 U22459 ( .A(n19359), .B(n19440), .ZN(n19361) );
  XNOR2_X1 U22460 ( .A(n29124), .B(n19361), .ZN(n19366) );
  XNOR2_X1 U22461 ( .A(n19584), .B(n2523), .ZN(n19364) );
  INV_X1 U22462 ( .A(n19362), .ZN(n19363) );
  XNOR2_X1 U22463 ( .A(n19364), .B(n19363), .ZN(n19365) );
  OAI21_X1 U22464 ( .B1(n20255), .B2(n20433), .A(n28894), .ZN(n19368) );
  NOR2_X1 U22465 ( .A1(n19920), .A2(n20617), .ZN(n19367) );
  AOI21_X2 U22466 ( .B1(n19369), .B2(n19368), .A(n19367), .ZN(n21366) );
  INV_X1 U22467 ( .A(n21366), .ZN(n21712) );
  AOI21_X1 U22468 ( .B1(n21712), .B2(n5772), .A(n21714), .ZN(n19419) );
  XNOR2_X1 U22469 ( .A(n19370), .B(n27452), .ZN(n19372) );
  XNOR2_X1 U22470 ( .A(n19372), .B(n19371), .ZN(n19375) );
  XNOR2_X1 U22471 ( .A(n19464), .B(n19373), .ZN(n19374) );
  XNOR2_X1 U22472 ( .A(n19375), .B(n19374), .ZN(n19380) );
  XNOR2_X1 U22473 ( .A(n19377), .B(n19376), .ZN(n19379) );
  XNOR2_X1 U22475 ( .A(n19380), .B(n19641), .ZN(n20033) );
  INV_X1 U22476 ( .A(n20033), .ZN(n20247) );
  XNOR2_X1 U22477 ( .A(n19726), .B(n19383), .ZN(n19386) );
  XNOR2_X1 U22478 ( .A(n19384), .B(n3067), .ZN(n19385) );
  XNOR2_X1 U22479 ( .A(n19386), .B(n19385), .ZN(n19387) );
  XNOR2_X1 U22480 ( .A(n19388), .B(n19635), .ZN(n19393) );
  XNOR2_X1 U22481 ( .A(n19389), .B(n2476), .ZN(n19390) );
  XNOR2_X1 U22482 ( .A(n19391), .B(n19390), .ZN(n19392) );
  XNOR2_X1 U22483 ( .A(n19393), .B(n19392), .ZN(n20453) );
  NOR2_X1 U22484 ( .A1(n20641), .A2(n20453), .ZN(n20689) );
  INV_X1 U22485 ( .A(n20689), .ZN(n19394) );
  NAND2_X1 U22486 ( .A1(n21364), .A2(n19394), .ZN(n19417) );
  XNOR2_X1 U22487 ( .A(n18927), .B(n2987), .ZN(n19396) );
  XNOR2_X1 U22488 ( .A(n19486), .B(n19616), .ZN(n19395) );
  XNOR2_X1 U22489 ( .A(n19396), .B(n19395), .ZN(n19401) );
  XNOR2_X1 U22490 ( .A(n19487), .B(n19397), .ZN(n19398) );
  XNOR2_X1 U22491 ( .A(n19399), .B(n19398), .ZN(n19400) );
  XNOR2_X1 U22492 ( .A(n19402), .B(n19651), .ZN(n19407) );
  XNOR2_X1 U22493 ( .A(n19403), .B(n19709), .ZN(n19405) );
  XNOR2_X1 U22494 ( .A(n19700), .B(n3463), .ZN(n19404) );
  XNOR2_X1 U22495 ( .A(n19405), .B(n19404), .ZN(n19406) );
  XNOR2_X1 U22496 ( .A(n19407), .B(n19406), .ZN(n19787) );
  XNOR2_X1 U22497 ( .A(n19409), .B(n19408), .ZN(n19411) );
  XNOR2_X1 U22498 ( .A(n19410), .B(n19411), .ZN(n19416) );
  XNOR2_X1 U22499 ( .A(n19695), .B(n27231), .ZN(n19414) );
  XNOR2_X1 U22500 ( .A(n19624), .B(n19414), .ZN(n19415) );
  INV_X1 U22501 ( .A(n20455), .ZN(n20639) );
  NOR2_X1 U22502 ( .A1(n21716), .A2(n21258), .ZN(n19460) );
  XNOR2_X1 U22503 ( .A(n19421), .B(n19686), .ZN(n19422) );
  XNOR2_X1 U22504 ( .A(n19632), .B(n1172), .ZN(n19425) );
  XNOR2_X1 U22505 ( .A(n19423), .B(n19481), .ZN(n19424) );
  XNOR2_X1 U22507 ( .A(n19428), .B(n19427), .ZN(n19429) );
  XNOR2_X1 U22508 ( .A(n19430), .B(n19429), .ZN(n19431) );
  XNOR2_X1 U22510 ( .A(n19433), .B(n19691), .ZN(n19435) );
  XNOR2_X1 U22511 ( .A(n19508), .B(n19626), .ZN(n19434) );
  XNOR2_X1 U22512 ( .A(n19435), .B(n19434), .ZN(n19437) );
  INV_X1 U22515 ( .A(n19438), .ZN(n19724) );
  XNOR2_X1 U22516 ( .A(n19724), .B(n19439), .ZN(n19444) );
  XNOR2_X1 U22517 ( .A(n19440), .B(n19644), .ZN(n19442) );
  XNOR2_X1 U22518 ( .A(n19475), .B(n2509), .ZN(n19441) );
  XNOR2_X1 U22519 ( .A(n19442), .B(n19441), .ZN(n19443) );
  XNOR2_X1 U22520 ( .A(n19484), .B(n19669), .ZN(n19446) );
  XNOR2_X1 U22521 ( .A(n19445), .B(n19446), .ZN(n19451) );
  INV_X1 U22522 ( .A(n19447), .ZN(n19714) );
  XNOR2_X1 U22523 ( .A(n19448), .B(n1215), .ZN(n19449) );
  XNOR2_X1 U22524 ( .A(n19714), .B(n19449), .ZN(n19450) );
  XNOR2_X1 U22525 ( .A(n19450), .B(n19451), .ZN(n20020) );
  INV_X1 U22526 ( .A(n20020), .ZN(n20520) );
  NOR2_X1 U22527 ( .A1(n20261), .A2(n20520), .ZN(n21360) );
  XNOR2_X1 U22528 ( .A(n19452), .B(n28623), .ZN(n19453) );
  XNOR2_X1 U22529 ( .A(n19454), .B(n19453), .ZN(n19456) );
  MUX2_X1 U22531 ( .A(n19457), .B(n21360), .S(n28586), .Z(n19459) );
  XNOR2_X1 U22533 ( .A(n22671), .B(n22698), .ZN(n22031) );
  INV_X1 U22534 ( .A(n22031), .ZN(n21756) );
  XNOR2_X1 U22535 ( .A(n29580), .B(n19462), .ZN(n19467) );
  XNOR2_X1 U22536 ( .A(n19464), .B(n19465), .ZN(n19466) );
  XNOR2_X1 U22537 ( .A(n19466), .B(n19467), .ZN(n19471) );
  INV_X1 U22538 ( .A(n27422), .ZN(n25250) );
  XNOR2_X1 U22539 ( .A(n19468), .B(n25250), .ZN(n19469) );
  XNOR2_X1 U22540 ( .A(n19474), .B(n19726), .ZN(n19477) );
  XNOR2_X1 U22541 ( .A(n19475), .B(n2982), .ZN(n19476) );
  XNOR2_X1 U22542 ( .A(n19477), .B(n19476), .ZN(n19478) );
  INV_X1 U22543 ( .A(n20130), .ZN(n19901) );
  MUX2_X1 U22544 ( .A(n20443), .B(n415), .S(n19901), .Z(n19506) );
  XNOR2_X1 U22545 ( .A(n19670), .B(n3673), .ZN(n19485) );
  XNOR2_X1 U22546 ( .A(n19484), .B(n19485), .ZN(n19489) );
  XNOR2_X1 U22547 ( .A(n19486), .B(n19487), .ZN(n19488) );
  XNOR2_X1 U22548 ( .A(n19489), .B(n19488), .ZN(n19494) );
  XNOR2_X1 U22549 ( .A(n19491), .B(n19490), .ZN(n19492) );
  INV_X1 U22550 ( .A(n19495), .ZN(n19497) );
  XNOR2_X1 U22551 ( .A(n19496), .B(n19497), .ZN(n19499) );
  XNOR2_X1 U22552 ( .A(n19498), .B(n19499), .ZN(n19504) );
  XNOR2_X1 U22553 ( .A(n19500), .B(n1161), .ZN(n19501) );
  XNOR2_X1 U22554 ( .A(n19502), .B(n19501), .ZN(n19503) );
  XNOR2_X1 U22555 ( .A(n19507), .B(n19508), .ZN(n19509) );
  XNOR2_X1 U22556 ( .A(n19510), .B(n19509), .ZN(n19515) );
  XNOR2_X1 U22557 ( .A(n19511), .B(n2577), .ZN(n19512) );
  XNOR2_X1 U22558 ( .A(n19513), .B(n19512), .ZN(n19514) );
  INV_X1 U22559 ( .A(n20125), .ZN(n20294) );
  INV_X1 U22560 ( .A(n20293), .ZN(n19814) );
  INV_X1 U22561 ( .A(n20123), .ZN(n19969) );
  INV_X1 U22562 ( .A(n20295), .ZN(n19818) );
  AOI21_X1 U22563 ( .B1(n20290), .B2(n19969), .A(n19818), .ZN(n19517) );
  NAND2_X1 U22564 ( .A1(n20123), .A2(n19814), .ZN(n19516) );
  XNOR2_X1 U22565 ( .A(n19519), .B(n19518), .ZN(n19524) );
  XNOR2_X1 U22566 ( .A(n19520), .B(n19611), .ZN(n19522) );
  XNOR2_X1 U22567 ( .A(n19617), .B(n3196), .ZN(n19521) );
  XNOR2_X1 U22568 ( .A(n19522), .B(n19521), .ZN(n19523) );
  XNOR2_X1 U22569 ( .A(n19524), .B(n19523), .ZN(n20647) );
  XNOR2_X1 U22570 ( .A(n19525), .B(n3644), .ZN(n19527) );
  XNOR2_X1 U22571 ( .A(n19526), .B(n19527), .ZN(n19531) );
  XNOR2_X1 U22572 ( .A(n19528), .B(n19529), .ZN(n19530) );
  XNOR2_X1 U22574 ( .A(n19533), .B(n19532), .ZN(n19539) );
  XNOR2_X1 U22575 ( .A(n19595), .B(n19534), .ZN(n19537) );
  XNOR2_X1 U22576 ( .A(n19535), .B(n3334), .ZN(n19536) );
  XNOR2_X1 U22577 ( .A(n19537), .B(n19536), .ZN(n19538) );
  INV_X1 U22578 ( .A(n19540), .ZN(n19542) );
  XNOR2_X1 U22579 ( .A(n19542), .B(n19541), .ZN(n19545) );
  INV_X1 U22580 ( .A(n19546), .ZN(n19547) );
  XNOR2_X1 U22581 ( .A(n19547), .B(n19548), .ZN(n19553) );
  XNOR2_X1 U22582 ( .A(n19727), .B(n19585), .ZN(n19551) );
  XNOR2_X1 U22583 ( .A(n19549), .B(n2441), .ZN(n19550) );
  XNOR2_X1 U22584 ( .A(n19551), .B(n19550), .ZN(n19552) );
  XNOR2_X1 U22585 ( .A(n19555), .B(n28143), .ZN(n19558) );
  XNOR2_X1 U22586 ( .A(n19557), .B(n19558), .ZN(n19572) );
  INV_X1 U22587 ( .A(n19559), .ZN(n19566) );
  NAND3_X1 U22588 ( .A1(n29125), .A2(n29044), .A3(n123), .ZN(n19563) );
  NAND2_X1 U22589 ( .A1(n19564), .A2(n19563), .ZN(n19565) );
  NOR2_X1 U22590 ( .A1(n19566), .A2(n19565), .ZN(n19567) );
  XNOR2_X1 U22591 ( .A(n19577), .B(n19567), .ZN(n19570) );
  XNOR2_X1 U22592 ( .A(n19570), .B(n19569), .ZN(n19571) );
  XNOR2_X1 U22593 ( .A(n19571), .B(n19572), .ZN(n19928) );
  OAI21_X1 U22594 ( .B1(n21807), .B2(n21806), .A(n21253), .ZN(n19735) );
  XNOR2_X1 U22595 ( .A(n19574), .B(n19575), .ZN(n19581) );
  XNOR2_X1 U22596 ( .A(n19637), .B(n29318), .ZN(n19579) );
  XNOR2_X1 U22597 ( .A(n19577), .B(n3528), .ZN(n19578) );
  XNOR2_X1 U22598 ( .A(n19579), .B(n19578), .ZN(n19580) );
  XNOR2_X1 U22599 ( .A(n19583), .B(n19582), .ZN(n19589) );
  XNOR2_X1 U22600 ( .A(n19584), .B(n3378), .ZN(n19587) );
  XNOR2_X1 U22601 ( .A(n19644), .B(n19585), .ZN(n19586) );
  XNOR2_X1 U22602 ( .A(n19586), .B(n19587), .ZN(n19588) );
  XNOR2_X1 U22603 ( .A(n19592), .B(n28693), .ZN(n19593) );
  NOR2_X1 U22604 ( .A1(n20109), .A2(n20319), .ZN(n19602) );
  XNOR2_X1 U22605 ( .A(n19595), .B(n3083), .ZN(n19596) );
  XNOR2_X1 U22606 ( .A(n19597), .B(n19596), .ZN(n19601) );
  XNOR2_X1 U22607 ( .A(n19599), .B(n19598), .ZN(n19600) );
  MUX2_X1 U22608 ( .A(n20323), .B(n19602), .S(n20322), .Z(n20694) );
  XNOR2_X1 U22609 ( .A(n18638), .B(n19603), .ZN(n19605) );
  XNOR2_X1 U22610 ( .A(n19605), .B(n19604), .ZN(n19610) );
  XNOR2_X1 U22611 ( .A(n19606), .B(n2996), .ZN(n19608) );
  XNOR2_X1 U22612 ( .A(n19607), .B(n19608), .ZN(n19609) );
  XNOR2_X2 U22613 ( .A(n19609), .B(n19610), .ZN(n20324) );
  INV_X1 U22614 ( .A(n19611), .ZN(n19612) );
  XNOR2_X1 U22615 ( .A(n19612), .B(n19669), .ZN(n19614) );
  XNOR2_X1 U22616 ( .A(n19614), .B(n19613), .ZN(n19621) );
  XNOR2_X1 U22617 ( .A(n19616), .B(n19615), .ZN(n19619) );
  XNOR2_X1 U22618 ( .A(n19617), .B(n2403), .ZN(n19618) );
  XNOR2_X1 U22619 ( .A(n19619), .B(n19618), .ZN(n19620) );
  XNOR2_X1 U22620 ( .A(n19620), .B(n19621), .ZN(n19955) );
  INV_X1 U22621 ( .A(n19955), .ZN(n19956) );
  NAND3_X1 U22622 ( .A1(n19956), .A2(n20320), .A3(n2180), .ZN(n20693) );
  NOR2_X1 U22623 ( .A1(n21809), .A2(n21810), .ZN(n21007) );
  XNOR2_X1 U22624 ( .A(n19622), .B(n3109), .ZN(n19623) );
  XNOR2_X1 U22625 ( .A(n19624), .B(n19623), .ZN(n19630) );
  XNOR2_X1 U22626 ( .A(n19625), .B(n19626), .ZN(n19627) );
  XOR2_X1 U22627 ( .A(n19628), .B(n19627), .Z(n19629) );
  XNOR2_X1 U22628 ( .A(n19630), .B(n19629), .ZN(n19810) );
  XNOR2_X1 U22629 ( .A(n19636), .B(n3695), .ZN(n19638) );
  XNOR2_X1 U22630 ( .A(n19638), .B(n19637), .ZN(n19640) );
  XNOR2_X1 U22631 ( .A(n19640), .B(n19639), .ZN(n19642) );
  XNOR2_X1 U22632 ( .A(n19642), .B(n19641), .ZN(n19938) );
  MUX2_X1 U22634 ( .A(n29166), .B(n29707), .S(n20281), .Z(n19677) );
  XNOR2_X1 U22635 ( .A(n19643), .B(n1928), .ZN(n19645) );
  XNOR2_X1 U22636 ( .A(n19645), .B(n19644), .ZN(n19647) );
  XNOR2_X1 U22637 ( .A(n19647), .B(n19646), .ZN(n19648) );
  INV_X1 U22638 ( .A(n19650), .ZN(n19652) );
  INV_X1 U22639 ( .A(n28516), .ZN(n19654) );
  XNOR2_X1 U22640 ( .A(n19655), .B(n19654), .ZN(n19663) );
  INV_X1 U22641 ( .A(n19659), .ZN(n19657) );
  NAND2_X1 U22642 ( .A1(n19657), .A2(n3386), .ZN(n19661) );
  OAI21_X1 U22643 ( .B1(n19656), .B2(n19659), .A(n19658), .ZN(n19660) );
  OAI21_X1 U22644 ( .B1(n19656), .B2(n19661), .A(n19660), .ZN(n19662) );
  XNOR2_X1 U22645 ( .A(n19663), .B(n19662), .ZN(n19664) );
  INV_X1 U22646 ( .A(n19665), .ZN(n19667) );
  XNOR2_X1 U22647 ( .A(n19667), .B(n19666), .ZN(n19674) );
  XNOR2_X1 U22648 ( .A(n19668), .B(n19669), .ZN(n19672) );
  XNOR2_X1 U22649 ( .A(n29554), .B(n28327), .ZN(n19671) );
  XNOR2_X1 U22650 ( .A(n19672), .B(n19671), .ZN(n19673) );
  INV_X1 U22651 ( .A(n20283), .ZN(n20285) );
  NAND2_X1 U22652 ( .A1(n20285), .A2(n20281), .ZN(n19675) );
  NAND2_X1 U22653 ( .A1(n20289), .A2(n19675), .ZN(n19676) );
  XNOR2_X1 U22654 ( .A(n19678), .B(n3223), .ZN(n19680) );
  XNOR2_X1 U22655 ( .A(n19680), .B(n19679), .ZN(n19682) );
  XNOR2_X1 U22656 ( .A(n19682), .B(n19681), .ZN(n19684) );
  INV_X1 U22658 ( .A(n20440), .ZN(n20608) );
  XNOR2_X1 U22659 ( .A(n19691), .B(n19692), .ZN(n19694) );
  XNOR2_X1 U22660 ( .A(n19695), .B(n19696), .ZN(n19699) );
  XNOR2_X1 U22661 ( .A(n19697), .B(n3527), .ZN(n19698) );
  MUX2_X1 U22662 ( .A(n29625), .B(n20608), .S(n20441), .Z(n19731) );
  XNOR2_X1 U22663 ( .A(n19701), .B(n19700), .ZN(n19703) );
  XNOR2_X1 U22664 ( .A(n19703), .B(n19702), .ZN(n19713) );
  INV_X1 U22665 ( .A(n19704), .ZN(n19705) );
  XNOR2_X1 U22666 ( .A(n19706), .B(n19705), .ZN(n19711) );
  XNOR2_X1 U22667 ( .A(n19707), .B(n2510), .ZN(n19708) );
  XNOR2_X1 U22668 ( .A(n19708), .B(n19709), .ZN(n19710) );
  XNOR2_X1 U22669 ( .A(n19710), .B(n19711), .ZN(n19712) );
  XNOR2_X1 U22670 ( .A(n19712), .B(n19713), .ZN(n20609) );
  XNOR2_X1 U22672 ( .A(n19714), .B(n19715), .ZN(n19722) );
  XNOR2_X1 U22673 ( .A(n19716), .B(n19717), .ZN(n19720) );
  XNOR2_X1 U22674 ( .A(n19718), .B(n2353), .ZN(n19719) );
  XNOR2_X1 U22675 ( .A(n19720), .B(n19719), .ZN(n19721) );
  XNOR2_X1 U22676 ( .A(n19726), .B(n28571), .ZN(n19729) );
  XNOR2_X1 U22677 ( .A(n19727), .B(n1062), .ZN(n19728) );
  XNOR2_X1 U22678 ( .A(n19729), .B(n19728), .ZN(n19730) );
  NOR2_X1 U22679 ( .A1(n21811), .A2(n21253), .ZN(n20698) );
  OAI211_X2 U22680 ( .C1(n21007), .C2(n19735), .A(n19734), .B(n19733), .ZN(
        n22295) );
  XNOR2_X1 U22681 ( .A(n22295), .B(n1133), .ZN(n19736) );
  XNOR2_X1 U22682 ( .A(n21756), .B(n19736), .ZN(n19737) );
  MUX2_X1 U22683 ( .A(n19739), .B(n20377), .S(n351), .Z(n19742) );
  MUX2_X1 U22684 ( .A(n20371), .B(n20373), .S(n20372), .Z(n19741) );
  INV_X1 U22685 ( .A(n20401), .ZN(n20558) );
  INV_X1 U22686 ( .A(n20208), .ZN(n20400) );
  OAI21_X1 U22687 ( .B1(n20558), .B2(n29041), .A(n20209), .ZN(n19746) );
  NAND2_X1 U22688 ( .A1(n20394), .A2(n20563), .ZN(n19744) );
  INV_X1 U22689 ( .A(n19851), .ZN(n20562) );
  MUX2_X1 U22690 ( .A(n19744), .B(n19743), .S(n20562), .Z(n19745) );
  INV_X1 U22691 ( .A(n19747), .ZN(n20417) );
  NAND2_X1 U22693 ( .A1(n20412), .A2(n20414), .ZN(n19749) );
  NAND2_X1 U22694 ( .A1(n503), .A2(n20577), .ZN(n19748) );
  INV_X1 U22695 ( .A(n22140), .ZN(n22142) );
  MUX2_X1 U22696 ( .A(n20383), .B(n19837), .S(n20567), .Z(n19751) );
  INV_X1 U22697 ( .A(n19836), .ZN(n19750) );
  INV_X1 U22698 ( .A(n28526), .ZN(n19844) );
  NOR2_X1 U22699 ( .A1(n18837), .A2(n19844), .ZN(n19754) );
  OAI211_X1 U22700 ( .C1(n6495), .C2(n29551), .A(n29582), .B(n20083), .ZN(
        n19753) );
  INV_X1 U22701 ( .A(n20041), .ZN(n20092) );
  NAND2_X1 U22702 ( .A1(n20092), .A2(n414), .ZN(n19756) );
  AOI21_X1 U22703 ( .B1(n19756), .B2(n19755), .A(n20039), .ZN(n19759) );
  NAND2_X1 U22704 ( .A1(n20041), .A2(n29114), .ZN(n19757) );
  MUX2_X1 U22705 ( .A(n29540), .B(n22145), .S(n22143), .Z(n19760) );
  NAND2_X1 U22706 ( .A1(n29540), .A2(n6532), .ZN(n21626) );
  NAND2_X1 U22707 ( .A1(n20069), .A2(n20049), .ZN(n19762) );
  NAND3_X1 U22708 ( .A1(n20048), .A2(n18765), .A3(n20049), .ZN(n19763) );
  INV_X1 U22709 ( .A(n19766), .ZN(n20146) );
  NOR2_X1 U22710 ( .A1(n20146), .A2(n28479), .ZN(n19767) );
  AOI22_X1 U22711 ( .A1(n20146), .A2(n29134), .B1(n19767), .B2(n20144), .ZN(
        n19768) );
  INV_X1 U22713 ( .A(n20158), .ZN(n20160) );
  OAI21_X1 U22716 ( .B1(n20163), .B2(n19769), .A(n28187), .ZN(n19772) );
  AOI21_X1 U22717 ( .B1(n19984), .B2(n20162), .A(n20159), .ZN(n19770) );
  OR2_X1 U22718 ( .A1(n19770), .A2(n20158), .ZN(n19771) );
  OAI21_X1 U22719 ( .B1(n28188), .B2(n19773), .A(n20043), .ZN(n19774) );
  OAI21_X1 U22720 ( .B1(n20092), .B2(n29114), .A(n20093), .ZN(n19777) );
  NOR2_X1 U22722 ( .A1(n20851), .A2(n21143), .ZN(n19783) );
  AND2_X1 U22723 ( .A1(n21118), .A2(n21143), .ZN(n19782) );
  XNOR2_X1 U22724 ( .A(n22194), .B(n22784), .ZN(n19805) );
  INV_X1 U22725 ( .A(n20349), .ZN(n19785) );
  NOR2_X1 U22726 ( .A1(n20013), .A2(n20342), .ZN(n19786) );
  INV_X1 U22727 ( .A(n20017), .ZN(n20345) );
  INV_X1 U22728 ( .A(n20343), .ZN(n20014) );
  NOR2_X1 U22729 ( .A1(n20247), .A2(n20453), .ZN(n19788) );
  OAI21_X1 U22731 ( .B1(n19788), .B2(n20032), .A(n20637), .ZN(n19790) );
  NAND2_X1 U22732 ( .A1(n20247), .A2(n28538), .ZN(n19789) );
  INV_X1 U22734 ( .A(n20481), .ZN(n20001) );
  NAND2_X1 U22735 ( .A1(n19793), .A2(n28155), .ZN(n19803) );
  INV_X1 U22736 ( .A(n21356), .ZN(n20023) );
  AND2_X1 U22738 ( .A1(n28610), .A2(n21355), .ZN(n20024) );
  INV_X1 U22739 ( .A(n21359), .ZN(n21354) );
  NAND2_X1 U22740 ( .A1(n21354), .A2(n19796), .ZN(n19797) );
  OAI21_X1 U22741 ( .B1(n20024), .B2(n21354), .A(n19797), .ZN(n19798) );
  NOR2_X1 U22742 ( .A1(n20498), .A2(n20499), .ZN(n19800) );
  NAND2_X1 U22744 ( .A1(n20333), .A2(n20334), .ZN(n20631) );
  INV_X1 U22745 ( .A(n20625), .ZN(n20628) );
  INV_X1 U22746 ( .A(n20626), .ZN(n20330) );
  NAND3_X1 U22747 ( .A1(n20628), .A2(n20005), .A3(n20330), .ZN(n19802) );
  XNOR2_X1 U22748 ( .A(n28449), .B(n27605), .ZN(n19804) );
  XNOR2_X1 U22749 ( .A(n19805), .B(n19804), .ZN(n19909) );
  INV_X1 U22750 ( .A(n20201), .ZN(n20305) );
  MUX2_X1 U22751 ( .A(n20202), .B(n20305), .S(n20200), .Z(n19807) );
  NOR2_X1 U22752 ( .A1(n416), .A2(n20200), .ZN(n19806) );
  NAND2_X1 U22753 ( .A1(n20205), .A2(n20302), .ZN(n20306) );
  NAND2_X1 U22754 ( .A1(n19810), .A2(n20284), .ZN(n19939) );
  INV_X1 U22755 ( .A(n19939), .ZN(n19809) );
  OAI21_X1 U22756 ( .B1(n2081), .B2(n19809), .A(n2152), .ZN(n19813) );
  INV_X1 U22757 ( .A(n19810), .ZN(n20286) );
  AOI21_X1 U22758 ( .B1(n20281), .B2(n20284), .A(n20286), .ZN(n19811) );
  NAND2_X1 U22759 ( .A1(n19967), .A2(n20123), .ZN(n20292) );
  INV_X1 U22760 ( .A(n19815), .ZN(n19968) );
  OAI22_X1 U22761 ( .A1(n20292), .A2(n19818), .B1(n19967), .B2(n20122), .ZN(
        n19817) );
  AND2_X1 U22762 ( .A1(n19818), .A2(n19815), .ZN(n20124) );
  INV_X1 U22763 ( .A(n20124), .ZN(n19816) );
  INV_X1 U22765 ( .A(n20546), .ZN(n20191) );
  NOR2_X1 U22766 ( .A1(n19820), .A2(n20389), .ZN(n19819) );
  AND2_X1 U22767 ( .A1(n20544), .A2(n20546), .ZN(n20190) );
  OAI21_X1 U22768 ( .B1(n20190), .B2(n20388), .A(n19820), .ZN(n19821) );
  INV_X1 U22769 ( .A(n20319), .ZN(n19940) );
  NAND2_X1 U22770 ( .A1(n19940), .A2(n20323), .ZN(n19822) );
  MUX2_X1 U22771 ( .A(n19822), .B(n20112), .S(n20324), .Z(n19826) );
  NOR2_X1 U22772 ( .A1(n20323), .A2(n20320), .ZN(n19824) );
  NOR2_X1 U22773 ( .A1(n19940), .A2(n20322), .ZN(n19823) );
  AOI22_X1 U22774 ( .A1(n19824), .A2(n19940), .B1(n19823), .B2(n502), .ZN(
        n19825) );
  NAND2_X1 U22775 ( .A1(n20311), .A2(n19949), .ZN(n19829) );
  INV_X1 U22776 ( .A(n20196), .ZN(n20588) );
  OR2_X1 U22777 ( .A1(n21495), .A2(n21496), .ZN(n19830) );
  NAND2_X1 U22778 ( .A1(n19834), .A2(n19838), .ZN(n19839) );
  OAI211_X1 U22779 ( .C1(n20379), .C2(n20373), .A(n351), .B(n20374), .ZN(
        n19842) );
  OAI21_X1 U22780 ( .B1(n6495), .B2(n20083), .A(n29582), .ZN(n19848) );
  NOR2_X1 U22781 ( .A1(n6495), .A2(n19844), .ZN(n19846) );
  AND2_X1 U22782 ( .A1(n19851), .A2(n20208), .ZN(n20396) );
  NAND2_X1 U22783 ( .A1(n20401), .A2(n20396), .ZN(n19854) );
  INV_X1 U22784 ( .A(n19849), .ZN(n19850) );
  NAND3_X1 U22785 ( .A1(n20209), .A2(n20562), .A3(n20563), .ZN(n19852) );
  NAND2_X1 U22786 ( .A1(n20749), .A2(n21574), .ZN(n21487) );
  MUX2_X1 U22787 ( .A(n20941), .B(n20577), .S(n28140), .Z(n19858) );
  XNOR2_X1 U22789 ( .A(n22661), .B(n21758), .ZN(n22575) );
  INV_X1 U22790 ( .A(n22575), .ZN(n19907) );
  OAI21_X1 U22793 ( .B1(n5303), .B2(n29616), .A(n20218), .ZN(n19864) );
  OAI21_X1 U22794 ( .B1(n19865), .B2(n20218), .A(n19864), .ZN(n19866) );
  INV_X1 U22795 ( .A(n21155), .ZN(n21158) );
  NAND2_X1 U22796 ( .A1(n19032), .A2(n382), .ZN(n20737) );
  INV_X1 U22797 ( .A(n20176), .ZN(n20054) );
  NOR2_X1 U22798 ( .A1(n19868), .A2(n20171), .ZN(n19869) );
  INV_X1 U22800 ( .A(n20144), .ZN(n20106) );
  NAND2_X1 U22801 ( .A1(n20527), .A2(n20858), .ZN(n19871) );
  INV_X1 U22802 ( .A(n20159), .ZN(n19981) );
  MUX2_X1 U22803 ( .A(n20160), .B(n20157), .S(n19981), .Z(n19876) );
  NOR2_X1 U22804 ( .A1(n19981), .A2(n29066), .ZN(n19873) );
  AOI22_X1 U22805 ( .A1(n19874), .A2(n19873), .B1(n19985), .B2(n19872), .ZN(
        n19875) );
  NAND2_X1 U22806 ( .A1(n494), .A2(n21159), .ZN(n21111) );
  OAI21_X1 U22808 ( .B1(n21111), .B2(n20858), .A(n19877), .ZN(n19878) );
  NOR2_X2 U22809 ( .A1(n19879), .A2(n19878), .ZN(n22218) );
  NAND2_X1 U22810 ( .A1(n20603), .A2(n1915), .ZN(n19880) );
  NOR2_X1 U22811 ( .A1(n20601), .A2(n20272), .ZN(n19883) );
  NOR2_X1 U22812 ( .A1(n20603), .A2(n20272), .ZN(n19882) );
  NOR3_X1 U22813 ( .A1(n19882), .A2(n28408), .A3(n19883), .ZN(n19884) );
  NOR2_X1 U22814 ( .A1(n19886), .A2(n20607), .ZN(n19888) );
  INV_X1 U22815 ( .A(n20618), .ZN(n19889) );
  AOI21_X1 U22816 ( .B1(n19889), .B2(n6567), .A(n20616), .ZN(n19891) );
  NOR2_X1 U22820 ( .A1(n20622), .A2(n19920), .ZN(n19893) );
  NOR2_X1 U22821 ( .A1(n20137), .A2(n19808), .ZN(n19895) );
  NOR2_X1 U22823 ( .A1(n20281), .A2(n20137), .ZN(n19897) );
  NOR2_X1 U22824 ( .A1(n20449), .A2(n20265), .ZN(n20450) );
  NAND2_X1 U22825 ( .A1(n20450), .A2(n5377), .ZN(n19900) );
  AOI211_X1 U22826 ( .C1(n415), .C2(n20444), .A(n3247), .B(n19901), .ZN(n19902) );
  INV_X1 U22827 ( .A(n21459), .ZN(n20842) );
  NAND2_X1 U22828 ( .A1(n1814), .A2(n20842), .ZN(n19904) );
  XNOR2_X1 U22830 ( .A(n22218), .B(n22279), .ZN(n19906) );
  XNOR2_X1 U22831 ( .A(n19907), .B(n19906), .ZN(n19908) );
  NOR2_X1 U22832 ( .A1(n23535), .A2(n23529), .ZN(n20473) );
  NAND2_X1 U22833 ( .A1(n22139), .A2(n22145), .ZN(n21029) );
  INV_X1 U22834 ( .A(n29540), .ZN(n22146) );
  NAND3_X1 U22835 ( .A1(n22146), .A2(n22139), .A3(n22143), .ZN(n19911) );
  NOR2_X1 U22836 ( .A1(n5939), .A2(n22139), .ZN(n21623) );
  MUX2_X1 U22838 ( .A(n20972), .B(n21217), .S(n21000), .Z(n19912) );
  NOR2_X1 U22839 ( .A1(n19912), .A2(n21220), .ZN(n19918) );
  NAND2_X1 U22841 ( .A1(n28980), .A2(n21218), .ZN(n19916) );
  NAND2_X1 U22842 ( .A1(n20966), .A2(n19914), .ZN(n20701) );
  OAI21_X1 U22843 ( .B1(n19916), .B2(n20701), .A(n19915), .ZN(n19917) );
  XNOR2_X1 U22844 ( .A(n21875), .B(n22330), .ZN(n19945) );
  NAND3_X1 U22845 ( .A1(n20255), .A2(n28894), .A3(n20616), .ZN(n19919) );
  OAI21_X1 U22846 ( .B1(n19901), .B2(n20443), .A(n19924), .ZN(n19925) );
  INV_X1 U22847 ( .A(n21748), .ZN(n21401) );
  NAND2_X1 U22849 ( .A1(n28555), .A2(n20440), .ZN(n19935) );
  NAND3_X1 U22850 ( .A1(n20441), .A2(n29508), .A3(n20607), .ZN(n19937) );
  NAND2_X1 U22851 ( .A1(n21642), .A2(n20658), .ZN(n21040) );
  AOI22_X1 U22852 ( .A1(n502), .A2(n20109), .B1(n20323), .B2(n20322), .ZN(
        n19942) );
  AND2_X1 U22853 ( .A1(n20109), .A2(n19955), .ZN(n20325) );
  OAI21_X1 U22854 ( .B1(n20325), .B2(n19940), .A(n2181), .ZN(n19941) );
  NAND2_X1 U22856 ( .A1(n20659), .A2(n497), .ZN(n19943) );
  XNOR2_X1 U22857 ( .A(n22265), .B(n2960), .ZN(n19944) );
  XNOR2_X1 U22858 ( .A(n19945), .B(n19944), .ZN(n20062) );
  NOR2_X1 U22859 ( .A1(n20205), .A2(n20302), .ZN(n19946) );
  INV_X1 U22860 ( .A(n20302), .ZN(n20119) );
  NOR2_X1 U22861 ( .A1(n19949), .A2(n20584), .ZN(n19950) );
  INV_X1 U22862 ( .A(n20585), .ZN(n20315) );
  MUX2_X1 U22863 ( .A(n20315), .B(n20196), .S(n20314), .Z(n19952) );
  NOR2_X1 U22864 ( .A1(n19952), .A2(n3973), .ZN(n19953) );
  NOR2_X1 U22865 ( .A1(n21472), .A2(n1930), .ZN(n21733) );
  NAND2_X1 U22866 ( .A1(n502), .A2(n20319), .ZN(n19957) );
  OAI21_X1 U22867 ( .B1(n20546), .B2(n20544), .A(n20188), .ZN(n19961) );
  AOI22_X2 U22868 ( .A1(n20392), .A2(n19961), .B1(n19960), .B2(n19959), .ZN(
        n21473) );
  MUX2_X1 U22869 ( .A(n21733), .B(n21388), .S(n21473), .Z(n19975) );
  INV_X1 U22870 ( .A(n19962), .ZN(n19966) );
  INV_X1 U22871 ( .A(n20405), .ZN(n20553) );
  NOR2_X1 U22872 ( .A1(n20556), .A2(n20553), .ZN(n19964) );
  OAI21_X1 U22873 ( .B1(n19964), .B2(n20404), .A(n505), .ZN(n21032) );
  OAI21_X1 U22874 ( .B1(n19968), .B2(n20125), .A(n19967), .ZN(n19972) );
  NOR2_X1 U22875 ( .A1(n19969), .A2(n20295), .ZN(n19970) );
  OAI21_X1 U22877 ( .B1(n21471), .B2(n21731), .A(n21477), .ZN(n19974) );
  INV_X1 U22878 ( .A(n20055), .ZN(n19980) );
  MUX2_X1 U22879 ( .A(n20178), .B(n20173), .S(n19976), .Z(n19978) );
  MUX2_X1 U22880 ( .A(n19978), .B(n19977), .S(n20054), .Z(n19979) );
  OAI21_X1 U22881 ( .B1(n19982), .B2(n19981), .A(n20164), .ZN(n19988) );
  AOI21_X1 U22882 ( .B1(n19985), .B2(n19984), .A(n19983), .ZN(n20047) );
  NOR2_X1 U22884 ( .A1(n297), .A2(n19989), .ZN(n19990) );
  NOR2_X1 U22885 ( .A1(n385), .A2(n19992), .ZN(n19994) );
  OAI211_X1 U22886 ( .C1(n20479), .C2(n19997), .A(n20475), .B(n383), .ZN(
        n19999) );
  NAND2_X1 U22887 ( .A1(n5408), .A2(n20478), .ZN(n19996) );
  NOR2_X1 U22888 ( .A1(n19996), .A2(n20477), .ZN(n19998) );
  NOR2_X1 U22889 ( .A1(n28620), .A2(n20000), .ZN(n20002) );
  AOI22_X1 U22890 ( .A1(n20002), .A2(n20001), .B1(n29527), .B2(n20485), .ZN(
        n20004) );
  XNOR2_X1 U22891 ( .A(n21956), .B(n22633), .ZN(n20060) );
  INV_X1 U22893 ( .A(n20623), .ZN(n20258) );
  NOR2_X1 U22895 ( .A1(n28515), .A2(n20012), .ZN(n20670) );
  NOR3_X1 U22896 ( .A1(n20675), .A2(n21638), .A3(n20670), .ZN(n20031) );
  INV_X1 U22897 ( .A(n20013), .ZN(n20344) );
  MUX2_X1 U22898 ( .A(n28489), .B(n19785), .S(n20344), .Z(n20016) );
  NOR2_X1 U22899 ( .A1(n20345), .A2(n20342), .ZN(n20015) );
  INV_X1 U22900 ( .A(n20347), .ZN(n20019) );
  NAND2_X1 U22901 ( .A1(n20511), .A2(n20349), .ZN(n20018) );
  NOR2_X1 U22902 ( .A1(n20019), .A2(n20018), .ZN(n20671) );
  NOR2_X2 U22903 ( .A1(n20669), .A2(n20671), .ZN(n21639) );
  MUX2_X1 U22905 ( .A(n20518), .B(n20021), .S(n21359), .Z(n20026) );
  NOR2_X1 U22906 ( .A1(n28610), .A2(n28491), .ZN(n20022) );
  AOI22_X1 U22907 ( .A1(n20024), .A2(n20023), .B1(n20022), .B2(n28586), .ZN(
        n20025) );
  NAND3_X1 U22908 ( .A1(n386), .A2(n20603), .A3(n20028), .ZN(n20029) );
  AND2_X1 U22909 ( .A1(n20033), .A2(n20453), .ZN(n20252) );
  NOR2_X1 U22912 ( .A1(n21092), .A2(n20146), .ZN(n20038) );
  NOR2_X1 U22913 ( .A1(n21091), .A2(n21095), .ZN(n20036) );
  AOI22_X1 U22914 ( .A1(n20038), .A2(n20148), .B1(n20036), .B2(n18919), .ZN(
        n20037) );
  NAND3_X1 U22916 ( .A1(n20045), .A2(n20158), .A3(n20044), .ZN(n20046) );
  OAI21_X1 U22917 ( .B1(n20047), .B2(n20163), .A(n20046), .ZN(n21211) );
  NAND2_X1 U22919 ( .A1(n20052), .A2(n28448), .ZN(n21209) );
  INV_X1 U22920 ( .A(n20053), .ZN(n20056) );
  NAND3_X1 U22921 ( .A1(n20056), .A2(n504), .A3(n20173), .ZN(n20057) );
  XNOR2_X1 U22922 ( .A(n22643), .B(n22690), .ZN(n20059) );
  XNOR2_X1 U22923 ( .A(n20060), .B(n20059), .ZN(n20061) );
  MUX2_X1 U22924 ( .A(n20065), .B(n20064), .S(n20063), .Z(n20067) );
  OAI21_X1 U22925 ( .B1(n351), .B2(n20374), .A(n20377), .ZN(n20072) );
  NAND2_X1 U22926 ( .A1(n20372), .A2(n20072), .ZN(n20073) );
  INV_X1 U22927 ( .A(n20075), .ZN(n20079) );
  NOR2_X1 U22928 ( .A1(n18837), .A2(n29315), .ZN(n20078) );
  NOR2_X1 U22930 ( .A1(n20081), .A2(n29551), .ZN(n20082) );
  AOI22_X1 U22931 ( .A1(n20084), .A2(n20083), .B1(n20082), .B2(n18837), .ZN(
        n20085) );
  NOR2_X1 U22932 ( .A1(n22013), .A2(n20532), .ZN(n21818) );
  NOR2_X1 U22933 ( .A1(n20155), .A2(n20096), .ZN(n20101) );
  NAND2_X1 U22934 ( .A1(n20097), .A2(n18887), .ZN(n20100) );
  NAND2_X1 U22935 ( .A1(n21078), .A2(n495), .ZN(n20108) );
  NAND2_X1 U22936 ( .A1(n18919), .A2(n20102), .ZN(n20107) );
  AOI21_X1 U22937 ( .B1(n29134), .B2(n20102), .A(n21091), .ZN(n20104) );
  NOR2_X1 U22938 ( .A1(n18919), .A2(n28479), .ZN(n20103) );
  OAI22_X1 U22939 ( .A1(n20104), .A2(n20103), .B1(n20102), .B2(n4877), .ZN(
        n20105) );
  NOR2_X1 U22940 ( .A1(n20320), .A2(n20319), .ZN(n20110) );
  NOR2_X1 U22941 ( .A1(n20112), .A2(n20324), .ZN(n20897) );
  NOR2_X1 U22942 ( .A1(n20607), .A2(n20440), .ZN(n20113) );
  NOR2_X1 U22943 ( .A1(n20113), .A2(n20441), .ZN(n20116) );
  NOR2_X1 U22944 ( .A1(n20441), .A2(n20440), .ZN(n20114) );
  NOR2_X1 U22945 ( .A1(n20609), .A2(n29508), .ZN(n20435) );
  OAI21_X1 U22946 ( .B1(n20114), .B2(n20435), .A(n20614), .ZN(n20115) );
  INV_X1 U22947 ( .A(n20898), .ZN(n20129) );
  INV_X1 U22948 ( .A(n20897), .ZN(n20118) );
  OAI21_X1 U22949 ( .B1(n20295), .B2(n20123), .A(n20122), .ZN(n20127) );
  NAND2_X1 U22950 ( .A1(n20125), .A2(n20124), .ZN(n20126) );
  INV_X1 U22951 ( .A(n20299), .ZN(n20131) );
  NOR2_X1 U22952 ( .A1(n20131), .A2(n20130), .ZN(n20132) );
  NOR2_X1 U22953 ( .A1(n20446), .A2(n20132), .ZN(n20134) );
  NAND3_X1 U22954 ( .A1(n19938), .A2(n19808), .A3(n20286), .ZN(n20136) );
  NAND2_X1 U22955 ( .A1(n20141), .A2(n20140), .ZN(n20142) );
  XNOR2_X1 U22956 ( .A(n22098), .B(n22270), .ZN(n20215) );
  NOR2_X1 U22957 ( .A1(n29134), .A2(n20144), .ZN(n21096) );
  NAND2_X1 U22958 ( .A1(n20149), .A2(n20148), .ZN(n21097) );
  INV_X1 U22959 ( .A(n21097), .ZN(n20953) );
  AOI21_X1 U22960 ( .B1(n20152), .B2(n20151), .A(n20150), .ZN(n20153) );
  NOR3_X1 U22961 ( .A1(n20954), .A2(n20953), .A3(n21932), .ZN(n20187) );
  NOR2_X1 U22962 ( .A1(n20165), .A2(n385), .ZN(n20170) );
  AND3_X1 U22963 ( .A1(n20166), .A2(n297), .A3(n20219), .ZN(n20167) );
  NOR2_X1 U22964 ( .A1(n20168), .A2(n20167), .ZN(n20169) );
  INV_X1 U22965 ( .A(n21089), .ZN(n20802) );
  NOR2_X1 U22966 ( .A1(n504), .A2(n20173), .ZN(n20175) );
  NAND2_X1 U22967 ( .A1(n20786), .A2(n21932), .ZN(n20951) );
  NAND2_X1 U22968 ( .A1(n20494), .A2(n20179), .ZN(n20181) );
  NAND2_X1 U22969 ( .A1(n21090), .A2(n21089), .ZN(n20466) );
  NAND2_X1 U22970 ( .A1(n20191), .A2(n20539), .ZN(n20189) );
  INV_X1 U22971 ( .A(n20388), .ZN(n20541) );
  NAND2_X1 U22973 ( .A1(n28779), .A2(n20416), .ZN(n20823) );
  NAND2_X1 U22974 ( .A1(n20823), .A2(n20418), .ZN(n20195) );
  NAND2_X1 U22975 ( .A1(n20192), .A2(n20193), .ZN(n20821) );
  NAND2_X1 U22976 ( .A1(n20193), .A2(n20580), .ZN(n20194) );
  NOR2_X1 U22977 ( .A1(n20413), .A2(n20194), .ZN(n20824) );
  NAND2_X1 U22978 ( .A1(n21675), .A2(n21677), .ZN(n21447) );
  MUX2_X1 U22979 ( .A(n20585), .B(n20311), .S(n29144), .Z(n20198) );
  NOR2_X1 U22980 ( .A1(n20585), .A2(n20196), .ZN(n20586) );
  NOR2_X1 U22981 ( .A1(n20315), .A2(n20314), .ZN(n20197) );
  AND2_X1 U22982 ( .A1(n20199), .A2(n20201), .ZN(n20303) );
  OAI21_X1 U22983 ( .B1(n6935), .B2(n20202), .A(n416), .ZN(n20203) );
  OAI21_X1 U22985 ( .B1(n20558), .B2(n20208), .A(n20560), .ZN(n20211) );
  OAI21_X1 U22986 ( .B1(n20209), .B2(n20563), .A(n20562), .ZN(n20210) );
  OAI22_X1 U22989 ( .A1(n21448), .A2(n21678), .B1(n21677), .B2(n21676), .ZN(
        n21004) );
  XNOR2_X1 U22990 ( .A(n20215), .B(n20214), .ZN(n20280) );
  NAND3_X1 U22991 ( .A1(n29488), .A2(n20878), .A3(n20875), .ZN(n20216) );
  XNOR2_X1 U22992 ( .A(n28483), .B(n1193), .ZN(n20278) );
  INV_X1 U22993 ( .A(n21655), .ZN(n21074) );
  NAND2_X1 U22994 ( .A1(n20498), .A2(n20504), .ZN(n20229) );
  NAND2_X1 U22995 ( .A1(n20226), .A2(n20503), .ZN(n20228) );
  NAND2_X1 U22997 ( .A1(n20480), .A2(n20475), .ZN(n20231) );
  OAI211_X1 U22998 ( .C1(n21074), .C2(n6275), .A(n21442), .B(n21654), .ZN(
        n20246) );
  INV_X1 U22999 ( .A(n20511), .ZN(n20235) );
  AOI21_X1 U23000 ( .B1(n20345), .B2(n20235), .A(n20349), .ZN(n20234) );
  NOR2_X1 U23001 ( .A1(n20014), .A2(n20510), .ZN(n20233) );
  OAI22_X1 U23002 ( .A1(n20234), .A2(n20233), .B1(n20344), .B2(n20235), .ZN(
        n20237) );
  NAND3_X1 U23003 ( .A1(n20235), .A2(n20342), .A3(n20510), .ZN(n20236) );
  AND2_X2 U23004 ( .A1(n20237), .A2(n20236), .ZN(n21653) );
  INV_X1 U23005 ( .A(n21442), .ZN(n21661) );
  NAND2_X1 U23007 ( .A1(n20488), .A2(n28620), .ZN(n20243) );
  AOI21_X1 U23008 ( .B1(n20240), .B2(n29527), .A(n20239), .ZN(n20242) );
  NOR2_X1 U23011 ( .A1(n20635), .A2(n20637), .ZN(n20250) );
  NOR2_X1 U23012 ( .A1(n20247), .A2(n28538), .ZN(n20249) );
  MUX2_X1 U23013 ( .A(n20250), .B(n20249), .S(n20248), .Z(n20254) );
  OAI21_X1 U23014 ( .B1(n20636), .B2(n20453), .A(n20635), .ZN(n20251) );
  NOR2_X1 U23017 ( .A1(n22402), .A2(n21429), .ZN(n20271) );
  NOR2_X1 U23018 ( .A1(n20630), .A2(n20334), .ZN(n20259) );
  NAND2_X1 U23019 ( .A1(n28515), .A2(n20259), .ZN(n20260) );
  NAND2_X1 U23020 ( .A1(n19795), .A2(n21359), .ZN(n20329) );
  AOI21_X1 U23021 ( .B1(n20329), .B2(n20262), .A(n20520), .ZN(n20264) );
  INV_X1 U23022 ( .A(n21067), .ZN(n20270) );
  NOR2_X1 U23023 ( .A1(n22397), .A2(n22401), .ZN(n20269) );
  NAND2_X1 U23025 ( .A1(n28552), .A2(n6203), .ZN(n21062) );
  OAI21_X1 U23026 ( .B1(n21061), .B2(n21063), .A(n21062), .ZN(n20268) );
  NAND2_X1 U23027 ( .A1(n20268), .A2(n21065), .ZN(n21665) );
  NOR2_X1 U23028 ( .A1(n28408), .A2(n20275), .ZN(n21431) );
  NOR2_X2 U23029 ( .A1(n21432), .A2(n21431), .ZN(n22404) );
  XNOR2_X1 U23030 ( .A(n20277), .B(n20278), .ZN(n20279) );
  MUX2_X1 U23031 ( .A(n20283), .B(n28657), .S(n20281), .Z(n20288) );
  NOR2_X1 U23032 ( .A1(n20285), .A2(n20284), .ZN(n20287) );
  AND2_X1 U23033 ( .A1(n20289), .A2(n2152), .ZN(n20766) );
  NOR2_X2 U23034 ( .A1(n20767), .A2(n20766), .ZN(n21304) );
  NAND2_X1 U23035 ( .A1(n20290), .A2(n20293), .ZN(n20291) );
  NAND2_X1 U23036 ( .A1(n20292), .A2(n20291), .ZN(n20297) );
  AOI21_X1 U23037 ( .B1(n3247), .B2(n19901), .A(n20299), .ZN(n20300) );
  NAND2_X1 U23038 ( .A1(n20303), .A2(n20302), .ZN(n20309) );
  NAND3_X1 U23039 ( .A1(n20306), .A2(n20305), .A3(n20304), .ZN(n20308) );
  NOR2_X1 U23040 ( .A1(n20587), .A2(n29144), .ZN(n20313) );
  NOR2_X1 U23041 ( .A1(n20311), .A2(n20584), .ZN(n20312) );
  MUX2_X1 U23042 ( .A(n20313), .B(n20312), .S(n20589), .Z(n20318) );
  NAND2_X1 U23043 ( .A1(n20315), .A2(n20314), .ZN(n20316) );
  OAI22_X1 U23044 ( .A1(n20316), .A2(n20589), .B1(n20588), .B2(n20584), .ZN(
        n20317) );
  OAI21_X1 U23045 ( .B1(n21311), .B2(n21309), .A(n21307), .ZN(n20326) );
  NAND2_X1 U23046 ( .A1(n20326), .A2(n20771), .ZN(n20327) );
  NAND2_X1 U23048 ( .A1(n1881), .A2(n20334), .ZN(n20332) );
  OAI21_X1 U23050 ( .B1(n28515), .B2(n20332), .A(n20331), .ZN(n20337) );
  NAND2_X1 U23051 ( .A1(n20335), .A2(n20334), .ZN(n20336) );
  NOR2_X1 U23052 ( .A1(n21550), .A2(n21177), .ZN(n20365) );
  MUX2_X1 U23053 ( .A(n20503), .B(n20504), .S(n20499), .Z(n20338) );
  NOR2_X1 U23055 ( .A1(n20500), .A2(n20498), .ZN(n20340) );
  MUX2_X1 U23056 ( .A(n20343), .B(n20342), .S(n20344), .Z(n20350) );
  AOI21_X1 U23057 ( .B1(n20345), .B2(n20344), .A(n19785), .ZN(n20346) );
  OAI21_X1 U23058 ( .B1(n20350), .B2(n20349), .A(n20348), .ZN(n20351) );
  OAI21_X1 U23059 ( .B1(n21549), .B2(n21177), .A(n21553), .ZN(n20364) );
  NOR2_X1 U23060 ( .A1(n20783), .A2(n21177), .ZN(n21520) );
  AOI21_X1 U23061 ( .B1(n20353), .B2(n20352), .A(n4557), .ZN(n20357) );
  OAI22_X1 U23062 ( .A1(n20355), .A2(n20354), .B1(n20480), .B2(n382), .ZN(
        n20356) );
  INV_X1 U23063 ( .A(n20782), .ZN(n21547) );
  INV_X1 U23064 ( .A(n20484), .ZN(n20358) );
  OAI21_X1 U23065 ( .B1(n20488), .B2(n20483), .A(n20358), .ZN(n20360) );
  AOI22_X1 U23066 ( .A1(n20361), .A2(n20360), .B1(n20481), .B2(n20359), .ZN(
        n21519) );
  XNOR2_X1 U23068 ( .A(n22301), .B(n22472), .ZN(n20424) );
  INV_X1 U23069 ( .A(n20848), .ZN(n20366) );
  NOR2_X1 U23070 ( .A1(n20366), .A2(n21576), .ZN(n20370) );
  AND2_X1 U23071 ( .A1(n20749), .A2(n21483), .ZN(n20367) );
  AOI22_X1 U23072 ( .A1(n5142), .A2(n20368), .B1(n20367), .B2(n21575), .ZN(
        n20369) );
  OAI21_X1 U23073 ( .B1(n5142), .B2(n20370), .A(n20369), .ZN(n22116) );
  MUX2_X1 U23074 ( .A(n20372), .B(n20371), .S(n20373), .Z(n20380) );
  NOR2_X1 U23075 ( .A1(n20374), .A2(n20373), .ZN(n20376) );
  INV_X1 U23078 ( .A(n20571), .ZN(n20387) );
  OAI21_X1 U23079 ( .B1(n20567), .B2(n20381), .A(n20383), .ZN(n20386) );
  INV_X1 U23080 ( .A(n20567), .ZN(n20382) );
  NAND2_X1 U23082 ( .A1(n20383), .A2(n97), .ZN(n20384) );
  OAI21_X1 U23084 ( .B1(n29644), .B2(n20389), .A(n20388), .ZN(n20390) );
  NAND2_X1 U23085 ( .A1(n20390), .A2(n20547), .ZN(n20391) );
  NOR2_X1 U23088 ( .A1(n6086), .A2(n505), .ZN(n20411) );
  OAI21_X1 U23089 ( .B1(n20552), .B2(n28501), .A(n20404), .ZN(n20410) );
  MUX2_X1 U23090 ( .A(n20408), .B(n20407), .S(n20551), .Z(n20409) );
  OAI21_X1 U23092 ( .B1(n21504), .B2(n21499), .A(n21503), .ZN(n20422) );
  INV_X1 U23093 ( .A(n20412), .ZN(n20413) );
  INV_X1 U23094 ( .A(n20583), .ZN(n20415) );
  NAND2_X1 U23095 ( .A1(n20577), .A2(n20414), .ZN(n20939) );
  MUX2_X1 U23096 ( .A(n20415), .B(n20939), .S(n20941), .Z(n20776) );
  NAND2_X1 U23097 ( .A1(n20419), .A2(n20823), .ZN(n20777) );
  AOI21_X1 U23098 ( .B1(n20776), .B2(n20777), .A(n28619), .ZN(n20420) );
  OAI21_X1 U23099 ( .B1(n21192), .B2(n20420), .A(n21539), .ZN(n20421) );
  AND2_X1 U23100 ( .A1(n20422), .A2(n20421), .ZN(n21949) );
  INV_X1 U23101 ( .A(n21949), .ZN(n22327) );
  XNOR2_X1 U23102 ( .A(n22327), .B(n22116), .ZN(n20423) );
  XNOR2_X1 U23103 ( .A(n20423), .B(n20424), .ZN(n20472) );
  NOR2_X1 U23104 ( .A1(n22012), .A2(n20934), .ZN(n20427) );
  NOR2_X1 U23107 ( .A1(n20618), .A2(n20617), .ZN(n20429) );
  INV_X1 U23108 ( .A(n20435), .ZN(n20439) );
  NAND2_X1 U23109 ( .A1(n20607), .A2(n20440), .ZN(n20438) );
  INV_X1 U23110 ( .A(n20614), .ZN(n20436) );
  NOR2_X1 U23111 ( .A1(n21514), .A2(n21513), .ZN(n21531) );
  AND3_X1 U23112 ( .A1(n20444), .A2(n19901), .A3(n20443), .ZN(n20445) );
  NOR2_X1 U23113 ( .A1(n20446), .A2(n20445), .ZN(n20447) );
  OAI21_X1 U23114 ( .B1(n20448), .B2(n415), .A(n20447), .ZN(n21199) );
  INV_X1 U23115 ( .A(n21199), .ZN(n21516) );
  NOR2_X1 U23116 ( .A1(n21531), .A2(n21516), .ZN(n20465) );
  NAND2_X1 U23117 ( .A1(n20634), .A2(n20453), .ZN(n20454) );
  NOR2_X1 U23118 ( .A1(n21516), .A2(n21513), .ZN(n20462) );
  OR2_X1 U23119 ( .A1(n20597), .A2(n1916), .ZN(n20457) );
  OAI21_X1 U23121 ( .B1(n20463), .B2(n20462), .A(n21509), .ZN(n20464) );
  XNOR2_X1 U23123 ( .A(n22302), .B(n28162), .ZN(n22157) );
  AND2_X1 U23124 ( .A1(n20951), .A2(n20466), .ZN(n20469) );
  OAI21_X1 U23125 ( .B1(n20955), .B2(n20802), .A(n21090), .ZN(n20467) );
  NAND2_X1 U23126 ( .A1(n20467), .A2(n29586), .ZN(n20468) );
  OAI21_X2 U23127 ( .B1(n21934), .B2(n20469), .A(n20468), .ZN(n22601) );
  XNOR2_X1 U23128 ( .A(n22601), .B(n2403), .ZN(n20470) );
  MUX2_X1 U23129 ( .A(n20473), .B(n23136), .S(n23531), .Z(n20657) );
  NAND3_X1 U23130 ( .A1(n20480), .A2(n20479), .A3(n20478), .ZN(n21330) );
  NAND2_X1 U23131 ( .A1(n20482), .A2(n20481), .ZN(n21610) );
  MUX2_X1 U23132 ( .A(n28620), .B(n20486), .S(n20483), .Z(n20489) );
  NOR3_X1 U23133 ( .A1(n20486), .A2(n20485), .A3(n20484), .ZN(n20487) );
  NAND2_X1 U23134 ( .A1(n20496), .A2(n20494), .ZN(n20490) );
  AOI21_X1 U23135 ( .B1(n20491), .B2(n20490), .A(n499), .ZN(n20492) );
  AOI21_X1 U23136 ( .B1(n20503), .B2(n20498), .A(n20504), .ZN(n20502) );
  NAND2_X1 U23137 ( .A1(n20500), .A2(n20499), .ZN(n20501) );
  NAND2_X1 U23138 ( .A1(n20502), .A2(n20501), .ZN(n20508) );
  NAND3_X1 U23139 ( .A1(n1624), .A2(n20504), .A3(n20503), .ZN(n20507) );
  OAI211_X1 U23140 ( .C1(n20511), .C2(n19785), .A(n20510), .B(n20509), .ZN(
        n20512) );
  NAND3_X1 U23142 ( .A1(n21610), .A2(n21611), .A3(n21612), .ZN(n20515) );
  NAND2_X1 U23143 ( .A1(n21618), .A2(n20515), .ZN(n20516) );
  NAND2_X1 U23144 ( .A1(n21619), .A2(n20516), .ZN(n20524) );
  NOR2_X1 U23145 ( .A1(n28610), .A2(n28586), .ZN(n20521) );
  AOI22_X1 U23146 ( .A1(n20521), .A2(n20520), .B1(n28133), .B2(n501), .ZN(
        n20522) );
  NAND2_X1 U23147 ( .A1(n21326), .A2(n21334), .ZN(n20523) );
  NOR2_X1 U23148 ( .A1(n20744), .A2(n21159), .ZN(n20531) );
  INV_X1 U23149 ( .A(n21159), .ZN(n20526) );
  NAND3_X1 U23150 ( .A1(n20526), .A2(n21157), .A3(n21155), .ZN(n20529) );
  INV_X1 U23151 ( .A(n20527), .ZN(n20528) );
  XNOR2_X1 U23153 ( .A(n22750), .B(n22609), .ZN(n22714) );
  INV_X1 U23154 ( .A(n20532), .ZN(n22011) );
  AND2_X1 U23155 ( .A1(n22011), .A2(n22013), .ZN(n20537) );
  NOR2_X1 U23156 ( .A1(n20933), .A2(n21078), .ZN(n20535) );
  NAND2_X1 U23157 ( .A1(n22011), .A2(n20533), .ZN(n20534) );
  MUX2_X1 U23160 ( .A(n20546), .B(n20547), .S(n29644), .Z(n20543) );
  NOR2_X1 U23161 ( .A1(n6261), .A2(n20539), .ZN(n20542) );
  INV_X1 U23162 ( .A(n20544), .ZN(n20545) );
  NOR2_X1 U23163 ( .A1(n21586), .A2(n21585), .ZN(n20889) );
  NAND2_X1 U23164 ( .A1(n20553), .A2(n20549), .ZN(n20550) );
  NAND3_X1 U23165 ( .A1(n20554), .A2(n20553), .A3(n20552), .ZN(n20555) );
  INV_X1 U23166 ( .A(n20559), .ZN(n20565) );
  OAI21_X1 U23167 ( .B1(n20563), .B2(n20562), .A(n20561), .ZN(n20564) );
  NAND2_X1 U23168 ( .A1(n6932), .A2(n97), .ZN(n20572) );
  NAND2_X1 U23169 ( .A1(n20574), .A2(n28508), .ZN(n20713) );
  NOR2_X1 U23170 ( .A1(n28779), .A2(n20941), .ZN(n20579) );
  INV_X1 U23171 ( .A(n21585), .ZN(n20591) );
  NOR2_X1 U23172 ( .A1(n3789), .A2(n21322), .ZN(n20593) );
  OAI21_X1 U23173 ( .B1(n20591), .B2(n21322), .A(n20886), .ZN(n20592) );
  NOR3_X1 U23174 ( .A1(n20594), .A2(n20593), .A3(n20592), .ZN(n20595) );
  NAND2_X1 U23178 ( .A1(n20601), .A2(n20597), .ZN(n20599) );
  MUX2_X1 U23179 ( .A(n20600), .B(n20599), .S(n28408), .Z(n20606) );
  NOR3_X1 U23180 ( .A1(n20601), .A2(n4569), .A3(n1915), .ZN(n20602) );
  AOI21_X1 U23181 ( .B1(n20604), .B2(n20603), .A(n20602), .ZN(n20605) );
  INV_X1 U23182 ( .A(n21599), .ZN(n21603) );
  AOI22_X1 U23183 ( .A1(n20609), .A2(n20611), .B1(n20608), .B2(n20607), .ZN(
        n20615) );
  NAND3_X1 U23184 ( .A1(n20614), .A2(n20611), .A3(n29625), .ZN(n20613) );
  INV_X1 U23185 ( .A(n21600), .ZN(n20720) );
  AND2_X1 U23186 ( .A1(n20617), .A2(n20616), .ZN(n20621) );
  MUX2_X1 U23187 ( .A(n20618), .B(n6567), .S(n20617), .Z(n20620) );
  INV_X1 U23188 ( .A(n20722), .ZN(n21316) );
  NOR2_X1 U23189 ( .A1(n1881), .A2(n20626), .ZN(n20627) );
  NAND2_X1 U23190 ( .A1(n20628), .A2(n20627), .ZN(n20629) );
  NAND2_X1 U23191 ( .A1(n21316), .A2(n21601), .ZN(n21138) );
  INV_X1 U23192 ( .A(n21138), .ZN(n20643) );
  INV_X1 U23193 ( .A(n28538), .ZN(n20642) );
  OAI21_X1 U23194 ( .B1(n20637), .B2(n20636), .A(n20635), .ZN(n20638) );
  OAI21_X1 U23195 ( .B1(n20642), .B2(n20641), .A(n20640), .ZN(n21314) );
  INV_X1 U23196 ( .A(n21314), .ZN(n21605) );
  NAND2_X1 U23197 ( .A1(n21314), .A2(n21601), .ZN(n20649) );
  NAND2_X1 U23198 ( .A1(n21308), .A2(n29531), .ZN(n21150) );
  XNOR2_X1 U23199 ( .A(n22681), .B(n22240), .ZN(n20655) );
  OAI21_X1 U23200 ( .B1(n21119), .B2(n21140), .A(n21143), .ZN(n20653) );
  NAND2_X1 U23201 ( .A1(n21141), .A2(n20650), .ZN(n20652) );
  NOR2_X1 U23202 ( .A1(n20851), .A2(n21118), .ZN(n20651) );
  AOI21_X2 U23203 ( .B1(n20652), .B2(n20653), .A(n20651), .ZN(n22855) );
  XNOR2_X1 U23204 ( .A(n22855), .B(n1079), .ZN(n20654) );
  XNOR2_X1 U23206 ( .A(n22227), .B(n3334), .ZN(n20660) );
  XNOR2_X1 U23207 ( .A(n20660), .B(n22773), .ZN(n20665) );
  OAI21_X1 U23210 ( .B1(n21472), .B2(n21473), .A(n21731), .ZN(n20661) );
  MUX2_X2 U23211 ( .A(n20662), .B(n20661), .S(n21471), .Z(n22697) );
  XNOR2_X1 U23212 ( .A(n22697), .B(n22882), .ZN(n20664) );
  XNOR2_X1 U23213 ( .A(n20665), .B(n20664), .ZN(n20682) );
  MUX2_X1 U23214 ( .A(n22286), .B(n22026), .S(n22023), .Z(n20667) );
  INV_X1 U23215 ( .A(n22286), .ZN(n22291) );
  NAND2_X1 U23218 ( .A1(n22286), .A2(n22290), .ZN(n21208) );
  NAND2_X1 U23220 ( .A1(n20668), .A2(n22294), .ZN(n22879) );
  INV_X1 U23221 ( .A(n22879), .ZN(n21848) );
  NOR2_X1 U23222 ( .A1(n21394), .A2(n21632), .ZN(n20679) );
  INV_X1 U23223 ( .A(n20669), .ZN(n20673) );
  NOR2_X1 U23224 ( .A1(n20671), .A2(n20670), .ZN(n20672) );
  NAND2_X1 U23225 ( .A1(n20673), .A2(n20672), .ZN(n20674) );
  OAI21_X1 U23226 ( .B1(n20675), .B2(n20674), .A(n21638), .ZN(n20678) );
  NAND2_X1 U23227 ( .A1(n21637), .A2(n21392), .ZN(n21226) );
  NAND2_X1 U23228 ( .A1(n21632), .A2(n21227), .ZN(n21393) );
  NAND2_X1 U23229 ( .A1(n21226), .A2(n21393), .ZN(n20676) );
  NAND2_X1 U23230 ( .A1(n20676), .A2(n21631), .ZN(n20677) );
  OAI21_X1 U23231 ( .B1(n20679), .B2(n20678), .A(n20677), .ZN(n22226) );
  INV_X1 U23232 ( .A(n22226), .ZN(n22073) );
  XNOR2_X1 U23233 ( .A(n21848), .B(n20680), .ZN(n20681) );
  INV_X1 U23234 ( .A(n22568), .ZN(n21841) );
  OAI21_X1 U23235 ( .B1(n29227), .B2(n6934), .A(n29526), .ZN(n20684) );
  AOI22_X1 U23236 ( .A1(n21704), .A2(n21273), .B1(n6934), .B2(n21703), .ZN(
        n20683) );
  NAND2_X1 U23237 ( .A1(n20684), .A2(n20683), .ZN(n22821) );
  XNOR2_X1 U23238 ( .A(n21841), .B(n22821), .ZN(n20687) );
  INV_X1 U23239 ( .A(n21287), .ZN(n20726) );
  NOR2_X1 U23240 ( .A1(n21288), .A2(n21291), .ZN(n20989) );
  OAI211_X1 U23241 ( .C1(n20914), .C2(n29313), .A(n21287), .B(n21292), .ZN(
        n20685) );
  XNOR2_X1 U23242 ( .A(n22890), .B(n3527), .ZN(n20686) );
  XNOR2_X1 U23243 ( .A(n20687), .B(n20686), .ZN(n20709) );
  OAI21_X1 U23244 ( .B1(n20688), .B2(n20689), .A(n5772), .ZN(n20975) );
  INV_X1 U23245 ( .A(n20975), .ZN(n21261) );
  INV_X1 U23246 ( .A(n20688), .ZN(n20691) );
  NOR2_X1 U23247 ( .A1(n20689), .A2(n21364), .ZN(n20690) );
  INV_X1 U23248 ( .A(n21717), .ZN(n21260) );
  NOR2_X1 U23249 ( .A1(n21714), .A2(n21713), .ZN(n21263) );
  OAI21_X1 U23250 ( .B1(n21260), .B2(n21258), .A(n21263), .ZN(n20692) );
  NAND2_X1 U23251 ( .A1(n21809), .A2(n21810), .ZN(n20699) );
  NAND2_X1 U23252 ( .A1(n20694), .A2(n20693), .ZN(n21250) );
  INV_X1 U23253 ( .A(n21250), .ZN(n20695) );
  INV_X1 U23254 ( .A(n21254), .ZN(n20696) );
  INV_X1 U23255 ( .A(n21806), .ZN(n21379) );
  AOI21_X1 U23256 ( .B1(n20696), .B2(n21379), .A(n21253), .ZN(n20697) );
  XNOR2_X1 U23257 ( .A(n22796), .B(n1858), .ZN(n22249) );
  NOR2_X1 U23258 ( .A1(n21346), .A2(n21343), .ZN(n21691) );
  NOR2_X1 U23261 ( .A1(n21695), .A2(n21242), .ZN(n20700) );
  INV_X1 U23262 ( .A(n21696), .ZN(n21348) );
  NOR2_X1 U23263 ( .A1(n20702), .A2(n20701), .ZN(n20969) );
  NAND2_X1 U23264 ( .A1(n20969), .A2(n20704), .ZN(n20707) );
  OAI21_X1 U23265 ( .B1(n20703), .B2(n381), .A(n21217), .ZN(n20706) );
  INV_X1 U23266 ( .A(n21218), .ZN(n20967) );
  XNOR2_X1 U23267 ( .A(n22798), .B(n22248), .ZN(n22486) );
  XOR2_X1 U23268 ( .A(n22249), .B(n22486), .Z(n20708) );
  INV_X1 U23269 ( .A(n20875), .ZN(n20710) );
  OAI21_X1 U23270 ( .B1(n21268), .B2(n20710), .A(n20878), .ZN(n20712) );
  NAND3_X1 U23271 ( .A1(n20816), .A2(n20878), .A3(n20875), .ZN(n20711) );
  XNOR2_X1 U23272 ( .A(n22327), .B(n22913), .ZN(n21838) );
  INV_X1 U23273 ( .A(n21591), .ZN(n20717) );
  AND2_X1 U23274 ( .A1(n21322), .A2(n5983), .ZN(n20716) );
  OAI21_X1 U23275 ( .B1(n20717), .B2(n20716), .A(n28584), .ZN(n20718) );
  AND2_X1 U23276 ( .A1(n21086), .A2(n21426), .ZN(n20719) );
  XNOR2_X1 U23277 ( .A(n22232), .B(n22759), .ZN(n22474) );
  XNOR2_X1 U23278 ( .A(n22474), .B(n21838), .ZN(n20735) );
  AOI21_X1 U23279 ( .B1(n21599), .B2(n20721), .A(n20720), .ZN(n20725) );
  NAND2_X1 U23280 ( .A1(n21598), .A2(n21601), .ZN(n20724) );
  NAND2_X1 U23281 ( .A1(n20916), .A2(n20726), .ZN(n20728) );
  INV_X1 U23282 ( .A(n20917), .ZN(n20727) );
  XNOR2_X1 U23283 ( .A(n22845), .B(n22762), .ZN(n22358) );
  NAND3_X1 U23287 ( .A1(n21326), .A2(n21327), .A3(n21612), .ZN(n20730) );
  XNOR2_X1 U23289 ( .A(n22763), .B(n2987), .ZN(n20733) );
  XNOR2_X1 U23290 ( .A(n22358), .B(n20733), .ZN(n20734) );
  INV_X1 U23291 ( .A(n20736), .ZN(n20738) );
  NAND2_X1 U23292 ( .A1(n20738), .A2(n20737), .ZN(n20742) );
  INV_X1 U23293 ( .A(n20739), .ZN(n20740) );
  NOR3_X1 U23294 ( .A1(n20742), .A2(n20741), .A3(n20740), .ZN(n20743) );
  NAND2_X1 U23295 ( .A1(n494), .A2(n21155), .ZN(n20745) );
  AOI21_X1 U23296 ( .B1(n20746), .B2(n20745), .A(n4960), .ZN(n20747) );
  NOR2_X2 U23297 ( .A1(n20748), .A2(n20747), .ZN(n22812) );
  INV_X1 U23298 ( .A(n22437), .ZN(n20750) );
  XNOR2_X1 U23299 ( .A(n20750), .B(n22812), .ZN(n20753) );
  NOR2_X1 U23300 ( .A1(n28789), .A2(n6752), .ZN(n20751) );
  AOI21_X1 U23301 ( .B1(n2037), .B2(n1946), .A(n21496), .ZN(n20752) );
  XNOR2_X1 U23302 ( .A(n22898), .B(n22245), .ZN(n22688) );
  XNOR2_X1 U23303 ( .A(n22688), .B(n20753), .ZN(n20761) );
  XNOR2_X1 U23304 ( .A(n21728), .B(n22330), .ZN(n20759) );
  XNOR2_X1 U23305 ( .A(n22778), .B(n135), .ZN(n20758) );
  XNOR2_X1 U23306 ( .A(n20759), .B(n20758), .ZN(n20760) );
  NOR2_X1 U23307 ( .A1(n20762), .A2(n4828), .ZN(n20764) );
  NOR3_X1 U23308 ( .A1(n22012), .A2(n22011), .A3(n22013), .ZN(n20763) );
  NOR3_X1 U23309 ( .A1(n22014), .A2(n20764), .A3(n20763), .ZN(n20765) );
  XNOR2_X1 U23310 ( .A(n20765), .B(n28499), .ZN(n21856) );
  INV_X1 U23312 ( .A(n21308), .ZN(n20769) );
  NOR2_X1 U23313 ( .A1(n20769), .A2(n29530), .ZN(n21305) );
  NOR2_X1 U23314 ( .A1(n21153), .A2(n21305), .ZN(n20775) );
  NAND2_X1 U23315 ( .A1(n20938), .A2(n21306), .ZN(n20770) );
  NAND2_X1 U23316 ( .A1(n21308), .A2(n20770), .ZN(n20772) );
  INV_X1 U23317 ( .A(n21500), .ZN(n21543) );
  AOI21_X1 U23319 ( .B1(n21500), .B2(n21539), .A(n21192), .ZN(n20778) );
  INV_X1 U23320 ( .A(n21539), .ZN(n20945) );
  INV_X1 U23321 ( .A(n28619), .ZN(n20948) );
  OAI21_X1 U23322 ( .B1(n20945), .B2(n20948), .A(n21192), .ZN(n20781) );
  INV_X1 U23323 ( .A(n21503), .ZN(n21540) );
  NOR3_X1 U23324 ( .A1(n21540), .A2(n21539), .A3(n28185), .ZN(n20780) );
  XNOR2_X1 U23325 ( .A(n20885), .B(n22219), .ZN(n22461) );
  INV_X1 U23327 ( .A(n22792), .ZN(n22086) );
  XNOR2_X1 U23328 ( .A(n22086), .B(n2961), .ZN(n20797) );
  NOR2_X1 U23329 ( .A1(n21930), .A2(n21932), .ZN(n20785) );
  NAND2_X1 U23330 ( .A1(n20785), .A2(n20954), .ZN(n20791) );
  INV_X1 U23331 ( .A(n20801), .ZN(n20788) );
  NOR2_X1 U23332 ( .A1(n21932), .A2(n21097), .ZN(n20787) );
  AOI22_X1 U23333 ( .A1(n20788), .A2(n21932), .B1(n20787), .B2(n20786), .ZN(
        n20790) );
  INV_X1 U23334 ( .A(n21513), .ZN(n21512) );
  NAND3_X1 U23335 ( .A1(n21534), .A2(n21530), .A3(n21509), .ZN(n20795) );
  INV_X1 U23336 ( .A(n21514), .ZN(n21533) );
  NAND3_X1 U23337 ( .A1(n21533), .A2(n21199), .A3(n21532), .ZN(n20794) );
  XNOR2_X1 U23338 ( .A(n22790), .B(n22835), .ZN(n22383) );
  NAND2_X1 U23339 ( .A1(n23353), .A2(n4231), .ZN(n20840) );
  INV_X1 U23340 ( .A(n20798), .ZN(n22340) );
  INV_X1 U23341 ( .A(n20954), .ZN(n20800) );
  XNOR2_X1 U23342 ( .A(n22340), .B(n22903), .ZN(n20813) );
  NAND2_X1 U23343 ( .A1(n20899), .A2(n21424), .ZN(n20808) );
  NAND2_X1 U23344 ( .A1(n21087), .A2(n21425), .ZN(n20806) );
  OAI21_X1 U23345 ( .B1(n28602), .B2(n20808), .A(n20807), .ZN(n22553) );
  INV_X1 U23346 ( .A(n21665), .ZN(n21015) );
  NAND3_X1 U23347 ( .A1(n22404), .A2(n21662), .A3(n22401), .ZN(n20811) );
  INV_X1 U23348 ( .A(n21018), .ZN(n20809) );
  NAND2_X1 U23349 ( .A1(n22402), .A2(n20809), .ZN(n20810) );
  AND3_X1 U23350 ( .A1(n20812), .A2(n20811), .A3(n20810), .ZN(n21805) );
  INV_X1 U23351 ( .A(n21805), .ZN(n22066) );
  XNOR2_X1 U23352 ( .A(n22066), .B(n22553), .ZN(n22748) );
  XNOR2_X1 U23353 ( .A(n20813), .B(n22748), .ZN(n20839) );
  NOR2_X1 U23354 ( .A1(n29488), .A2(n20816), .ZN(n20815) );
  INV_X1 U23355 ( .A(n20816), .ZN(n20874) );
  NAND3_X1 U23356 ( .A1(n21268), .A2(n20874), .A3(n20875), .ZN(n20817) );
  NAND2_X1 U23357 ( .A1(n21272), .A2(n20817), .ZN(n20820) );
  INV_X1 U23358 ( .A(n20878), .ZN(n21267) );
  AOI21_X1 U23359 ( .B1(n20818), .B2(n21267), .A(n21268), .ZN(n20819) );
  INV_X1 U23360 ( .A(n21676), .ZN(n21673) );
  INV_X1 U23361 ( .A(n20821), .ZN(n20822) );
  NOR2_X1 U23362 ( .A1(n20823), .A2(n20822), .ZN(n20828) );
  INV_X1 U23363 ( .A(n20824), .ZN(n20825) );
  NAND2_X1 U23364 ( .A1(n20825), .A2(n20418), .ZN(n20827) );
  OAI21_X1 U23365 ( .B1(n20828), .B2(n20827), .A(n28215), .ZN(n20829) );
  XNOR2_X1 U23366 ( .A(n22718), .B(n22426), .ZN(n22497) );
  INV_X1 U23367 ( .A(n21653), .ZN(n21660) );
  XNOR2_X1 U23371 ( .A(n22497), .B(n20837), .ZN(n20838) );
  NAND3_X1 U23372 ( .A1(n21125), .A2(n21458), .A3(n21567), .ZN(n20845) );
  XNOR2_X1 U23373 ( .A(n22703), .B(n22033), .ZN(n20850) );
  XNOR2_X1 U23374 ( .A(n22773), .B(n20850), .ZN(n20873) );
  INV_X1 U23375 ( .A(n21118), .ZN(n20854) );
  MUX2_X1 U23376 ( .A(n20854), .B(n20851), .S(n21119), .Z(n20856) );
  OAI21_X1 U23378 ( .B1(n494), .B2(n20858), .A(n20857), .ZN(n20859) );
  AOI21_X1 U23379 ( .B1(n21158), .B2(n20858), .A(n20859), .ZN(n20860) );
  XNOR2_X1 U23380 ( .A(n22670), .B(n22526), .ZN(n21339) );
  XNOR2_X1 U23381 ( .A(n22387), .B(n3081), .ZN(n20870) );
  MUX2_X1 U23382 ( .A(n21497), .B(n21495), .S(n20864), .Z(n20869) );
  NOR2_X1 U23383 ( .A1(n28789), .A2(n21496), .ZN(n20866) );
  XNOR2_X1 U23386 ( .A(n20870), .B(n22523), .ZN(n20871) );
  XNOR2_X1 U23387 ( .A(n20871), .B(n21339), .ZN(n20872) );
  OR3_X1 U23388 ( .A1(n21269), .A2(n20874), .A3(n21266), .ZN(n20884) );
  NAND3_X1 U23389 ( .A1(n21269), .A2(n21268), .A3(n20878), .ZN(n20883) );
  NOR2_X1 U23390 ( .A1(n20876), .A2(n20875), .ZN(n20881) );
  NOR2_X1 U23391 ( .A1(n21268), .A2(n21267), .ZN(n20880) );
  INV_X1 U23392 ( .A(n20890), .ZN(n20893) );
  INV_X1 U23393 ( .A(n20891), .ZN(n20892) );
  NOR4_X1 U23394 ( .A1(n20898), .A2(n20897), .A3(n20893), .A4(n20892), .ZN(
        n20894) );
  NAND2_X1 U23395 ( .A1(n1925), .A2(n21085), .ZN(n20901) );
  NOR3_X1 U23396 ( .A1(n20898), .A2(n20897), .A3(n21424), .ZN(n21084) );
  INV_X1 U23397 ( .A(n20899), .ZN(n20900) );
  XNOR2_X1 U23398 ( .A(n21760), .B(n22545), .ZN(n20925) );
  OAI21_X1 U23399 ( .B1(n28442), .B2(n21600), .A(n21316), .ZN(n20904) );
  INV_X1 U23400 ( .A(n21601), .ZN(n21315) );
  NOR2_X1 U23401 ( .A1(n21598), .A2(n21601), .ZN(n21320) );
  INV_X1 U23402 ( .A(n21320), .ZN(n20902) );
  OAI211_X1 U23403 ( .C1(n20905), .C2(n21315), .A(n1941), .B(n20902), .ZN(
        n20903) );
  INV_X1 U23405 ( .A(n20906), .ZN(n20908) );
  NOR2_X1 U23406 ( .A1(n20908), .A2(n20907), .ZN(n20912) );
  INV_X1 U23407 ( .A(n21334), .ZN(n21607) );
  INV_X1 U23408 ( .A(n21612), .ZN(n21609) );
  AOI22_X1 U23409 ( .A1(n20910), .A2(n21163), .B1(n20909), .B2(n21609), .ZN(
        n20911) );
  NAND2_X1 U23410 ( .A1(n20915), .A2(n20914), .ZN(n20920) );
  NAND3_X1 U23411 ( .A1(n21292), .A2(n20916), .A3(n20986), .ZN(n20919) );
  NAND4_X2 U23412 ( .A1(n20918), .A2(n20921), .A3(n20920), .A4(n20919), .ZN(
        n22664) );
  XNOR2_X1 U23413 ( .A(n22664), .B(n27298), .ZN(n20922) );
  XNOR2_X1 U23414 ( .A(n20923), .B(n20922), .ZN(n20924) );
  XNOR2_X1 U23415 ( .A(n20925), .B(n20924), .ZN(n23167) );
  NOR2_X1 U23416 ( .A1(n28457), .A2(n23167), .ZN(n21027) );
  MUX2_X1 U23417 ( .A(n21530), .B(n21514), .S(n21513), .Z(n20928) );
  NAND2_X1 U23419 ( .A1(n21516), .A2(n21514), .ZN(n20926) );
  MUX2_X1 U23420 ( .A(n21535), .B(n20926), .S(n21530), .Z(n20927) );
  NAND2_X1 U23421 ( .A1(n20931), .A2(n21549), .ZN(n20929) );
  INV_X1 U23422 ( .A(n22689), .ZN(n20937) );
  INV_X1 U23423 ( .A(n20934), .ZN(n20935) );
  XNOR2_X1 U23424 ( .A(n22897), .B(n22437), .ZN(n20936) );
  XNOR2_X1 U23425 ( .A(n20937), .B(n20936), .ZN(n20960) );
  INV_X1 U23426 ( .A(n21192), .ZN(n21538) );
  NAND2_X1 U23427 ( .A1(n21500), .A2(n28611), .ZN(n20950) );
  INV_X1 U23429 ( .A(n20939), .ZN(n20942) );
  NOR2_X1 U23430 ( .A1(n503), .A2(n20941), .ZN(n20940) );
  AOI22_X1 U23431 ( .A1(n20942), .A2(n20941), .B1(n20940), .B2(n20413), .ZN(
        n20943) );
  NAND2_X1 U23432 ( .A1(n20777), .A2(n20943), .ZN(n20944) );
  NOR3_X1 U23436 ( .A1(n20954), .A2(n28916), .A3(n20953), .ZN(n20956) );
  XNOR2_X1 U23437 ( .A(n22811), .B(n730), .ZN(n20958) );
  XNOR2_X1 U23438 ( .A(n22502), .B(n20958), .ZN(n20959) );
  NAND2_X1 U23441 ( .A1(n21347), .A2(n20961), .ZN(n20965) );
  NOR3_X1 U23442 ( .A1(n3260), .A2(n28440), .A3(n21692), .ZN(n20964) );
  NOR3_X2 U23443 ( .A1(n20965), .A2(n20964), .A3(n20963), .ZN(n22338) );
  NOR2_X1 U23444 ( .A1(n20999), .A2(n21221), .ZN(n20971) );
  OAI21_X1 U23445 ( .B1(n20969), .B2(n20968), .A(n20967), .ZN(n20970) );
  OAI21_X1 U23446 ( .B1(n20972), .B2(n20971), .A(n20970), .ZN(n22717) );
  XNOR2_X1 U23447 ( .A(n29562), .B(n3134), .ZN(n20973) );
  XNOR2_X1 U23448 ( .A(n22519), .B(n20973), .ZN(n20997) );
  NAND2_X1 U23449 ( .A1(n21713), .A2(n20976), .ZN(n20974) );
  AOI21_X1 U23450 ( .B1(n20975), .B2(n20974), .A(n21260), .ZN(n20979) );
  OAI22_X1 U23451 ( .A1(n20977), .A2(n21717), .B1(n20976), .B2(n21712), .ZN(
        n20978) );
  NOR2_X1 U23452 ( .A1(n20979), .A2(n20978), .ZN(n22104) );
  INV_X1 U23454 ( .A(n21811), .ZN(n20982) );
  NOR2_X1 U23455 ( .A1(n21809), .A2(n21806), .ZN(n21380) );
  INV_X1 U23456 ( .A(n21380), .ZN(n20984) );
  XNOR2_X1 U23457 ( .A(n22713), .B(n29591), .ZN(n20995) );
  NOR2_X1 U23458 ( .A1(n20988), .A2(n21291), .ZN(n20987) );
  OAI21_X1 U23459 ( .B1(n20987), .B2(n20986), .A(n20985), .ZN(n20991) );
  OAI21_X1 U23460 ( .B1(n20989), .B2(n6911), .A(n20988), .ZN(n20990) );
  INV_X1 U23461 ( .A(n21703), .ZN(n20992) );
  NAND2_X1 U23462 ( .A1(n20992), .A2(n29526), .ZN(n21281) );
  INV_X1 U23463 ( .A(n21372), .ZN(n21702) );
  NAND3_X1 U23464 ( .A1(n21705), .A2(n20992), .A3(n21372), .ZN(n20993) );
  XNOR2_X1 U23465 ( .A(n22006), .B(n22856), .ZN(n21470) );
  XNOR2_X1 U23466 ( .A(n21470), .B(n20995), .ZN(n20996) );
  XNOR2_X1 U23467 ( .A(n20996), .B(n20997), .ZN(n23168) );
  NOR2_X1 U23468 ( .A1(n23683), .A2(n23168), .ZN(n21026) );
  NAND2_X1 U23469 ( .A1(n20998), .A2(n21221), .ZN(n21003) );
  INV_X1 U23470 ( .A(n20999), .ZN(n21002) );
  NAND3_X1 U23471 ( .A1(n21221), .A2(n21000), .A3(n21218), .ZN(n21001) );
  XNOR2_X1 U23472 ( .A(n22759), .B(n22912), .ZN(n21766) );
  INV_X1 U23473 ( .A(n21004), .ZN(n21006) );
  NOR2_X1 U23474 ( .A1(n21675), .A2(n21677), .ZN(n21079) );
  OAI21_X1 U23475 ( .B1(n21079), .B2(n21676), .A(n21448), .ZN(n21005) );
  AND2_X1 U23476 ( .A1(n21808), .A2(n19732), .ZN(n21011) );
  NOR2_X1 U23477 ( .A1(n19732), .A2(n21806), .ZN(n21010) );
  INV_X1 U23478 ( .A(n21810), .ZN(n21008) );
  NAND3_X1 U23479 ( .A1(n21811), .A2(n21008), .A3(n21379), .ZN(n21009) );
  XNOR2_X1 U23480 ( .A(n22910), .B(n22734), .ZN(n22532) );
  XNOR2_X1 U23481 ( .A(n22532), .B(n21766), .ZN(n21025) );
  XNOR2_X1 U23482 ( .A(n22731), .B(n22735), .ZN(n21023) );
  OAI21_X1 U23483 ( .B1(n22291), .B2(n29364), .A(n21213), .ZN(n21021) );
  INV_X1 U23484 ( .A(n22290), .ZN(n21019) );
  INV_X1 U23485 ( .A(n21917), .ZN(n22844) );
  XNOR2_X1 U23486 ( .A(n22844), .B(n3423), .ZN(n21022) );
  XNOR2_X1 U23487 ( .A(n21023), .B(n21022), .ZN(n21024) );
  XNOR2_X2 U23488 ( .A(n21025), .B(n21024), .ZN(n23016) );
  INV_X1 U23490 ( .A(n23168), .ZN(n23682) );
  NOR2_X1 U23491 ( .A1(n22140), .A2(n22139), .ZN(n21106) );
  NOR2_X1 U23492 ( .A1(n21030), .A2(n5339), .ZN(n21031) );
  NAND2_X1 U23493 ( .A1(n21736), .A2(n21389), .ZN(n21033) );
  XNOR2_X1 U23494 ( .A(n22271), .B(n22888), .ZN(n22511) );
  XNOR2_X1 U23495 ( .A(n22798), .B(n3586), .ZN(n21035) );
  XNOR2_X1 U23496 ( .A(n22511), .B(n21035), .ZN(n21057) );
  NOR2_X1 U23497 ( .A1(n21639), .A2(n21036), .ZN(n21038) );
  NAND2_X1 U23498 ( .A1(n21227), .A2(n21392), .ZN(n21395) );
  NAND2_X1 U23499 ( .A1(n21395), .A2(n21638), .ZN(n21037) );
  INV_X1 U23500 ( .A(n21040), .ZN(n21041) );
  NAND2_X1 U23501 ( .A1(n21041), .A2(n21400), .ZN(n21045) );
  NAND3_X1 U23502 ( .A1(n21042), .A2(n21402), .A3(n21750), .ZN(n21044) );
  NAND2_X1 U23503 ( .A1(n21410), .A2(n21409), .ZN(n21051) );
  AND2_X1 U23505 ( .A1(n21408), .A2(n21171), .ZN(n21413) );
  NAND2_X1 U23507 ( .A1(n21053), .A2(n21187), .ZN(n21054) );
  NAND2_X1 U23508 ( .A1(n21055), .A2(n21054), .ZN(n22509) );
  XNOR2_X1 U23509 ( .A(n22820), .B(n22509), .ZN(n21525) );
  XNOR2_X1 U23510 ( .A(n22727), .B(n21525), .ZN(n21056) );
  NAND2_X1 U23511 ( .A1(n23679), .A2(n23168), .ZN(n21058) );
  NOR2_X2 U23513 ( .A1(n21060), .A2(n21059), .ZN(n24617) );
  NAND2_X1 U23515 ( .A1(n21061), .A2(n21062), .ZN(n21066) );
  NAND2_X1 U23516 ( .A1(n21063), .A2(n21062), .ZN(n21064) );
  INV_X1 U23517 ( .A(n21663), .ZN(n21433) );
  AND2_X1 U23518 ( .A1(n21433), .A2(n22401), .ZN(n21068) );
  NAND2_X1 U23519 ( .A1(n22404), .A2(n21067), .ZN(n22403) );
  NAND2_X1 U23520 ( .A1(n21656), .A2(n21657), .ZN(n21075) );
  NAND3_X1 U23521 ( .A1(n21654), .A2(n6275), .A3(n21012), .ZN(n21072) );
  NAND2_X1 U23522 ( .A1(n20833), .A2(n21657), .ZN(n21071) );
  AND2_X1 U23523 ( .A1(n21077), .A2(n21076), .ZN(n21819) );
  XNOR2_X1 U23524 ( .A(n21847), .B(n22594), .ZN(n21105) );
  INV_X1 U23525 ( .A(n21079), .ZN(n21082) );
  AOI21_X1 U23526 ( .B1(n21675), .B2(n21673), .A(n21678), .ZN(n21081) );
  INV_X1 U23527 ( .A(n21448), .ZN(n21680) );
  XNOR2_X1 U23528 ( .A(n22199), .B(n2986), .ZN(n21083) );
  OAI211_X1 U23529 ( .C1(n21087), .C2(n21425), .A(n21424), .B(n21086), .ZN(
        n21088) );
  AOI21_X1 U23530 ( .B1(n4877), .B2(n21091), .A(n28479), .ZN(n21094) );
  NAND2_X1 U23531 ( .A1(n29134), .A2(n18919), .ZN(n21093) );
  AOI22_X1 U23532 ( .A1(n21096), .A2(n28479), .B1(n21094), .B2(n21093), .ZN(
        n21098) );
  NAND2_X1 U23533 ( .A1(n21098), .A2(n21097), .ZN(n21099) );
  XNOR2_X1 U23534 ( .A(n22298), .B(n22768), .ZN(n21946) );
  NAND3_X1 U23536 ( .A1(n22141), .A2(n22145), .A3(n6532), .ZN(n21108) );
  NAND2_X1 U23537 ( .A1(n21106), .A2(n22141), .ZN(n21107) );
  INV_X1 U23538 ( .A(n22116), .ZN(n21871) );
  XNOR2_X1 U23539 ( .A(n21871), .B(n22052), .ZN(n21116) );
  NAND3_X1 U23540 ( .A1(n21156), .A2(n21155), .A3(n21159), .ZN(n21110) );
  OAI21_X1 U23541 ( .B1(n21111), .B2(n4960), .A(n21110), .ZN(n21112) );
  NAND2_X1 U23542 ( .A1(n21113), .A2(n21464), .ZN(n21564) );
  XNOR2_X1 U23544 ( .A(n28486), .B(n22410), .ZN(n22159) );
  XNOR2_X1 U23545 ( .A(n22159), .B(n21116), .ZN(n21133) );
  AOI21_X1 U23546 ( .B1(n21143), .B2(n21140), .A(n21119), .ZN(n21123) );
  AOI22_X1 U23547 ( .A1(n21119), .A2(n21118), .B1(n21144), .B2(n21140), .ZN(
        n21121) );
  OAI22_X1 U23548 ( .A1(n21123), .A2(n21122), .B1(n21121), .B2(n21120), .ZN(
        n22760) );
  INV_X1 U23549 ( .A(n22760), .ZN(n22328) );
  XNOR2_X1 U23550 ( .A(n22328), .B(n3374), .ZN(n21131) );
  NAND3_X1 U23551 ( .A1(n1832), .A2(n21496), .A3(n21495), .ZN(n21128) );
  XNOR2_X1 U23553 ( .A(n22409), .B(n22414), .ZN(n21130) );
  XNOR2_X1 U23554 ( .A(n21131), .B(n21130), .ZN(n21132) );
  XNOR2_X1 U23555 ( .A(n21133), .B(n21132), .ZN(n23678) );
  NOR2_X1 U23556 ( .A1(n23360), .A2(n23678), .ZN(n23367) );
  XNOR2_X1 U23557 ( .A(n22418), .B(n22822), .ZN(n21149) );
  NOR2_X1 U23558 ( .A1(n21140), .A2(n21143), .ZN(n21142) );
  NOR2_X1 U23559 ( .A1(n21142), .A2(n21141), .ZN(n21147) );
  XNOR2_X1 U23560 ( .A(n22059), .B(n26680), .ZN(n21148) );
  XNOR2_X1 U23561 ( .A(n21149), .B(n21148), .ZN(n21170) );
  NAND2_X1 U23562 ( .A1(n21311), .A2(n21309), .ZN(n21152) );
  INV_X1 U23564 ( .A(n22419), .ZN(n21154) );
  XNOR2_X1 U23565 ( .A(n22098), .B(n21154), .ZN(n21168) );
  NAND3_X1 U23566 ( .A1(n21156), .A2(n4960), .A3(n21155), .ZN(n21161) );
  INV_X1 U23567 ( .A(n21618), .ZN(n21166) );
  AND2_X1 U23568 ( .A1(n21162), .A2(n21613), .ZN(n21165) );
  INV_X1 U23569 ( .A(n21326), .ZN(n21608) );
  XNOR2_X1 U23570 ( .A(n22656), .B(n22506), .ZN(n22801) );
  INV_X1 U23571 ( .A(n22801), .ZN(n21167) );
  XNOR2_X1 U23572 ( .A(n21167), .B(n21168), .ZN(n21169) );
  NAND3_X1 U23573 ( .A1(n21412), .A2(n21414), .A3(n28184), .ZN(n21175) );
  AND2_X1 U23574 ( .A1(n21410), .A2(n21171), .ZN(n21173) );
  INV_X1 U23575 ( .A(n21410), .ZN(n21172) );
  AOI22_X1 U23576 ( .A1(n21414), .A2(n21173), .B1(n21172), .B2(n21408), .ZN(
        n21174) );
  NAND2_X1 U23578 ( .A1(n21549), .A2(n1875), .ZN(n21179) );
  NAND3_X1 U23579 ( .A1(n21180), .A2(n21549), .A3(n21547), .ZN(n21178) );
  XNOR2_X1 U23580 ( .A(n21182), .B(n22678), .ZN(n22752) );
  INV_X1 U23581 ( .A(n22752), .ZN(n21191) );
  NOR2_X1 U23582 ( .A1(n1832), .A2(n28789), .ZN(n21184) );
  NAND2_X1 U23584 ( .A1(n22286), .A2(n21213), .ZN(n21189) );
  XNOR2_X1 U23585 ( .A(n22427), .B(n22068), .ZN(n21190) );
  XNOR2_X1 U23586 ( .A(n21191), .B(n21190), .ZN(n21206) );
  NAND2_X1 U23588 ( .A1(n21503), .A2(n21500), .ZN(n21196) );
  NOR2_X1 U23589 ( .A1(n21503), .A2(n28619), .ZN(n21194) );
  XNOR2_X1 U23591 ( .A(n29489), .B(n22855), .ZN(n21204) );
  AOI22_X1 U23592 ( .A1(n21198), .A2(n21532), .B1(n21514), .B2(n21512), .ZN(
        n21202) );
  NOR2_X1 U23593 ( .A1(n21514), .A2(n21530), .ZN(n21200) );
  AOI22_X1 U23594 ( .A1(n21200), .A2(n21509), .B1(n21533), .B2(n21199), .ZN(
        n21201) );
  XNOR2_X1 U23595 ( .A(n22854), .B(n900), .ZN(n21203) );
  XNOR2_X1 U23596 ( .A(n21204), .B(n21203), .ZN(n21205) );
  NOR2_X1 U23597 ( .A1(n23672), .A2(n23131), .ZN(n21207) );
  NOR2_X1 U23598 ( .A1(n23367), .A2(n21207), .ZN(n23108) );
  INV_X1 U23599 ( .A(n23678), .ZN(n23363) );
  OAI21_X1 U23600 ( .B1(n28790), .B2(n22286), .A(n21208), .ZN(n21214) );
  AOI21_X1 U23601 ( .B1(n21210), .B2(n21209), .A(n22290), .ZN(n21212) );
  AND2_X1 U23602 ( .A1(n21215), .A2(n21221), .ZN(n21225) );
  OR2_X1 U23603 ( .A1(n21220), .A2(n21216), .ZN(n21224) );
  NAND2_X1 U23604 ( .A1(n21220), .A2(n381), .ZN(n21222) );
  NAND2_X1 U23605 ( .A1(n21218), .A2(n21217), .ZN(n21219) );
  OAI22_X1 U23606 ( .A1(n21222), .A2(n21221), .B1(n21220), .B2(n21219), .ZN(
        n21223) );
  XNOR2_X1 U23607 ( .A(n29079), .B(n28517), .ZN(n21671) );
  XNOR2_X1 U23608 ( .A(n22164), .B(n21671), .ZN(n21241) );
  XNOR2_X1 U23609 ( .A(n22194), .B(n2465), .ZN(n21239) );
  INV_X1 U23610 ( .A(n21472), .ZN(n21478) );
  MUX2_X1 U23611 ( .A(n1930), .B(n21471), .S(n21478), .Z(n21234) );
  NOR2_X1 U23612 ( .A1(n21389), .A2(n21473), .ZN(n21231) );
  NAND2_X1 U23613 ( .A1(n21231), .A2(n1930), .ZN(n21232) );
  NAND2_X1 U23615 ( .A1(n21748), .A2(n20658), .ZN(n21235) );
  NAND2_X1 U23616 ( .A1(n21645), .A2(n21400), .ZN(n21646) );
  OAI22_X1 U23617 ( .A1(n21235), .A2(n21749), .B1(n20658), .B2(n21646), .ZN(
        n21238) );
  NAND2_X1 U23618 ( .A1(n21402), .A2(n497), .ZN(n21236) );
  XNOR2_X1 U23619 ( .A(n22195), .B(n22278), .ZN(n22442) );
  XNOR2_X1 U23620 ( .A(n22442), .B(n21239), .ZN(n21240) );
  XNOR2_X1 U23621 ( .A(n21241), .B(n21240), .ZN(n23673) );
  NOR2_X1 U23622 ( .A1(n21346), .A2(n29101), .ZN(n21244) );
  NOR2_X1 U23623 ( .A1(n21242), .A2(n21698), .ZN(n21243) );
  NOR2_X1 U23624 ( .A1(n21348), .A2(n28440), .ZN(n21245) );
  NAND3_X1 U23626 ( .A1(n21251), .A2(n21250), .A3(n21249), .ZN(n21252) );
  OAI211_X1 U23627 ( .C1(n21254), .C2(n21253), .A(n19732), .B(n21252), .ZN(
        n21256) );
  OAI211_X1 U23628 ( .C1(n21808), .C2(n19732), .A(n21256), .B(n21255), .ZN(
        n21955) );
  XNOR2_X1 U23629 ( .A(n22204), .B(n21955), .ZN(n22436) );
  INV_X1 U23630 ( .A(n21713), .ZN(n21257) );
  NOR3_X1 U23631 ( .A1(n21714), .A2(n21366), .A3(n21258), .ZN(n21259) );
  AOI21_X1 U23632 ( .B1(n21261), .B2(n21260), .A(n21259), .ZN(n21262) );
  XNOR2_X1 U23633 ( .A(n22093), .B(n22561), .ZN(n22810) );
  XNOR2_X1 U23635 ( .A(n28432), .B(n22436), .ZN(n21300) );
  INV_X1 U23636 ( .A(n21269), .ZN(n21270) );
  XNOR2_X1 U23637 ( .A(n22363), .B(n3516), .ZN(n21298) );
  NAND2_X1 U23639 ( .A1(n21274), .A2(n29227), .ZN(n21285) );
  INV_X1 U23640 ( .A(n21275), .ZN(n21276) );
  NAND2_X1 U23641 ( .A1(n29526), .A2(n21276), .ZN(n21282) );
  NAND2_X1 U23642 ( .A1(n21372), .A2(n496), .ZN(n21279) );
  NAND2_X1 U23643 ( .A1(n21279), .A2(n21278), .ZN(n21280) );
  OAI211_X1 U23644 ( .C1(n21283), .C2(n21282), .A(n21281), .B(n21280), .ZN(
        n21284) );
  NAND2_X1 U23645 ( .A1(n21288), .A2(n21287), .ZN(n21294) );
  NAND2_X1 U23646 ( .A1(n21294), .A2(n29313), .ZN(n21296) );
  NAND2_X1 U23647 ( .A1(n21291), .A2(n21290), .ZN(n21293) );
  MUX2_X1 U23648 ( .A(n21294), .B(n21293), .S(n21292), .Z(n21295) );
  XNOR2_X1 U23649 ( .A(n22501), .B(n22644), .ZN(n22776) );
  XNOR2_X1 U23650 ( .A(n22776), .B(n21298), .ZN(n21299) );
  OAI211_X1 U23652 ( .C1(n23363), .C2(n23673), .A(n23672), .B(n28604), .ZN(
        n21301) );
  OAI21_X1 U23653 ( .B1(n21302), .B2(n23108), .A(n21301), .ZN(n24748) );
  INV_X1 U23654 ( .A(n24748), .ZN(n21303) );
  INV_X1 U23655 ( .A(n22594), .ZN(n22077) );
  OAI21_X1 U23656 ( .B1(n29328), .B2(n21307), .A(n21311), .ZN(n21313) );
  NOR2_X1 U23657 ( .A1(n21308), .A2(n29531), .ZN(n21312) );
  NAND3_X1 U23658 ( .A1(n21316), .A2(n21315), .A3(n21314), .ZN(n21318) );
  NAND3_X1 U23659 ( .A1(n21603), .A2(n21601), .A3(n21600), .ZN(n21317) );
  AOI21_X1 U23660 ( .B1(n21613), .B2(n21327), .A(n21326), .ZN(n21337) );
  NAND2_X1 U23661 ( .A1(n21328), .A2(n21327), .ZN(n21333) );
  NAND3_X1 U23662 ( .A1(n21331), .A2(n20497), .A3(n21330), .ZN(n21332) );
  XNOR2_X1 U23663 ( .A(n29514), .B(n3276), .ZN(n21338) );
  XNOR2_X1 U23664 ( .A(n21339), .B(n21338), .ZN(n21340) );
  XNOR2_X1 U23665 ( .A(n22664), .B(n3049), .ZN(n21342) );
  XNOR2_X1 U23666 ( .A(n21342), .B(n28517), .ZN(n21371) );
  NAND2_X1 U23667 ( .A1(n21692), .A2(n28440), .ZN(n21345) );
  OAI21_X1 U23668 ( .B1(n21346), .B2(n21345), .A(n21344), .ZN(n21352) );
  NOR2_X1 U23670 ( .A1(n21348), .A2(n21698), .ZN(n21349) );
  NOR2_X2 U23672 ( .A1(n21352), .A2(n21351), .ZN(n22380) );
  MUX2_X1 U23673 ( .A(n21713), .B(n21714), .S(n21366), .Z(n21369) );
  NAND2_X1 U23674 ( .A1(n28491), .A2(n21354), .ZN(n21358) );
  NAND2_X1 U23675 ( .A1(n28126), .A2(n21354), .ZN(n21357) );
  MUX2_X1 U23676 ( .A(n21358), .B(n21357), .S(n28133), .Z(n21363) );
  NAND2_X1 U23677 ( .A1(n21360), .A2(n28586), .ZN(n21361) );
  NAND3_X1 U23678 ( .A1(n21363), .A2(n21362), .A3(n21361), .ZN(n21365) );
  AND2_X1 U23679 ( .A1(n21364), .A2(n21365), .ZN(n21368) );
  XNOR2_X1 U23680 ( .A(n22380), .B(n22628), .ZN(n21370) );
  XNOR2_X1 U23681 ( .A(n21371), .B(n21370), .ZN(n21386) );
  MUX2_X1 U23682 ( .A(n21373), .B(n21372), .S(n21704), .Z(n21376) );
  INV_X1 U23685 ( .A(n22625), .ZN(n21383) );
  XNOR2_X1 U23686 ( .A(n21384), .B(n21383), .ZN(n21385) );
  INV_X1 U23687 ( .A(n21389), .ZN(n21476) );
  NAND2_X1 U23688 ( .A1(n1930), .A2(n21476), .ZN(n21390) );
  XNOR2_X1 U23689 ( .A(n22326), .B(n22052), .ZN(n21407) );
  NOR3_X1 U23690 ( .A1(n21394), .A2(n21638), .A3(n21639), .ZN(n21397) );
  NOR2_X1 U23691 ( .A1(n21639), .A2(n21395), .ZN(n21396) );
  NOR2_X1 U23692 ( .A1(n21397), .A2(n21396), .ZN(n21398) );
  NAND3_X1 U23693 ( .A1(n21401), .A2(n21400), .A3(n21399), .ZN(n21405) );
  OAI21_X1 U23694 ( .B1(n21749), .B2(n20658), .A(n21748), .ZN(n21404) );
  NOR3_X1 U23695 ( .A1(n21749), .A2(n21402), .A3(n497), .ZN(n21403) );
  XNOR2_X1 U23696 ( .A(n22158), .B(n22411), .ZN(n22325) );
  INV_X1 U23697 ( .A(n22325), .ZN(n21406) );
  XNOR2_X1 U23698 ( .A(n21407), .B(n21406), .ZN(n21419) );
  OAI21_X1 U23699 ( .B1(n21410), .B2(n21409), .A(n21408), .ZN(n21411) );
  XNOR2_X1 U23700 ( .A(n22912), .B(n22473), .ZN(n21417) );
  XNOR2_X1 U23701 ( .A(n22844), .B(n1179), .ZN(n21416) );
  XNOR2_X1 U23702 ( .A(n21417), .B(n21416), .ZN(n21418) );
  OAI21_X1 U23704 ( .B1(n23344), .B2(n23338), .A(n28570), .ZN(n21529) );
  NAND2_X1 U23705 ( .A1(n21421), .A2(n21425), .ZN(n21423) );
  NAND2_X1 U23706 ( .A1(n21423), .A2(n21422), .ZN(n21427) );
  XNOR2_X1 U23707 ( .A(n22897), .B(n22434), .ZN(n21446) );
  MUX2_X1 U23708 ( .A(n21664), .B(n22398), .S(n21429), .Z(n21430) );
  NOR2_X1 U23709 ( .A1(n21430), .A2(n22404), .ZN(n21434) );
  NOR2_X1 U23710 ( .A1(n21014), .A2(n21433), .ZN(n22396) );
  NAND2_X1 U23711 ( .A1(n21653), .A2(n21657), .ZN(n21445) );
  INV_X1 U23712 ( .A(n21435), .ZN(n21436) );
  NOR2_X1 U23713 ( .A1(n21437), .A2(n21436), .ZN(n21438) );
  NAND2_X1 U23714 ( .A1(n21443), .A2(n21656), .ZN(n21444) );
  XNOR2_X1 U23715 ( .A(n22333), .B(n22479), .ZN(n21876) );
  XNOR2_X1 U23716 ( .A(n21446), .B(n21876), .ZN(n21456) );
  INV_X1 U23717 ( .A(n21447), .ZN(n21452) );
  OAI21_X1 U23718 ( .B1(n21677), .B2(n21674), .A(n21680), .ZN(n21451) );
  NOR2_X1 U23719 ( .A1(n21673), .A2(n21674), .ZN(n21450) );
  INV_X1 U23720 ( .A(n891), .ZN(n27788) );
  XNOR2_X1 U23721 ( .A(n22334), .B(n27788), .ZN(n21453) );
  XNOR2_X1 U23722 ( .A(n21454), .B(n21453), .ZN(n21455) );
  XNOR2_X1 U23725 ( .A(n22605), .B(n22677), .ZN(n21970) );
  XNOR2_X1 U23726 ( .A(n21470), .B(n21970), .ZN(n21492) );
  NAND2_X1 U23727 ( .A1(n21473), .A2(n21472), .ZN(n21474) );
  NAND2_X1 U23728 ( .A1(n21475), .A2(n21474), .ZN(n21480) );
  NAND2_X1 U23729 ( .A1(n21477), .A2(n21476), .ZN(n21479) );
  XNOR2_X1 U23730 ( .A(n22610), .B(n22068), .ZN(n21490) );
  XNOR2_X1 U23734 ( .A(n21889), .B(n2912), .ZN(n21489) );
  XNOR2_X1 U23735 ( .A(n21490), .B(n21489), .ZN(n21491) );
  AOI21_X1 U23737 ( .B1(n21501), .B2(n21500), .A(n21499), .ZN(n21508) );
  NOR2_X1 U23739 ( .A1(n21503), .A2(n28185), .ZN(n21506) );
  INV_X1 U23740 ( .A(n21504), .ZN(n21505) );
  XNOR2_X1 U23742 ( .A(n22374), .B(n22619), .ZN(n21523) );
  NAND3_X1 U23743 ( .A1(n21509), .A2(n21513), .A3(n21514), .ZN(n21510) );
  NAND2_X1 U23744 ( .A1(n21511), .A2(n21510), .ZN(n21518) );
  NAND2_X1 U23745 ( .A1(n21520), .A2(n21551), .ZN(n21521) );
  INV_X1 U23746 ( .A(n22567), .ZN(n22487) );
  XNOR2_X1 U23747 ( .A(n22487), .B(n22615), .ZN(n21881) );
  XNOR2_X1 U23748 ( .A(n21881), .B(n21523), .ZN(n21527) );
  XNOR2_X1 U23749 ( .A(n22059), .B(n5490), .ZN(n21524) );
  XNOR2_X1 U23750 ( .A(n21525), .B(n21524), .ZN(n21526) );
  XNOR2_X1 U23751 ( .A(n21527), .B(n21526), .ZN(n23138) );
  OAI21_X1 U23752 ( .B1(n29108), .B2(n28659), .A(n23139), .ZN(n21528) );
  XNOR2_X1 U23753 ( .A(n22522), .B(n21537), .ZN(n21546) );
  NAND2_X1 U23754 ( .A1(n21540), .A2(n21539), .ZN(n21542) );
  XNOR2_X1 U23755 ( .A(n22594), .B(n21980), .ZN(n21545) );
  OAI21_X1 U23757 ( .B1(n21551), .B2(n21550), .A(n21549), .ZN(n21555) );
  INV_X1 U23758 ( .A(n21552), .ZN(n21554) );
  XNOR2_X1 U23759 ( .A(n22768), .B(n22829), .ZN(n22313) );
  XNOR2_X1 U23760 ( .A(n21982), .B(n22033), .ZN(n21557) );
  XNOR2_X1 U23761 ( .A(n22313), .B(n21557), .ZN(n21558) );
  XNOR2_X2 U23762 ( .A(n21558), .B(n21559), .ZN(n23662) );
  AND2_X1 U23763 ( .A1(n21561), .A2(n21560), .ZN(n21562) );
  XNOR2_X1 U23764 ( .A(n22887), .B(n27894), .ZN(n21566) );
  INV_X1 U23765 ( .A(n21568), .ZN(n21569) );
  XNOR2_X1 U23766 ( .A(n22656), .B(n22891), .ZN(n21573) );
  NOR2_X1 U23767 ( .A1(n21575), .A2(n21574), .ZN(n21578) );
  XNOR2_X1 U23768 ( .A(n21987), .B(n22059), .ZN(n21582) );
  XNOR2_X1 U23769 ( .A(n21582), .B(n22619), .ZN(n21583) );
  INV_X1 U23770 ( .A(n22644), .ZN(n21593) );
  XNOR2_X1 U23771 ( .A(n21998), .B(n21593), .ZN(n21595) );
  XNOR2_X1 U23772 ( .A(n22692), .B(n2544), .ZN(n21594) );
  XNOR2_X1 U23773 ( .A(n21595), .B(n21594), .ZN(n21622) );
  NOR2_X1 U23774 ( .A1(n21601), .A2(n21600), .ZN(n21602) );
  NAND2_X1 U23775 ( .A1(n21603), .A2(n21602), .ZN(n21604) );
  NAND3_X1 U23776 ( .A1(n21608), .A2(n21607), .A3(n21613), .ZN(n21617) );
  INV_X1 U23777 ( .A(n21611), .ZN(n21615) );
  NAND2_X1 U23778 ( .A1(n21613), .A2(n21612), .ZN(n21614) );
  XNOR2_X1 U23779 ( .A(n22500), .B(n22813), .ZN(n22899) );
  XNOR2_X1 U23780 ( .A(n22899), .B(n21620), .ZN(n21621) );
  XNOR2_X1 U23781 ( .A(n21621), .B(n21622), .ZN(n23162) );
  AOI21_X1 U23782 ( .B1(n22146), .B2(n22145), .A(n21623), .ZN(n21628) );
  INV_X1 U23783 ( .A(n22717), .ZN(n21800) );
  XNOR2_X1 U23784 ( .A(n21800), .B(n22606), .ZN(n21630) );
  XNOR2_X1 U23785 ( .A(n22068), .B(n2389), .ZN(n21629) );
  XNOR2_X1 U23786 ( .A(n21630), .B(n21629), .ZN(n21652) );
  NOR2_X1 U23787 ( .A1(n21633), .A2(n21632), .ZN(n21636) );
  AOI21_X1 U23788 ( .B1(n21639), .B2(n21636), .A(n21635), .ZN(n21641) );
  OR3_X1 U23789 ( .A1(n21639), .A2(n21638), .A3(n21637), .ZN(n21640) );
  XNOR2_X1 U23790 ( .A(n22180), .B(n22678), .ZN(n22341) );
  NAND2_X1 U23791 ( .A1(n21042), .A2(n21642), .ZN(n21644) );
  NAND2_X1 U23792 ( .A1(n21750), .A2(n21645), .ZN(n21647) );
  XNOR2_X1 U23793 ( .A(n22067), .B(n21649), .ZN(n22181) );
  INV_X1 U23794 ( .A(n22181), .ZN(n21650) );
  XNOR2_X1 U23795 ( .A(n22341), .B(n21650), .ZN(n21651) );
  XNOR2_X1 U23796 ( .A(n21651), .B(n21652), .ZN(n23006) );
  INV_X1 U23797 ( .A(n23006), .ZN(n23665) );
  OAI21_X1 U23798 ( .B1(n23666), .B2(n23162), .A(n23665), .ZN(n21690) );
  NOR2_X1 U23799 ( .A1(n23666), .A2(n23006), .ZN(n23164) );
  NOR2_X1 U23800 ( .A1(n21654), .A2(n21653), .ZN(n21659) );
  NOR2_X1 U23801 ( .A1(n21656), .A2(n21655), .ZN(n21658) );
  NOR2_X1 U23802 ( .A1(n21662), .A2(n22401), .ZN(n21668) );
  NOR2_X1 U23803 ( .A1(n21664), .A2(n21663), .ZN(n21669) );
  NOR2_X1 U23804 ( .A1(n21665), .A2(n22397), .ZN(n21666) );
  NOR2_X1 U23805 ( .A1(n21669), .A2(n21666), .ZN(n21667) );
  XNOR2_X1 U23807 ( .A(n22574), .B(n22542), .ZN(n22193) );
  XNOR2_X1 U23808 ( .A(n21671), .B(n22193), .ZN(n21689) );
  XNOR2_X1 U23809 ( .A(n22710), .B(n22625), .ZN(n21687) );
  INV_X1 U23810 ( .A(n21672), .ZN(n21685) );
  OAI21_X1 U23811 ( .B1(n21675), .B2(n21674), .A(n21673), .ZN(n21684) );
  NAND2_X1 U23812 ( .A1(n21677), .A2(n21676), .ZN(n21682) );
  NAND2_X1 U23813 ( .A1(n21679), .A2(n21678), .ZN(n21681) );
  MUX2_X1 U23814 ( .A(n21682), .B(n21681), .S(n21680), .Z(n21683) );
  XNOR2_X1 U23815 ( .A(n22221), .B(n3787), .ZN(n21686) );
  XNOR2_X1 U23816 ( .A(n21687), .B(n21686), .ZN(n21688) );
  XNOR2_X1 U23817 ( .A(n21689), .B(n21688), .ZN(n23163) );
  AOI22_X1 U23818 ( .A1(n23662), .A2(n21690), .B1(n23164), .B2(n23163), .ZN(
        n21725) );
  INV_X1 U23819 ( .A(n21691), .ZN(n21693) );
  INV_X1 U23820 ( .A(n21692), .ZN(n21694) );
  NOR2_X1 U23821 ( .A1(n21693), .A2(n21694), .ZN(n21701) );
  NOR2_X1 U23822 ( .A1(n21695), .A2(n21694), .ZN(n21700) );
  AOI21_X1 U23823 ( .B1(n21698), .B2(n21697), .A(n3260), .ZN(n21699) );
  XNOR2_X1 U23824 ( .A(n21872), .B(n22734), .ZN(n21719) );
  NAND3_X1 U23825 ( .A1(n21705), .A2(n21704), .A3(n21703), .ZN(n21706) );
  NOR2_X1 U23826 ( .A1(n21709), .A2(n21708), .ZN(n21710) );
  NOR2_X2 U23827 ( .A1(n21711), .A2(n21710), .ZN(n22589) );
  AOI21_X1 U23828 ( .B1(n21714), .B2(n21713), .A(n21712), .ZN(n21715) );
  OAI22_X1 U23829 ( .A1(n21718), .A2(n21717), .B1(n21716), .B2(n21715), .ZN(
        n22535) );
  XNOR2_X1 U23830 ( .A(n22589), .B(n22535), .ZN(n22908) );
  XNOR2_X1 U23831 ( .A(n22908), .B(n21719), .ZN(n21723) );
  XNOR2_X1 U23832 ( .A(n22052), .B(n22411), .ZN(n21721) );
  INV_X1 U23833 ( .A(n3212), .ZN(n27936) );
  XNOR2_X1 U23834 ( .A(n22328), .B(n27936), .ZN(n21720) );
  XNOR2_X1 U23835 ( .A(n21720), .B(n21721), .ZN(n21722) );
  XNOR2_X1 U23836 ( .A(n21723), .B(n21722), .ZN(n23525) );
  NAND2_X1 U23837 ( .A1(n29123), .A2(n23163), .ZN(n21898) );
  MUX2_X1 U23839 ( .A(n493), .B(n29314), .S(n1930), .Z(n21737) );
  INV_X1 U23840 ( .A(n21731), .ZN(n21732) );
  NAND2_X1 U23841 ( .A1(n21732), .A2(n21736), .ZN(n21735) );
  NAND2_X1 U23842 ( .A1(n21733), .A2(n493), .ZN(n21734) );
  OAI211_X1 U23843 ( .C1(n21737), .C2(n21736), .A(n21735), .B(n21734), .ZN(
        n21738) );
  XNOR2_X1 U23844 ( .A(n22643), .B(n3323), .ZN(n21740) );
  XNOR2_X1 U23845 ( .A(n21739), .B(n21740), .ZN(n21741) );
  XNOR2_X1 U23846 ( .A(n21741), .B(n21742), .ZN(n23783) );
  INV_X1 U23847 ( .A(n23783), .ZN(n23785) );
  INV_X1 U23848 ( .A(n22426), .ZN(n21743) );
  XNOR2_X1 U23849 ( .A(n21743), .B(n21801), .ZN(n22749) );
  XNOR2_X1 U23850 ( .A(n22609), .B(n22553), .ZN(n22037) );
  XNOR2_X1 U23851 ( .A(n22749), .B(n22037), .ZN(n21747) );
  XNOR2_X1 U23852 ( .A(n22681), .B(n29490), .ZN(n21745) );
  INV_X1 U23853 ( .A(n22006), .ZN(n22515) );
  INV_X1 U23854 ( .A(n2441), .ZN(n26314) );
  XNOR2_X1 U23855 ( .A(n22515), .B(n26314), .ZN(n21744) );
  XNOR2_X1 U23856 ( .A(n21745), .B(n21744), .ZN(n21746) );
  INV_X1 U23858 ( .A(n21825), .ZN(n22285) );
  XNOR2_X1 U23859 ( .A(n22285), .B(n22526), .ZN(n21755) );
  MUX2_X1 U23860 ( .A(n21749), .B(n21042), .S(n21748), .Z(n21752) );
  MUX2_X1 U23861 ( .A(n21752), .B(n21751), .S(n21750), .Z(n22584) );
  XNOR2_X1 U23862 ( .A(n22199), .B(n2476), .ZN(n21753) );
  XNOR2_X1 U23863 ( .A(n21753), .B(n22584), .ZN(n21754) );
  XNOR2_X1 U23864 ( .A(n21755), .B(n21754), .ZN(n21757) );
  INV_X1 U23865 ( .A(n21758), .ZN(n22786) );
  INV_X1 U23866 ( .A(n22195), .ZN(n21759) );
  XNOR2_X1 U23867 ( .A(n22786), .B(n21759), .ZN(n21761) );
  XNOR2_X1 U23868 ( .A(n22218), .B(n22790), .ZN(n22015) );
  XNOR2_X1 U23869 ( .A(n28449), .B(n72), .ZN(n21762) );
  XNOR2_X1 U23870 ( .A(n22015), .B(n21762), .ZN(n21763) );
  XNOR2_X1 U23871 ( .A(n21764), .B(n21763), .ZN(n23784) );
  XNOR2_X1 U23872 ( .A(n22409), .B(n3087), .ZN(n21765) );
  XNOR2_X1 U23873 ( .A(n22601), .B(n28589), .ZN(n21767) );
  XNOR2_X1 U23874 ( .A(n22472), .B(n21767), .ZN(n22048) );
  XNOR2_X1 U23875 ( .A(n21768), .B(n22048), .ZN(n21775) );
  INV_X1 U23876 ( .A(n22798), .ZN(n22422) );
  XNOR2_X1 U23877 ( .A(n22422), .B(n22418), .ZN(n21770) );
  XNOR2_X1 U23878 ( .A(n22796), .B(n21959), .ZN(n22569) );
  XNOR2_X1 U23879 ( .A(n21770), .B(n22569), .ZN(n21774) );
  XNOR2_X1 U23880 ( .A(n28492), .B(n1123), .ZN(n21772) );
  XNOR2_X1 U23882 ( .A(n22509), .B(n22724), .ZN(n21771) );
  XNOR2_X1 U23883 ( .A(n21772), .B(n21771), .ZN(n21773) );
  XNOR2_X1 U23884 ( .A(n21774), .B(n21773), .ZN(n23786) );
  INV_X1 U23885 ( .A(n23786), .ZN(n23005) );
  INV_X1 U23886 ( .A(n21775), .ZN(n23482) );
  AOI211_X1 U23887 ( .C1(n23005), .C2(n23482), .A(n23484), .B(n23036), .ZN(
        n21776) );
  XNOR2_X1 U23888 ( .A(n22710), .B(n22086), .ZN(n21778) );
  XNOR2_X1 U23889 ( .A(n28517), .B(n22786), .ZN(n21777) );
  XNOR2_X1 U23890 ( .A(n21778), .B(n21777), .ZN(n21782) );
  INV_X1 U23891 ( .A(n22835), .ZN(n21995) );
  XNOR2_X1 U23892 ( .A(n21995), .B(n22219), .ZN(n21780) );
  XNOR2_X1 U23893 ( .A(n21780), .B(n21779), .ZN(n21781) );
  XNOR2_X1 U23894 ( .A(n22757), .B(n22052), .ZN(n21784) );
  XNOR2_X1 U23895 ( .A(n28461), .B(n22734), .ZN(n21783) );
  XNOR2_X1 U23896 ( .A(n21784), .B(n21783), .ZN(n21788) );
  XNOR2_X1 U23897 ( .A(n22763), .B(n3650), .ZN(n21785) );
  XNOR2_X1 U23898 ( .A(n21786), .B(n21785), .ZN(n21787) );
  XNOR2_X2 U23899 ( .A(n21788), .B(n21787), .ZN(n23765) );
  AND2_X1 U23900 ( .A1(n23767), .A2(n23765), .ZN(n21829) );
  XNOR2_X1 U23901 ( .A(n21789), .B(n22245), .ZN(n21792) );
  INV_X1 U23902 ( .A(n22363), .ZN(n21790) );
  XNOR2_X1 U23903 ( .A(n21956), .B(n21790), .ZN(n21791) );
  XNOR2_X1 U23904 ( .A(n22812), .B(n22692), .ZN(n21794) );
  XNOR2_X1 U23905 ( .A(n22778), .B(n2602), .ZN(n21793) );
  XNOR2_X1 U23906 ( .A(n21794), .B(n21793), .ZN(n21795) );
  XNOR2_X1 U23907 ( .A(n22821), .B(n22059), .ZN(n22617) );
  XNOR2_X1 U23908 ( .A(n22728), .B(n22617), .ZN(n21799) );
  XNOR2_X1 U23909 ( .A(n21959), .B(n1859), .ZN(n21797) );
  XNOR2_X1 U23910 ( .A(n22488), .B(n3770), .ZN(n21796) );
  XNOR2_X1 U23911 ( .A(n21797), .B(n21796), .ZN(n21798) );
  XNOR2_X1 U23912 ( .A(n22068), .B(n2404), .ZN(n21804) );
  XNOR2_X1 U23913 ( .A(n21800), .B(n21801), .ZN(n22259) );
  INV_X1 U23914 ( .A(n22718), .ZN(n21802) );
  XNOR2_X1 U23915 ( .A(n22259), .B(n21802), .ZN(n21803) );
  NAND3_X1 U23916 ( .A1(n21808), .A2(n21807), .A3(n21806), .ZN(n21815) );
  OAI21_X1 U23917 ( .B1(n21811), .B2(n21810), .A(n21809), .ZN(n21814) );
  INV_X1 U23918 ( .A(n21812), .ZN(n21813) );
  AOI21_X1 U23919 ( .B1(n21815), .B2(n21814), .A(n21813), .ZN(n22370) );
  XNOR2_X1 U23920 ( .A(n21816), .B(n22370), .ZN(n22008) );
  INV_X1 U23921 ( .A(n22703), .ZN(n21817) );
  INV_X1 U23923 ( .A(n21818), .ZN(n21822) );
  NOR2_X1 U23924 ( .A1(n491), .A2(n22013), .ZN(n21820) );
  AOI22_X1 U23925 ( .A1(n21823), .A2(n21820), .B1(n21819), .B2(n22013), .ZN(
        n21821) );
  OAI21_X1 U23926 ( .B1(n21823), .B2(n21822), .A(n21821), .ZN(n21824) );
  XNOR2_X1 U23927 ( .A(n21979), .B(n21824), .ZN(n22390) );
  INV_X1 U23928 ( .A(n22390), .ZN(n21828) );
  XNOR2_X1 U23929 ( .A(n22033), .B(n22226), .ZN(n22524) );
  XNOR2_X1 U23930 ( .A(n22524), .B(n21826), .ZN(n21827) );
  NOR2_X1 U23931 ( .A1(n23501), .A2(n23499), .ZN(n21830) );
  XNOR2_X1 U23932 ( .A(n22204), .B(n22265), .ZN(n22642) );
  XNOR2_X1 U23933 ( .A(n28387), .B(n22898), .ZN(n21831) );
  XNOR2_X1 U23934 ( .A(n22642), .B(n21831), .ZN(n21835) );
  XNOR2_X1 U23935 ( .A(n22330), .B(n22501), .ZN(n21833) );
  XNOR2_X1 U23936 ( .A(n22334), .B(n3386), .ZN(n21832) );
  XNOR2_X1 U23937 ( .A(n21833), .B(n21832), .ZN(n21834) );
  XNOR2_X1 U23939 ( .A(n22326), .B(n2353), .ZN(n21836) );
  XNOR2_X1 U23941 ( .A(n22302), .B(n22409), .ZN(n22650) );
  XNOR2_X1 U23942 ( .A(n21838), .B(n22650), .ZN(n21839) );
  XNOR2_X1 U23943 ( .A(n22374), .B(n21841), .ZN(n21842) );
  XNOR2_X1 U23944 ( .A(n22100), .B(n21842), .ZN(n21846) );
  XNOR2_X1 U23945 ( .A(n22822), .B(n22890), .ZN(n21844) );
  XNOR2_X1 U23946 ( .A(n22506), .B(n3211), .ZN(n21843) );
  XNOR2_X1 U23947 ( .A(n21844), .B(n21843), .ZN(n21845) );
  NOR2_X1 U23948 ( .A1(n339), .A2(n23772), .ZN(n21853) );
  XNOR2_X1 U23949 ( .A(n22386), .B(n3083), .ZN(n21849) );
  XNOR2_X1 U23950 ( .A(n22199), .B(n21850), .ZN(n22675) );
  INV_X1 U23951 ( .A(n22675), .ZN(n21851) );
  INV_X1 U23952 ( .A(n23156), .ZN(n23512) );
  AOI22_X1 U23953 ( .A1(n23488), .A2(n23513), .B1(n21853), .B2(n23512), .ZN(
        n21864) );
  XNOR2_X1 U23954 ( .A(n22240), .B(n29489), .ZN(n21854) );
  XNOR2_X1 U23955 ( .A(n21854), .B(n22340), .ZN(n22684) );
  XNOR2_X1 U23956 ( .A(n22514), .B(n22854), .ZN(n21855) );
  XNOR2_X1 U23957 ( .A(n22164), .B(n21856), .ZN(n21860) );
  XNOR2_X1 U23958 ( .A(n22380), .B(n27422), .ZN(n21858) );
  INV_X1 U23959 ( .A(n22279), .ZN(n21857) );
  XNOR2_X1 U23960 ( .A(n22195), .B(n21857), .ZN(n22663) );
  XNOR2_X1 U23961 ( .A(n22663), .B(n21858), .ZN(n21859) );
  XNOR2_X1 U23962 ( .A(n21859), .B(n21860), .ZN(n23771) );
  INV_X1 U23963 ( .A(n23771), .ZN(n23487) );
  NOR2_X1 U23964 ( .A1(n23487), .A2(n23772), .ZN(n21861) );
  XNOR2_X1 U23967 ( .A(n22194), .B(n22221), .ZN(n21912) );
  XNOR2_X1 U23968 ( .A(n22278), .B(n22380), .ZN(n22839) );
  XNOR2_X1 U23969 ( .A(n22839), .B(n21912), .ZN(n21868) );
  XNOR2_X1 U23970 ( .A(n22464), .B(n22784), .ZN(n22578) );
  XNOR2_X1 U23971 ( .A(n22628), .B(n21865), .ZN(n21866) );
  XNOR2_X1 U23972 ( .A(n22578), .B(n21866), .ZN(n21867) );
  XNOR2_X1 U23973 ( .A(n21868), .B(n21867), .ZN(n23802) );
  INV_X1 U23974 ( .A(n23802), .ZN(n23541) );
  XNOR2_X1 U23975 ( .A(n22158), .B(n3336), .ZN(n21870) );
  XNOR2_X1 U23976 ( .A(n22326), .B(n22414), .ZN(n22843) );
  XNOR2_X1 U23978 ( .A(n21870), .B(n28613), .ZN(n21874) );
  XNOR2_X1 U23979 ( .A(n21871), .B(n21872), .ZN(n21918) );
  XNOR2_X1 U23980 ( .A(n28162), .B(n22473), .ZN(n22588) );
  XNOR2_X1 U23981 ( .A(n22588), .B(n21918), .ZN(n21873) );
  XNOR2_X1 U23982 ( .A(n21998), .B(n21875), .ZN(n21940) );
  INV_X1 U23983 ( .A(n21940), .ZN(n21877) );
  XNOR2_X1 U23984 ( .A(n22690), .B(n29247), .ZN(n21878) );
  XNOR2_X1 U23985 ( .A(n21987), .B(n22098), .ZN(n21880) );
  XNOR2_X1 U23986 ( .A(n22723), .B(n2511), .ZN(n21879) );
  XNOR2_X1 U23987 ( .A(n21880), .B(n21879), .ZN(n21883) );
  XNOR2_X1 U23988 ( .A(n22374), .B(n22419), .ZN(n22819) );
  INV_X1 U23989 ( .A(n22819), .ZN(n22057) );
  XNOR2_X1 U23990 ( .A(n22057), .B(n21881), .ZN(n21882) );
  XNOR2_X1 U23991 ( .A(n22298), .B(n22386), .ZN(n22827) );
  XNOR2_X1 U23992 ( .A(n22827), .B(n21884), .ZN(n21887) );
  XNOR2_X1 U23993 ( .A(n21980), .B(n3554), .ZN(n21885) );
  XNOR2_X1 U23994 ( .A(n22152), .B(n29514), .ZN(n21947) );
  XNOR2_X1 U23995 ( .A(n21885), .B(n21947), .ZN(n21886) );
  XNOR2_X2 U23996 ( .A(n21887), .B(n21886), .ZN(n23689) );
  XNOR2_X1 U23997 ( .A(n22606), .B(n22855), .ZN(n21888) );
  XNOR2_X1 U23998 ( .A(n21970), .B(n21888), .ZN(n21892) );
  INV_X1 U23999 ( .A(n22852), .ZN(n22065) );
  XNOR2_X1 U24000 ( .A(n22750), .B(n3062), .ZN(n21890) );
  XNOR2_X1 U24001 ( .A(n22065), .B(n21890), .ZN(n21891) );
  INV_X1 U24002 ( .A(n23800), .ZN(n21893) );
  OAI22_X1 U24003 ( .A1(n21895), .A2(n23690), .B1(n23803), .B2(n21894), .ZN(
        n23932) );
  INV_X1 U24004 ( .A(n23932), .ZN(n24728) );
  OR2_X1 U24005 ( .A1(n24596), .A2(n24728), .ZN(n24732) );
  INV_X1 U24007 ( .A(n23666), .ZN(n21896) );
  NAND2_X1 U24008 ( .A1(n28577), .A2(n21896), .ZN(n21897) );
  MUX2_X1 U24009 ( .A(n21898), .B(n21897), .S(n23162), .Z(n21901) );
  NOR2_X1 U24010 ( .A1(n23163), .A2(n23663), .ZN(n21899) );
  NOR2_X1 U24011 ( .A1(n23162), .A2(n23006), .ZN(n23669) );
  AOI21_X1 U24012 ( .B1(n23662), .B2(n21899), .A(n23669), .ZN(n21900) );
  NAND2_X1 U24013 ( .A1(n21901), .A2(n21900), .ZN(n24595) );
  INV_X1 U24014 ( .A(n24595), .ZN(n24288) );
  NAND2_X1 U24015 ( .A1(n24732), .A2(n24724), .ZN(n21943) );
  XNOR2_X1 U24016 ( .A(n22820), .B(n22891), .ZN(n22061) );
  XNOR2_X1 U24017 ( .A(n22061), .B(n22098), .ZN(n22213) );
  XNOR2_X1 U24018 ( .A(n21902), .B(n22888), .ZN(n21904) );
  XNOR2_X1 U24019 ( .A(n21904), .B(n22620), .ZN(n21905) );
  XNOR2_X1 U24020 ( .A(n29591), .B(n22606), .ZN(n21907) );
  XNOR2_X1 U24021 ( .A(n22338), .B(n22067), .ZN(n22905) );
  INV_X1 U24022 ( .A(n22905), .ZN(n21906) );
  XNOR2_X1 U24023 ( .A(n21906), .B(n21907), .ZN(n21911) );
  XNOR2_X1 U24024 ( .A(n22718), .B(n22856), .ZN(n21909) );
  XNOR2_X1 U24025 ( .A(n22855), .B(n27105), .ZN(n21908) );
  XNOR2_X1 U24026 ( .A(n21909), .B(n21908), .ZN(n21910) );
  XNOR2_X1 U24027 ( .A(n22320), .B(n22542), .ZN(n22920) );
  XNOR2_X1 U24028 ( .A(n21912), .B(n22920), .ZN(n21916) );
  XNOR2_X1 U24029 ( .A(n22123), .B(n22219), .ZN(n21914) );
  XNOR2_X1 U24030 ( .A(n22664), .B(n1247), .ZN(n21913) );
  XNOR2_X1 U24031 ( .A(n21914), .B(n21913), .ZN(n21915) );
  XNOR2_X1 U24034 ( .A(n21917), .B(n22535), .ZN(n22187) );
  XNOR2_X1 U24035 ( .A(n21918), .B(n22187), .ZN(n21922) );
  XNOR2_X1 U24036 ( .A(n22731), .B(n28461), .ZN(n21920) );
  XNOR2_X1 U24037 ( .A(n28472), .B(n3035), .ZN(n21919) );
  XNOR2_X1 U24038 ( .A(n21920), .B(n21919), .ZN(n21921) );
  XNOR2_X1 U24039 ( .A(n21922), .B(n21921), .ZN(n23793) );
  XNOR2_X1 U24040 ( .A(n22697), .B(n22523), .ZN(n21924) );
  XNOR2_X1 U24041 ( .A(n22828), .B(n21924), .ZN(n21928) );
  XNOR2_X1 U24042 ( .A(n21980), .B(n22387), .ZN(n22595) );
  INV_X1 U24043 ( .A(n22595), .ZN(n21926) );
  XNOR2_X1 U24044 ( .A(n22522), .B(n3565), .ZN(n21925) );
  XNOR2_X1 U24045 ( .A(n21926), .B(n21925), .ZN(n21927) );
  NAND2_X1 U24046 ( .A1(n29586), .A2(n21932), .ZN(n21933) );
  OAI22_X1 U24047 ( .A1(n21934), .A2(n21933), .B1(n21932), .B2(n21931), .ZN(
        n21935) );
  INV_X1 U24048 ( .A(n22205), .ZN(n22080) );
  XNOR2_X1 U24049 ( .A(n22094), .B(n22245), .ZN(n21938) );
  XNOR2_X1 U24050 ( .A(n22080), .B(n21938), .ZN(n21942) );
  XNOR2_X1 U24051 ( .A(n22896), .B(n2598), .ZN(n21939) );
  XOR2_X1 U24052 ( .A(n21940), .B(n21939), .Z(n21941) );
  XNOR2_X1 U24055 ( .A(n22582), .B(n21946), .ZN(n21948) );
  XNOR2_X1 U24056 ( .A(n22158), .B(n22760), .ZN(n22117) );
  XNOR2_X1 U24057 ( .A(n21949), .B(n22301), .ZN(n22587) );
  XNOR2_X1 U24058 ( .A(n22117), .B(n22587), .ZN(n21953) );
  XNOR2_X1 U24059 ( .A(n22535), .B(n22473), .ZN(n21951) );
  XNOR2_X1 U24060 ( .A(n22414), .B(n1215), .ZN(n21950) );
  XNOR2_X1 U24061 ( .A(n21951), .B(n21950), .ZN(n21952) );
  NAND2_X1 U24063 ( .A1(n23606), .A2(n23247), .ZN(n23211) );
  XNOR2_X1 U24065 ( .A(n22479), .B(n22330), .ZN(n22641) );
  XNOR2_X1 U24066 ( .A(n22500), .B(n3463), .ZN(n21954) );
  XNOR2_X1 U24067 ( .A(n22641), .B(n21954), .ZN(n21958) );
  XNOR2_X1 U24068 ( .A(n21956), .B(n21955), .ZN(n22264) );
  XNOR2_X1 U24069 ( .A(n22333), .B(n22644), .ZN(n22092) );
  XNOR2_X1 U24070 ( .A(n22264), .B(n22092), .ZN(n21957) );
  XNOR2_X1 U24071 ( .A(n21957), .B(n21958), .ZN(n23245) );
  XNOR2_X1 U24072 ( .A(n22419), .B(n21959), .ZN(n22272) );
  XNOR2_X1 U24073 ( .A(n22272), .B(n22350), .ZN(n21963) );
  XNOR2_X1 U24074 ( .A(n22567), .B(n22891), .ZN(n21961) );
  XNOR2_X1 U24075 ( .A(n28483), .B(n3728), .ZN(n21960) );
  XNOR2_X1 U24076 ( .A(n21961), .B(n21960), .ZN(n21962) );
  XNOR2_X1 U24077 ( .A(n21963), .B(n21962), .ZN(n23246) );
  INV_X1 U24078 ( .A(n23246), .ZN(n23603) );
  XNOR2_X1 U24081 ( .A(n22278), .B(n22542), .ZN(n21967) );
  INV_X1 U24082 ( .A(n2477), .ZN(n26287) );
  XNOR2_X1 U24083 ( .A(n22464), .B(n26287), .ZN(n21966) );
  XNOR2_X1 U24084 ( .A(n21967), .B(n21966), .ZN(n21969) );
  XNOR2_X1 U24085 ( .A(n22783), .B(n22628), .ZN(n22318) );
  XNOR2_X1 U24086 ( .A(n22575), .B(n22318), .ZN(n21968) );
  INV_X1 U24087 ( .A(n23607), .ZN(n22985) );
  INV_X1 U24088 ( .A(n23247), .ZN(n23578) );
  XNOR2_X1 U24089 ( .A(n21970), .B(n21971), .ZN(n21975) );
  XNOR2_X1 U24090 ( .A(n22678), .B(n22067), .ZN(n21973) );
  XNOR2_X1 U24091 ( .A(n6504), .B(n1062), .ZN(n21972) );
  XNOR2_X1 U24092 ( .A(n21973), .B(n21972), .ZN(n21974) );
  XNOR2_X1 U24093 ( .A(n21974), .B(n21975), .ZN(n23602) );
  INV_X1 U24094 ( .A(n23602), .ZN(n23583) );
  OAI21_X1 U24095 ( .B1(n22985), .B2(n23578), .A(n23583), .ZN(n21976) );
  NAND2_X1 U24096 ( .A1(n21976), .A2(n23577), .ZN(n21977) );
  XNOR2_X1 U24099 ( .A(n22671), .B(n25044), .ZN(n21984) );
  XNOR2_X1 U24100 ( .A(n21982), .B(n22226), .ZN(n21983) );
  XNOR2_X1 U24101 ( .A(n21984), .B(n21983), .ZN(n21985) );
  XNOR2_X1 U24102 ( .A(n21987), .B(n22509), .ZN(n22252) );
  XNOR2_X1 U24103 ( .A(n22252), .B(n22821), .ZN(n22886) );
  XNOR2_X1 U24104 ( .A(n22488), .B(n1858), .ZN(n21988) );
  XNOR2_X1 U24105 ( .A(n22886), .B(n21989), .ZN(n23258) );
  XNOR2_X1 U24106 ( .A(n22411), .B(n22735), .ZN(n22188) );
  XNOR2_X1 U24107 ( .A(n22599), .B(n22188), .ZN(n21993) );
  INV_X1 U24108 ( .A(n22472), .ZN(n22300) );
  XNOR2_X1 U24109 ( .A(n22300), .B(n4029), .ZN(n21991) );
  XNOR2_X1 U24110 ( .A(n22533), .B(n21991), .ZN(n21992) );
  XNOR2_X1 U24111 ( .A(n22459), .B(n22625), .ZN(n22192) );
  XNOR2_X1 U24112 ( .A(n21994), .B(n22792), .ZN(n22220) );
  XNOR2_X1 U24113 ( .A(n22192), .B(n22220), .ZN(n21997) );
  XNOR2_X1 U24114 ( .A(n21995), .B(n22221), .ZN(n22922) );
  NAND2_X1 U24115 ( .A1(n23735), .A2(n23227), .ZN(n23734) );
  INV_X1 U24116 ( .A(n21998), .ZN(n21999) );
  XNOR2_X1 U24117 ( .A(n22000), .B(n21789), .ZN(n22001) );
  XNOR2_X1 U24118 ( .A(n29136), .B(n22001), .ZN(n22005) );
  XNOR2_X1 U24119 ( .A(n22643), .B(n22434), .ZN(n22003) );
  XNOR2_X1 U24120 ( .A(n22778), .B(n2916), .ZN(n22002) );
  XNOR2_X1 U24121 ( .A(n22003), .B(n22002), .ZN(n22004) );
  XNOR2_X1 U24122 ( .A(n22606), .B(n22006), .ZN(n22238) );
  XNOR2_X1 U24123 ( .A(n22681), .B(n26825), .ZN(n22007) );
  AOI21_X1 U24124 ( .B1(n22010), .B2(n23734), .A(n22009), .ZN(n23962) );
  AND2_X1 U24125 ( .A1(n24583), .A2(n23962), .ZN(n24586) );
  XNOR2_X1 U24126 ( .A(n22923), .B(n22015), .ZN(n22018) );
  XNOR2_X1 U24127 ( .A(n28450), .B(n24897), .ZN(n22016) );
  XNOR2_X1 U24128 ( .A(n22017), .B(n22018), .ZN(n22976) );
  INV_X1 U24129 ( .A(n22976), .ZN(n23408) );
  XNOR2_X1 U24130 ( .A(n22633), .B(n28387), .ZN(n22020) );
  XNOR2_X1 U24131 ( .A(n21728), .B(n3036), .ZN(n22019) );
  XNOR2_X1 U24132 ( .A(n22020), .B(n22019), .ZN(n22021) );
  OAI211_X1 U24136 ( .C1(n489), .C2(n21019), .A(n22291), .B(n22025), .ZN(
        n22030) );
  INV_X1 U24138 ( .A(n1927), .ZN(n28108) );
  OAI21_X1 U24139 ( .B1(n22027), .B2(n22028), .A(n28108), .ZN(n22029) );
  XNOR2_X1 U24140 ( .A(n22031), .B(n22032), .ZN(n22036) );
  XNOR2_X1 U24141 ( .A(n22830), .B(n22033), .ZN(n22034) );
  XNOR2_X1 U24142 ( .A(n22034), .B(n22523), .ZN(n22035) );
  XNOR2_X1 U24143 ( .A(n22036), .B(n22035), .ZN(n22977) );
  MUX2_X1 U24144 ( .A(n23408), .B(n23406), .S(n23252), .Z(n22051) );
  XNOR2_X1 U24146 ( .A(n22495), .B(n22037), .ZN(n22040) );
  XNOR2_X1 U24147 ( .A(n22854), .B(n3154), .ZN(n22038) );
  XNOR2_X1 U24148 ( .A(n22519), .B(n22038), .ZN(n22039) );
  XNOR2_X1 U24149 ( .A(n22040), .B(n22039), .ZN(n22979) );
  XNOR2_X1 U24150 ( .A(n22041), .B(n22511), .ZN(n22045) );
  XNOR2_X1 U24151 ( .A(n22796), .B(n22822), .ZN(n22043) );
  XNOR2_X1 U24152 ( .A(n22890), .B(n3029), .ZN(n22042) );
  XNOR2_X1 U24153 ( .A(n22043), .B(n22042), .ZN(n22044) );
  XNOR2_X1 U24154 ( .A(n22045), .B(n22044), .ZN(n23213) );
  INV_X1 U24155 ( .A(n23213), .ZN(n22980) );
  MUX2_X1 U24156 ( .A(n22979), .B(n22980), .S(n28527), .Z(n22050) );
  XNOR2_X1 U24157 ( .A(n29519), .B(n1225), .ZN(n22046) );
  XNOR2_X1 U24158 ( .A(n22046), .B(n22913), .ZN(n22047) );
  XNOR2_X1 U24159 ( .A(n22532), .B(n22047), .ZN(n22049) );
  INV_X1 U24160 ( .A(n24584), .ZN(n24581) );
  XNOR2_X1 U24161 ( .A(n29087), .B(n22187), .ZN(n22056) );
  XNOR2_X1 U24162 ( .A(n22763), .B(n3508), .ZN(n22055) );
  XNOR2_X1 U24163 ( .A(n22057), .B(n22058), .ZN(n22063) );
  XNOR2_X1 U24164 ( .A(n22059), .B(n3109), .ZN(n22060) );
  XNOR2_X1 U24165 ( .A(n22061), .B(n22060), .ZN(n22062) );
  XNOR2_X1 U24166 ( .A(n22063), .B(n22062), .ZN(n23706) );
  XNOR2_X1 U24167 ( .A(n22856), .B(n1248), .ZN(n22064) );
  XNOR2_X1 U24168 ( .A(n22065), .B(n22064), .ZN(n22071) );
  XNOR2_X1 U24169 ( .A(n22066), .B(n22067), .ZN(n22518) );
  INV_X1 U24170 ( .A(n22518), .ZN(n22069) );
  XNOR2_X1 U24171 ( .A(n22068), .B(n22104), .ZN(n22607) );
  XNOR2_X1 U24172 ( .A(n22069), .B(n22607), .ZN(n22070) );
  XNOR2_X1 U24173 ( .A(n22387), .B(n22072), .ZN(n22074) );
  XNOR2_X1 U24174 ( .A(n22074), .B(n22073), .ZN(n22075) );
  XNOR2_X1 U24175 ( .A(n22827), .B(n22075), .ZN(n22079) );
  XNOR2_X1 U24176 ( .A(n22670), .B(n22522), .ZN(n22076) );
  XNOR2_X1 U24177 ( .A(n22077), .B(n22076), .ZN(n22078) );
  XNOR2_X1 U24178 ( .A(n22079), .B(n22078), .ZN(n22451) );
  XNOR2_X1 U24180 ( .A(n22363), .B(n22094), .ZN(n22634) );
  XNOR2_X1 U24181 ( .A(n22080), .B(n22634), .ZN(n22083) );
  XNOR2_X1 U24182 ( .A(n22778), .B(n2510), .ZN(n22081) );
  XNOR2_X1 U24183 ( .A(n22081), .B(n22809), .ZN(n22082) );
  XNOR2_X1 U24185 ( .A(n22086), .B(n22542), .ZN(n22088) );
  XNOR2_X1 U24186 ( .A(n22123), .B(n28517), .ZN(n22626) );
  XNOR2_X1 U24187 ( .A(n22626), .B(n22088), .ZN(n22091) );
  XNOR2_X1 U24188 ( .A(n22664), .B(n1246), .ZN(n22089) );
  XNOR2_X1 U24189 ( .A(n22839), .B(n22089), .ZN(n22090) );
  XNOR2_X1 U24190 ( .A(n22091), .B(n22090), .ZN(n22452) );
  INV_X1 U24191 ( .A(n22452), .ZN(n23220) );
  XNOR2_X1 U24192 ( .A(n22642), .B(n22092), .ZN(n22097) );
  XNOR2_X1 U24193 ( .A(n22093), .B(n22813), .ZN(n22207) );
  XNOR2_X1 U24194 ( .A(n22094), .B(n3598), .ZN(n22095) );
  XNOR2_X1 U24195 ( .A(n22207), .B(n22095), .ZN(n22096) );
  XNOR2_X1 U24196 ( .A(n22097), .B(n22096), .ZN(n22953) );
  XNOR2_X1 U24197 ( .A(n28409), .B(n22099), .ZN(n22818) );
  XNOR2_X1 U24198 ( .A(n22100), .B(n22818), .ZN(n22103) );
  XNOR2_X1 U24199 ( .A(n22350), .B(n22101), .ZN(n22102) );
  XNOR2_X1 U24200 ( .A(n22103), .B(n22102), .ZN(n22455) );
  XNOR2_X1 U24201 ( .A(n22104), .B(n22240), .ZN(n22105) );
  XNOR2_X1 U24202 ( .A(n22341), .B(n22105), .ZN(n22109) );
  XNOR2_X1 U24203 ( .A(n22428), .B(n22605), .ZN(n22107) );
  XNOR2_X1 U24204 ( .A(n22855), .B(n26214), .ZN(n22106) );
  XNOR2_X1 U24205 ( .A(n22107), .B(n22106), .ZN(n22108) );
  XNOR2_X1 U24206 ( .A(n22109), .B(n22108), .ZN(n23843) );
  INV_X1 U24208 ( .A(n22199), .ZN(n22110) );
  XNOR2_X1 U24209 ( .A(n22313), .B(n22111), .ZN(n22115) );
  XNOR2_X1 U24210 ( .A(n22387), .B(n22295), .ZN(n22113) );
  XNOR2_X1 U24211 ( .A(n22152), .B(n1172), .ZN(n22112) );
  XNOR2_X1 U24212 ( .A(n22113), .B(n22112), .ZN(n22114) );
  XNOR2_X1 U24214 ( .A(n22589), .B(n22116), .ZN(n22842) );
  INV_X1 U24215 ( .A(n22842), .ZN(n22118) );
  XNOR2_X1 U24217 ( .A(n22731), .B(n2381), .ZN(n22119) );
  XNOR2_X1 U24218 ( .A(n22119), .B(n22650), .ZN(n22120) );
  INV_X1 U24221 ( .A(n22455), .ZN(n23722) );
  XNOR2_X1 U24222 ( .A(n22194), .B(n3662), .ZN(n22122) );
  XNOR2_X1 U24223 ( .A(n22663), .B(n22122), .ZN(n22126) );
  XNOR2_X1 U24224 ( .A(n22574), .B(n22123), .ZN(n22124) );
  XNOR2_X1 U24225 ( .A(n22318), .B(n22124), .ZN(n22125) );
  XNOR2_X1 U24226 ( .A(n22126), .B(n22125), .ZN(n22954) );
  NAND2_X1 U24227 ( .A1(n22127), .A2(n23845), .ZN(n22128) );
  INV_X1 U24229 ( .A(n24577), .ZN(n23963) );
  MUX2_X1 U24230 ( .A(n24586), .B(n22130), .S(n23963), .Z(n22179) );
  XNOR2_X1 U24231 ( .A(n22615), .B(n22270), .ZN(n22131) );
  XNOR2_X1 U24232 ( .A(n22486), .B(n22131), .ZN(n22135) );
  XNOR2_X1 U24233 ( .A(n22506), .B(n2894), .ZN(n22133) );
  XNOR2_X1 U24234 ( .A(n22571), .B(n22133), .ZN(n22134) );
  XNOR2_X1 U24235 ( .A(n22134), .B(n22135), .ZN(n22174) );
  INV_X1 U24236 ( .A(n22174), .ZN(n23710) );
  XNOR2_X1 U24237 ( .A(n22514), .B(n22240), .ZN(n22261) );
  XNOR2_X1 U24238 ( .A(n22497), .B(n22261), .ZN(n22138) );
  XNOR2_X1 U24239 ( .A(n22605), .B(n2505), .ZN(n22136) );
  XNOR2_X1 U24240 ( .A(n22854), .B(n22750), .ZN(n22558) );
  XNOR2_X1 U24241 ( .A(n22136), .B(n22558), .ZN(n22137) );
  INV_X1 U24242 ( .A(n23712), .ZN(n22971) );
  OAI21_X1 U24243 ( .B1(n22140), .B2(n5339), .A(n22139), .ZN(n22149) );
  NOR2_X1 U24244 ( .A1(n22142), .A2(n22141), .ZN(n22148) );
  NAND2_X1 U24245 ( .A1(n22146), .A2(n22143), .ZN(n22144) );
  OAI211_X1 U24246 ( .C1(n22146), .C2(n22145), .A(n22144), .B(n21624), .ZN(
        n22147) );
  XNOR2_X1 U24247 ( .A(n22295), .B(n22525), .ZN(n22150) );
  XNOR2_X1 U24248 ( .A(n22151), .B(n22150), .ZN(n22156) );
  XNOR2_X1 U24249 ( .A(n22830), .B(n29548), .ZN(n22154) );
  XNOR2_X1 U24250 ( .A(n22152), .B(n3385), .ZN(n22153) );
  XNOR2_X1 U24251 ( .A(n22154), .B(n22153), .ZN(n22155) );
  XNOR2_X1 U24252 ( .A(n22157), .B(n22474), .ZN(n22162) );
  XNOR2_X1 U24253 ( .A(n22158), .B(n2306), .ZN(n22160) );
  XNOR2_X1 U24254 ( .A(n22159), .B(n22160), .ZN(n22161) );
  XNOR2_X1 U24255 ( .A(n22162), .B(n22161), .ZN(n23262) );
  XNOR2_X1 U24257 ( .A(n22164), .B(n22461), .ZN(n22168) );
  XNOR2_X1 U24258 ( .A(n22279), .B(n22628), .ZN(n22166) );
  XNOR2_X1 U24259 ( .A(n22784), .B(n3491), .ZN(n22165) );
  XNOR2_X1 U24260 ( .A(n22166), .B(n22165), .ZN(n22167) );
  XNOR2_X1 U24261 ( .A(n22168), .B(n22167), .ZN(n23233) );
  INV_X1 U24262 ( .A(n23233), .ZN(n23585) );
  XNOR2_X1 U24263 ( .A(n22333), .B(n22169), .ZN(n22170) );
  XNOR2_X1 U24264 ( .A(n22265), .B(n2995), .ZN(n22171) );
  XNOR2_X1 U24265 ( .A(n22172), .B(n22245), .ZN(n22483) );
  OAI211_X1 U24266 ( .C1(n23716), .C2(n23585), .A(n23715), .B(n23260), .ZN(
        n22175) );
  MUX2_X1 U24267 ( .A(n24584), .B(n24054), .S(n29026), .Z(n22177) );
  XNOR2_X1 U24269 ( .A(n22713), .B(n22180), .ZN(n22182) );
  XNOR2_X1 U24270 ( .A(n22181), .B(n22182), .ZN(n22186) );
  XNOR2_X1 U24271 ( .A(n22428), .B(n22856), .ZN(n22184) );
  XNOR2_X1 U24272 ( .A(n22855), .B(Key[19]), .ZN(n22183) );
  XNOR2_X1 U24273 ( .A(n22184), .B(n22183), .ZN(n22185) );
  XNOR2_X1 U24274 ( .A(n22186), .B(n22185), .ZN(n23266) );
  XNOR2_X1 U24275 ( .A(n22188), .B(n22187), .ZN(n22191) );
  XNOR2_X1 U24276 ( .A(n22409), .B(n3673), .ZN(n22189) );
  XNOR2_X1 U24277 ( .A(n22842), .B(n22189), .ZN(n22190) );
  XNOR2_X1 U24278 ( .A(n22193), .B(n22192), .ZN(n22198) );
  XNOR2_X1 U24279 ( .A(n22664), .B(n22194), .ZN(n22837) );
  XNOR2_X1 U24280 ( .A(n22195), .B(n3695), .ZN(n22196) );
  XNOR2_X1 U24281 ( .A(n22837), .B(n22196), .ZN(n22197) );
  XNOR2_X1 U24282 ( .A(n22198), .B(n22197), .ZN(n23267) );
  XNOR2_X1 U24283 ( .A(n22828), .B(n22395), .ZN(n22203) );
  XNOR2_X1 U24284 ( .A(n22522), .B(n355), .ZN(n22201) );
  XNOR2_X1 U24285 ( .A(n22703), .B(n3633), .ZN(n22200) );
  XNOR2_X1 U24286 ( .A(n22201), .B(n22200), .ZN(n22202) );
  MUX2_X1 U24287 ( .A(n379), .B(n23217), .S(n406), .Z(n22217) );
  XNOR2_X1 U24288 ( .A(n28514), .B(n22206), .ZN(n22210) );
  XNOR2_X1 U24289 ( .A(n22434), .B(n2996), .ZN(n22208) );
  XNOR2_X1 U24290 ( .A(n22208), .B(n22207), .ZN(n22209) );
  INV_X1 U24291 ( .A(n23562), .ZN(n23615) );
  OAI22_X1 U24292 ( .A1(n23615), .A2(n406), .B1(n23267), .B2(n23266), .ZN(
        n22215) );
  XNOR2_X1 U24293 ( .A(n22488), .B(n6319), .ZN(n22211) );
  XNOR2_X1 U24294 ( .A(n22211), .B(n22418), .ZN(n22212) );
  XNOR2_X1 U24295 ( .A(n22619), .B(n28409), .ZN(n22348) );
  XNOR2_X1 U24296 ( .A(n22212), .B(n22348), .ZN(n22214) );
  XNOR2_X1 U24297 ( .A(n22213), .B(n22214), .ZN(n23611) );
  INV_X1 U24298 ( .A(n23611), .ZN(n23216) );
  NAND2_X1 U24299 ( .A1(n22215), .A2(n23216), .ZN(n22216) );
  INV_X1 U24301 ( .A(n24735), .ZN(n24280) );
  INV_X1 U24302 ( .A(n22218), .ZN(n22624) );
  INV_X1 U24304 ( .A(n22220), .ZN(n22546) );
  XNOR2_X1 U24305 ( .A(n22712), .B(n22546), .ZN(n22225) );
  XNOR2_X1 U24306 ( .A(n22221), .B(n22790), .ZN(n22223) );
  XNOR2_X1 U24307 ( .A(n22279), .B(n27956), .ZN(n22222) );
  XNOR2_X1 U24308 ( .A(n22223), .B(n22222), .ZN(n22224) );
  XNOR2_X1 U24309 ( .A(n22225), .B(n22224), .ZN(n23563) );
  XNOR2_X1 U24310 ( .A(n22226), .B(n22227), .ZN(n22772) );
  XNOR2_X1 U24311 ( .A(n22880), .B(n22772), .ZN(n22231) );
  XNOR2_X1 U24312 ( .A(n22295), .B(n22697), .ZN(n22229) );
  XNOR2_X1 U24313 ( .A(n22698), .B(n3752), .ZN(n22228) );
  XNOR2_X1 U24314 ( .A(n22229), .B(n22228), .ZN(n22230) );
  XNOR2_X1 U24315 ( .A(n22232), .B(n22601), .ZN(n22733) );
  INV_X1 U24316 ( .A(n22733), .ZN(n22233) );
  XNOR2_X1 U24317 ( .A(n22533), .B(n22233), .ZN(n22237) );
  XNOR2_X1 U24318 ( .A(n22762), .B(Key[66]), .ZN(n22234) );
  XNOR2_X1 U24319 ( .A(n22235), .B(n22234), .ZN(n22236) );
  INV_X1 U24320 ( .A(n22609), .ZN(n22239) );
  XNOR2_X1 U24321 ( .A(n22240), .B(n22239), .ZN(n22242) );
  XNOR2_X1 U24322 ( .A(n22718), .B(n2981), .ZN(n22241) );
  XNOR2_X1 U24323 ( .A(n22242), .B(n22241), .ZN(n22243) );
  XNOR2_X1 U24324 ( .A(n22633), .B(n22778), .ZN(n22247) );
  XNOR2_X1 U24325 ( .A(n22247), .B(n22897), .ZN(n22504) );
  XNOR2_X1 U24327 ( .A(n22248), .B(n22270), .ZN(n22250) );
  XNOR2_X1 U24328 ( .A(n22249), .B(n22250), .ZN(n22254) );
  XNOR2_X1 U24329 ( .A(n22724), .B(n2984), .ZN(n22251) );
  XNOR2_X1 U24330 ( .A(n22251), .B(n22252), .ZN(n22253) );
  INV_X1 U24332 ( .A(n23640), .ZN(n23314) );
  NAND2_X1 U24333 ( .A1(n2138), .A2(n23640), .ZN(n22255) );
  OAI211_X1 U24335 ( .C1(n28963), .C2(n23564), .A(n22258), .B(n22257), .ZN(
        n22311) );
  NOR2_X1 U24336 ( .A1(n24280), .A2(n22311), .ZN(n24737) );
  XNOR2_X1 U24337 ( .A(n22495), .B(n22259), .ZN(n22263) );
  XNOR2_X1 U24338 ( .A(n6504), .B(n3067), .ZN(n22260) );
  XNOR2_X1 U24339 ( .A(n22261), .B(n22260), .ZN(n22262) );
  XNOR2_X1 U24340 ( .A(n22263), .B(n22262), .ZN(n23309) );
  INV_X1 U24341 ( .A(n23309), .ZN(n23632) );
  XNOR2_X1 U24342 ( .A(n22264), .B(n22481), .ZN(n22269) );
  XNOR2_X1 U24343 ( .A(n22501), .B(n2402), .ZN(n22267) );
  XNOR2_X1 U24344 ( .A(n22265), .B(n22692), .ZN(n22266) );
  XNOR2_X1 U24345 ( .A(n22267), .B(n22266), .ZN(n22268) );
  XNOR2_X1 U24346 ( .A(n22271), .B(n22270), .ZN(n22274) );
  INV_X1 U24347 ( .A(n22272), .ZN(n22273) );
  XNOR2_X1 U24348 ( .A(n22273), .B(n22274), .ZN(n22276) );
  XNOR2_X1 U24349 ( .A(n22506), .B(n22890), .ZN(n22485) );
  XNOR2_X1 U24350 ( .A(n28492), .B(n3751), .ZN(n22275) );
  XNOR2_X1 U24352 ( .A(n22786), .B(n22278), .ZN(n22281) );
  XNOR2_X1 U24353 ( .A(n22279), .B(n22791), .ZN(n22280) );
  XNOR2_X1 U24354 ( .A(n22281), .B(n22280), .ZN(n22282) );
  XNOR2_X1 U24355 ( .A(n22283), .B(n22282), .ZN(n23630) );
  XNOR2_X1 U24356 ( .A(n22285), .B(n22525), .ZN(n22771) );
  AOI21_X1 U24357 ( .B1(n22286), .B2(n28790), .A(n22290), .ZN(n22287) );
  OAI21_X1 U24358 ( .B1(n28790), .B2(n22288), .A(n22287), .ZN(n22293) );
  NAND3_X1 U24359 ( .A1(n22291), .A2(n489), .A3(n22290), .ZN(n22292) );
  NAND3_X1 U24360 ( .A1(n22294), .A2(n22293), .A3(n22292), .ZN(n22699) );
  XNOR2_X1 U24361 ( .A(n22699), .B(n22295), .ZN(n22297) );
  XNOR2_X1 U24362 ( .A(n22671), .B(n2527), .ZN(n22296) );
  XNOR2_X1 U24363 ( .A(n22033), .B(n22394), .ZN(n22299) );
  MUX2_X1 U24364 ( .A(n23630), .B(n23558), .S(n23557), .Z(n22310) );
  XNOR2_X1 U24365 ( .A(n22300), .B(n22734), .ZN(n22304) );
  XNOR2_X1 U24366 ( .A(n22301), .B(n22302), .ZN(n22303) );
  XNOR2_X1 U24367 ( .A(n22304), .B(n22303), .ZN(n22309) );
  XNOR2_X1 U24368 ( .A(n22913), .B(n22414), .ZN(n22307) );
  INV_X1 U24369 ( .A(n22756), .ZN(n22305) );
  XNOR2_X1 U24370 ( .A(n22305), .B(n1196), .ZN(n22306) );
  XNOR2_X1 U24371 ( .A(n22307), .B(n22306), .ZN(n22308) );
  XNOR2_X1 U24372 ( .A(n22309), .B(n22308), .ZN(n23631) );
  INV_X1 U24373 ( .A(n23631), .ZN(n23629) );
  INV_X1 U24374 ( .A(n22311), .ZN(n24736) );
  XNOR2_X1 U24375 ( .A(n22312), .B(n22523), .ZN(n22314) );
  XNOR2_X1 U24376 ( .A(n22314), .B(n22313), .ZN(n22317) );
  INV_X1 U24377 ( .A(n22315), .ZN(n22316) );
  XNOR2_X1 U24378 ( .A(n22574), .B(n22625), .ZN(n22319) );
  XNOR2_X1 U24379 ( .A(n22319), .B(n22318), .ZN(n22324) );
  XNOR2_X1 U24380 ( .A(n22380), .B(n3483), .ZN(n22322) );
  XNOR2_X1 U24381 ( .A(n22379), .B(n28499), .ZN(n22321) );
  XNOR2_X1 U24382 ( .A(n22321), .B(n22322), .ZN(n22323) );
  XNOR2_X1 U24383 ( .A(n22326), .B(n22910), .ZN(n22357) );
  XNOR2_X1 U24384 ( .A(n22357), .B(n22325), .ZN(n22329) );
  OAI21_X1 U24386 ( .B1(n23761), .B2(n23762), .A(n23474), .ZN(n22346) );
  XNOR2_X1 U24387 ( .A(n22330), .B(n22644), .ZN(n22332) );
  XNOR2_X1 U24388 ( .A(n22813), .B(n3232), .ZN(n22331) );
  XNOR2_X1 U24389 ( .A(n22332), .B(n22331), .ZN(n22336) );
  XNOR2_X1 U24390 ( .A(n22333), .B(n22434), .ZN(n22635) );
  XNOR2_X1 U24391 ( .A(n22635), .B(n22362), .ZN(n22335) );
  XNOR2_X1 U24393 ( .A(n22338), .B(n22337), .ZN(n22369) );
  XNOR2_X1 U24394 ( .A(n22610), .B(n27462), .ZN(n22339) );
  XNOR2_X1 U24395 ( .A(n22339), .B(n22369), .ZN(n22345) );
  XNOR2_X1 U24396 ( .A(n22605), .B(n22340), .ZN(n22343) );
  INV_X1 U24397 ( .A(n22341), .ZN(n22342) );
  XNOR2_X1 U24398 ( .A(n22342), .B(n22343), .ZN(n22344) );
  NAND2_X1 U24400 ( .A1(n22346), .A2(n23475), .ZN(n22355) );
  NAND2_X1 U24401 ( .A1(n23762), .A2(n23760), .ZN(n22354) );
  XNOR2_X1 U24402 ( .A(n22374), .B(n22888), .ZN(n22347) );
  XNOR2_X1 U24403 ( .A(n22348), .B(n22347), .ZN(n22352) );
  XNOR2_X1 U24404 ( .A(n28483), .B(n3625), .ZN(n22349) );
  XNOR2_X1 U24405 ( .A(n22350), .B(n22349), .ZN(n22351) );
  XNOR2_X1 U24406 ( .A(n22351), .B(n22352), .ZN(n23326) );
  INV_X1 U24407 ( .A(n23762), .ZN(n23034) );
  AOI22_X1 U24409 ( .A1(n22356), .A2(n24735), .B1(n24736), .B2(n24602), .ZN(
        n22450) );
  XNOR2_X1 U24410 ( .A(n22735), .B(n26531), .ZN(n22359) );
  XNOR2_X1 U24411 ( .A(n22358), .B(n22359), .ZN(n22360) );
  XNOR2_X1 U24412 ( .A(n22689), .B(n22362), .ZN(n22367) );
  XNOR2_X1 U24413 ( .A(n22363), .B(n22812), .ZN(n22365) );
  XNOR2_X1 U24414 ( .A(n21728), .B(n1119), .ZN(n22364) );
  XNOR2_X1 U24415 ( .A(n22365), .B(n22364), .ZN(n22366) );
  XNOR2_X1 U24416 ( .A(n22369), .B(n22368), .ZN(n22373) );
  XNOR2_X1 U24417 ( .A(n22370), .B(n22553), .ZN(n22371) );
  XNOR2_X1 U24418 ( .A(n22607), .B(n22371), .ZN(n22372) );
  XNOR2_X1 U24419 ( .A(n22372), .B(n22373), .ZN(n23620) );
  NAND2_X1 U24420 ( .A1(n23621), .A2(n23620), .ZN(n23273) );
  XNOR2_X1 U24421 ( .A(n22374), .B(n3660), .ZN(n22375) );
  XNOR2_X1 U24422 ( .A(n22617), .B(n22375), .ZN(n22378) );
  XNOR2_X1 U24423 ( .A(n22796), .B(n22888), .ZN(n22376) );
  XNOR2_X1 U24424 ( .A(n22727), .B(n22376), .ZN(n22377) );
  XNOR2_X1 U24425 ( .A(n22377), .B(n22378), .ZN(n23619) );
  INV_X1 U24426 ( .A(n23619), .ZN(n22987) );
  OAI21_X1 U24427 ( .B1(n23620), .B2(n22987), .A(n23273), .ZN(n22392) );
  XNOR2_X1 U24428 ( .A(n22379), .B(n22380), .ZN(n22381) );
  XNOR2_X1 U24429 ( .A(n22626), .B(n22381), .ZN(n22385) );
  XNOR2_X1 U24430 ( .A(n22383), .B(n22382), .ZN(n22384) );
  NAND2_X1 U24432 ( .A1(n23622), .A2(n23566), .ZN(n22391) );
  XNOR2_X1 U24433 ( .A(n22386), .B(n22584), .ZN(n22389) );
  XNOR2_X1 U24434 ( .A(n22387), .B(n3722), .ZN(n22388) );
  INV_X1 U24435 ( .A(n23618), .ZN(n23567) );
  OAI21_X1 U24436 ( .B1(n23622), .B2(n23273), .A(n22393), .ZN(n24739) );
  INV_X1 U24437 ( .A(n24739), .ZN(n24282) );
  AND2_X1 U24438 ( .A1(n3310), .A2(n22311), .ZN(n24603) );
  INV_X1 U24439 ( .A(n22396), .ZN(n22400) );
  NAND2_X1 U24440 ( .A1(n22402), .A2(n22397), .ZN(n22399) );
  AOI21_X1 U24441 ( .B1(n22400), .B2(n22399), .A(n22398), .ZN(n22406) );
  OAI21_X1 U24442 ( .B1(n6940), .B2(n22404), .A(n22403), .ZN(n22405) );
  NOR2_X1 U24443 ( .A1(n22406), .A2(n22405), .ZN(n22407) );
  INV_X1 U24444 ( .A(n22581), .ZN(n22408) );
  INV_X1 U24445 ( .A(n23049), .ZN(n23472) );
  XNOR2_X1 U24446 ( .A(n22759), .B(n22409), .ZN(n22413) );
  XNOR2_X1 U24447 ( .A(n22414), .B(n22473), .ZN(n22415) );
  XNOR2_X1 U24448 ( .A(n28162), .B(n22415), .ZN(n22416) );
  XNOR2_X1 U24449 ( .A(n22418), .B(n2577), .ZN(n22421) );
  XNOR2_X1 U24450 ( .A(n22567), .B(n22419), .ZN(n22420) );
  XNOR2_X1 U24451 ( .A(n22421), .B(n22420), .ZN(n22425) );
  XNOR2_X1 U24452 ( .A(n22422), .B(n22619), .ZN(n22423) );
  XNOR2_X1 U24453 ( .A(n22423), .B(n22571), .ZN(n22424) );
  XNOR2_X1 U24454 ( .A(n22610), .B(n29562), .ZN(n22430) );
  XNOR2_X1 U24455 ( .A(n29490), .B(n22427), .ZN(n22429) );
  INV_X1 U24456 ( .A(n3378), .ZN(n26545) );
  XNOR2_X1 U24457 ( .A(n22556), .B(n26545), .ZN(n22431) );
  XNOR2_X1 U24458 ( .A(n22558), .B(n22431), .ZN(n22432) );
  OAI21_X1 U24459 ( .B1(n23318), .B2(n23472), .A(n22433), .ZN(n23473) );
  INV_X1 U24460 ( .A(n23473), .ZN(n22448) );
  XNOR2_X1 U24461 ( .A(n22561), .B(n22434), .ZN(n22435) );
  XNOR2_X1 U24462 ( .A(n22436), .B(n22435), .ZN(n22440) );
  XNOR2_X1 U24463 ( .A(n22690), .B(n22437), .ZN(n22780) );
  XNOR2_X1 U24464 ( .A(n22479), .B(n1046), .ZN(n22438) );
  XNOR2_X1 U24465 ( .A(n22780), .B(n22438), .ZN(n22439) );
  XNOR2_X1 U24466 ( .A(n22784), .B(n3422), .ZN(n22441) );
  XNOR2_X1 U24467 ( .A(n22443), .B(n22442), .ZN(n22446) );
  XNOR2_X1 U24468 ( .A(n22464), .B(n22787), .ZN(n22444) );
  XNOR2_X1 U24469 ( .A(n22444), .B(n22625), .ZN(n22445) );
  XNOR2_X1 U24470 ( .A(n22446), .B(n22445), .ZN(n23648) );
  AOI22_X1 U24471 ( .A1(n24744), .A2(n24604), .B1(n24603), .B2(n24734), .ZN(
        n22449) );
  OAI21_X1 U24472 ( .B1(n24737), .B2(n22450), .A(n22449), .ZN(n25428) );
  XNOR2_X1 U24473 ( .A(n26044), .B(n25428), .ZN(n25803) );
  XNOR2_X1 U24474 ( .A(n24885), .B(n25803), .ZN(n22943) );
  OAI21_X1 U24476 ( .B1(n29618), .B2(n23700), .A(n23705), .ZN(n22453) );
  NOR2_X1 U24477 ( .A1(n22953), .A2(n22455), .ZN(n23396) );
  NOR2_X1 U24478 ( .A1(n23396), .A2(n23726), .ZN(n22458) );
  NOR2_X1 U24479 ( .A1(n28484), .A2(n23843), .ZN(n22456) );
  AOI22_X1 U24480 ( .A1(n23396), .A2(n23845), .B1(n22456), .B2(n22455), .ZN(
        n22457) );
  XNOR2_X1 U24482 ( .A(n22791), .B(n3607), .ZN(n22460) );
  XNOR2_X1 U24483 ( .A(n22460), .B(n22459), .ZN(n22462) );
  XNOR2_X1 U24484 ( .A(n22462), .B(n22461), .ZN(n22466) );
  XNOR2_X1 U24485 ( .A(n22464), .B(n28450), .ZN(n22666) );
  XNOR2_X1 U24486 ( .A(n22923), .B(n22666), .ZN(n22465) );
  XNOR2_X1 U24487 ( .A(n22703), .B(n2889), .ZN(n22467) );
  XNOR2_X1 U24488 ( .A(n22671), .B(n29514), .ZN(n22469) );
  XNOR2_X1 U24489 ( .A(n22472), .B(n22473), .ZN(n22652) );
  XNOR2_X1 U24490 ( .A(n22652), .B(n22474), .ZN(n22478) );
  XNOR2_X1 U24491 ( .A(n22913), .B(n22735), .ZN(n22476) );
  XNOR2_X1 U24492 ( .A(n28486), .B(n26665), .ZN(n22475) );
  XNOR2_X1 U24493 ( .A(n22476), .B(n22475), .ZN(n22477) );
  INV_X1 U24494 ( .A(n22494), .ZN(n23837) );
  XNOR2_X1 U24496 ( .A(n22479), .B(n3114), .ZN(n22480) );
  XNOR2_X1 U24497 ( .A(n22480), .B(n21789), .ZN(n22482) );
  XNOR2_X1 U24498 ( .A(n22481), .B(n22482), .ZN(n22484) );
  XNOR2_X1 U24499 ( .A(n22485), .B(n22486), .ZN(n22493) );
  XNOR2_X1 U24500 ( .A(n22487), .B(n22488), .ZN(n22491) );
  XNOR2_X1 U24501 ( .A(n22657), .B(n22489), .ZN(n22490) );
  XNOR2_X1 U24502 ( .A(n22491), .B(n22490), .ZN(n22492) );
  XNOR2_X1 U24503 ( .A(n22493), .B(n22492), .ZN(n23078) );
  INV_X1 U24504 ( .A(n23078), .ZN(n23390) );
  XNOR2_X1 U24505 ( .A(n22514), .B(n22713), .ZN(n22496) );
  XNOR2_X1 U24506 ( .A(n22556), .B(n3191), .ZN(n22498) );
  NAND3_X1 U24507 ( .A1(n28460), .A2(n23839), .A3(n28418), .ZN(n22499) );
  MUX2_X1 U24508 ( .A(n24614), .B(n24610), .S(n29109), .Z(n22640) );
  XNOR2_X1 U24509 ( .A(n22503), .B(n22502), .ZN(n22505) );
  XNOR2_X1 U24510 ( .A(n22891), .B(n22724), .ZN(n22508) );
  XNOR2_X1 U24511 ( .A(n22506), .B(n3654), .ZN(n22507) );
  XNOR2_X1 U24512 ( .A(n22508), .B(n22507), .ZN(n22513) );
  XNOR2_X1 U24513 ( .A(n1858), .B(n22509), .ZN(n22510) );
  XNOR2_X1 U24514 ( .A(n22514), .B(n22609), .ZN(n22517) );
  XNOR2_X1 U24515 ( .A(n22515), .B(n5059), .ZN(n22516) );
  XNOR2_X1 U24516 ( .A(n22517), .B(n22516), .ZN(n22521) );
  XNOR2_X1 U24517 ( .A(n22519), .B(n22518), .ZN(n22520) );
  XNOR2_X1 U24518 ( .A(n22520), .B(n22521), .ZN(n23295) );
  MUX2_X1 U24519 ( .A(n22531), .B(n23077), .S(n23295), .Z(n22552) );
  XNOR2_X1 U24520 ( .A(n22523), .B(n22522), .ZN(n22884) );
  XNOR2_X1 U24521 ( .A(n22884), .B(n22524), .ZN(n22530) );
  XNOR2_X1 U24522 ( .A(n22526), .B(n22525), .ZN(n22528) );
  XNOR2_X1 U24523 ( .A(n22698), .B(n3493), .ZN(n22527) );
  XNOR2_X1 U24524 ( .A(n22528), .B(n22527), .ZN(n22529) );
  INV_X1 U24525 ( .A(n23297), .ZN(n22962) );
  INV_X1 U24526 ( .A(n23295), .ZN(n23832) );
  XNOR2_X1 U24527 ( .A(n22532), .B(n22533), .ZN(n22540) );
  XNOR2_X1 U24528 ( .A(n28486), .B(n22534), .ZN(n22538) );
  INV_X1 U24529 ( .A(n22601), .ZN(n22536) );
  XNOR2_X1 U24530 ( .A(n22536), .B(n22535), .ZN(n22537) );
  XNOR2_X1 U24531 ( .A(n22537), .B(n22538), .ZN(n22539) );
  NAND2_X1 U24532 ( .A1(n23832), .A2(n29602), .ZN(n22541) );
  NOR2_X1 U24533 ( .A1(n23833), .A2(n22541), .ZN(n22550) );
  NOR2_X1 U24534 ( .A1(n29020), .A2(n29602), .ZN(n22549) );
  XNOR2_X1 U24535 ( .A(n22624), .B(n22542), .ZN(n22544) );
  XNOR2_X1 U24536 ( .A(n22791), .B(n3528), .ZN(n22543) );
  XNOR2_X1 U24537 ( .A(n22544), .B(n22543), .ZN(n22548) );
  XNOR2_X1 U24538 ( .A(n22546), .B(n22545), .ZN(n22547) );
  XNOR2_X1 U24539 ( .A(n22547), .B(n22548), .ZN(n22864) );
  INV_X1 U24540 ( .A(n23831), .ZN(n23296) );
  OAI21_X1 U24541 ( .B1(n22550), .B2(n22549), .A(n23298), .ZN(n22551) );
  OAI21_X1 U24542 ( .B1(n22552), .B2(n22962), .A(n22551), .ZN(n24017) );
  XNOR2_X1 U24543 ( .A(n22180), .B(n22553), .ZN(n22554) );
  XNOR2_X1 U24544 ( .A(n22555), .B(n22554), .ZN(n22560) );
  XNOR2_X1 U24545 ( .A(n22556), .B(n1184), .ZN(n22557) );
  XNOR2_X1 U24546 ( .A(n22558), .B(n22557), .ZN(n22559) );
  XNOR2_X1 U24548 ( .A(n22813), .B(n2325), .ZN(n22562) );
  XNOR2_X1 U24550 ( .A(n22567), .B(n22568), .ZN(n22655) );
  XNOR2_X1 U24551 ( .A(n22569), .B(n22655), .ZN(n22573) );
  XNOR2_X1 U24552 ( .A(n28409), .B(n3003), .ZN(n22570) );
  XNOR2_X1 U24553 ( .A(n22571), .B(n22570), .ZN(n22572) );
  XNOR2_X1 U24554 ( .A(n22575), .B(n22838), .ZN(n22580) );
  INV_X1 U24555 ( .A(n22790), .ZN(n22576) );
  XNOR2_X1 U24556 ( .A(n22576), .B(n3180), .ZN(n22577) );
  XNOR2_X1 U24557 ( .A(n22578), .B(n22577), .ZN(n22579) );
  XNOR2_X2 U24558 ( .A(n22579), .B(n22580), .ZN(n23382) );
  XNOR2_X1 U24559 ( .A(n22582), .B(n22581), .ZN(n22586) );
  INV_X1 U24560 ( .A(n22829), .ZN(n22881) );
  XNOR2_X1 U24561 ( .A(n22881), .B(n3457), .ZN(n22583) );
  XNOR2_X1 U24562 ( .A(n22584), .B(n22583), .ZN(n22585) );
  XNOR2_X1 U24563 ( .A(n22586), .B(n22585), .ZN(n22946) );
  XNOR2_X1 U24564 ( .A(n22589), .B(n28589), .ZN(n22591) );
  XNOR2_X1 U24565 ( .A(n22410), .B(n2541), .ZN(n22590) );
  MUX2_X1 U24566 ( .A(n24017), .B(n29109), .S(n24612), .Z(n22639) );
  XNOR2_X1 U24567 ( .A(n22596), .B(n22595), .ZN(n22597) );
  XNOR2_X1 U24568 ( .A(n22598), .B(n22597), .ZN(n22742) );
  INV_X1 U24569 ( .A(n22599), .ZN(n22909) );
  XNOR2_X1 U24570 ( .A(n22909), .B(n22600), .ZN(n22604) );
  XNOR2_X1 U24571 ( .A(n22601), .B(n3015), .ZN(n22602) );
  XNOR2_X1 U24572 ( .A(n22325), .B(n22602), .ZN(n22603) );
  XNOR2_X1 U24574 ( .A(n22605), .B(n22606), .ZN(n22608) );
  XNOR2_X1 U24575 ( .A(n22607), .B(n22608), .ZN(n22614) );
  XNOR2_X1 U24576 ( .A(n22610), .B(n2982), .ZN(n22611) );
  XNOR2_X1 U24577 ( .A(n22611), .B(n22612), .ZN(n22613) );
  XNOR2_X1 U24578 ( .A(n22613), .B(n22614), .ZN(n23810) );
  XNOR2_X1 U24579 ( .A(n22615), .B(n3644), .ZN(n22616) );
  XNOR2_X1 U24580 ( .A(n22617), .B(n22616), .ZN(n22623) );
  XNOR2_X1 U24581 ( .A(n22618), .B(n22619), .ZN(n22621) );
  XNOR2_X1 U24582 ( .A(n22620), .B(n22621), .ZN(n22622) );
  XNOR2_X1 U24583 ( .A(n22624), .B(n22625), .ZN(n22627) );
  XNOR2_X1 U24584 ( .A(n22626), .B(n22627), .ZN(n22631) );
  XNOR2_X1 U24585 ( .A(n22628), .B(n27452), .ZN(n22629) );
  XNOR2_X1 U24586 ( .A(n22922), .B(n22629), .ZN(n22630) );
  XNOR2_X1 U24587 ( .A(n22630), .B(n22631), .ZN(n23285) );
  XNOR2_X1 U24588 ( .A(n22635), .B(n22634), .ZN(n22636) );
  XNOR2_X1 U24589 ( .A(n22637), .B(n22636), .ZN(n22877) );
  INV_X1 U24590 ( .A(n22877), .ZN(n23074) );
  MUX2_X1 U24591 ( .A(n22640), .B(n22639), .S(n5137), .Z(n25727) );
  XNOR2_X1 U24592 ( .A(n22641), .B(n22642), .ZN(n22648) );
  XNOR2_X1 U24593 ( .A(n22811), .B(n22643), .ZN(n22646) );
  XNOR2_X1 U24594 ( .A(n22644), .B(n1887), .ZN(n22645) );
  XNOR2_X1 U24595 ( .A(n22646), .B(n22645), .ZN(n22647) );
  XNOR2_X1 U24596 ( .A(n22844), .B(n857), .ZN(n22649) );
  XNOR2_X1 U24597 ( .A(n22650), .B(n22649), .ZN(n22654) );
  XNOR2_X1 U24598 ( .A(n22651), .B(n22652), .ZN(n22653) );
  XNOR2_X1 U24599 ( .A(n22656), .B(n22820), .ZN(n22659) );
  XNOR2_X1 U24600 ( .A(n28492), .B(n3697), .ZN(n22658) );
  XNOR2_X1 U24601 ( .A(n22659), .B(n22658), .ZN(n22660) );
  MUX2_X1 U24602 ( .A(n1829), .B(n22686), .S(n408), .Z(n22676) );
  XNOR2_X1 U24603 ( .A(n22661), .B(n29079), .ZN(n22662) );
  XNOR2_X1 U24604 ( .A(n22663), .B(n22662), .ZN(n22667) );
  XNOR2_X1 U24605 ( .A(n22664), .B(n27225), .ZN(n22665) );
  XNOR2_X1 U24606 ( .A(n22668), .B(n3537), .ZN(n22669) );
  XNOR2_X1 U24607 ( .A(n22670), .B(n22669), .ZN(n22673) );
  XNOR2_X1 U24608 ( .A(n22768), .B(n22671), .ZN(n22672) );
  XNOR2_X1 U24609 ( .A(n22673), .B(n22672), .ZN(n22674) );
  XNOR2_X1 U24610 ( .A(n22674), .B(n22675), .ZN(n23302) );
  INV_X1 U24611 ( .A(n22678), .ZN(n22679) );
  XNOR2_X1 U24612 ( .A(n22679), .B(n22680), .ZN(n22683) );
  XNOR2_X1 U24613 ( .A(n22681), .B(n22856), .ZN(n22682) );
  XNOR2_X1 U24614 ( .A(n22683), .B(n22682), .ZN(n22685) );
  XNOR2_X1 U24615 ( .A(n22685), .B(n22684), .ZN(n23433) );
  XNOR2_X1 U24616 ( .A(n22688), .B(n22689), .ZN(n22696) );
  XNOR2_X1 U24617 ( .A(n22691), .B(n22690), .ZN(n22694) );
  XNOR2_X1 U24618 ( .A(n22692), .B(n1161), .ZN(n22693) );
  XNOR2_X1 U24619 ( .A(n22694), .B(n22693), .ZN(n22695) );
  INV_X1 U24621 ( .A(n23450), .ZN(n23447) );
  XNOR2_X1 U24622 ( .A(n22697), .B(n22033), .ZN(n22702) );
  XNOR2_X1 U24625 ( .A(n22701), .B(n22702), .ZN(n22709) );
  XNOR2_X1 U24626 ( .A(n22703), .B(n22387), .ZN(n22707) );
  XNOR2_X1 U24627 ( .A(n22707), .B(n22706), .ZN(n22708) );
  XNOR2_X1 U24628 ( .A(n22784), .B(n3223), .ZN(n22711) );
  XNOR2_X1 U24629 ( .A(n22713), .B(n22903), .ZN(n22715) );
  XNOR2_X1 U24630 ( .A(n22715), .B(n22714), .ZN(n22722) );
  XNOR2_X1 U24631 ( .A(n22717), .B(n29591), .ZN(n22720) );
  XNOR2_X1 U24632 ( .A(n22718), .B(n3414), .ZN(n22719) );
  XNOR2_X1 U24633 ( .A(n22720), .B(n22719), .ZN(n22721) );
  XNOR2_X1 U24634 ( .A(n22722), .B(n22721), .ZN(n22935) );
  INV_X1 U24635 ( .A(n22935), .ZN(n23109) );
  AOI22_X1 U24636 ( .A1(n23447), .A2(n23442), .B1(n23370), .B2(n23109), .ZN(
        n22741) );
  XNOR2_X1 U24637 ( .A(n22723), .B(n28693), .ZN(n22726) );
  XNOR2_X1 U24638 ( .A(n22724), .B(n22890), .ZN(n22725) );
  XNOR2_X1 U24639 ( .A(n22725), .B(n22726), .ZN(n22730) );
  XNOR2_X2 U24640 ( .A(n22729), .B(n22730), .ZN(n23445) );
  XNOR2_X1 U24641 ( .A(n22731), .B(n28162), .ZN(n22732) );
  XNOR2_X1 U24642 ( .A(n22732), .B(n22733), .ZN(n22739) );
  XNOR2_X1 U24643 ( .A(n22735), .B(n22734), .ZN(n22737) );
  XNOR2_X1 U24644 ( .A(n22913), .B(n3196), .ZN(n22736) );
  XNOR2_X1 U24645 ( .A(n22736), .B(n22737), .ZN(n22738) );
  INV_X1 U24646 ( .A(n24552), .ZN(n23205) );
  INV_X1 U24647 ( .A(n23809), .ZN(n23075) );
  INV_X1 U24648 ( .A(n24551), .ZN(n22746) );
  NOR2_X1 U24649 ( .A1(n22747), .A2(n22746), .ZN(n22872) );
  XNOR2_X1 U24650 ( .A(n22748), .B(n22749), .ZN(n22754) );
  XNOR2_X1 U24651 ( .A(n22750), .B(n2385), .ZN(n22751) );
  XNOR2_X1 U24652 ( .A(n22752), .B(n22751), .ZN(n22753) );
  XNOR2_X1 U24653 ( .A(n22754), .B(n22753), .ZN(n23099) );
  XNOR2_X1 U24654 ( .A(n22756), .B(n22755), .ZN(n22758) );
  XNOR2_X1 U24655 ( .A(n22759), .B(n22760), .ZN(n22761) );
  XNOR2_X1 U24656 ( .A(n22763), .B(n28589), .ZN(n22764) );
  XNOR2_X1 U24657 ( .A(n28162), .B(n22764), .ZN(n22766) );
  XNOR2_X2 U24658 ( .A(n22767), .B(n22766), .ZN(n23419) );
  XNOR2_X1 U24659 ( .A(n22769), .B(n22768), .ZN(n22770) );
  XNOR2_X1 U24660 ( .A(n22770), .B(n22771), .ZN(n22775) );
  XNOR2_X1 U24661 ( .A(n22773), .B(n22772), .ZN(n22774) );
  XNOR2_X1 U24662 ( .A(n22777), .B(n22776), .ZN(n22782) );
  XNOR2_X1 U24663 ( .A(n22778), .B(n3244), .ZN(n22779) );
  XNOR2_X1 U24664 ( .A(n22780), .B(n22779), .ZN(n22781) );
  XNOR2_X1 U24665 ( .A(n22782), .B(n22781), .ZN(n23073) );
  INV_X1 U24666 ( .A(n23073), .ZN(n23417) );
  XNOR2_X1 U24667 ( .A(n22785), .B(n22784), .ZN(n22789) );
  XNOR2_X1 U24668 ( .A(n22787), .B(n22786), .ZN(n22788) );
  XNOR2_X1 U24669 ( .A(n22789), .B(n22788), .ZN(n22795) );
  XNOR2_X1 U24670 ( .A(n22791), .B(n22790), .ZN(n22793) );
  XNOR2_X1 U24671 ( .A(n22792), .B(n22793), .ZN(n22794) );
  INV_X1 U24672 ( .A(n22796), .ZN(n22797) );
  XNOR2_X1 U24673 ( .A(n22797), .B(n22798), .ZN(n22799) );
  XNOR2_X1 U24674 ( .A(n22799), .B(n22800), .ZN(n22804) );
  XNOR2_X1 U24675 ( .A(n1859), .B(n3164), .ZN(n22802) );
  XNOR2_X1 U24676 ( .A(n22801), .B(n22802), .ZN(n22803) );
  NAND2_X1 U24677 ( .A1(n480), .A2(n23418), .ZN(n22805) );
  MUX2_X1 U24678 ( .A(n22806), .B(n22805), .S(n23415), .Z(n22807) );
  NOR2_X1 U24680 ( .A1(n24556), .A2(n24552), .ZN(n23207) );
  INV_X1 U24681 ( .A(n23207), .ZN(n22870) );
  XNOR2_X1 U24682 ( .A(n22810), .B(n22809), .ZN(n22817) );
  XNOR2_X1 U24683 ( .A(n22811), .B(n22812), .ZN(n22815) );
  XNOR2_X1 U24684 ( .A(n22813), .B(n2446), .ZN(n22814) );
  XNOR2_X1 U24685 ( .A(n22815), .B(n22814), .ZN(n22816) );
  XNOR2_X1 U24686 ( .A(n22819), .B(n22818), .ZN(n22826) );
  XNOR2_X1 U24687 ( .A(n22820), .B(n22821), .ZN(n22824) );
  XNOR2_X1 U24688 ( .A(n22822), .B(n2973), .ZN(n22823) );
  XNOR2_X1 U24689 ( .A(n22824), .B(n22823), .ZN(n22825) );
  XNOR2_X1 U24690 ( .A(n22826), .B(n22825), .ZN(n22931) );
  NOR2_X1 U24691 ( .A1(n23820), .A2(n22931), .ZN(n22851) );
  XNOR2_X1 U24692 ( .A(n22828), .B(n22827), .ZN(n22834) );
  XNOR2_X1 U24693 ( .A(n355), .B(n22882), .ZN(n22832) );
  XNOR2_X1 U24694 ( .A(n22830), .B(n26909), .ZN(n22831) );
  XNOR2_X1 U24695 ( .A(n22832), .B(n22831), .ZN(n22833) );
  XNOR2_X1 U24696 ( .A(n22835), .B(n2946), .ZN(n22836) );
  XNOR2_X1 U24697 ( .A(n22837), .B(n22836), .ZN(n22841) );
  XNOR2_X1 U24699 ( .A(n22842), .B(n22843), .ZN(n22850) );
  XNOR2_X1 U24700 ( .A(n22844), .B(n22845), .ZN(n22848) );
  XNOR2_X1 U24701 ( .A(n22410), .B(n3256), .ZN(n22847) );
  XNOR2_X1 U24702 ( .A(n22848), .B(n22847), .ZN(n22849) );
  XNOR2_X1 U24703 ( .A(n22852), .B(n22902), .ZN(n22860) );
  INV_X1 U24704 ( .A(n2509), .ZN(n22853) );
  XNOR2_X1 U24705 ( .A(n22854), .B(n22853), .ZN(n22858) );
  XNOR2_X1 U24706 ( .A(n22856), .B(n22855), .ZN(n22857) );
  XNOR2_X1 U24707 ( .A(n22858), .B(n22857), .ZN(n22859) );
  XNOR2_X1 U24708 ( .A(n22860), .B(n22859), .ZN(n23291) );
  MUX2_X1 U24709 ( .A(n23290), .B(n23291), .S(n28182), .Z(n22861) );
  INV_X1 U24710 ( .A(n22864), .ZN(n23835) );
  NAND2_X1 U24711 ( .A1(n23835), .A2(n29602), .ZN(n22865) );
  AOI21_X1 U24712 ( .B1(n22865), .B2(n23295), .A(n23833), .ZN(n22866) );
  INV_X1 U24714 ( .A(n24555), .ZN(n24178) );
  OAI22_X1 U24715 ( .A1(n22870), .A2(n22869), .B1(n22868), .B2(n24178), .ZN(
        n22871) );
  XNOR2_X1 U24716 ( .A(n28576), .B(n25727), .ZN(n22941) );
  NOR2_X1 U24717 ( .A1(n1829), .A2(n23433), .ZN(n22874) );
  NOR2_X1 U24718 ( .A1(n23302), .A2(n4020), .ZN(n22873) );
  MUX2_X1 U24719 ( .A(n22874), .B(n22873), .S(n23431), .Z(n22876) );
  INV_X1 U24720 ( .A(n23430), .ZN(n23301) );
  INV_X1 U24721 ( .A(n24592), .ZN(n23929) );
  XNOR2_X1 U24722 ( .A(n22879), .B(n22880), .ZN(n22885) );
  XNOR2_X1 U24723 ( .A(n22881), .B(n3482), .ZN(n22883) );
  INV_X1 U24724 ( .A(n23145), .ZN(n23465) );
  INV_X1 U24725 ( .A(n22886), .ZN(n22895) );
  XNOR2_X1 U24726 ( .A(n22887), .B(n27231), .ZN(n22889) );
  XNOR2_X1 U24727 ( .A(n22889), .B(n22888), .ZN(n22893) );
  XNOR2_X1 U24728 ( .A(n22891), .B(n22890), .ZN(n22892) );
  XNOR2_X1 U24729 ( .A(n22893), .B(n22892), .ZN(n22894) );
  XNOR2_X1 U24730 ( .A(n22895), .B(n22894), .ZN(n23148) );
  XNOR2_X1 U24731 ( .A(n22898), .B(n1923), .ZN(n22900) );
  XNOR2_X1 U24732 ( .A(n22900), .B(n22899), .ZN(n22901) );
  XNOR2_X1 U24733 ( .A(n22903), .B(n2523), .ZN(n22904) );
  XNOR2_X1 U24734 ( .A(n22905), .B(n22904), .ZN(n22906) );
  XNOR2_X1 U24735 ( .A(n22907), .B(n22906), .ZN(n23454) );
  AOI21_X1 U24736 ( .B1(n23455), .B2(n23456), .A(n23454), .ZN(n22926) );
  XNOR2_X1 U24737 ( .A(n22909), .B(n22908), .ZN(n22917) );
  INV_X1 U24738 ( .A(n28472), .ZN(n22911) );
  XNOR2_X1 U24739 ( .A(n22912), .B(n22911), .ZN(n22915) );
  XNOR2_X1 U24740 ( .A(n22913), .B(n2411), .ZN(n22914) );
  XNOR2_X1 U24741 ( .A(n22915), .B(n22914), .ZN(n22916) );
  NOR2_X1 U24742 ( .A1(n23454), .A2(n23148), .ZN(n22925) );
  XNOR2_X1 U24743 ( .A(n22919), .B(n22918), .ZN(n22921) );
  XNOR2_X1 U24744 ( .A(n22921), .B(n22920), .ZN(n22924) );
  NOR2_X1 U24745 ( .A1(n23099), .A2(n23073), .ZN(n22927) );
  MUX2_X1 U24746 ( .A(n22928), .B(n22927), .S(n23419), .Z(n22930) );
  INV_X1 U24749 ( .A(n24593), .ZN(n23853) );
  NOR2_X1 U24750 ( .A1(n23289), .A2(n28182), .ZN(n22934) );
  NOR2_X1 U24753 ( .A1(n23290), .A2(n28609), .ZN(n23818) );
  AND3_X1 U24754 ( .A1(n22931), .A2(n28609), .A3(n23291), .ZN(n22932) );
  NOR2_X1 U24755 ( .A1(n23818), .A2(n22932), .ZN(n22933) );
  OAI21_X1 U24756 ( .B1(n22934), .B2(n23090), .A(n22933), .ZN(n24141) );
  INV_X1 U24757 ( .A(n23442), .ZN(n23446) );
  MUX2_X1 U24758 ( .A(n292), .B(n23446), .S(n29296), .Z(n22939) );
  NAND2_X1 U24759 ( .A1(n23370), .A2(n292), .ZN(n22937) );
  NAND2_X1 U24760 ( .A1(n23445), .A2(n23449), .ZN(n22936) );
  MUX2_X1 U24761 ( .A(n22937), .B(n22936), .S(n23442), .Z(n22938) );
  XNOR2_X1 U24762 ( .A(n25369), .B(n3527), .ZN(n22940) );
  XNOR2_X1 U24763 ( .A(n22941), .B(n22940), .ZN(n22942) );
  NOR2_X1 U24765 ( .A1(n885), .A2(n23382), .ZN(n22945) );
  NOR2_X1 U24766 ( .A1(n24542), .A2(n2823), .ZN(n22952) );
  INV_X1 U24767 ( .A(n23733), .ZN(n23257) );
  AOI21_X1 U24768 ( .B1(n23399), .B2(n23228), .A(n23257), .ZN(n22951) );
  NOR2_X1 U24769 ( .A1(n22949), .A2(n23736), .ZN(n23401) );
  INV_X1 U24770 ( .A(n24001), .ZN(n24541) );
  NOR2_X1 U24771 ( .A1(n22952), .A2(n24541), .ZN(n22970) );
  INV_X1 U24772 ( .A(n22953), .ZN(n23721) );
  INV_X1 U24773 ( .A(n22954), .ZN(n23849) );
  INV_X1 U24774 ( .A(n23843), .ZN(n23720) );
  NOR2_X1 U24775 ( .A1(n23846), .A2(n23720), .ZN(n22955) );
  NAND2_X1 U24776 ( .A1(n23846), .A2(n28484), .ZN(n23724) );
  INV_X1 U24777 ( .A(n24547), .ZN(n22969) );
  MUX2_X1 U24778 ( .A(n6279), .B(n23839), .S(n487), .Z(n22961) );
  NAND2_X1 U24780 ( .A1(n28551), .A2(n23839), .ZN(n22959) );
  NAND2_X1 U24781 ( .A1(n23280), .A2(n23078), .ZN(n22958) );
  NAND2_X1 U24782 ( .A1(n22962), .A2(n23831), .ZN(n22964) );
  NAND2_X1 U24783 ( .A1(n23832), .A2(n23077), .ZN(n22963) );
  NAND2_X1 U24784 ( .A1(n22531), .A2(n23077), .ZN(n23294) );
  NAND2_X1 U24785 ( .A1(n23294), .A2(n23832), .ZN(n22965) );
  NOR2_X1 U24786 ( .A1(n24547), .A2(n24019), .ZN(n22967) );
  NAND2_X1 U24787 ( .A1(n24538), .A2(n24001), .ZN(n23127) );
  INV_X1 U24788 ( .A(n22972), .ZN(n22975) );
  OAI21_X1 U24789 ( .B1(n23260), .B2(n22971), .A(n380), .ZN(n22974) );
  NAND2_X1 U24790 ( .A1(n23585), .A2(n23587), .ZN(n23586) );
  MUX2_X1 U24791 ( .A(n23586), .B(n22972), .S(n23716), .Z(n22973) );
  NOR2_X1 U24792 ( .A1(n22977), .A2(n22976), .ZN(n23251) );
  INV_X1 U24793 ( .A(n23251), .ZN(n22978) );
  NAND2_X1 U24794 ( .A1(n22980), .A2(n22979), .ZN(n23747) );
  NAND2_X1 U24795 ( .A1(n22980), .A2(n28527), .ZN(n22981) );
  AOI21_X1 U24796 ( .B1(n22979), .B2(n22981), .A(n23252), .ZN(n22982) );
  INV_X1 U24798 ( .A(n22984), .ZN(n23208) );
  INV_X1 U24799 ( .A(n23245), .ZN(n23604) );
  INV_X1 U24800 ( .A(n23621), .ZN(n23270) );
  NAND2_X1 U24801 ( .A1(n23270), .A2(n22987), .ZN(n23624) );
  OR2_X1 U24802 ( .A1(n23624), .A2(n22986), .ZN(n22990) );
  INV_X1 U24803 ( .A(n23620), .ZN(n23569) );
  OAI22_X1 U24804 ( .A1(n23618), .A2(n23622), .B1(n22987), .B2(n23569), .ZN(
        n23184) );
  INV_X1 U24805 ( .A(n23184), .ZN(n22989) );
  INV_X1 U24806 ( .A(n23626), .ZN(n22988) );
  NAND2_X1 U24808 ( .A1(n22991), .A2(n1838), .ZN(n23183) );
  INV_X1 U24809 ( .A(n23183), .ZN(n22994) );
  INV_X1 U24810 ( .A(n23563), .ZN(n23317) );
  NAND2_X1 U24812 ( .A1(n23180), .A2(n29074), .ZN(n22998) );
  NOR2_X1 U24814 ( .A1(n23615), .A2(n23216), .ZN(n23000) );
  INV_X1 U24815 ( .A(n23267), .ZN(n23610) );
  NOR2_X1 U24816 ( .A1(n23610), .A2(n406), .ZN(n22999) );
  MUX2_X1 U24817 ( .A(n23000), .B(n22999), .S(n28581), .Z(n23003) );
  NOR2_X1 U24818 ( .A1(n23001), .A2(n760), .ZN(n23002) );
  NOR2_X2 U24819 ( .A1(n23003), .A2(n23002), .ZN(n24435) );
  AND3_X1 U24820 ( .A1(n29128), .A2(n24437), .A3(n24434), .ZN(n23004) );
  XNOR2_X1 U24821 ( .A(n28645), .B(n25681), .ZN(n24834) );
  NOR2_X1 U24822 ( .A1(n23787), .A2(n23786), .ZN(n23480) );
  OAI21_X1 U24823 ( .B1(n23486), .B2(n23480), .A(n473), .ZN(n24686) );
  INV_X1 U24824 ( .A(n23162), .ZN(n23522) );
  NOR2_X1 U24825 ( .A1(n23006), .A2(n23522), .ZN(n23007) );
  INV_X1 U24826 ( .A(n23662), .ZN(n23667) );
  INV_X1 U24830 ( .A(n23014), .ZN(n23015) );
  INV_X1 U24831 ( .A(n23016), .ZN(n23680) );
  INV_X1 U24832 ( .A(n23134), .ZN(n23019) );
  NOR2_X1 U24833 ( .A1(n23516), .A2(n23680), .ZN(n23018) );
  NAND2_X1 U24834 ( .A1(n24682), .A2(n24688), .ZN(n23020) );
  NAND2_X1 U24835 ( .A1(n23513), .A2(n29641), .ZN(n23022) );
  MUX2_X1 U24836 ( .A(n23022), .B(n23021), .S(n23512), .Z(n24684) );
  NOR2_X1 U24837 ( .A1(n23512), .A2(n339), .ZN(n23023) );
  OAI21_X1 U24838 ( .B1(n23023), .B2(n23488), .A(n6424), .ZN(n24685) );
  NAND2_X1 U24839 ( .A1(n24684), .A2(n24685), .ZN(n24310) );
  NAND2_X1 U24840 ( .A1(n24391), .A2(n24688), .ZN(n23025) );
  AOI21_X1 U24841 ( .B1(n24682), .B2(n23025), .A(n24390), .ZN(n23026) );
  AND2_X1 U24842 ( .A1(n23764), .A2(n23763), .ZN(n23028) );
  NAND2_X1 U24843 ( .A1(n23028), .A2(n23767), .ZN(n23031) );
  NAND2_X1 U24844 ( .A1(n23028), .A2(n23766), .ZN(n23030) );
  NAND3_X1 U24845 ( .A1(n23769), .A2(n23765), .A3(n28554), .ZN(n23029) );
  NOR2_X1 U24846 ( .A1(n23768), .A2(n23765), .ZN(n23151) );
  INV_X1 U24847 ( .A(n23190), .ZN(n23035) );
  INV_X1 U24848 ( .A(n23326), .ZN(n23759) );
  INV_X1 U24849 ( .A(n23474), .ZN(n23033) );
  NOR2_X1 U24850 ( .A1(n23036), .A2(n473), .ZN(n23154) );
  AOI21_X1 U24851 ( .B1(n23785), .B2(n23787), .A(n23484), .ZN(n23038) );
  NAND2_X1 U24852 ( .A1(n23783), .A2(n473), .ZN(n23037) );
  AOI21_X1 U24853 ( .B1(n24706), .B2(n29043), .A(n24707), .ZN(n23051) );
  INV_X1 U24854 ( .A(n23793), .ZN(n23493) );
  NAND2_X1 U24855 ( .A1(n23795), .A2(n23493), .ZN(n23321) );
  INV_X1 U24856 ( .A(n23799), .ZN(n23497) );
  NOR2_X1 U24857 ( .A1(n23799), .A2(n23789), .ZN(n23039) );
  INV_X1 U24858 ( .A(n23555), .ZN(n23045) );
  NAND2_X1 U24859 ( .A1(n23041), .A2(n477), .ZN(n23044) );
  INV_X1 U24860 ( .A(n23630), .ZN(n23559) );
  NAND2_X1 U24861 ( .A1(n23559), .A2(n29061), .ZN(n23042) );
  INV_X1 U24862 ( .A(n23194), .ZN(n23046) );
  AOI21_X1 U24863 ( .B1(n23470), .B2(n23472), .A(n23046), .ZN(n23047) );
  MUX2_X1 U24864 ( .A(n23048), .B(n23047), .S(n23469), .Z(n24339) );
  NOR2_X1 U24865 ( .A1(n23648), .A2(n661), .ZN(n23050) );
  NAND2_X1 U24866 ( .A1(n23193), .A2(n23050), .ZN(n24334) );
  XNOR2_X1 U24867 ( .A(n25910), .B(n28593), .ZN(n24890) );
  XNOR2_X1 U24868 ( .A(n24834), .B(n24890), .ZN(n23125) );
  NAND2_X1 U24869 ( .A1(n29295), .A2(n23445), .ZN(n23052) );
  AOI21_X1 U24870 ( .B1(n23052), .B2(n23442), .A(n292), .ZN(n23056) );
  INV_X1 U24871 ( .A(n23445), .ZN(n23053) );
  NAND3_X1 U24872 ( .A1(n23109), .A2(n23053), .A3(n292), .ZN(n23055) );
  NAND3_X1 U24873 ( .A1(n23370), .A2(n29295), .A3(n23445), .ZN(n23054) );
  INV_X1 U24874 ( .A(n23138), .ZN(n23057) );
  NAND2_X1 U24875 ( .A1(n28570), .A2(n23057), .ZN(n23058) );
  AND2_X1 U24876 ( .A1(n23341), .A2(n23058), .ZN(n23061) );
  NOR2_X1 U24877 ( .A1(n28570), .A2(n28659), .ZN(n23059) );
  NAND2_X1 U24878 ( .A1(n23416), .A2(n485), .ZN(n23062) );
  AOI21_X1 U24879 ( .B1(n24713), .B2(n24716), .A(n4136), .ZN(n23072) );
  MUX2_X1 U24880 ( .A(n23454), .B(n23148), .S(n23456), .Z(n23066) );
  INV_X1 U24881 ( .A(n23456), .ZN(n23147) );
  MUX2_X2 U24882 ( .A(n23066), .B(n23065), .S(n23460), .Z(n24712) );
  INV_X1 U24883 ( .A(n23676), .ZN(n23364) );
  INV_X1 U24884 ( .A(n23672), .ZN(n23366) );
  INV_X1 U24885 ( .A(n23673), .ZN(n23107) );
  NOR2_X1 U24886 ( .A1(n23107), .A2(n23363), .ZN(n23068) );
  NOR2_X1 U24887 ( .A1(n28604), .A2(n23131), .ZN(n23674) );
  AND2_X1 U24888 ( .A1(n24409), .A2(n24711), .ZN(n24351) );
  INV_X1 U24889 ( .A(n24711), .ZN(n24715) );
  XNOR2_X1 U24891 ( .A(n28769), .B(n27737), .ZN(n23123) );
  AND2_X1 U24892 ( .A1(n28653), .A2(n23285), .ZN(n23805) );
  INV_X1 U24893 ( .A(n23810), .ZN(n23807) );
  NAND2_X1 U24894 ( .A1(n22877), .A2(n23806), .ZN(n23286) );
  INV_X1 U24895 ( .A(n24374), .ZN(n24372) );
  NOR2_X1 U24896 ( .A1(n24373), .A2(n24372), .ZN(n23083) );
  OAI211_X1 U24897 ( .C1(n23392), .C2(n23839), .A(n487), .B(n28418), .ZN(
        n23080) );
  OAI21_X1 U24898 ( .B1(n28551), .B2(n23078), .A(n28460), .ZN(n23079) );
  NOR2_X1 U24899 ( .A1(n23995), .A2(n23994), .ZN(n23082) );
  NOR2_X1 U24900 ( .A1(n23301), .A2(n23433), .ZN(n23085) );
  NOR2_X1 U24901 ( .A1(n4178), .A2(n4020), .ZN(n23084) );
  MUX2_X1 U24902 ( .A(n23085), .B(n23084), .S(n201), .Z(n23088) );
  MUX2_X1 U24903 ( .A(n1829), .B(n408), .S(n23433), .Z(n23086) );
  NOR2_X1 U24904 ( .A1(n23086), .A2(n5699), .ZN(n23087) );
  NAND2_X1 U24905 ( .A1(n22931), .A2(n28609), .ZN(n23089) );
  NAND3_X1 U24906 ( .A1(n23441), .A2(n23090), .A3(n23089), .ZN(n23091) );
  OAI211_X1 U24908 ( .C1(n23994), .C2(n23906), .A(n23093), .B(n24372), .ZN(
        n23094) );
  OAI21_X1 U24910 ( .B1(n23415), .B2(n23419), .A(n23101), .ZN(n23968) );
  INV_X1 U24911 ( .A(n23968), .ZN(n23972) );
  NOR2_X1 U24912 ( .A1(n1829), .A2(n29018), .ZN(n23103) );
  NOR2_X1 U24913 ( .A1(n23302), .A2(n23102), .ZN(n23434) );
  OAI21_X1 U24914 ( .B1(n23103), .B2(n23434), .A(n4020), .ZN(n23104) );
  INV_X1 U24915 ( .A(n24209), .ZN(n24046) );
  AOI21_X1 U24916 ( .B1(n23364), .B2(n23366), .A(n23131), .ZN(n23106) );
  NAND2_X1 U24917 ( .A1(n29296), .A2(n23109), .ZN(n23110) );
  NOR2_X1 U24918 ( .A1(n469), .A2(n24479), .ZN(n23970) );
  INV_X1 U24919 ( .A(n23422), .ZN(n23428) );
  INV_X1 U24920 ( .A(n23338), .ZN(n23426) );
  MUX2_X1 U24921 ( .A(n23138), .B(n23427), .S(n28659), .Z(n23114) );
  INV_X1 U24922 ( .A(n23343), .ZN(n23339) );
  NOR2_X1 U24924 ( .A1(n23339), .A2(n28122), .ZN(n23113) );
  INV_X1 U24925 ( .A(n29108), .ZN(n23112) );
  AOI22_X1 U24926 ( .A1(n23344), .A2(n23114), .B1(n23113), .B2(n23112), .ZN(
        n23115) );
  OAI21_X1 U24927 ( .B1(n23116), .B2(n23970), .A(n24483), .ZN(n23121) );
  NOR2_X1 U24929 ( .A1(n23456), .A2(n29042), .ZN(n23117) );
  INV_X1 U24930 ( .A(n23460), .ZN(n23458) );
  AND2_X1 U24931 ( .A1(n23455), .A2(n23460), .ZN(n23355) );
  NAND2_X1 U24932 ( .A1(n24484), .A2(n24209), .ZN(n23119) );
  XNOR2_X1 U24933 ( .A(n28628), .B(n25845), .ZN(n23122) );
  XNOR2_X1 U24934 ( .A(n23122), .B(n23123), .ZN(n23124) );
  INV_X1 U24935 ( .A(n26789), .ZN(n26575) );
  NAND2_X1 U24936 ( .A1(n24542), .A2(n2823), .ZN(n24540) );
  OAI21_X1 U24937 ( .B1(n24540), .B2(n24160), .A(n23128), .ZN(n23130) );
  INV_X1 U24939 ( .A(n23683), .ZN(n23517) );
  NOR2_X1 U24940 ( .A1(n4232), .A2(n4231), .ZN(n23142) );
  INV_X1 U24941 ( .A(n24891), .ZN(n23144) );
  NAND2_X1 U24942 ( .A1(n24631), .A2(n24629), .ZN(n24530) );
  OAI21_X1 U24943 ( .B1(n1837), .B2(n23461), .A(n23458), .ZN(n23146) );
  NAND2_X1 U24944 ( .A1(n29042), .A2(n23456), .ZN(n23457) );
  INV_X1 U24945 ( .A(n23767), .ZN(n23329) );
  OAI21_X1 U24946 ( .B1(n23764), .B2(n23763), .A(n23769), .ZN(n23152) );
  NAND2_X1 U24947 ( .A1(n23768), .A2(n23152), .ZN(n23153) );
  INV_X1 U24948 ( .A(n24642), .ZN(n24568) );
  NAND3_X1 U24949 ( .A1(n23785), .A2(n475), .A3(n23788), .ZN(n23155) );
  NAND2_X1 U24950 ( .A1(n24568), .A2(n24237), .ZN(n24641) );
  NAND2_X1 U24951 ( .A1(n23156), .A2(n23771), .ZN(n23157) );
  INV_X1 U24952 ( .A(n23157), .ZN(n23489) );
  OAI21_X1 U24953 ( .B1(n23779), .B2(n23776), .A(n23772), .ZN(n23161) );
  NOR2_X1 U24954 ( .A1(n23514), .A2(n23776), .ZN(n23159) );
  AND2_X1 U24955 ( .A1(n23666), .A2(n23162), .ZN(n23527) );
  OAI21_X1 U24956 ( .B1(n29123), .B2(n23163), .A(n23527), .ZN(n23166) );
  NAND2_X1 U24957 ( .A1(n23164), .A2(n23663), .ZN(n23165) );
  OAI211_X1 U24958 ( .C1(n23662), .C2(n23663), .A(n23166), .B(n23165), .ZN(
        n24638) );
  NAND2_X1 U24959 ( .A1(n23169), .A2(n23016), .ZN(n23171) );
  AOI21_X1 U24962 ( .B1(n23801), .B2(n23800), .A(n1913), .ZN(n23174) );
  NOR2_X1 U24963 ( .A1(n23537), .A2(n28444), .ZN(n23172) );
  NOR3_X1 U24965 ( .A1(n29074), .A2(n23177), .A3(n23563), .ZN(n23179) );
  NAND2_X1 U24966 ( .A1(n23621), .A2(n23619), .ZN(n23568) );
  NAND2_X1 U24967 ( .A1(n23568), .A2(n23620), .ZN(n23185) );
  NAND2_X1 U24968 ( .A1(n23185), .A2(n726), .ZN(n23186) );
  NOR2_X1 U24969 ( .A1(n24241), .A2(n24240), .ZN(n23990) );
  NOR2_X1 U24970 ( .A1(n5775), .A2(n23629), .ZN(n23187) );
  NOR2_X1 U24971 ( .A1(n23309), .A2(n28644), .ZN(n23188) );
  MUX2_X1 U24973 ( .A(n23193), .B(n23649), .S(n23651), .Z(n23195) );
  NAND2_X1 U24974 ( .A1(n23196), .A2(n23492), .ZN(n23197) );
  NAND2_X1 U24975 ( .A1(n23197), .A2(n23792), .ZN(n23200) );
  NAND2_X1 U24979 ( .A1(n24239), .A2(n25794), .ZN(n23201) );
  XNOR2_X1 U24980 ( .A(n25775), .B(n26004), .ZN(n25216) );
  XNOR2_X1 U24981 ( .A(n25216), .B(n25563), .ZN(n23244) );
  AOI21_X1 U24982 ( .B1(n23202), .B2(n1883), .A(n24377), .ZN(n23204) );
  NOR3_X1 U24983 ( .A1(n24373), .A2(n24374), .A3(n1883), .ZN(n23203) );
  NAND2_X1 U24984 ( .A1(n23936), .A2(n24553), .ZN(n23206) );
  XNOR2_X1 U24985 ( .A(n29534), .B(n25565), .ZN(n23242) );
  NOR2_X1 U24986 ( .A1(n23607), .A2(n23247), .ZN(n23209) );
  NAND2_X1 U24988 ( .A1(n23602), .A2(n23246), .ZN(n23210) );
  OAI21_X1 U24989 ( .B1(n23606), .B2(n23578), .A(n23210), .ZN(n23608) );
  INV_X1 U24990 ( .A(n23406), .ZN(n23214) );
  OAI21_X1 U24991 ( .B1(n23403), .B2(n23250), .A(n23252), .ZN(n23215) );
  AOI22_X1 U24992 ( .A1(n23615), .A2(n23216), .B1(n28225), .B2(n28544), .ZN(
        n23219) );
  NAND2_X1 U24996 ( .A1(n1862), .A2(n23398), .ZN(n23230) );
  INV_X1 U24997 ( .A(n23736), .ZN(n23228) );
  NAND2_X1 U24999 ( .A1(n24524), .A2(n28481), .ZN(n23238) );
  NAND2_X1 U25000 ( .A1(n380), .A2(n23714), .ZN(n23713) );
  NAND2_X1 U25004 ( .A1(n23238), .A2(n24245), .ZN(n23239) );
  NOR2_X2 U25005 ( .A1(n23240), .A2(n23239), .ZN(n25346) );
  XNOR2_X1 U25006 ( .A(n25346), .B(n1079), .ZN(n23241) );
  XNOR2_X1 U25007 ( .A(n23242), .B(n23241), .ZN(n23243) );
  MUX2_X1 U25008 ( .A(n23602), .B(n23246), .S(n23245), .Z(n23248) );
  AND2_X1 U25009 ( .A1(n23406), .A2(n22979), .ZN(n23254) );
  NOR2_X1 U25010 ( .A1(n23213), .A2(n22979), .ZN(n23253) );
  INV_X1 U25011 ( .A(n23258), .ZN(n23256) );
  NAND2_X1 U25012 ( .A1(n23732), .A2(n23257), .ZN(n23259) );
  NOR2_X1 U25014 ( .A1(n28528), .A2(n28415), .ZN(n23269) );
  AOI21_X1 U25015 ( .B1(n23267), .B2(n28582), .A(n29115), .ZN(n23268) );
  NOR2_X1 U25016 ( .A1(n24368), .A2(n24369), .ZN(n24064) );
  OAI21_X1 U25019 ( .B1(n29564), .B2(n23382), .A(n23825), .ZN(n23276) );
  AOI21_X1 U25020 ( .B1(n23385), .B2(n23382), .A(n23276), .ZN(n23279) );
  NAND3_X1 U25021 ( .A1(n28181), .A2(n23382), .A3(n2187), .ZN(n23277) );
  OAI21_X1 U25022 ( .B1(n23738), .B2(n28181), .A(n23277), .ZN(n23278) );
  INV_X1 U25024 ( .A(n24083), .ZN(n24084) );
  INV_X1 U25025 ( .A(n23281), .ZN(n23282) );
  INV_X1 U25026 ( .A(n23285), .ZN(n23287) );
  MUX2_X1 U25027 ( .A(n24084), .B(n6265), .S(n24403), .Z(n23307) );
  INV_X1 U25028 ( .A(n23291), .ZN(n23816) );
  NOR3_X1 U25029 ( .A1(n4950), .A2(n28182), .A3(n23290), .ZN(n23292) );
  OAI22_X1 U25030 ( .A1(n23292), .A2(n23821), .B1(n23819), .B2(n5591), .ZN(
        n23293) );
  INV_X1 U25031 ( .A(n23294), .ZN(n23300) );
  OAI21_X1 U25032 ( .B1(n22531), .B2(n23295), .A(n29602), .ZN(n23299) );
  OAI21_X1 U25033 ( .B1(n23301), .B2(n29018), .A(n5530), .ZN(n23304) );
  XNOR2_X1 U25034 ( .A(n26011), .B(n25884), .ZN(n23337) );
  NOR2_X1 U25035 ( .A1(n23637), .A2(n23630), .ZN(n23308) );
  OAI21_X1 U25036 ( .B1(n23309), .B2(n5775), .A(n477), .ZN(n23311) );
  NAND2_X1 U25038 ( .A1(n22992), .A2(n23640), .ZN(n23313) );
  OAI21_X1 U25039 ( .B1(n22996), .B2(n23314), .A(n1838), .ZN(n23316) );
  NOR2_X1 U25041 ( .A1(n24395), .A2(n28635), .ZN(n24068) );
  NOR2_X1 U25042 ( .A1(n23320), .A2(n23792), .ZN(n23322) );
  NOR2_X1 U25043 ( .A1(n24678), .A2(n24672), .ZN(n23324) );
  NOR2_X1 U25044 ( .A1(n24068), .A2(n23324), .ZN(n23334) );
  INV_X1 U25045 ( .A(n28635), .ZN(n24676) );
  MUX2_X1 U25046 ( .A(n23758), .B(n23326), .S(n29131), .Z(n23327) );
  NAND2_X1 U25048 ( .A1(n4759), .A2(n23769), .ZN(n23332) );
  NAND2_X1 U25049 ( .A1(n23764), .A2(n28554), .ZN(n23330) );
  MUX2_X1 U25050 ( .A(n23330), .B(n23501), .S(n23767), .Z(n23331) );
  AND2_X1 U25052 ( .A1(n29471), .A2(n24688), .ZN(n23335) );
  AOI22_X1 U25053 ( .A1(n466), .A2(n23335), .B1(n24682), .B2(n24391), .ZN(
        n23336) );
  XNOR2_X1 U25054 ( .A(n25761), .B(n25444), .ZN(n25234) );
  XNOR2_X1 U25055 ( .A(n25234), .B(n23337), .ZN(n23414) );
  NAND2_X1 U25056 ( .A1(n23339), .A2(n23338), .ZN(n23342) );
  NOR3_X1 U25057 ( .A1(n23344), .A2(n29108), .A3(n28570), .ZN(n23345) );
  MUX2_X1 U25059 ( .A(n23535), .B(n5030), .S(n28164), .Z(n23350) );
  NAND2_X1 U25060 ( .A1(n23696), .A2(n23529), .ZN(n23347) );
  MUX2_X1 U25061 ( .A(n23348), .B(n23347), .S(n23535), .Z(n23349) );
  INV_X1 U25062 ( .A(n24665), .ZN(n24382) );
  AOI21_X1 U25063 ( .B1(n23657), .B2(n23351), .A(n29583), .ZN(n23352) );
  NAND2_X1 U25064 ( .A1(n4605), .A2(n4195), .ZN(n23375) );
  NAND2_X1 U25065 ( .A1(n23355), .A2(n29042), .ZN(n23359) );
  INV_X1 U25066 ( .A(n23356), .ZN(n23358) );
  NOR2_X1 U25067 ( .A1(n24665), .A2(n24666), .ZN(n23373) );
  MUX2_X1 U25069 ( .A(n23362), .B(n23361), .S(n23360), .Z(n23369) );
  AOI21_X1 U25070 ( .B1(n23367), .B2(n23366), .A(n23365), .ZN(n23368) );
  NOR2_X1 U25071 ( .A1(n24382), .A2(n24668), .ZN(n24073) );
  INV_X1 U25072 ( .A(n23370), .ZN(n23371) );
  NAND2_X1 U25073 ( .A1(n24316), .A2(n24383), .ZN(n23372) );
  AOI21_X1 U25075 ( .B1(n24374), .B2(n1828), .A(n24373), .ZN(n23376) );
  NAND2_X1 U25076 ( .A1(n23906), .A2(n24376), .ZN(n23380) );
  NAND2_X1 U25077 ( .A1(n1828), .A2(n24380), .ZN(n23378) );
  XNOR2_X1 U25078 ( .A(n25933), .B(n25931), .ZN(n23412) );
  NAND2_X1 U25079 ( .A1(n23738), .A2(n23827), .ZN(n23384) );
  OAI21_X1 U25080 ( .B1(n22451), .B2(n29618), .A(n23702), .ZN(n23388) );
  OAI21_X1 U25081 ( .B1(n23722), .B2(n28484), .A(n23726), .ZN(n23395) );
  NOR2_X1 U25082 ( .A1(n28484), .A2(n23720), .ZN(n23394) );
  INV_X1 U25083 ( .A(n24388), .ZN(n23911) );
  OAI211_X1 U25084 ( .C1(n23228), .C2(n23399), .A(n23398), .B(n23397), .ZN(
        n23400) );
  NOR2_X1 U25085 ( .A1(n23403), .A2(n28527), .ZN(n23404) );
  NAND3_X1 U25086 ( .A1(n24133), .A2(n24388), .A3(n24078), .ZN(n23409) );
  XNOR2_X1 U25087 ( .A(n25179), .B(n622), .ZN(n23411) );
  XNOR2_X1 U25088 ( .A(n23412), .B(n23411), .ZN(n23413) );
  NAND2_X1 U25090 ( .A1(n23422), .A2(n28659), .ZN(n23423) );
  NAND2_X1 U25091 ( .A1(n23424), .A2(n23423), .ZN(n23429) );
  NOR2_X1 U25092 ( .A1(n1829), .A2(n408), .ZN(n23437) );
  NAND2_X1 U25093 ( .A1(n4020), .A2(n23431), .ZN(n23436) );
  OAI21_X1 U25094 ( .B1(n23433), .B2(n29018), .A(n23431), .ZN(n23435) );
  NAND2_X1 U25095 ( .A1(n4950), .A2(n28182), .ZN(n23440) );
  NAND3_X1 U25096 ( .A1(n2281), .A2(n4950), .A3(n22931), .ZN(n23438) );
  NOR2_X1 U25097 ( .A1(n23445), .A2(n23442), .ZN(n23443) );
  NAND3_X1 U25098 ( .A1(n23447), .A2(n23446), .A3(n23445), .ZN(n23452) );
  NAND3_X1 U25099 ( .A1(n29296), .A2(n23449), .A3(n292), .ZN(n23451) );
  MUX2_X1 U25100 ( .A(n23456), .B(n23455), .S(n23454), .Z(n23466) );
  INV_X1 U25101 ( .A(n23457), .ZN(n23459) );
  AND2_X1 U25102 ( .A1(n23460), .A2(n23461), .ZN(n23462) );
  NAND2_X1 U25103 ( .A1(n23462), .A2(n23465), .ZN(n23463) );
  OR2_X1 U25105 ( .A1(n24012), .A2(n23597), .ZN(n23468) );
  INV_X1 U25106 ( .A(n23475), .ZN(n23479) );
  OAI21_X1 U25107 ( .B1(n23758), .B2(n23759), .A(n23761), .ZN(n23478) );
  MUX2_X1 U25108 ( .A(n23476), .B(n23475), .S(n23474), .Z(n23477) );
  NOR2_X1 U25109 ( .A1(n24775), .A2(n470), .ZN(n23502) );
  INV_X1 U25110 ( .A(n23480), .ZN(n23481) );
  NOR2_X1 U25111 ( .A1(n23481), .A2(n23788), .ZN(n23485) );
  NAND2_X1 U25112 ( .A1(n23482), .A2(n23784), .ZN(n23483) );
  INV_X1 U25113 ( .A(n24777), .ZN(n24780) );
  OAI22_X1 U25114 ( .A1(n23157), .A2(n23778), .B1(n23514), .B2(n29641), .ZN(
        n23490) );
  NAND3_X1 U25115 ( .A1(n23493), .A2(n23789), .A3(n23492), .ZN(n23494) );
  OAI21_X1 U25116 ( .B1(n23495), .B2(n23795), .A(n23494), .ZN(n23496) );
  AOI21_X2 U25117 ( .B1(n23498), .B2(n23497), .A(n23496), .ZN(n24776) );
  NOR2_X1 U25118 ( .A1(n23946), .A2(n24776), .ZN(n24454) );
  OAI21_X1 U25119 ( .B1(n23499), .B2(n23765), .A(n23764), .ZN(n23500) );
  XNOR2_X1 U25120 ( .A(n25282), .B(n26029), .ZN(n23511) );
  NAND2_X1 U25121 ( .A1(n24083), .A2(n24408), .ZN(n23504) );
  MUX2_X1 U25122 ( .A(n23504), .B(n23503), .S(n24404), .Z(n23505) );
  MUX2_X1 U25123 ( .A(n24077), .B(n24388), .S(n24387), .Z(n23510) );
  XNOR2_X1 U25125 ( .A(n25324), .B(n25751), .ZN(n24307) );
  XNOR2_X1 U25126 ( .A(n23511), .B(n24307), .ZN(n23596) );
  MUX2_X2 U25128 ( .A(n23521), .B(n23520), .S(n23016), .Z(n24772) );
  MUX2_X1 U25130 ( .A(n23524), .B(n23523), .S(n23663), .Z(n23528) );
  NOR2_X1 U25131 ( .A1(n23666), .A2(n23525), .ZN(n23526) );
  MUX2_X1 U25132 ( .A(n24697), .B(n24772), .S(n24765), .Z(n23550) );
  NAND2_X1 U25133 ( .A1(n23531), .A2(n23697), .ZN(n23534) );
  INV_X1 U25135 ( .A(n23689), .ZN(n23539) );
  INV_X1 U25136 ( .A(n23540), .ZN(n23542) );
  NOR2_X1 U25138 ( .A1(n24769), .A2(n29624), .ZN(n23547) );
  AOI21_X2 U25139 ( .B1(n23550), .B2(n28598), .A(n23549), .ZN(n25037) );
  INV_X1 U25142 ( .A(n24484), .ZN(n24213) );
  NAND3_X1 U25143 ( .A1(n24213), .A2(n29597), .A3(n24209), .ZN(n23552) );
  NAND3_X1 U25144 ( .A1(n24480), .A2(n24210), .A3(n24483), .ZN(n23551) );
  OAI211_X2 U25145 ( .C1(n24482), .C2(n23553), .A(n23552), .B(n23551), .ZN(
        n25209) );
  XNOR2_X1 U25146 ( .A(n25037), .B(n25209), .ZN(n25939) );
  NAND2_X1 U25147 ( .A1(n23559), .A2(n23558), .ZN(n23560) );
  NOR3_X1 U25148 ( .A1(n29115), .A2(n379), .A3(n28225), .ZN(n23955) );
  INV_X1 U25149 ( .A(n23955), .ZN(n24218) );
  NAND2_X1 U25150 ( .A1(n24447), .A2(n24218), .ZN(n23576) );
  NAND2_X1 U25151 ( .A1(n23641), .A2(n23563), .ZN(n23646) );
  NOR2_X1 U25152 ( .A1(n23618), .A2(n23621), .ZN(n23574) );
  OAI21_X1 U25153 ( .B1(n23567), .B2(n23566), .A(n23622), .ZN(n23573) );
  INV_X1 U25154 ( .A(n23568), .ZN(n23571) );
  NOR2_X1 U25155 ( .A1(n23621), .A2(n23569), .ZN(n23570) );
  INV_X1 U25156 ( .A(n24760), .ZN(n23588) );
  AOI21_X1 U25157 ( .B1(n29592), .B2(n24761), .A(n23588), .ZN(n23575) );
  MUX2_X1 U25158 ( .A(n5347), .B(n23578), .S(n23577), .Z(n23582) );
  NAND2_X1 U25159 ( .A1(n23583), .A2(n23603), .ZN(n23580) );
  NAND2_X1 U25160 ( .A1(n23607), .A2(n23578), .ZN(n23579) );
  MUX2_X1 U25161 ( .A(n23580), .B(n23579), .S(n5347), .Z(n23581) );
  INV_X1 U25162 ( .A(n24757), .ZN(n24220) );
  OAI21_X1 U25163 ( .B1(n24220), .B2(n24756), .A(n23588), .ZN(n23591) );
  INV_X1 U25164 ( .A(n23956), .ZN(n23589) );
  AOI21_X1 U25165 ( .B1(n23589), .B2(n24218), .A(n28509), .ZN(n23590) );
  INV_X1 U25167 ( .A(n2544), .ZN(n23593) );
  XNOR2_X1 U25168 ( .A(n25785), .B(n23593), .ZN(n23594) );
  XNOR2_X1 U25169 ( .A(n25939), .B(n23594), .ZN(n23595) );
  XNOR2_X1 U25170 ( .A(n23595), .B(n23596), .ZN(n26791) );
  NOR2_X1 U25172 ( .A1(n24972), .A2(n24256), .ZN(n23598) );
  OAI21_X1 U25173 ( .B1(n23604), .B2(n23603), .A(n23602), .ZN(n23605) );
  NAND3_X1 U25175 ( .A1(n4599), .A2(n23610), .A3(n28581), .ZN(n23617) );
  MUX2_X1 U25176 ( .A(n23611), .B(n23615), .S(n379), .Z(n23613) );
  NOR2_X1 U25177 ( .A1(n24790), .A2(n24791), .ZN(n24507) );
  AOI21_X1 U25178 ( .B1(n23622), .B2(n23619), .A(n23618), .ZN(n23625) );
  NOR2_X1 U25179 ( .A1(n23621), .A2(n23620), .ZN(n23623) );
  INV_X1 U25180 ( .A(n24790), .ZN(n24792) );
  AOI21_X1 U25181 ( .B1(n23630), .B2(n23629), .A(n23628), .ZN(n23635) );
  NOR2_X1 U25182 ( .A1(n23632), .A2(n28644), .ZN(n23634) );
  MUX2_X1 U25183 ( .A(n23635), .B(n23634), .S(n29061), .Z(n23639) );
  NOR2_X1 U25184 ( .A1(n23637), .A2(n23636), .ZN(n23638) );
  OR2_X2 U25185 ( .A1(n23639), .A2(n23638), .ZN(n24269) );
  NOR2_X1 U25186 ( .A1(n23641), .A2(n23640), .ZN(n23644) );
  NAND2_X1 U25187 ( .A1(n23648), .A2(n23647), .ZN(n23650) );
  XNOR2_X1 U25188 ( .A(n25944), .B(n25826), .ZN(n23756) );
  NOR2_X1 U25189 ( .A1(n23656), .A2(n23657), .ZN(n23660) );
  NOR2_X1 U25190 ( .A1(n23662), .A2(n28577), .ZN(n23664) );
  NOR2_X1 U25191 ( .A1(n23666), .A2(n23665), .ZN(n23668) );
  NOR3_X1 U25192 ( .A1(n23669), .A2(n23668), .A3(n23667), .ZN(n23670) );
  NOR2_X1 U25194 ( .A1(n23673), .A2(n23672), .ZN(n23675) );
  AOI21_X1 U25195 ( .B1(n28604), .B2(n23675), .A(n23674), .ZN(n23677) );
  INV_X1 U25196 ( .A(n23681), .ZN(n23685) );
  NOR2_X1 U25197 ( .A1(n23016), .A2(n23682), .ZN(n23684) );
  NOR2_X1 U25198 ( .A1(n24808), .A2(n24817), .ZN(n23691) );
  OAI21_X1 U25199 ( .B1(n23801), .B2(n23687), .A(n23800), .ZN(n23688) );
  MUX2_X1 U25200 ( .A(n23692), .B(n23691), .S(n5004), .Z(n23699) );
  INV_X1 U25201 ( .A(n24817), .ZN(n24461) );
  NAND2_X1 U25202 ( .A1(n484), .A2(n23067), .ZN(n23695) );
  NOR2_X2 U25203 ( .A1(n23699), .A2(n23698), .ZN(n25943) );
  NOR2_X1 U25204 ( .A1(n22084), .A2(n23700), .ZN(n23703) );
  MUX2_X1 U25205 ( .A(n23704), .B(n23703), .S(n23387), .Z(n23709) );
  NOR2_X2 U25206 ( .A1(n23709), .A2(n23708), .ZN(n24111) );
  INV_X1 U25207 ( .A(n24111), .ZN(n24179) );
  NAND2_X1 U25208 ( .A1(n23714), .A2(n23710), .ZN(n23711) );
  MUX2_X1 U25209 ( .A(n23712), .B(n23711), .S(n23715), .Z(n23719) );
  OAI21_X1 U25210 ( .B1(n23715), .B2(n23714), .A(n23713), .ZN(n23717) );
  NAND2_X1 U25211 ( .A1(n23717), .A2(n23716), .ZN(n23718) );
  INV_X1 U25212 ( .A(n24517), .ZN(n24113) );
  MUX2_X1 U25213 ( .A(n23722), .B(n23721), .S(n23720), .Z(n23723) );
  NOR2_X1 U25214 ( .A1(n23724), .A2(n23843), .ZN(n23729) );
  NOR2_X1 U25215 ( .A1(n23849), .A2(n28484), .ZN(n23727) );
  INV_X1 U25217 ( .A(n23745), .ZN(n24515) );
  NOR2_X1 U25218 ( .A1(n24520), .A2(n24515), .ZN(n23744) );
  INV_X1 U25219 ( .A(n23738), .ZN(n23739) );
  OAI21_X1 U25220 ( .B1(n28181), .B2(n23827), .A(n23739), .ZN(n23740) );
  OAI21_X2 U25221 ( .B1(n23743), .B2(n23382), .A(n23742), .ZN(n24514) );
  NAND2_X1 U25222 ( .A1(n24515), .A2(n24514), .ZN(n24424) );
  NOR2_X1 U25223 ( .A1(n24516), .A2(n24111), .ZN(n23752) );
  INV_X1 U25224 ( .A(n23746), .ZN(n23751) );
  XNOR2_X1 U25226 ( .A(n25943), .B(n26056), .ZN(n23755) );
  XNOR2_X1 U25227 ( .A(n23756), .B(n23755), .ZN(n23861) );
  NAND2_X1 U25228 ( .A1(n23764), .A2(n23765), .ZN(n23770) );
  NOR2_X1 U25229 ( .A1(n339), .A2(n23771), .ZN(n23775) );
  NOR2_X1 U25230 ( .A1(n29641), .A2(n23772), .ZN(n23774) );
  MUX2_X1 U25231 ( .A(n23775), .B(n23774), .S(n23776), .Z(n23782) );
  AOI21_X1 U25232 ( .B1(n23780), .B2(n23779), .A(n23778), .ZN(n23781) );
  MUX2_X1 U25234 ( .A(n24162), .B(n24503), .S(n24801), .Z(n23804) );
  MUX2_X1 U25236 ( .A(n23790), .B(n23789), .S(n23791), .Z(n23798) );
  NAND3_X1 U25237 ( .A1(n6608), .A2(n23792), .A3(n23791), .ZN(n23794) );
  OAI21_X1 U25238 ( .B1(n23796), .B2(n23795), .A(n23794), .ZN(n23797) );
  NOR2_X1 U25239 ( .A1(n22742), .A2(n23808), .ZN(n23812) );
  OAI21_X1 U25240 ( .B1(n23812), .B2(n23811), .A(n23810), .ZN(n23813) );
  NOR2_X1 U25241 ( .A1(n23819), .A2(n23816), .ZN(n23817) );
  AND2_X1 U25244 ( .A1(n23842), .A2(n24472), .ZN(n24475) );
  OAI211_X1 U25245 ( .C1(n23829), .C2(n482), .A(n28181), .B(n23827), .ZN(
        n24091) );
  NOR2_X1 U25246 ( .A1(n23832), .A2(n29602), .ZN(n23834) );
  NOR2_X1 U25247 ( .A1(n24471), .A2(n29051), .ZN(n23841) );
  NAND3_X1 U25248 ( .A1(n6279), .A2(n28460), .A3(n23839), .ZN(n23840) );
  INV_X1 U25249 ( .A(n23842), .ZN(n24100) );
  XNOR2_X1 U25250 ( .A(n24949), .B(n26054), .ZN(n23859) );
  NOR2_X1 U25251 ( .A1(n23853), .A2(n24141), .ZN(n23857) );
  INV_X1 U25252 ( .A(n24591), .ZN(n24143) );
  NOR2_X1 U25253 ( .A1(n24143), .A2(n24592), .ZN(n23854) );
  XNOR2_X1 U25254 ( .A(n25858), .B(n3081), .ZN(n23858) );
  XNOR2_X1 U25255 ( .A(n23858), .B(n23859), .ZN(n23860) );
  INV_X1 U25256 ( .A(n26793), .ZN(n26572) );
  NOR2_X1 U25257 ( .A1(n23863), .A2(n6826), .ZN(n23864) );
  INV_X1 U25258 ( .A(n307), .ZN(n24364) );
  INV_X1 U25259 ( .A(n24767), .ZN(n24426) );
  MUX2_X1 U25260 ( .A(n1856), .B(n24426), .S(n24765), .Z(n23866) );
  MUX2_X1 U25261 ( .A(n24765), .B(n24427), .S(n24772), .Z(n23865) );
  MUX2_X1 U25262 ( .A(n24711), .B(n24716), .S(n24712), .Z(n23868) );
  INV_X1 U25263 ( .A(n24409), .ZN(n24720) );
  INV_X1 U25265 ( .A(n24514), .ZN(n24421) );
  NOR2_X1 U25266 ( .A1(n24111), .A2(n24420), .ZN(n24518) );
  INV_X1 U25267 ( .A(n24518), .ZN(n23871) );
  XNOR2_X1 U25270 ( .A(n26073), .B(n26040), .ZN(n25687) );
  XNOR2_X1 U25271 ( .A(n25687), .B(n25260), .ZN(n23893) );
  INV_X1 U25272 ( .A(n23874), .ZN(n24474) );
  NAND2_X1 U25273 ( .A1(n24474), .A2(n24471), .ZN(n24490) );
  INV_X1 U25274 ( .A(n24490), .ZN(n23879) );
  INV_X1 U25275 ( .A(n24472), .ZN(n24491) );
  NAND2_X1 U25276 ( .A1(n24491), .A2(n24100), .ZN(n23876) );
  MUX2_X1 U25277 ( .A(n24408), .B(n24085), .S(n24405), .Z(n23883) );
  NAND2_X1 U25278 ( .A1(n24403), .A2(n24084), .ZN(n23881) );
  MUX2_X1 U25279 ( .A(n23881), .B(n23880), .S(n24405), .Z(n23882) );
  OAI21_X2 U25280 ( .B1(n23883), .B2(n24403), .A(n23882), .ZN(n26045) );
  XNOR2_X1 U25281 ( .A(n1922), .B(n26045), .ZN(n23891) );
  NAND2_X1 U25282 ( .A1(n24347), .A2(n29726), .ZN(n23884) );
  XNOR2_X1 U25284 ( .A(n28540), .B(n624), .ZN(n23890) );
  XNOR2_X1 U25285 ( .A(n23891), .B(n23890), .ZN(n23892) );
  INV_X1 U25286 ( .A(n26179), .ZN(n26456) );
  NAND2_X1 U25287 ( .A1(n24323), .A2(n28635), .ZN(n23896) );
  NAND2_X1 U25288 ( .A1(n24678), .A2(n24672), .ZN(n24396) );
  NAND2_X1 U25289 ( .A1(n24396), .A2(n6944), .ZN(n23894) );
  NAND2_X1 U25290 ( .A1(n24068), .A2(n24677), .ZN(n23895) );
  AND3_X1 U25291 ( .A1(n24369), .A2(n24304), .A3(n25005), .ZN(n23898) );
  XNOR2_X1 U25292 ( .A(n25532), .B(n25855), .ZN(n25150) );
  INV_X1 U25293 ( .A(n24691), .ZN(n23899) );
  NOR2_X1 U25295 ( .A1(n24682), .A2(n24391), .ZN(n23902) );
  NOR2_X1 U25296 ( .A1(n466), .A2(n29567), .ZN(n23901) );
  NOR2_X1 U25297 ( .A1(n23905), .A2(n24372), .ZN(n23907) );
  XNOR2_X1 U25298 ( .A(n25246), .B(n26055), .ZN(n23908) );
  XNOR2_X1 U25299 ( .A(n25150), .B(n23908), .ZN(n23920) );
  XNOR2_X1 U25300 ( .A(n25375), .B(n27978), .ZN(n23918) );
  INV_X1 U25301 ( .A(n24387), .ZN(n24079) );
  NOR2_X1 U25302 ( .A1(n28424), .A2(n24072), .ZN(n23917) );
  NAND2_X1 U25303 ( .A1(n23914), .A2(n4195), .ZN(n23916) );
  NAND2_X1 U25304 ( .A1(n24668), .A2(n24383), .ZN(n23913) );
  XNOR2_X1 U25306 ( .A(n26060), .B(n25372), .ZN(n25698) );
  XNOR2_X1 U25307 ( .A(n23918), .B(n25698), .ZN(n23919) );
  NAND2_X1 U25308 ( .A1(n26456), .A2(n26449), .ZN(n25622) );
  INV_X1 U25309 ( .A(n24610), .ZN(n23953) );
  OAI21_X1 U25310 ( .B1(n23953), .B2(n24057), .A(n24614), .ZN(n23923) );
  XNOR2_X1 U25311 ( .A(n25848), .B(n29543), .ZN(n25310) );
  NOR2_X1 U25313 ( .A1(n24617), .A2(n24747), .ZN(n24022) );
  NOR2_X1 U25314 ( .A1(n21303), .A2(n24617), .ZN(n23926) );
  AOI22_X1 U25315 ( .A1(n28223), .A2(n24022), .B1(n23926), .B2(n24751), .ZN(
        n23927) );
  OAI21_X1 U25316 ( .B1(n24593), .B2(n24277), .A(n24590), .ZN(n23930) );
  XNOR2_X1 U25317 ( .A(n25328), .B(n25249), .ZN(n26021) );
  XNOR2_X1 U25318 ( .A(n26021), .B(n25310), .ZN(n23941) );
  OAI21_X1 U25319 ( .B1(n24596), .B2(n24597), .A(n24595), .ZN(n23934) );
  XNOR2_X1 U25320 ( .A(n25808), .B(n2477), .ZN(n23939) );
  INV_X1 U25321 ( .A(n24734), .ZN(n24601) );
  OAI21_X1 U25322 ( .B1(n24601), .B2(n24736), .A(n24602), .ZN(n23935) );
  OAI21_X1 U25324 ( .B1(n24555), .B2(n24551), .A(n28519), .ZN(n23937) );
  XNOR2_X1 U25325 ( .A(n25133), .B(n25396), .ZN(n23938) );
  XNOR2_X1 U25326 ( .A(n23939), .B(n23938), .ZN(n23940) );
  INV_X1 U25327 ( .A(n24471), .ZN(n23942) );
  NOR2_X1 U25329 ( .A1(n23945), .A2(n29308), .ZN(n24040) );
  INV_X1 U25330 ( .A(n24040), .ZN(n24456) );
  OAI21_X1 U25331 ( .B1(n23946), .B2(n24777), .A(n29308), .ZN(n23947) );
  NAND2_X1 U25332 ( .A1(n24456), .A2(n23947), .ZN(n23949) );
  OAI211_X1 U25333 ( .C1(n24779), .C2(n24775), .A(n24777), .B(n24776), .ZN(
        n23948) );
  XNOR2_X1 U25334 ( .A(n25708), .B(n25922), .ZN(n23952) );
  AOI21_X1 U25335 ( .B1(n5004), .B2(n24808), .A(n24499), .ZN(n23950) );
  XNOR2_X1 U25337 ( .A(n23952), .B(n29111), .ZN(n25258) );
  OAI211_X1 U25338 ( .C1(n5168), .C2(n24017), .A(n24057), .B(n23953), .ZN(
        n23954) );
  AOI21_X1 U25339 ( .B1(n24220), .B2(n28509), .A(n378), .ZN(n23959) );
  AND2_X1 U25340 ( .A1(n24760), .A2(n24756), .ZN(n24450) );
  INV_X1 U25341 ( .A(n24450), .ZN(n23957) );
  XNOR2_X1 U25342 ( .A(n25868), .B(n27515), .ZN(n23960) );
  XNOR2_X1 U25343 ( .A(n23960), .B(n25773), .ZN(n23961) );
  INV_X1 U25344 ( .A(n23962), .ZN(n24467) );
  INV_X1 U25347 ( .A(n24055), .ZN(n23966) );
  MUX2_X1 U25349 ( .A(n24484), .B(n469), .S(n23968), .Z(n24050) );
  NAND2_X1 U25350 ( .A1(n24050), .A2(n23969), .ZN(n23975) );
  INV_X1 U25351 ( .A(n23970), .ZN(n23974) );
  INV_X1 U25352 ( .A(n24483), .ZN(n23971) );
  AND3_X1 U25353 ( .A1(n23972), .A2(n24480), .A3(n23971), .ZN(n23973) );
  XNOR2_X1 U25355 ( .A(n25187), .B(n28485), .ZN(n25713) );
  INV_X1 U25356 ( .A(n24556), .ZN(n24174) );
  NOR2_X1 U25357 ( .A1(n24174), .A2(n24552), .ZN(n23977) );
  MUX2_X1 U25358 ( .A(n24555), .B(n24551), .S(n24173), .Z(n23976) );
  NAND2_X1 U25359 ( .A1(n23981), .A2(n23980), .ZN(n25270) );
  NAND2_X1 U25361 ( .A1(n29642), .A2(n24642), .ZN(n24639) );
  NOR2_X1 U25362 ( .A1(n24237), .A2(n24644), .ZN(n24231) );
  NAND2_X1 U25363 ( .A1(n24231), .A2(n24568), .ZN(n23987) );
  INV_X1 U25364 ( .A(n24645), .ZN(n24232) );
  NAND2_X1 U25365 ( .A1(n2209), .A2(n24638), .ZN(n23985) );
  OAI211_X1 U25366 ( .C1(n24232), .C2(n2209), .A(n29645), .B(n23985), .ZN(
        n23986) );
  OAI211_X1 U25367 ( .C1(n2209), .C2(n24639), .A(n23987), .B(n23986), .ZN(
        n24984) );
  XNOR2_X1 U25368 ( .A(n28534), .B(n25781), .ZN(n23988) );
  XNOR2_X1 U25369 ( .A(n25056), .B(n23988), .ZN(n24011) );
  INV_X1 U25370 ( .A(n24634), .ZN(n24557) );
  NOR2_X1 U25371 ( .A1(n24637), .A2(n23990), .ZN(n23991) );
  NOR2_X2 U25372 ( .A1(n23992), .A2(n23991), .ZN(n25516) );
  NAND2_X1 U25373 ( .A1(n24380), .A2(n24372), .ZN(n23993) );
  OAI21_X1 U25374 ( .B1(n24373), .B2(n24380), .A(n23993), .ZN(n23999) );
  NAND2_X1 U25375 ( .A1(n24373), .A2(n24374), .ZN(n23997) );
  XNOR2_X1 U25378 ( .A(n28654), .B(n2996), .ZN(n24000) );
  XNOR2_X1 U25379 ( .A(n25516), .B(n24000), .ZN(n24009) );
  MUX2_X1 U25380 ( .A(n24542), .B(n2823), .S(n24541), .Z(n24004) );
  OAI22_X1 U25381 ( .A1(n24547), .A2(n24002), .B1(n24542), .B2(n24159), .ZN(
        n24003) );
  XNOR2_X1 U25384 ( .A(n26109), .B(n25577), .ZN(n24008) );
  XNOR2_X1 U25385 ( .A(n24009), .B(n24008), .ZN(n24010) );
  XNOR2_X1 U25386 ( .A(n24011), .B(n24010), .ZN(n26454) );
  NAND2_X1 U25387 ( .A1(n26452), .A2(n26454), .ZN(n25415) );
  NOR2_X1 U25388 ( .A1(n26456), .A2(n25415), .ZN(n24038) );
  NOR2_X1 U25389 ( .A1(n24972), .A2(n471), .ZN(n24974) );
  INV_X1 U25390 ( .A(n24012), .ZN(n24980) );
  AOI21_X1 U25391 ( .B1(n24976), .B2(n24974), .A(n24980), .ZN(n24013) );
  OAI21_X1 U25392 ( .B1(n24014), .B2(n23597), .A(n24013), .ZN(n24018) );
  MUX2_X1 U25393 ( .A(n24610), .B(n24614), .S(n24613), .Z(n24015) );
  INV_X1 U25394 ( .A(n24015), .ZN(n24016) );
  INV_X1 U25395 ( .A(n24017), .ZN(n24609) );
  XNOR2_X1 U25396 ( .A(n24018), .B(n24852), .ZN(n26013) );
  XNOR2_X1 U25398 ( .A(n25381), .B(n2522), .ZN(n24021) );
  XNOR2_X1 U25399 ( .A(n26013), .B(n24021), .ZN(n24036) );
  NAND2_X1 U25402 ( .A1(n462), .A2(n24751), .ZN(n24618) );
  OAI21_X1 U25403 ( .B1(n28223), .B2(n24024), .A(n24618), .ZN(n24025) );
  INV_X1 U25404 ( .A(n28785), .ZN(n24029) );
  AOI21_X1 U25405 ( .B1(n1955), .B2(n24792), .A(n24507), .ZN(n24034) );
  MUX2_X1 U25406 ( .A(n24789), .B(n24794), .S(n28455), .Z(n24033) );
  NOR2_X1 U25407 ( .A1(n28455), .A2(n24791), .ZN(n24032) );
  XNOR2_X1 U25409 ( .A(n25703), .B(n29073), .ZN(n25408) );
  XNOR2_X1 U25410 ( .A(n25412), .B(n25408), .ZN(n24035) );
  XNOR2_X1 U25411 ( .A(n24035), .B(n24036), .ZN(n26450) );
  INV_X1 U25412 ( .A(n26450), .ZN(n26162) );
  NAND3_X1 U25413 ( .A1(n26162), .A2(n26448), .A3(n26449), .ZN(n24037) );
  MUX2_X1 U25414 ( .A(n29308), .B(n24776), .S(n24777), .Z(n24043) );
  NAND2_X1 U25415 ( .A1(n24040), .A2(n24779), .ZN(n24042) );
  NAND3_X1 U25416 ( .A1(n23946), .A2(n24776), .A3(n29308), .ZN(n24041) );
  OAI211_X1 U25417 ( .C1(n24043), .C2(n463), .A(n24042), .B(n24041), .ZN(
        n26084) );
  XNOR2_X1 U25418 ( .A(n26084), .B(n25943), .ZN(n25569) );
  NAND2_X1 U25419 ( .A1(n24758), .A2(n29592), .ZN(n24449) );
  INV_X1 U25420 ( .A(n24449), .ZN(n24045) );
  OAI21_X1 U25421 ( .B1(n29592), .B2(n24756), .A(n23588), .ZN(n24044) );
  NAND2_X1 U25422 ( .A1(n24479), .A2(n24483), .ZN(n24048) );
  OAI21_X2 U25424 ( .B1(n24050), .B2(n24479), .A(n24049), .ZN(n25454) );
  XNOR2_X1 U25425 ( .A(n25454), .B(n26053), .ZN(n24051) );
  XNOR2_X1 U25426 ( .A(n25569), .B(n24051), .ZN(n24063) );
  NOR2_X1 U25427 ( .A1(n24584), .A2(n24582), .ZN(n24053) );
  NOR2_X1 U25428 ( .A1(n24583), .A2(n29025), .ZN(n24052) );
  NAND2_X1 U25429 ( .A1(n24577), .A2(n24584), .ZN(n24466) );
  MUX2_X1 U25431 ( .A(n24057), .B(n23922), .S(n24610), .Z(n24058) );
  XNOR2_X1 U25433 ( .A(n25722), .B(n24061), .ZN(n24062) );
  NOR2_X1 U25435 ( .A1(n25006), .A2(n25005), .ZN(n24366) );
  NOR2_X1 U25436 ( .A1(n24366), .A2(n24304), .ZN(n24066) );
  OAI21_X1 U25437 ( .B1(n23897), .B2(n24066), .A(n24065), .ZN(n26019) );
  XNOR2_X1 U25438 ( .A(n26019), .B(n25190), .ZN(n24070) );
  XNOR2_X1 U25439 ( .A(n25910), .B(n25809), .ZN(n25590) );
  XNOR2_X1 U25440 ( .A(n25590), .B(n24070), .ZN(n24089) );
  NOR2_X1 U25441 ( .A1(n24666), .A2(n24072), .ZN(n24071) );
  INV_X1 U25442 ( .A(n24074), .ZN(n24669) );
  AOI22_X1 U25443 ( .A1(n28424), .A2(n24075), .B1(n24383), .B2(n24669), .ZN(
        n24076) );
  AOI21_X1 U25444 ( .B1(n24077), .B2(n24388), .A(n24079), .ZN(n24082) );
  XNOR2_X1 U25445 ( .A(n25398), .B(n25251), .ZN(n25743) );
  OAI21_X1 U25446 ( .B1(n24403), .B2(n24408), .A(n24084), .ZN(n24086) );
  INV_X1 U25447 ( .A(n2961), .ZN(n27333) );
  XNOR2_X1 U25448 ( .A(n29039), .B(n27333), .ZN(n24087) );
  XNOR2_X1 U25449 ( .A(n24087), .B(n25743), .ZN(n24088) );
  INV_X1 U25450 ( .A(n24090), .ZN(n24098) );
  INV_X1 U25451 ( .A(n24093), .ZN(n24094) );
  XNOR2_X1 U25452 ( .A(n25037), .B(n25509), .ZN(n24110) );
  INV_X1 U25453 ( .A(n24712), .ZN(n24104) );
  AOI21_X1 U25454 ( .B1(n24720), .B2(n24711), .A(n24104), .ZN(n24108) );
  AOI21_X1 U25455 ( .B1(n4136), .B2(n24412), .A(n24712), .ZN(n24107) );
  NOR2_X1 U25456 ( .A1(n24716), .A2(n4136), .ZN(n24105) );
  XNOR2_X1 U25457 ( .A(n25385), .B(n2960), .ZN(n24109) );
  XNOR2_X1 U25458 ( .A(n24110), .B(n24109), .ZN(n24131) );
  NOR2_X1 U25459 ( .A1(n24520), .A2(n24516), .ZN(n24112) );
  NOR2_X1 U25460 ( .A1(n24111), .A2(n24517), .ZN(n24180) );
  MUX2_X1 U25461 ( .A(n24112), .B(n24180), .S(n24514), .Z(n24116) );
  OAI21_X1 U25462 ( .B1(n24420), .B2(n24113), .A(n24516), .ZN(n24114) );
  NOR2_X1 U25463 ( .A1(n24180), .A2(n24114), .ZN(n24115) );
  XNOR2_X1 U25464 ( .A(n28402), .B(n25751), .ZN(n24129) );
  NAND2_X1 U25465 ( .A1(n24347), .A2(n24433), .ZN(n24119) );
  INV_X1 U25466 ( .A(n24434), .ZN(n24117) );
  NAND2_X1 U25467 ( .A1(n24338), .A2(n29043), .ZN(n24123) );
  NAND3_X1 U25468 ( .A1(n24707), .A2(n24417), .A3(n5571), .ZN(n24126) );
  XNOR2_X1 U25469 ( .A(n25513), .B(n26110), .ZN(n25387) );
  XNOR2_X1 U25470 ( .A(n25387), .B(n24129), .ZN(n24130) );
  XNOR2_X1 U25471 ( .A(n24130), .B(n24131), .ZN(n25317) );
  INV_X1 U25472 ( .A(n25317), .ZN(n26181) );
  NOR2_X1 U25473 ( .A1(n811), .A2(n29470), .ZN(n24136) );
  XNOR2_X1 U25474 ( .A(n25563), .B(n24137), .ZN(n24152) );
  NOR2_X1 U25475 ( .A1(n24367), .A2(n24369), .ZN(n25009) );
  AOI211_X1 U25476 ( .C1(n24369), .C2(n24368), .A(n28415), .B(n24138), .ZN(
        n24140) );
  NAND2_X1 U25477 ( .A1(n24278), .A2(n24141), .ZN(n24588) );
  INV_X1 U25478 ( .A(n24142), .ZN(n24146) );
  NOR2_X1 U25479 ( .A1(n22356), .A2(n24735), .ZN(n24740) );
  OAI211_X1 U25480 ( .C1(n29050), .C2(n24280), .A(n24736), .B(n24601), .ZN(
        n24150) );
  XNOR2_X1 U25481 ( .A(n25735), .B(n26007), .ZN(n24151) );
  XNOR2_X1 U25482 ( .A(n24151), .B(n24152), .ZN(n25666) );
  INV_X1 U25483 ( .A(n25666), .ZN(n26180) );
  NAND3_X1 U25484 ( .A1(n26181), .A2(n26180), .A3(n28561), .ZN(n24202) );
  NOR2_X1 U25485 ( .A1(n26186), .A2(n29528), .ZN(n24171) );
  INV_X1 U25486 ( .A(n24256), .ZN(n24508) );
  MUX2_X1 U25487 ( .A(n24651), .B(n28785), .S(n24653), .Z(n24156) );
  INV_X1 U25488 ( .A(n24248), .ZN(n24526) );
  OAI21_X1 U25489 ( .B1(n24526), .B2(n28785), .A(n24249), .ZN(n24649) );
  MUX2_X1 U25490 ( .A(n24794), .B(n24789), .S(n28455), .Z(n24158) );
  MUX2_X1 U25491 ( .A(n24793), .B(n24791), .S(n1955), .Z(n24157) );
  XNOR2_X1 U25492 ( .A(n25901), .B(n26041), .ZN(n25015) );
  XNOR2_X1 U25493 ( .A(n25903), .B(n25727), .ZN(n24168) );
  NOR2_X1 U25497 ( .A1(n29120), .A2(n24162), .ZN(n24163) );
  NAND2_X1 U25498 ( .A1(n24163), .A2(n6600), .ZN(n24164) );
  XNOR2_X1 U25499 ( .A(n26039), .B(n24166), .ZN(n24167) );
  XNOR2_X1 U25500 ( .A(n24167), .B(n24168), .ZN(n24169) );
  NAND2_X1 U25501 ( .A1(n24171), .A2(n28547), .ZN(n24201) );
  NOR2_X1 U25502 ( .A1(n28519), .A2(n24552), .ZN(n24554) );
  AOI21_X1 U25503 ( .B1(n24174), .B2(n24173), .A(n24554), .ZN(n24177) );
  OAI22_X1 U25504 ( .A1(n24175), .A2(n24178), .B1(n24556), .B2(n24553), .ZN(
        n24176) );
  NAND2_X1 U25506 ( .A1(n24179), .A2(n24514), .ZN(n24185) );
  NOR2_X1 U25507 ( .A1(n24179), .A2(n24420), .ZN(n24181) );
  AOI21_X1 U25508 ( .B1(n24181), .B2(n24520), .A(n24180), .ZN(n24184) );
  AND2_X1 U25509 ( .A1(n24516), .A2(n24514), .ZN(n24182) );
  NAND2_X1 U25510 ( .A1(n24520), .A2(n24182), .ZN(n24183) );
  OAI211_X1 U25511 ( .C1(n24520), .C2(n24185), .A(n24184), .B(n24183), .ZN(
        n25932) );
  XNOR2_X1 U25512 ( .A(n25932), .B(n28520), .ZN(n24187) );
  XNOR2_X1 U25513 ( .A(n25931), .B(n2274), .ZN(n24186) );
  XNOR2_X1 U25514 ( .A(n24187), .B(n24186), .ZN(n24199) );
  MUX2_X1 U25515 ( .A(n24436), .B(n24437), .S(n24347), .Z(n24191) );
  OAI21_X1 U25516 ( .B1(n403), .B2(n29726), .A(n24188), .ZN(n24190) );
  NAND2_X1 U25518 ( .A1(n2619), .A2(n24434), .ZN(n24189) );
  XNOR2_X1 U25519 ( .A(n25179), .B(n25440), .ZN(n25763) );
  INV_X1 U25520 ( .A(n24241), .ZN(n24242) );
  MUX2_X1 U25521 ( .A(n24557), .B(n24192), .S(n24633), .Z(n24193) );
  OAI21_X2 U25522 ( .B1(n24194), .B2(n25794), .A(n24193), .ZN(n25702) );
  XNOR2_X1 U25523 ( .A(n26102), .B(n25702), .ZN(n26015) );
  XNOR2_X1 U25524 ( .A(n25763), .B(n26015), .ZN(n24198) );
  OAI21_X1 U25525 ( .B1(n24204), .B2(n26181), .A(n24203), .ZN(n27032) );
  INV_X1 U25526 ( .A(n24205), .ZN(n24460) );
  NOR2_X1 U25528 ( .A1(n24816), .A2(n24817), .ZN(n24206) );
  AOI21_X2 U25529 ( .B1(n24207), .B2(n24208), .A(n24206), .ZN(n26046) );
  XNOR2_X1 U25530 ( .A(n26046), .B(n25107), .ZN(n25429) );
  INV_X1 U25531 ( .A(n24776), .ZN(n24457) );
  XNOR2_X1 U25532 ( .A(n25429), .B(n25081), .ZN(n24226) );
  XNOR2_X1 U25533 ( .A(n26044), .B(n25727), .ZN(n24224) );
  NOR2_X1 U25534 ( .A1(n24758), .A2(n24216), .ZN(n24222) );
  NOR2_X1 U25535 ( .A1(n24222), .A2(n24221), .ZN(n25498) );
  XNOR2_X1 U25536 ( .A(n25498), .B(n3211), .ZN(n24223) );
  XNOR2_X1 U25537 ( .A(n24224), .B(n24223), .ZN(n24225) );
  XNOR2_X2 U25538 ( .A(n24226), .B(n24225), .ZN(n27395) );
  INV_X1 U25539 ( .A(n27395), .ZN(n26195) );
  OAI21_X1 U25540 ( .B1(n24630), .B2(n24293), .A(n24295), .ZN(n24228) );
  XNOR2_X1 U25542 ( .A(n26023), .B(n25134), .ZN(n25806) );
  XNOR2_X1 U25543 ( .A(n28628), .B(n25396), .ZN(n24230) );
  XNOR2_X1 U25544 ( .A(n25806), .B(n24230), .ZN(n24255) );
  NAND2_X1 U25545 ( .A1(n24231), .A2(n24642), .ZN(n24235) );
  INV_X1 U25546 ( .A(n24638), .ZN(n24564) );
  OAI21_X1 U25547 ( .B1(n24232), .B2(n24564), .A(n24643), .ZN(n24233) );
  NAND2_X1 U25548 ( .A1(n24233), .A2(n29645), .ZN(n24234) );
  OAI21_X1 U25550 ( .B1(n24633), .B2(n465), .A(n24634), .ZN(n24238) );
  XNOR2_X1 U25552 ( .A(n25065), .B(n25745), .ZN(n25449) );
  NAND2_X1 U25553 ( .A1(n24247), .A2(n28481), .ZN(n24252) );
  NAND2_X1 U25554 ( .A1(n24249), .A2(n24248), .ZN(n24250) );
  INV_X1 U25555 ( .A(n24653), .ZN(n24655) );
  NAND2_X1 U25556 ( .A1(n24250), .A2(n24655), .ZN(n24251) );
  NAND2_X1 U25557 ( .A1(n24252), .A2(n24251), .ZN(n24963) );
  XNOR2_X1 U25558 ( .A(n26120), .B(n26701), .ZN(n24253) );
  XNOR2_X1 U25559 ( .A(n25449), .B(n24253), .ZN(n24254) );
  XNOR2_X1 U25560 ( .A(n25346), .B(n25059), .ZN(n25772) );
  XNOR2_X1 U25561 ( .A(n25773), .B(n300), .ZN(n24264) );
  XNOR2_X1 U25562 ( .A(n25772), .B(n24264), .ZN(n24276) );
  NAND3_X1 U25563 ( .A1(n24748), .A2(n24751), .A3(n24747), .ZN(n24267) );
  OAI211_X1 U25564 ( .C1(n28550), .C2(n24747), .A(n24267), .B(n24266), .ZN(
        n25736) );
  XNOR2_X1 U25565 ( .A(n25738), .B(n29017), .ZN(n24274) );
  INV_X1 U25566 ( .A(n24791), .ZN(n24268) );
  OAI211_X1 U25567 ( .C1(n24792), .C2(n24268), .A(n24793), .B(n24789), .ZN(
        n24271) );
  NAND3_X1 U25568 ( .A1(n28512), .A2(n24269), .A3(n4576), .ZN(n24270) );
  NAND3_X1 U25569 ( .A1(n24271), .A2(n24270), .A3(n6943), .ZN(n24272) );
  XNOR2_X1 U25570 ( .A(n26095), .B(n6653), .ZN(n24273) );
  XNOR2_X1 U25571 ( .A(n24274), .B(n24273), .ZN(n24275) );
  XNOR2_X1 U25572 ( .A(n24276), .B(n24275), .ZN(n26464) );
  NOR2_X1 U25573 ( .A1(n24593), .A2(n24278), .ZN(n24589) );
  XNOR2_X1 U25574 ( .A(n26011), .B(n25820), .ZN(n25277) );
  NAND2_X1 U25575 ( .A1(n24282), .A2(n24280), .ZN(n24284) );
  NAND2_X1 U25576 ( .A1(n22311), .A2(n24602), .ZN(n24600) );
  NAND3_X1 U25577 ( .A1(n24282), .A2(n24736), .A3(n24734), .ZN(n24283) );
  OAI211_X1 U25578 ( .C1(n22356), .C2(n24284), .A(n24600), .B(n24283), .ZN(
        n24286) );
  XNOR2_X1 U25580 ( .A(n25381), .B(n25341), .ZN(n24287) );
  XNOR2_X1 U25581 ( .A(n24287), .B(n25277), .ZN(n24302) );
  AOI22_X1 U25582 ( .A1(n24596), .A2(n24728), .B1(n24730), .B2(n24729), .ZN(
        n24292) );
  INV_X1 U25583 ( .A(n24598), .ZN(n24289) );
  NAND2_X1 U25585 ( .A1(n4364), .A2(n24295), .ZN(n24296) );
  XNOR2_X1 U25586 ( .A(n25760), .B(n25890), .ZN(n24300) );
  XNOR2_X1 U25587 ( .A(n25179), .B(n3423), .ZN(n24299) );
  XNOR2_X1 U25588 ( .A(n24300), .B(n24299), .ZN(n24301) );
  XNOR2_X1 U25590 ( .A(n24306), .B(n25782), .ZN(n24308) );
  XNOR2_X1 U25591 ( .A(n24308), .B(n24307), .ZN(n24329) );
  NAND2_X1 U25593 ( .A1(n29567), .A2(n24310), .ZN(n24312) );
  NOR2_X1 U25596 ( .A1(n24668), .A2(n24383), .ZN(n24317) );
  INV_X1 U25598 ( .A(n24383), .ZN(n24318) );
  NAND3_X1 U25599 ( .A1(n24667), .A2(n24669), .A3(n24318), .ZN(n24319) );
  XNOR2_X1 U25600 ( .A(n25386), .B(n25780), .ZN(n24328) );
  NOR3_X1 U25601 ( .A1(n29555), .A2(n24677), .A3(n24676), .ZN(n24325) );
  NOR2_X2 U25602 ( .A1(n24326), .A2(n24325), .ZN(n26108) );
  INV_X1 U25603 ( .A(n26108), .ZN(n24327) );
  XNOR2_X1 U25604 ( .A(n24328), .B(n24327), .ZN(n25040) );
  XNOR2_X1 U25605 ( .A(n24329), .B(n25040), .ZN(n26194) );
  INV_X1 U25606 ( .A(n26194), .ZN(n25404) );
  INV_X1 U25608 ( .A(n25375), .ZN(n24330) );
  INV_X1 U25609 ( .A(n24772), .ZN(n24331) );
  NOR2_X1 U25610 ( .A1(n24697), .A2(n29624), .ZN(n24332) );
  AOI22_X1 U25611 ( .A1(n24699), .A2(n24768), .B1(n24765), .B2(n24332), .ZN(
        n24333) );
  INV_X1 U25612 ( .A(n24334), .ZN(n24335) );
  NOR3_X1 U25613 ( .A1(n24337), .A2(n24336), .A3(n24335), .ZN(n24340) );
  NAND3_X1 U25614 ( .A1(n24341), .A2(n24417), .A3(n29043), .ZN(n24343) );
  XNOR2_X1 U25617 ( .A(n25458), .B(n24345), .ZN(n24360) );
  AND3_X2 U25620 ( .A1(n24349), .A2(n24348), .A3(n6945), .ZN(n25535) );
  XNOR2_X1 U25621 ( .A(n24949), .B(n25535), .ZN(n24358) );
  NOR2_X1 U25622 ( .A1(n24714), .A2(n24713), .ZN(n24350) );
  MUX2_X1 U25623 ( .A(n24351), .B(n24350), .S(n24712), .Z(n24355) );
  XNOR2_X1 U25624 ( .A(n25149), .B(n24356), .ZN(n24357) );
  XNOR2_X1 U25625 ( .A(n24358), .B(n24357), .ZN(n24359) );
  OAI21_X1 U25627 ( .B1(n25404), .B2(n26469), .A(n27394), .ZN(n24361) );
  OAI211_X1 U25628 ( .C1(n26195), .C2(n25406), .A(n24362), .B(n24361), .ZN(
        n27026) );
  NAND2_X1 U25629 ( .A1(n27032), .A2(n27026), .ZN(n24363) );
  NAND2_X1 U25630 ( .A1(n26705), .A2(n26819), .ZN(n24828) );
  INV_X1 U25631 ( .A(n27026), .ZN(n26817) );
  NOR2_X1 U25632 ( .A1(n24366), .A2(n24365), .ZN(n24371) );
  MUX2_X1 U25633 ( .A(n25005), .B(n24368), .S(n24367), .Z(n24370) );
  NOR2_X1 U25635 ( .A1(n29340), .A2(n24374), .ZN(n24379) );
  XNOR2_X1 U25636 ( .A(n25352), .B(n25430), .ZN(n24389) );
  MUX2_X1 U25637 ( .A(n24667), .B(n4605), .S(n24669), .Z(n24385) );
  XNOR2_X1 U25639 ( .A(n24389), .B(n25541), .ZN(n24402) );
  MUX2_X1 U25640 ( .A(n466), .B(n29471), .S(n24390), .Z(n24394) );
  INV_X1 U25641 ( .A(n24682), .ZN(n24392) );
  INV_X1 U25642 ( .A(n24688), .ZN(n24681) );
  OAI21_X1 U25644 ( .B1(n24397), .B2(n24678), .A(n24396), .ZN(n24398) );
  XNOR2_X1 U25645 ( .A(n25689), .B(n25900), .ZN(n25354) );
  XNOR2_X1 U25646 ( .A(n26045), .B(n3109), .ZN(n24400) );
  XNOR2_X1 U25647 ( .A(n25354), .B(n24400), .ZN(n24401) );
  OR2_X1 U25648 ( .A1(n24405), .A2(n24404), .ZN(n24406) );
  NAND2_X1 U25649 ( .A1(n24720), .A2(n24713), .ZN(n24414) );
  XNOR2_X1 U25651 ( .A(n25550), .B(n25345), .ZN(n26091) );
  NAND2_X1 U25652 ( .A1(n24416), .A2(n24415), .ZN(n24419) );
  AND2_X1 U25653 ( .A1(n24420), .A2(n24514), .ZN(n24423) );
  XNOR2_X1 U25654 ( .A(n25737), .B(n25864), .ZN(n24425) );
  XNOR2_X1 U25655 ( .A(n26091), .B(n24425), .ZN(n24446) );
  XNOR2_X1 U25656 ( .A(n25867), .B(n25708), .ZN(n24444) );
  NOR2_X1 U25657 ( .A1(n24434), .A2(n24433), .ZN(n24441) );
  OR2_X1 U25658 ( .A1(n24435), .A2(n29726), .ZN(n24440) );
  NAND3_X1 U25659 ( .A1(n29726), .A2(n24437), .A3(n29128), .ZN(n24439) );
  XNOR2_X1 U25660 ( .A(n25564), .B(n26825), .ZN(n24443) );
  XNOR2_X1 U25661 ( .A(n24444), .B(n24443), .ZN(n24445) );
  XNOR2_X1 U25662 ( .A(n24446), .B(n24445), .ZN(n26559) );
  NOR2_X1 U25663 ( .A1(n28385), .A2(n26559), .ZN(n24576) );
  NAND2_X1 U25664 ( .A1(n24449), .A2(n24448), .ZN(n24452) );
  AOI21_X1 U25665 ( .B1(n24757), .B2(n24756), .A(n24450), .ZN(n24451) );
  AOI22_X1 U25666 ( .A1(n24452), .A2(n24451), .B1(n24758), .B2(n24757), .ZN(
        n25182) );
  XNOR2_X1 U25667 ( .A(n24453), .B(n25441), .ZN(n24465) );
  NAND2_X1 U25668 ( .A1(n24780), .A2(n24776), .ZN(n24455) );
  NAND2_X1 U25669 ( .A1(n1426), .A2(n24779), .ZN(n24459) );
  AND3_X1 U25670 ( .A1(n24457), .A2(n24775), .A3(n24779), .ZN(n24458) );
  NAND2_X1 U25671 ( .A1(n24812), .A2(n24460), .ZN(n24464) );
  NOR2_X1 U25672 ( .A1(n24812), .A2(n24814), .ZN(n24498) );
  OAI21_X1 U25673 ( .B1(n24498), .B2(n24808), .A(n24817), .ZN(n24463) );
  XNOR2_X1 U25675 ( .A(n25889), .B(n29155), .ZN(n25340) );
  XNOR2_X1 U25676 ( .A(n24465), .B(n25340), .ZN(n24488) );
  NAND2_X1 U25677 ( .A1(n24583), .A2(n24467), .ZN(n24469) );
  NAND3_X1 U25678 ( .A1(n24471), .A2(n24470), .A3(n24491), .ZN(n24478) );
  AOI22_X1 U25679 ( .A1(n24473), .A2(n23842), .B1(n24474), .B2(n24489), .ZN(
        n24477) );
  NAND2_X1 U25680 ( .A1(n24475), .A2(n24474), .ZN(n24476) );
  NOR2_X1 U25681 ( .A1(n24479), .A2(n24483), .ZN(n24481) );
  XNOR2_X1 U25683 ( .A(n24487), .B(n26100), .ZN(n25529) );
  AOI21_X1 U25684 ( .B1(n24493), .B2(n24492), .A(n24491), .ZN(n24494) );
  INV_X1 U25685 ( .A(n24808), .ZN(n24497) );
  NAND2_X1 U25686 ( .A1(n24498), .A2(n220), .ZN(n24501) );
  NOR2_X1 U25687 ( .A1(n24503), .A2(n24801), .ZN(n24504) );
  NOR2_X1 U25688 ( .A1(n24504), .A2(n24802), .ZN(n24505) );
  XNOR2_X1 U25689 ( .A(n25844), .B(n25914), .ZN(n25330) );
  AOI21_X1 U25690 ( .B1(n24972), .B2(n24509), .A(n24508), .ZN(n24510) );
  NOR2_X1 U25691 ( .A1(n23467), .A2(n24510), .ZN(n24511) );
  NOR2_X2 U25692 ( .A1(n24512), .A2(n24511), .ZN(n26115) );
  OAI21_X1 U25693 ( .B1(n24518), .B2(n24517), .A(n24516), .ZN(n24519) );
  XNOR2_X1 U25694 ( .A(n26115), .B(n25909), .ZN(n24521) );
  XNOR2_X1 U25695 ( .A(n25330), .B(n24521), .ZN(n24522) );
  OAI21_X1 U25696 ( .B1(n24523), .B2(n3061), .A(n24653), .ZN(n24525) );
  NOR2_X1 U25697 ( .A1(n3061), .A2(n28785), .ZN(n24527) );
  NAND2_X1 U25698 ( .A1(n24527), .A2(n24526), .ZN(n24528) );
  XNOR2_X1 U25699 ( .A(n24529), .B(n26055), .ZN(n24549) );
  NOR2_X1 U25700 ( .A1(n23144), .A2(n24631), .ZN(n24893) );
  NAND2_X1 U25701 ( .A1(n4366), .A2(n24533), .ZN(n24628) );
  INV_X1 U25702 ( .A(n24628), .ZN(n24534) );
  NAND2_X1 U25703 ( .A1(n24534), .A2(n24631), .ZN(n24535) );
  AOI21_X1 U25705 ( .B1(n24542), .B2(n24541), .A(n23126), .ZN(n24546) );
  XNOR2_X1 U25707 ( .A(n26080), .B(n29606), .ZN(n25287) );
  XNOR2_X1 U25708 ( .A(n24549), .B(n25287), .ZN(n24574) );
  NOR2_X1 U25710 ( .A1(n24559), .A2(n24633), .ZN(n24636) );
  AOI22_X1 U25711 ( .A1(n24561), .A2(n24560), .B1(n24636), .B2(n465), .ZN(
        n24562) );
  NOR2_X1 U25712 ( .A1(n24644), .A2(n24564), .ZN(n24566) );
  NOR2_X1 U25713 ( .A1(n24644), .A2(n24638), .ZN(n24565) );
  AOI22_X1 U25714 ( .A1(n24566), .A2(n24642), .B1(n24565), .B2(n29643), .ZN(
        n24570) );
  NOR2_X1 U25715 ( .A1(n29643), .A2(n24643), .ZN(n24567) );
  NAND2_X1 U25716 ( .A1(n24568), .A2(n24567), .ZN(n24569) );
  XNOR2_X1 U25718 ( .A(n25696), .B(n25947), .ZN(n24572) );
  XNOR2_X1 U25719 ( .A(n26083), .B(n24572), .ZN(n24573) );
  NOR2_X1 U25720 ( .A1(n24578), .A2(n29026), .ZN(n24580) );
  NOR2_X1 U25721 ( .A1(n24583), .A2(n24582), .ZN(n24585) );
  OAI21_X1 U25722 ( .B1(n24586), .B2(n24585), .A(n24584), .ZN(n24587) );
  OAI21_X1 U25725 ( .B1(n24601), .B2(n24602), .A(n24744), .ZN(n24606) );
  AOI22_X1 U25726 ( .A1(n22356), .A2(n24604), .B1(n24603), .B2(n24602), .ZN(
        n24605) );
  XNOR2_X1 U25728 ( .A(n24608), .B(n29518), .ZN(n24625) );
  NOR3_X1 U25729 ( .A1(n459), .A2(n24609), .A3(n5168), .ZN(n24615) );
  MUX2_X1 U25730 ( .A(n24610), .B(n29109), .S(n24614), .Z(n24611) );
  AOI21_X1 U25731 ( .B1(n21303), .B2(n2879), .A(n24616), .ZN(n24623) );
  NOR2_X1 U25732 ( .A1(n24618), .A2(n24747), .ZN(n24619) );
  NOR2_X1 U25733 ( .A1(n24620), .A2(n24619), .ZN(n24621) );
  OAI21_X1 U25734 ( .B1(n24623), .B2(n28223), .A(n24621), .ZN(n25165) );
  NOR2_X1 U25736 ( .A1(n26457), .A2(n28578), .ZN(n26563) );
  NAND2_X1 U25737 ( .A1(n26563), .A2(n28385), .ZN(n24627) );
  NOR2_X1 U25738 ( .A1(n26458), .A2(n28578), .ZN(n25614) );
  NAND2_X1 U25739 ( .A1(n25614), .A2(n26559), .ZN(n24626) );
  OAI21_X1 U25740 ( .B1(n24630), .B2(n24629), .A(n24628), .ZN(n24632) );
  INV_X1 U25741 ( .A(n29645), .ZN(n24640) );
  OAI22_X1 U25742 ( .A1(n24641), .A2(n24640), .B1(n24639), .B2(n24638), .ZN(
        n24648) );
  MUX2_X1 U25743 ( .A(n24644), .B(n24643), .S(n24642), .Z(n24646) );
  NOR2_X1 U25744 ( .A1(n24646), .A2(n29642), .ZN(n24647) );
  XNOR2_X1 U25745 ( .A(n29069), .B(n25542), .ZN(n25294) );
  XNOR2_X1 U25746 ( .A(n25294), .B(n25207), .ZN(n24664) );
  NAND3_X1 U25747 ( .A1(n24649), .A2(n3697), .A3(n3061), .ZN(n24659) );
  XNOR2_X1 U25748 ( .A(n28785), .B(n629), .ZN(n24654) );
  NOR2_X1 U25749 ( .A1(n24653), .A2(n3697), .ZN(n24652) );
  AOI22_X1 U25750 ( .A1(n24654), .A2(n24653), .B1(n24652), .B2(n28481), .ZN(
        n24657) );
  NAND3_X1 U25751 ( .A1(n24660), .A2(n24659), .A3(n24658), .ZN(n24661) );
  XNOR2_X1 U25752 ( .A(n25352), .B(n24661), .ZN(n24662) );
  XNOR2_X1 U25753 ( .A(n28576), .B(n24662), .ZN(n24663) );
  XNOR2_X2 U25754 ( .A(n24664), .B(n24663), .ZN(n26927) );
  XNOR2_X1 U25755 ( .A(n25215), .B(n24671), .ZN(n24696) );
  XNOR2_X1 U25756 ( .A(n25345), .B(n29534), .ZN(n24694) );
  OAI211_X1 U25757 ( .C1(n24678), .C2(n404), .A(n24677), .B(n24676), .ZN(
        n24679) );
  NAND2_X1 U25758 ( .A1(n24680), .A2(n24679), .ZN(n25562) );
  AOI21_X1 U25759 ( .B1(n24683), .B2(n24682), .A(n24681), .ZN(n24693) );
  NAND4_X1 U25760 ( .A1(n24687), .A2(n24686), .A3(n24685), .A4(n24684), .ZN(
        n24690) );
  AOI21_X1 U25761 ( .B1(n24690), .B2(n29471), .A(n24688), .ZN(n24692) );
  OAI21_X1 U25762 ( .B1(n24693), .B2(n24692), .A(n24691), .ZN(n25549) );
  XNOR2_X1 U25763 ( .A(n25562), .B(n25549), .ZN(n25304) );
  XNOR2_X1 U25764 ( .A(n25304), .B(n24694), .ZN(n24695) );
  AND2_X1 U25767 ( .A1(n24765), .A2(n24768), .ZN(n24701) );
  XNOR2_X1 U25768 ( .A(n25927), .B(n25884), .ZN(n25298) );
  XNOR2_X1 U25769 ( .A(n25298), .B(n24703), .ZN(n24723) );
  MUX2_X1 U25770 ( .A(n24712), .B(n24714), .S(n24711), .Z(n24721) );
  NAND3_X1 U25771 ( .A1(n24715), .A2(n24714), .A3(n24713), .ZN(n24719) );
  NAND2_X1 U25772 ( .A1(n28416), .A2(n24716), .ZN(n24718) );
  OAI211_X2 U25773 ( .C1(n24721), .C2(n24720), .A(n24719), .B(n24718), .ZN(
        n25885) );
  XNOR2_X1 U25774 ( .A(n25932), .B(n25885), .ZN(n25486) );
  XNOR2_X1 U25775 ( .A(n25486), .B(n25113), .ZN(n24722) );
  XNOR2_X2 U25776 ( .A(n24722), .B(n24723), .ZN(n26933) );
  NOR2_X1 U25777 ( .A1(n24726), .A2(n24725), .ZN(n24727) );
  NAND2_X1 U25778 ( .A1(n24729), .A2(n24728), .ZN(n24731) );
  AOI21_X1 U25779 ( .B1(n24732), .B2(n24731), .A(n24730), .ZN(n24733) );
  NAND2_X1 U25780 ( .A1(n24740), .A2(n24739), .ZN(n24741) );
  XNOR2_X1 U25782 ( .A(n25531), .B(n29563), .ZN(n25288) );
  OAI21_X1 U25783 ( .B1(n28550), .B2(n24748), .A(n24747), .ZN(n24750) );
  XNOR2_X1 U25784 ( .A(n25288), .B(n25479), .ZN(n24755) );
  XNOR2_X1 U25785 ( .A(n28630), .B(n1187), .ZN(n24752) );
  XNOR2_X1 U25786 ( .A(n24753), .B(n24752), .ZN(n24754) );
  XNOR2_X1 U25787 ( .A(n24755), .B(n24754), .ZN(n26579) );
  NAND3_X1 U25788 ( .A1(n26927), .A2(n24788), .A3(n5505), .ZN(n24825) );
  XNOR2_X1 U25789 ( .A(n26115), .B(n29614), .ZN(n24764) );
  NAND2_X1 U25790 ( .A1(n24761), .A2(n24760), .ZN(n24762) );
  XNOR2_X1 U25791 ( .A(n25251), .B(n25810), .ZN(n25089) );
  XNOR2_X1 U25792 ( .A(n24764), .B(n25089), .ZN(n24787) );
  OAI21_X1 U25793 ( .B1(n24765), .B2(n1856), .A(n29624), .ZN(n24766) );
  OAI21_X1 U25794 ( .B1(n24772), .B2(n24771), .A(n24770), .ZN(n24773) );
  XNOR2_X1 U25795 ( .A(n29047), .B(n25845), .ZN(n24785) );
  NOR2_X1 U25796 ( .A1(n24777), .A2(n24776), .ZN(n24778) );
  OAI21_X1 U25797 ( .B1(n24778), .B2(n23946), .A(n463), .ZN(n24782) );
  XNOR2_X1 U25798 ( .A(n24785), .B(n24784), .ZN(n24786) );
  XNOR2_X1 U25799 ( .A(n24787), .B(n24786), .ZN(n25364) );
  INV_X1 U25800 ( .A(n25364), .ZN(n26926) );
  NAND2_X1 U25802 ( .A1(n26929), .A2(n24788), .ZN(n24824) );
  XNOR2_X1 U25803 ( .A(n25282), .B(n27730), .ZN(n24798) );
  OAI21_X1 U25804 ( .B1(n1955), .B2(n24791), .A(n28512), .ZN(n24796) );
  OAI21_X1 U25805 ( .B1(n24794), .B2(n24793), .A(n24792), .ZN(n24795) );
  XNOR2_X1 U25806 ( .A(n24797), .B(n25463), .ZN(n25753) );
  XNOR2_X1 U25807 ( .A(n24798), .B(n25753), .ZN(n24822) );
  OAI21_X1 U25808 ( .B1(n24801), .B2(n24800), .A(n28919), .ZN(n24807) );
  MUX2_X1 U25809 ( .A(n24809), .B(n24817), .S(n24808), .Z(n24811) );
  XNOR2_X1 U25810 ( .A(n25322), .B(n25509), .ZN(n25153) );
  XNOR2_X1 U25811 ( .A(n24923), .B(n25153), .ZN(n24821) );
  XNOR2_X1 U25812 ( .A(n24821), .B(n24822), .ZN(n26581) );
  XNOR2_X1 U25813 ( .A(n24829), .B(n622), .ZN(Ciphertext[31]) );
  XNOR2_X1 U25814 ( .A(n25366), .B(n26045), .ZN(n25080) );
  XNOR2_X1 U25815 ( .A(n25803), .B(n25080), .ZN(n24833) );
  XNOR2_X1 U25816 ( .A(n25901), .B(n25836), .ZN(n24831) );
  XNOR2_X1 U25817 ( .A(n26039), .B(n3751), .ZN(n24830) );
  XNOR2_X1 U25818 ( .A(n24831), .B(n24830), .ZN(n24832) );
  XNOR2_X1 U25819 ( .A(n24833), .B(n24832), .ZN(n26425) );
  XNOR2_X1 U25820 ( .A(n24834), .B(n25590), .ZN(n24837) );
  XNOR2_X1 U25821 ( .A(n29047), .B(n3695), .ZN(n24835) );
  XNOR2_X1 U25822 ( .A(n25069), .B(n24835), .ZN(n24836) );
  XNOR2_X1 U25823 ( .A(n24837), .B(n24836), .ZN(n26382) );
  INV_X1 U25824 ( .A(n26382), .ZN(n26361) );
  XNOR2_X1 U25825 ( .A(n25569), .B(n24948), .ZN(n24841) );
  XNOR2_X1 U25826 ( .A(n25826), .B(n29613), .ZN(n24839) );
  XNOR2_X1 U25827 ( .A(n26055), .B(n3752), .ZN(n24838) );
  XNOR2_X1 U25828 ( .A(n24839), .B(n24838), .ZN(n24840) );
  XNOR2_X1 U25829 ( .A(n25708), .B(n25346), .ZN(n26006) );
  XNOR2_X1 U25830 ( .A(n25391), .B(n25869), .ZN(n24938) );
  XNOR2_X1 U25831 ( .A(n24938), .B(n26006), .ZN(n24845) );
  XNOR2_X1 U25832 ( .A(n26093), .B(n25775), .ZN(n24843) );
  XNOR2_X1 U25833 ( .A(n25921), .B(n3378), .ZN(n24842) );
  XNOR2_X1 U25834 ( .A(n24843), .B(n24842), .ZN(n24844) );
  XNOR2_X1 U25835 ( .A(n24845), .B(n24844), .ZN(n26378) );
  NOR2_X1 U25836 ( .A1(n26426), .A2(n26378), .ZN(n24846) );
  XNOR2_X1 U25837 ( .A(n25037), .B(n25785), .ZN(n24913) );
  XNOR2_X1 U25838 ( .A(n24913), .B(n25056), .ZN(n24850) );
  XNOR2_X1 U25839 ( .A(n24847), .B(n25385), .ZN(n24848) );
  XNOR2_X1 U25840 ( .A(n26110), .B(n25324), .ZN(n26034) );
  XNOR2_X1 U25841 ( .A(n26034), .B(n24848), .ZN(n24849) );
  XNOR2_X1 U25842 ( .A(n24850), .B(n24849), .ZN(n26431) );
  XNOR2_X1 U25843 ( .A(n26011), .B(n25885), .ZN(n24851) );
  XNOR2_X1 U25844 ( .A(n26102), .B(n25444), .ZN(n25821) );
  XNOR2_X1 U25845 ( .A(n25821), .B(n24851), .ZN(n24855) );
  XNOR2_X1 U25846 ( .A(n25445), .B(n24852), .ZN(n25071) );
  XNOR2_X1 U25847 ( .A(n25931), .B(n3035), .ZN(n24853) );
  XNOR2_X1 U25848 ( .A(n25071), .B(n24853), .ZN(n24854) );
  XNOR2_X1 U25849 ( .A(n24854), .B(n24855), .ZN(n26381) );
  OAI21_X1 U25850 ( .B1(n26380), .B2(n26381), .A(n26426), .ZN(n24856) );
  INV_X1 U25852 ( .A(n27646), .ZN(n26978) );
  XNOR2_X1 U25853 ( .A(n25913), .B(n24858), .ZN(n25492) );
  XNOR2_X1 U25854 ( .A(n25492), .B(n25330), .ZN(n24862) );
  XNOR2_X1 U25855 ( .A(n28771), .B(n3787), .ZN(n24860) );
  XNOR2_X1 U25856 ( .A(n25808), .B(n26118), .ZN(n24859) );
  XNOR2_X1 U25857 ( .A(n24860), .B(n24859), .ZN(n24861) );
  XNOR2_X1 U25858 ( .A(n24862), .B(n24861), .ZN(n27178) );
  XNOR2_X1 U25859 ( .A(n25165), .B(n24984), .ZN(n26106) );
  XNOR2_X1 U25860 ( .A(n29518), .B(n26106), .ZN(n24866) );
  XNOR2_X1 U25861 ( .A(n25577), .B(n25509), .ZN(n24864) );
  INV_X1 U25862 ( .A(n730), .ZN(n27879) );
  XNOR2_X1 U25863 ( .A(n25209), .B(n27879), .ZN(n24863) );
  XNOR2_X1 U25864 ( .A(n24864), .B(n24863), .ZN(n24865) );
  XNOR2_X1 U25865 ( .A(n24866), .B(n24865), .ZN(n26129) );
  INV_X1 U25867 ( .A(n26264), .ZN(n27130) );
  XNOR2_X1 U25868 ( .A(n25790), .B(n26713), .ZN(n24867) );
  XNOR2_X1 U25869 ( .A(n25583), .B(n25903), .ZN(n25128) );
  XNOR2_X1 U25870 ( .A(n24867), .B(n25128), .ZN(n24869) );
  XNOR2_X1 U25871 ( .A(n26071), .B(n25369), .ZN(n25105) );
  XNOR2_X1 U25872 ( .A(n25105), .B(n25354), .ZN(n24868) );
  XNOR2_X1 U25873 ( .A(n24870), .B(n25855), .ZN(n25570) );
  XNOR2_X1 U25874 ( .A(n29094), .B(n25947), .ZN(n24871) );
  XNOR2_X1 U25875 ( .A(n24871), .B(n25570), .ZN(n24875) );
  XNOR2_X1 U25876 ( .A(n26080), .B(n25696), .ZN(n24872) );
  XNOR2_X1 U25877 ( .A(n24873), .B(n24872), .ZN(n24874) );
  XNOR2_X2 U25878 ( .A(n24875), .B(n24874), .ZN(n27175) );
  XNOR2_X1 U25879 ( .A(n25932), .B(n29073), .ZN(n25141) );
  XNOR2_X1 U25880 ( .A(n25112), .B(n25141), .ZN(n24879) );
  INV_X1 U25881 ( .A(n2411), .ZN(n27766) );
  XNOR2_X1 U25882 ( .A(n29053), .B(n27766), .ZN(n24876) );
  XNOR2_X1 U25883 ( .A(n24877), .B(n24876), .ZN(n24878) );
  XNOR2_X1 U25884 ( .A(n24879), .B(n24878), .ZN(n27177) );
  XNOR2_X1 U25885 ( .A(n25867), .B(n25737), .ZN(n25348) );
  XNOR2_X1 U25886 ( .A(n29067), .B(n25565), .ZN(n25102) );
  XNOR2_X1 U25887 ( .A(n25348), .B(n25102), .ZN(n24882) );
  XNOR2_X1 U25888 ( .A(n29634), .B(n4501), .ZN(n24880) );
  XNOR2_X1 U25889 ( .A(n25145), .B(n24880), .ZN(n24881) );
  MUX2_X1 U25890 ( .A(n27175), .B(n27178), .S(n26263), .Z(n24883) );
  NAND2_X1 U25891 ( .A1(n28392), .A2(n24883), .ZN(n24884) );
  XNOR2_X1 U25892 ( .A(n25262), .B(n25107), .ZN(n25791) );
  XNOR2_X1 U25893 ( .A(n24885), .B(n25791), .ZN(n24889) );
  XNOR2_X1 U25894 ( .A(n25542), .B(n25261), .ZN(n24887) );
  XNOR2_X1 U25895 ( .A(n25428), .B(n6319), .ZN(n24886) );
  XNOR2_X1 U25896 ( .A(n24887), .B(n24886), .ZN(n24888) );
  XNOR2_X2 U25897 ( .A(n24889), .B(n24888), .ZN(n27193) );
  AOI22_X1 U25898 ( .A1(n24894), .A2(n24893), .B1(n24892), .B2(n24891), .ZN(
        n24896) );
  NAND2_X1 U25899 ( .A1(n24896), .A2(n24895), .ZN(n25066) );
  XNOR2_X1 U25900 ( .A(n25251), .B(n25066), .ZN(n24899) );
  XNOR2_X1 U25901 ( .A(n24899), .B(n24898), .ZN(n24900) );
  XNOR2_X1 U25902 ( .A(n25549), .B(n365), .ZN(n24901) );
  XNOR2_X1 U25903 ( .A(n25099), .B(n24901), .ZN(n24905) );
  INV_X1 U25904 ( .A(n3369), .ZN(n24902) );
  XNOR2_X1 U25905 ( .A(n25921), .B(n24902), .ZN(n24903) );
  XNOR2_X1 U25906 ( .A(n25216), .B(n24903), .ZN(n24904) );
  XNOR2_X1 U25907 ( .A(n24905), .B(n24904), .ZN(n27190) );
  XNOR2_X1 U25908 ( .A(n25927), .B(n25381), .ZN(n24908) );
  XNOR2_X1 U25909 ( .A(n25440), .B(n24906), .ZN(n24907) );
  XNOR2_X1 U25910 ( .A(n24908), .B(n24907), .ZN(n24910) );
  XNOR2_X1 U25911 ( .A(n25820), .B(n25931), .ZN(n25029) );
  XNOR2_X1 U25912 ( .A(n25234), .B(n25029), .ZN(n24909) );
  INV_X1 U25914 ( .A(n2995), .ZN(n27444) );
  XNOR2_X1 U25915 ( .A(n25465), .B(n27444), .ZN(n24911) );
  XNOR2_X1 U25916 ( .A(n24911), .B(n25515), .ZN(n24912) );
  XNOR2_X1 U25917 ( .A(n25780), .B(n28402), .ZN(n25271) );
  XNOR2_X1 U25918 ( .A(n24912), .B(n25271), .ZN(n24915) );
  XNOR2_X1 U25919 ( .A(n24913), .B(n26029), .ZN(n24914) );
  AOI21_X1 U25921 ( .B1(n26140), .B2(n26290), .A(n27124), .ZN(n24922) );
  XNOR2_X1 U25922 ( .A(n29103), .B(n3372), .ZN(n24917) );
  XNOR2_X1 U25923 ( .A(n25375), .B(n24916), .ZN(n25456) );
  XNOR2_X1 U25924 ( .A(n25456), .B(n24917), .ZN(n24919) );
  XNOR2_X1 U25925 ( .A(n26054), .B(n25826), .ZN(n25225) );
  XNOR2_X1 U25926 ( .A(n25943), .B(n25149), .ZN(n25020) );
  XNOR2_X1 U25927 ( .A(n25225), .B(n25020), .ZN(n24918) );
  AOI21_X1 U25928 ( .B1(n24920), .B2(n27191), .A(n27193), .ZN(n24921) );
  NOR2_X2 U25929 ( .A1(n24922), .A2(n24921), .ZN(n27641) );
  AOI21_X1 U25930 ( .B1(n27637), .B2(n28466), .A(n27641), .ZN(n27640) );
  OAI21_X1 U25931 ( .B1(n3606), .B2(n26978), .A(n27640), .ZN(n24999) );
  XNOR2_X1 U25932 ( .A(n25786), .B(n25714), .ZN(n24924) );
  XNOR2_X1 U25933 ( .A(n25751), .B(n25385), .ZN(n24926) );
  XNOR2_X1 U25934 ( .A(n363), .B(n25909), .ZN(n24927) );
  XNOR2_X1 U25935 ( .A(n25810), .B(n28628), .ZN(n25589) );
  XNOR2_X1 U25936 ( .A(n25589), .B(n24927), .ZN(n24931) );
  XNOR2_X1 U25937 ( .A(n25398), .B(n3422), .ZN(n24929) );
  XNOR2_X1 U25938 ( .A(n29046), .B(n25191), .ZN(n24928) );
  XNOR2_X1 U25939 ( .A(n24929), .B(n24928), .ZN(n24930) );
  XNOR2_X1 U25941 ( .A(n24932), .B(n25885), .ZN(n24935) );
  INV_X1 U25942 ( .A(n3336), .ZN(n24933) );
  XNOR2_X1 U25943 ( .A(n28520), .B(n24933), .ZN(n24934) );
  XNOR2_X1 U25944 ( .A(n24935), .B(n24934), .ZN(n24937) );
  XNOR2_X1 U25945 ( .A(n25179), .B(n25819), .ZN(n24936) );
  XNOR2_X1 U25946 ( .A(n24936), .B(n25441), .ZN(n25560) );
  XNOR2_X1 U25947 ( .A(n25304), .B(n24938), .ZN(n24941) );
  XNOR2_X1 U25948 ( .A(n25738), .B(n25564), .ZN(n25188) );
  XNOR2_X1 U25949 ( .A(n25867), .B(n26314), .ZN(n24939) );
  XNOR2_X1 U25950 ( .A(n25188), .B(n24939), .ZN(n24940) );
  XNOR2_X1 U25951 ( .A(n24941), .B(n24940), .ZN(n27161) );
  XNOR2_X1 U25953 ( .A(n25430), .B(n25727), .ZN(n25174) );
  XNOR2_X1 U25954 ( .A(n25294), .B(n25174), .ZN(n24945) );
  XNOR2_X1 U25955 ( .A(n25366), .B(n25836), .ZN(n24943) );
  XNOR2_X1 U25956 ( .A(n25689), .B(n3770), .ZN(n24942) );
  XNOR2_X1 U25957 ( .A(n24943), .B(n24942), .ZN(n24944) );
  XNOR2_X2 U25958 ( .A(n24945), .B(n24944), .ZN(n27701) );
  XNOR2_X1 U25960 ( .A(n25288), .B(n24948), .ZN(n24952) );
  XNOR2_X1 U25961 ( .A(n24949), .B(n25948), .ZN(n25572) );
  XNOR2_X1 U25962 ( .A(n25696), .B(n3565), .ZN(n24950) );
  XNOR2_X1 U25963 ( .A(n25572), .B(n24950), .ZN(n24951) );
  XNOR2_X2 U25964 ( .A(n24952), .B(n24951), .ZN(n27704) );
  AND2_X1 U25965 ( .A1(n27704), .A2(n27702), .ZN(n26128) );
  INV_X1 U25966 ( .A(n27703), .ZN(n26350) );
  NAND2_X1 U25967 ( .A1(n27650), .A2(n27641), .ZN(n25001) );
  INV_X1 U25968 ( .A(n25001), .ZN(n25004) );
  INV_X1 U25969 ( .A(n25736), .ZN(n24954) );
  XNOR2_X1 U25970 ( .A(n25187), .B(n24954), .ZN(n26008) );
  XNOR2_X1 U25971 ( .A(n29533), .B(n29634), .ZN(n24955) );
  XNOR2_X1 U25972 ( .A(n25864), .B(n2982), .ZN(n24956) );
  XNOR2_X1 U25973 ( .A(n24272), .B(n25922), .ZN(n25547) );
  XNOR2_X1 U25974 ( .A(n24956), .B(n25547), .ZN(n24957) );
  INV_X1 U25975 ( .A(n26384), .ZN(n26387) );
  XNOR2_X1 U25976 ( .A(n25293), .B(n26040), .ZN(n25172) );
  XNOR2_X1 U25977 ( .A(n25260), .B(n25172), .ZN(n24962) );
  XNOR2_X1 U25978 ( .A(n26046), .B(n24959), .ZN(n24960) );
  INV_X1 U25979 ( .A(n25498), .ZN(n25351) );
  XNOR2_X1 U25980 ( .A(n25082), .B(n24960), .ZN(n24961) );
  XNOR2_X1 U25981 ( .A(n25133), .B(n25808), .ZN(n25254) );
  XNOR2_X1 U25982 ( .A(n25849), .B(n24963), .ZN(n25521) );
  XNOR2_X1 U25983 ( .A(n25254), .B(n25521), .ZN(n24967) );
  XNOR2_X1 U25984 ( .A(n25328), .B(n25845), .ZN(n24965) );
  INV_X1 U25985 ( .A(n3223), .ZN(n27263) );
  XNOR2_X1 U25986 ( .A(n25745), .B(n27263), .ZN(n24964) );
  XNOR2_X1 U25987 ( .A(n24965), .B(n24964), .ZN(n24966) );
  XNOR2_X2 U25988 ( .A(n24967), .B(n24966), .ZN(n27165) );
  MUX2_X1 U25989 ( .A(n26387), .B(n28572), .S(n27165), .Z(n24993) );
  XNOR2_X1 U25990 ( .A(n29094), .B(n25535), .ZN(n26086) );
  XNOR2_X1 U25991 ( .A(n25532), .B(n25534), .ZN(n25856) );
  XNOR2_X1 U25992 ( .A(n26086), .B(n25856), .ZN(n24971) );
  XNOR2_X1 U25993 ( .A(n26059), .B(n28630), .ZN(n24969) );
  XNOR2_X1 U25994 ( .A(n28465), .B(n27324), .ZN(n24968) );
  XNOR2_X1 U25995 ( .A(n24969), .B(n24968), .ZN(n24970) );
  NAND2_X1 U25996 ( .A1(n24973), .A2(n24972), .ZN(n24978) );
  NOR2_X1 U25997 ( .A1(n24975), .A2(n24974), .ZN(n24977) );
  XNOR2_X1 U26000 ( .A(n25341), .B(n25884), .ZN(n25485) );
  XNOR2_X1 U26001 ( .A(n25411), .B(n25485), .ZN(n24983) );
  NAND2_X1 U26002 ( .A1(n28642), .A2(n26386), .ZN(n24991) );
  XNOR2_X1 U26003 ( .A(n24984), .B(n3244), .ZN(n24985) );
  XNOR2_X1 U26004 ( .A(n25386), .B(n24985), .ZN(n24986) );
  XNOR2_X1 U26005 ( .A(n24986), .B(n25516), .ZN(n24989) );
  INV_X1 U26006 ( .A(n26028), .ZN(n24987) );
  XNOR2_X1 U26007 ( .A(n24987), .B(n25282), .ZN(n25167) );
  XNOR2_X1 U26008 ( .A(n25508), .B(n25876), .ZN(n25054) );
  XNOR2_X1 U26009 ( .A(n25167), .B(n25054), .ZN(n24988) );
  MUX2_X1 U26010 ( .A(n24991), .B(n24990), .S(n27165), .Z(n24992) );
  NOR2_X1 U26012 ( .A1(n29532), .A2(n25044), .ZN(n25003) );
  INV_X1 U26014 ( .A(n27640), .ZN(n24996) );
  NAND2_X1 U26015 ( .A1(n28466), .A2(n3606), .ZN(n25047) );
  INV_X1 U26016 ( .A(n25047), .ZN(n24994) );
  NAND3_X1 U26017 ( .A1(n24994), .A2(n27638), .A3(n29532), .ZN(n24995) );
  INV_X1 U26018 ( .A(n26671), .ZN(n27645) );
  NAND3_X1 U26019 ( .A1(n25001), .A2(n27645), .A3(n25044), .ZN(n25050) );
  NOR3_X1 U26020 ( .A1(n27637), .A2(n26978), .A3(n27645), .ZN(n25002) );
  AOI21_X1 U26021 ( .B1(n25004), .B2(n25003), .A(n25002), .ZN(n25049) );
  XNOR2_X1 U26022 ( .A(n1514), .B(n26119), .ZN(n25680) );
  INV_X1 U26024 ( .A(n25134), .ZN(n25010) );
  XNOR2_X1 U26025 ( .A(n28565), .B(n25010), .ZN(n25011) );
  XNOR2_X1 U26026 ( .A(n25680), .B(n25011), .ZN(n25014) );
  XNOR2_X1 U26027 ( .A(n25910), .B(n3180), .ZN(n25012) );
  XNOR2_X1 U26028 ( .A(n25449), .B(n25012), .ZN(n25013) );
  XNOR2_X1 U26030 ( .A(n25081), .B(n25015), .ZN(n25019) );
  XNOR2_X1 U26031 ( .A(n25352), .B(n26046), .ZN(n25017) );
  XNOR2_X1 U26032 ( .A(n29129), .B(n6016), .ZN(n25016) );
  XNOR2_X1 U26033 ( .A(n25017), .B(n25016), .ZN(n25018) );
  XNOR2_X1 U26034 ( .A(n25019), .B(n25018), .ZN(n25119) );
  XNOR2_X1 U26035 ( .A(n25020), .B(n25533), .ZN(n25023) );
  XNOR2_X1 U26036 ( .A(n26059), .B(n25361), .ZN(n25021) );
  XNOR2_X1 U26037 ( .A(n25697), .B(n25372), .ZN(n26081) );
  XNOR2_X1 U26038 ( .A(n26081), .B(n25021), .ZN(n25022) );
  INV_X1 U26040 ( .A(n27181), .ZN(n26396) );
  XNOR2_X1 U26041 ( .A(n25345), .B(n365), .ZN(n25024) );
  XNOR2_X1 U26042 ( .A(n300), .B(n25546), .ZN(n25711) );
  XNOR2_X1 U26043 ( .A(n25024), .B(n25711), .ZN(n25028) );
  XNOR2_X1 U26044 ( .A(n26094), .B(n25736), .ZN(n25026) );
  XNOR2_X1 U26045 ( .A(n25921), .B(n3154), .ZN(n25025) );
  XNOR2_X1 U26046 ( .A(n25026), .B(n25025), .ZN(n25027) );
  XNOR2_X1 U26047 ( .A(n25028), .B(n25027), .ZN(n25034) );
  INV_X1 U26048 ( .A(n25034), .ZN(n27183) );
  XNOR2_X1 U26049 ( .A(n25029), .B(n26101), .ZN(n25033) );
  XNOR2_X1 U26050 ( .A(n25890), .B(n25702), .ZN(n25031) );
  XNOR2_X1 U26051 ( .A(n25760), .B(n1215), .ZN(n25030) );
  XNOR2_X1 U26052 ( .A(n25031), .B(n25030), .ZN(n25032) );
  XNOR2_X1 U26053 ( .A(n25033), .B(n25032), .ZN(n25124) );
  NAND2_X1 U26055 ( .A1(n25035), .A2(n25034), .ZN(n25043) );
  INV_X1 U26056 ( .A(n3598), .ZN(n26814) );
  XNOR2_X1 U26057 ( .A(n25268), .B(n26814), .ZN(n25036) );
  XNOR2_X1 U26058 ( .A(n26109), .B(n25036), .ZN(n25039) );
  XNOR2_X1 U26059 ( .A(n25037), .B(n25322), .ZN(n25038) );
  XNOR2_X1 U26060 ( .A(n25039), .B(n25038), .ZN(n25041) );
  XNOR2_X1 U26061 ( .A(n25041), .B(n25040), .ZN(n25120) );
  INV_X1 U26062 ( .A(n25120), .ZN(n26356) );
  NAND3_X1 U26063 ( .A1(n27183), .A2(n28651), .A3(n26356), .ZN(n25042) );
  INV_X1 U26064 ( .A(n27639), .ZN(n26980) );
  NOR3_X1 U26065 ( .A1(n26980), .A2(n28466), .A3(n3606), .ZN(n25046) );
  NOR2_X1 U26066 ( .A1(n27639), .A2(n25044), .ZN(n25045) );
  OAI21_X1 U26067 ( .B1(n25046), .B2(n25045), .A(n29532), .ZN(n25048) );
  XNOR2_X1 U26070 ( .A(n25780), .B(n3036), .ZN(n25053) );
  XNOR2_X1 U26071 ( .A(n25385), .B(n25781), .ZN(n25055) );
  XNOR2_X1 U26072 ( .A(n25056), .B(n25055), .ZN(n25057) );
  XNOR2_X1 U26073 ( .A(n365), .B(n300), .ZN(n25061) );
  XNOR2_X1 U26074 ( .A(n25391), .B(n29111), .ZN(n25060) );
  XNOR2_X1 U26075 ( .A(n25708), .B(n25864), .ZN(n25063) );
  INV_X1 U26076 ( .A(Key[19]), .ZN(n25991) );
  XNOR2_X1 U26077 ( .A(n26095), .B(n25991), .ZN(n25062) );
  XNOR2_X1 U26078 ( .A(n25063), .B(n25062), .ZN(n25064) );
  NOR2_X1 U26079 ( .A1(n26172), .A2(n26173), .ZN(n25079) );
  XNOR2_X1 U26080 ( .A(n26114), .B(n25066), .ZN(n25068) );
  XNOR2_X1 U26081 ( .A(n25808), .B(n3622), .ZN(n25067) );
  XNOR2_X1 U26082 ( .A(n25068), .B(n25067), .ZN(n25070) );
  INV_X1 U26083 ( .A(Key[66]), .ZN(n27742) );
  XNOR2_X1 U26084 ( .A(n25341), .B(n25072), .ZN(n26104) );
  XNOR2_X1 U26085 ( .A(n25454), .B(n26055), .ZN(n25074) );
  XNOR2_X1 U26086 ( .A(n26086), .B(n25074), .ZN(n25078) );
  XNOR2_X1 U26087 ( .A(n25149), .B(n25534), .ZN(n25076) );
  XNOR2_X1 U26088 ( .A(n25697), .B(n3385), .ZN(n25075) );
  XNOR2_X1 U26089 ( .A(n25076), .B(n25075), .ZN(n25077) );
  XNOR2_X1 U26090 ( .A(n25081), .B(n25080), .ZN(n25085) );
  XNOR2_X1 U26091 ( .A(n25790), .B(n3728), .ZN(n25083) );
  XNOR2_X1 U26092 ( .A(n25082), .B(n25083), .ZN(n25084) );
  NOR2_X1 U26093 ( .A1(n26917), .A2(n26172), .ZN(n26781) );
  XNOR2_X1 U26094 ( .A(n25507), .B(n25753), .ZN(n25088) );
  XNOR2_X1 U26095 ( .A(n28654), .B(n25209), .ZN(n25388) );
  XNOR2_X1 U26096 ( .A(n29599), .B(n3323), .ZN(n25086) );
  XNOR2_X1 U26097 ( .A(n25388), .B(n25086), .ZN(n25087) );
  XNOR2_X1 U26098 ( .A(n25088), .B(n25087), .ZN(n26280) );
  XNOR2_X1 U26099 ( .A(n26020), .B(n29046), .ZN(n25493) );
  XNOR2_X1 U26100 ( .A(n25493), .B(n25089), .ZN(n25093) );
  XNOR2_X1 U26101 ( .A(n28769), .B(n3742), .ZN(n25091) );
  XNOR2_X1 U26102 ( .A(n26118), .B(n25396), .ZN(n25090) );
  XNOR2_X1 U26103 ( .A(n25091), .B(n25090), .ZN(n25092) );
  XNOR2_X1 U26106 ( .A(n25094), .B(n25456), .ZN(n25098) );
  XNOR2_X1 U26107 ( .A(n26054), .B(n29563), .ZN(n25096) );
  XNOR2_X1 U26108 ( .A(n3083), .B(n26080), .ZN(n25095) );
  XNOR2_X1 U26109 ( .A(n25095), .B(n25096), .ZN(n25097) );
  XNOR2_X1 U26112 ( .A(n26004), .B(n25562), .ZN(n25734) );
  XNOR2_X1 U26113 ( .A(n25099), .B(n25734), .ZN(n25104) );
  INV_X1 U26114 ( .A(n2389), .ZN(n25100) );
  XNOR2_X1 U26115 ( .A(n25869), .B(n25100), .ZN(n25101) );
  XNOR2_X1 U26116 ( .A(n25102), .B(n25101), .ZN(n25103) );
  XNOR2_X1 U26117 ( .A(n25104), .B(n25103), .ZN(n26278) );
  XNOR2_X1 U26118 ( .A(n25836), .B(n26038), .ZN(n25106) );
  XNOR2_X1 U26119 ( .A(n25105), .B(n25106), .ZN(n25111) );
  XNOR2_X1 U26120 ( .A(n29069), .B(n25261), .ZN(n25109) );
  XNOR2_X1 U26121 ( .A(n1922), .B(n2511), .ZN(n25108) );
  XNOR2_X1 U26122 ( .A(n25109), .B(n25108), .ZN(n25110) );
  XNOR2_X1 U26123 ( .A(n25112), .B(n25113), .ZN(n25117) );
  XNOR2_X1 U26124 ( .A(n25381), .B(n2987), .ZN(n25115) );
  XNOR2_X1 U26125 ( .A(n25761), .B(n25885), .ZN(n25114) );
  XNOR2_X1 U26126 ( .A(n25115), .B(n25114), .ZN(n25116) );
  XNOR2_X1 U26127 ( .A(n25116), .B(n25117), .ZN(n26797) );
  INV_X1 U26128 ( .A(n26797), .ZN(n26362) );
  INV_X1 U26129 ( .A(n25119), .ZN(n26397) );
  NOR2_X1 U26130 ( .A1(n26397), .A2(n27181), .ZN(n25123) );
  AND2_X1 U26131 ( .A1(n27182), .A2(n28467), .ZN(n25122) );
  NAND2_X1 U26132 ( .A1(n26357), .A2(n25124), .ZN(n26399) );
  INV_X1 U26133 ( .A(n27203), .ZN(n27538) );
  XNOR2_X1 U26134 ( .A(n26040), .B(n25262), .ZN(n25126) );
  XNOR2_X1 U26135 ( .A(n25689), .B(n25543), .ZN(n25839) );
  XNOR2_X1 U26136 ( .A(n25126), .B(n25839), .ZN(n25130) );
  XNOR2_X1 U26137 ( .A(n25352), .B(n28007), .ZN(n25127) );
  XNOR2_X1 U26138 ( .A(n25128), .B(n25127), .ZN(n25129) );
  XNOR2_X1 U26140 ( .A(n28565), .B(n363), .ZN(n25132) );
  XNOR2_X1 U26141 ( .A(n25132), .B(n25492), .ZN(n25138) );
  INV_X1 U26143 ( .A(n2946), .ZN(n26601) );
  XNOR2_X1 U26144 ( .A(n25328), .B(n26601), .ZN(n25135) );
  XNOR2_X1 U26145 ( .A(n25136), .B(n25135), .ZN(n25137) );
  XNOR2_X1 U26146 ( .A(n25889), .B(n25820), .ZN(n25139) );
  XNOR2_X1 U26147 ( .A(n25411), .B(n25139), .ZN(n25144) );
  XNOR2_X1 U26148 ( .A(n25140), .B(n25928), .ZN(n25142) );
  XNOR2_X1 U26149 ( .A(n25142), .B(n25141), .ZN(n25143) );
  XNOR2_X1 U26150 ( .A(n25143), .B(n25144), .ZN(n26769) );
  INV_X1 U26151 ( .A(n26769), .ZN(n26937) );
  XNOR2_X1 U26152 ( .A(n25922), .B(n25345), .ZN(n25146) );
  XNOR2_X1 U26153 ( .A(n28496), .B(n25146), .ZN(n25147) );
  XNOR2_X1 U26154 ( .A(n25148), .B(n25147), .ZN(n26936) );
  INV_X1 U26155 ( .A(n26772), .ZN(n25152) );
  INV_X1 U26156 ( .A(n25696), .ZN(n25151) );
  XNOR2_X1 U26157 ( .A(n25151), .B(n26083), .ZN(n25336) );
  INV_X1 U26158 ( .A(n26935), .ZN(n26944) );
  XNOR2_X1 U26159 ( .A(n25516), .B(n25714), .ZN(n25874) );
  XNOR2_X1 U26160 ( .A(n25874), .B(n25153), .ZN(n25157) );
  XNOR2_X1 U26161 ( .A(n28534), .B(n25577), .ZN(n25155) );
  XNOR2_X1 U26162 ( .A(n25780), .B(n28294), .ZN(n25154) );
  XNOR2_X1 U26163 ( .A(n25155), .B(n25154), .ZN(n25156) );
  XNOR2_X1 U26164 ( .A(n25157), .B(n25156), .ZN(n26943) );
  INV_X1 U26165 ( .A(n26943), .ZN(n26771) );
  INV_X1 U26166 ( .A(n26436), .ZN(n26768) );
  XNOR2_X1 U26167 ( .A(n25531), .B(n25947), .ZN(n25160) );
  XNOR2_X1 U26168 ( .A(n25160), .B(n25572), .ZN(n25164) );
  XNOR2_X1 U26169 ( .A(n26080), .B(n28630), .ZN(n25162) );
  XNOR2_X1 U26170 ( .A(n28465), .B(n3276), .ZN(n25161) );
  XNOR2_X1 U26171 ( .A(n25162), .B(n25161), .ZN(n25163) );
  XNOR2_X1 U26173 ( .A(n29599), .B(n25751), .ZN(n25166) );
  XNOR2_X1 U26174 ( .A(n25167), .B(n25166), .ZN(n25171) );
  XNOR2_X1 U26175 ( .A(n25754), .B(n25515), .ZN(n25169) );
  XNOR2_X1 U26176 ( .A(n25169), .B(n25168), .ZN(n25170) );
  INV_X1 U26178 ( .A(n25172), .ZN(n25173) );
  XNOR2_X1 U26179 ( .A(n25173), .B(n25174), .ZN(n25178) );
  XNOR2_X1 U26180 ( .A(n26071), .B(n25900), .ZN(n25176) );
  XNOR2_X1 U26181 ( .A(n25542), .B(n27231), .ZN(n25175) );
  XNOR2_X1 U26182 ( .A(n25176), .B(n25175), .ZN(n25177) );
  MUX2_X1 U26183 ( .A(n29071), .B(n29631), .S(n26950), .Z(n25197) );
  XNOR2_X1 U26184 ( .A(n25180), .B(n26100), .ZN(n25181) );
  XNOR2_X1 U26185 ( .A(n25411), .B(n25181), .ZN(n25184) );
  XNOR2_X1 U26186 ( .A(n25759), .B(n25182), .ZN(n25929) );
  XNOR2_X1 U26187 ( .A(n25929), .B(n25298), .ZN(n25183) );
  XNOR2_X1 U26188 ( .A(n25184), .B(n25183), .ZN(n26951) );
  INV_X1 U26189 ( .A(n26951), .ZN(n26948) );
  XNOR2_X1 U26190 ( .A(n25550), .B(n3414), .ZN(n25185) );
  XNOR2_X1 U26191 ( .A(n25185), .B(n29533), .ZN(n25186) );
  XNOR2_X1 U26192 ( .A(n25737), .B(n25549), .ZN(n25920) );
  XNOR2_X1 U26193 ( .A(n25186), .B(n25920), .ZN(n25189) );
  MUX2_X1 U26194 ( .A(n26948), .B(n28542), .S(n29071), .Z(n25196) );
  XNOR2_X1 U26195 ( .A(n25190), .B(n25914), .ZN(n25744) );
  XNOR2_X1 U26196 ( .A(n25191), .B(n25845), .ZN(n25312) );
  XNOR2_X1 U26197 ( .A(n25312), .B(n25744), .ZN(n25195) );
  XNOR2_X1 U26198 ( .A(n25328), .B(n25909), .ZN(n25193) );
  XNOR2_X1 U26199 ( .A(n26118), .B(n27605), .ZN(n25192) );
  XNOR2_X1 U26200 ( .A(n25193), .B(n25192), .ZN(n25194) );
  XNOR2_X1 U26201 ( .A(n25195), .B(n25194), .ZN(n26440) );
  INV_X1 U26203 ( .A(n26431), .ZN(n26275) );
  NAND3_X1 U26204 ( .A1(n26426), .A2(n26382), .A3(n26381), .ZN(n25198) );
  OAI21_X1 U26205 ( .B1(n26430), .B2(n26275), .A(n25198), .ZN(n25201) );
  INV_X1 U26206 ( .A(n26378), .ZN(n26427) );
  MUX2_X1 U26207 ( .A(n26427), .B(n26426), .S(n26381), .Z(n25199) );
  NOR2_X1 U26208 ( .A1(n26425), .A2(n25199), .ZN(n25200) );
  AOI22_X1 U26209 ( .A1(n27200), .A2(n27203), .B1(n27199), .B2(n27547), .ZN(
        n25202) );
  NAND2_X1 U26210 ( .A1(n25203), .A2(n25202), .ZN(n25204) );
  XNOR2_X1 U26211 ( .A(n25204), .B(n2912), .ZN(Ciphertext[74]) );
  XNOR2_X1 U26212 ( .A(n25205), .B(n25428), .ZN(n25206) );
  XNOR2_X1 U26213 ( .A(n25898), .B(n25206), .ZN(n25208) );
  XOR2_X1 U26214 ( .A(n25209), .B(n25509), .Z(n25210) );
  XNOR2_X1 U26215 ( .A(n25876), .B(n2446), .ZN(n25211) );
  XNOR2_X1 U26216 ( .A(n25864), .B(n25565), .ZN(n25214) );
  XNOR2_X1 U26217 ( .A(n25564), .B(n3191), .ZN(n25213) );
  XNOR2_X1 U26218 ( .A(n25214), .B(n25213), .ZN(n25218) );
  XNOR2_X1 U26219 ( .A(n25216), .B(n25215), .ZN(n25217) );
  NOR2_X1 U26220 ( .A1(n26731), .A2(n28560), .ZN(n25224) );
  XNOR2_X1 U26221 ( .A(n25681), .B(n29614), .ZN(n25219) );
  XNOR2_X1 U26222 ( .A(n25493), .B(n25219), .ZN(n25223) );
  XNOR2_X1 U26223 ( .A(n28771), .B(n27225), .ZN(n25221) );
  XNOR2_X1 U26224 ( .A(n25849), .B(n25909), .ZN(n25220) );
  XNOR2_X1 U26225 ( .A(n25220), .B(n25221), .ZN(n25222) );
  NOR2_X1 U26226 ( .A1(n25224), .A2(n1622), .ZN(n25231) );
  XNOR2_X1 U26227 ( .A(n25225), .B(n25479), .ZN(n25229) );
  XNOR2_X1 U26228 ( .A(n25944), .B(n29606), .ZN(n25227) );
  XNOR2_X1 U26229 ( .A(n25948), .B(n3321), .ZN(n25226) );
  XNOR2_X1 U26230 ( .A(n25227), .B(n25226), .ZN(n25228) );
  NOR2_X1 U26231 ( .A1(n25628), .A2(n29579), .ZN(n25230) );
  INV_X1 U26232 ( .A(n26729), .ZN(n26484) );
  XNOR2_X1 U26233 ( .A(n25441), .B(n25891), .ZN(n25232) );
  XNOR2_X1 U26234 ( .A(n25486), .B(n25232), .ZN(n25236) );
  INV_X1 U26235 ( .A(n2381), .ZN(n27961) );
  XNOR2_X1 U26236 ( .A(n25933), .B(n27961), .ZN(n25233) );
  XNOR2_X1 U26237 ( .A(n25234), .B(n25233), .ZN(n25235) );
  NOR3_X1 U26238 ( .A1(n26484), .A2(n29501), .A3(n1622), .ZN(n25237) );
  NOR2_X1 U26239 ( .A1(n26194), .A2(n25406), .ZN(n27393) );
  INV_X1 U26241 ( .A(n26466), .ZN(n25239) );
  XNOR2_X1 U26244 ( .A(n25532), .B(n27669), .ZN(n25244) );
  XNOR2_X1 U26245 ( .A(n26055), .B(n26053), .ZN(n25694) );
  XNOR2_X1 U26246 ( .A(n25245), .B(n25694), .ZN(n25248) );
  XNOR2_X1 U26247 ( .A(n25246), .B(n25149), .ZN(n25247) );
  XNOR2_X1 U26248 ( .A(n29612), .B(n25247), .ZN(n25830) );
  INV_X1 U26249 ( .A(n26754), .ZN(n26237) );
  XNOR2_X1 U26250 ( .A(n25249), .B(n26019), .ZN(n25253) );
  XNOR2_X1 U26251 ( .A(n25251), .B(n25250), .ZN(n25252) );
  XNOR2_X1 U26252 ( .A(n25253), .B(n25252), .ZN(n25256) );
  XNOR2_X1 U26253 ( .A(n25806), .B(n25254), .ZN(n25255) );
  XNOR2_X1 U26254 ( .A(n25255), .B(n25256), .ZN(n25267) );
  XNOR2_X1 U26256 ( .A(n26041), .B(n26045), .ZN(n25688) );
  XNOR2_X1 U26257 ( .A(n25260), .B(n25688), .ZN(n25266) );
  XNOR2_X1 U26258 ( .A(n28475), .B(n3586), .ZN(n25264) );
  XNOR2_X1 U26259 ( .A(n25261), .B(n25262), .ZN(n25263) );
  XNOR2_X1 U26260 ( .A(n25264), .B(n25263), .ZN(n25265) );
  INV_X1 U26261 ( .A(n25267), .ZN(n26241) );
  INV_X1 U26262 ( .A(n25268), .ZN(n25269) );
  XNOR2_X1 U26263 ( .A(n25270), .B(n25269), .ZN(n26030) );
  XNOR2_X1 U26264 ( .A(n25271), .B(n26030), .ZN(n25275) );
  XNOR2_X1 U26265 ( .A(n25324), .B(n29247), .ZN(n25272) );
  XNOR2_X1 U26266 ( .A(n25272), .B(n25781), .ZN(n25273) );
  XNOR2_X1 U26267 ( .A(n25273), .B(n25516), .ZN(n25274) );
  XNOR2_X1 U26268 ( .A(n25274), .B(n25275), .ZN(n26755) );
  XNOR2_X1 U26269 ( .A(n25412), .B(n25277), .ZN(n25281) );
  XNOR2_X1 U26270 ( .A(n24852), .B(n3374), .ZN(n25279) );
  XNOR2_X1 U26271 ( .A(n25702), .B(n25440), .ZN(n25278) );
  XNOR2_X1 U26272 ( .A(n25279), .B(n25278), .ZN(n25280) );
  XNOR2_X1 U26273 ( .A(n25281), .B(n25280), .ZN(n26240) );
  NAND2_X1 U26274 ( .A1(n26237), .A2(n25603), .ZN(n25357) );
  XNOR2_X1 U26275 ( .A(n25517), .B(n25875), .ZN(n25286) );
  XNOR2_X1 U26276 ( .A(n25786), .B(n25515), .ZN(n25284) );
  XNOR2_X1 U26277 ( .A(n1871), .B(n2916), .ZN(n25283) );
  XNOR2_X1 U26278 ( .A(n25284), .B(n25283), .ZN(n25285) );
  XNOR2_X1 U26279 ( .A(n25287), .B(n25288), .ZN(n25292) );
  XNOR2_X1 U26280 ( .A(n28630), .B(n25855), .ZN(n25290) );
  XNOR2_X1 U26281 ( .A(n25372), .B(n1927), .ZN(n25289) );
  XNOR2_X1 U26282 ( .A(n25290), .B(n25289), .ZN(n25291) );
  XNOR2_X1 U26283 ( .A(n25583), .B(n25293), .ZN(n25840) );
  XNOR2_X1 U26284 ( .A(n25294), .B(n25840), .ZN(n25297) );
  XNOR2_X1 U26285 ( .A(n29129), .B(n2894), .ZN(n25295) );
  XNOR2_X1 U26286 ( .A(n25541), .B(n25295), .ZN(n25296) );
  INV_X1 U26288 ( .A(n25659), .ZN(n26716) );
  XNOR2_X1 U26289 ( .A(n25298), .B(n25408), .ZN(n25302) );
  XNOR2_X1 U26290 ( .A(n26100), .B(n25819), .ZN(n25300) );
  XNOR2_X1 U26291 ( .A(n25891), .B(n26531), .ZN(n25299) );
  XNOR2_X1 U26292 ( .A(n25300), .B(n25299), .ZN(n25301) );
  XNOR2_X1 U26293 ( .A(n25302), .B(n25301), .ZN(n26718) );
  INV_X1 U26294 ( .A(n25868), .ZN(n25303) );
  XNOR2_X1 U26295 ( .A(n25303), .B(n29533), .ZN(n25474) );
  XNOR2_X1 U26296 ( .A(n25304), .B(n25474), .ZN(n25308) );
  XNOR2_X1 U26297 ( .A(n25864), .B(n28485), .ZN(n25306) );
  XNOR2_X1 U26298 ( .A(n29067), .B(n1062), .ZN(n25305) );
  XNOR2_X1 U26299 ( .A(n25306), .B(n25305), .ZN(n25307) );
  MUX2_X1 U26300 ( .A(n26718), .B(n28459), .S(n26717), .Z(n25315) );
  XNOR2_X1 U26301 ( .A(n25810), .B(n1246), .ZN(n25309) );
  XNOR2_X1 U26302 ( .A(n25310), .B(n25309), .ZN(n25314) );
  XNOR2_X1 U26303 ( .A(n25312), .B(n25311), .ZN(n25313) );
  NAND2_X1 U26305 ( .A1(n28503), .A2(n29528), .ZN(n25319) );
  NAND2_X1 U26306 ( .A1(n25666), .A2(n28525), .ZN(n25318) );
  MUX2_X1 U26307 ( .A(n25319), .B(n25318), .S(n28547), .Z(n25320) );
  XNOR2_X1 U26308 ( .A(n26107), .B(n29518), .ZN(n25327) );
  XNOR2_X1 U26309 ( .A(n1871), .B(n26028), .ZN(n25717) );
  XNOR2_X1 U26310 ( .A(n25324), .B(n2402), .ZN(n25325) );
  XNOR2_X1 U26311 ( .A(n25717), .B(n25325), .ZN(n25326) );
  XNOR2_X1 U26312 ( .A(n26115), .B(n25328), .ZN(n25329) );
  XNOR2_X1 U26313 ( .A(n25330), .B(n25329), .ZN(n25334) );
  XNOR2_X1 U26314 ( .A(n28645), .B(n29543), .ZN(n25332) );
  XNOR2_X1 U26315 ( .A(n26120), .B(n27956), .ZN(n25331) );
  XNOR2_X1 U26316 ( .A(n25332), .B(n25331), .ZN(n25333) );
  XNOR2_X1 U26317 ( .A(n25334), .B(n25333), .ZN(n25344) );
  INV_X1 U26318 ( .A(n25344), .ZN(n26235) );
  XNOR2_X1 U26319 ( .A(n25947), .B(n29612), .ZN(n25335) );
  XNOR2_X1 U26320 ( .A(n25336), .B(n25335), .ZN(n25339) );
  XNOR2_X1 U26321 ( .A(n25535), .B(n3686), .ZN(n25337) );
  XNOR2_X1 U26322 ( .A(n25698), .B(n25337), .ZN(n25338) );
  XNOR2_X1 U26323 ( .A(n25338), .B(n25339), .ZN(n25654) );
  XNOR2_X1 U26325 ( .A(n26011), .B(n3087), .ZN(n25342) );
  INV_X1 U26326 ( .A(n25341), .ZN(n25526) );
  XNOR2_X1 U26327 ( .A(n25526), .B(n25342), .ZN(n25343) );
  NOR2_X1 U26329 ( .A1(n26230), .A2(n26737), .ZN(n25349) );
  XNOR2_X1 U26330 ( .A(n26095), .B(Key[151]), .ZN(n25347) );
  XNOR2_X1 U26331 ( .A(n26077), .B(n25687), .ZN(n25356) );
  XNOR2_X1 U26332 ( .A(n28475), .B(n28097), .ZN(n25353) );
  XNOR2_X1 U26333 ( .A(n25354), .B(n25353), .ZN(n25355) );
  XNOR2_X1 U26334 ( .A(n25356), .B(n25355), .ZN(n25597) );
  INV_X1 U26335 ( .A(n25597), .ZN(n26200) );
  INV_X1 U26336 ( .A(n25357), .ZN(n25358) );
  XNOR2_X1 U26340 ( .A(n25367), .B(n25366), .ZN(n25368) );
  XNOR2_X1 U26341 ( .A(n26041), .B(n25369), .ZN(n25370) );
  XNOR2_X1 U26342 ( .A(n26039), .B(n25370), .ZN(n25371) );
  XNOR2_X1 U26343 ( .A(n25944), .B(n26053), .ZN(n25374) );
  XNOR2_X1 U26344 ( .A(n25372), .B(n2804), .ZN(n25373) );
  XNOR2_X1 U26345 ( .A(n25374), .B(n25373), .ZN(n25377) );
  XNOR2_X1 U26346 ( .A(n25454), .B(n26059), .ZN(n25721) );
  XNOR2_X1 U26347 ( .A(n25375), .B(n26084), .ZN(n25828) );
  XNOR2_X1 U26348 ( .A(n25721), .B(n25828), .ZN(n25376) );
  XNOR2_X1 U26349 ( .A(n25376), .B(n25377), .ZN(n26420) );
  INV_X1 U26350 ( .A(n26420), .ZN(n26567) );
  XNOR2_X1 U26351 ( .A(n25445), .B(n25703), .ZN(n25380) );
  XNOR2_X1 U26352 ( .A(n25933), .B(n25378), .ZN(n25379) );
  XNOR2_X1 U26353 ( .A(n25380), .B(n25379), .ZN(n25384) );
  INV_X1 U26354 ( .A(n25381), .ZN(n25382) );
  XNOR2_X1 U26355 ( .A(n25760), .B(n25382), .ZN(n25442) );
  XNOR2_X1 U26356 ( .A(n25442), .B(n26015), .ZN(n25383) );
  XNOR2_X1 U26357 ( .A(n25383), .B(n25384), .ZN(n26786) );
  XNOR2_X1 U26358 ( .A(n25386), .B(n25385), .ZN(n25756) );
  XNOR2_X1 U26359 ( .A(n25387), .B(n25756), .ZN(n25390) );
  XNOR2_X1 U26360 ( .A(n26109), .B(n1046), .ZN(n25389) );
  XNOR2_X1 U26361 ( .A(n25773), .B(n29017), .ZN(n25436) );
  XNOR2_X1 U26362 ( .A(n26094), .B(n2404), .ZN(n25393) );
  XNOR2_X1 U26363 ( .A(n25391), .B(n25565), .ZN(n25392) );
  XNOR2_X1 U26364 ( .A(n25393), .B(n25392), .ZN(n25394) );
  XNOR2_X1 U26365 ( .A(n28769), .B(n25396), .ZN(n25397) );
  XNOR2_X1 U26366 ( .A(n25680), .B(n25397), .ZN(n25401) );
  XNOR2_X1 U26367 ( .A(n25809), .B(n25745), .ZN(n26025) );
  XNOR2_X1 U26368 ( .A(n25398), .B(n3451), .ZN(n25399) );
  XNOR2_X1 U26369 ( .A(n26025), .B(n25399), .ZN(n25400) );
  NOR2_X1 U26370 ( .A1(n26912), .A2(n26914), .ZN(n26788) );
  NAND3_X1 U26372 ( .A1(n29617), .A2(n29028), .A3(n25239), .ZN(n25405) );
  XNOR2_X1 U26375 ( .A(n24852), .B(n2522), .ZN(n25410) );
  XNOR2_X1 U26376 ( .A(n25408), .B(n25381), .ZN(n25409) );
  XNOR2_X1 U26377 ( .A(n25410), .B(n25409), .ZN(n25414) );
  XNOR2_X1 U26378 ( .A(n25412), .B(n25411), .ZN(n25413) );
  NAND2_X1 U26379 ( .A1(n26179), .A2(n26448), .ZN(n26455) );
  AND2_X1 U26380 ( .A1(n26447), .A2(n26449), .ZN(n25416) );
  NOR2_X1 U26382 ( .A1(n26576), .A2(n28710), .ZN(n25419) );
  INV_X1 U26383 ( .A(n26576), .ZN(n25421) );
  NOR3_X1 U26384 ( .A1(n25421), .A2(n29576), .A3(n28711), .ZN(n25422) );
  NOR2_X1 U26386 ( .A1(n25426), .A2(n25425), .ZN(n25427) );
  XNOR2_X1 U26387 ( .A(n25427), .B(n3565), .ZN(Ciphertext[40]) );
  XNOR2_X1 U26388 ( .A(n25428), .B(n26070), .ZN(n25691) );
  XNOR2_X1 U26389 ( .A(n25429), .B(n25691), .ZN(n25434) );
  INV_X1 U26390 ( .A(n25430), .ZN(n25431) );
  XNOR2_X1 U26391 ( .A(n25431), .B(n3164), .ZN(n25432) );
  XNOR2_X2 U26392 ( .A(n25434), .B(n25433), .ZN(n26222) );
  XNOR2_X1 U26393 ( .A(n25564), .B(n3501), .ZN(n25435) );
  XNOR2_X1 U26394 ( .A(n25436), .B(n25435), .ZN(n25439) );
  XNOR2_X1 U26395 ( .A(n25775), .B(n300), .ZN(n25437) );
  XNOR2_X1 U26396 ( .A(n25735), .B(n25437), .ZN(n25438) );
  NOR2_X1 U26398 ( .A1(n26222), .A2(n29100), .ZN(n25462) );
  XNOR2_X1 U26399 ( .A(n25441), .B(n25440), .ZN(n25443) );
  XNOR2_X1 U26400 ( .A(n25442), .B(n25443), .ZN(n25448) );
  XNOR2_X1 U26401 ( .A(n25890), .B(n25444), .ZN(n25701) );
  XNOR2_X1 U26402 ( .A(n28520), .B(n3015), .ZN(n25446) );
  XNOR2_X1 U26403 ( .A(n25446), .B(n25701), .ZN(n25447) );
  XNOR2_X1 U26404 ( .A(n25807), .B(n25449), .ZN(n25452) );
  XNOR2_X1 U26405 ( .A(n25909), .B(n3049), .ZN(n25450) );
  XNOR2_X1 U26406 ( .A(n25743), .B(n25450), .ZN(n25451) );
  XNOR2_X1 U26407 ( .A(n25452), .B(n25451), .ZN(n26749) );
  INV_X1 U26408 ( .A(n26749), .ZN(n25453) );
  XNOR2_X1 U26409 ( .A(n25826), .B(n25454), .ZN(n25455) );
  XNOR2_X1 U26410 ( .A(n25456), .B(n25455), .ZN(n25460) );
  XNOR2_X1 U26411 ( .A(n25948), .B(n3643), .ZN(n25457) );
  XNOR2_X1 U26412 ( .A(n25458), .B(n25457), .ZN(n25459) );
  XNOR2_X1 U26413 ( .A(n25459), .B(n25460), .ZN(n26746) );
  XNOR2_X1 U26415 ( .A(n28402), .B(n26108), .ZN(n25464) );
  XNOR2_X1 U26416 ( .A(n25756), .B(n25464), .ZN(n25469) );
  XNOR2_X1 U26417 ( .A(n25782), .B(n1923), .ZN(n25466) );
  XNOR2_X1 U26418 ( .A(n25467), .B(n25466), .ZN(n25468) );
  NOR2_X1 U26419 ( .A1(n29159), .A2(n26747), .ZN(n25645) );
  NAND2_X1 U26420 ( .A1(n25645), .A2(n26222), .ZN(n25471) );
  XNOR2_X1 U26421 ( .A(n26004), .B(n25737), .ZN(n25473) );
  XNOR2_X1 U26422 ( .A(n25474), .B(n25473), .ZN(n25478) );
  XNOR2_X1 U26423 ( .A(n25869), .B(n2981), .ZN(n25476) );
  XNOR2_X1 U26427 ( .A(n25947), .B(n26054), .ZN(n25724) );
  XNOR2_X1 U26428 ( .A(n25724), .B(n25479), .ZN(n25483) );
  XNOR2_X1 U26429 ( .A(n25855), .B(n25535), .ZN(n25481) );
  XNOR2_X1 U26430 ( .A(n25858), .B(n3633), .ZN(n25480) );
  XNOR2_X1 U26431 ( .A(n25481), .B(n25480), .ZN(n25482) );
  XNOR2_X1 U26433 ( .A(n25486), .B(n25485), .ZN(n25491) );
  INV_X1 U26434 ( .A(n25886), .ZN(n25487) );
  XNOR2_X1 U26435 ( .A(n29154), .B(n25487), .ZN(n25489) );
  XNOR2_X1 U26436 ( .A(n25761), .B(n3462), .ZN(n25488) );
  XNOR2_X1 U26437 ( .A(n25489), .B(n25488), .ZN(n25490) );
  XNOR2_X1 U26438 ( .A(n25491), .B(n25490), .ZN(n27014) );
  NAND2_X1 U26439 ( .A1(n26623), .A2(n27014), .ZN(n25505) );
  XNOR2_X1 U26440 ( .A(n25493), .B(n25492), .ZN(n25497) );
  XNOR2_X1 U26441 ( .A(n25914), .B(n25845), .ZN(n25495) );
  XNOR2_X1 U26442 ( .A(n26120), .B(n3491), .ZN(n25494) );
  XNOR2_X1 U26443 ( .A(n25495), .B(n25494), .ZN(n25496) );
  XNOR2_X1 U26445 ( .A(n25498), .B(n3660), .ZN(n25499) );
  XNOR2_X1 U26446 ( .A(n25499), .B(n25900), .ZN(n25500) );
  XNOR2_X1 U26447 ( .A(n25840), .B(n25500), .ZN(n25501) );
  NAND2_X1 U26448 ( .A1(n28639), .A2(n27052), .ZN(n25506) );
  NOR2_X1 U26449 ( .A1(n27052), .A2(n27013), .ZN(n25504) );
  XNOR2_X1 U26450 ( .A(n25507), .B(n25875), .ZN(n25512) );
  XNOR2_X1 U26451 ( .A(n25508), .B(n3463), .ZN(n25510) );
  XNOR2_X1 U26452 ( .A(n29485), .B(n25509), .ZN(n25940) );
  XNOR2_X1 U26453 ( .A(n25510), .B(n25940), .ZN(n25511) );
  NOR2_X1 U26454 ( .A1(n29160), .A2(n28025), .ZN(n28039) );
  XNOR2_X1 U26455 ( .A(n25513), .B(n2598), .ZN(n25514) );
  XNOR2_X1 U26456 ( .A(n26107), .B(n25514), .ZN(n25519) );
  XNOR2_X1 U26457 ( .A(n25516), .B(n25515), .ZN(n25942) );
  XNOR2_X1 U26458 ( .A(n25517), .B(n25942), .ZN(n25518) );
  XNOR2_X1 U26459 ( .A(n25518), .B(n25519), .ZN(n27043) );
  XNOR2_X1 U26460 ( .A(n26118), .B(n3483), .ZN(n25520) );
  XNOR2_X1 U26461 ( .A(n25521), .B(n25520), .ZN(n25524) );
  XNOR2_X1 U26462 ( .A(n26115), .B(n26019), .ZN(n25522) );
  XNOR2_X1 U26463 ( .A(n25915), .B(n25522), .ZN(n25523) );
  XNOR2_X1 U26464 ( .A(n25702), .B(n3212), .ZN(n25525) );
  XNOR2_X1 U26465 ( .A(n25927), .B(n25525), .ZN(n25528) );
  XNOR2_X1 U26466 ( .A(n25526), .B(n25928), .ZN(n25527) );
  XNOR2_X1 U26467 ( .A(n25528), .B(n25527), .ZN(n25530) );
  XNOR2_X1 U26468 ( .A(n25529), .B(n25530), .ZN(n27048) );
  INV_X1 U26469 ( .A(n29570), .ZN(n27004) );
  XNOR2_X1 U26470 ( .A(n29103), .B(n25532), .ZN(n25945) );
  XNOR2_X1 U26471 ( .A(n25945), .B(n25533), .ZN(n25539) );
  XNOR2_X1 U26472 ( .A(n25535), .B(n29606), .ZN(n25537) );
  XNOR2_X1 U26473 ( .A(n26080), .B(n3380), .ZN(n25536) );
  XNOR2_X1 U26474 ( .A(n25536), .B(n25537), .ZN(n25538) );
  OAI21_X1 U26476 ( .B1(n27001), .B2(n27004), .A(n28783), .ZN(n25556) );
  XNOR2_X1 U26477 ( .A(n26041), .B(n1123), .ZN(n25540) );
  XNOR2_X1 U26478 ( .A(n25541), .B(n25540), .ZN(n25545) );
  XNOR2_X1 U26479 ( .A(n25542), .B(n25543), .ZN(n25899) );
  XNOR2_X1 U26480 ( .A(n26077), .B(n25899), .ZN(n25544) );
  XNOR2_X1 U26481 ( .A(n25546), .B(n25345), .ZN(n25548) );
  XNOR2_X1 U26482 ( .A(n25548), .B(n25547), .ZN(n25554) );
  XNOR2_X1 U26483 ( .A(n25864), .B(n25549), .ZN(n25552) );
  XNOR2_X1 U26484 ( .A(n29067), .B(n1175), .ZN(n25551) );
  XNOR2_X1 U26485 ( .A(n25552), .B(n25551), .ZN(n25553) );
  NOR2_X1 U26488 ( .A1(n28039), .A2(n29031), .ZN(n25607) );
  XNOR2_X1 U26489 ( .A(n26102), .B(n25931), .ZN(n25558) );
  XNOR2_X1 U26490 ( .A(n25559), .B(n25558), .ZN(n25561) );
  XNOR2_X1 U26491 ( .A(n26093), .B(n25562), .ZN(n25771) );
  XNOR2_X1 U26492 ( .A(n25771), .B(n25563), .ZN(n25568) );
  XNOR2_X1 U26493 ( .A(n25565), .B(n25564), .ZN(n25919) );
  XNOR2_X1 U26494 ( .A(n25868), .B(n1248), .ZN(n25566) );
  XNOR2_X1 U26495 ( .A(n25919), .B(n25566), .ZN(n25567) );
  INV_X1 U26497 ( .A(n26998), .ZN(n25575) );
  XNOR2_X1 U26498 ( .A(n25569), .B(n25570), .ZN(n25574) );
  XNOR2_X1 U26499 ( .A(n25825), .B(n3457), .ZN(n25571) );
  XNOR2_X1 U26500 ( .A(n25572), .B(n25571), .ZN(n25573) );
  INV_X1 U26503 ( .A(n26997), .ZN(n25588) );
  XNOR2_X1 U26504 ( .A(n25939), .B(n25576), .ZN(n25581) );
  XNOR2_X1 U26505 ( .A(n25786), .B(n25577), .ZN(n25579) );
  XNOR2_X1 U26506 ( .A(n26110), .B(n25751), .ZN(n25578) );
  XNOR2_X1 U26507 ( .A(n25579), .B(n25578), .ZN(n25580) );
  XNOR2_X1 U26508 ( .A(n25581), .B(n25580), .ZN(n26733) );
  XNOR2_X1 U26509 ( .A(n25901), .B(n25727), .ZN(n25582) );
  XNOR2_X1 U26510 ( .A(n25898), .B(n25582), .ZN(n25587) );
  XNOR2_X1 U26511 ( .A(n25729), .B(n28540), .ZN(n25585) );
  XNOR2_X1 U26512 ( .A(n26039), .B(n3710), .ZN(n25584) );
  XNOR2_X1 U26513 ( .A(n25585), .B(n25584), .ZN(n25586) );
  MUX2_X1 U26514 ( .A(n25588), .B(n26733), .S(n26995), .Z(n25595) );
  XNOR2_X1 U26515 ( .A(n25589), .B(n25590), .ZN(n25594) );
  XNOR2_X1 U26516 ( .A(n25848), .B(n25909), .ZN(n25592) );
  XNOR2_X1 U26517 ( .A(n28771), .B(n3528), .ZN(n25591) );
  XNOR2_X1 U26518 ( .A(n25592), .B(n25591), .ZN(n25593) );
  INV_X1 U26519 ( .A(n25654), .ZN(n26203) );
  OAI22_X1 U26520 ( .A1(n26204), .A2(n26230), .B1(n26203), .B2(n26229), .ZN(
        n25598) );
  INV_X1 U26521 ( .A(n26204), .ZN(n26228) );
  AOI22_X1 U26522 ( .A1(n26741), .A2(n26228), .B1(n26230), .B2(n26200), .ZN(
        n25599) );
  INV_X1 U26524 ( .A(n28038), .ZN(n25601) );
  AOI21_X1 U26525 ( .B1(n26237), .B2(n25603), .A(n25602), .ZN(n25605) );
  NAND2_X1 U26526 ( .A1(n26753), .A2(n26755), .ZN(n25604) );
  OAI21_X1 U26527 ( .B1(n25605), .B2(n26753), .A(n25604), .ZN(n25606) );
  INV_X1 U26528 ( .A(n25649), .ZN(n26242) );
  NOR2_X1 U26529 ( .A1(n25606), .A2(n26242), .ZN(n26658) );
  NOR2_X1 U26530 ( .A1(n26760), .A2(n26240), .ZN(n26659) );
  NOR2_X1 U26531 ( .A1(n26658), .A2(n26659), .ZN(n26602) );
  OAI22_X1 U26532 ( .A1(n25607), .A2(n28035), .B1(n26664), .B2(n26602), .ZN(
        n25608) );
  XNOR2_X1 U26533 ( .A(n25608), .B(n2117), .ZN(Ciphertext[179]) );
  INV_X1 U26534 ( .A(n28547), .ZN(n25670) );
  NAND2_X1 U26535 ( .A1(n26181), .A2(n28503), .ZN(n26477) );
  NOR2_X1 U26536 ( .A1(n25670), .A2(n26477), .ZN(n25612) );
  OAI21_X1 U26537 ( .B1(n26186), .B2(n26185), .A(n26476), .ZN(n25609) );
  AOI21_X1 U26538 ( .B1(n26182), .B2(n28503), .A(n25609), .ZN(n25610) );
  INV_X1 U26539 ( .A(n27407), .ZN(n27402) );
  NOR2_X1 U26540 ( .A1(n28476), .A2(n28434), .ZN(n25613) );
  NOR2_X1 U26541 ( .A1(n25614), .A2(n25613), .ZN(n26159) );
  OAI21_X1 U26542 ( .B1(n26560), .B2(n28434), .A(n377), .ZN(n25615) );
  NAND2_X1 U26543 ( .A1(n28385), .A2(n25615), .ZN(n25616) );
  NAND2_X1 U26545 ( .A1(n27402), .A2(n27386), .ZN(n27404) );
  INV_X1 U26548 ( .A(n25622), .ZN(n25624) );
  OAI21_X1 U26549 ( .B1(n26448), .B2(n26449), .A(n26162), .ZN(n25623) );
  NOR2_X1 U26550 ( .A1(n25624), .A2(n25623), .ZN(n25626) );
  NOR2_X1 U26551 ( .A1(n26454), .A2(n26448), .ZN(n25625) );
  OAI211_X1 U26552 ( .C1(n27404), .C2(n28607), .A(n25627), .B(n1175), .ZN(
        n25634) );
  NAND2_X1 U26553 ( .A1(n28548), .A2(n29560), .ZN(n25665) );
  INV_X1 U26554 ( .A(n26715), .ZN(n26209) );
  INV_X1 U26556 ( .A(n26721), .ZN(n26208) );
  INV_X1 U26557 ( .A(n26718), .ZN(n26215) );
  OAI21_X1 U26558 ( .B1(n26723), .B2(n26208), .A(n26215), .ZN(n25631) );
  NAND2_X1 U26559 ( .A1(n27402), .A2(n27387), .ZN(n25636) );
  NOR2_X1 U26560 ( .A1(n26960), .A2(n1175), .ZN(n25635) );
  OAI211_X1 U26561 ( .C1(n27410), .C2(n27402), .A(n25636), .B(n25635), .ZN(
        n25637) );
  NAND2_X1 U26562 ( .A1(n25638), .A2(n25637), .ZN(n25639) );
  NOR2_X1 U26563 ( .A1(n25640), .A2(n25639), .ZN(Ciphertext[20]) );
  NOR2_X1 U26564 ( .A1(n29501), .A2(n28560), .ZN(n25641) );
  NAND2_X1 U26565 ( .A1(n25453), .A2(n26747), .ZN(n25647) );
  NAND2_X1 U26566 ( .A1(n29099), .A2(n26747), .ZN(n25642) );
  NAND2_X1 U26567 ( .A1(n5760), .A2(n25642), .ZN(n25643) );
  OAI21_X1 U26568 ( .B1(n25645), .B2(n25644), .A(n25643), .ZN(n25646) );
  OAI21_X1 U26569 ( .B1(n5035), .B2(n25647), .A(n25646), .ZN(n27354) );
  INV_X1 U26570 ( .A(n27354), .ZN(n25657) );
  NOR2_X1 U26571 ( .A1(n27340), .A2(n25657), .ZN(n25658) );
  INV_X1 U26573 ( .A(n25650), .ZN(n25653) );
  NOR2_X1 U26574 ( .A1(n26761), .A2(n26237), .ZN(n25652) );
  NAND2_X1 U26575 ( .A1(n26241), .A2(n26755), .ZN(n25651) );
  AOI22_X2 U26576 ( .A1(n25975), .A2(n25653), .B1(n25652), .B2(n25651), .ZN(
        n27358) );
  INV_X1 U26577 ( .A(n27358), .ZN(n27350) );
  INV_X1 U26578 ( .A(n26742), .ZN(n25656) );
  NOR2_X1 U26579 ( .A1(n26204), .A2(n25597), .ZN(n26738) );
  NOR2_X1 U26580 ( .A1(n26203), .A2(n26740), .ZN(n25655) );
  NOR2_X1 U26581 ( .A1(n28473), .A2(n25654), .ZN(n26739) );
  INV_X1 U26584 ( .A(n26717), .ZN(n26210) );
  NOR2_X1 U26585 ( .A1(n29560), .A2(n26718), .ZN(n25661) );
  NOR2_X1 U26587 ( .A1(n28548), .A2(n28459), .ZN(n25662) );
  NAND2_X1 U26588 ( .A1(n25662), .A2(n283), .ZN(n25663) );
  NAND3_X1 U26589 ( .A1(n27350), .A2(n29052), .A3(n28549), .ZN(n25672) );
  OR2_X1 U26590 ( .A1(n27340), .A2(n27352), .ZN(n25957) );
  NOR2_X1 U26591 ( .A1(n26186), .A2(n26182), .ZN(n26472) );
  NOR2_X1 U26592 ( .A1(n25666), .A2(n26185), .ZN(n25667) );
  NOR2_X1 U26593 ( .A1(n26472), .A2(n25667), .ZN(n26474) );
  INV_X1 U26594 ( .A(n28561), .ZN(n25668) );
  AOI21_X1 U26595 ( .B1(n26180), .B2(n25668), .A(n28525), .ZN(n25669) );
  INV_X1 U26597 ( .A(n1046), .ZN(n25674) );
  XNOR2_X1 U26598 ( .A(n25675), .B(n25674), .ZN(Ciphertext[5]) );
  NOR2_X1 U26599 ( .A1(n27048), .A2(n28130), .ZN(n25968) );
  INV_X1 U26600 ( .A(n27044), .ZN(n27002) );
  AOI21_X1 U26601 ( .B1(n28783), .B2(n27002), .A(n27048), .ZN(n25677) );
  OR2_X1 U26602 ( .A1(n25677), .A2(n27041), .ZN(n25678) );
  NAND2_X1 U26603 ( .A1(n25679), .A2(n25678), .ZN(n26539) );
  INV_X1 U26604 ( .A(n26539), .ZN(n27865) );
  XNOR2_X1 U26605 ( .A(n26021), .B(n25680), .ZN(n25686) );
  INV_X1 U26606 ( .A(n25681), .ZN(n25682) );
  XNOR2_X1 U26607 ( .A(n363), .B(n25682), .ZN(n25684) );
  XNOR2_X1 U26608 ( .A(n26114), .B(n27298), .ZN(n25683) );
  XNOR2_X1 U26609 ( .A(n25683), .B(n25684), .ZN(n25685) );
  XNOR2_X1 U26610 ( .A(n25685), .B(n25686), .ZN(n26614) );
  XNOR2_X1 U26611 ( .A(n25687), .B(n25688), .ZN(n25693) );
  XNOR2_X1 U26612 ( .A(n25689), .B(n26680), .ZN(n25690) );
  XNOR2_X1 U26613 ( .A(n25691), .B(n25690), .ZN(n25692) );
  XNOR2_X1 U26614 ( .A(n25826), .B(n1133), .ZN(n25695) );
  XNOR2_X1 U26615 ( .A(n25694), .B(n25695), .ZN(n25700) );
  XNOR2_X1 U26616 ( .A(n25697), .B(n25696), .ZN(n25859) );
  XNOR2_X1 U26617 ( .A(n25698), .B(n25859), .ZN(n25699) );
  XNOR2_X1 U26619 ( .A(n25701), .B(n26013), .ZN(n25707) );
  XNOR2_X1 U26620 ( .A(n25702), .B(n29053), .ZN(n25705) );
  XNOR2_X1 U26621 ( .A(n25703), .B(n3196), .ZN(n25704) );
  XNOR2_X1 U26622 ( .A(n25705), .B(n25704), .ZN(n25706) );
  XNOR2_X1 U26623 ( .A(n25775), .B(n25867), .ZN(n25710) );
  XNOR2_X1 U26624 ( .A(n25708), .B(n2912), .ZN(n25709) );
  XNOR2_X1 U26625 ( .A(n25710), .B(n25709), .ZN(n25712) );
  XNOR2_X1 U26626 ( .A(n25714), .B(n26108), .ZN(n25715) );
  XNOR2_X1 U26627 ( .A(n26030), .B(n25715), .ZN(n25719) );
  XNOR2_X1 U26628 ( .A(n25785), .B(n135), .ZN(n25716) );
  XNOR2_X1 U26629 ( .A(n25717), .B(n25716), .ZN(n25718) );
  NOR2_X1 U26631 ( .A1(n27865), .A2(n27877), .ZN(n26594) );
  XNOR2_X1 U26632 ( .A(n25722), .B(n25721), .ZN(n25726) );
  XNOR2_X1 U26633 ( .A(n29563), .B(n3606), .ZN(n25723) );
  XNOR2_X1 U26634 ( .A(n25724), .B(n25723), .ZN(n25725) );
  XNOR2_X1 U26635 ( .A(n25726), .B(n25725), .ZN(n26988) );
  INV_X1 U26636 ( .A(n26988), .ZN(n26991) );
  XNOR2_X1 U26637 ( .A(n25727), .B(n26038), .ZN(n25728) );
  XNOR2_X1 U26638 ( .A(n25900), .B(n440), .ZN(n25731) );
  XNOR2_X1 U26639 ( .A(n25729), .B(n26046), .ZN(n25730) );
  XNOR2_X1 U26640 ( .A(n25730), .B(n25731), .ZN(n25732) );
  XNOR2_X2 U26641 ( .A(n25733), .B(n25732), .ZN(n27074) );
  XNOR2_X1 U26642 ( .A(n25735), .B(n25734), .ZN(n25742) );
  XNOR2_X1 U26643 ( .A(n25737), .B(n29017), .ZN(n25740) );
  XNOR2_X1 U26644 ( .A(n25738), .B(n2505), .ZN(n25739) );
  XNOR2_X1 U26645 ( .A(n25740), .B(n25739), .ZN(n25741) );
  XNOR2_X1 U26647 ( .A(n28593), .B(n25810), .ZN(n25747) );
  XNOR2_X1 U26648 ( .A(n25745), .B(n3662), .ZN(n25746) );
  XNOR2_X1 U26650 ( .A(n26029), .B(n25751), .ZN(n25752) );
  XNOR2_X1 U26651 ( .A(n25752), .B(n25753), .ZN(n25758) );
  XNOR2_X1 U26652 ( .A(n25754), .B(n2510), .ZN(n25755) );
  XNOR2_X1 U26653 ( .A(n25756), .B(n25755), .ZN(n25757) );
  INV_X1 U26654 ( .A(n26322), .ZN(n27077) );
  NOR2_X1 U26655 ( .A1(n27074), .A2(n27077), .ZN(n25768) );
  XNOR2_X1 U26656 ( .A(n29155), .B(n25819), .ZN(n25762) );
  XNOR2_X1 U26657 ( .A(n25760), .B(n25761), .ZN(n26014) );
  XNOR2_X1 U26658 ( .A(n26014), .B(n25762), .ZN(n25766) );
  XNOR2_X1 U26659 ( .A(n25445), .B(n3673), .ZN(n25764) );
  XNOR2_X1 U26660 ( .A(n25763), .B(n25764), .ZN(n25765) );
  NOR2_X1 U26661 ( .A1(n26991), .A2(n26989), .ZN(n25767) );
  INV_X1 U26662 ( .A(n29623), .ZN(n27317) );
  XNOR2_X1 U26663 ( .A(n25772), .B(n25771), .ZN(n25779) );
  XNOR2_X1 U26664 ( .A(n29634), .B(n25773), .ZN(n25777) );
  INV_X1 U26665 ( .A(Key[13]), .ZN(n25774) );
  XNOR2_X1 U26666 ( .A(n25775), .B(n25774), .ZN(n25776) );
  XNOR2_X1 U26667 ( .A(n25777), .B(n25776), .ZN(n25778) );
  XNOR2_X1 U26668 ( .A(n25779), .B(n25778), .ZN(n25815) );
  XNOR2_X1 U26669 ( .A(n25781), .B(n25780), .ZN(n25784) );
  XNOR2_X1 U26670 ( .A(n25782), .B(n1887), .ZN(n25783) );
  XNOR2_X1 U26671 ( .A(n25783), .B(n25784), .ZN(n25789) );
  XNOR2_X1 U26672 ( .A(n25786), .B(n25785), .ZN(n25787) );
  XNOR2_X1 U26673 ( .A(n26034), .B(n25787), .ZN(n25788) );
  XNOR2_X1 U26674 ( .A(n25789), .B(n25788), .ZN(n27018) );
  XNOR2_X1 U26676 ( .A(n25790), .B(n26039), .ZN(n26076) );
  XNOR2_X1 U26677 ( .A(n26076), .B(n25791), .ZN(n25805) );
  INV_X1 U26678 ( .A(n25797), .ZN(n25792) );
  NAND2_X1 U26679 ( .A1(n25792), .A2(n3644), .ZN(n25801) );
  INV_X1 U26680 ( .A(n25793), .ZN(n25796) );
  NOR2_X1 U26681 ( .A1(n25794), .A2(n3644), .ZN(n25795) );
  NAND2_X1 U26682 ( .A1(n25796), .A2(n25795), .ZN(n25799) );
  INV_X1 U26683 ( .A(n3644), .ZN(n26257) );
  NAND2_X1 U26684 ( .A1(n25797), .A2(n26257), .ZN(n25798) );
  OAI211_X1 U26685 ( .C1(n25801), .C2(n25800), .A(n25799), .B(n25798), .ZN(
        n25802) );
  XNOR2_X1 U26686 ( .A(n25803), .B(n25802), .ZN(n25804) );
  MUX2_X1 U26687 ( .A(n25815), .B(n28640), .S(n26841), .Z(n25814) );
  XNOR2_X1 U26688 ( .A(n25806), .B(n25807), .ZN(n25813) );
  XNOR2_X1 U26689 ( .A(n25809), .B(n25808), .ZN(n26116) );
  XNOR2_X1 U26690 ( .A(n25810), .B(n3317), .ZN(n25811) );
  XNOR2_X1 U26691 ( .A(n26116), .B(n25811), .ZN(n25812) );
  NOR2_X1 U26692 ( .A1(n26841), .A2(n27086), .ZN(n25833) );
  XNOR2_X1 U26693 ( .A(n26011), .B(n2541), .ZN(n25818) );
  XNOR2_X1 U26694 ( .A(n25818), .B(n25817), .ZN(n25824) );
  XNOR2_X1 U26695 ( .A(n25820), .B(n25819), .ZN(n25822) );
  XNOR2_X1 U26696 ( .A(n25821), .B(n25822), .ZN(n25823) );
  NOR2_X1 U26697 ( .A1(n26507), .A2(n26840), .ZN(n25832) );
  XNOR2_X1 U26698 ( .A(n25825), .B(n26909), .ZN(n25827) );
  XNOR2_X1 U26699 ( .A(n25826), .B(n25827), .ZN(n25829) );
  XNOR2_X1 U26700 ( .A(n25829), .B(n25828), .ZN(n25831) );
  XNOR2_X1 U26701 ( .A(n25831), .B(n25830), .ZN(n27081) );
  INV_X1 U26702 ( .A(n27081), .ZN(n26842) );
  XNOR2_X1 U26703 ( .A(n26070), .B(n25836), .ZN(n25838) );
  XNOR2_X1 U26704 ( .A(n25838), .B(n25837), .ZN(n25842) );
  XNOR2_X1 U26705 ( .A(n25839), .B(n25840), .ZN(n25841) );
  XNOR2_X1 U26706 ( .A(n25133), .B(n363), .ZN(n25847) );
  XNOR2_X1 U26707 ( .A(n26114), .B(n25845), .ZN(n25846) );
  XNOR2_X1 U26708 ( .A(n25846), .B(n25847), .ZN(n25854) );
  XNOR2_X1 U26709 ( .A(n25849), .B(n25848), .ZN(n25852) );
  XNOR2_X1 U26710 ( .A(n29046), .B(n72), .ZN(n25851) );
  XNOR2_X1 U26711 ( .A(n25852), .B(n25851), .ZN(n25853) );
  NOR2_X1 U26712 ( .A1(n27120), .A2(n26837), .ZN(n26516) );
  XNOR2_X1 U26713 ( .A(n25856), .B(n25857), .ZN(n25862) );
  XNOR2_X1 U26714 ( .A(n25858), .B(n3554), .ZN(n25860) );
  XNOR2_X1 U26715 ( .A(n25859), .B(n25860), .ZN(n25861) );
  XNOR2_X1 U26717 ( .A(n29534), .B(n300), .ZN(n25866) );
  XNOR2_X1 U26718 ( .A(n25864), .B(n25922), .ZN(n25865) );
  XNOR2_X1 U26719 ( .A(n25866), .B(n25865), .ZN(n25873) );
  XNOR2_X1 U26720 ( .A(n25868), .B(n25867), .ZN(n25871) );
  XNOR2_X1 U26721 ( .A(n25869), .B(n27643), .ZN(n25870) );
  XNOR2_X1 U26722 ( .A(n25871), .B(n25870), .ZN(n25872) );
  XNOR2_X1 U26723 ( .A(n25873), .B(n25872), .ZN(n26835) );
  XNOR2_X1 U26724 ( .A(n25875), .B(n25874), .ZN(n25880) );
  XNOR2_X1 U26725 ( .A(n25876), .B(n3386), .ZN(n25878) );
  XNOR2_X1 U26726 ( .A(n25878), .B(n25877), .ZN(n25879) );
  XNOR2_X1 U26727 ( .A(n25880), .B(n25879), .ZN(n27121) );
  NAND2_X1 U26728 ( .A1(n6951), .A2(n27121), .ZN(n25883) );
  NAND2_X1 U26729 ( .A1(n28631), .A2(n28437), .ZN(n25881) );
  INV_X1 U26730 ( .A(n27121), .ZN(n26334) );
  NAND2_X1 U26731 ( .A1(n25881), .A2(n26334), .ZN(n25882) );
  OAI21_X1 U26732 ( .B1(n26516), .B2(n25883), .A(n25882), .ZN(n25896) );
  XNOR2_X1 U26733 ( .A(n25928), .B(n25884), .ZN(n25888) );
  XNOR2_X1 U26734 ( .A(n29073), .B(n25885), .ZN(n25887) );
  XNOR2_X1 U26735 ( .A(n25888), .B(n25887), .ZN(n25895) );
  XNOR2_X1 U26736 ( .A(n25890), .B(n29053), .ZN(n25893) );
  XNOR2_X1 U26737 ( .A(n25891), .B(n2403), .ZN(n25892) );
  XNOR2_X1 U26738 ( .A(n25893), .B(n25892), .ZN(n25894) );
  XNOR2_X1 U26739 ( .A(n25895), .B(n25894), .ZN(n26512) );
  NAND2_X1 U26740 ( .A1(n27118), .A2(n26512), .ZN(n26302) );
  NAND2_X1 U26741 ( .A1(n25896), .A2(n26302), .ZN(n27862) );
  XNOR2_X1 U26742 ( .A(n25898), .B(n25899), .ZN(n25907) );
  XNOR2_X1 U26743 ( .A(n25901), .B(n25900), .ZN(n25905) );
  XNOR2_X1 U26744 ( .A(n25903), .B(n25902), .ZN(n25904) );
  XNOR2_X1 U26745 ( .A(n25905), .B(n25904), .ZN(n25906) );
  XNOR2_X1 U26746 ( .A(n28771), .B(n3219), .ZN(n25912) );
  XNOR2_X1 U26747 ( .A(n25910), .B(n25909), .ZN(n25911) );
  XNOR2_X1 U26748 ( .A(n25912), .B(n25911), .ZN(n25918) );
  XNOR2_X1 U26749 ( .A(n29039), .B(n25914), .ZN(n25916) );
  XNOR2_X1 U26750 ( .A(n25915), .B(n25916), .ZN(n25917) );
  XNOR2_X1 U26751 ( .A(n25920), .B(n25919), .ZN(n25926) );
  XNOR2_X1 U26752 ( .A(n25921), .B(n27462), .ZN(n25924) );
  XNOR2_X1 U26753 ( .A(n25924), .B(n25923), .ZN(n25925) );
  XNOR2_X1 U26754 ( .A(n25926), .B(n25925), .ZN(n26848) );
  XNOR2_X1 U26755 ( .A(n25927), .B(n25928), .ZN(n25930) );
  XNOR2_X1 U26756 ( .A(n25929), .B(n25930), .ZN(n25937) );
  XNOR2_X1 U26757 ( .A(n25932), .B(n25931), .ZN(n25935) );
  XNOR2_X1 U26758 ( .A(n25933), .B(n3650), .ZN(n25934) );
  XNOR2_X1 U26759 ( .A(n25935), .B(n25934), .ZN(n25936) );
  AOI22_X1 U26760 ( .A1(n26510), .A2(n26849), .B1(n26848), .B2(n27056), .ZN(
        n26301) );
  INV_X1 U26761 ( .A(n26850), .ZN(n27898) );
  XNOR2_X1 U26762 ( .A(n25939), .B(n25938), .ZN(n25941) );
  XNOR2_X1 U26763 ( .A(n25943), .B(n25944), .ZN(n25946) );
  XNOR2_X1 U26764 ( .A(n25946), .B(n25945), .ZN(n25952) );
  INV_X1 U26765 ( .A(n2527), .ZN(n27915) );
  XNOR2_X1 U26766 ( .A(n25948), .B(n27915), .ZN(n25949) );
  XNOR2_X1 U26767 ( .A(n25950), .B(n25949), .ZN(n25951) );
  XNOR2_X2 U26768 ( .A(n25952), .B(n25951), .ZN(n27902) );
  OAI21_X1 U26770 ( .B1(n26849), .B2(n29536), .A(n26852), .ZN(n25953) );
  MUX2_X1 U26771 ( .A(n27865), .B(n27872), .S(n27871), .Z(n25954) );
  XNOR2_X1 U26772 ( .A(n25955), .B(n6016), .ZN(Ciphertext[147]) );
  OAI21_X1 U26773 ( .B1(n27358), .B2(n27354), .A(n29052), .ZN(n25956) );
  NAND2_X1 U26774 ( .A1(n27355), .A2(n27354), .ZN(n27330) );
  MUX2_X1 U26775 ( .A(n27357), .B(n25956), .S(n27330), .Z(n25959) );
  NOR2_X1 U26776 ( .A1(n27340), .A2(n27357), .ZN(n27328) );
  NAND2_X1 U26777 ( .A1(n25959), .A2(n25958), .ZN(n25961) );
  INV_X1 U26778 ( .A(n3081), .ZN(n25960) );
  XNOR2_X1 U26779 ( .A(n25961), .B(n25960), .ZN(Ciphertext[4]) );
  NAND2_X1 U26780 ( .A1(n27066), .A2(n25963), .ZN(n25966) );
  NOR2_X1 U26781 ( .A1(n922), .A2(n28452), .ZN(n25964) );
  OR2_X1 U26782 ( .A1(n25964), .A2(n29520), .ZN(n25965) );
  OAI211_X1 U26784 ( .C1(n29524), .C2(n29058), .A(n28130), .B(n398), .ZN(
        n25969) );
  NAND2_X1 U26785 ( .A1(n25970), .A2(n25969), .ZN(n28017) );
  INV_X1 U26786 ( .A(n28017), .ZN(n28001) );
  NOR2_X1 U26787 ( .A1(n29482), .A2(n26733), .ZN(n26734) );
  NOR2_X1 U26788 ( .A1(n26997), .A2(n26998), .ZN(n28099) );
  INV_X1 U26790 ( .A(n26755), .ZN(n26236) );
  OR2_X1 U26791 ( .A1(n29479), .A2(n28575), .ZN(n25973) );
  AOI21_X1 U26792 ( .B1(n25973), .B2(n25603), .A(n26753), .ZN(n25974) );
  NOR2_X1 U26794 ( .A1(n29099), .A2(n26748), .ZN(n25977) );
  NOR2_X1 U26795 ( .A1(n5035), .A2(n25977), .ZN(n25982) );
  INV_X1 U26796 ( .A(n26747), .ZN(n26223) );
  AOI21_X1 U26797 ( .B1(n26223), .B2(n29159), .A(n26222), .ZN(n25981) );
  AOI22_X1 U26798 ( .A1(n26222), .A2(n25979), .B1(n25453), .B2(n25978), .ZN(
        n25980) );
  OAI21_X1 U26799 ( .B1(n25982), .B2(n25981), .A(n25980), .ZN(n28021) );
  NOR2_X1 U26800 ( .A1(n26984), .A2(n28021), .ZN(n27034) );
  MUX2_X1 U26801 ( .A(n27014), .B(n26623), .S(n29062), .Z(n25986) );
  INV_X1 U26802 ( .A(n29062), .ZN(n25983) );
  INV_X1 U26803 ( .A(n27010), .ZN(n27053) );
  NOR2_X1 U26804 ( .A1(n28446), .A2(n27053), .ZN(n25984) );
  NOR2_X1 U26805 ( .A1(n27017), .A2(n25984), .ZN(n25985) );
  NAND2_X1 U26806 ( .A1(n27034), .A2(n28019), .ZN(n25989) );
  NOR2_X1 U26807 ( .A1(n28019), .A2(n28411), .ZN(n25987) );
  NAND2_X1 U26808 ( .A1(n25987), .A2(n28003), .ZN(n25988) );
  NAND3_X1 U26809 ( .A1(n25990), .A2(n25989), .A3(n25988), .ZN(n25993) );
  XNOR2_X1 U26810 ( .A(n25993), .B(n25992), .ZN(Ciphertext[170]) );
  INV_X1 U26811 ( .A(n27371), .ZN(n26497) );
  INV_X1 U26812 ( .A(n26808), .ZN(n25994) );
  XNOR2_X1 U26813 ( .A(n25996), .B(n857), .ZN(Ciphertext[7]) );
  NOR2_X1 U26814 ( .A1(n29538), .A2(n28562), .ZN(n25999) );
  NOR2_X1 U26815 ( .A1(n25994), .A2(n27371), .ZN(n27365) );
  AOI22_X1 U26816 ( .A1(n25999), .A2(n27362), .B1(n27365), .B2(n27368), .ZN(
        n26001) );
  NAND2_X1 U26817 ( .A1(n27366), .A2(n27368), .ZN(n26000) );
  INV_X1 U26818 ( .A(n3622), .ZN(n26003) );
  XNOR2_X1 U26819 ( .A(n26004), .B(n26214), .ZN(n26005) );
  XNOR2_X1 U26820 ( .A(n26006), .B(n26005), .ZN(n26010) );
  INV_X1 U26821 ( .A(n27155), .ZN(n26018) );
  XNOR2_X1 U26822 ( .A(n26011), .B(n4029), .ZN(n26012) );
  XNOR2_X1 U26823 ( .A(n26013), .B(n26012), .ZN(n26017) );
  XNOR2_X1 U26824 ( .A(n26014), .B(n26015), .ZN(n26016) );
  XNOR2_X1 U26825 ( .A(n26016), .B(n26017), .ZN(n26867) );
  INV_X1 U26826 ( .A(n26867), .ZN(n27153) );
  NOR2_X1 U26827 ( .A1(n26018), .A2(n27153), .ZN(n26052) );
  XNOR2_X1 U26828 ( .A(n26020), .B(n26019), .ZN(n26022) );
  XNOR2_X1 U26829 ( .A(n26021), .B(n26022), .ZN(n26027) );
  XNOR2_X1 U26830 ( .A(n26023), .B(n27452), .ZN(n26024) );
  XNOR2_X1 U26831 ( .A(n26025), .B(n26024), .ZN(n26026) );
  XNOR2_X1 U26832 ( .A(n28534), .B(n26029), .ZN(n26031) );
  XNOR2_X1 U26833 ( .A(n26030), .B(n26031), .ZN(n26037) );
  XNOR2_X1 U26834 ( .A(n25386), .B(n26032), .ZN(n26035) );
  XNOR2_X1 U26835 ( .A(n26034), .B(n26035), .ZN(n26036) );
  XNOR2_X1 U26836 ( .A(n26037), .B(n26036), .ZN(n26868) );
  XNOR2_X1 U26838 ( .A(n26039), .B(n26038), .ZN(n26043) );
  XNOR2_X1 U26839 ( .A(n26041), .B(n26040), .ZN(n26042) );
  XNOR2_X1 U26841 ( .A(n28475), .B(n3003), .ZN(n26048) );
  XNOR2_X1 U26842 ( .A(n26046), .B(n26045), .ZN(n26047) );
  XNOR2_X1 U26843 ( .A(n26047), .B(n26048), .ZN(n26049) );
  XNOR2_X1 U26845 ( .A(n26054), .B(n26053), .ZN(n26058) );
  XNOR2_X1 U26846 ( .A(n29613), .B(n26055), .ZN(n26057) );
  XNOR2_X1 U26847 ( .A(n26057), .B(n26058), .ZN(n26064) );
  XNOR2_X1 U26848 ( .A(n26084), .B(n26059), .ZN(n26062) );
  XNOR2_X1 U26849 ( .A(n26060), .B(n2889), .ZN(n26061) );
  XNOR2_X1 U26850 ( .A(n26062), .B(n26061), .ZN(n26063) );
  NOR2_X1 U26852 ( .A1(n29474), .A2(n29048), .ZN(n26066) );
  NOR2_X1 U26856 ( .A1(n26067), .A2(n26867), .ZN(n26068) );
  INV_X1 U26857 ( .A(n27728), .ZN(n26126) );
  XNOR2_X1 U26858 ( .A(n26071), .B(n26070), .ZN(n26075) );
  INV_X1 U26859 ( .A(n28693), .ZN(n26072) );
  XNOR2_X1 U26860 ( .A(n29129), .B(n26072), .ZN(n26074) );
  XNOR2_X1 U26861 ( .A(n26075), .B(n26074), .ZN(n26079) );
  XNOR2_X1 U26862 ( .A(n26080), .B(n3482), .ZN(n26082) );
  XNOR2_X1 U26863 ( .A(n26082), .B(n26081), .ZN(n26088) );
  XNOR2_X1 U26864 ( .A(n26084), .B(n26083), .ZN(n26085) );
  XNOR2_X1 U26865 ( .A(n26086), .B(n26085), .ZN(n26087) );
  XNOR2_X1 U26866 ( .A(n300), .B(n26089), .ZN(n26092) );
  XNOR2_X1 U26867 ( .A(n26091), .B(n26092), .ZN(n26099) );
  XNOR2_X1 U26868 ( .A(n26094), .B(n26093), .ZN(n26097) );
  INV_X1 U26869 ( .A(n2385), .ZN(n27887) );
  XNOR2_X1 U26870 ( .A(n26095), .B(n27887), .ZN(n26096) );
  XNOR2_X1 U26871 ( .A(n26097), .B(n26096), .ZN(n26098) );
  INV_X1 U26872 ( .A(n27137), .ZN(n26858) );
  XNOR2_X1 U26874 ( .A(n26105), .B(n26104), .ZN(n26518) );
  XNOR2_X1 U26875 ( .A(n1871), .B(n26108), .ZN(n26112) );
  XNOR2_X1 U26876 ( .A(n26110), .B(n27788), .ZN(n26111) );
  XNOR2_X1 U26877 ( .A(n26112), .B(n26111), .ZN(n26113) );
  XNOR2_X1 U26878 ( .A(n26114), .B(n26115), .ZN(n26117) );
  XNOR2_X1 U26879 ( .A(n26117), .B(n26116), .ZN(n26124) );
  XNOR2_X1 U26880 ( .A(n29543), .B(n26118), .ZN(n26122) );
  INV_X1 U26881 ( .A(n2465), .ZN(n28050) );
  XNOR2_X1 U26882 ( .A(n26120), .B(n28050), .ZN(n26121) );
  XNOR2_X1 U26883 ( .A(n26122), .B(n26121), .ZN(n26123) );
  INV_X1 U26885 ( .A(n26518), .ZN(n27142) );
  NOR2_X1 U26886 ( .A1(n26350), .A2(n27704), .ZN(n26127) );
  NOR2_X1 U26888 ( .A1(n27691), .A2(n27707), .ZN(n27727) );
  NAND2_X1 U26889 ( .A1(n6953), .A2(n27727), .ZN(n26148) );
  INV_X1 U26890 ( .A(n27178), .ZN(n27129) );
  NOR2_X1 U26891 ( .A1(n27175), .A2(n28536), .ZN(n26130) );
  OAI21_X1 U26892 ( .B1(n26130), .B2(n28392), .A(n27178), .ZN(n26131) );
  INV_X1 U26893 ( .A(n26386), .ZN(n26132) );
  NOR2_X1 U26894 ( .A1(n26260), .A2(n26133), .ZN(n26137) );
  AND2_X1 U26896 ( .A1(n26384), .A2(n1907), .ZN(n26135) );
  OAI21_X1 U26897 ( .B1(n27171), .B2(n26135), .A(n28535), .ZN(n26136) );
  NAND2_X1 U26899 ( .A1(n27193), .A2(n28595), .ZN(n26139) );
  MUX2_X1 U26900 ( .A(n26139), .B(n26138), .S(n27123), .Z(n26144) );
  NOR3_X1 U26901 ( .A1(n27193), .A2(n4109), .A3(n27124), .ZN(n26142) );
  NOR2_X1 U26902 ( .A1(n26140), .A2(n28595), .ZN(n26141) );
  NOR2_X1 U26906 ( .A1(n26576), .A2(n26789), .ZN(n26924) );
  NAND2_X1 U26907 ( .A1(n26924), .A2(n26791), .ZN(n26154) );
  INV_X1 U26911 ( .A(n26458), .ZN(n26461) );
  NOR2_X1 U26912 ( .A1(n26461), .A2(n28578), .ZN(n26562) );
  NAND2_X1 U26913 ( .A1(n28578), .A2(n26457), .ZN(n26157) );
  NAND3_X1 U26914 ( .A1(n26157), .A2(n26560), .A3(n28434), .ZN(n26158) );
  INV_X1 U26916 ( .A(n27460), .ZN(n27467) );
  INV_X1 U26917 ( .A(n26455), .ZN(n26161) );
  INV_X1 U26919 ( .A(n26454), .ZN(n26177) );
  NOR2_X1 U26920 ( .A1(n29105), .A2(n26454), .ZN(n26163) );
  OAI21_X1 U26921 ( .B1(n26163), .B2(n26162), .A(n29467), .ZN(n26164) );
  OAI21_X1 U26922 ( .B1(n27465), .B2(n27467), .A(n29468), .ZN(n26170) );
  AND2_X1 U26923 ( .A1(n28435), .A2(n27463), .ZN(n27236) );
  INV_X1 U26924 ( .A(n26914), .ZN(n26568) );
  MUX2_X1 U26925 ( .A(n29610), .B(n26568), .S(n26567), .Z(n26169) );
  NOR2_X1 U26926 ( .A1(n5625), .A2(n26786), .ZN(n26168) );
  INV_X1 U26927 ( .A(n27457), .ZN(n27235) );
  AOI22_X1 U26928 ( .A1(n26170), .A2(n27458), .B1(n27236), .B2(n27235), .ZN(
        n26175) );
  NAND2_X1 U26929 ( .A1(n26920), .A2(n4820), .ZN(n26171) );
  INV_X1 U26930 ( .A(n26782), .ZN(n26174) );
  NOR2_X1 U26931 ( .A1(n27457), .A2(n27447), .ZN(n26606) );
  NOR2_X1 U26932 ( .A1(n26180), .A2(n26476), .ZN(n26184) );
  NOR2_X1 U26933 ( .A1(n26181), .A2(n28503), .ZN(n26183) );
  MUX2_X1 U26934 ( .A(n26184), .B(n26183), .S(n28547), .Z(n26190) );
  NAND3_X1 U26936 ( .A1(n28561), .A2(n28503), .A3(n28525), .ZN(n26187) );
  OAI21_X1 U26937 ( .B1(n29596), .B2(n26475), .A(n26187), .ZN(n26189) );
  NAND2_X1 U26938 ( .A1(n26464), .A2(n26191), .ZN(n26193) );
  AOI21_X1 U26939 ( .B1(n26193), .B2(n26192), .A(n27395), .ZN(n26197) );
  AND3_X1 U26940 ( .A1(n28908), .A2(n280), .A3(n26469), .ZN(n26196) );
  MUX2_X1 U26941 ( .A(n28560), .B(n26728), .S(n26729), .Z(n26198) );
  NAND2_X1 U26942 ( .A1(n26198), .A2(n1622), .ZN(n26199) );
  NAND3_X1 U26943 ( .A1(n26200), .A2(n26204), .A3(n26737), .ZN(n26207) );
  NOR2_X1 U26944 ( .A1(n26204), .A2(n26235), .ZN(n26201) );
  NAND2_X1 U26945 ( .A1(n26201), .A2(n1874), .ZN(n26206) );
  NAND2_X1 U26946 ( .A1(n28473), .A2(n1874), .ZN(n26234) );
  NAND3_X1 U26947 ( .A1(n26204), .A2(n26203), .A3(n26740), .ZN(n26205) );
  AND4_X1 U26948 ( .A1(n26207), .A2(n26206), .A3(n26234), .A4(n26205), .ZN(
        n27379) );
  INV_X1 U26949 ( .A(n26217), .ZN(n26213) );
  AND2_X1 U26950 ( .A1(n26715), .A2(n26718), .ZN(n26216) );
  NAND2_X1 U26951 ( .A1(n26216), .A2(n26208), .ZN(n26212) );
  AOI21_X1 U26953 ( .B1(n283), .B2(n28459), .A(n26215), .ZN(n26219) );
  NOR2_X1 U26955 ( .A1(n26222), .A2(n5760), .ZN(n26221) );
  AOI21_X1 U26956 ( .B1(n26223), .B2(n26222), .A(n26221), .ZN(n26226) );
  INV_X1 U26957 ( .A(n29100), .ZN(n26224) );
  INV_X1 U26959 ( .A(n28069), .ZN(n26227) );
  NAND2_X1 U26960 ( .A1(n26231), .A2(n26234), .ZN(n26232) );
  NAND2_X1 U26961 ( .A1(n26236), .A2(n26757), .ZN(n26239) );
  MUX2_X1 U26962 ( .A(n26239), .B(n26238), .S(n26753), .Z(n26244) );
  AND2_X1 U26963 ( .A1(n28575), .A2(n26240), .ZN(n26758) );
  AOI22_X1 U26964 ( .A1(n26242), .A2(n26761), .B1(n26758), .B2(n26241), .ZN(
        n26243) );
  INV_X1 U26965 ( .A(n27014), .ZN(n27049) );
  NAND2_X1 U26966 ( .A1(n29062), .A2(n27049), .ZN(n26245) );
  NAND2_X1 U26967 ( .A1(n26246), .A2(n26245), .ZN(n26249) );
  OAI21_X1 U26968 ( .B1(n27053), .B2(n399), .A(n28639), .ZN(n26248) );
  NOR2_X1 U26969 ( .A1(n27010), .A2(n27050), .ZN(n26247) );
  NOR3_X1 U26970 ( .A1(n28543), .A2(n28065), .A3(n28063), .ZN(n26250) );
  AOI21_X1 U26971 ( .B1(n28055), .B2(n28067), .A(n26250), .ZN(n26256) );
  NAND2_X1 U26972 ( .A1(n26632), .A2(n26998), .ZN(n26251) );
  OAI21_X1 U26973 ( .B1(n29481), .B2(n5389), .A(n28099), .ZN(n26252) );
  INV_X1 U26974 ( .A(n28066), .ZN(n28044) );
  OAI21_X1 U26975 ( .B1(n28044), .B2(n28063), .A(n28069), .ZN(n26254) );
  NOR2_X1 U26976 ( .A1(n28543), .A2(n28066), .ZN(n28053) );
  NAND2_X1 U26977 ( .A1(n26256), .A2(n26255), .ZN(n26258) );
  XNOR2_X1 U26978 ( .A(n26258), .B(n26257), .ZN(Ciphertext[183]) );
  NOR2_X1 U26979 ( .A1(n28535), .A2(n28572), .ZN(n26261) );
  INV_X1 U26980 ( .A(n27165), .ZN(n27168) );
  INV_X1 U26981 ( .A(n26129), .ZN(n27131) );
  MUX2_X1 U26982 ( .A(n29071), .B(n26950), .S(n26949), .Z(n26269) );
  MUX2_X1 U26983 ( .A(n26267), .B(n26948), .S(n26952), .Z(n26268) );
  AOI21_X1 U26985 ( .B1(n1901), .B2(n27585), .A(n28179), .ZN(n26286) );
  OAI21_X1 U26986 ( .B1(n28650), .B2(n27183), .A(n26270), .ZN(n26271) );
  NAND2_X1 U26987 ( .A1(n26271), .A2(n26397), .ZN(n26274) );
  AND3_X1 U26988 ( .A1(n28651), .A2(n27181), .A3(n25124), .ZN(n26272) );
  AOI21_X1 U26989 ( .B1(n28652), .B2(n26357), .A(n26272), .ZN(n26273) );
  MUX2_X2 U26990 ( .A(n26277), .B(n26276), .S(n26361), .Z(n27596) );
  NAND2_X1 U26991 ( .A1(n26798), .A2(n26362), .ZN(n26804) );
  INV_X1 U26992 ( .A(n26392), .ZN(n26279) );
  AOI22_X1 U26994 ( .A1(n26279), .A2(n28470), .B1(n26800), .B2(n29573), .ZN(
        n26282) );
  OR3_X1 U26995 ( .A1(n26798), .A2(n26280), .A3(n26799), .ZN(n26281) );
  OAI211_X1 U26996 ( .C1(n29573), .C2(n26804), .A(n26282), .B(n26281), .ZN(
        n27590) );
  INV_X1 U26997 ( .A(n27590), .ZN(n26284) );
  NOR2_X1 U26998 ( .A1(n26284), .A2(n27586), .ZN(n26285) );
  INV_X1 U26999 ( .A(n2598), .ZN(n26288) );
  MUX2_X1 U27000 ( .A(n28487), .B(n29621), .S(n27137), .Z(n26289) );
  AND2_X1 U27001 ( .A1(n29621), .A2(n27141), .ZN(n26326) );
  INV_X1 U27002 ( .A(n26290), .ZN(n26291) );
  INV_X1 U27003 ( .A(n26292), .ZN(n26293) );
  NOR2_X1 U27004 ( .A1(n29070), .A2(n27768), .ZN(n27782) );
  NAND2_X1 U27005 ( .A1(n27700), .A2(n27702), .ZN(n26297) );
  NAND2_X1 U27006 ( .A1(n26350), .A2(n27704), .ZN(n26296) );
  INV_X1 U27007 ( .A(n27161), .ZN(n26352) );
  OAI21_X1 U27008 ( .B1(n400), .B2(n26352), .A(n455), .ZN(n26295) );
  NOR2_X1 U27009 ( .A1(n27782), .A2(n26298), .ZN(n26315) );
  AOI21_X1 U27011 ( .B1(n27902), .B2(n26848), .A(n28600), .ZN(n26300) );
  NAND2_X1 U27012 ( .A1(n26315), .A2(n29537), .ZN(n26313) );
  INV_X1 U27013 ( .A(n26302), .ZN(n26305) );
  INV_X1 U27014 ( .A(n27120), .ZN(n26303) );
  NOR2_X1 U27015 ( .A1(n26303), .A2(n27121), .ZN(n26304) );
  MUX2_X1 U27016 ( .A(n26305), .B(n26304), .S(n26837), .Z(n26308) );
  INV_X1 U27017 ( .A(n26512), .ZN(n27117) );
  MUX2_X1 U27018 ( .A(n28631), .B(n402), .S(n27117), .Z(n26306) );
  NOR2_X1 U27019 ( .A1(n26306), .A2(n29016), .ZN(n26307) );
  NOR2_X1 U27020 ( .A1(n26308), .A2(n26307), .ZN(n27762) );
  INV_X1 U27021 ( .A(n27111), .ZN(n27154) );
  AOI21_X1 U27022 ( .B1(n27110), .B2(n27154), .A(n26865), .ZN(n26311) );
  NOR2_X1 U27023 ( .A1(n27762), .A2(n27777), .ZN(n27771) );
  OAI21_X1 U27025 ( .B1(n26317), .B2(n2441), .A(n26316), .ZN(n26318) );
  NOR2_X1 U27026 ( .A1(n26319), .A2(n26318), .ZN(Ciphertext[122]) );
  INV_X1 U27027 ( .A(n27074), .ZN(n26321) );
  INV_X1 U27028 ( .A(n26989), .ZN(n26320) );
  MUX2_X1 U27029 ( .A(n26989), .B(n26323), .S(n27074), .Z(n26324) );
  INV_X1 U27031 ( .A(n27140), .ZN(n26855) );
  NOR2_X1 U27032 ( .A1(n29621), .A2(n27137), .ZN(n26325) );
  NAND2_X1 U27033 ( .A1(n27136), .A2(n26326), .ZN(n26327) );
  NOR2_X1 U27034 ( .A1(n29232), .A2(n27807), .ZN(n26339) );
  INV_X1 U27035 ( .A(n27902), .ZN(n27836) );
  AND2_X1 U27036 ( .A1(n27902), .A2(n27898), .ZN(n26511) );
  AOI21_X1 U27037 ( .B1(n26510), .B2(n27836), .A(n26511), .ZN(n26329) );
  NOR2_X1 U27038 ( .A1(n29497), .A2(n26848), .ZN(n26328) );
  NOR2_X1 U27042 ( .A1(n27155), .A2(n26867), .ZN(n27151) );
  NAND2_X1 U27043 ( .A1(n27154), .A2(n27155), .ZN(n27109) );
  NOR2_X1 U27044 ( .A1(n29060), .A2(n26865), .ZN(n26332) );
  INV_X1 U27046 ( .A(n27118), .ZN(n26836) );
  AND2_X1 U27047 ( .A1(n26837), .A2(n27117), .ZN(n26333) );
  NAND2_X1 U27048 ( .A1(n26516), .A2(n26334), .ZN(n26335) );
  AOI22_X1 U27049 ( .A1(n26339), .A2(n27800), .B1(n27819), .B2(n27812), .ZN(
        n26341) );
  OAI21_X1 U27051 ( .B1(n27795), .B2(n29469), .A(n27818), .ZN(n26338) );
  INV_X1 U27052 ( .A(n27807), .ZN(n27821) );
  INV_X1 U27053 ( .A(n27791), .ZN(n26344) );
  NAND2_X1 U27054 ( .A1(n27800), .A2(n28403), .ZN(n26343) );
  AND2_X1 U27055 ( .A1(n27819), .A2(n27818), .ZN(n26342) );
  AOI22_X1 U27056 ( .A1(n27823), .A2(n26344), .B1(n26343), .B2(n26342), .ZN(
        n26345) );
  XNOR2_X1 U27057 ( .A(n26345), .B(n3673), .ZN(Ciphertext[127]) );
  MUX2_X1 U27058 ( .A(n27597), .B(n26346), .S(n27596), .Z(n26348) );
  NOR2_X1 U27059 ( .A1(n27582), .A2(n27594), .ZN(n27265) );
  AND2_X1 U27060 ( .A1(n27582), .A2(n27590), .ZN(n27593) );
  NOR2_X1 U27061 ( .A1(n27265), .A2(n27593), .ZN(n26347) );
  XNOR2_X1 U27063 ( .A(n26349), .B(n1079), .ZN(Ciphertext[86]) );
  NAND2_X1 U27066 ( .A1(n26397), .A2(n27181), .ZN(n26401) );
  NAND2_X1 U27067 ( .A1(n26357), .A2(n26356), .ZN(n27188) );
  MUX2_X1 U27069 ( .A(n27183), .B(n25124), .S(n27181), .Z(n26359) );
  INV_X1 U27070 ( .A(n28650), .ZN(n26358) );
  INV_X1 U27071 ( .A(n27630), .ZN(n27619) );
  AND2_X1 U27072 ( .A1(n26427), .A2(n26381), .ZN(n26432) );
  MUX2_X1 U27073 ( .A(n26798), .B(n26362), .S(n26799), .Z(n26365) );
  OR2_X1 U27075 ( .A1(n26799), .A2(n26280), .ZN(n26363) );
  OAI22_X1 U27076 ( .A1(n27626), .A2(n27619), .B1(n27627), .B2(n27632), .ZN(
        n27610) );
  NAND2_X1 U27077 ( .A1(n27175), .A2(n27177), .ZN(n27134) );
  NAND2_X1 U27078 ( .A1(n27129), .A2(n29132), .ZN(n26366) );
  AOI21_X1 U27080 ( .B1(n27165), .B2(n26384), .A(n28572), .ZN(n26367) );
  INV_X1 U27081 ( .A(n26367), .ZN(n26369) );
  NOR2_X1 U27082 ( .A1(n26385), .A2(n27168), .ZN(n26368) );
  INV_X1 U27083 ( .A(n27625), .ZN(n27613) );
  OAI21_X1 U27084 ( .B1(n27627), .B2(n27613), .A(n3366), .ZN(n26370) );
  AOI22_X1 U27085 ( .A1(n27610), .A2(n27628), .B1(n26370), .B2(n27619), .ZN(
        n26371) );
  XNOR2_X1 U27086 ( .A(n26371), .B(n3232), .ZN(Ciphertext[95]) );
  NOR2_X1 U27087 ( .A1(n28646), .A2(n26775), .ZN(n26373) );
  AOI21_X1 U27088 ( .B1(n26949), .B2(n26440), .A(n26952), .ZN(n26372) );
  INV_X1 U27090 ( .A(n27571), .ZN(n27552) );
  NAND2_X1 U27091 ( .A1(n26935), .A2(n26936), .ZN(n26376) );
  AOI21_X1 U27092 ( .B1(n26772), .B2(n26376), .A(n26943), .ZN(n26377) );
  MUX2_X1 U27093 ( .A(n26382), .B(n26426), .S(n26378), .Z(n26379) );
  OAI21_X1 U27095 ( .B1(n28573), .B2(n27165), .A(n27166), .ZN(n26390) );
  OAI21_X1 U27096 ( .B1(n26387), .B2(n1907), .A(n26385), .ZN(n26389) );
  AOI22_X2 U27097 ( .A1(n27169), .A2(n26390), .B1(n26389), .B2(n28573), .ZN(
        n27562) );
  OAI21_X1 U27098 ( .B1(n28470), .B2(n26797), .A(n29573), .ZN(n26410) );
  NAND2_X1 U27099 ( .A1(n26392), .A2(n26799), .ZN(n26394) );
  NOR2_X1 U27100 ( .A1(n26800), .A2(n29573), .ZN(n26413) );
  MUX2_X1 U27101 ( .A(n26394), .B(n26280), .S(n26413), .Z(n26395) );
  AOI21_X1 U27102 ( .B1(n28651), .B2(n26396), .A(n25124), .ZN(n26402) );
  NAND3_X1 U27103 ( .A1(n26397), .A2(n28650), .A3(n27182), .ZN(n26398) );
  OAI21_X1 U27104 ( .B1(n26399), .B2(n25034), .A(n26398), .ZN(n26400) );
  NAND2_X1 U27105 ( .A1(n27561), .A2(n27562), .ZN(n27567) );
  NAND2_X1 U27106 ( .A1(n27572), .A2(n27567), .ZN(n26403) );
  OAI21_X1 U27107 ( .B1(n27149), .B2(n29085), .A(n26403), .ZN(n26404) );
  XNOR2_X1 U27109 ( .A(n26406), .B(n1062), .ZN(Ciphertext[80]) );
  NAND2_X1 U27110 ( .A1(n28035), .A2(n28038), .ZN(n28037) );
  NOR2_X1 U27111 ( .A1(n29161), .A2(n29032), .ZN(n28028) );
  INV_X1 U27112 ( .A(n28028), .ZN(n26408) );
  INV_X1 U27113 ( .A(n3372), .ZN(n26409) );
  INV_X1 U27114 ( .A(n26410), .ZN(n26414) );
  AND2_X1 U27115 ( .A1(n26280), .A2(n29330), .ZN(n26412) );
  NOR3_X1 U27116 ( .A1(n26414), .A2(n26413), .A3(n26412), .ZN(n26417) );
  MUX2_X1 U27117 ( .A(n26799), .B(n26798), .S(n26797), .Z(n26415) );
  NOR2_X1 U27118 ( .A1(n26415), .A2(n26800), .ZN(n26416) );
  NAND2_X1 U27120 ( .A1(n26565), .A2(n26420), .ZN(n26418) );
  OAI21_X1 U27121 ( .B1(n29610), .B2(n1872), .A(n26418), .ZN(n26419) );
  NOR2_X1 U27122 ( .A1(n26419), .A2(n26914), .ZN(n27305) );
  NOR2_X1 U27123 ( .A1(n26565), .A2(n26911), .ZN(n26421) );
  NOR2_X2 U27124 ( .A1(n27305), .A2(n27304), .ZN(n27308) );
  INV_X1 U27125 ( .A(n26920), .ZN(n26422) );
  OAI21_X1 U27126 ( .B1(n26172), .B2(n26919), .A(n26422), .ZN(n26424) );
  NAND2_X1 U27127 ( .A1(n26782), .A2(n454), .ZN(n26423) );
  MUX2_X1 U27128 ( .A(n26424), .B(n26423), .S(n4820), .Z(n27302) );
  NAND2_X1 U27129 ( .A1(n26917), .A2(n26919), .ZN(n27303) );
  NAND2_X1 U27130 ( .A1(n27302), .A2(n27303), .ZN(n26879) );
  NAND2_X1 U27132 ( .A1(n26430), .A2(n26429), .ZN(n26434) );
  NAND2_X1 U27133 ( .A1(n26432), .A2(n4679), .ZN(n26433) );
  INV_X1 U27134 ( .A(n26936), .ZN(n26435) );
  NAND3_X1 U27135 ( .A1(n28541), .A2(n26943), .A3(n26768), .ZN(n26437) );
  OAI22_X1 U27136 ( .A1(n27308), .A2(n28510), .B1(n29493), .B2(n27301), .ZN(
        n26887) );
  INV_X1 U27137 ( .A(n26952), .ZN(n26439) );
  MUX2_X1 U27138 ( .A(n26439), .B(n26440), .S(n28542), .Z(n26444) );
  NAND2_X1 U27139 ( .A1(n28646), .A2(n26439), .ZN(n26441) );
  MUX2_X1 U27140 ( .A(n26442), .B(n26441), .S(n26440), .Z(n26443) );
  XNOR2_X1 U27144 ( .A(n26446), .B(n3386), .ZN(Ciphertext[71]) );
  NAND2_X1 U27145 ( .A1(n29105), .A2(n26451), .ZN(n26453) );
  NOR2_X1 U27146 ( .A1(n28385), .A2(n26457), .ZN(n26460) );
  NAND2_X1 U27147 ( .A1(n26464), .A2(n26466), .ZN(n26465) );
  OAI21_X1 U27148 ( .B1(n28908), .B2(n280), .A(n26465), .ZN(n26468) );
  INV_X1 U27149 ( .A(n26468), .ZN(n26470) );
  MUX2_X2 U27150 ( .A(n26471), .B(n26470), .S(n26469), .Z(n27429) );
  MUX2_X1 U27151 ( .A(n29542), .B(n27426), .S(n27429), .Z(n26494) );
  NOR2_X1 U27152 ( .A1(n26472), .A2(n28503), .ZN(n26473) );
  NOR2_X1 U27153 ( .A1(n26474), .A2(n26473), .ZN(n26479) );
  AND3_X1 U27154 ( .A1(n28561), .A2(n26477), .A3(n26475), .ZN(n26478) );
  NOR2_X2 U27155 ( .A1(n26479), .A2(n26478), .ZN(n27428) );
  NAND3_X1 U27156 ( .A1(n26482), .A2(n28560), .A3(n26480), .ZN(n26488) );
  NOR2_X1 U27157 ( .A1(n26482), .A2(n26727), .ZN(n26483) );
  NOR2_X1 U27158 ( .A1(n26927), .A2(n25364), .ZN(n26582) );
  NOR2_X1 U27159 ( .A1(n26489), .A2(n26933), .ZN(n26490) );
  NOR2_X1 U27160 ( .A1(n26582), .A2(n26490), .ZN(n26493) );
  OAI21_X1 U27161 ( .B1(n26928), .B2(n26933), .A(n26927), .ZN(n26492) );
  NOR2_X1 U27162 ( .A1(n28477), .A2(n26933), .ZN(n26491) );
  OAI22_X2 U27163 ( .A1(n26493), .A2(n26581), .B1(n26492), .B2(n26491), .ZN(
        n27425) );
  XNOR2_X1 U27164 ( .A(n26495), .B(n3191), .ZN(Ciphertext[26]) );
  NOR2_X1 U27165 ( .A1(n27366), .A2(n29541), .ZN(n26498) );
  NAND2_X1 U27168 ( .A1(n29075), .A2(n27063), .ZN(n26501) );
  INV_X1 U27169 ( .A(n27088), .ZN(n26506) );
  NOR2_X1 U27171 ( .A1(n28458), .A2(n27085), .ZN(n26504) );
  NOR2_X1 U27172 ( .A1(n27086), .A2(n26840), .ZN(n26503) );
  NOR2_X1 U27173 ( .A1(n26504), .A2(n26503), .ZN(n26505) );
  NOR2_X1 U27174 ( .A1(n26841), .A2(n28640), .ZN(n26509) );
  AND2_X1 U27175 ( .A1(n27085), .A2(n26840), .ZN(n26508) );
  NOR3_X1 U27176 ( .A1(n27852), .A2(n26638), .A3(n26639), .ZN(n27849) );
  NAND2_X1 U27178 ( .A1(n27849), .A2(n447), .ZN(n26525) );
  NOR2_X1 U27179 ( .A1(n402), .A2(n28631), .ZN(n26513) );
  OAI21_X1 U27180 ( .B1(n26334), .B2(n28437), .A(n26513), .ZN(n26515) );
  NOR2_X1 U27181 ( .A1(n27136), .A2(n29621), .ZN(n26857) );
  AND2_X1 U27182 ( .A1(n27137), .A2(n27141), .ZN(n26517) );
  OAI21_X1 U27183 ( .B1(n26857), .B2(n26517), .A(n27147), .ZN(n26521) );
  OAI21_X1 U27184 ( .B1(n26519), .B2(n27138), .A(n27139), .ZN(n26520) );
  INV_X1 U27185 ( .A(n26641), .ZN(n27851) );
  AOI21_X1 U27186 ( .B1(n27855), .B2(n27851), .A(n27847), .ZN(n26522) );
  OAI21_X1 U27187 ( .B1(n27855), .B2(n5295), .A(n26522), .ZN(n26524) );
  NAND2_X1 U27188 ( .A1(n27855), .A2(n6907), .ZN(n26523) );
  INV_X1 U27189 ( .A(n27425), .ZN(n27418) );
  INV_X1 U27192 ( .A(n26669), .ZN(n26529) );
  INV_X1 U27193 ( .A(n26531), .ZN(n26528) );
  INV_X1 U27194 ( .A(n27426), .ZN(n26668) );
  AND2_X1 U27195 ( .A1(n27424), .A2(n27428), .ZN(n26530) );
  OAI21_X1 U27196 ( .B1(n26668), .B2(n27425), .A(n26530), .ZN(n26532) );
  AND3_X1 U27197 ( .A1(n26529), .A2(n26528), .A3(n26532), .ZN(n26536) );
  NAND2_X1 U27198 ( .A1(n27429), .A2(n27425), .ZN(n27417) );
  OAI21_X1 U27202 ( .B1(n27875), .B2(n27866), .A(n3378), .ZN(n26538) );
  INV_X1 U27203 ( .A(n26538), .ZN(n26543) );
  INV_X1 U27205 ( .A(n27864), .ZN(n26540) );
  NAND3_X1 U27206 ( .A1(n27875), .A2(n27872), .A3(n26540), .ZN(n26542) );
  NAND3_X1 U27207 ( .A1(n27872), .A2(n27873), .A3(n27864), .ZN(n26541) );
  NAND4_X1 U27208 ( .A1(n26544), .A2(n26543), .A3(n26542), .A4(n26541), .ZN(
        n26551) );
  AOI22_X1 U27209 ( .A1(n27317), .A2(n27313), .B1(n27864), .B2(n27862), .ZN(
        n26548) );
  INV_X1 U27210 ( .A(n27872), .ZN(n26595) );
  AOI21_X1 U27211 ( .B1(n26595), .B2(n27875), .A(n3378), .ZN(n26547) );
  INV_X1 U27212 ( .A(n27327), .ZN(n26546) );
  NAND3_X1 U27213 ( .A1(n26548), .A2(n26547), .A3(n26546), .ZN(n26549) );
  AND3_X1 U27214 ( .A1(n26551), .A2(n26550), .A3(n26549), .ZN(Ciphertext[146])
         );
  AND2_X1 U27215 ( .A1(n26920), .A2(n26782), .ZN(n26554) );
  MUX2_X1 U27216 ( .A(n26554), .B(n26553), .S(n454), .Z(n26557) );
  MUX2_X1 U27217 ( .A(n4820), .B(n26920), .S(n26782), .Z(n26555) );
  NOR2_X1 U27218 ( .A1(n26917), .A2(n26555), .ZN(n26556) );
  NOR2_X2 U27219 ( .A1(n26557), .A2(n26556), .ZN(n27492) );
  AND2_X1 U27220 ( .A1(n26560), .A2(n26559), .ZN(n26561) );
  OAI21_X1 U27221 ( .B1(n26563), .B2(n377), .A(n28482), .ZN(n26564) );
  NAND2_X1 U27222 ( .A1(n26568), .A2(n1872), .ZN(n26566) );
  NOR3_X1 U27223 ( .A1(n26568), .A2(n26567), .A3(n26786), .ZN(n26569) );
  AOI21_X1 U27224 ( .B1(n26788), .B2(n5625), .A(n26569), .ZN(n26570) );
  OR2_X1 U27227 ( .A1(n26791), .A2(n26575), .ZN(n26922) );
  NOR2_X1 U27228 ( .A1(n29552), .A2(n26922), .ZN(n26577) );
  NAND3_X1 U27229 ( .A1(n27492), .A2(n29093), .A3(n27497), .ZN(n26589) );
  NAND2_X1 U27230 ( .A1(n26928), .A2(n29054), .ZN(n26586) );
  NOR2_X1 U27231 ( .A1(n28477), .A2(n26928), .ZN(n26584) );
  NAND2_X1 U27232 ( .A1(n26581), .A2(n29054), .ZN(n26583) );
  AOI21_X1 U27233 ( .B1(n26584), .B2(n26583), .A(n26582), .ZN(n26585) );
  OAI21_X1 U27234 ( .B1(n26933), .B2(n26586), .A(n26585), .ZN(n27493) );
  INV_X1 U27235 ( .A(n27493), .ZN(n26965) );
  NOR2_X1 U27236 ( .A1(n29522), .A2(n26965), .ZN(n26587) );
  NAND2_X1 U27237 ( .A1(n27492), .A2(n26587), .ZN(n26588) );
  INV_X1 U27238 ( .A(n3483), .ZN(n26590) );
  INV_X1 U27239 ( .A(n2404), .ZN(n26592) );
  XNOR2_X1 U27240 ( .A(n26593), .B(n26592), .ZN(Ciphertext[32]) );
  NOR2_X1 U27241 ( .A1(n27873), .A2(n27872), .ZN(n27311) );
  INV_X1 U27242 ( .A(n27311), .ZN(n26600) );
  NAND3_X1 U27243 ( .A1(n27872), .A2(n27877), .A3(n27863), .ZN(n26599) );
  NAND2_X1 U27244 ( .A1(n26595), .A2(n26594), .ZN(n26598) );
  INV_X1 U27245 ( .A(n27877), .ZN(n26596) );
  NOR2_X1 U27247 ( .A1(n28035), .A2(n29032), .ZN(n28026) );
  INV_X1 U27248 ( .A(n26602), .ZN(n28030) );
  MUX2_X1 U27249 ( .A(n29032), .B(n29160), .S(n28025), .Z(n26603) );
  INV_X1 U27250 ( .A(n3770), .ZN(n26604) );
  MUX2_X1 U27251 ( .A(n27465), .B(n27447), .S(n28435), .Z(n26608) );
  XNOR2_X1 U27254 ( .A(n26609), .B(n440), .ZN(Ciphertext[45]) );
  INV_X1 U27255 ( .A(n27379), .ZN(n27377) );
  OAI21_X1 U27256 ( .B1(n27209), .B2(n28393), .A(n27377), .ZN(n26613) );
  OAI21_X1 U27257 ( .B1(n5581), .B2(n446), .A(n27379), .ZN(n26612) );
  NOR2_X1 U27258 ( .A1(n295), .A2(n27382), .ZN(n26611) );
  NOR2_X1 U27259 ( .A1(n26614), .A2(n28452), .ZN(n26615) );
  NAND2_X1 U27260 ( .A1(n26616), .A2(n26615), .ZN(n26619) );
  NOR2_X1 U27261 ( .A1(n28545), .A2(n29520), .ZN(n26617) );
  NAND2_X1 U27262 ( .A1(n26617), .A2(n27066), .ZN(n26618) );
  MUX2_X1 U27263 ( .A(n26841), .B(n27085), .S(n27018), .Z(n26622) );
  NOR2_X1 U27264 ( .A1(n27018), .A2(n25815), .ZN(n26620) );
  MUX2_X1 U27265 ( .A(n26840), .B(n26620), .S(n26842), .Z(n26621) );
  NOR2_X1 U27266 ( .A1(n27050), .A2(n27014), .ZN(n26625) );
  MUX2_X1 U27268 ( .A(n26995), .B(n29481), .S(n28532), .Z(n26631) );
  NOR2_X1 U27270 ( .A1(n26632), .A2(n26998), .ZN(n26628) );
  INV_X1 U27274 ( .A(n29095), .ZN(n26640) );
  NAND2_X1 U27275 ( .A1(n6907), .A2(n26640), .ZN(n26644) );
  XNOR2_X1 U27276 ( .A(n26645), .B(n2804), .ZN(Ciphertext[142]) );
  OR2_X1 U27277 ( .A1(n29095), .A2(n27847), .ZN(n27858) );
  NAND2_X1 U27278 ( .A1(n27851), .A2(n27854), .ZN(n26646) );
  AOI21_X1 U27279 ( .B1(n27636), .B2(n27641), .A(n27639), .ZN(n26649) );
  OAI22_X1 U27280 ( .A1(n29532), .A2(n27641), .B1(n26978), .B2(n26980), .ZN(
        n27649) );
  INV_X1 U27281 ( .A(n27641), .ZN(n26648) );
  AOI22_X1 U27282 ( .A1(n26649), .A2(n27637), .B1(n27649), .B2(n26979), .ZN(
        n26650) );
  XNOR2_X1 U27283 ( .A(n26650), .B(n3256), .ZN(Ciphertext[97]) );
  NOR2_X1 U27284 ( .A1(n27202), .A2(n27203), .ZN(n26651) );
  AOI21_X1 U27285 ( .B1(n27539), .B2(n27202), .A(n26651), .ZN(n26655) );
  NOR2_X1 U27286 ( .A1(n27549), .A2(n27203), .ZN(n27541) );
  NOR2_X1 U27287 ( .A1(n27539), .A2(n28468), .ZN(n26653) );
  OAI21_X1 U27288 ( .B1(n26655), .B2(n27547), .A(n26654), .ZN(n26657) );
  XNOR2_X1 U27289 ( .A(n26657), .B(n26656), .ZN(Ciphertext[75]) );
  INV_X1 U27290 ( .A(n26658), .ZN(n26662) );
  INV_X1 U27291 ( .A(n26659), .ZN(n26660) );
  AND2_X1 U27292 ( .A1(n28038), .A2(n26660), .ZN(n26661) );
  NAND3_X1 U27293 ( .A1(n28036), .A2(n29160), .A3(n28025), .ZN(n26663) );
  OAI21_X1 U27294 ( .B1(n26664), .B2(n28026), .A(n26663), .ZN(n26666) );
  XNOR2_X1 U27295 ( .A(n26666), .B(n630), .ZN(Ciphertext[175]) );
  INV_X1 U27296 ( .A(n27427), .ZN(n27430) );
  OAI21_X1 U27297 ( .B1(n27428), .B2(n29542), .A(n27430), .ZN(n26667) );
  AOI22_X1 U27298 ( .A1(n26669), .A2(n26668), .B1(n27429), .B2(n26667), .ZN(
        n26670) );
  XNOR2_X1 U27299 ( .A(n26670), .B(n2996), .ZN(Ciphertext[29]) );
  NAND2_X1 U27300 ( .A1(n26978), .A2(n27641), .ZN(n26673) );
  OAI22_X1 U27301 ( .A1(n26979), .A2(n27636), .B1(n26673), .B2(n27638), .ZN(
        n26674) );
  NOR2_X1 U27302 ( .A1(n26675), .A2(n26674), .ZN(n26676) );
  XNOR2_X1 U27303 ( .A(n26676), .B(n2577), .ZN(Ciphertext[99]) );
  INV_X1 U27305 ( .A(n27818), .ZN(n27790) );
  INV_X1 U27306 ( .A(n27800), .ZN(n27822) );
  INV_X1 U27307 ( .A(n26680), .ZN(n26681) );
  INV_X1 U27308 ( .A(n26830), .ZN(n27438) );
  INV_X1 U27309 ( .A(n27442), .ZN(n26831) );
  OAI21_X1 U27310 ( .B1(n27442), .B2(n26710), .A(n25417), .ZN(n26683) );
  NAND2_X1 U27311 ( .A1(n26683), .A2(n27439), .ZN(n26684) );
  XNOR2_X1 U27312 ( .A(n26685), .B(n633), .ZN(Ciphertext[36]) );
  NOR2_X1 U27313 ( .A1(n27308), .A2(n27300), .ZN(n27310) );
  NOR2_X1 U27314 ( .A1(n27310), .A2(n29493), .ZN(n26687) );
  NAND2_X1 U27315 ( .A1(n26687), .A2(n26686), .ZN(n26688) );
  OAI21_X1 U27316 ( .B1(n26689), .B2(n26880), .A(n26688), .ZN(n26690) );
  XNOR2_X1 U27317 ( .A(n26690), .B(n3369), .ZN(Ciphertext[68]) );
  NAND2_X1 U27318 ( .A1(n27025), .A2(n29588), .ZN(n26691) );
  NOR2_X1 U27319 ( .A1(n26692), .A2(n27025), .ZN(n26693) );
  NOR2_X1 U27320 ( .A1(n26694), .A2(n26693), .ZN(n26695) );
  XNOR2_X1 U27321 ( .A(n26695), .B(n3607), .ZN(Ciphertext[30]) );
  NOR2_X1 U27322 ( .A1(n27859), .A2(n27847), .ZN(n26697) );
  AOI21_X1 U27323 ( .B1(n29095), .B2(n26697), .A(n26696), .ZN(n26700) );
  NAND3_X1 U27324 ( .A1(n27855), .A2(n29095), .A3(n27854), .ZN(n26699) );
  OAI211_X1 U27325 ( .C1(n27855), .C2(n27858), .A(n26700), .B(n26699), .ZN(
        n26702) );
  XNOR2_X1 U27326 ( .A(n26702), .B(n26701), .ZN(Ciphertext[138]) );
  NAND2_X1 U27327 ( .A1(n29093), .A2(n27497), .ZN(n27478) );
  INV_X1 U27328 ( .A(n3586), .ZN(n26703) );
  XNOR2_X1 U27329 ( .A(n26704), .B(n26703), .ZN(Ciphertext[51]) );
  OAI21_X1 U27330 ( .B1(n27025), .B2(n26817), .A(n27032), .ZN(n26706) );
  NOR2_X1 U27332 ( .A1(n27439), .A2(n26708), .ZN(n26709) );
  AOI21_X1 U27333 ( .B1(n26830), .B2(n27439), .A(n26709), .ZN(n27435) );
  NOR2_X1 U27334 ( .A1(n27433), .A2(n26710), .ZN(n26828) );
  AOI22_X1 U27335 ( .A1(n26831), .A2(n26833), .B1(n26828), .B2(n27438), .ZN(
        n26711) );
  OAI21_X1 U27336 ( .B1(n26712), .B2(n27435), .A(n26711), .ZN(n26714) );
  XNOR2_X1 U27337 ( .A(n26714), .B(n26713), .ZN(Ciphertext[39]) );
  NOR2_X1 U27338 ( .A1(n26716), .A2(n28459), .ZN(n26720) );
  NOR3_X1 U27340 ( .A1(n26723), .A2(n28548), .A3(n29560), .ZN(n26724) );
  OAI21_X1 U27342 ( .B1(n29579), .B2(n26727), .A(n26726), .ZN(n26732) );
  NOR2_X1 U27343 ( .A1(n28115), .A2(n28794), .ZN(n28094) );
  MUX2_X1 U27345 ( .A(n26742), .B(n26741), .S(n26740), .Z(n26743) );
  AOI21_X1 U27348 ( .B1(n29159), .B2(n26747), .A(n28563), .ZN(n26752) );
  AND2_X1 U27349 ( .A1(n29159), .A2(n26748), .ZN(n26751) );
  MUX2_X1 U27350 ( .A(n26752), .B(n26751), .S(n29099), .Z(n28103) );
  INV_X1 U27351 ( .A(n28089), .ZN(n28112) );
  AOI21_X1 U27352 ( .B1(n28591), .B2(n28112), .A(n29056), .ZN(n26763) );
  NAND2_X1 U27353 ( .A1(n26758), .A2(n26757), .ZN(n26759) );
  NAND3_X1 U27355 ( .A1(n28107), .A2(n28590), .A3(n29121), .ZN(n26762) );
  OAI21_X1 U27356 ( .B1(n26764), .B2(n26763), .A(n26762), .ZN(n26766) );
  INV_X1 U27357 ( .A(n3491), .ZN(n26765) );
  XNOR2_X1 U27358 ( .A(n26766), .B(n26765), .ZN(Ciphertext[186]) );
  MUX2_X1 U27359 ( .A(n26935), .B(n26768), .S(n26936), .Z(n26767) );
  NOR2_X1 U27360 ( .A1(n26767), .A2(n28541), .ZN(n26774) );
  NOR2_X2 U27363 ( .A1(n26774), .A2(n26773), .ZN(n27275) );
  MUX2_X1 U27364 ( .A(n26950), .B(n26775), .S(n29071), .Z(n26779) );
  NOR2_X1 U27365 ( .A1(n26949), .A2(n26775), .ZN(n26777) );
  NOR2_X1 U27366 ( .A1(n26948), .A2(n28542), .ZN(n26776) );
  MUX2_X1 U27367 ( .A(n26777), .B(n26776), .S(n26950), .Z(n26778) );
  AOI21_X2 U27368 ( .B1(n26948), .B2(n26779), .A(n26778), .ZN(n27291) );
  NOR2_X1 U27369 ( .A1(n457), .A2(n26920), .ZN(n26780) );
  NOR2_X1 U27370 ( .A1(n26781), .A2(n26780), .ZN(n26784) );
  MUX2_X1 U27371 ( .A(n26782), .B(n4820), .S(n26920), .Z(n26783) );
  MUX2_X1 U27372 ( .A(n27275), .B(n27291), .S(n27282), .Z(n26806) );
  NAND2_X1 U27373 ( .A1(n28471), .A2(n26911), .ZN(n26785) );
  AND3_X1 U27374 ( .A1(n26914), .A2(n5625), .A3(n26786), .ZN(n26787) );
  NOR2_X1 U27375 ( .A1(n25418), .A2(n26789), .ZN(n26790) );
  MUX2_X1 U27379 ( .A(n27286), .B(n27287), .S(n27275), .Z(n26805) );
  XNOR2_X1 U27383 ( .A(n26807), .B(n3414), .ZN(Ciphertext[62]) );
  XNOR2_X1 U27384 ( .A(n26810), .B(n3244), .ZN(Ciphertext[11]) );
  INV_X1 U27385 ( .A(n27277), .ZN(n27288) );
  NOR2_X1 U27386 ( .A1(n27282), .A2(n27288), .ZN(n26812) );
  NOR2_X1 U27388 ( .A1(n26812), .A2(n26811), .ZN(n26897) );
  INV_X1 U27389 ( .A(n27275), .ZN(n27290) );
  AOI21_X1 U27390 ( .B1(n27280), .B2(n27290), .A(n27287), .ZN(n26813) );
  OAI22_X1 U27391 ( .A1(n26897), .A2(n27291), .B1(n27278), .B2(n26813), .ZN(
        n26815) );
  XNOR2_X1 U27392 ( .A(n26815), .B(n26814), .ZN(Ciphertext[65]) );
  NOR2_X1 U27393 ( .A1(n27032), .A2(n306), .ZN(n26818) );
  NAND2_X1 U27394 ( .A1(n27025), .A2(n26818), .ZN(n26820) );
  INV_X1 U27395 ( .A(n3728), .ZN(n26821) );
  MUX2_X1 U27396 ( .A(n27354), .B(n29052), .S(n27357), .Z(n26824) );
  NAND2_X1 U27397 ( .A1(n27358), .A2(n28549), .ZN(n26822) );
  MUX2_X1 U27398 ( .A(n26822), .B(n27348), .S(n27357), .Z(n26823) );
  OAI21_X1 U27399 ( .B1(n26824), .B2(n27355), .A(n26823), .ZN(n26826) );
  XNOR2_X1 U27400 ( .A(n26826), .B(n26825), .ZN(Ciphertext[2]) );
  NOR2_X1 U27401 ( .A1(n25417), .A2(n26830), .ZN(n26827) );
  NOR2_X1 U27402 ( .A1(n26828), .A2(n26827), .ZN(n27443) );
  OAI211_X1 U27403 ( .C1(n26831), .C2(n27434), .A(n26830), .B(n26829), .ZN(
        n26832) );
  XNOR2_X1 U27405 ( .A(n26834), .B(n5892), .ZN(Ciphertext[37]) );
  MUX2_X1 U27406 ( .A(n27117), .B(n26835), .S(n28631), .Z(n26839) );
  MUX2_X1 U27407 ( .A(n27121), .B(n26836), .S(n27120), .Z(n26838) );
  INV_X1 U27408 ( .A(n27843), .ZN(n26846) );
  OAI21_X1 U27409 ( .B1(n26842), .B2(n25815), .A(n26840), .ZN(n26843) );
  NAND2_X1 U27410 ( .A1(n26843), .A2(n27088), .ZN(n26844) );
  OAI21_X1 U27412 ( .B1(n26849), .B2(n29575), .A(n29497), .ZN(n26853) );
  OAI21_X1 U27413 ( .B1(n26853), .B2(n26852), .A(n26851), .ZN(n26854) );
  AOI21_X1 U27414 ( .B1(n27137), .B2(n27138), .A(n26855), .ZN(n26856) );
  NOR2_X1 U27415 ( .A1(n26857), .A2(n26856), .ZN(n27830) );
  NAND2_X1 U27416 ( .A1(n28487), .A2(n26858), .ZN(n26859) );
  NOR2_X1 U27417 ( .A1(n26860), .A2(n26859), .ZN(n27829) );
  MUX2_X1 U27418 ( .A(n27074), .B(n27076), .S(n26991), .Z(n26864) );
  NAND2_X1 U27419 ( .A1(n26992), .A2(n27076), .ZN(n26861) );
  MUX2_X1 U27420 ( .A(n26862), .B(n26861), .S(n27074), .Z(n26863) );
  OAI21_X1 U27421 ( .B1(n26864), .B2(n28521), .A(n26863), .ZN(n27826) );
  NAND2_X1 U27422 ( .A1(n26866), .A2(n26865), .ZN(n27834) );
  NAND2_X1 U27423 ( .A1(n26867), .A2(n29048), .ZN(n26871) );
  INV_X1 U27424 ( .A(n26868), .ZN(n27159) );
  OAI21_X1 U27426 ( .B1(n27155), .B2(n29060), .A(n27154), .ZN(n26869) );
  OAI21_X1 U27427 ( .B1(n26871), .B2(n26870), .A(n26869), .ZN(n27831) );
  NAND2_X1 U27428 ( .A1(n27834), .A2(n27831), .ZN(n27841) );
  AOI21_X1 U27429 ( .B1(n27826), .B2(n27827), .A(n27841), .ZN(n26872) );
  XNOR2_X1 U27430 ( .A(n26873), .B(n625), .ZN(Ciphertext[132]) );
  MUX2_X1 U27431 ( .A(n27825), .B(n27101), .S(n27100), .Z(n26876) );
  NAND2_X1 U27432 ( .A1(n26902), .A2(n27826), .ZN(n26874) );
  OAI211_X1 U27433 ( .C1(n26876), .C2(n27828), .A(n26875), .B(n26874), .ZN(
        n26878) );
  XNOR2_X1 U27434 ( .A(n26878), .B(n26877), .ZN(Ciphertext[135]) );
  NOR2_X1 U27435 ( .A1(n27300), .A2(n26879), .ZN(n26886) );
  OAI21_X1 U27436 ( .B1(n26880), .B2(n28510), .A(n444), .ZN(n26883) );
  OAI211_X1 U27437 ( .C1(n26886), .C2(n26883), .A(n26882), .B(n26881), .ZN(
        n26884) );
  XNOR2_X1 U27438 ( .A(n26884), .B(n6174), .ZN(Ciphertext[69]) );
  NAND2_X1 U27439 ( .A1(n29493), .A2(n27255), .ZN(n26885) );
  XNOR2_X1 U27440 ( .A(n26888), .B(n3336), .ZN(Ciphertext[67]) );
  INV_X1 U27441 ( .A(n27727), .ZN(n26894) );
  INV_X1 U27442 ( .A(n326), .ZN(n27715) );
  OAI21_X1 U27443 ( .B1(n27714), .B2(n27715), .A(n26889), .ZN(n26893) );
  NOR2_X1 U27444 ( .A1(n324), .A2(n27728), .ZN(n27681) );
  NOR2_X1 U27445 ( .A1(n27725), .A2(n27711), .ZN(n26890) );
  AOI22_X1 U27446 ( .A1(n27691), .A2(n27681), .B1(n325), .B2(n26890), .ZN(
        n26892) );
  NAND2_X1 U27447 ( .A1(n27681), .A2(n27707), .ZN(n26891) );
  NAND2_X1 U27448 ( .A1(n27282), .A2(n27277), .ZN(n27285) );
  INV_X1 U27449 ( .A(n27285), .ZN(n26898) );
  INV_X1 U27450 ( .A(n27291), .ZN(n26895) );
  OAI211_X1 U27451 ( .C1(n26895), .C2(n27277), .A(n27275), .B(n27286), .ZN(
        n26896) );
  OAI21_X1 U27452 ( .B1(n26898), .B2(n26897), .A(n26896), .ZN(n26900) );
  XNOR2_X1 U27453 ( .A(n26900), .B(n26899), .ZN(Ciphertext[61]) );
  INV_X1 U27454 ( .A(n27841), .ZN(n26901) );
  INV_X1 U27455 ( .A(n26902), .ZN(n26905) );
  AND2_X1 U27456 ( .A1(n27101), .A2(n27100), .ZN(n26904) );
  NOR2_X1 U27457 ( .A1(n27826), .A2(n27827), .ZN(n27102) );
  INV_X1 U27458 ( .A(n27102), .ZN(n26903) );
  AOI22_X1 U27459 ( .A1(n26905), .A2(n27249), .B1(n26904), .B2(n26903), .ZN(
        n26906) );
  XNOR2_X1 U27460 ( .A(n26906), .B(n3374), .ZN(Ciphertext[133]) );
  NAND2_X1 U27461 ( .A1(n27235), .A2(n27447), .ZN(n26908) );
  INV_X1 U27462 ( .A(n27447), .ZN(n27472) );
  INV_X1 U27463 ( .A(n26909), .ZN(n26910) );
  MUX2_X1 U27464 ( .A(n26911), .B(n28423), .S(n28471), .Z(n26916) );
  INV_X1 U27465 ( .A(n27531), .ZN(n27506) );
  NAND2_X1 U27466 ( .A1(n26922), .A2(n26921), .ZN(n26923) );
  OAI21_X1 U27467 ( .B1(n26925), .B2(n26924), .A(n26923), .ZN(n27528) );
  INV_X1 U27468 ( .A(n27528), .ZN(n27502) );
  AOI22_X1 U27469 ( .A1(n26928), .A2(n5505), .B1(n26927), .B2(n1279), .ZN(
        n26932) );
  INV_X1 U27470 ( .A(n26929), .ZN(n26931) );
  MUX2_X1 U27471 ( .A(n26932), .B(n26931), .S(n26930), .Z(n26934) );
  OAI21_X1 U27472 ( .B1(n27520), .B2(n27502), .A(n27527), .ZN(n26958) );
  AND2_X1 U27473 ( .A1(n6768), .A2(n26935), .ZN(n26939) );
  NOR2_X1 U27474 ( .A1(n6768), .A2(n26936), .ZN(n26938) );
  OAI21_X1 U27475 ( .B1(n26939), .B2(n26938), .A(n28541), .ZN(n26946) );
  NOR2_X1 U27476 ( .A1(n28541), .A2(n26940), .ZN(n26942) );
  INV_X1 U27478 ( .A(n26950), .ZN(n26954) );
  AOI21_X1 U27479 ( .B1(n29071), .B2(n28542), .A(n28646), .ZN(n26953) );
  NAND3_X1 U27481 ( .A1(n27527), .A2(n27528), .A3(n27525), .ZN(n26956) );
  OAI21_X1 U27482 ( .B1(n27506), .B2(n27221), .A(n26956), .ZN(n26957) );
  AOI21_X1 U27483 ( .B1(n27506), .B2(n26958), .A(n26957), .ZN(n26959) );
  XNOR2_X1 U27484 ( .A(n26959), .B(n2544), .ZN(Ciphertext[59]) );
  OAI21_X1 U27485 ( .B1(n27386), .B2(n27410), .A(n28177), .ZN(n26962) );
  OAI21_X1 U27486 ( .B1(n27400), .B2(n27387), .A(n27390), .ZN(n26961) );
  NAND2_X1 U27488 ( .A1(n27496), .A2(n27493), .ZN(n26964) );
  OAI21_X1 U27489 ( .B1(n27494), .B2(n27480), .A(n26964), .ZN(n27477) );
  INV_X1 U27490 ( .A(n27498), .ZN(n27487) );
  OAI21_X1 U27491 ( .B1(n27487), .B2(n26965), .A(n27496), .ZN(n26966) );
  AOI22_X1 U27492 ( .A1(n5368), .A2(n27477), .B1(n26966), .B2(n29093), .ZN(
        n26967) );
  XNOR2_X1 U27493 ( .A(n26967), .B(n2916), .ZN(Ciphertext[53]) );
  OAI21_X1 U27494 ( .B1(n27417), .B2(n27426), .A(n26968), .ZN(n26971) );
  NAND2_X1 U27496 ( .A1(n29529), .A2(n27425), .ZN(n26969) );
  INV_X1 U27497 ( .A(n27424), .ZN(n27420) );
  NOR2_X1 U27498 ( .A1(n26971), .A2(n26970), .ZN(n26972) );
  INV_X1 U27500 ( .A(n27629), .ZN(n26973) );
  OAI21_X1 U27501 ( .B1(n26973), .B2(n27627), .A(n27630), .ZN(n26974) );
  NOR2_X1 U27502 ( .A1(n27614), .A2(n27625), .ZN(n27609) );
  NAND2_X1 U27503 ( .A1(n1912), .A2(n27632), .ZN(n27601) );
  OAI22_X1 U27504 ( .A1(n26974), .A2(n27609), .B1(n27601), .B2(n27625), .ZN(
        n26976) );
  NOR2_X1 U27505 ( .A1(n1912), .A2(n27630), .ZN(n27607) );
  AND2_X1 U27506 ( .A1(n27607), .A2(n27628), .ZN(n26975) );
  NOR2_X1 U27507 ( .A1(n26976), .A2(n26975), .ZN(n26977) );
  XNOR2_X1 U27508 ( .A(n26977), .B(n2973), .ZN(Ciphertext[93]) );
  OAI21_X1 U27509 ( .B1(n27636), .B2(n27641), .A(n26978), .ZN(n26982) );
  OAI21_X1 U27510 ( .B1(n26980), .B2(n27638), .A(n26979), .ZN(n26981) );
  XNOR2_X1 U27512 ( .A(n26983), .B(Key[173]), .ZN(Ciphertext[96]) );
  INV_X1 U27515 ( .A(n28021), .ZN(n28006) );
  OAI21_X1 U27516 ( .B1(n28006), .B2(n28003), .A(n28015), .ZN(n26985) );
  AOI22_X1 U27517 ( .A1(n26986), .A2(n28006), .B1(n28411), .B2(n26985), .ZN(
        n26987) );
  XNOR2_X1 U27518 ( .A(n26987), .B(n1919), .ZN(Ciphertext[168]) );
  INV_X1 U27520 ( .A(n27944), .ZN(n27927) );
  MUX2_X1 U27521 ( .A(n29500), .B(n27069), .S(n28660), .Z(n27000) );
  MUX2_X1 U27522 ( .A(n28452), .B(n29076), .S(n28545), .Z(n26999) );
  MUX2_X1 U27523 ( .A(n27000), .B(n26999), .S(n29520), .Z(n27925) );
  NOR2_X1 U27524 ( .A1(n27004), .A2(n29058), .ZN(n27005) );
  NAND2_X1 U27525 ( .A1(n27005), .A2(n398), .ZN(n27008) );
  AND2_X1 U27526 ( .A1(n28783), .A2(n28130), .ZN(n27006) );
  NAND2_X1 U27527 ( .A1(n27041), .A2(n27006), .ZN(n27007) );
  NOR2_X1 U27529 ( .A1(n26623), .A2(n27014), .ZN(n27012) );
  NOR2_X1 U27530 ( .A1(n27010), .A2(n28639), .ZN(n27011) );
  NAND2_X1 U27531 ( .A1(n29062), .A2(n27013), .ZN(n27015) );
  NAND2_X1 U27532 ( .A1(n27015), .A2(n27014), .ZN(n27016) );
  NOR2_X1 U27533 ( .A1(n26507), .A2(n27018), .ZN(n27089) );
  NOR3_X1 U27534 ( .A1(n27089), .A2(n27086), .A3(n27085), .ZN(n27019) );
  AOI21_X1 U27535 ( .B1(n27927), .B2(n27023), .A(n27022), .ZN(n27024) );
  XNOR2_X1 U27536 ( .A(n27024), .B(n3643), .ZN(Ciphertext[160]) );
  NOR2_X1 U27537 ( .A1(n27032), .A2(n29588), .ZN(n27027) );
  NAND2_X1 U27538 ( .A1(n27027), .A2(n28592), .ZN(n27031) );
  NOR2_X1 U27539 ( .A1(n6568), .A2(n306), .ZN(n27030) );
  INV_X1 U27540 ( .A(n27034), .ZN(n27035) );
  AOI22_X1 U27541 ( .A1(n27035), .A2(n28000), .B1(n28005), .B2(n28022), .ZN(
        n27036) );
  XNOR2_X1 U27542 ( .A(n27036), .B(n2353), .ZN(Ciphertext[169]) );
  OAI21_X1 U27543 ( .B1(n27382), .B2(n28393), .A(n27379), .ZN(n27037) );
  XNOR2_X1 U27544 ( .A(n27039), .B(n3787), .ZN(Ciphertext[12]) );
  NAND2_X1 U27545 ( .A1(n27048), .A2(n28130), .ZN(n27046) );
  MUX2_X1 U27546 ( .A(n4497), .B(n27046), .S(n27045), .Z(n27047) );
  AOI21_X1 U27548 ( .B1(n29062), .B2(n26623), .A(n27049), .ZN(n27051) );
  OR2_X1 U27549 ( .A1(n29536), .A2(n27898), .ZN(n27058) );
  OAI211_X1 U27550 ( .C1(n29536), .C2(n27056), .A(n27902), .B(n27055), .ZN(
        n27057) );
  OAI21_X1 U27551 ( .B1(n29497), .B2(n27058), .A(n27057), .ZN(n27062) );
  NOR2_X1 U27552 ( .A1(n27902), .A2(n29575), .ZN(n27903) );
  AND2_X1 U27553 ( .A1(n27903), .A2(n27060), .ZN(n27061) );
  NOR2_X1 U27554 ( .A1(n922), .A2(n27063), .ZN(n27064) );
  NOR2_X1 U27555 ( .A1(n27065), .A2(n27064), .ZN(n27073) );
  INV_X1 U27556 ( .A(n27066), .ZN(n27072) );
  NOR2_X1 U27557 ( .A1(n28228), .A2(n28545), .ZN(n27071) );
  NOR2_X1 U27558 ( .A1(n27069), .A2(n29076), .ZN(n27070) );
  OAI211_X1 U27559 ( .C1(n27092), .C2(n27908), .A(n27905), .B(n27080), .ZN(
        n27094) );
  NAND2_X1 U27560 ( .A1(n27077), .A2(n27076), .ZN(n27078) );
  AND2_X1 U27561 ( .A1(n27079), .A2(n27078), .ZN(n27899) );
  INV_X1 U27563 ( .A(n28453), .ZN(n27918) );
  OAI21_X1 U27564 ( .B1(n27919), .B2(n27920), .A(n27918), .ZN(n27093) );
  AOI21_X1 U27565 ( .B1(n27084), .B2(n28458), .A(n27081), .ZN(n27083) );
  OAI21_X1 U27566 ( .B1(n27088), .B2(n27084), .A(n27083), .ZN(n27091) );
  OAI21_X1 U27567 ( .B1(n27087), .B2(n27086), .A(n27085), .ZN(n27090) );
  INV_X1 U27568 ( .A(n27271), .ZN(n27913) );
  AOI22_X1 U27569 ( .A1(n27094), .A2(n27093), .B1(n27889), .B2(n27092), .ZN(
        n27095) );
  XNOR2_X1 U27570 ( .A(n27095), .B(n3422), .ZN(Ciphertext[150]) );
  OAI21_X1 U27571 ( .B1(n27520), .B2(n27528), .A(n27096), .ZN(n27097) );
  XNOR2_X1 U27572 ( .A(n27098), .B(n3109), .ZN(Ciphertext[57]) );
  NAND2_X1 U27573 ( .A1(n27825), .A2(n27099), .ZN(n27104) );
  NAND2_X1 U27574 ( .A1(n27102), .A2(n27828), .ZN(n27103) );
  NAND2_X1 U27575 ( .A1(n27703), .A2(n27161), .ZN(n27106) );
  INV_X1 U27577 ( .A(n27755), .ZN(n27745) );
  AOI21_X1 U27578 ( .B1(n27155), .B2(n29474), .A(n27152), .ZN(n27116) );
  INV_X1 U27579 ( .A(n27109), .ZN(n27115) );
  NOR2_X1 U27580 ( .A1(n29474), .A2(n27159), .ZN(n27113) );
  NOR2_X1 U27581 ( .A1(n27153), .A2(n29048), .ZN(n27112) );
  NAND2_X1 U27583 ( .A1(n27745), .A2(n29049), .ZN(n27227) );
  AOI21_X1 U27584 ( .B1(n28631), .B2(n402), .A(n27117), .ZN(n27119) );
  INV_X1 U27585 ( .A(n27128), .ZN(n27732) );
  MUX2_X1 U27586 ( .A(n27124), .B(n27123), .S(n27193), .Z(n27127) );
  NAND2_X1 U27587 ( .A1(n27130), .A2(n27175), .ZN(n27133) );
  NAND3_X1 U27588 ( .A1(n27173), .A2(n27131), .A3(n28536), .ZN(n27132) );
  AOI21_X1 U27589 ( .B1(n27137), .B2(n27142), .A(n27136), .ZN(n27145) );
  NAND2_X1 U27590 ( .A1(n27139), .A2(n27138), .ZN(n27144) );
  NOR3_X1 U27591 ( .A1(n27142), .A2(n28487), .A3(n29621), .ZN(n27143) );
  AOI21_X1 U27592 ( .B1(n27145), .B2(n27144), .A(n27143), .ZN(n27146) );
  OAI21_X1 U27593 ( .B1(n27690), .B2(n27147), .A(n27146), .ZN(n27739) );
  INV_X1 U27594 ( .A(n27739), .ZN(n27757) );
  NOR2_X1 U27595 ( .A1(n27551), .A2(n29085), .ZN(n27148) );
  NOR2_X1 U27596 ( .A1(n27572), .A2(n27562), .ZN(n27576) );
  MUX2_X1 U27597 ( .A(n27148), .B(n27576), .S(n27552), .Z(n27150) );
  NOR2_X1 U27598 ( .A1(n27561), .A2(n27562), .ZN(n27554) );
  OAI21_X1 U27599 ( .B1(n27155), .B2(n27154), .A(n27153), .ZN(n27156) );
  OR2_X1 U27601 ( .A1(n27704), .A2(n27703), .ZN(n27162) );
  OAI21_X1 U27602 ( .B1(n27169), .B2(n27168), .A(n27167), .ZN(n27170) );
  NOR2_X1 U27603 ( .A1(n28392), .A2(n29132), .ZN(n27172) );
  AOI21_X1 U27604 ( .B1(n28392), .B2(n27173), .A(n27172), .ZN(n27180) );
  MUX2_X1 U27605 ( .A(n27177), .B(n28536), .S(n27175), .Z(n27179) );
  INV_X1 U27606 ( .A(n27661), .ZN(n27674) );
  NAND2_X1 U27607 ( .A1(n26396), .A2(n25124), .ZN(n27185) );
  OAI21_X1 U27608 ( .B1(n27183), .B2(n27182), .A(n27181), .ZN(n27184) );
  OAI21_X1 U27609 ( .B1(n28652), .B2(n27185), .A(n27184), .ZN(n27187) );
  OAI21_X1 U27610 ( .B1(n28650), .B2(n27188), .A(n27187), .ZN(n27671) );
  NOR2_X1 U27612 ( .A1(n27652), .A2(n27676), .ZN(n27194) );
  AOI211_X1 U27613 ( .C1(n27196), .C2(n27674), .A(n27195), .B(n27194), .ZN(
        n27197) );
  XNOR2_X1 U27614 ( .A(n27197), .B(n3164), .ZN(Ciphertext[105]) );
  NAND2_X1 U27615 ( .A1(n27537), .A2(n27202), .ZN(n27198) );
  OAI21_X1 U27617 ( .B1(n27537), .B2(n27538), .A(n28386), .ZN(n27201) );
  NOR2_X1 U27618 ( .A1(n27201), .A2(n27200), .ZN(n27207) );
  NAND2_X1 U27619 ( .A1(n27547), .A2(n27548), .ZN(n27205) );
  NAND2_X1 U27621 ( .A1(n394), .A2(n27203), .ZN(n27204) );
  NOR2_X1 U27623 ( .A1(n295), .A2(n446), .ZN(n27211) );
  AND2_X1 U27624 ( .A1(n27208), .A2(n27379), .ZN(n27210) );
  XNOR2_X1 U27626 ( .A(n27215), .B(n28693), .ZN(Ciphertext[15]) );
  NOR2_X1 U27627 ( .A1(n27572), .A2(n27561), .ZN(n27216) );
  XNOR2_X1 U27629 ( .A(n27220), .B(n2986), .ZN(Ciphertext[82]) );
  NOR3_X1 U27630 ( .A1(n27531), .A2(n27505), .A3(n29556), .ZN(n27224) );
  INV_X1 U27631 ( .A(n27527), .ZN(n27222) );
  NAND2_X1 U27632 ( .A1(n27755), .A2(n397), .ZN(n27226) );
  INV_X1 U27633 ( .A(n27759), .ZN(n27749) );
  AOI21_X1 U27634 ( .B1(n27227), .B2(n27226), .A(n27749), .ZN(n27230) );
  NAND2_X1 U27636 ( .A1(n28445), .A2(n27732), .ZN(n27228) );
  XNOR2_X1 U27637 ( .A(n27232), .B(n27231), .ZN(Ciphertext[117]) );
  AOI21_X1 U27638 ( .B1(n27762), .B2(n27777), .A(n6419), .ZN(n27233) );
  XNOR2_X1 U27639 ( .A(n27234), .B(n3180), .ZN(Ciphertext[120]) );
  OAI211_X1 U27640 ( .C1(n27235), .C2(n27472), .A(n27465), .B(n27467), .ZN(
        n27238) );
  NAND2_X1 U27641 ( .A1(n27447), .A2(n27236), .ZN(n27237) );
  OAI211_X1 U27642 ( .C1(n27458), .C2(n27447), .A(n27238), .B(n27237), .ZN(
        n27240) );
  INV_X1 U27643 ( .A(n2403), .ZN(n27239) );
  XNOR2_X1 U27644 ( .A(n27240), .B(n27239), .ZN(Ciphertext[43]) );
  OAI21_X1 U27645 ( .B1(n27400), .B2(n27386), .A(n27241), .ZN(n27243) );
  INV_X1 U27646 ( .A(n27387), .ZN(n27242) );
  MUX2_X1 U27647 ( .A(n27246), .B(n27245), .S(n28441), .Z(n27247) );
  XNOR2_X1 U27648 ( .A(n27247), .B(n2981), .ZN(Ciphertext[158]) );
  NAND2_X1 U27649 ( .A1(n27248), .A2(n27841), .ZN(n27250) );
  AOI21_X1 U27652 ( .B1(n27278), .B2(n27253), .A(n27252), .ZN(n27254) );
  XNOR2_X1 U27653 ( .A(n27254), .B(n2511), .ZN(Ciphertext[63]) );
  OAI21_X1 U27655 ( .B1(n6910), .B2(n395), .A(n29619), .ZN(n27262) );
  NOR2_X1 U27656 ( .A1(n28510), .A2(n27300), .ZN(n27260) );
  OAI21_X1 U27657 ( .B1(n27260), .B2(n27259), .A(n27255), .ZN(n27261) );
  NAND2_X1 U27658 ( .A1(n27262), .A2(n27261), .ZN(n27264) );
  XNOR2_X1 U27659 ( .A(n27264), .B(n27263), .ZN(Ciphertext[66]) );
  INV_X1 U27660 ( .A(n27265), .ZN(n27266) );
  INV_X1 U27661 ( .A(n27596), .ZN(n27588) );
  NOR3_X1 U27662 ( .A1(n27588), .A2(n27597), .A3(n27585), .ZN(n27268) );
  NOR3_X1 U27663 ( .A1(n27596), .A2(n28429), .A3(n28179), .ZN(n27267) );
  NOR3_X1 U27664 ( .A1(n27269), .A2(n27268), .A3(n27267), .ZN(n27270) );
  XNOR2_X1 U27665 ( .A(n27270), .B(n3385), .ZN(Ciphertext[88]) );
  INV_X1 U27666 ( .A(n27889), .ZN(n27273) );
  OAI22_X1 U27667 ( .A1(n27919), .A2(n27905), .B1(n27923), .B2(n27908), .ZN(
        n27921) );
  INV_X1 U27668 ( .A(n27919), .ZN(n27272) );
  NOR2_X1 U27669 ( .A1(n27272), .A2(n27080), .ZN(n27893) );
  AOI22_X1 U27670 ( .A1(n27273), .A2(n27921), .B1(n27883), .B2(n27893), .ZN(
        n27274) );
  XNOR2_X1 U27671 ( .A(n27274), .B(Key[126]), .ZN(Ciphertext[151]) );
  MUX2_X1 U27672 ( .A(n27277), .B(n27282), .S(n27275), .Z(n27276) );
  NAND2_X1 U27673 ( .A1(n27276), .A2(n27281), .ZN(n27284) );
  NOR2_X1 U27674 ( .A1(n27291), .A2(n27277), .ZN(n27279) );
  NAND2_X1 U27675 ( .A1(n27279), .A2(n27278), .ZN(n27283) );
  OAI21_X1 U27676 ( .B1(n27286), .B2(n27290), .A(n27285), .ZN(n27292) );
  OAI21_X1 U27677 ( .B1(n27291), .B2(n2438), .A(n27287), .ZN(n27289) );
  AOI22_X1 U27678 ( .A1(n27292), .A2(n27291), .B1(n27290), .B2(n27289), .ZN(
        n27293) );
  XNOR2_X1 U27679 ( .A(n27293), .B(n3451), .ZN(Ciphertext[60]) );
  NAND2_X1 U27680 ( .A1(n28655), .A2(n27663), .ZN(n27295) );
  AOI21_X1 U27681 ( .B1(n27676), .B2(n27672), .A(n27673), .ZN(n27294) );
  AOI21_X1 U27682 ( .B1(n29091), .B2(n27295), .A(n27294), .ZN(n27297) );
  INV_X1 U27683 ( .A(n27664), .ZN(n27668) );
  NOR2_X1 U27684 ( .A1(n27652), .A2(n28655), .ZN(n27296) );
  NOR3_X1 U27685 ( .A1(n27297), .A2(n27668), .A3(n27296), .ZN(n27299) );
  XNOR2_X1 U27686 ( .A(n27299), .B(n27298), .ZN(Ciphertext[102]) );
  INV_X1 U27687 ( .A(n27303), .ZN(n27306) );
  NOR2_X1 U27688 ( .A1(n27317), .A2(n27324), .ZN(n27314) );
  INV_X1 U27689 ( .A(n27313), .ZN(n27319) );
  NOR2_X1 U27690 ( .A1(n27875), .A2(n27324), .ZN(n27316) );
  AOI22_X1 U27691 ( .A1(n27314), .A2(n27319), .B1(n27311), .B2(n27316), .ZN(
        n27326) );
  NOR3_X1 U27692 ( .A1(n27875), .A2(n3537), .A3(n27871), .ZN(n27312) );
  NOR2_X1 U27693 ( .A1(n27875), .A2(n27872), .ZN(n27315) );
  OAI21_X1 U27694 ( .B1(n27315), .B2(n3537), .A(n27862), .ZN(n27322) );
  NAND2_X1 U27695 ( .A1(n27316), .A2(n29504), .ZN(n27321) );
  NOR2_X1 U27696 ( .A1(n27317), .A2(n3537), .ZN(n27318) );
  NAND2_X1 U27697 ( .A1(n27319), .A2(n27318), .ZN(n27320) );
  INV_X1 U27699 ( .A(n27328), .ZN(n27332) );
  OAI22_X1 U27700 ( .A1(n5421), .A2(n27357), .B1(n27358), .B2(n27355), .ZN(
        n27329) );
  NAND2_X1 U27701 ( .A1(n27329), .A2(n27340), .ZN(n27331) );
  OAI211_X1 U27702 ( .C1(n27332), .C2(n27353), .A(n27331), .B(n27330), .ZN(
        n27334) );
  XNOR2_X1 U27703 ( .A(n27334), .B(n27333), .ZN(Ciphertext[0]) );
  AND2_X1 U27704 ( .A1(n27358), .A2(n2522), .ZN(n27343) );
  XNOR2_X1 U27705 ( .A(n27354), .B(n2522), .ZN(n27335) );
  OAI21_X1 U27706 ( .B1(n27335), .B2(n27358), .A(n27357), .ZN(n27336) );
  AOI21_X1 U27707 ( .B1(n27340), .B2(n27343), .A(n27336), .ZN(n27347) );
  INV_X1 U27708 ( .A(n2522), .ZN(n27337) );
  OAI21_X1 U27709 ( .B1(n27358), .B2(n27337), .A(n27351), .ZN(n27339) );
  OR2_X1 U27710 ( .A1(n27351), .A2(n27337), .ZN(n27338) );
  AOI21_X1 U27711 ( .B1(n27339), .B2(n27338), .A(n27357), .ZN(n27346) );
  INV_X1 U27712 ( .A(n27340), .ZN(n27342) );
  INV_X1 U27713 ( .A(n27357), .ZN(n27349) );
  NOR3_X1 U27714 ( .A1(n27350), .A2(n2522), .A3(n28549), .ZN(n27341) );
  OAI21_X1 U27715 ( .B1(n27342), .B2(n27349), .A(n27341), .ZN(n27345) );
  OAI211_X1 U27716 ( .C1(n27351), .C2(n27357), .A(n27343), .B(n28549), .ZN(
        n27344) );
  OAI211_X1 U27717 ( .C1(n27347), .C2(n27346), .A(n27345), .B(n27344), .ZN(
        Ciphertext[1]) );
  INV_X1 U27718 ( .A(n27348), .ZN(n27360) );
  OAI21_X1 U27719 ( .B1(n27351), .B2(n27350), .A(n27349), .ZN(n27359) );
  NOR2_X1 U27720 ( .A1(n27354), .A2(n28549), .ZN(n27356) );
  XNOR2_X1 U27721 ( .A(n27361), .B(n629), .ZN(Ciphertext[3]) );
  AOI211_X1 U27722 ( .C1(n29541), .C2(n27362), .A(n3751), .B(n27364), .ZN(
        n27367) );
  NAND2_X1 U27723 ( .A1(n27365), .A2(n27364), .ZN(n27375) );
  NAND2_X1 U27725 ( .A1(n27368), .A2(n27370), .ZN(n27369) );
  NAND3_X1 U27726 ( .A1(n28494), .A2(n27372), .A3(n29541), .ZN(n27374) );
  OAI21_X1 U27728 ( .B1(n27380), .B2(n27379), .A(n295), .ZN(n27381) );
  XNOR2_X1 U27730 ( .A(n27385), .B(n27384), .ZN(Ciphertext[17]) );
  OAI22_X1 U27731 ( .A1(n27400), .A2(n28177), .B1(n27386), .B2(n342), .ZN(
        n27411) );
  NOR2_X1 U27732 ( .A1(n25629), .A2(n27387), .ZN(n27389) );
  AOI22_X1 U27733 ( .A1(n27411), .A2(n27390), .B1(n27389), .B2(n27388), .ZN(
        n27391) );
  XNOR2_X1 U27734 ( .A(n27391), .B(n3196), .ZN(Ciphertext[19]) );
  NOR2_X1 U27735 ( .A1(n27408), .A2(n27392), .ZN(n27399) );
  INV_X1 U27736 ( .A(n27393), .ZN(n27397) );
  MUX2_X1 U27737 ( .A(n27397), .B(n27396), .S(n27395), .Z(n27398) );
  AOI22_X1 U27738 ( .A1(n27400), .A2(n28177), .B1(n27399), .B2(n27398), .ZN(
        n27401) );
  OAI222_X1 U27739 ( .A1(n27404), .A2(n27410), .B1(n27403), .B2(n28177), .C1(
        n27402), .C2(n27401), .ZN(n27406) );
  INV_X1 U27740 ( .A(n3457), .ZN(n27405) );
  XNOR2_X1 U27741 ( .A(n27406), .B(n27405), .ZN(Ciphertext[22]) );
  OAI21_X1 U27742 ( .B1(n27409), .B2(n28177), .A(n342), .ZN(n27413) );
  NAND2_X1 U27743 ( .A1(n27411), .A2(n4922), .ZN(n27412) );
  NAND2_X1 U27744 ( .A1(n27413), .A2(n27412), .ZN(n27414) );
  XNOR2_X1 U27745 ( .A(n27414), .B(n4222), .ZN(Ciphertext[23]) );
  OAI21_X1 U27748 ( .B1(n27426), .B2(n6738), .A(n27427), .ZN(n27419) );
  AOI22_X1 U27749 ( .A1(n27421), .A2(n27426), .B1(n27420), .B2(n27419), .ZN(
        n27423) );
  XNOR2_X1 U27750 ( .A(n27423), .B(n27422), .ZN(Ciphertext[24]) );
  INV_X1 U27752 ( .A(n2982), .ZN(n27436) );
  XNOR2_X1 U27753 ( .A(n27437), .B(n27436), .ZN(Ciphertext[38]) );
  AOI21_X1 U27754 ( .B1(n27439), .B2(n27438), .A(n25417), .ZN(n27440) );
  OAI22_X1 U27755 ( .A1(n27443), .A2(n27442), .B1(n27441), .B2(n27440), .ZN(
        n27445) );
  XNOR2_X1 U27756 ( .A(n27445), .B(n27444), .ZN(Ciphertext[41]) );
  NAND3_X1 U27757 ( .A1(n27458), .A2(n27457), .A3(n27472), .ZN(n27451) );
  INV_X1 U27758 ( .A(n27446), .ZN(n27450) );
  OR3_X1 U27759 ( .A1(n27465), .A2(n27447), .A3(n27457), .ZN(n27449) );
  NAND3_X1 U27760 ( .A1(n27457), .A2(n27465), .A3(n28435), .ZN(n27448) );
  INV_X1 U27761 ( .A(n27452), .ZN(n27453) );
  INV_X1 U27762 ( .A(n27462), .ZN(n27466) );
  NOR2_X1 U27763 ( .A1(n27465), .A2(n27466), .ZN(n27461) );
  AND2_X1 U27764 ( .A1(n27465), .A2(n27466), .ZN(n27454) );
  NOR2_X1 U27765 ( .A1(n27461), .A2(n27454), .ZN(n27456) );
  AOI21_X1 U27767 ( .B1(n27456), .B2(n4823), .A(n27472), .ZN(n27474) );
  XNOR2_X1 U27768 ( .A(n27457), .B(n27462), .ZN(n27459) );
  NAND2_X1 U27769 ( .A1(n27459), .A2(n27458), .ZN(n27473) );
  NAND2_X1 U27770 ( .A1(n27461), .A2(n28435), .ZN(n27470) );
  XNOR2_X1 U27771 ( .A(n27463), .B(n27462), .ZN(n27464) );
  NAND2_X1 U27772 ( .A1(n27464), .A2(n27465), .ZN(n27469) );
  NAND3_X1 U27773 ( .A1(n449), .A2(n27467), .A3(n27466), .ZN(n27468) );
  NAND3_X1 U27774 ( .A1(n27470), .A2(n27469), .A3(n27468), .ZN(n27471) );
  AOI22_X1 U27775 ( .A1(n27474), .A2(n27473), .B1(n27472), .B2(n27471), .ZN(
        Ciphertext[44]) );
  AOI22_X1 U27777 ( .A1(n27478), .A2(n27477), .B1(n27476), .B2(n27475), .ZN(
        n27479) );
  XNOR2_X1 U27778 ( .A(n27479), .B(n1225), .ZN(Ciphertext[49]) );
  XNOR2_X1 U27779 ( .A(n27492), .B(n3501), .ZN(n27484) );
  NAND2_X1 U27780 ( .A1(n29093), .A2(n27480), .ZN(n27483) );
  XNOR2_X1 U27781 ( .A(n29523), .B(n5513), .ZN(n27482) );
  OR2_X1 U27782 ( .A1(n29093), .A2(n27497), .ZN(n27481) );
  OAI22_X1 U27783 ( .A1(n27484), .A2(n27483), .B1(n27482), .B2(n27481), .ZN(
        n27491) );
  XNOR2_X1 U27784 ( .A(n27496), .B(n3501), .ZN(n27485) );
  OAI21_X1 U27785 ( .B1(n27485), .B2(n29522), .A(n27497), .ZN(n27489) );
  XNOR2_X1 U27786 ( .A(n27493), .B(n3501), .ZN(n27486) );
  NOR2_X1 U27787 ( .A1(n27487), .A2(n27486), .ZN(n27488) );
  NOR2_X1 U27788 ( .A1(n27489), .A2(n27488), .ZN(n27490) );
  NOR2_X1 U27789 ( .A1(n27491), .A2(n27490), .ZN(Ciphertext[50]) );
  NOR2_X1 U27791 ( .A1(n27496), .A2(n27493), .ZN(n27495) );
  NAND3_X1 U27792 ( .A1(n29522), .A2(n27497), .A3(n27496), .ZN(n27499) );
  XNOR2_X1 U27793 ( .A(n27501), .B(n628), .ZN(Ciphertext[52]) );
  NAND3_X1 U27794 ( .A1(n27520), .A2(n27502), .A3(n27510), .ZN(n27504) );
  NAND3_X1 U27795 ( .A1(n27527), .A2(n27526), .A3(n27528), .ZN(n27503) );
  OAI211_X1 U27796 ( .C1(n27506), .C2(n27505), .A(n27504), .B(n27503), .ZN(
        n27507) );
  XNOR2_X1 U27797 ( .A(n27507), .B(n632), .ZN(Ciphertext[55]) );
  INV_X1 U27798 ( .A(n27509), .ZN(n27512) );
  AOI21_X1 U27799 ( .B1(n27531), .B2(n27512), .A(n27511), .ZN(n27514) );
  NOR3_X1 U27800 ( .A1(n27526), .A2(n27520), .A3(n27528), .ZN(n27516) );
  NAND2_X1 U27801 ( .A1(n27516), .A2(n27515), .ZN(n27517) );
  AND3_X1 U27802 ( .A1(n27518), .A2(n27519), .A3(n27517), .ZN(Ciphertext[56])
         );
  INV_X1 U27803 ( .A(n27531), .ZN(n27521) );
  AOI21_X1 U27804 ( .B1(n27524), .B2(n27523), .A(n27522), .ZN(n27533) );
  AND2_X1 U27805 ( .A1(n27526), .A2(n27525), .ZN(n27530) );
  NOR3_X1 U27806 ( .A1(n27531), .A2(n27528), .A3(n27527), .ZN(n27529) );
  AOI21_X1 U27807 ( .B1(n27531), .B2(n27530), .A(n27529), .ZN(n27532) );
  OAI21_X1 U27810 ( .B1(n27541), .B2(n28386), .A(n27539), .ZN(n27542) );
  OAI21_X1 U27811 ( .B1(n27543), .B2(n394), .A(n27542), .ZN(n27544) );
  XNOR2_X1 U27812 ( .A(n27544), .B(n621), .ZN(Ciphertext[72]) );
  INV_X1 U27813 ( .A(n3114), .ZN(n27550) );
  AOI22_X1 U27814 ( .A1(n27551), .A2(n27552), .B1(n29085), .B2(n2433), .ZN(
        n27556) );
  INV_X1 U27815 ( .A(n27561), .ZN(n27575) );
  NOR2_X1 U27816 ( .A1(n27554), .A2(n27553), .ZN(n27555) );
  OAI22_X1 U27817 ( .A1(n27556), .A2(n27575), .B1(n27551), .B2(n27555), .ZN(
        n27558) );
  INV_X1 U27818 ( .A(n3049), .ZN(n27557) );
  XNOR2_X1 U27819 ( .A(n27558), .B(n27557), .ZN(Ciphertext[78]) );
  AOI21_X1 U27820 ( .B1(n27571), .B2(n27551), .A(n27576), .ZN(n27566) );
  NOR2_X1 U27821 ( .A1(n27571), .A2(n27573), .ZN(n27577) );
  AOI21_X1 U27822 ( .B1(n27577), .B2(n29158), .A(n3087), .ZN(n27559) );
  NAND2_X1 U27823 ( .A1(n27566), .A2(n27559), .ZN(n27570) );
  AND3_X1 U27824 ( .A1(n27562), .A2(n27561), .A3(n27560), .ZN(n27565) );
  NAND2_X1 U27825 ( .A1(n27562), .A2(n3087), .ZN(n27563) );
  NAND2_X1 U27826 ( .A1(n27577), .A2(n27563), .ZN(n27564) );
  OAI21_X1 U27827 ( .B1(n27577), .B2(n27565), .A(n27564), .ZN(n27569) );
  INV_X1 U27828 ( .A(n27566), .ZN(n27568) );
  NOR2_X1 U27829 ( .A1(n27551), .A2(n27571), .ZN(n27574) );
  OAI21_X1 U27830 ( .B1(n27574), .B2(n29578), .A(n29085), .ZN(n27579) );
  OAI21_X1 U27831 ( .B1(n27577), .B2(n27576), .A(n27575), .ZN(n27578) );
  NAND2_X1 U27832 ( .A1(n27578), .A2(n27579), .ZN(n27581) );
  INV_X1 U27833 ( .A(n2602), .ZN(n27580) );
  XNOR2_X1 U27834 ( .A(n27581), .B(n27580), .ZN(Ciphertext[83]) );
  OAI21_X1 U27835 ( .B1(n1901), .B2(n27585), .A(n27589), .ZN(n27583) );
  OAI21_X1 U27836 ( .B1(n27598), .B2(n27592), .A(n27583), .ZN(n27584) );
  XNOR2_X1 U27837 ( .A(n27584), .B(n22534), .ZN(Ciphertext[85]) );
  NOR2_X1 U27838 ( .A1(n930), .A2(n27593), .ZN(n27595) );
  OAI22_X1 U27839 ( .A1(n27598), .A2(n27597), .B1(n27596), .B2(n27595), .ZN(
        n27600) );
  INV_X1 U27840 ( .A(n28294), .ZN(n27599) );
  XNOR2_X1 U27841 ( .A(n27600), .B(n27599), .ZN(Ciphertext[89]) );
  NAND2_X1 U27842 ( .A1(n27601), .A2(n27625), .ZN(n27604) );
  NOR2_X1 U27843 ( .A1(n27628), .A2(n3366), .ZN(n27603) );
  NOR2_X1 U27844 ( .A1(n27627), .A2(n27625), .ZN(n27602) );
  XNOR2_X1 U27845 ( .A(n27606), .B(n27605), .ZN(Ciphertext[90]) );
  NAND2_X1 U27847 ( .A1(n27626), .A2(n27617), .ZN(n27608) );
  AOI22_X1 U27848 ( .A1(n27610), .A2(n28505), .B1(n27609), .B2(n27608), .ZN(
        n27612) );
  XNOR2_X1 U27849 ( .A(n27612), .B(n3035), .ZN(Ciphertext[91]) );
  MUX2_X1 U27850 ( .A(n27614), .B(n3366), .S(n27613), .Z(n27615) );
  XNOR2_X1 U27852 ( .A(n27625), .B(n28213), .ZN(n27616) );
  NAND3_X1 U27853 ( .A1(n27619), .A2(n27617), .A3(n3154), .ZN(n27621) );
  NAND3_X1 U27854 ( .A1(n27619), .A2(n28213), .A3(n27628), .ZN(n27620) );
  NOR3_X1 U27855 ( .A1(n27624), .A2(n27623), .A3(n27622), .ZN(Ciphertext[92])
         );
  NAND2_X1 U27856 ( .A1(n1912), .A2(n27628), .ZN(n27631) );
  INV_X1 U27857 ( .A(n3334), .ZN(n27633) );
  XNOR2_X1 U27858 ( .A(n27634), .B(n27633), .ZN(Ciphertext[94]) );
  MUX2_X1 U27859 ( .A(n27637), .B(n27636), .S(n29532), .Z(n27642) );
  NAND2_X1 U27860 ( .A1(n27639), .A2(n27638), .ZN(n27647) );
  AOI21_X1 U27863 ( .B1(n27647), .B2(n28466), .A(n27645), .ZN(n27648) );
  AOI21_X1 U27864 ( .B1(n27650), .B2(n27649), .A(n27648), .ZN(n27651) );
  XNOR2_X1 U27865 ( .A(n27651), .B(n1887), .ZN(Ciphertext[101]) );
  INV_X1 U27866 ( .A(n27652), .ZN(n27655) );
  AOI22_X1 U27867 ( .A1(n27674), .A2(n27663), .B1(n27672), .B2(n27671), .ZN(
        n27677) );
  INV_X1 U27868 ( .A(n29091), .ZN(n27653) );
  OAI21_X1 U27869 ( .B1(n27655), .B2(n27677), .A(n27654), .ZN(n27657) );
  XNOR2_X1 U27870 ( .A(n27657), .B(n27656), .ZN(Ciphertext[103]) );
  MUX2_X1 U27871 ( .A(n29091), .B(n28655), .S(n27661), .Z(n27659) );
  MUX2_X1 U27872 ( .A(n27659), .B(n27658), .S(n27663), .Z(n27660) );
  XNOR2_X1 U27873 ( .A(n27660), .B(n4503), .ZN(Ciphertext[104]) );
  XNOR2_X1 U27877 ( .A(n27670), .B(n27669), .ZN(Ciphertext[106]) );
  AOI21_X1 U27878 ( .B1(n29090), .B2(n27672), .A(n85), .ZN(n27675) );
  OAI22_X1 U27879 ( .A1(n27677), .A2(n27676), .B1(n27675), .B2(n27674), .ZN(
        n27679) );
  XNOR2_X1 U27880 ( .A(n27679), .B(n27678), .ZN(Ciphertext[107]) );
  NOR2_X1 U27882 ( .A1(n27714), .A2(n27725), .ZN(n27680) );
  NAND2_X1 U27883 ( .A1(n1826), .A2(n27680), .ZN(n27683) );
  OAI21_X1 U27884 ( .B1(n27681), .B2(n27711), .A(n27725), .ZN(n27682) );
  OAI211_X1 U27885 ( .C1(n27727), .C2(n27684), .A(n27683), .B(n27682), .ZN(
        n27686) );
  INV_X1 U27886 ( .A(n1246), .ZN(n27685) );
  XNOR2_X1 U27887 ( .A(n27686), .B(n27685), .ZN(Ciphertext[108]) );
  INV_X1 U27888 ( .A(n27707), .ZN(n27689) );
  NAND2_X1 U27889 ( .A1(n27689), .A2(n27687), .ZN(n27693) );
  NAND3_X1 U27890 ( .A1(n27690), .A2(n27689), .A3(n27688), .ZN(n27692) );
  AOI21_X1 U27891 ( .B1(n27693), .B2(n27692), .A(n27691), .ZN(n27695) );
  INV_X1 U27892 ( .A(n27711), .ZN(n27723) );
  NOR2_X1 U27893 ( .A1(n27695), .A2(n27694), .ZN(n27729) );
  NOR2_X1 U27894 ( .A1(n27727), .A2(n326), .ZN(n27697) );
  OAI21_X1 U27895 ( .B1(n28396), .B2(n27697), .A(n27696), .ZN(n27698) );
  XNOR2_X1 U27896 ( .A(n27698), .B(n22755), .ZN(Ciphertext[109]) );
  NOR2_X1 U27897 ( .A1(n27701), .A2(n27704), .ZN(n27699) );
  AOI211_X1 U27898 ( .C1(n27701), .C2(n27700), .A(n27702), .B(n27699), .ZN(
        n27709) );
  NAND2_X1 U27899 ( .A1(n27703), .A2(n27702), .ZN(n27705) );
  NOR2_X1 U27900 ( .A1(n27705), .A2(n27704), .ZN(n27706) );
  OR2_X1 U27901 ( .A1(n27707), .A2(n27706), .ZN(n27708) );
  NOR2_X1 U27902 ( .A1(n27709), .A2(n27708), .ZN(n27716) );
  INV_X1 U27905 ( .A(n27725), .ZN(n27712) );
  NAND2_X1 U27906 ( .A1(n27713), .A2(n27712), .ZN(n27721) );
  NAND3_X1 U27907 ( .A1(n27715), .A2(n27714), .A3(n27725), .ZN(n27720) );
  INV_X1 U27908 ( .A(n27716), .ZN(n27717) );
  NAND3_X1 U27909 ( .A1(n1826), .A2(n324), .A3(n27717), .ZN(n27719) );
  XNOR2_X1 U27911 ( .A(n27722), .B(n3062), .ZN(Ciphertext[110]) );
  AOI21_X1 U27912 ( .B1(n27725), .B2(n27724), .A(n27723), .ZN(n27726) );
  OAI22_X1 U27913 ( .A1(n27729), .A2(n1826), .B1(n27727), .B2(n27726), .ZN(
        n27731) );
  XNOR2_X1 U27914 ( .A(n27731), .B(n27730), .ZN(Ciphertext[113]) );
  INV_X1 U27915 ( .A(n29049), .ZN(n27746) );
  AOI21_X1 U27916 ( .B1(n27739), .B2(n28430), .A(n27744), .ZN(n27736) );
  NOR2_X1 U27917 ( .A1(n27745), .A2(n29049), .ZN(n27734) );
  NOR2_X1 U27918 ( .A1(n27739), .A2(n27732), .ZN(n27733) );
  XNOR2_X1 U27919 ( .A(n27738), .B(n27737), .ZN(Ciphertext[114]) );
  OR2_X1 U27920 ( .A1(n29049), .A2(n27755), .ZN(n27741) );
  NOR2_X1 U27921 ( .A1(n27739), .A2(n28430), .ZN(n27740) );
  AOI22_X1 U27922 ( .A1(n27755), .A2(n27744), .B1(n27759), .B2(n397), .ZN(
        n27758) );
  XNOR2_X1 U27923 ( .A(n27743), .B(n27742), .ZN(Ciphertext[115]) );
  NOR2_X1 U27924 ( .A1(n27745), .A2(n27744), .ZN(n27747) );
  OAI22_X1 U27925 ( .A1(n27747), .A2(n27759), .B1(n27746), .B2(n28445), .ZN(
        n27752) );
  NOR3_X1 U27926 ( .A1(n27757), .A2(n27749), .A3(n397), .ZN(n27751) );
  NOR2_X1 U27927 ( .A1(n28445), .A2(n397), .ZN(n27748) );
  OAI211_X1 U27928 ( .C1(n27757), .C2(n27749), .A(n27748), .B(n29049), .ZN(
        n27750) );
  AOI21_X1 U27931 ( .B1(n29049), .B2(n27755), .A(n28445), .ZN(n27760) );
  OAI22_X1 U27932 ( .A1(n27760), .A2(n27759), .B1(n27758), .B2(n27757), .ZN(
        n27761) );
  XNOR2_X1 U27933 ( .A(n27761), .B(n4882), .ZN(Ciphertext[119]) );
  OAI211_X1 U27935 ( .C1(n29027), .C2(n29537), .A(n29070), .B(n29118), .ZN(
        n27765) );
  INV_X1 U27936 ( .A(n27784), .ZN(n27764) );
  NOR2_X1 U27937 ( .A1(n28414), .A2(n29117), .ZN(n27785) );
  XNOR2_X1 U27938 ( .A(n27767), .B(n27766), .ZN(Ciphertext[121]) );
  OAI211_X1 U27939 ( .C1(n27777), .C2(n27776), .A(n27775), .B(n27774), .ZN(
        n27779) );
  XNOR2_X1 U27940 ( .A(n27779), .B(n27778), .ZN(Ciphertext[124]) );
  OAI21_X1 U27941 ( .B1(n27782), .B2(n28414), .A(n27780), .ZN(n27787) );
  OAI21_X1 U27942 ( .B1(n27785), .B2(n27784), .A(n29027), .ZN(n27786) );
  NAND2_X1 U27943 ( .A1(n27787), .A2(n27786), .ZN(n27789) );
  XNOR2_X1 U27944 ( .A(n27789), .B(n27788), .ZN(Ciphertext[125]) );
  NAND2_X1 U27946 ( .A1(n27790), .A2(n27817), .ZN(n27793) );
  OAI211_X1 U27947 ( .C1(n27800), .C2(n29535), .A(n27793), .B(n27792), .ZN(
        n27794) );
  XNOR2_X1 U27948 ( .A(n27794), .B(n4070), .ZN(Ciphertext[126]) );
  NAND2_X1 U27949 ( .A1(n28403), .A2(n3380), .ZN(n27799) );
  AND2_X1 U27950 ( .A1(n27817), .A2(n3380), .ZN(n27806) );
  OAI21_X1 U27951 ( .B1(n27795), .B2(n3380), .A(n27807), .ZN(n27796) );
  AOI21_X1 U27952 ( .B1(n27812), .B2(n27806), .A(n27796), .ZN(n27798) );
  NAND2_X1 U27953 ( .A1(n27800), .A2(n27811), .ZN(n27797) );
  OAI211_X1 U27954 ( .C1(n27800), .C2(n27799), .A(n27798), .B(n27797), .ZN(
        n27816) );
  NAND2_X1 U27955 ( .A1(n29469), .A2(n27811), .ZN(n27805) );
  AOI21_X1 U27956 ( .B1(n27819), .B2(n3380), .A(n27807), .ZN(n27804) );
  NAND2_X1 U27957 ( .A1(n27818), .A2(n27811), .ZN(n27802) );
  NAND2_X1 U27958 ( .A1(n27802), .A2(n27817), .ZN(n27803) );
  OAI211_X1 U27959 ( .C1(n27819), .C2(n27805), .A(n27804), .B(n27803), .ZN(
        n27815) );
  INV_X1 U27960 ( .A(n27806), .ZN(n27808) );
  NOR3_X1 U27961 ( .A1(n27808), .A2(n27818), .A3(n27807), .ZN(n27809) );
  NAND2_X1 U27962 ( .A1(n29535), .A2(n27809), .ZN(n27814) );
  NAND3_X1 U27963 ( .A1(n27812), .A2(n27811), .A3(n27817), .ZN(n27813) );
  NAND4_X1 U27964 ( .A1(n27816), .A2(n27815), .A3(n27814), .A4(n27813), .ZN(
        Ciphertext[130]) );
  OAI21_X1 U27965 ( .B1(n27819), .B2(n27818), .A(n27817), .ZN(n27820) );
  AOI22_X1 U27966 ( .A1(n27823), .A2(n27822), .B1(n27821), .B2(n27820), .ZN(
        n27824) );
  XNOR2_X1 U27967 ( .A(n27824), .B(n3463), .ZN(Ciphertext[131]) );
  INV_X1 U27968 ( .A(n27829), .ZN(n27833) );
  INV_X1 U27969 ( .A(n27830), .ZN(n27832) );
  NAND4_X1 U27970 ( .A1(n27834), .A2(n27833), .A3(n27832), .A4(n27831), .ZN(
        n27845) );
  MUX2_X1 U27971 ( .A(n27898), .B(n27836), .S(n29575), .Z(n27837) );
  NOR2_X1 U27972 ( .A1(n27837), .A2(n5299), .ZN(n27840) );
  NOR3_X1 U27973 ( .A1(n27840), .A2(n27839), .A3(n27838), .ZN(n27842) );
  NAND2_X1 U27974 ( .A1(n27842), .A2(n27841), .ZN(n27844) );
  AOI21_X1 U27975 ( .B1(n27845), .B2(n27844), .A(n27843), .ZN(n27846) );
  NOR2_X1 U27976 ( .A1(n27851), .A2(n27852), .ZN(n27853) );
  AOI22_X1 U27977 ( .A1(n27855), .A2(n27853), .B1(n27859), .B2(n6949), .ZN(
        n27857) );
  OAI211_X1 U27978 ( .C1(n27859), .C2(n27858), .A(n27857), .B(n27856), .ZN(
        n27861) );
  INV_X1 U27979 ( .A(n3527), .ZN(n27860) );
  XNOR2_X1 U27980 ( .A(n27861), .B(n27860), .ZN(Ciphertext[141]) );
  AOI22_X1 U27981 ( .A1(n27875), .A2(n27864), .B1(n27862), .B2(n27863), .ZN(
        n27878) );
  NOR2_X1 U27982 ( .A1(n27875), .A2(n26540), .ZN(n27868) );
  NAND3_X1 U27983 ( .A1(n27872), .A2(n27871), .A3(n27866), .ZN(n27867) );
  OAI21_X1 U27984 ( .B1(n27878), .B2(n27868), .A(n27867), .ZN(n27870) );
  INV_X1 U27985 ( .A(n2987), .ZN(n27869) );
  XNOR2_X1 U27986 ( .A(n27870), .B(n27869), .ZN(Ciphertext[145]) );
  NOR2_X1 U27987 ( .A1(n27872), .A2(n27871), .ZN(n27874) );
  NOR2_X1 U27988 ( .A1(n27874), .A2(n27873), .ZN(n27876) );
  OAI22_X1 U27989 ( .A1(n27878), .A2(n27877), .B1(n27876), .B2(n27875), .ZN(
        n27880) );
  XNOR2_X1 U27990 ( .A(n27880), .B(n27879), .ZN(Ciphertext[149]) );
  NAND2_X1 U27991 ( .A1(n27919), .A2(n27080), .ZN(n27882) );
  OAI21_X1 U27992 ( .B1(n27905), .B2(n27908), .A(n27918), .ZN(n27881) );
  OAI21_X1 U27993 ( .B1(n27882), .B2(n27908), .A(n27881), .ZN(n27886) );
  NAND2_X1 U27994 ( .A1(n27908), .A2(n27923), .ZN(n27885) );
  INV_X1 U27995 ( .A(n27883), .ZN(n27884) );
  XNOR2_X1 U27996 ( .A(n27888), .B(n27887), .ZN(Ciphertext[152]) );
  INV_X1 U27997 ( .A(n27908), .ZN(n27909) );
  OAI21_X1 U27998 ( .B1(n27919), .B2(n27909), .A(n1843), .ZN(n27892) );
  NAND3_X1 U27999 ( .A1(n27918), .A2(n27908), .A3(n27905), .ZN(n27891) );
  NAND2_X1 U28000 ( .A1(n27889), .A2(n27920), .ZN(n27890) );
  OAI21_X1 U28004 ( .B1(n27060), .B2(n27898), .A(n28600), .ZN(n27901) );
  AOI211_X1 U28005 ( .C1(n27902), .C2(n27901), .A(n27900), .B(n27899), .ZN(
        n27907) );
  OAI21_X1 U28006 ( .B1(n27904), .B2(n27903), .A(n27060), .ZN(n27906) );
  INV_X1 U28007 ( .A(n27905), .ZN(n27917) );
  NAND3_X1 U28008 ( .A1(n27920), .A2(n27908), .A3(n1843), .ZN(n27912) );
  NAND3_X1 U28009 ( .A1(n27080), .A2(n27909), .A3(n27917), .ZN(n27911) );
  OAI211_X1 U28010 ( .C1(n27914), .C2(n1843), .A(n27912), .B(n27911), .ZN(
        n27916) );
  XNOR2_X1 U28011 ( .A(n27916), .B(n27915), .ZN(Ciphertext[154]) );
  OAI21_X1 U28012 ( .B1(n27919), .B2(n27918), .A(n27917), .ZN(n27922) );
  AOI22_X1 U28013 ( .A1(n27923), .A2(n27922), .B1(n27921), .B2(n27920), .ZN(
        n27924) );
  XNOR2_X1 U28014 ( .A(n27924), .B(n2510), .ZN(Ciphertext[155]) );
  INV_X1 U28015 ( .A(n27925), .ZN(n27950) );
  INV_X1 U28016 ( .A(n27934), .ZN(n27942) );
  OAI21_X1 U28018 ( .B1(n27948), .B2(n27927), .A(n27926), .ZN(n27929) );
  OAI211_X1 U28019 ( .C1(n27942), .C2(n28451), .A(n27929), .B(n27928), .ZN(
        n27931) );
  INV_X1 U28020 ( .A(n3317), .ZN(n27930) );
  XNOR2_X1 U28021 ( .A(n27931), .B(n27930), .ZN(Ciphertext[156]) );
  NOR2_X1 U28022 ( .A1(n27944), .A2(n27938), .ZN(n27947) );
  NOR2_X1 U28023 ( .A1(n27244), .A2(n27947), .ZN(n27935) );
  NAND2_X1 U28024 ( .A1(n27941), .A2(n28441), .ZN(n27932) );
  OAI21_X1 U28025 ( .B1(n27935), .B2(n27934), .A(n27933), .ZN(n27937) );
  XNOR2_X1 U28026 ( .A(n27937), .B(n27936), .ZN(Ciphertext[157]) );
  XNOR2_X1 U28027 ( .A(n27943), .B(n5802), .ZN(Ciphertext[159]) );
  AOI21_X1 U28028 ( .B1(n27926), .B2(n4998), .A(n27944), .ZN(n27951) );
  AOI22_X1 U28029 ( .A1(n27948), .A2(n27950), .B1(n27947), .B2(n28451), .ZN(
        n27949) );
  OAI21_X1 U28030 ( .B1(n27951), .B2(n27950), .A(n27949), .ZN(n27953) );
  XNOR2_X1 U28031 ( .A(n27953), .B(n27952), .ZN(Ciphertext[161]) );
  NOR2_X1 U28032 ( .A1(n27972), .A2(n27996), .ZN(n27965) );
  AND2_X1 U28034 ( .A1(n29021), .A2(n27977), .ZN(n27954) );
  INV_X1 U28035 ( .A(n27956), .ZN(n27957) );
  INV_X1 U28038 ( .A(n27997), .ZN(n27964) );
  OAI211_X1 U28040 ( .C1(n27964), .C2(n29092), .A(n27977), .B(n27979), .ZN(
        n27960) );
  OAI21_X1 U28041 ( .B1(n27998), .B2(n27965), .A(n27960), .ZN(n27962) );
  XNOR2_X1 U28042 ( .A(n27962), .B(n27961), .ZN(Ciphertext[163]) );
  MUX2_X1 U28043 ( .A(n27970), .B(n27977), .S(n27979), .Z(n27967) );
  INV_X1 U28044 ( .A(n27996), .ZN(n27983) );
  AND2_X1 U28045 ( .A1(n27977), .A2(n27972), .ZN(n27963) );
  AOI22_X1 U28046 ( .A1(n27965), .A2(n27964), .B1(n27963), .B2(n28456), .ZN(
        n27966) );
  OAI21_X1 U28047 ( .B1(n27967), .B2(n27983), .A(n27966), .ZN(n27969) );
  INV_X1 U28048 ( .A(n3211), .ZN(n27968) );
  XNOR2_X1 U28049 ( .A(n27969), .B(n27968), .ZN(Ciphertext[165]) );
  NOR2_X1 U28050 ( .A1(n28456), .A2(n27977), .ZN(n27987) );
  INV_X1 U28051 ( .A(n27987), .ZN(n27971) );
  NOR2_X1 U28052 ( .A1(n27971), .A2(n27970), .ZN(n27991) );
  AND2_X1 U28053 ( .A1(n27972), .A2(n3722), .ZN(n27976) );
  INV_X1 U28054 ( .A(n27976), .ZN(n27975) );
  AOI21_X1 U28055 ( .B1(n28636), .B2(n27978), .A(n27983), .ZN(n27974) );
  NAND2_X1 U28056 ( .A1(n29092), .A2(n27978), .ZN(n27985) );
  OAI211_X1 U28057 ( .C1(n28636), .C2(n27975), .A(n27974), .B(n27985), .ZN(
        n27990) );
  AND2_X1 U28058 ( .A1(n27987), .A2(n27976), .ZN(n27984) );
  NAND2_X1 U28059 ( .A1(n27977), .A2(n27978), .ZN(n27982) );
  XNOR2_X1 U28060 ( .A(n27979), .B(n27978), .ZN(n27980) );
  INV_X1 U28061 ( .A(n27985), .ZN(n27986) );
  NAND2_X1 U28062 ( .A1(n27987), .A2(n27986), .ZN(n27988) );
  OAI211_X1 U28063 ( .C1(n27991), .C2(n27990), .A(n27989), .B(n27988), .ZN(
        Ciphertext[166]) );
  AOI21_X1 U28064 ( .B1(n29021), .B2(n29063), .A(n28456), .ZN(n27995) );
  OAI22_X1 U28065 ( .A1(n27998), .A2(n28636), .B1(n27996), .B2(n27995), .ZN(
        n27999) );
  XNOR2_X1 U28066 ( .A(n27999), .B(n635), .ZN(Ciphertext[167]) );
  NAND3_X1 U28067 ( .A1(n445), .A2(n28003), .A3(n28015), .ZN(n28004) );
  INV_X1 U28068 ( .A(n28015), .ZN(n28008) );
  NAND3_X1 U28069 ( .A1(n28411), .A2(n28008), .A3(n26984), .ZN(n28011) );
  NAND2_X1 U28070 ( .A1(n6955), .A2(n443), .ZN(n28010) );
  XNOR2_X1 U28071 ( .A(n28014), .B(n28013), .ZN(Ciphertext[172]) );
  NAND2_X1 U28072 ( .A1(n28017), .A2(n28016), .ZN(n28018) );
  NAND2_X1 U28073 ( .A1(n28008), .A2(n28018), .ZN(n28020) );
  AOI22_X1 U28074 ( .A1(n28022), .A2(n28021), .B1(n28020), .B2(n28019), .ZN(
        n28023) );
  XNOR2_X1 U28075 ( .A(n28023), .B(n3323), .ZN(Ciphertext[173]) );
  AOI22_X1 U28076 ( .A1(n28030), .A2(n28028), .B1(n28034), .B2(n28027), .ZN(
        n28029) );
  OAI21_X1 U28077 ( .B1(n28031), .B2(n28030), .A(n28029), .ZN(n28033) );
  INV_X1 U28078 ( .A(n3695), .ZN(n28032) );
  XNOR2_X1 U28079 ( .A(n28033), .B(n28032), .ZN(Ciphertext[174]) );
  NOR3_X1 U28080 ( .A1(n28040), .A2(n28039), .A3(n28038), .ZN(n28041) );
  NOR2_X1 U28081 ( .A1(n28042), .A2(n28041), .ZN(n28043) );
  XNOR2_X1 U28082 ( .A(n28043), .B(n4501), .ZN(Ciphertext[176]) );
  NOR2_X1 U28083 ( .A1(n28044), .A2(n28543), .ZN(n28046) );
  INV_X1 U28084 ( .A(n28067), .ZN(n28045) );
  OAI21_X1 U28085 ( .B1(n28055), .B2(n28046), .A(n28045), .ZN(n28049) );
  OAI21_X1 U28086 ( .B1(n28047), .B2(n28065), .A(n28543), .ZN(n28048) );
  NAND2_X1 U28087 ( .A1(n28049), .A2(n28048), .ZN(n28051) );
  XNOR2_X1 U28088 ( .A(n28051), .B(n28050), .ZN(Ciphertext[180]) );
  NOR2_X1 U28089 ( .A1(n28052), .A2(n28063), .ZN(n28056) );
  OAI21_X1 U28090 ( .B1(n28067), .B2(n28063), .A(n28053), .ZN(n28054) );
  OAI21_X1 U28091 ( .B1(n28056), .B2(n28055), .A(n28054), .ZN(n28058) );
  INV_X1 U28092 ( .A(n3650), .ZN(n28057) );
  XNOR2_X1 U28093 ( .A(n28058), .B(n28057), .ZN(Ciphertext[181]) );
  MUX2_X1 U28094 ( .A(n28067), .B(n28543), .S(n28069), .Z(n28060) );
  MUX2_X1 U28095 ( .A(n28060), .B(n28059), .S(n28063), .Z(n28062) );
  INV_X1 U28096 ( .A(n2505), .ZN(n28061) );
  XNOR2_X1 U28097 ( .A(n28062), .B(n28061), .ZN(Ciphertext[182]) );
  INV_X1 U28098 ( .A(n28063), .ZN(n28068) );
  MUX2_X1 U28099 ( .A(n28069), .B(n28068), .S(n28543), .Z(n28072) );
  OR2_X1 U28100 ( .A1(n28066), .A2(n28065), .ZN(n28070) );
  XNOR2_X1 U28101 ( .A(n28074), .B(n28073), .ZN(Ciphertext[184]) );
  INV_X1 U28103 ( .A(n28115), .ZN(n28075) );
  OAI211_X1 U28104 ( .C1(n28075), .C2(n29121), .A(n28089), .B(n28090), .ZN(
        n28076) );
  INV_X1 U28106 ( .A(n3015), .ZN(n28078) );
  XNOR2_X1 U28107 ( .A(n28079), .B(n28078), .ZN(Ciphertext[187]) );
  NAND2_X1 U28109 ( .A1(n28590), .A2(n28794), .ZN(n28081) );
  OAI21_X1 U28111 ( .B1(n29480), .B2(n28081), .A(n28080), .ZN(n28087) );
  NAND2_X1 U28112 ( .A1(n28090), .A2(n28794), .ZN(n28084) );
  NAND3_X1 U28113 ( .A1(n28111), .A2(n28090), .A3(n29121), .ZN(n28083) );
  OAI211_X1 U28114 ( .C1(n28107), .C2(n28084), .A(n1928), .B(n28083), .ZN(
        n28086) );
  NOR2_X1 U28115 ( .A1(n28111), .A2(n28794), .ZN(n28105) );
  AND2_X1 U28116 ( .A1(n28087), .A2(n4359), .ZN(n28088) );
  NAND2_X1 U28117 ( .A1(n29056), .A2(n28089), .ZN(n28096) );
  NOR3_X1 U28118 ( .A1(n28107), .A2(n28089), .A3(n28794), .ZN(n28093) );
  AND3_X1 U28119 ( .A1(n28111), .A2(n28794), .A3(n28090), .ZN(n28092) );
  NOR2_X1 U28120 ( .A1(n28093), .A2(n28092), .ZN(n28095) );
  AOI21_X1 U28122 ( .B1(n29056), .B2(n28112), .A(n28111), .ZN(n28114) );
  INV_X1 U28123 ( .A(n2446), .ZN(n28116) );
  NAND2_X2 U6151 ( .A1(n5663), .A2(n5665), .ZN(n22434) );
  XNOR2_X2 U3467 ( .A(Key[105]), .B(Plaintext[105]), .ZN(n8231) );
  OAI21_X2 U2036 ( .B1(n6976), .B2(n8231), .A(n6975), .ZN(n5945) );
  BUF_X1 U1808 ( .A(n7560), .Z(n8044) );
  NOR2_X2 U5612 ( .A1(n26355), .A2(n26354), .ZN(n1912) );
  INV_X1 U14802 ( .A(n7198), .ZN(n8281) );
  XNOR2_X2 U3188 ( .A(n9769), .B(n9768), .ZN(n3441) );
  OAI211_X2 U1772 ( .C1(n20932), .C2(n20931), .A(n20930), .B(n20929), .ZN(
        n22094) );
  XNOR2_X2 U14624 ( .A(n7077), .B(Key[185]), .ZN(n7093) );
  BUF_X1 U775 ( .A(n24205), .Z(n24814) );
  XNOR2_X1 U1023 ( .A(n15043), .B(n15044), .ZN(n337) );
  NOR2_X1 U10135 ( .A1(n3991), .A2(n10050), .ZN(n11855) );
  XNOR2_X2 U2015 ( .A(n4506), .B(n4505), .ZN(n11209) );
  AND2_X2 U2541 ( .A1(n20402), .A2(n5871), .ZN(n21539) );
  NOR2_X2 U1999 ( .A1(n11405), .A2(n11403), .ZN(n11848) );
  OAI21_X1 U1253 ( .B1(n11952), .B2(n11665), .A(n5901), .ZN(n11668) );
  NAND3_X2 U3263 ( .A1(n3296), .A2(n8406), .A3(n8405), .ZN(n10128) );
  NAND3_X2 U2202 ( .A1(n24884), .A2(n2615), .A3(n1995), .ZN(n27638) );
  OAI21_X1 U462 ( .B1(n11784), .B2(n666), .A(n667), .ZN(n12542) );
  OAI21_X2 U2363 ( .B1(n23574), .B2(n23573), .A(n23572), .ZN(n24760) );
  AND3_X2 U1864 ( .A1(n873), .A2(n5350), .A3(n5348), .ZN(n25681) );
  NAND2_X2 U21 ( .A1(n24090), .A2(n24091), .ZN(n24471) );
  BUF_X1 U27204 ( .A(n26539), .Z(n27864) );
  MUX2_X2 U1879 ( .A(n23249), .B(n23248), .S(n23247), .Z(n24367) );
  XNOR2_X1 U248 ( .A(n24301), .B(n24302), .ZN(n26191) );
  XNOR2_X2 U4391 ( .A(n19204), .B(n19205), .ZN(n20349) );
  INV_X1 U445 ( .A(n17780), .ZN(n18168) );
  XNOR2_X2 U20591 ( .A(n16276), .B(n16275), .ZN(n17148) );
  BUF_X1 U2038 ( .A(n7371), .Z(n8222) );
  XNOR2_X1 U12034 ( .A(n4753), .B(n16342), .ZN(n17179) );
  AOI22_X1 U219 ( .A1(n28807), .A2(n125), .B1(n11611), .B2(n11767), .ZN(n12548) );
  CLKBUF_X1 U2052 ( .A(Key[92]), .Z(n3164) );
  CLKBUF_X1 U3493 ( .A(Key[158]), .Z(n3644) );
  CLKBUF_X1 U3450 ( .A(Key[111]), .Z(n26909) );
  CLKBUF_X1 U113 ( .A(Key[125]), .Z(n2946) );
  XNOR2_X1 U821 ( .A(Key[28]), .B(Plaintext[28]), .ZN(n8151) );
  CLKBUF_X1 U642 ( .A(Key[138]), .Z(n2403) );
  CLKBUF_X1 U1045 ( .A(Key[152]), .Z(n3527) );
  CLKBUF_X1 U3483 ( .A(Key[77]), .Z(n2961) );
  CLKBUF_X1 U228 ( .A(Key[99]), .Z(n2527) );
  CLKBUF_X1 U115 ( .A(Key[95]), .Z(n72) );
  XNOR2_X1 U14797 ( .A(Key[138]), .B(Plaintext[138]), .ZN(n8275) );
  AND2_X1 U846 ( .A1(n7857), .A2(n7858), .ZN(n9015) );
  NAND3_X1 U3381 ( .A1(n7323), .A2(n7280), .A3(n2716), .ZN(n8889) );
  OAI211_X1 U6648 ( .C1(n5559), .C2(n5558), .A(n7305), .B(n7304), .ZN(n9421)
         );
  NAND2_X1 U8556 ( .A1(n7246), .A2(n2470), .ZN(n8749) );
  OAI211_X1 U1321 ( .C1(n7967), .C2(n7188), .A(n7962), .B(n5470), .ZN(n8809)
         );
  OAI211_X1 U4350 ( .C1(n4939), .C2(n1700), .A(n1404), .B(n7091), .ZN(n8586)
         );
  NAND2_X1 U423 ( .A1(n7078), .A2(n2507), .ZN(n8521) );
  INV_X1 U6673 ( .A(n8589), .ZN(n8594) );
  NAND2_X1 U2032 ( .A1(n6382), .A2(n6381), .ZN(n8610) );
  NAND2_X1 U391 ( .A1(n2388), .A2(n2080), .ZN(n9202) );
  OR2_X1 U1191 ( .A1(n8439), .A2(n8720), .ZN(n224) );
  BUF_X1 U715 ( .A(n8230), .Z(n8961) );
  BUF_X1 U16085 ( .A(n9306), .Z(n9725) );
  AND3_X1 U889 ( .A1(n9365), .A2(n3273), .A3(n3272), .ZN(n10352) );
  NAND3_X1 U3264 ( .A1(n1118), .A2(n9048), .A3(n1117), .ZN(n10435) );
  NAND2_X1 U3258 ( .A1(n8083), .A2(n8082), .ZN(n10289) );
  XNOR2_X1 U3233 ( .A(n10262), .B(n10261), .ZN(n10876) );
  XNOR2_X1 U10153 ( .A(n9554), .B(n9553), .ZN(n11275) );
  XNOR2_X1 U4315 ( .A(n5185), .B(n10058), .ZN(n11154) );
  XNOR2_X1 U15875 ( .A(n8922), .B(n8923), .ZN(n10810) );
  NAND4_X1 U469 ( .A1(n4146), .A2(n10527), .A3(n10526), .A4(n10838), .ZN(
        n11747) );
  AND3_X1 U940 ( .A1(n11080), .A2(n11079), .A3(n11078), .ZN(n12270) );
  AOI21_X1 U408 ( .B1(n10807), .B2(n7814), .A(n6347), .ZN(n12145) );
  NAND2_X1 U783 ( .A1(n139), .A2(n5902), .ZN(n11951) );
  INV_X1 U2007 ( .A(n11473), .ZN(n431) );
  OR2_X1 U3073 ( .A1(n12148), .A2(n5636), .ZN(n12559) );
  XNOR2_X1 U233 ( .A(n12854), .B(n13484), .ZN(n13347) );
  XNOR2_X1 U18835 ( .A(n13477), .B(n13476), .ZN(n13719) );
  XNOR2_X1 U3028 ( .A(n11511), .B(n11510), .ZN(n14240) );
  XNOR2_X1 U17990 ( .A(n12393), .B(n12392), .ZN(n14406) );
  INV_X1 U282 ( .A(n12607), .ZN(n14294) );
  OR2_X1 U854 ( .A1(n14165), .A2(n14484), .ZN(n14483) );
  NOR2_X1 U404 ( .A1(n14483), .A2(n14164), .ZN(n14660) );
  NOR2_X1 U10190 ( .A1(n14290), .A2(n14289), .ZN(n15054) );
  NAND3_X1 U2968 ( .A1(n6234), .A2(n6235), .A3(n6233), .ZN(n15370) );
  BUF_X1 U836 ( .A(n14600), .Z(n14845) );
  MUX2_X1 U1347 ( .A(n13940), .B(n13939), .S(n14253), .Z(n15300) );
  AOI22_X1 U5630 ( .A1(n13960), .A2(n13959), .B1(n13961), .B2(n14437), .ZN(
        n15323) );
  NAND3_X1 U186 ( .A1(n2742), .A2(n2745), .A3(n2743), .ZN(n15790) );
  AND3_X1 U342 ( .A1(n36), .A2(n5093), .A3(n5092), .ZN(n16393) );
  XNOR2_X1 U973 ( .A(n15604), .B(n15603), .ZN(n17386) );
  XNOR2_X1 U474 ( .A(n4215), .B(n15614), .ZN(n16878) );
  XNOR2_X1 U10808 ( .A(n3677), .B(n5828), .ZN(n17261) );
  XNOR2_X1 U19212 ( .A(n14028), .B(n14027), .ZN(n17428) );
  XNOR2_X1 U567 ( .A(n15573), .B(n15574), .ZN(n17155) );
  BUF_X1 U511 ( .A(n17255), .Z(n1880) );
  AND3_X2 U241 ( .A1(n6800), .A2(n6799), .A3(n5986), .ZN(n18506) );
  CLKBUF_X1 U14303 ( .A(n16693), .Z(n17948) );
  BUF_X2 U2735 ( .A(n16685), .Z(n514) );
  BUF_X1 U904 ( .A(n15810), .Z(n18064) );
  NAND3_X1 U1090 ( .A1(n1480), .A2(n4244), .A3(n4191), .ZN(n19534) );
  AND3_X1 U40 ( .A1(n1170), .A2(n3933), .A3(n3931), .ZN(n19243) );
  AOI22_X1 U8922 ( .A1(n17748), .A2(n3239), .B1(n17747), .B2(n18195), .ZN(
        n18856) );
  OAI211_X1 U5418 ( .C1(n1759), .C2(n1758), .A(n17247), .B(n4761), .ZN(n19246)
         );
  NAND4_X1 U9607 ( .A1(n17578), .A2(n3086), .A3(n3085), .A4(n3084), .ZN(n19373) );
  AOI22_X1 U609 ( .A1(n18103), .A2(n18104), .B1(n1143), .B2(n106), .ZN(n19004)
         );
  NAND2_X1 U1323 ( .A1(n6342), .A2(n16873), .ZN(n19686) );
  AND2_X1 U2639 ( .A1(n5492), .A2(n19172), .ZN(n19692) );
  INV_X1 U2652 ( .A(n19245), .ZN(n19348) );
  XNOR2_X1 U1563 ( .A(n4339), .B(n18086), .ZN(n20205) );
  AOI21_X1 U1149 ( .B1(n6261), .B2(n20546), .A(n19958), .ZN(n20392) );
  NAND2_X1 U1550 ( .A1(n3473), .A2(n19821), .ZN(n21495) );
  AOI21_X1 U1289 ( .B1(n20195), .B2(n20821), .A(n20824), .ZN(n21677) );
  AND2_X1 U1381 ( .A1(n20891), .A2(n20890), .ZN(n21087) );
  OR2_X1 U2542 ( .A1(n2529), .A2(n2528), .ZN(n20688) );
  NAND3_X1 U12584 ( .A1(n5252), .A2(n19881), .A3(n5253), .ZN(n21713) );
  OAI22_X1 U883 ( .A1(n28797), .A2(n21039), .B1(n21038), .B2(n21037), .ZN(
        n21903) );
  AND3_X1 U2485 ( .A1(n1940), .A2(n2041), .A3(n1948), .ZN(n22194) );
  AND3_X1 U881 ( .A1(n658), .A2(n5128), .A3(n656), .ZN(n22898) );
  XNOR2_X1 U6159 ( .A(n22643), .B(n22898), .ZN(n22481) );
  XNOR2_X1 U1669 ( .A(n20708), .B(n20709), .ZN(n23351) );
  OAI21_X1 U197 ( .B1(n23401), .B2(n23402), .A(n23400), .ZN(n24077) );
  MUX2_X1 U14074 ( .A(n24158), .B(n24157), .S(n28512), .Z(n26041) );
  AND3_X1 U12962 ( .A1(n5654), .A2(n5655), .A3(n5653), .ZN(n25714) );
  XNOR2_X1 U519 ( .A(n5755), .B(n5754), .ZN(n27700) );
  XNOR2_X1 U13844 ( .A(n25058), .B(n25057), .ZN(n26172) );
  BUF_X1 U5574 ( .A(n26436), .Z(n26940) );
  NAND4_X1 U8458 ( .A1(n27135), .A2(n27134), .A3(n27133), .A4(n27132), .ZN(
        n27744) );
  AND2_X1 U1358 ( .A1(n26521), .A2(n26520), .ZN(n26641) );
  AND2_X1 U1384 ( .A1(n3376), .A2(n3397), .ZN(n27591) );
  AND3_X1 U970 ( .A1(n26486), .A2(n26488), .A3(n26487), .ZN(n27427) );
  NOR2_X1 U853 ( .A1(n27877), .A2(n26539), .ZN(n27313) );
  CLKBUF_X1 U3484 ( .A(Key[1]), .Z(n27462) );
  CLKBUF_X1 U3456 ( .A(Key[117]), .Z(n3385) );
  CLKBUF_X1 U760 ( .A(Key[166]), .Z(n135) );
  NOR2_X1 U5163 ( .A1(n9184), .A2(n9007), .ZN(n2250) );
  INV_X1 U3364 ( .A(n9425), .ZN(n604) );
  AND2_X1 U661 ( .A1(n8109), .A2(n9041), .ZN(n9042) );
  AND2_X1 U8339 ( .A1(n7490), .A2(n9084), .ZN(n8724) );
  NAND2_X1 U999 ( .A1(n8483), .A2(n8484), .ZN(n10250) );
  INV_X1 U3239 ( .A(n11000), .ZN(n592) );
  INV_X1 U2014 ( .A(n10687), .ZN(n10959) );
  CLKBUF_X1 U1106 ( .A(n10668), .Z(n11048) );
  AND2_X1 U10428 ( .A1(n11881), .A2(n11875), .ZN(n11883) );
  AOI22_X1 U1362 ( .A1(n2430), .A2(n10870), .B1(n1630), .B2(n11883), .ZN(
        n13195) );
  NAND3_X1 U4337 ( .A1(n3020), .A2(n3021), .A3(n11513), .ZN(n13137) );
  INV_X1 U19201 ( .A(n14132), .ZN(n14341) );
  INV_X1 U11243 ( .A(n5584), .ZN(n14411) );
  INV_X1 U13346 ( .A(n13920), .ZN(n14033) );
  BUF_X1 U612 ( .A(n13677), .Z(n14466) );
  OAI21_X1 U1457 ( .B1(n13813), .B2(n14411), .A(n5542), .ZN(n14904) );
  NAND3_X1 U744 ( .A1(n6433), .A2(n13712), .A3(n13713), .ZN(n15135) );
  INV_X1 U1963 ( .A(n17389), .ZN(n424) );
  BUF_X1 U20851 ( .A(n16712), .Z(n17379) );
  NOR2_X1 U10285 ( .A1(n16803), .A2(n17474), .ZN(n17475) );
  AND3_X1 U536 ( .A1(n16972), .A2(n16971), .A3(n17267), .ZN(n18285) );
  INV_X1 U6061 ( .A(n18476), .ZN(n18480) );
  OAI211_X1 U4403 ( .C1(n17950), .C2(n17906), .A(n17949), .B(n6387), .ZN(
        n19622) );
  OAI211_X1 U2670 ( .C1(n18423), .C2(n18044), .A(n5496), .B(n5495), .ZN(n19389) );
  OR2_X1 U2492 ( .A1(n21227), .A2(n21632), .ZN(n21036) );
  INV_X1 U8131 ( .A(n23789), .ZN(n23792) );
  OR2_X1 U1118 ( .A1(n23375), .A2(n24072), .ZN(n205) );
  OR2_X1 U155 ( .A1(n23916), .A2(n23917), .ZN(n985) );
  XNOR2_X1 U26486 ( .A(n25554), .B(n25553), .ZN(n27044) );
  XNOR2_X1 U4317 ( .A(n25496), .B(n25497), .ZN(n27013) );
  NAND2_X1 U14388 ( .A1(n26623), .A2(n27013), .ZN(n26624) );
  AOI22_X1 U26586 ( .A1(n26217), .A2(n28459), .B1(n26210), .B2(n25661), .ZN(
        n25664) );
  AND2_X2 U11169 ( .A1(n3928), .A2(n3927), .ZN(n15343) );
  OR2_X2 U9574 ( .A1(n7699), .A2(n7698), .ZN(n9034) );
  AND3_X2 U4450 ( .A1(n3709), .A2(n3823), .A3(n3825), .ZN(n19228) );
  OR2_X2 U3816 ( .A1(n24336), .A2(n24337), .ZN(n24341) );
  BUF_X2 U624 ( .A(n14061), .Z(n14064) );
  OR2_X2 U708 ( .A1(n8172), .A2(n8171), .ZN(n8984) );
  BUF_X2 U2251 ( .A(n26518), .Z(n27138) );
  MUX2_X2 U1333 ( .A(n15450), .B(n15449), .S(n15448), .Z(n16557) );
  OR2_X2 U779 ( .A1(n19918), .A2(n19917), .ZN(n21875) );
  AND2_X2 U543 ( .A1(n4209), .A2(n3402), .ZN(n18913) );
  AND3_X2 U11200 ( .A1(n3956), .A2(n3960), .A3(n3955), .ZN(n13175) );
  OAI21_X2 U11407 ( .B1(n10862), .B2(n11512), .A(n4140), .ZN(n12566) );
  AND3_X2 U13213 ( .A1(n5906), .A2(n5908), .A3(n5907), .ZN(n19251) );
  AOI21_X2 U17368 ( .B1(n11327), .B2(n11328), .A(n11326), .ZN(n11801) );
  XNOR2_X2 U4110 ( .A(n19515), .B(n19514), .ZN(n20299) );
  OAI211_X2 U72 ( .C1(n15507), .C2(n15506), .A(n15505), .B(n15504), .ZN(n16607) );
  AND3_X2 U1105 ( .A1(n14130), .A2(n14129), .A3(n14128), .ZN(n14752) );
  XNOR2_X2 U8465 ( .A(Key[111]), .B(Plaintext[111]), .ZN(n7626) );
  AND3_X2 U8079 ( .A1(n2049), .A2(n20984), .A3(n21812), .ZN(n22713) );
  NAND2_X2 U4045 ( .A1(n910), .A2(n5547), .ZN(n23467) );
  BUF_X1 U3426 ( .A(n7017), .Z(n8245) );
  OR2_X2 U1101 ( .A1(n8684), .A2(n8683), .ZN(n9949) );
  NAND2_X2 U1697 ( .A1(n6444), .A2(n6443), .ZN(n19025) );
  MUX2_X2 U2035 ( .A(n7820), .B(n7819), .S(n8243), .Z(n9016) );
  OR2_X2 U938 ( .A1(n17585), .A2(n1376), .ZN(n19245) );
  AND2_X2 U849 ( .A1(n17705), .A2(n17704), .ZN(n19603) );
  NAND3_X2 U10806 ( .A1(n3676), .A2(n3675), .A3(n7227), .ZN(n9971) );
  MUX2_X2 U9935 ( .A(n7081), .B(n7080), .S(n8812), .Z(n10037) );
  NAND2_X2 U1437 ( .A1(n5034), .A2(n5033), .ZN(n21932) );
  NAND2_X2 U348 ( .A1(n2678), .A2(n10857), .ZN(n12241) );
  MUX2_X2 U10408 ( .A(n26839), .B(n26838), .S(n26837), .Z(n27843) );
  OR2_X2 U24797 ( .A1(n22983), .A2(n22982), .ZN(n24433) );
  BUF_X2 U1533 ( .A(n8847), .Z(n12205) );
  AND3_X2 U2465 ( .A1(n20796), .A2(n20795), .A3(n20794), .ZN(n22790) );
  MUX2_X2 U12 ( .A(n24371), .B(n24370), .S(n24369), .Z(n25430) );
  NAND3_X2 U4745 ( .A1(n23439), .A2(n1228), .A3(n23438), .ZN(n24256) );
  BUF_X1 U1568 ( .A(n20224), .Z(n296) );
  NAND2_X2 U684 ( .A1(n11296), .A2(n3556), .ZN(n12841) );
  NAND2_X2 U11437 ( .A1(n26934), .A2(n6950), .ZN(n27527) );
  XNOR2_X2 U2043 ( .A(n7138), .B(Key[48]), .ZN(n8013) );
  NAND2_X2 U10033 ( .A1(n24333), .A2(n3696), .ZN(n26059) );
  XNOR2_X2 U3215 ( .A(n9804), .B(n9803), .ZN(n10992) );
  MUX2_X2 U22792 ( .A(n19862), .B(n19861), .S(n385), .Z(n20744) );
  OAI211_X2 U19927 ( .C1(n15495), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        n16309) );
  OAI21_X2 U9185 ( .B1(n8743), .B2(n8742), .A(n2859), .ZN(n10265) );
  NOR2_X1 U8068 ( .A1(n7569), .A2(n8326), .ZN(n8581) );
  AOI21_X2 U1548 ( .B1(n9145), .B2(n9144), .A(n9143), .ZN(n10159) );
  BUF_X1 U3202 ( .A(n10482), .Z(n11258) );
  AND2_X1 U5280 ( .A1(n1663), .A2(n11974), .ZN(n1664) );
  BUF_X1 U1754 ( .A(n18522), .Z(n374) );
  OAI21_X1 U2570 ( .B1(n20694), .B2(n6730), .A(n20693), .ZN(n21810) );
  BUF_X1 U5902 ( .A(n23702), .Z(n23387) );
  NAND3_X1 U4140 ( .A1(n24342), .A2(n2460), .A3(n24343), .ZN(n25697) );
  XNOR2_X1 U47 ( .A(n6447), .B(n16080), .ZN(n16812) );
  BUF_X1 U77 ( .A(n8151), .Z(n28149) );
  NAND3_X2 U118 ( .A1(n28306), .A2(n15038), .A3(n28305), .ZN(n15989) );
  NAND3_X2 U126 ( .A1(n4550), .A2(n4551), .A3(n7826), .ZN(n9012) );
  NAND3_X2 U135 ( .A1(n28707), .A2(n3499), .A3(n5387), .ZN(n24697) );
  OAI21_X2 U194 ( .B1(n19857), .B2(n20556), .A(n19856), .ZN(n21481) );
  BUF_X1 U216 ( .A(n1308), .Z(n28407) );
  OR2_X2 U235 ( .A1(n14269), .A2(n14270), .ZN(n15260) );
  XNOR2_X1 U293 ( .A(n26064), .B(n26063), .ZN(n27111) );
  OAI21_X2 U307 ( .B1(n4351), .B2(n10871), .A(n4350), .ZN(n12236) );
  AND3_X2 U323 ( .A1(n3023), .A2(n4045), .A3(n4171), .ZN(n11430) );
  XNOR2_X1 U335 ( .A(n12458), .B(n12457), .ZN(n14416) );
  NOR2_X1 U353 ( .A1(n14036), .A2(n13719), .ZN(n28121) );
  XOR2_X1 U378 ( .A(n21492), .B(n21491), .Z(n28122) );
  XNOR2_X2 U383 ( .A(n24522), .B(n4643), .ZN(n28578) );
  INV_X1 U396 ( .A(n17696), .ZN(n16898) );
  XNOR2_X1 U429 ( .A(n19432), .B(n19431), .ZN(n21355) );
  NAND2_X2 U444 ( .A1(n4609), .A2(n4608), .ZN(n14733) );
  XNOR2_X2 U471 ( .A(n4764), .B(n25928), .ZN(n25412) );
  NOR2_X2 U500 ( .A1(n20596), .A2(n20595), .ZN(n21801) );
  OAI21_X2 U507 ( .B1(n7578), .B2(n7577), .A(n7576), .ZN(n8717) );
  BUF_X2 U525 ( .A(n21356), .Z(n28133) );
  XNOR2_X1 U527 ( .A(n19437), .B(n19436), .ZN(n21356) );
  XNOR2_X2 U551 ( .A(n25098), .B(n25097), .ZN(n26799) );
  XNOR2_X2 U562 ( .A(n9093), .B(n9092), .ZN(n11192) );
  XNOR2_X2 U566 ( .A(n15628), .B(n15627), .ZN(n17359) );
  XNOR2_X1 U587 ( .A(n22049), .B(n22048), .ZN(n23250) );
  NOR2_X2 U592 ( .A1(n13313), .A2(n13312), .ZN(n16346) );
  XNOR2_X2 U601 ( .A(n6074), .B(n21757), .ZN(n23036) );
  OAI21_X2 U608 ( .B1(n17778), .B2(n17980), .A(n6264), .ZN(n19685) );
  AOI21_X2 U623 ( .B1(n26249), .B2(n26248), .A(n26247), .ZN(n28065) );
  OAI211_X2 U634 ( .C1(n21187), .C2(n22288), .A(n1694), .B(n1692), .ZN(n22690)
         );
  OR2_X2 U636 ( .A1(n3486), .A2(n21592), .ZN(n21998) );
  OAI21_X2 U670 ( .B1(n18627), .B2(n20381), .A(n18626), .ZN(n21218) );
  NOR2_X2 U695 ( .A1(n20898), .A2(n20897), .ZN(n1925) );
  XNOR2_X2 U697 ( .A(n13047), .B(n13046), .ZN(n14354) );
  XNOR2_X2 U718 ( .A(n15820), .B(n15821), .ZN(n17555) );
  OAI21_X2 U721 ( .B1(n7923), .B2(n8234), .A(n7922), .ZN(n9108) );
  OR2_X2 U735 ( .A1(n20138), .A2(n20139), .ZN(n21425) );
  NOR2_X1 U746 ( .A1(n17010), .A2(n17011), .ZN(n18601) );
  INV_X1 U753 ( .A(n13842), .ZN(n14345) );
  NOR2_X1 U756 ( .A1(n18543), .A2(n28339), .ZN(n19556) );
  AND2_X2 U757 ( .A1(n11134), .A2(n11775), .ZN(n11551) );
  BUF_X2 U766 ( .A(n20354), .Z(n383) );
  XNOR2_X2 U778 ( .A(n13515), .B(n13514), .ZN(n13587) );
  NOR2_X2 U785 ( .A1(n3243), .A2(n19975), .ZN(n21956) );
  CLKBUF_X1 U794 ( .A(n11275), .Z(n28147) );
  XNOR2_X2 U831 ( .A(n4747), .B(n4745), .ZN(n20494) );
  AND3_X2 U857 ( .A1(n23379), .A2(n23381), .A3(n23380), .ZN(n25933) );
  XNOR2_X2 U882 ( .A(n25286), .B(n25285), .ZN(n26723) );
  XNOR2_X2 U896 ( .A(n7105), .B(Key[186]), .ZN(n7312) );
  INV_X1 U905 ( .A(n10544), .ZN(n10742) );
  AND3_X2 U911 ( .A1(n1105), .A2(n19919), .A3(n4658), .ZN(n20658) );
  XNOR2_X2 U964 ( .A(n6980), .B(Key[96]), .ZN(n7828) );
  XNOR2_X2 U968 ( .A(n23861), .B(n23860), .ZN(n25418) );
  XNOR2_X2 U1058 ( .A(n7003), .B(Key[72]), .ZN(n7250) );
  NAND2_X2 U1067 ( .A1(n5619), .A2(n5618), .ZN(n24408) );
  OAI211_X2 U1077 ( .C1(n8823), .C2(n7529), .A(n8475), .B(n7528), .ZN(n10395)
         );
  BUF_X2 U1091 ( .A(n21565), .Z(n28155) );
  OAI211_X1 U1096 ( .C1(n19792), .C2(n20488), .A(n5208), .B(n2383), .ZN(n21565) );
  CLKBUF_X1 U1143 ( .A(n7141), .Z(n28161) );
  AOI22_X2 U1155 ( .A1(n2220), .A2(n11750), .B1(n28698), .B2(n11501), .ZN(
        n12965) );
  NOR3_X1 U1183 ( .A1(n20428), .A2(n20427), .A3(n20426), .ZN(n22765) );
  XNOR2_X2 U1203 ( .A(n15540), .B(n15539), .ZN(n17025) );
  AND3_X2 U1207 ( .A1(n17468), .A2(n3981), .A3(n3980), .ZN(n18500) );
  AND2_X2 U1228 ( .A1(n1539), .A2(n1542), .ZN(n22522) );
  INV_X1 U1281 ( .A(n10830), .ZN(n11338) );
  NOR2_X2 U1305 ( .A1(n24026), .A2(n24025), .ZN(n4764) );
  AND2_X2 U1324 ( .A1(n4177), .A2(n3204), .ZN(n24405) );
  OAI211_X2 U1325 ( .C1(n12587), .C2(n13711), .A(n12586), .B(n12585), .ZN(
        n15094) );
  OAI211_X2 U1326 ( .C1(n3880), .C2(n1581), .A(n3878), .B(n3879), .ZN(n18421)
         );
  AND2_X2 U1342 ( .A1(n2942), .A2(n2941), .ZN(n9140) );
  AOI21_X2 U1348 ( .B1(n21234), .B2(n21389), .A(n21233), .ZN(n22195) );
  XNOR2_X2 U1353 ( .A(n19471), .B(n19470), .ZN(n20443) );
  OAI21_X2 U1364 ( .B1(n5863), .B2(n24146), .A(n24145), .ZN(n25391) );
  XNOR2_X2 U1391 ( .A(n4430), .B(n5184), .ZN(n4086) );
  OAI22_X2 U1393 ( .A1(n4661), .A2(n4660), .B1(n14580), .B2(n15095), .ZN(
        n16494) );
  XNOR2_X2 U1394 ( .A(n9288), .B(n9287), .ZN(n10942) );
  XNOR2_X2 U1415 ( .A(n12530), .B(n12531), .ZN(n13872) );
  AOI21_X2 U1422 ( .B1(n792), .B2(n17226), .A(n4763), .ZN(n18431) );
  BUF_X2 U1488 ( .A(n24074), .Z(n24072) );
  AND2_X1 U1529 ( .A1(n17423), .A2(n17421), .ZN(n28739) );
  BUF_X1 U1530 ( .A(n17452), .Z(n28193) );
  BUF_X1 U1532 ( .A(n15980), .Z(n17275) );
  INV_X1 U1545 ( .A(n13730), .ZN(n28171) );
  INV_X1 U1559 ( .A(n10957), .ZN(n28173) );
  INV_X1 U1572 ( .A(n11045), .ZN(n28174) );
  INV_X1 U1573 ( .A(n11158), .ZN(n28175) );
  INV_X1 U1574 ( .A(n10703), .ZN(n28176) );
  AND2_X1 U1579 ( .A1(n9196), .A2(n9197), .ZN(n231) );
  AND3_X1 U1608 ( .A1(n2432), .A2(n28341), .A3(n2434), .ZN(n27220) );
  AOI22_X1 U1609 ( .A1(n29021), .A2(n27958), .B1(n29092), .B2(n27996), .ZN(
        n27998) );
  NAND3_X1 U1611 ( .A1(n27009), .A2(n27008), .A3(n27007), .ZN(n27926) );
  OAI21_X1 U1613 ( .B1(n24857), .B2(n4679), .A(n24856), .ZN(n28466) );
  AND3_X1 U1625 ( .A1(n28216), .A2(n28238), .A3(n28237), .ZN(n27800) );
  INV_X1 U1632 ( .A(n27594), .ZN(n28179) );
  OR3_X1 U1634 ( .A1(n26129), .A2(n28392), .A3(n27129), .ZN(n27135) );
  XNOR2_X1 U1644 ( .A(n25478), .B(n28230), .ZN(n26623) );
  INV_X1 U1645 ( .A(n29474), .ZN(n28180) );
  AND2_X1 U1657 ( .A1(n24102), .A2(n24101), .ZN(n28256) );
  NOR2_X1 U1658 ( .A1(n22177), .A2(n24468), .ZN(n22178) );
  OR2_X1 U1659 ( .A1(n24583), .A2(n24584), .ZN(n28315) );
  BUF_X1 U1663 ( .A(n24790), .Z(n28512) );
  OR2_X1 U1673 ( .A1(n29567), .A2(n24391), .ZN(n2648) );
  CLKBUF_X1 U1676 ( .A(n24717), .Z(n28416) );
  AND4_X1 U1679 ( .A1(n6154), .A2(n4234), .A3(n4233), .A4(n6153), .ZN(n28509)
         );
  AND2_X1 U1680 ( .A1(n23783), .A2(n23787), .ZN(n21769) );
  OR2_X1 U1684 ( .A1(n23772), .A2(n23771), .ZN(n23021) );
  INV_X1 U1692 ( .A(n22566), .ZN(n28181) );
  XNOR2_X1 U1698 ( .A(n22850), .B(n22849), .ZN(n28609) );
  OR2_X1 U1699 ( .A1(n23769), .A2(n23763), .ZN(n28354) );
  INV_X1 U1702 ( .A(n23725), .ZN(n28183) );
  AOI22_X1 U1717 ( .A1(n28750), .A2(n28749), .B1(n22012), .B2(n20537), .ZN(
        n20798) );
  INV_X1 U1718 ( .A(n21068), .ZN(n28301) );
  INV_X1 U1719 ( .A(n20853), .ZN(n20852) );
  OR2_X1 U1723 ( .A1(n21581), .A2(n21481), .ZN(n28723) );
  BUF_X1 U1729 ( .A(n21343), .Z(n28440) );
  INV_X1 U1730 ( .A(n20663), .ZN(n28184) );
  INV_X1 U1734 ( .A(n21541), .ZN(n28185) );
  OAI21_X1 U1736 ( .B1(n2715), .B2(n18831), .A(n19773), .ZN(n28326) );
  INV_X1 U1738 ( .A(n20162), .ZN(n28187) );
  INV_X1 U1742 ( .A(n20099), .ZN(n28188) );
  XNOR2_X1 U1746 ( .A(n6157), .B(n19135), .ZN(n20506) );
  INV_X1 U1755 ( .A(n19413), .ZN(n18628) );
  NOR2_X1 U1764 ( .A1(n17724), .A2(n373), .ZN(n19659) );
  OR2_X1 U1765 ( .A1(n18291), .A2(n18292), .ZN(n3768) );
  INV_X1 U1767 ( .A(n18493), .ZN(n18487) );
  OR2_X1 U1777 ( .A1(n18387), .A2(n18393), .ZN(n686) );
  OR2_X1 U1787 ( .A1(n4732), .A2(n526), .ZN(n17330) );
  OR2_X1 U1794 ( .A1(n18193), .A2(n16718), .ZN(n1025) );
  NAND2_X1 U1796 ( .A1(n1592), .A2(n1591), .ZN(n18493) );
  OR2_X1 U1801 ( .A1(n526), .A2(n18144), .ZN(n193) );
  INV_X1 U1803 ( .A(n17762), .ZN(n28191) );
  OR2_X1 U1848 ( .A1(n28323), .A2(n4270), .ZN(n2858) );
  AND2_X1 U1880 ( .A1(n17355), .A2(n17357), .ZN(n16713) );
  XNOR2_X1 U1889 ( .A(n15699), .B(n15700), .ZN(n17368) );
  INV_X1 U1893 ( .A(n17426), .ZN(n28194) );
  INV_X1 U1947 ( .A(n14942), .ZN(n28195) );
  AND2_X1 U1991 ( .A1(n12414), .A2(n12415), .ZN(n14906) );
  INV_X1 U2008 ( .A(n15060), .ZN(n28197) );
  INV_X1 U2021 ( .A(n14695), .ZN(n28198) );
  OR2_X1 U2031 ( .A1(n28569), .A2(n13587), .ZN(n28257) );
  INV_X1 U2104 ( .A(n13703), .ZN(n28199) );
  INV_X1 U2144 ( .A(n14438), .ZN(n28200) );
  INV_X1 U2148 ( .A(n12696), .ZN(n12861) );
  NAND3_X1 U2174 ( .A1(n28682), .A2(n3987), .A3(n11391), .ZN(n4474) );
  OR2_X1 U2201 ( .A1(n12081), .A2(n3558), .ZN(n28703) );
  INV_X1 U2249 ( .A(n12232), .ZN(n28201) );
  INV_X1 U2255 ( .A(n12211), .ZN(n28203) );
  AND2_X1 U2258 ( .A1(n4352), .A2(n10666), .ZN(n28363) );
  INV_X1 U2259 ( .A(n10668), .ZN(n28204) );
  INV_X1 U2263 ( .A(n11113), .ZN(n28205) );
  INV_X1 U2281 ( .A(n11145), .ZN(n28206) );
  XNOR2_X1 U2286 ( .A(n6891), .B(n9309), .ZN(n28608) );
  INV_X1 U2307 ( .A(n10467), .ZN(n28208) );
  AND3_X1 U2345 ( .A1(n1045), .A2(n28352), .A3(n5130), .ZN(n9323) );
  AOI21_X1 U2357 ( .B1(n9419), .B2(n604), .A(n9420), .ZN(n2290) );
  INV_X1 U2414 ( .A(n9028), .ZN(n28210) );
  INV_X1 U2422 ( .A(n8109), .ZN(n28211) );
  INV_X1 U2442 ( .A(n9075), .ZN(n28212) );
  OR2_X1 U2446 ( .A1(n6988), .A2(n7822), .ZN(n7426) );
  OR2_X1 U2452 ( .A1(n7935), .A2(n7933), .ZN(n7616) );
  INV_X1 U2466 ( .A(n3154), .ZN(n28213) );
  CLKBUF_X1 U2467 ( .A(Key[172]), .Z(n28294) );
  INV_X1 U2503 ( .A(n7822), .ZN(n3821) );
  INV_X1 U2526 ( .A(n441), .ZN(n7870) );
  OAI21_X1 U2544 ( .B1(n627), .B2(n8217), .A(n7925), .ZN(n6961) );
  BUF_X1 U2557 ( .A(n7093), .Z(n7309) );
  OR2_X1 U2565 ( .A1(n9009), .A2(n9007), .ZN(n9189) );
  INV_X1 U2585 ( .A(n8440), .ZN(n28743) );
  OR2_X1 U2590 ( .A1(n7952), .A2(n8258), .ZN(n117) );
  AND3_X1 U2603 ( .A1(n1418), .A2(n1417), .A3(n7574), .ZN(n28281) );
  OR2_X1 U2605 ( .A1(n8351), .A2(n8353), .ZN(n238) );
  BUF_X1 U2620 ( .A(n7665), .Z(n8265) );
  NAND2_X1 U2656 ( .A1(n4673), .A2(n4674), .ZN(n8192) );
  OR2_X1 U2657 ( .A1(n8976), .A2(n8819), .ZN(n142) );
  OR2_X1 U2660 ( .A1(n10406), .A2(n3787), .ZN(n2891) );
  OR2_X1 U2674 ( .A1(n8575), .A2(n9421), .ZN(n28352) );
  OR2_X1 U2684 ( .A1(n9139), .A2(n8185), .ZN(n8187) );
  AOI21_X1 U2710 ( .B1(n8738), .B2(n8731), .A(n8730), .ZN(n8374) );
  AND2_X1 U2717 ( .A1(n8702), .A2(n8700), .ZN(n105) );
  INV_X1 U2747 ( .A(n8077), .ZN(n8431) );
  NOR2_X1 U2756 ( .A1(n8491), .A2(n8666), .ZN(n8495) );
  OR2_X1 U2792 ( .A1(n8598), .A2(n9062), .ZN(n8402) );
  XNOR2_X1 U2799 ( .A(n9635), .B(n9634), .ZN(n11047) );
  OR2_X1 U2822 ( .A1(n10942), .A2(n10703), .ZN(n28310) );
  MUX2_X1 U2831 ( .A(n11034), .B(n10671), .S(n28147), .Z(n10672) );
  NOR2_X1 U2836 ( .A1(n11106), .A2(n10871), .ZN(n10280) );
  INV_X1 U2855 ( .A(n10482), .ZN(n4296) );
  NOR2_X1 U2886 ( .A1(n4389), .A2(n10741), .ZN(n4390) );
  XNOR2_X1 U2900 ( .A(n2662), .B(n1988), .ZN(n10930) );
  AND2_X1 U2927 ( .A1(n6703), .A2(n2063), .ZN(n28336) );
  AND2_X1 U2932 ( .A1(n11888), .A2(n12328), .ZN(n28260) );
  OR2_X1 U2934 ( .A1(n349), .A2(n11933), .ZN(n11594) );
  INV_X1 U2935 ( .A(n11377), .ZN(n12167) );
  OAI211_X1 U2959 ( .C1(n11799), .C2(n12289), .A(n11798), .B(n11797), .ZN(
        n12734) );
  INV_X1 U2975 ( .A(n12589), .ZN(n13539) );
  AND2_X1 U2981 ( .A1(n14295), .A2(n14293), .ZN(n28322) );
  AND2_X1 U2983 ( .A1(n14304), .A2(n5341), .ZN(n28273) );
  XNOR2_X1 U2986 ( .A(n11866), .B(n11865), .ZN(n14252) );
  OAI21_X1 U3037 ( .B1(n12122), .B2(n12121), .A(n14487), .ZN(n141) );
  NAND2_X1 U3044 ( .A1(n1389), .A2(n57), .ZN(n14971) );
  OR2_X1 U3085 ( .A1(n14583), .A2(n14971), .ZN(n14886) );
  OAI211_X1 U3098 ( .C1(n13651), .C2(n14302), .A(n13650), .B(n13649), .ZN(
        n15117) );
  OR2_X1 U3116 ( .A1(n15351), .A2(n15343), .ZN(n150) );
  CLKBUF_X1 U3147 ( .A(n14826), .Z(n15030) );
  AND2_X1 U3163 ( .A1(n15009), .A2(n15370), .ZN(n15376) );
  OAI21_X1 U3170 ( .B1(n1662), .B2(n15376), .A(n15371), .ZN(n5) );
  XNOR2_X1 U3191 ( .A(n6080), .B(n16494), .ZN(n15903) );
  AND2_X1 U3214 ( .A1(n5714), .A2(n17304), .ZN(n28233) );
  NOR2_X1 U3228 ( .A1(n28233), .A2(n16968), .ZN(n28232) );
  OR2_X1 U3265 ( .A1(n17139), .A2(n16887), .ZN(n17135) );
  NOR2_X1 U3279 ( .A1(n16706), .A2(n16884), .ZN(n16430) );
  AND2_X1 U3303 ( .A1(n18181), .A2(n18180), .ZN(n17738) );
  OR2_X1 U3342 ( .A1(n517), .A2(n17762), .ZN(n66) );
  OR2_X1 U3412 ( .A1(n1384), .A2(n18467), .ZN(n17917) );
  AND2_X1 U3420 ( .A1(n18458), .A2(n18106), .ZN(n28241) );
  OR2_X1 U3496 ( .A1(n2853), .A2(n18430), .ZN(n18147) );
  BUF_X1 U3502 ( .A(n18708), .Z(n28558) );
  OR2_X1 U3507 ( .A1(n17814), .A2(n420), .ZN(n17247) );
  INV_X1 U3518 ( .A(n18423), .ZN(n512) );
  OR2_X1 U3519 ( .A1(n5203), .A2(n18171), .ZN(n17785) );
  XNOR2_X1 U3532 ( .A(n18737), .B(n19475), .ZN(n19040) );
  OR2_X1 U3541 ( .A1(n18019), .A2(n28370), .ZN(n3070) );
  XNOR2_X1 U3570 ( .A(n18926), .B(n18925), .ZN(n28479) );
  AND2_X1 U3578 ( .A1(n21088), .A2(n628), .ZN(n28275) );
  NOR2_X1 U3584 ( .A1(n20382), .A2(n28508), .ZN(n20385) );
  OR2_X1 U3593 ( .A1(n21227), .A2(n21392), .ZN(n3418) );
  AND2_X1 U3615 ( .A1(n21171), .A2(n21047), .ZN(n28287) );
  OR2_X1 U3616 ( .A1(n21144), .A2(n21118), .ZN(n20853) );
  XNOR2_X1 U3641 ( .A(n1859), .B(n5803), .ZN(n22058) );
  OR2_X1 U3642 ( .A1(n4104), .A2(n43), .ZN(n4203) );
  AND3_X1 U3655 ( .A1(n20532), .A2(n20933), .A3(n20533), .ZN(n20426) );
  INV_X1 U3682 ( .A(n4872), .ZN(n23150) );
  OR2_X1 U3701 ( .A1(n23712), .A2(n22174), .ZN(n22163) );
  NOR2_X1 U3716 ( .A1(n23629), .A2(n23630), .ZN(n23555) );
  XNOR2_X1 U3723 ( .A(n22115), .B(n22114), .ZN(n23726) );
  OR2_X1 U3729 ( .A1(n23647), .A2(n2779), .ZN(n640) );
  XNOR2_X1 U3739 ( .A(n22083), .B(n22082), .ZN(n23386) );
  XNOR2_X1 U3745 ( .A(n21104), .B(n21105), .ZN(n23360) );
  AND2_X1 U3760 ( .A1(n23147), .A2(n23461), .ZN(n4872) );
  OR2_X1 U3772 ( .A1(n23465), .A2(n22926), .ZN(n28317) );
  OR2_X1 U3850 ( .A1(n23388), .A2(n23704), .ZN(n28695) );
  OR2_X1 U3856 ( .A1(n22867), .A2(n22866), .ZN(n28519) );
  OR2_X1 U3866 ( .A1(n23373), .A2(n24316), .ZN(n28681) );
  NOR2_X1 U3871 ( .A1(n24816), .A2(n24461), .ZN(n28678) );
  AND2_X1 U3893 ( .A1(n23590), .A2(n24447), .ZN(n28330) );
  XNOR2_X1 U3906 ( .A(n25693), .B(n25692), .ZN(n28545) );
  BUF_X1 U3912 ( .A(n26941), .Z(n28541) );
  AOI21_X1 U3943 ( .B1(n28289), .B2(n28288), .A(n26352), .ZN(n26354) );
  XNOR2_X1 U3994 ( .A(n25854), .B(n25853), .ZN(n26837) );
  NOR2_X1 U4001 ( .A1(n25814), .A2(n27087), .ZN(n28249) );
  NOR2_X1 U4032 ( .A1(n27038), .A2(n27379), .ZN(n26610) );
  AND3_X1 U4118 ( .A1(n3390), .A2(n6634), .A3(n6633), .ZN(n27548) );
  INV_X1 U4131 ( .A(n26696), .ZN(n28248) );
  NAND3_X1 U4135 ( .A1(n6755), .A2(n5391), .A3(n5390), .ZN(n27244) );
  CLKBUF_X1 U4144 ( .A(Key[151]), .Z(n27105) );
  CLKBUF_X1 U4146 ( .A(Key[154]), .Z(n2510) );
  AND2_X1 U4151 ( .A1(n29537), .A2(n26314), .ZN(n28214) );
  NAND3_X1 U4160 ( .A1(n29644), .A2(n20191), .A3(n20541), .ZN(n28215) );
  OR3_X1 U4162 ( .A1(n5299), .A2(n27060), .A3(n26849), .ZN(n28216) );
  OR2_X1 U4190 ( .A1(n28228), .A2(n29076), .ZN(n28217) );
  INV_X1 U4198 ( .A(n7424), .ZN(n28721) );
  AND2_X1 U4201 ( .A1(n7837), .A2(n7700), .ZN(n28218) );
  AND2_X1 U4202 ( .A1(n7492), .A2(n8850), .ZN(n28219) );
  INV_X1 U4229 ( .A(n10929), .ZN(n10927) );
  INV_X1 U4247 ( .A(n12042), .ZN(n28726) );
  AND2_X1 U4265 ( .A1(n14455), .A2(n14200), .ZN(n28220) );
  INV_X1 U4266 ( .A(n14696), .ZN(n15288) );
  OR2_X1 U4268 ( .A1(n15081), .A2(n15082), .ZN(n28221) );
  NOR2_X1 U4279 ( .A1(n14763), .A2(n15260), .ZN(n28222) );
  INV_X1 U4281 ( .A(n17294), .ZN(n28729) );
  INV_X1 U4282 ( .A(n15691), .ZN(n28666) );
  INV_X1 U4308 ( .A(n18020), .ZN(n28370) );
  NAND4_X2 U4323 ( .A1(n4189), .A2(n4190), .A3(n6410), .A4(n6409), .ZN(n22290)
         );
  OR2_X1 U4335 ( .A1(n20657), .A2(n20656), .ZN(n28223) );
  NAND3_X1 U4351 ( .A1(n23326), .A2(n23034), .A3(n23760), .ZN(n28224) );
  XOR2_X1 U4360 ( .A(n22191), .B(n22190), .Z(n28225) );
  XOR2_X1 U4387 ( .A(n24962), .B(n24961), .Z(n28226) );
  AND2_X1 U4393 ( .A1(n24668), .A2(n24665), .ZN(n28227) );
  XOR2_X1 U4394 ( .A(n25719), .B(n25718), .Z(n28228) );
  INV_X1 U4421 ( .A(n23862), .ZN(n28710) );
  AND2_X1 U4423 ( .A1(n29060), .A2(n29474), .ZN(n28229) );
  XOR2_X1 U4428 ( .A(n25476), .B(n25475), .Z(n28230) );
  NAND2_X1 U4511 ( .A1(n4543), .A2(n6053), .ZN(n4542) );
  NAND2_X1 U4550 ( .A1(n28232), .A2(n28231), .ZN(n6224) );
  NAND2_X1 U4551 ( .A1(n28768), .A2(n1738), .ZN(n28231) );
  NAND2_X1 U4572 ( .A1(n20377), .A2(n20371), .ZN(n28235) );
  NAND2_X1 U4583 ( .A1(n20376), .A2(n351), .ZN(n28236) );
  NAND2_X1 U4593 ( .A1(n26328), .A2(n28600), .ZN(n28237) );
  NAND2_X1 U4597 ( .A1(n26329), .A2(n27056), .ZN(n28238) );
  NAND2_X1 U4603 ( .A1(n6931), .A2(n19951), .ZN(n28244) );
  NAND2_X1 U4616 ( .A1(n28240), .A2(n20192), .ZN(n3016) );
  NOR2_X1 U4642 ( .A1(n503), .A2(n20416), .ZN(n28240) );
  NAND3_X1 U4651 ( .A1(n4033), .A2(n28393), .A3(n4236), .ZN(n4032) );
  NAND2_X1 U4664 ( .A1(n17729), .A2(n18109), .ZN(n3849) );
  NAND2_X1 U4710 ( .A1(n28242), .A2(n5822), .ZN(n5820) );
  NAND2_X1 U4733 ( .A1(n5804), .A2(n13935), .ZN(n28242) );
  NAND2_X1 U4741 ( .A1(n28243), .A2(n5943), .ZN(n21581) );
  NAND3_X1 U4742 ( .A1(n19839), .A2(n5100), .A3(n5099), .ZN(n28243) );
  NOR2_X1 U4764 ( .A1(n19953), .A2(n28244), .ZN(n21729) );
  NAND3_X1 U4767 ( .A1(n28641), .A2(n27862), .A3(n27324), .ZN(n27325) );
  NAND2_X1 U4778 ( .A1(n24241), .A2(n24559), .ZN(n5332) );
  AOI21_X1 U4786 ( .B1(n15267), .B2(n15266), .A(n15506), .ZN(n28245) );
  NAND2_X1 U4925 ( .A1(n1483), .A2(n24780), .ZN(n24781) );
  NAND2_X1 U4945 ( .A1(n28246), .A2(n8204), .ZN(n8206) );
  NOR2_X2 U4977 ( .A1(n5289), .A2(n28247), .ZN(n4384) );
  NOR2_X1 U4996 ( .A1(n24058), .A2(n459), .ZN(n28247) );
  OR2_X1 U4998 ( .A1(n20381), .A2(n20573), .ZN(n19834) );
  NAND3_X1 U4999 ( .A1(n447), .A2(n3681), .A3(n28248), .ZN(n26643) );
  NOR2_X2 U5011 ( .A1(n25834), .A2(n28249), .ZN(n27872) );
  NOR2_X2 U5049 ( .A1(n28251), .A2(n28250), .ZN(n18802) );
  OAI22_X1 U5063 ( .A1(n18013), .A2(n18480), .B1(n18012), .B2(n18011), .ZN(
        n28250) );
  NAND2_X1 U5067 ( .A1(n6574), .A2(n6575), .ZN(n28251) );
  NAND2_X1 U5113 ( .A1(n28894), .A2(n20430), .ZN(n28252) );
  NAND2_X1 U5118 ( .A1(n24590), .A2(n831), .ZN(n4692) );
  NAND2_X2 U5131 ( .A1(n28317), .A2(n5269), .ZN(n831) );
  OAI21_X2 U5149 ( .B1(n12310), .B2(n28253), .A(n12309), .ZN(n13419) );
  NOR2_X1 U5153 ( .A1(n12299), .A2(n12303), .ZN(n28253) );
  NAND3_X1 U5154 ( .A1(n26930), .A2(n26927), .A3(n26926), .ZN(n1277) );
  NAND2_X1 U5180 ( .A1(n1561), .A2(n18172), .ZN(n28254) );
  NAND2_X1 U5183 ( .A1(n24099), .A2(n53), .ZN(n28255) );
  OAI21_X1 U5195 ( .B1(n14976), .B2(n14974), .A(n14973), .ZN(n14975) );
  NAND2_X1 U5196 ( .A1(n14971), .A2(n13789), .ZN(n14974) );
  NAND2_X1 U5244 ( .A1(n21440), .A2(n6275), .ZN(n28258) );
  NAND2_X1 U5246 ( .A1(n20244), .A2(n21661), .ZN(n28259) );
  AOI21_X1 U5254 ( .B1(n12333), .B2(n12332), .A(n28260), .ZN(n11748) );
  OAI21_X1 U5299 ( .B1(n6097), .B2(n24493), .A(n28261), .ZN(n690) );
  NAND3_X1 U5300 ( .A1(n24470), .A2(n23942), .A3(n29033), .ZN(n28261) );
  NAND2_X1 U5301 ( .A1(n26573), .A2(n29576), .ZN(n28284) );
  NAND2_X1 U5318 ( .A1(n28263), .A2(n28262), .ZN(n24393) );
  NAND2_X1 U5320 ( .A1(n24392), .A2(n29471), .ZN(n28263) );
  NAND3_X2 U5376 ( .A1(n11620), .A2(n28265), .A3(n28264), .ZN(n13055) );
  NAND2_X1 U5379 ( .A1(n11618), .A2(n5637), .ZN(n28264) );
  INV_X1 U5388 ( .A(n11989), .ZN(n28265) );
  NAND2_X1 U5425 ( .A1(n28268), .A2(n28266), .ZN(n8815) );
  NAND2_X1 U5441 ( .A1(n8814), .A2(n28267), .ZN(n28266) );
  INV_X1 U5465 ( .A(n8812), .ZN(n28267) );
  NAND2_X1 U5483 ( .A1(n8681), .A2(n8810), .ZN(n8814) );
  NAND2_X1 U5498 ( .A1(n8813), .A2(n8812), .ZN(n28268) );
  AOI21_X1 U5503 ( .B1(n10569), .B2(n4101), .A(n28270), .ZN(n28269) );
  INV_X1 U5511 ( .A(n10795), .ZN(n28270) );
  NAND2_X1 U5523 ( .A1(n17833), .A2(n17832), .ZN(n17838) );
  XNOR2_X1 U5524 ( .A(n28271), .B(n26214), .ZN(Ciphertext[14]) );
  NAND2_X1 U5540 ( .A1(n4032), .A2(n4034), .ZN(n28271) );
  NAND3_X1 U5555 ( .A1(n27721), .A2(n27719), .A3(n27720), .ZN(n27722) );
  OAI21_X2 U5584 ( .B1(n11209), .B2(n10656), .A(n10655), .ZN(n375) );
  NAND2_X1 U5597 ( .A1(n2196), .A2(n8359), .ZN(n9948) );
  OAI21_X2 U5598 ( .B1(n20116), .B2(n20117), .A(n20115), .ZN(n21424) );
  NAND2_X1 U5626 ( .A1(n1422), .A2(n1426), .ZN(n28274) );
  NAND2_X1 U5632 ( .A1(n1420), .A2(n23946), .ZN(n1425) );
  NAND2_X1 U5677 ( .A1(n11220), .A2(n11223), .ZN(n11106) );
  NAND2_X1 U5681 ( .A1(n3237), .A2(n28275), .ZN(n1267) );
  NAND3_X1 U5711 ( .A1(n28276), .A2(n1606), .A3(n7354), .ZN(n9139) );
  NAND2_X1 U5740 ( .A1(n1608), .A2(n7353), .ZN(n28276) );
  NAND2_X1 U5743 ( .A1(n13829), .A2(n14360), .ZN(n14075) );
  XNOR2_X1 U5764 ( .A(n28277), .B(n27643), .ZN(Ciphertext[98]) );
  AOI22_X1 U5797 ( .A1(n27642), .A2(n27641), .B1(n27647), .B2(n27640), .ZN(
        n28277) );
  OAI21_X1 U5810 ( .B1(n20078), .B2(n20079), .A(n20077), .ZN(n20086) );
  NOR2_X1 U5828 ( .A1(n7454), .A2(n28278), .ZN(n7461) );
  INV_X1 U5831 ( .A(n7984), .ZN(n28278) );
  NAND2_X1 U5839 ( .A1(n7643), .A2(n7456), .ZN(n7984) );
  INV_X1 U5867 ( .A(n9575), .ZN(n8715) );
  NAND2_X1 U5939 ( .A1(n1251), .A2(n3121), .ZN(n24154) );
  OR2_X1 U5942 ( .A1(n7164), .A2(n7320), .ZN(n3167) );
  NAND2_X1 U5983 ( .A1(n3809), .A2(n3808), .ZN(n19962) );
  NAND2_X1 U5984 ( .A1(n28279), .A2(n28737), .ZN(n23842) );
  NOR2_X1 U5991 ( .A1(n23822), .A2(n23821), .ZN(n28279) );
  OR2_X1 U5997 ( .A1(n5918), .A2(n14039), .ZN(n59) );
  NAND3_X1 U6024 ( .A1(n16940), .A2(n211), .A3(n16939), .ZN(n42) );
  OAI22_X1 U6037 ( .A1(n8268), .A2(n8267), .B1(n341), .B2(n8270), .ZN(n8272)
         );
  XNOR2_X1 U6180 ( .A(n28280), .B(n26681), .ZN(Ciphertext[129]) );
  NAND3_X1 U6192 ( .A1(n3561), .A2(n26678), .A3(n6902), .ZN(n28280) );
  NAND2_X1 U6230 ( .A1(n1355), .A2(n28281), .ZN(n1884) );
  NAND3_X1 U6271 ( .A1(n24422), .A2(n24421), .A3(n24517), .ZN(n903) );
  NAND2_X1 U6394 ( .A1(n11774), .A2(n10497), .ZN(n28282) );
  INV_X1 U6411 ( .A(n10716), .ZN(n28283) );
  NAND2_X1 U6463 ( .A1(n26574), .A2(n28286), .ZN(n28285) );
  INV_X1 U6484 ( .A(n26575), .ZN(n28286) );
  NAND2_X1 U6524 ( .A1(n3803), .A2(n3802), .ZN(n3800) );
  NAND2_X1 U6526 ( .A1(n8438), .A2(n224), .ZN(n8441) );
  NAND2_X1 U6536 ( .A1(n28184), .A2(n28287), .ZN(n5477) );
  NAND2_X1 U6559 ( .A1(n400), .A2(n27703), .ZN(n28288) );
  NAND2_X1 U6561 ( .A1(n27701), .A2(n27704), .ZN(n28289) );
  NAND2_X1 U6579 ( .A1(n5651), .A2(n5652), .ZN(n5650) );
  NAND2_X1 U6590 ( .A1(n7932), .A2(n7613), .ZN(n8310) );
  NAND3_X1 U6604 ( .A1(n28290), .A2(n20901), .A3(n5830), .ZN(n5014) );
  NAND2_X1 U6684 ( .A1(n20896), .A2(n21426), .ZN(n28290) );
  NAND2_X1 U6718 ( .A1(n28291), .A2(n15288), .ZN(n1392) );
  NAND2_X1 U6766 ( .A1(n1394), .A2(n756), .ZN(n28291) );
  NAND2_X1 U6795 ( .A1(n29023), .A2(n17592), .ZN(n28292) );
  AOI22_X1 U6830 ( .A1(n26981), .A2(n27636), .B1(n26982), .B2(n27638), .ZN(
        n26983) );
  NAND2_X1 U6852 ( .A1(n8271), .A2(n8270), .ZN(n7210) );
  NAND2_X1 U6855 ( .A1(n18490), .A2(n18488), .ZN(n18291) );
  NAND2_X1 U6872 ( .A1(n52), .A2(n54), .ZN(n51) );
  XNOR2_X1 U7082 ( .A(n21817), .B(n22882), .ZN(n21979) );
  NAND2_X1 U7162 ( .A1(n2250), .A2(n8784), .ZN(n1566) );
  INV_X1 U7243 ( .A(n7775), .ZN(n28692) );
  OAI22_X1 U7251 ( .A1(n27418), .A2(n27429), .B1(n27428), .B2(n27427), .ZN(
        n26669) );
  XNOR2_X1 U7254 ( .A(n13432), .B(n12919), .ZN(n12921) );
  OAI21_X2 U7340 ( .B1(n11748), .B2(n6432), .A(n3281), .ZN(n13432) );
  NOR2_X1 U7353 ( .A1(n20251), .A2(n20252), .ZN(n28295) );
  INV_X1 U7389 ( .A(n11271), .ZN(n652) );
  NAND2_X1 U7400 ( .A1(n279), .A2(n11038), .ZN(n11271) );
  OAI21_X1 U7433 ( .B1(n8720), .B2(n8718), .A(n28296), .ZN(n8413) );
  NAND2_X1 U7458 ( .A1(n8718), .A2(n8788), .ZN(n28296) );
  OAI21_X1 U7468 ( .B1(n28298), .B2(n28532), .A(n28297), .ZN(n25596) );
  NAND2_X1 U7470 ( .A1(n25575), .A2(n28532), .ZN(n28297) );
  INV_X1 U7520 ( .A(n26996), .ZN(n28298) );
  NAND2_X1 U7521 ( .A1(n11574), .A2(n12264), .ZN(n5963) );
  AND3_X2 U7546 ( .A1(n11041), .A2(n11040), .A3(n11042), .ZN(n11574) );
  NAND3_X1 U7579 ( .A1(n21069), .A2(n22403), .A3(n28299), .ZN(n22830) );
  NAND2_X1 U7605 ( .A1(n28301), .A2(n28300), .ZN(n28299) );
  NOR2_X1 U7635 ( .A1(n22402), .A2(n22404), .ZN(n28300) );
  NAND2_X1 U7637 ( .A1(n27715), .A2(n1826), .ZN(n27684) );
  NAND4_X2 U7645 ( .A1(n28302), .A2(n3512), .A3(n1522), .A4(n3514), .ZN(n26011) );
  NAND2_X1 U7678 ( .A1(n28419), .A2(n24368), .ZN(n28302) );
  XNOR2_X1 U7684 ( .A(n2813), .B(n28303), .ZN(n26230) );
  INV_X1 U7702 ( .A(n2812), .ZN(n28303) );
  NAND2_X1 U7711 ( .A1(n27977), .A2(n28456), .ZN(n28355) );
  NAND2_X1 U7756 ( .A1(n18433), .A2(n18430), .ZN(n17815) );
  OAI21_X2 U7779 ( .B1(n17218), .B2(n17217), .A(n17216), .ZN(n18430) );
  NAND2_X1 U7782 ( .A1(n2576), .A2(n6023), .ZN(n14936) );
  BUF_X1 U7817 ( .A(n22991), .Z(n23180) );
  NAND2_X1 U7837 ( .A1(n15040), .A2(n14517), .ZN(n28305) );
  NAND3_X1 U7852 ( .A1(n5811), .A2(n14971), .A3(n14793), .ZN(n5810) );
  NOR2_X2 U7871 ( .A1(n28307), .A2(n5201), .ZN(n18114) );
  OAI21_X1 U7916 ( .B1(n1708), .B2(n5203), .A(n853), .ZN(n28307) );
  NAND2_X1 U7920 ( .A1(n4419), .A2(n4420), .ZN(n28308) );
  OAI21_X1 U7973 ( .B1(n27711), .B2(n27714), .A(n26146), .ZN(n26145) );
  NAND2_X1 U8011 ( .A1(n27725), .A2(n27711), .ZN(n26146) );
  AND2_X1 U8018 ( .A1(n14400), .A2(n29628), .ZN(n13962) );
  OAI21_X1 U8019 ( .B1(n6128), .B2(n16790), .A(n28309), .ZN(n6126) );
  NAND3_X1 U8027 ( .A1(n28768), .A2(n17421), .A3(n17012), .ZN(n28309) );
  NOR2_X1 U8052 ( .A1(n15222), .A2(n15223), .ZN(n5238) );
  NAND2_X1 U8060 ( .A1(n10940), .A2(n10942), .ZN(n10702) );
  XNOR2_X1 U8073 ( .A(n13442), .B(n13443), .ZN(n28311) );
  NOR2_X1 U8074 ( .A1(n21349), .A2(n28312), .ZN(n21351) );
  NAND2_X1 U8080 ( .A1(n21346), .A2(n21347), .ZN(n28312) );
  NAND2_X1 U8094 ( .A1(n6314), .A2(n21698), .ZN(n21347) );
  NAND2_X1 U8095 ( .A1(n14677), .A2(n3315), .ZN(n6681) );
  NAND2_X1 U8101 ( .A1(n14902), .A2(n15097), .ZN(n14677) );
  NAND2_X1 U8103 ( .A1(n28313), .A2(n18078), .ZN(n18080) );
  OAI22_X1 U8106 ( .A1(n18076), .A2(n18075), .B1(n18074), .B2(n5814), .ZN(
        n28313) );
  NAND2_X1 U8110 ( .A1(n24557), .A2(n24633), .ZN(n24558) );
  NAND2_X1 U8111 ( .A1(n24461), .A2(n28314), .ZN(n24462) );
  AND2_X1 U8112 ( .A1(n24812), .A2(n24809), .ZN(n28314) );
  BUF_X2 U8123 ( .A(n21729), .Z(n1930) );
  AND3_X2 U8143 ( .A1(n6518), .A2(n6519), .A3(n11542), .ZN(n13273) );
  NAND2_X1 U8164 ( .A1(n28316), .A2(n28315), .ZN(n23921) );
  NAND2_X1 U8187 ( .A1(n6740), .A2(n24583), .ZN(n28316) );
  NAND2_X1 U8223 ( .A1(n24592), .A2(n831), .ZN(n24142) );
  OAI21_X1 U8282 ( .B1(n4370), .B2(n7977), .A(n7976), .ZN(n7978) );
  NAND2_X1 U8297 ( .A1(n28320), .A2(n28319), .ZN(n26069) );
  NAND2_X1 U8298 ( .A1(n401), .A2(n28229), .ZN(n28319) );
  NAND2_X1 U8326 ( .A1(n26052), .A2(n28180), .ZN(n28320) );
  XNOR2_X1 U8349 ( .A(n28321), .B(n22841), .ZN(n23289) );
  XNOR2_X1 U8351 ( .A(n22839), .B(n22838), .ZN(n28321) );
  NAND2_X1 U8376 ( .A1(n28322), .A2(n14294), .ZN(n14296) );
  NAND3_X1 U8403 ( .A1(n5198), .A2(n15154), .A3(n5199), .ZN(n5197) );
  INV_X1 U8427 ( .A(n520), .ZN(n5690) );
  NAND2_X1 U8429 ( .A1(n28324), .A2(n2938), .ZN(n2442) );
  NAND2_X1 U8431 ( .A1(n2937), .A2(n23655), .ZN(n28324) );
  NAND3_X1 U8475 ( .A1(n772), .A2(n1458), .A3(n770), .ZN(n25205) );
  OR2_X1 U8481 ( .A1(n2096), .A2(n20170), .ZN(n4640) );
  NAND3_X1 U8514 ( .A1(n27621), .A2(n27620), .A3(n1912), .ZN(n1186) );
  NAND3_X1 U8516 ( .A1(n29126), .A2(n23619), .A3(n23270), .ZN(n23271) );
  NAND3_X1 U8523 ( .A1(n7939), .A2(n7657), .A3(n8301), .ZN(n7658) );
  NAND2_X1 U8538 ( .A1(n24484), .A2(n24483), .ZN(n967) );
  NAND2_X1 U8598 ( .A1(n2283), .A2(n28329), .ZN(n10270) );
  NAND2_X1 U8604 ( .A1(n10872), .A2(n11219), .ZN(n28329) );
  AOI21_X2 U8608 ( .B1(n28331), .B2(n23591), .A(n28330), .ZN(n25785) );
  NAND2_X1 U8609 ( .A1(n23575), .A2(n2079), .ZN(n28331) );
  NAND3_X1 U8610 ( .A1(n14379), .A2(n14005), .A3(n14007), .ZN(n6106) );
  XNOR2_X2 U8616 ( .A(n12247), .B(n12248), .ZN(n14259) );
  NAND2_X1 U8658 ( .A1(n28333), .A2(n11338), .ZN(n28332) );
  NAND2_X1 U8710 ( .A1(n11336), .A2(n11176), .ZN(n28333) );
  NAND2_X1 U8714 ( .A1(n11178), .A2(n10830), .ZN(n28334) );
  NAND2_X1 U8716 ( .A1(n14550), .A2(n14549), .ZN(n15476) );
  AND2_X2 U8744 ( .A1(n28335), .A2(n87), .ZN(n9233) );
  NAND2_X1 U8758 ( .A1(n6963), .A2(n6962), .ZN(n28335) );
  NAND2_X1 U8771 ( .A1(n471), .A2(n24972), .ZN(n1251) );
  NAND2_X1 U8775 ( .A1(n10694), .A2(n10985), .ZN(n10695) );
  NAND2_X1 U8821 ( .A1(n6704), .A2(n28336), .ZN(n11599) );
  NAND2_X1 U8822 ( .A1(n8064), .A2(n582), .ZN(n6704) );
  NAND2_X1 U8907 ( .A1(n17379), .A2(n17179), .ZN(n17177) );
  NOR2_X1 U8921 ( .A1(n26953), .A2(n26954), .ZN(n28337) );
  OR2_X1 U8927 ( .A1(n7145), .A2(n7146), .ZN(n28674) );
  NAND2_X1 U8941 ( .A1(n6284), .A2(n6285), .ZN(n28339) );
  NOR2_X1 U8959 ( .A1(n28094), .A2(n28340), .ZN(n26764) );
  NAND2_X1 U8972 ( .A1(n29056), .A2(n28111), .ZN(n28340) );
  NAND2_X1 U9030 ( .A1(n27219), .A2(n27572), .ZN(n28341) );
  XNOR2_X2 U9065 ( .A(n12617), .B(n12618), .ZN(n14295) );
  NAND2_X1 U9125 ( .A1(n5624), .A2(n28343), .ZN(n26682) );
  AOI21_X1 U9184 ( .B1(n26788), .B2(n1872), .A(n28344), .ZN(n28343) );
  AND2_X1 U9195 ( .A1(n26912), .A2(n28423), .ZN(n28344) );
  NAND2_X1 U9225 ( .A1(n14487), .A2(n14481), .ZN(n14169) );
  OAI211_X1 U9237 ( .C1(n3976), .C2(n14761), .A(n15055), .B(n28345), .ZN(n3979) );
  NAND2_X1 U9246 ( .A1(n4162), .A2(n14761), .ZN(n28345) );
  NAND2_X1 U9309 ( .A1(n507), .A2(n20133), .ZN(n19903) );
  NAND2_X1 U9401 ( .A1(n85), .A2(n27672), .ZN(n28347) );
  NAND2_X1 U9405 ( .A1(n28348), .A2(n18658), .ZN(n20966) );
  OAI21_X1 U9435 ( .B1(n20559), .B2(n18650), .A(n20563), .ZN(n28348) );
  AND2_X1 U9453 ( .A1(n9421), .A2(n8327), .ZN(n1386) );
  NAND3_X1 U9487 ( .A1(n24261), .A2(n24503), .A3(n24801), .ZN(n24262) );
  AND2_X2 U9527 ( .A1(n7259), .A2(n3683), .ZN(n9562) );
  INV_X1 U9597 ( .A(n12512), .ZN(n28349) );
  NOR2_X2 U9609 ( .A1(n2655), .A2(n10102), .ZN(n12512) );
  NAND2_X1 U9686 ( .A1(n14299), .A2(n13816), .ZN(n28351) );
  OR2_X1 U9740 ( .A1(n430), .A2(n12991), .ZN(n28677) );
  NAND2_X1 U9743 ( .A1(n24814), .A2(n24812), .ZN(n2246) );
  NAND3_X1 U9784 ( .A1(n23332), .A2(n23768), .A3(n28354), .ZN(n28353) );
  OAI21_X1 U9799 ( .B1(n21012), .B2(n21443), .A(n20833), .ZN(n20836) );
  OAI21_X1 U9815 ( .B1(n27977), .B2(n29021), .A(n28355), .ZN(n26637) );
  OR2_X2 U9829 ( .A1(n6060), .A2(n28357), .ZN(n9073) );
  AOI21_X1 U9833 ( .B1(n7430), .B2(n7431), .A(n8234), .ZN(n28357) );
  XNOR2_X1 U9924 ( .A(n28359), .B(n18579), .ZN(n18834) );
  XNOR2_X1 U9971 ( .A(n18576), .B(n19693), .ZN(n28359) );
  OAI21_X1 U9982 ( .B1(n4819), .B2(n26174), .A(n28360), .ZN(n4817) );
  NAND3_X1 U10020 ( .A1(n26172), .A2(n26917), .A3(n26919), .ZN(n28360) );
  NAND3_X1 U10062 ( .A1(n24422), .A2(n24515), .A3(n24421), .ZN(n28361) );
  NAND3_X1 U10126 ( .A1(n23871), .A2(n23870), .A3(n24514), .ZN(n28362) );
  MUX2_X1 U10141 ( .A(n12280), .B(n11357), .S(n12404), .Z(n11358) );
  NAND2_X1 U10147 ( .A1(n12281), .A2(n12407), .ZN(n12404) );
  OR2_X1 U10193 ( .A1(n10667), .A2(n11077), .ZN(n28364) );
  NAND2_X1 U10198 ( .A1(n28722), .A2(n14109), .ZN(n14517) );
  NAND2_X1 U10199 ( .A1(n28218), .A2(n439), .ZN(n28365) );
  NAND4_X2 U10235 ( .A1(n24319), .A2(n28369), .A3(n28368), .A4(n28367), .ZN(
        n25780) );
  NAND2_X1 U10255 ( .A1(n24317), .A2(n24316), .ZN(n28367) );
  NAND2_X1 U10259 ( .A1(n28227), .A2(n24072), .ZN(n28368) );
  NAND2_X1 U10296 ( .A1(n24315), .A2(n24669), .ZN(n28369) );
  NAND2_X1 U10299 ( .A1(n17771), .A2(n17772), .ZN(n18019) );
  NAND2_X1 U10300 ( .A1(n9124), .A2(n8899), .ZN(n1651) );
  NAND3_X1 U10311 ( .A1(n618), .A2(n7521), .A3(n8030), .ZN(n8031) );
  NAND3_X1 U10335 ( .A1(n149), .A2(n2940), .A3(n2939), .ZN(n851) );
  NAND2_X1 U10347 ( .A1(n28371), .A2(n485), .ZN(n1676) );
  OAI22_X1 U10360 ( .A1(n28626), .A2(n23417), .B1(n480), .B2(n23416), .ZN(
        n28371) );
  NAND2_X1 U10424 ( .A1(n8008), .A2(n8504), .ZN(n28372) );
  AND2_X1 U10504 ( .A1(n19827), .A2(n20311), .ZN(n5826) );
  NAND2_X1 U10526 ( .A1(n6752), .A2(n21495), .ZN(n21127) );
  NAND2_X1 U10586 ( .A1(n28377), .A2(n28376), .ZN(n27214) );
  NAND2_X1 U10587 ( .A1(n27209), .A2(n27210), .ZN(n28376) );
  NAND2_X1 U10601 ( .A1(n27211), .A2(n27038), .ZN(n28377) );
  INV_X1 U10602 ( .A(n27209), .ZN(n28378) );
  NAND2_X1 U10665 ( .A1(n28381), .A2(n28379), .ZN(n10218) );
  INV_X1 U10704 ( .A(n28380), .ZN(n28379) );
  OAI21_X1 U10711 ( .B1(n9000), .B2(n329), .A(n9001), .ZN(n28380) );
  OAI211_X1 U10728 ( .C1(n329), .C2(n9202), .A(n8779), .B(n28862), .ZN(n28381)
         );
  NAND2_X1 U10812 ( .A1(n25470), .A2(n25471), .ZN(n28670) );
  NAND2_X1 U10852 ( .A1(n18835), .A2(n29582), .ZN(n28383) );
  NAND2_X1 U10859 ( .A1(n18836), .A2(n29315), .ZN(n28384) );
  NAND2_X1 U10862 ( .A1(n4672), .A2(n23835), .ZN(n6557) );
  INV_X1 U10889 ( .A(n10844), .ZN(n1812) );
  NAND2_X1 U10895 ( .A1(n11272), .A2(n11269), .ZN(n10844) );
  XNOR2_X1 U10911 ( .A(n24402), .B(n24401), .ZN(n28385) );
  NAND3_X1 U10968 ( .A1(n3390), .A2(n6634), .A3(n6633), .ZN(n28386) );
  NAND2_X1 U10969 ( .A1(n21262), .A2(n3318), .ZN(n28387) );
  XNOR2_X1 U10970 ( .A(n28388), .B(n22562), .ZN(n22564) );
  XOR2_X1 U10981 ( .A(n22561), .B(n22690), .Z(n28388) );
  NAND2_X1 U10991 ( .A1(n21262), .A2(n3318), .ZN(n22561) );
  XOR2_X1 U11015 ( .A(n10306), .B(n8477), .Z(n8479) );
  NAND2_X1 U11031 ( .A1(n23972), .A2(n24209), .ZN(n4754) );
  XNOR2_X1 U11051 ( .A(n22231), .B(n22230), .ZN(n28390) );
  INV_X1 U11088 ( .A(n23193), .ZN(n28391) );
  XNOR2_X1 U11105 ( .A(n24868), .B(n24869), .ZN(n28392) );
  AND2_X1 U11127 ( .A1(n6125), .A2(n6124), .ZN(n28393) );
  AND2_X1 U11191 ( .A1(n6125), .A2(n6124), .ZN(n28394) );
  AND2_X1 U11229 ( .A1(n6125), .A2(n6124), .ZN(n27208) );
  OAI21_X1 U11267 ( .B1(n14888), .B2(n14889), .A(n14887), .ZN(n28395) );
  XOR2_X1 U11276 ( .A(n16555), .B(n16026), .Z(n16030) );
  OAI21_X1 U11295 ( .B1(n14888), .B2(n14889), .A(n14887), .ZN(n3792) );
  AOI21_X1 U11307 ( .B1(n18346), .B2(n514), .A(n18344), .ZN(n17950) );
  NOR2_X1 U11343 ( .A1(n27695), .A2(n27694), .ZN(n28396) );
  XOR2_X1 U11363 ( .A(n28397), .B(n3321), .Z(Ciphertext[136]) );
  NAND3_X1 U11377 ( .A1(n2765), .A2(n2764), .A3(n2763), .ZN(n28397) );
  MUX2_X1 U11388 ( .A(n28399), .B(n28400), .S(n27701), .Z(n28398) );
  OR2_X1 U11434 ( .A1(n27702), .A2(n27700), .ZN(n28399) );
  OR2_X1 U11441 ( .A1(n27703), .A2(n27161), .ZN(n28400) );
  NOR2_X1 U11459 ( .A1(n6277), .A2(n6278), .ZN(n28401) );
  NOR2_X1 U11478 ( .A1(n24116), .A2(n24115), .ZN(n28402) );
  NOR2_X1 U11498 ( .A1(n1008), .A2(n26324), .ZN(n28403) );
  NOR2_X1 U11499 ( .A1(n24116), .A2(n24115), .ZN(n25463) );
  OR2_X1 U11509 ( .A1(n3283), .A2(n18376), .ZN(n28404) );
  XOR2_X1 U11510 ( .A(n13420), .B(n13067), .Z(n12943) );
  XNOR2_X1 U11532 ( .A(n9394), .B(n9395), .ZN(n11004) );
  XNOR2_X1 U11593 ( .A(n9408), .B(n9407), .ZN(n1308) );
  XNOR2_X1 U11628 ( .A(n19282), .B(n19281), .ZN(n28408) );
  NAND2_X1 U11658 ( .A1(n3758), .A2(n1050), .ZN(n28409) );
  NAND2_X1 U11699 ( .A1(n3758), .A2(n1050), .ZN(n22887) );
  NAND3_X1 U11716 ( .A1(n664), .A2(n25971), .A3(n663), .ZN(n28411) );
  NAND3_X1 U11724 ( .A1(n664), .A2(n25971), .A3(n663), .ZN(n28016) );
  CLKBUF_X1 U11729 ( .A(Key[44]), .Z(n27894) );
  NAND2_X1 U11761 ( .A1(n28412), .A2(n28413), .ZN(n994) );
  OR2_X1 U11837 ( .A1(n17659), .A2(n18467), .ZN(n28412) );
  OR2_X1 U11874 ( .A1(n18464), .A2(n1383), .ZN(n28413) );
  BUF_X1 U11875 ( .A(n11739), .Z(n11742) );
  AND2_X1 U11902 ( .A1(n6025), .A2(n6024), .ZN(n28414) );
  XOR2_X1 U11908 ( .A(n19269), .B(n18858), .Z(n18861) );
  AOI22_X1 U11971 ( .A1(n456), .A2(n26436), .B1(n26937), .B2(n26936), .ZN(
        n5546) );
  OAI21_X1 U12005 ( .B1(n6091), .B2(n23419), .A(n23063), .ZN(n24717) );
  XNOR2_X1 U12012 ( .A(n19545), .B(n19544), .ZN(n28417) );
  XNOR2_X1 U12023 ( .A(n6846), .B(n6847), .ZN(n23280) );
  NOR2_X1 U12025 ( .A1(n24369), .A2(n23897), .ZN(n28419) );
  NAND2_X1 U12026 ( .A1(n20605), .A2(n20606), .ZN(n21599) );
  XNOR2_X1 U12029 ( .A(n25862), .B(n25861), .ZN(n28631) );
  AND2_X1 U12038 ( .A1(n28420), .A2(n23211), .ZN(n21978) );
  OR2_X1 U12041 ( .A1(n23577), .A2(n23603), .ZN(n28420) );
  INV_X1 U12046 ( .A(n26937), .ZN(n28421) );
  AND2_X1 U12076 ( .A1(n25159), .A2(n25158), .ZN(n28422) );
  XOR2_X1 U12101 ( .A(n25383), .B(n25384), .Z(n28423) );
  MUX2_X1 U12105 ( .A(n26805), .B(n26806), .S(n2438), .Z(n26807) );
  OAI21_X1 U12134 ( .B1(n480), .B2(n22808), .A(n22807), .ZN(n24556) );
  INV_X1 U12149 ( .A(n24382), .ZN(n28424) );
  XNOR2_X1 U12150 ( .A(n28425), .B(n28426), .ZN(n5306) );
  XNOR2_X1 U12169 ( .A(n25743), .B(n25744), .ZN(n28425) );
  XOR2_X1 U12192 ( .A(n25747), .B(n25746), .Z(n28426) );
  OAI21_X1 U12222 ( .B1(n23350), .B2(n4429), .A(n23349), .ZN(n24665) );
  XNOR2_X1 U12318 ( .A(n22070), .B(n22071), .ZN(n23700) );
  BUF_X1 U12397 ( .A(n27590), .Z(n28429) );
  INV_X1 U12418 ( .A(n27732), .ZN(n28430) );
  XOR2_X1 U12444 ( .A(n9648), .B(n9899), .Z(n10156) );
  XOR2_X1 U12477 ( .A(n13565), .B(n12834), .Z(n12381) );
  XOR2_X1 U12482 ( .A(n22070), .B(n22071), .Z(n28431) );
  OR2_X1 U12483 ( .A1(n24560), .A2(n23990), .ZN(n28687) );
  XOR2_X1 U12515 ( .A(n22093), .B(n28387), .Z(n28432) );
  AOI21_X1 U12518 ( .B1(n219), .B2(n28679), .A(n28678), .ZN(n28433) );
  AOI21_X1 U12519 ( .B1(n219), .B2(n28679), .A(n28678), .ZN(n4263) );
  XOR2_X1 U12520 ( .A(n24446), .B(n24445), .Z(n28434) );
  BUF_X1 U12525 ( .A(n27460), .Z(n28435) );
  OAI21_X1 U12527 ( .B1(n26159), .B2(n26562), .A(n26158), .ZN(n27460) );
  BUF_X1 U12548 ( .A(n11787), .Z(n28436) );
  XOR2_X1 U12551 ( .A(n25854), .B(n25853), .Z(n28437) );
  OAI21_X1 U12558 ( .B1(n10729), .B2(n10730), .A(n10728), .ZN(n11787) );
  MUX2_X2 U12574 ( .A(n26783), .B(n26784), .S(n454), .Z(n27282) );
  AND3_X1 U12604 ( .A1(n27009), .A2(n27008), .A3(n27007), .ZN(n28438) );
  AND3_X1 U12605 ( .A1(n27009), .A2(n27008), .A3(n27007), .ZN(n28439) );
  AOI22_X1 U12620 ( .A1(n18546), .A2(n19967), .B1(n18547), .B2(n20123), .ZN(
        n21343) );
  AND3_X1 U12634 ( .A1(n6755), .A2(n5391), .A3(n5390), .ZN(n28441) );
  NAND2_X1 U12641 ( .A1(n5779), .A2(n5780), .ZN(n28442) );
  XOR2_X1 U12708 ( .A(n12383), .B(n12087), .Z(n12119) );
  XNOR2_X1 U12714 ( .A(n21882), .B(n21883), .ZN(n28444) );
  AND4_X1 U12740 ( .A1(n27135), .A2(n27134), .A3(n27133), .A4(n27132), .ZN(
        n28445) );
  XNOR2_X1 U12759 ( .A(n21882), .B(n21883), .ZN(n23687) );
  XNOR2_X1 U12786 ( .A(n25502), .B(n25501), .ZN(n27052) );
  CLKBUF_X1 U12804 ( .A(n22205), .Z(n28514) );
  NOR2_X1 U12832 ( .A1(n17817), .A2(n17816), .ZN(n28447) );
  INV_X1 U12847 ( .A(n20049), .ZN(n28448) );
  XNOR2_X1 U12848 ( .A(n22053), .B(n22052), .ZN(n22600) );
  XNOR2_X1 U12858 ( .A(n25823), .B(n25824), .ZN(n26840) );
  NAND3_X1 U12864 ( .A1(n2299), .A2(n19803), .A3(n4225), .ZN(n28449) );
  BUF_X1 U12952 ( .A(n1534), .Z(n28451) );
  NAND2_X1 U12959 ( .A1(n25001), .A2(n25003), .ZN(n894) );
  XNOR2_X1 U12997 ( .A(n25719), .B(n25718), .ZN(n28452) );
  OAI211_X1 U12999 ( .C1(n27073), .C2(n27072), .A(n3786), .B(n3785), .ZN(
        n28453) );
  INV_X1 U13018 ( .A(n16693), .ZN(n18343) );
  XNOR2_X1 U13067 ( .A(n15786), .B(n15785), .ZN(n17541) );
  OAI211_X1 U13070 ( .C1(n29126), .C2(n23626), .A(n5554), .B(n5556), .ZN(
        n28455) );
  OAI211_X1 U13110 ( .C1(n29126), .C2(n23626), .A(n5554), .B(n5556), .ZN(
        n23655) );
  XNOR2_X1 U13133 ( .A(n20872), .B(n20873), .ZN(n28457) );
  XOR2_X1 U13142 ( .A(n25823), .B(n25824), .Z(n28458) );
  XNOR2_X1 U13143 ( .A(n20872), .B(n20873), .ZN(n23686) );
  XNOR2_X1 U13148 ( .A(n25308), .B(n25307), .ZN(n28459) );
  XNOR2_X1 U13187 ( .A(n25308), .B(n25307), .ZN(n26715) );
  INV_X1 U13188 ( .A(n7298), .ZN(n8162) );
  AOI22_X1 U13189 ( .A1(n25632), .A2(n26723), .B1(n26717), .B2(n25631), .ZN(
        n27408) );
  BUF_X1 U13202 ( .A(n22232), .Z(n28461) );
  OAI22_X1 U13234 ( .A1(n20719), .A2(n28602), .B1(n5622), .B2(n20899), .ZN(
        n22232) );
  AOI21_X1 U13262 ( .B1(n3950), .B2(n14345), .A(n3947), .ZN(n28462) );
  AOI21_X1 U13289 ( .B1(n3950), .B2(n14345), .A(n3947), .ZN(n15175) );
  OR2_X1 U13290 ( .A1(n10828), .A2(n11337), .ZN(n1190) );
  OR2_X1 U13345 ( .A1(n24056), .A2(n5507), .ZN(n24916) );
  NAND2_X1 U13376 ( .A1(n23915), .A2(n985), .ZN(n28465) );
  NAND2_X1 U13385 ( .A1(n985), .A2(n23915), .ZN(n26060) );
  OAI21_X1 U13398 ( .B1(n24857), .B2(n4679), .A(n24856), .ZN(n27646) );
  XOR2_X1 U13400 ( .A(n25697), .B(n26059), .Z(n25458) );
  XOR2_X1 U13417 ( .A(n22218), .B(n22219), .Z(n22712) );
  XNOR2_X1 U13418 ( .A(n1502), .B(n1055), .ZN(n23370) );
  XOR2_X1 U13442 ( .A(n25033), .B(n25032), .Z(n28467) );
  INV_X1 U13466 ( .A(n27203), .ZN(n28468) );
  XOR2_X1 U13547 ( .A(n25098), .B(n25097), .Z(n28470) );
  XNOR2_X1 U13548 ( .A(n25376), .B(n25377), .ZN(n28471) );
  OAI211_X1 U13567 ( .C1(n21011), .C2(n21010), .A(n21009), .B(n2343), .ZN(
        n28472) );
  OAI211_X1 U13598 ( .C1(n21011), .C2(n21010), .A(n21009), .B(n2343), .ZN(
        n22910) );
  XNOR2_X1 U13647 ( .A(n2813), .B(n2812), .ZN(n28473) );
  OR2_X1 U13676 ( .A1(n11322), .A2(n29316), .ZN(n22) );
  INV_X1 U13682 ( .A(n29157), .ZN(n28474) );
  NOR2_X1 U13696 ( .A1(n22178), .A2(n22179), .ZN(n28475) );
  NOR2_X1 U13704 ( .A1(n22178), .A2(n22179), .ZN(n26044) );
  XNOR2_X1 U13710 ( .A(n3596), .B(n25258), .ZN(n26447) );
  XNOR2_X1 U13718 ( .A(n13276), .B(n13275), .ZN(n28478) );
  XNOR2_X1 U13719 ( .A(n18926), .B(n18925), .ZN(n21095) );
  XOR2_X1 U13729 ( .A(n24879), .B(n24878), .Z(n28480) );
  OAI21_X1 U13874 ( .B1(n23232), .B2(n1862), .A(n23231), .ZN(n28481) );
  XOR2_X1 U13875 ( .A(n24574), .B(n24573), .Z(n28482) );
  AND2_X1 U13879 ( .A1(n9207), .A2(n41), .ZN(n9437) );
  NAND4_X1 U13898 ( .A1(n6425), .A2(n6427), .A3(n6426), .A4(n20216), .ZN(
        n28483) );
  NAND4_X1 U13917 ( .A1(n6425), .A2(n6427), .A3(n6426), .A4(n20216), .ZN(
        n22568) );
  NOR2_X1 U13925 ( .A1(n23967), .A2(n23966), .ZN(n28485) );
  XNOR2_X1 U13935 ( .A(n22121), .B(n22120), .ZN(n23725) );
  NOR2_X1 U13936 ( .A1(n23967), .A2(n23966), .ZN(n26094) );
  NOR2_X1 U13969 ( .A1(n21112), .A2(n4755), .ZN(n28486) );
  XOR2_X1 U13970 ( .A(n22159), .B(n21836), .Z(n21840) );
  NOR2_X1 U13973 ( .A1(n21112), .A2(n4755), .ZN(n22756) );
  XNOR2_X1 U13977 ( .A(n26087), .B(n26088), .ZN(n28487) );
  XNOR2_X1 U13980 ( .A(n26087), .B(n26088), .ZN(n27141) );
  XNOR2_X1 U13982 ( .A(n25561), .B(n25560), .ZN(n26632) );
  BUF_X1 U14077 ( .A(n27972), .Z(n27970) );
  INV_X1 U14098 ( .A(n4950), .ZN(n28738) );
  OR2_X1 U14099 ( .A1(n15787), .A2(n17542), .ZN(n16940) );
  OAI211_X1 U14107 ( .C1(n9167), .C2(n9163), .A(n8317), .B(n8316), .ZN(n9921)
         );
  NAND2_X1 U14130 ( .A1(n1810), .A2(n20276), .ZN(n28492) );
  OR2_X1 U14274 ( .A1(n17415), .A2(n17413), .ZN(n17301) );
  AND2_X1 U14306 ( .A1(n25359), .A2(n25357), .ZN(n28494) );
  XNOR2_X1 U14316 ( .A(n9270), .B(n9269), .ZN(n28495) );
  CLKBUF_X1 U14322 ( .A(n25187), .Z(n28496) );
  XNOR2_X1 U14340 ( .A(n9270), .B(n9269), .ZN(n10941) );
  NOR2_X1 U14423 ( .A1(n4466), .A2(n4465), .ZN(n28499) );
  NAND2_X1 U14510 ( .A1(n7482), .A2(n7483), .ZN(n9080) );
  XNOR2_X1 U14511 ( .A(n16871), .B(n16870), .ZN(n28501) );
  XNOR2_X1 U14537 ( .A(n24088), .B(n24089), .ZN(n28503) );
  NAND2_X1 U14625 ( .A1(n23293), .A2(n4175), .ZN(n3797) );
  NAND3_X1 U14633 ( .A1(n5427), .A2(n24030), .A3(n24031), .ZN(n25703) );
  XOR2_X1 U14666 ( .A(n24931), .B(n24930), .Z(n28504) );
  OR2_X1 U14747 ( .A1(n1912), .A2(n27630), .ZN(n28505) );
  MUX2_X2 U14786 ( .A(n26360), .B(n26359), .S(n26358), .Z(n27630) );
  XOR2_X1 U14843 ( .A(n5702), .B(n5703), .Z(n28506) );
  INV_X1 U14848 ( .A(n14358), .ZN(n28507) );
  OR2_X1 U14907 ( .A1(n29037), .A2(n13672), .ZN(n2965) );
  XNOR2_X1 U15011 ( .A(n5703), .B(n5702), .ZN(n23801) );
  CLKBUF_X1 U15032 ( .A(n20573), .Z(n28508) );
  XNOR2_X1 U15033 ( .A(n18609), .B(n19683), .ZN(n20573) );
  AND2_X1 U15037 ( .A1(n27302), .A2(n27303), .ZN(n28510) );
  MUX2_X2 U15073 ( .A(n25316), .B(n25315), .S(n29560), .Z(n27364) );
  XNOR2_X1 U15128 ( .A(n24918), .B(n24919), .ZN(n28513) );
  AOI22_X1 U15131 ( .A1(n23608), .A2(n23607), .B1(n23605), .B2(n23606), .ZN(
        n24790) );
  CLKBUF_X1 U15132 ( .A(n20333), .Z(n28515) );
  XNOR2_X1 U15138 ( .A(n19288), .B(n19287), .ZN(n20333) );
  OAI22_X1 U15238 ( .A1(n23108), .A2(n23107), .B1(n23106), .B2(n486), .ZN(
        n24211) );
  OAI21_X1 U15286 ( .B1(n14004), .B2(n13575), .A(n13574), .ZN(n28518) );
  OAI21_X1 U15305 ( .B1(n14004), .B2(n13575), .A(n13574), .ZN(n14942) );
  AOI21_X1 U15309 ( .B1(n24177), .B2(n24178), .A(n24176), .ZN(n28520) );
  XNOR2_X1 U15315 ( .A(n25766), .B(n25765), .ZN(n28521) );
  AOI21_X1 U15373 ( .B1(n24177), .B2(n24178), .A(n24176), .ZN(n25445) );
  XNOR2_X2 U15492 ( .A(n24841), .B(n24840), .ZN(n26426) );
  NOR2_X1 U15493 ( .A1(n6599), .A2(n23797), .ZN(n28522) );
  NOR2_X1 U15508 ( .A1(n6599), .A2(n23797), .ZN(n28523) );
  NOR2_X1 U15511 ( .A1(n6599), .A2(n23797), .ZN(n24803) );
  OAI211_X1 U15516 ( .C1(n23694), .C2(n23135), .A(n6442), .B(n6441), .ZN(
        n24409) );
  XNOR2_X1 U15528 ( .A(n24198), .B(n24199), .ZN(n28525) );
  XNOR2_X1 U15535 ( .A(n24198), .B(n24199), .ZN(n26185) );
  XNOR2_X1 U15572 ( .A(n22022), .B(n22021), .ZN(n28527) );
  OR2_X1 U15617 ( .A1(n5320), .A2(n23255), .ZN(n28528) );
  XNOR2_X1 U15620 ( .A(n22022), .B(n22021), .ZN(n23406) );
  XNOR2_X2 U15625 ( .A(n24625), .B(n24624), .ZN(n26457) );
  NOR2_X1 U15640 ( .A1(n4803), .A2(n174), .ZN(n28530) );
  NOR2_X1 U15722 ( .A1(n4803), .A2(n174), .ZN(n19636) );
  INV_X1 U15759 ( .A(n24697), .ZN(n28531) );
  XNOR2_X1 U15779 ( .A(n25574), .B(n25573), .ZN(n28532) );
  XNOR2_X1 U15804 ( .A(n25574), .B(n25573), .ZN(n26997) );
  XNOR2_X1 U15828 ( .A(n24882), .B(n24881), .ZN(n28536) );
  XNOR2_X1 U15995 ( .A(n19416), .B(n19415), .ZN(n28538) );
  XNOR2_X1 U15996 ( .A(n19416), .B(n19415), .ZN(n20634) );
  XNOR2_X1 U16017 ( .A(n22210), .B(n22209), .ZN(n23562) );
  OAI211_X1 U16066 ( .C1(n17897), .C2(n18268), .A(n1718), .B(n1716), .ZN(
        n18928) );
  OAI22_X1 U16088 ( .A1(n23889), .A2(n23888), .B1(n23887), .B2(n24434), .ZN(
        n28540) );
  OAI22_X1 U16159 ( .A1(n23889), .A2(n23888), .B1(n23887), .B2(n24434), .ZN(
        n25583) );
  XNOR2_X1 U16245 ( .A(n25129), .B(n25130), .ZN(n26941) );
  XNOR2_X1 U16380 ( .A(n25189), .B(n6789), .ZN(n28542) );
  XNOR2_X1 U16535 ( .A(n25189), .B(n6789), .ZN(n26266) );
  XOR2_X1 U16536 ( .A(n16566), .B(n15256), .Z(n15257) );
  NAND2_X1 U16829 ( .A1(n26243), .A2(n26244), .ZN(n28064) );
  INV_X1 U16831 ( .A(n4599), .ZN(n28544) );
  XNOR2_X1 U16952 ( .A(n25693), .B(n25692), .ZN(n27067) );
  XNOR2_X1 U16961 ( .A(n24170), .B(n24169), .ZN(n28547) );
  XNOR2_X1 U16965 ( .A(n24170), .B(n24169), .ZN(n26182) );
  XNOR2_X1 U17022 ( .A(n25296), .B(n25297), .ZN(n28548) );
  NAND3_X1 U17039 ( .A1(n25664), .A2(n6288), .A3(n25663), .ZN(n28549) );
  NAND3_X1 U17040 ( .A1(n25664), .A2(n6288), .A3(n25663), .ZN(n27355) );
  XOR2_X1 U17051 ( .A(n25901), .B(n26038), .Z(n24885) );
  CLKBUF_X3 U17098 ( .A(n26537), .Z(n27875) );
  XNOR2_X1 U17103 ( .A(n25171), .B(n25170), .ZN(n26949) );
  XOR2_X1 U17208 ( .A(n22466), .B(n22465), .Z(n28551) );
  XNOR2_X1 U17328 ( .A(n19524), .B(n19523), .ZN(n28552) );
  XOR2_X1 U17523 ( .A(n19713), .B(n19712), .Z(n28555) );
  OAI211_X1 U17611 ( .C1(n24743), .C2(n24744), .A(n24742), .B(n24741), .ZN(
        n25825) );
  AOI22_X1 U17664 ( .A1(n14114), .A2(n15116), .B1(n13668), .B2(n1001), .ZN(
        n28557) );
  AOI22_X1 U17689 ( .A1(n14114), .A2(n15116), .B1(n13668), .B2(n1001), .ZN(
        n16039) );
  AOI22_X1 U17776 ( .A1(n17380), .A2(n4295), .B1(n17378), .B2(n17379), .ZN(
        n18708) );
  CLKBUF_X1 U17840 ( .A(n10556), .Z(n28559) );
  BUF_X1 U17841 ( .A(n26481), .Z(n28560) );
  XNOR2_X1 U17844 ( .A(n25217), .B(n25218), .ZN(n26481) );
  OR2_X1 U17856 ( .A1(n7164), .A2(n7770), .ZN(n7323) );
  XNOR2_X1 U17893 ( .A(n24063), .B(n24062), .ZN(n28561) );
  BUF_X1 U17939 ( .A(n26808), .Z(n28562) );
  XNOR2_X1 U17944 ( .A(n24063), .B(n24062), .ZN(n26476) );
  OAI21_X1 U17980 ( .B1(n25321), .B2(n28525), .A(n25320), .ZN(n26808) );
  OR3_X1 U17981 ( .A1(n17259), .A2(n17260), .A3(n17262), .ZN(n3587) );
  XNOR2_X1 U18075 ( .A(n15564), .B(n6929), .ZN(n28564) );
  OR2_X1 U18110 ( .A1(n24512), .A2(n24511), .ZN(n28565) );
  XOR2_X1 U18211 ( .A(n6212), .B(n21728), .Z(n28566) );
  OR2_X1 U18328 ( .A1(n22948), .A2(n22947), .ZN(n28567) );
  NOR2_X2 U18329 ( .A1(n24648), .A2(n24647), .ZN(n25542) );
  XNOR2_X1 U18438 ( .A(n9714), .B(n6916), .ZN(n28568) );
  XNOR2_X1 U18458 ( .A(n19282), .B(n19281), .ZN(n20598) );
  OR2_X1 U18477 ( .A1(n23683), .A2(n23686), .ZN(n3434) );
  XNOR2_X1 U18854 ( .A(n13483), .B(n6651), .ZN(n28569) );
  XNOR2_X1 U18911 ( .A(n21419), .B(n21418), .ZN(n28570) );
  XNOR2_X1 U18915 ( .A(n13483), .B(n6651), .ZN(n14039) );
  XNOR2_X1 U18959 ( .A(n21419), .B(n21418), .ZN(n23343) );
  INV_X1 U18983 ( .A(n17012), .ZN(n16968) );
  NAND2_X1 U18984 ( .A1(n5228), .A2(n17863), .ZN(n28571) );
  NAND2_X1 U19007 ( .A1(n5228), .A2(n17863), .ZN(n19725) );
  XNOR2_X1 U19010 ( .A(n24962), .B(n24961), .ZN(n28572) );
  XNOR2_X1 U19044 ( .A(n24962), .B(n24961), .ZN(n28573) );
  NOR2_X1 U19059 ( .A1(n28226), .A2(n27165), .ZN(n27171) );
  XOR2_X1 U19065 ( .A(n6870), .B(n6869), .Z(n28574) );
  XNOR2_X1 U19131 ( .A(n25830), .B(n25248), .ZN(n28575) );
  OR2_X1 U19284 ( .A1(n20494), .A2(n20493), .ZN(n19867) );
  XOR2_X1 U19386 ( .A(n21689), .B(n21688), .Z(n28577) );
  NAND2_X1 U19419 ( .A1(n3344), .A2(n13988), .ZN(n28579) );
  NAND2_X1 U19477 ( .A1(n3967), .A2(n19798), .ZN(n28580) );
  XNOR2_X1 U19672 ( .A(n22191), .B(n22190), .ZN(n28581) );
  XNOR2_X1 U19699 ( .A(n22191), .B(n22190), .ZN(n28582) );
  XOR2_X1 U19726 ( .A(n25448), .B(n25447), .Z(n28583) );
  XOR2_X1 U19728 ( .A(n22698), .B(n22699), .Z(n22701) );
  BUF_X1 U19805 ( .A(n13566), .Z(n28587) );
  XOR2_X1 U19826 ( .A(n11866), .B(n11865), .Z(n28588) );
  OAI21_X1 U19866 ( .B1(n11863), .B2(n11862), .A(n1526), .ZN(n13566) );
  NAND2_X1 U19871 ( .A1(n3531), .A2(n3530), .ZN(n28589) );
  NAND2_X1 U19942 ( .A1(n3531), .A2(n3530), .ZN(n22762) );
  NOR2_X1 U20053 ( .A1(n26725), .A2(n26724), .ZN(n28591) );
  OAI21_X1 U20146 ( .B1(n24038), .B2(n24039), .A(n24037), .ZN(n27029) );
  XNOR2_X1 U20172 ( .A(n19379), .B(n19378), .ZN(n19641) );
  NAND2_X1 U20226 ( .A1(n6513), .A2(n1223), .ZN(n28593) );
  XOR2_X1 U20358 ( .A(n22598), .B(n22597), .Z(n28594) );
  XOR2_X1 U20400 ( .A(n24905), .B(n24904), .Z(n28595) );
  NOR2_X1 U20423 ( .A1(n23083), .A2(n23082), .ZN(n28596) );
  OAI21_X1 U20425 ( .B1(n14669), .B2(n15304), .A(n14668), .ZN(n28597) );
  INV_X1 U20426 ( .A(n24426), .ZN(n28598) );
  OAI21_X1 U20645 ( .B1(n14669), .B2(n15304), .A(n14668), .ZN(n16470) );
  OAI21_X1 U20745 ( .B1(n23535), .B2(n23534), .A(n6942), .ZN(n24767) );
  NAND2_X1 U20809 ( .A1(n6513), .A2(n1223), .ZN(n26020) );
  XOR2_X1 U20853 ( .A(n25937), .B(n25936), .Z(n28600) );
  XOR2_X1 U20908 ( .A(n12773), .B(n12772), .Z(n28601) );
  BUF_X1 U20940 ( .A(n1925), .Z(n28602) );
  NOR2_X1 U20944 ( .A1(n12185), .A2(n12184), .ZN(n28603) );
  XNOR2_X1 U21033 ( .A(n21300), .B(n21299), .ZN(n28604) );
  XNOR2_X1 U21048 ( .A(n21300), .B(n21299), .ZN(n23676) );
  OR2_X1 U21119 ( .A1(n29629), .A2(n7257), .ZN(n7512) );
  XNOR2_X1 U21125 ( .A(n6977), .B(Key[101]), .ZN(n28605) );
  OR2_X1 U21158 ( .A1(n20480), .A2(n19995), .ZN(n20230) );
  NOR2_X1 U21159 ( .A1(n20357), .A2(n20356), .ZN(n20782) );
  INV_X1 U21237 ( .A(n27242), .ZN(n28607) );
  NOR2_X1 U21290 ( .A1(n3445), .A2(n155), .ZN(n9081) );
  XNOR2_X1 U21318 ( .A(n6891), .B(n9309), .ZN(n10948) );
  XOR2_X1 U21330 ( .A(n19444), .B(n19443), .Z(n28610) );
  INV_X1 U21334 ( .A(n20393), .ZN(n28611) );
  XOR2_X1 U21376 ( .A(n9527), .B(n9526), .Z(n28612) );
  XOR2_X1 U21395 ( .A(n22326), .B(n22414), .Z(n28613) );
  MUX2_X1 U21419 ( .A(n7616), .B(n7615), .S(n29135), .Z(n7617) );
  XNOR2_X1 U21424 ( .A(n7219), .B(Key[128]), .ZN(n28614) );
  XNOR2_X1 U21440 ( .A(n7219), .B(Key[128]), .ZN(n28615) );
  XNOR2_X1 U21463 ( .A(n7219), .B(Key[128]), .ZN(n8256) );
  AND2_X1 U21495 ( .A1(n20573), .A2(n19838), .ZN(n19833) );
  OR2_X1 U21498 ( .A1(n12057), .A2(n12320), .ZN(n28747) );
  XNOR2_X1 U21514 ( .A(n7220), .B(Key[129]), .ZN(n28617) );
  XNOR2_X1 U21549 ( .A(n7220), .B(Key[129]), .ZN(n28618) );
  AOI22_X1 U21550 ( .A1(n20387), .A2(n20386), .B1(n20385), .B2(n20384), .ZN(
        n28619) );
  XNOR2_X1 U21554 ( .A(n7220), .B(Key[129]), .ZN(n8263) );
  AOI22_X1 U21784 ( .A1(n20387), .A2(n20386), .B1(n20385), .B2(n20384), .ZN(
        n21501) );
  XNOR2_X1 U21803 ( .A(n19080), .B(n19081), .ZN(n28620) );
  XNOR2_X1 U21817 ( .A(n19081), .B(n19080), .ZN(n20485) );
  XOR2_X1 U21819 ( .A(n19121), .B(n19120), .Z(n28621) );
  NOR2_X1 U21900 ( .A1(n2205), .A2(n24559), .ZN(n24561) );
  NOR2_X1 U21910 ( .A1(n19656), .A2(n19659), .ZN(n28623) );
  XNOR2_X1 U22058 ( .A(n10125), .B(n10124), .ZN(n28624) );
  XNOR2_X1 U22085 ( .A(n10124), .B(n10125), .ZN(n11210) );
  XOR2_X1 U22105 ( .A(n12897), .B(n12898), .Z(n28625) );
  XNOR2_X1 U22116 ( .A(n22775), .B(n22774), .ZN(n28626) );
  XNOR2_X1 U22120 ( .A(n22775), .B(n22774), .ZN(n2452) );
  XNOR2_X1 U22305 ( .A(n7811), .B(n7812), .ZN(n28627) );
  XNOR2_X1 U22412 ( .A(n7811), .B(n7812), .ZN(n11145) );
  OAI21_X1 U22413 ( .B1(n1777), .B2(n1828), .A(n23094), .ZN(n25190) );
  OAI211_X1 U22509 ( .C1(n23857), .C2(n23856), .A(n841), .B(n840), .ZN(n28630)
         );
  OAI211_X1 U22513 ( .C1(n23857), .C2(n23856), .A(n841), .B(n840), .ZN(n25858)
         );
  XNOR2_X1 U22671 ( .A(n25862), .B(n25861), .ZN(n27118) );
  BUF_X1 U22715 ( .A(n18492), .Z(n28633) );
  AOI22_X1 U22737 ( .A1(n16878), .A2(n15616), .B1(n15615), .B2(n424), .ZN(
        n18492) );
  OAI211_X1 U22764 ( .C1(n9106), .C2(n8512), .A(n9105), .B(n8072), .ZN(n28634)
         );
  OAI211_X1 U22883 ( .C1(n9106), .C2(n8512), .A(n9105), .B(n8072), .ZN(n10145)
         );
  AOI21_X1 U23009 ( .B1(n26632), .B2(n26631), .A(n26630), .ZN(n27997) );
  XNOR2_X1 U23010 ( .A(n18586), .B(n18585), .ZN(n28637) );
  XNOR2_X1 U23015 ( .A(n18586), .B(n18585), .ZN(n19836) );
  XNOR2_X1 U23016 ( .A(n8520), .B(n8519), .ZN(n28638) );
  XOR2_X1 U23067 ( .A(n25496), .B(n25497), .Z(n28639) );
  XNOR2_X1 U23076 ( .A(n8520), .B(n8519), .ZN(n10814) );
  XOR2_X1 U23077 ( .A(n25789), .B(n25788), .Z(n28640) );
  INV_X1 U23081 ( .A(n26546), .ZN(n28641) );
  NOR2_X1 U23091 ( .A1(n27865), .A2(n27872), .ZN(n27327) );
  XNOR2_X1 U23105 ( .A(n24982), .B(n24983), .ZN(n28642) );
  OAI21_X1 U23106 ( .B1(n7161), .B2(n7160), .A(n7159), .ZN(n28643) );
  CLKBUF_X1 U23122 ( .A(n23631), .Z(n28644) );
  OAI21_X1 U23158 ( .B1(n22970), .B2(n22969), .A(n22968), .ZN(n28645) );
  BUF_X1 U23159 ( .A(n26951), .Z(n28646) );
  XNOR2_X1 U23175 ( .A(n12480), .B(n12479), .ZN(n28647) );
  XNOR2_X1 U23205 ( .A(n12480), .B(n12479), .ZN(n28648) );
  INV_X1 U23259 ( .A(n4044), .ZN(n28649) );
  XNOR2_X1 U23318 ( .A(n12480), .B(n12479), .ZN(n14444) );
  NOR2_X1 U23368 ( .A1(n17781), .A2(n17782), .ZN(n18174) );
  OR2_X1 U23377 ( .A1(n14845), .A2(n15284), .ZN(n14849) );
  XNOR2_X1 U23418 ( .A(n25014), .B(n25013), .ZN(n28650) );
  XNOR2_X1 U23428 ( .A(n25014), .B(n25013), .ZN(n28651) );
  NOR2_X1 U23433 ( .A1(n26356), .A2(n28650), .ZN(n28652) );
  XNOR2_X1 U23552 ( .A(n22604), .B(n22603), .ZN(n28653) );
  AOI21_X1 U23614 ( .B1(n24376), .B2(n23999), .A(n23998), .ZN(n28654) );
  XNOR2_X1 U23625 ( .A(n22604), .B(n22603), .ZN(n23809) );
  AOI21_X1 U23634 ( .B1(n24376), .B2(n23999), .A(n23998), .ZN(n25465) );
  OAI211_X1 U23651 ( .C1(n27192), .C2(n27193), .A(n4108), .B(n4110), .ZN(
        n28655) );
  OAI211_X1 U23669 ( .C1(n27192), .C2(n27193), .A(n4108), .B(n4110), .ZN(
        n27662) );
  BUF_X1 U23671 ( .A(n17872), .Z(n28656) );
  BUF_X1 U23703 ( .A(n20282), .Z(n28657) );
  XOR2_X1 U23736 ( .A(n18568), .B(n18567), .Z(n28658) );
  XNOR2_X1 U23838 ( .A(n21492), .B(n21491), .ZN(n28659) );
  XNOR2_X1 U23857 ( .A(n25699), .B(n25700), .ZN(n28660) );
  XNOR2_X1 U23922 ( .A(n19128), .B(n19127), .ZN(n20225) );
  NOR2_X1 U23977 ( .A1(n20583), .A2(n20582), .ZN(n28661) );
  NAND2_X1 U24006 ( .A1(n2372), .A2(n2371), .ZN(n28662) );
  AOI21_X1 U24054 ( .B1(n28663), .B2(n3771), .A(n5263), .ZN(n1008) );
  NAND2_X1 U24064 ( .A1(n26320), .A2(n26992), .ZN(n28663) );
  OAI21_X2 U24097 ( .B1(n8122), .B2(n8351), .A(n8121), .ZN(n10088) );
  OR2_X1 U24133 ( .A1(n20248), .A2(n20033), .ZN(n20641) );
  OAI21_X1 U24179 ( .B1(n15689), .B2(n28666), .A(n28665), .ZN(n15693) );
  NAND2_X1 U24213 ( .A1(n15689), .A2(n15690), .ZN(n28665) );
  NOR2_X1 U24219 ( .A1(n20044), .A2(n20158), .ZN(n19982) );
  NAND2_X1 U24220 ( .A1(n17762), .A2(n17942), .ZN(n17761) );
  NAND2_X1 U24408 ( .A1(n15388), .A2(n15144), .ZN(n15390) );
  NAND2_X1 U24475 ( .A1(n27107), .A2(n28667), .ZN(n27755) );
  NAND2_X1 U24547 ( .A1(n4794), .A2(n23370), .ZN(n2119) );
  XNOR2_X1 U24549 ( .A(n28668), .B(n3083), .ZN(Ciphertext[118]) );
  OAI21_X1 U24573 ( .B1(n27752), .B2(n27751), .A(n27750), .ZN(n28668) );
  OAI21_X1 U24698 ( .B1(n20362), .B2(n21520), .A(n21180), .ZN(n20363) );
  NOR2_X1 U24748 ( .A1(n8509), .A2(n8510), .ZN(n9431) );
  NAND2_X1 U24752 ( .A1(n28671), .A2(n17849), .ZN(n6444) );
  NAND2_X1 U24779 ( .A1(n2719), .A2(n17845), .ZN(n28671) );
  NAND3_X1 U24923 ( .A1(n11661), .A2(n2142), .A3(n12163), .ZN(n12104) );
  NAND2_X1 U24993 ( .A1(n12167), .A2(n11376), .ZN(n11381) );
  NAND2_X1 U24995 ( .A1(n5234), .A2(n18388), .ZN(n28672) );
  AND4_X2 U24998 ( .A1(n1556), .A2(n1555), .A3(n4994), .A4(n1558), .ZN(n24633)
         );
  NAND2_X1 U25074 ( .A1(n24460), .A2(n24808), .ZN(n24816) );
  INV_X1 U25166 ( .A(n5759), .ZN(n5245) );
  NAND2_X1 U25171 ( .A1(n5758), .A2(n5756), .ZN(n5759) );
  INV_X1 U25174 ( .A(n21634), .ZN(n21635) );
  NAND2_X1 U25283 ( .A1(n12149), .A2(n12991), .ZN(n28676) );
  NAND2_X1 U25328 ( .A1(n24811), .A2(n24810), .ZN(n28679) );
  NAND2_X1 U25348 ( .A1(n21013), .A2(n2639), .ZN(n22053) );
  NAND2_X1 U25376 ( .A1(n25966), .A2(n25965), .ZN(n28680) );
  NAND3_X1 U25377 ( .A1(n8630), .A2(n8627), .A3(n8664), .ZN(n8629) );
  NAND3_X1 U25397 ( .A1(n24372), .A2(n23994), .A3(n23995), .ZN(n28717) );
  NAND2_X1 U25423 ( .A1(n7968), .A2(n1938), .ZN(n7970) );
  NAND2_X1 U25432 ( .A1(n20948), .A2(n21499), .ZN(n20949) );
  OAI21_X1 U25434 ( .B1(n24073), .B2(n23372), .A(n28681), .ZN(n23374) );
  NAND2_X1 U25505 ( .A1(n3989), .A2(n11548), .ZN(n28682) );
  OAI211_X2 U25517 ( .C1(n14511), .C2(n14512), .A(n14509), .B(n28683), .ZN(
        n16023) );
  NAND2_X1 U25527 ( .A1(n14512), .A2(n15251), .ZN(n28683) );
  NAND3_X1 U25592 ( .A1(n12278), .A2(n11801), .A3(n12280), .ZN(n2288) );
  AOI21_X2 U25595 ( .B1(n8118), .B2(n8653), .A(n5819), .ZN(n10087) );
  NAND2_X1 U25615 ( .A1(n981), .A2(n28685), .ZN(n28684) );
  NOR2_X1 U25616 ( .A1(n14204), .A2(n28220), .ZN(n28685) );
  NAND3_X2 U25643 ( .A1(n28687), .A2(n23201), .A3(n28686), .ZN(n25775) );
  INV_X1 U25650 ( .A(n24561), .ZN(n28686) );
  NAND2_X1 U25674 ( .A1(n6046), .A2(n3881), .ZN(n6044) );
  OAI21_X1 U25682 ( .B1(n29547), .B2(n18410), .A(n28688), .ZN(n17820) );
  NAND2_X1 U25709 ( .A1(n18028), .A2(n18410), .ZN(n28688) );
  NAND2_X1 U25735 ( .A1(n7755), .A2(n887), .ZN(n28689) );
  NAND2_X1 U25781 ( .A1(n28690), .A2(n23751), .ZN(n2818) );
  NAND2_X1 U25851 ( .A1(n23747), .A2(n409), .ZN(n28690) );
  OAI21_X1 U25940 ( .B1(n28692), .B2(n7890), .A(n28691), .ZN(n7090) );
  NAND2_X1 U25952 ( .A1(n7315), .A2(n7890), .ZN(n28691) );
  NAND2_X1 U26013 ( .A1(n11114), .A2(n10490), .ZN(n10547) );
  NAND2_X1 U26023 ( .A1(n22971), .A2(n6728), .ZN(n4233) );
  NAND2_X1 U26029 ( .A1(n24712), .A2(n28524), .ZN(n24410) );
  NAND2_X1 U26054 ( .A1(n15362), .A2(n15363), .ZN(n15364) );
  NAND2_X1 U26139 ( .A1(n28694), .A2(n27417), .ZN(n27421) );
  NAND2_X1 U26304 ( .A1(n29529), .A2(n29542), .ZN(n28694) );
  NAND3_X1 U26371 ( .A1(n7293), .A2(n8156), .A3(n7781), .ZN(n28696) );
  INV_X1 U26424 ( .A(n19881), .ZN(n20604) );
  NAND2_X1 U26425 ( .A1(n20598), .A2(n4569), .ZN(n19881) );
  NAND2_X1 U26426 ( .A1(n14885), .A2(n14972), .ZN(n14582) );
  NAND2_X1 U26444 ( .A1(n14971), .A2(n14969), .ZN(n14885) );
  NAND2_X1 U26501 ( .A1(n390), .A2(n11751), .ZN(n28698) );
  NAND2_X1 U26502 ( .A1(n12219), .A2(n12218), .ZN(n12222) );
  OAI21_X1 U26630 ( .B1(n8718), .B2(n8717), .A(n28699), .ZN(n8442) );
  NAND2_X1 U26646 ( .A1(n8718), .A2(n8719), .ZN(n28699) );
  NAND2_X1 U26789 ( .A1(n28702), .A2(n10717), .ZN(n28701) );
  INV_X1 U26793 ( .A(n11793), .ZN(n28702) );
  NAND2_X1 U26837 ( .A1(n21698), .A2(n21696), .ZN(n21695) );
  NAND3_X1 U26844 ( .A1(n3016), .A2(n2019), .A3(n17754), .ZN(n21698) );
  NAND3_X2 U26851 ( .A1(n5543), .A2(n28704), .A3(n28703), .ZN(n13447) );
  NAND2_X1 U26895 ( .A1(n12083), .A2(n12289), .ZN(n28704) );
  NAND2_X1 U26898 ( .A1(n7591), .A2(n441), .ZN(n5483) );
  AND2_X1 U26915 ( .A1(n21503), .A2(n21539), .ZN(n20947) );
  NAND3_X1 U26952 ( .A1(n28706), .A2(n29552), .A3(n26151), .ZN(n26153) );
  NAND2_X1 U26954 ( .A1(n28710), .A2(n26789), .ZN(n28706) );
  NAND2_X1 U26984 ( .A1(n3459), .A2(n23779), .ZN(n28707) );
  OAI21_X1 U26993 ( .B1(n26792), .B2(n28709), .A(n28708), .ZN(n26795) );
  NAND2_X1 U27010 ( .A1(n26792), .A2(n26793), .ZN(n28708) );
  INV_X1 U27039 ( .A(n26791), .ZN(n28711) );
  NAND2_X1 U27045 ( .A1(n1764), .A2(n1763), .ZN(n28712) );
  NAND2_X1 U27065 ( .A1(n28714), .A2(n28713), .ZN(n26796) );
  NAND2_X1 U27131 ( .A1(n26790), .A2(n26791), .ZN(n28713) );
  NAND2_X1 U27170 ( .A1(n26924), .A2(n28711), .ZN(n28714) );
  NAND2_X1 U27191 ( .A1(n28715), .A2(n8176), .ZN(n2659) );
  NAND2_X1 U27201 ( .A1(n7763), .A2(n7347), .ZN(n28715) );
  AOI21_X1 U27226 ( .B1(n28716), .B2(n7313), .A(n7176), .ZN(n7112) );
  NAND2_X1 U27267 ( .A1(n7896), .A2(n7895), .ZN(n28716) );
  OAI21_X1 U27341 ( .B1(n1828), .B2(n23997), .A(n28717), .ZN(n23998) );
  NAND2_X1 U27346 ( .A1(n23819), .A2(n23820), .ZN(n23090) );
  NAND2_X1 U27376 ( .A1(n17316), .A2(n4220), .ZN(n16836) );
  AOI22_X1 U27377 ( .A1(n28718), .A2(n27382), .B1(n27037), .B2(n28378), .ZN(
        n27039) );
  NAND2_X1 U27382 ( .A1(n27212), .A2(n5312), .ZN(n28718) );
  XNOR2_X1 U27477 ( .A(n12861), .B(n3871), .ZN(n253) );
  NAND2_X1 U27480 ( .A1(n11569), .A2(n11568), .ZN(n28719) );
  NAND2_X1 U27511 ( .A1(n11570), .A2(n4341), .ZN(n28720) );
  NAND2_X1 U27528 ( .A1(n28721), .A2(n7822), .ZN(n7823) );
  NAND3_X1 U27562 ( .A1(n16804), .A2(n16802), .A3(n16801), .ZN(n17780) );
  NAND3_X1 U27576 ( .A1(n26), .A2(n11469), .A3(n11468), .ZN(n25) );
  NAND2_X1 U27616 ( .A1(n14104), .A2(n14103), .ZN(n28722) );
  NOR2_X1 U27620 ( .A1(n21484), .A2(n28723), .ZN(n19859) );
  NAND2_X1 U27625 ( .A1(n1528), .A2(n1529), .ZN(n1527) );
  NAND2_X1 U27628 ( .A1(n18111), .A2(n17902), .ZN(n17905) );
  NAND2_X1 U27654 ( .A1(n11965), .A2(n28726), .ZN(n28725) );
  NAND2_X1 U27698 ( .A1(n17487), .A2(n17076), .ZN(n17486) );
  OR2_X1 U27724 ( .A1(n14947), .A2(n6855), .ZN(n28727) );
  OR2_X1 U27766 ( .A1(n20577), .A2(n20580), .ZN(n5545) );
  NAND3_X1 U27851 ( .A1(n28730), .A2(n9244), .A3(n9410), .ZN(n9251) );
  NAND2_X1 U27861 ( .A1(n28211), .A2(n9243), .ZN(n28730) );
  NAND2_X1 U27862 ( .A1(n17804), .A2(n16898), .ZN(n28) );
  OR2_X1 U27876 ( .A1(n7266), .A2(n7265), .ZN(n8029) );
  NAND2_X1 U27881 ( .A1(n2170), .A2(n4129), .ZN(n7259) );
  NAND2_X1 U27903 ( .A1(n342), .A2(n26960), .ZN(n27390) );
  NAND2_X1 U27929 ( .A1(n28732), .A2(n2954), .ZN(n11058) );
  OAI21_X1 U27930 ( .B1(n11030), .B2(n11031), .A(n11283), .ZN(n28732) );
  NAND3_X1 U28002 ( .A1(n28404), .A2(n18349), .A3(n17646), .ZN(n28733) );
  INV_X1 U28003 ( .A(n13857), .ZN(n13856) );
  NAND2_X1 U28017 ( .A1(n13673), .A2(n13855), .ZN(n13857) );
  NAND2_X1 U28037 ( .A1(n28734), .A2(n6465), .ZN(n16667) );
  OAI21_X1 U28039 ( .B1(n17277), .B2(n17278), .A(n16844), .ZN(n28734) );
  NAND3_X2 U28121 ( .A1(n2645), .A2(n14700), .A3(n2642), .ZN(n16216) );
  NAND2_X1 U28126 ( .A1(n6097), .A2(n6098), .ZN(n23878) );
  OAI21_X1 U28127 ( .B1(n7964), .B2(n7963), .A(n28736), .ZN(n7578) );
  NAND2_X1 U28128 ( .A1(n7964), .A2(n7965), .ZN(n28736) );
  XNOR2_X1 U28129 ( .A(n22681), .B(n22903), .ZN(n22495) );
  OAI21_X1 U28130 ( .B1(n23817), .B2(n23818), .A(n28738), .ZN(n28737) );
  INV_X1 U28131 ( .A(n15617), .ZN(n15106) );
  NOR2_X1 U28133 ( .A1(n16965), .A2(n28739), .ZN(n16966) );
  AOI22_X2 U28135 ( .A1(n5407), .A2(n14780), .B1(n14683), .B2(n14684), .ZN(
        n15909) );
  NAND2_X1 U28138 ( .A1(n28741), .A2(n26946), .ZN(n27525) );
  AOI22_X1 U28139 ( .A1(n6948), .A2(n26944), .B1(n26942), .B2(n26943), .ZN(
        n28741) );
  NAND2_X1 U28140 ( .A1(n28744), .A2(n28742), .ZN(n9916) );
  NAND2_X1 U28141 ( .A1(n8442), .A2(n28743), .ZN(n28742) );
  NAND2_X1 U28142 ( .A1(n8441), .A2(n8440), .ZN(n28744) );
  INV_X1 U28143 ( .A(n18292), .ZN(n28745) );
  NOR2_X1 U28144 ( .A1(n1630), .A2(n567), .ZN(n2542) );
  OAI211_X2 U28145 ( .C1(n13781), .C2(n14254), .A(n13779), .B(n28746), .ZN(
        n15208) );
  NAND3_X1 U28146 ( .A1(n14253), .A2(n14254), .A3(n29312), .ZN(n28746) );
  NAND2_X1 U28147 ( .A1(n307), .A2(n27029), .ZN(n26819) );
  NAND3_X2 U28148 ( .A1(n14726), .A2(n3605), .A3(n14727), .ZN(n16280) );
  NAND3_X1 U28149 ( .A1(n6678), .A2(n6680), .A3(n28747), .ZN(n12589) );
  NAND2_X1 U28150 ( .A1(n28748), .A2(n5889), .ZN(n3781) );
  NAND2_X1 U28151 ( .A1(n9025), .A2(n9024), .ZN(n28748) );
  NAND2_X1 U28152 ( .A1(n697), .A2(n18322), .ZN(n17714) );
  NAND2_X1 U28155 ( .A1(n20535), .A2(n20934), .ZN(n28749) );
  NAND2_X1 U28156 ( .A1(n20534), .A2(n21078), .ZN(n28750) );
  NAND2_X1 U28157 ( .A1(n2697), .A2(n405), .ZN(n4686) );
  INV_X1 U28158 ( .A(n28752), .ZN(n28751) );
  OAI21_X1 U28159 ( .B1(n7423), .B2(n370), .A(n7422), .ZN(n28752) );
  NAND2_X1 U28162 ( .A1(n28121), .A2(n58), .ZN(n28753) );
  OR2_X1 U28163 ( .A1(n13898), .A2(n58), .ZN(n28754) );
  NAND3_X2 U28165 ( .A1(n1463), .A2(n1468), .A3(n17448), .ZN(n18942) );
  OAI211_X1 U28167 ( .C1(n28015), .C2(n28411), .A(n26984), .B(n28018), .ZN(
        n25990) );
  NAND3_X1 U28168 ( .A1(n1802), .A2(n1800), .A3(n1801), .ZN(n1798) );
  NAND3_X1 U28170 ( .A1(n17803), .A2(n3994), .A3(n18277), .ZN(n27) );
  NAND2_X1 U28171 ( .A1(n416), .A2(n19946), .ZN(n3809) );
  NAND2_X1 U28172 ( .A1(n17106), .A2(n17470), .ZN(n17515) );
  XNOR2_X2 U28174 ( .A(n12086), .B(n12085), .ZN(n14484) );
  NAND2_X1 U28175 ( .A1(n26315), .A2(n28214), .ZN(n26316) );
  NAND3_X1 U28178 ( .A1(n7464), .A2(n7618), .A3(n7463), .ZN(n7469) );
  NAND2_X1 U28179 ( .A1(n8246), .A2(n7690), .ZN(n3510) );
  NAND2_X1 U28181 ( .A1(n3658), .A2(n698), .ZN(n22835) );
  NAND2_X1 U28182 ( .A1(n4048), .A2(n4050), .ZN(n15047) );
  NAND2_X1 U28183 ( .A1(n693), .A2(n695), .ZN(n15341) );
  NAND2_X1 U28184 ( .A1(n18500), .A2(n520), .ZN(n4707) );
  NAND2_X1 U28185 ( .A1(n12079), .A2(n12058), .ZN(n5543) );
  OAI22_X1 U28186 ( .A1(n12291), .A2(n12080), .B1(n29324), .B2(n11795), .ZN(
        n12079) );
  NAND3_X1 U28188 ( .A1(n15205), .A2(n15203), .A3(n15204), .ZN(n28756) );
  NAND3_X1 U28191 ( .A1(n28757), .A2(n217), .A3(n15509), .ZN(n4708) );
  NAND2_X1 U28192 ( .A1(n2347), .A2(n15515), .ZN(n28757) );
  NAND3_X1 U28194 ( .A1(n18509), .A2(n510), .A3(n18510), .ZN(n6255) );
  NAND3_X1 U28195 ( .A1(n28759), .A2(n3690), .A3(n2463), .ZN(n1688) );
  OAI21_X1 U28196 ( .B1(n1691), .B2(n1690), .A(n28107), .ZN(n28759) );
  OR3_X1 U28198 ( .A1(n16992), .A2(n29299), .A3(n17263), .ZN(n16771) );
  NAND2_X1 U28200 ( .A1(n4892), .A2(n4872), .ZN(n4871) );
  OAI22_X1 U28201 ( .A1(n27113), .A2(n401), .B1(n26865), .B2(n27112), .ZN(
        n27114) );
  OAI211_X2 U28202 ( .C1(n8738), .C2(n8739), .A(n8737), .B(n8736), .ZN(n9931)
         );
  AND2_X1 U28203 ( .A1(n1876), .A2(n14432), .ZN(n28761) );
  AND2_X1 U28204 ( .A1(n15374), .A2(n14863), .ZN(n28762) );
  NAND2_X1 U28206 ( .A1(n18506), .A2(n18213), .ZN(n28763) );
  CLKBUF_X1 U28207 ( .A(n20425), .Z(n22012) );
  OAI211_X2 U28208 ( .C1(n5826), .C2(n6914), .A(n19828), .B(n1972), .ZN(n21496) );
  OR2_X1 U28209 ( .A1(n23194), .A2(n23647), .ZN(n28764) );
  NAND2_X2 U28210 ( .A1(n5309), .A2(n1162), .ZN(n6348) );
  OR2_X1 U28212 ( .A1(n23183), .A2(n23641), .ZN(n28765) );
  OR2_X2 U28215 ( .A1(n26190), .A2(n26189), .ZN(n27038) );
  OR2_X2 U1524 ( .A1(n28308), .A2(n17893), .ZN(n18691) );
  XNOR2_X2 U627 ( .A(n22917), .B(n22916), .ZN(n23460) );
  XNOR2_X2 U2310 ( .A(n10155), .B(n10154), .ZN(n11086) );
  MUX2_X2 U932 ( .A(n8660), .B(n8659), .S(n8658), .Z(n9915) );
  AND2_X2 U1752 ( .A1(n669), .A2(n670), .ZN(n19331) );
  AND2_X2 U1204 ( .A1(n5791), .A2(n5792), .ZN(n18471) );
  OAI21_X2 U12394 ( .B1(n22939), .B2(n23449), .A(n22938), .ZN(n24591) );
  AND2_X2 U4286 ( .A1(n1189), .A2(n1188), .ZN(n21657) );
  OAI21_X2 U5085 ( .B1(n23111), .B2(n29295), .A(n1498), .ZN(n24479) );
  NAND2_X2 U9238 ( .A1(n3850), .A2(n14208), .ZN(n15334) );
  XNOR2_X2 U18658 ( .A(n13188), .B(n13187), .ZN(n14031) );
  OR2_X2 U11500 ( .A1(n17817), .A2(n17816), .ZN(n19500) );
  AND2_X2 U1453 ( .A1(n9865), .A2(n12194), .ZN(n2483) );
  NAND2_X2 U2217 ( .A1(n11693), .A2(n11694), .ZN(n12219) );
  MUX2_X2 U1269 ( .A(n8435), .B(n8434), .S(n9034), .Z(n10295) );
  AND3_X2 U2252 ( .A1(n6373), .A2(n10112), .A3(n10111), .ZN(n10863) );
  BUF_X1 U19384 ( .A(n25293), .Z(n28576) );
  XNOR2_X2 U3435 ( .A(n7140), .B(Key[49]), .ZN(n7743) );
  BUF_X2 U907 ( .A(n12166), .Z(n1931) );
  AND2_X2 U8002 ( .A1(n20095), .A2(n20094), .ZN(n21078) );
  BUF_X1 U2344 ( .A(n23599), .Z(n24973) );
  MUX2_X2 U930 ( .A(n8070), .B(n8069), .S(n8501), .Z(n10219) );
  OR2_X2 U9983 ( .A1(n6516), .A2(n6514), .ZN(n12233) );
  NAND2_X2 U231 ( .A1(n3574), .A2(n3577), .ZN(n16416) );
  XNOR2_X2 U22399 ( .A(n19266), .B(n19265), .ZN(n19271) );
  AND2_X2 U292 ( .A1(n6103), .A2(n6101), .ZN(n19584) );
  OR2_X2 U10925 ( .A1(n8728), .A2(n8727), .ZN(n10264) );
  BUF_X1 U3427 ( .A(n7377), .Z(n7818) );
  OAI211_X2 U17446 ( .C1(n12334), .C2(n12327), .A(n11452), .B(n11451), .ZN(
        n13278) );
  OR2_X1 U1237 ( .A1(n6034), .A2(n23167), .ZN(n23681) );
  BUF_X1 U754 ( .A(n19556), .Z(n28143) );
  BUF_X1 U1199 ( .A(n27718), .Z(n324) );
  OR2_X2 U685 ( .A1(n21437), .A2(n5274), .ZN(n20833) );
  INV_X2 U3463 ( .A(n18469), .ZN(n6079) );
  MUX2_X2 U60 ( .A(n16228), .B(n16227), .S(n17138), .Z(n18469) );
  NAND3_X2 U4047 ( .A1(n4127), .A2(n1525), .A3(n4128), .ZN(n11867) );
  OAI211_X2 U3087 ( .C1(n11883), .C2(n11882), .A(n2349), .B(n2348), .ZN(n13478) );
  OAI211_X2 U15571 ( .C1(n22404), .C2(n21018), .A(n1720), .B(n21017), .ZN(
        n22735) );
  NAND4_X2 U5769 ( .A1(n7683), .A2(n7682), .A3(n7680), .A4(n7681), .ZN(n10322)
         );
  AND3_X2 U1110 ( .A1(n20884), .A2(n20883), .A3(n20882), .ZN(n21994) );
  MUX2_X2 U1933 ( .A(n16493), .B(n16492), .S(n18464), .Z(n18912) );
  MUX2_X2 U9665 ( .A(n9091), .B(n9090), .S(n2320), .Z(n10344) );
  OAI211_X2 U1894 ( .C1(n15288), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        n16017) );
  OAI21_X2 U3359 ( .B1(n7677), .B2(n7678), .A(n6540), .ZN(n9434) );
  OAI211_X2 U12642 ( .C1(n21138), .C2(n21605), .A(n21604), .B(n5719), .ZN(
        n22500) );
  AOI22_X1 U13340 ( .A1(n24580), .A2(n24581), .B1(n6056), .B2(n24467), .ZN(
        n6055) );
  XNOR2_X1 U12485 ( .A(n23125), .B(n23124), .ZN(n26789) );
  OAI21_X1 U5199 ( .B1(n1596), .B2(n16951), .A(n16950), .ZN(n18538) );
  AOI22_X1 U5477 ( .A1(n20271), .A2(n20270), .B1(n20269), .B2(n21665), .ZN(
        n1810) );
  MUX2_X2 U2671 ( .A(n17821), .B(n17820), .S(n18418), .Z(n19706) );
  OAI21_X1 U1294 ( .B1(n24297), .B2(n24894), .A(n24296), .ZN(n24298) );
  MUX2_X2 U6738 ( .A(n3863), .B(n10463), .S(n11137), .Z(n10766) );
  AOI22_X1 U4670 ( .A1(n21021), .A2(n22023), .B1(n21053), .B2(n22026), .ZN(
        n21917) );
  AND3_X2 U23577 ( .A1(n21176), .A2(n21175), .A3(n21174), .ZN(n22678) );
  XNOR2_X1 U8743 ( .A(n9276), .B(n9275), .ZN(n10703) );
  MUX2_X2 U1214 ( .A(n12046), .B(n12045), .S(n12219), .Z(n13525) );
  AND2_X2 U4815 ( .A1(n4153), .A2(n1282), .ZN(n25322) );
  BUF_X1 U3948 ( .A(n26125), .Z(n27147) );
  NAND4_X2 U2559 ( .A1(n20030), .A2(n20029), .A3(n4933), .A4(n4567), .ZN(
        n21392) );
  AND4_X2 U2918 ( .A1(n2068), .A2(n5848), .A3(n5886), .A4(n5845), .ZN(n14810)
         );
  OAI21_X1 U22015 ( .B1(n21220), .B2(n21215), .A(n18786), .ZN(n18787) );
  NAND2_X1 U232 ( .A1(n3030), .A2(n7247), .ZN(n8941) );
  XNOR2_X1 U5741 ( .A(n22213), .B(n21905), .ZN(n23790) );
  XNOR2_X1 U20810 ( .A(n4453), .B(n4452), .ZN(n17271) );
  MUX2_X2 U164 ( .A(n21944), .B(n21943), .S(n24729), .Z(n26038) );
  XNOR2_X1 U1957 ( .A(n3938), .B(n3937), .ZN(n16879) );
  OAI21_X2 U563 ( .B1(n23207), .B2(n24550), .A(n23206), .ZN(n25565) );
  BUF_X1 U1635 ( .A(n27718), .Z(n325) );
  XNOR2_X2 U2842 ( .A(n16466), .B(n16465), .ZN(n17506) );
  INV_X1 U23512 ( .A(n23686), .ZN(n23516) );
  NAND2_X2 U2668 ( .A1(n18112), .A2(n3074), .ZN(n19700) );
  MUX2_X1 U279 ( .A(n19926), .B(n19925), .S(n5935), .Z(n21748) );
  CLKBUF_X1 U2125 ( .A(Key[150]), .Z(n3673) );
  CLKBUF_X1 U1597 ( .A(Key[112]), .Z(n2916) );
  CLKBUF_X1 U1589 ( .A(Key[4]), .Z(n3598) );
  CLKBUF_X1 U1817 ( .A(Key[105]), .Z(n3081) );
  CLKBUF_X1 U2127 ( .A(Key[29]), .Z(n3483) );
  CLKBUF_X1 U76 ( .A(Key[116]), .Z(n3654) );
  CLKBUF_X1 U1826 ( .A(Key[47]), .Z(n3695) );
  XNOR2_X1 U14714 ( .A(n7139), .B(Key[52]), .ZN(n7533) );
  BUF_X1 U6646 ( .A(n7191), .Z(n7642) );
  NAND3_X1 U512 ( .A1(n7918), .A2(n2569), .A3(n2568), .ZN(n9116) );
  OAI211_X1 U9155 ( .C1(n8039), .C2(n8038), .A(n8037), .B(n2841), .ZN(n9123)
         );
  AND2_X1 U3349 ( .A1(n7567), .A2(n7566), .ZN(n9064) );
  AND2_X1 U192 ( .A1(n7277), .A2(n7276), .ZN(n8886) );
  INV_X1 U902 ( .A(n9245), .ZN(n9410) );
  NAND3_X1 U3367 ( .A1(n3034), .A2(n7602), .A3(n7603), .ZN(n8787) );
  OAI211_X1 U302 ( .C1(n7297), .C2(n8159), .A(n7158), .B(n7296), .ZN(n9243) );
  NAND2_X1 U371 ( .A1(n1033), .A2(n1032), .ZN(n8977) );
  NAND2_X1 U4523 ( .A1(n1139), .A2(n5989), .ZN(n8873) );
  INV_X1 U249 ( .A(n8635), .ZN(n8653) );
  INV_X1 U15171 ( .A(n7679), .ZN(n9438) );
  INV_X1 U2030 ( .A(n8735), .ZN(n8731) );
  AND2_X1 U768 ( .A1(n7066), .A2(n7065), .ZN(n2238) );
  AOI21_X1 U201 ( .B1(n7860), .B2(n7859), .A(n1614), .ZN(n10353) );
  AND3_X1 U3283 ( .A1(n9251), .A2(n9250), .A3(n9249), .ZN(n9785) );
  OAI21_X1 U3284 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(n10391) );
  AND3_X1 U3286 ( .A1(n3718), .A2(n4932), .A3(n1047), .ZN(n9446) );
  OAI21_X1 U4464 ( .B1(n9174), .B2(n8963), .A(n8470), .ZN(n10263) );
  NAND2_X1 U1317 ( .A1(n3101), .A2(n240), .ZN(n10202) );
  MUX2_X1 U8678 ( .A(n8668), .B(n8667), .S(n8666), .Z(n10133) );
  OR2_X1 U3260 ( .A1(n8633), .A2(n8632), .ZN(n9986) );
  OR2_X1 U5590 ( .A1(n8374), .A2(n8373), .ZN(n1895) );
  NAND2_X1 U9241 ( .A1(n8815), .A2(n2899), .ZN(n9852) );
  XNOR2_X1 U3247 ( .A(n748), .B(n10064), .ZN(n10332) );
  NAND2_X1 U3252 ( .A1(n8571), .A2(n9378), .ZN(n10311) );
  XNOR2_X1 U11328 ( .A(n10341), .B(n10340), .ZN(n11282) );
  XNOR2_X1 U16033 ( .A(n9263), .B(n9264), .ZN(n10592) );
  XNOR2_X1 U11514 ( .A(n9394), .B(n9395), .ZN(n28405) );
  CLKBUF_X1 U3211 ( .A(n9608), .Z(n10476) );
  BUF_X2 U683 ( .A(n10522), .Z(n10523) );
  OR2_X1 U14235 ( .A1(n11127), .A2(n11123), .ZN(n10760) );
  OR2_X1 U8939 ( .A1(n28204), .A2(n11045), .ZN(n11262) );
  AND2_X1 U311 ( .A1(n4405), .A2(n11494), .ZN(n12307) );
  NAND2_X1 U3131 ( .A1(n11658), .A2(n11657), .ZN(n12162) );
  NAND2_X1 U2239 ( .A1(n6248), .A2(n10100), .ZN(n3653) );
  NAND2_X1 U10478 ( .A1(n10584), .A2(n3533), .ZN(n12354) );
  OR2_X1 U8188 ( .A1(n11279), .A2(n11278), .ZN(n11795) );
  INV_X1 U17369 ( .A(n11801), .ZN(n12286) );
  OR3_X1 U5650 ( .A1(n4844), .A2(n12200), .A3(n12202), .ZN(n5524) );
  CLKBUF_X1 U1454 ( .A(n12286), .Z(n12401) );
  OAI22_X1 U3089 ( .A1(n5079), .A2(n11673), .B1(n11848), .B2(n11672), .ZN(
        n11846) );
  NAND2_X1 U234 ( .A1(n11936), .A2(n11935), .ZN(n13265) );
  OR2_X1 U3102 ( .A1(n1493), .A2(n11550), .ZN(n11160) );
  OAI211_X1 U79 ( .C1(n11518), .C2(n11674), .A(n11517), .B(n11516), .ZN(n12780) );
  AND2_X1 U1990 ( .A1(n2355), .A2(n4711), .ZN(n6645) );
  OAI21_X1 U1410 ( .B1(n11846), .B2(n11679), .A(n11678), .ZN(n13553) );
  AND2_X1 U256 ( .A1(n11504), .A2(n11503), .ZN(n12722) );
  XNOR2_X1 U2081 ( .A(n13123), .B(n13124), .ZN(n14131) );
  XNOR2_X1 U1985 ( .A(n13135), .B(n3097), .ZN(n14325) );
  XNOR2_X1 U417 ( .A(n13399), .B(n2875), .ZN(n2974) );
  XNOR2_X1 U18094 ( .A(n12494), .B(n12493), .ZN(n14429) );
  NAND3_X1 U18469 ( .A1(n28625), .A2(n14286), .A3(n14281), .ZN(n12936) );
  XNOR2_X1 U18167 ( .A(n12565), .B(n12564), .ZN(n14318) );
  OR2_X1 U2980 ( .A1(n14350), .A2(n13825), .ZN(n1748) );
  OR2_X1 U1980 ( .A1(n14240), .A2(n563), .ZN(n14244) );
  OR2_X1 U10034 ( .A1(n14244), .A2(n15199), .ZN(n14245) );
  OAI21_X1 U819 ( .B1(n4122), .B2(n4121), .A(n13125), .ZN(n15073) );
  AOI21_X1 U372 ( .B1(n14067), .B2(n14328), .A(n14066), .ZN(n15285) );
  OAI211_X1 U19343 ( .C1(n14386), .C2(n14385), .A(n14384), .B(n14383), .ZN(
        n15275) );
  CLKBUF_X1 U14236 ( .A(n14806), .Z(n28493) );
  NAND3_X1 U420 ( .A1(n645), .A2(n643), .A3(n642), .ZN(n15438) );
  OR2_X1 U6879 ( .A1(n5635), .A2(n15456), .ZN(n14797) );
  BUF_X1 U4646 ( .A(n13979), .Z(n14740) );
  NAND2_X1 U2921 ( .A1(n974), .A2(n973), .ZN(n15185) );
  MUX2_X1 U10271 ( .A(n14988), .B(n14987), .S(n15155), .Z(n16519) );
  OAI211_X1 U1639 ( .C1(n14559), .C2(n14558), .A(n14557), .B(n14556), .ZN(
        n16618) );
  AND2_X1 U686 ( .A1(n6673), .A2(n6672), .ZN(n16467) );
  OR2_X1 U2872 ( .A1(n13984), .A2(n13983), .ZN(n15788) );
  OAI21_X1 U19692 ( .B1(n1809), .B2(n14958), .A(n14957), .ZN(n16296) );
  NAND3_X1 U6796 ( .A1(n150), .A2(n14758), .A3(n14759), .ZN(n16578) );
  INV_X1 U2866 ( .A(n15618), .ZN(n16400) );
  NAND3_X1 U214 ( .A1(n5), .A2(n14867), .A3(n2), .ZN(n16456) );
  NOR2_X1 U11559 ( .A1(n5596), .A2(n15172), .ZN(n16264) );
  XNOR2_X1 U5849 ( .A(n15838), .B(n15837), .ZN(n17556) );
  XNOR2_X1 U4538 ( .A(n16158), .B(n16157), .ZN(n17464) );
  XNOR2_X1 U1053 ( .A(n4588), .B(n16055), .ZN(n17283) );
  BUF_X1 U20127 ( .A(n16943), .Z(n17549) );
  INV_X1 U2814 ( .A(n17433), .ZN(n17440) );
  XNOR2_X1 U965 ( .A(n15258), .B(n15257), .ZN(n6002) );
  BUF_X1 U2783 ( .A(n16883), .Z(n17527) );
  OR2_X1 U328 ( .A1(n17432), .A2(n17431), .ZN(n31) );
  OR2_X1 U6976 ( .A1(n17781), .A2(n17782), .ZN(n4044) );
  AND2_X1 U1267 ( .A1(n16966), .A2(n6224), .ZN(n17858) );
  NOR2_X1 U20249 ( .A1(n18063), .A2(n18064), .ZN(n15939) );
  OR2_X1 U6428 ( .A1(n18186), .A2(n527), .ZN(n2135) );
  OR2_X1 U2685 ( .A1(n757), .A2(n18343), .ZN(n4077) );
  OAI211_X1 U8519 ( .C1(n17676), .C2(n18487), .A(n17675), .B(n2459), .ZN(n3444) );
  OAI211_X1 U2680 ( .C1(n4943), .C2(n5223), .A(n3349), .B(n3350), .ZN(n16990)
         );
  NOR2_X1 U731 ( .A1(n18714), .A2(n18713), .ZN(n19075) );
  AND2_X1 U524 ( .A1(n17723), .A2(n17722), .ZN(n19656) );
  NAND3_X1 U2659 ( .A1(n18436), .A2(n18435), .A3(n18434), .ZN(n19207) );
  XNOR2_X1 U2629 ( .A(n5523), .B(n5520), .ZN(n20295) );
  XNOR2_X1 U2630 ( .A(n18775), .B(n6667), .ZN(n19761) );
  XNOR2_X1 U22372 ( .A(n19223), .B(n19224), .ZN(n20342) );
  XNOR2_X1 U21923 ( .A(n18673), .B(n18674), .ZN(n20374) );
  XNOR2_X1 U2614 ( .A(n5224), .B(n17171), .ZN(n20404) );
  XNOR2_X1 U691 ( .A(n18694), .B(n18693), .ZN(n20373) );
  OR2_X1 U6105 ( .A1(n4245), .A2(n19928), .ZN(n20645) );
  OR2_X1 U7077 ( .A1(n20645), .A2(n5783), .ZN(n5781) );
  NAND3_X1 U2533 ( .A1(n20257), .A2(n20256), .A3(n1564), .ZN(n21429) );
  INV_X1 U2543 ( .A(n20966), .ZN(n21217) );
  OAI21_X1 U22855 ( .B1(n19942), .B2(n19955), .A(n19941), .ZN(n21400) );
  INV_X1 U23260 ( .A(n21343), .ZN(n21242) );
  BUF_X1 U2506 ( .A(n21014), .Z(n22402) );
  NAND2_X1 U1904 ( .A1(n20058), .A2(n20057), .ZN(n21213) );
  OR2_X1 U2514 ( .A1(n19893), .A2(n19894), .ZN(n21567) );
  AND3_X1 U2481 ( .A1(n6733), .A2(n20768), .A3(n6731), .ZN(n22240) );
  XNOR2_X1 U24385 ( .A(n22327), .B(n22328), .ZN(n22651) );
  XNOR2_X1 U24216 ( .A(n22118), .B(n22117), .ZN(n22121) );
  BUF_X1 U2424 ( .A(n23102), .Z(n23431) );
  XNOR2_X1 U227 ( .A(n22484), .B(n22483), .ZN(n28460) );
  XNOR2_X1 U5614 ( .A(n21873), .B(n21874), .ZN(n1914) );
  XNOR2_X1 U1895 ( .A(n21057), .B(n21056), .ZN(n23679) );
  BUF_X1 U161 ( .A(n23213), .Z(n23403) );
  XNOR2_X1 U488 ( .A(n21928), .B(n21927), .ZN(n23799) );
  OAI21_X1 U22929 ( .B1(n28390), .B2(n2138), .A(n23313), .ZN(n23565) );
  AND2_X1 U1678 ( .A1(n23264), .A2(n23265), .ZN(n25005) );
  MUX2_X1 U24827 ( .A(n23007), .B(n23524), .S(n23663), .Z(n23009) );
  NAND2_X1 U11924 ( .A1(n23264), .A2(n23265), .ZN(n28415) );
  NOR2_X1 U25233 ( .A1(n23782), .A2(n23781), .ZN(n24801) );
  OAI21_X1 U168 ( .B1(n23232), .B2(n1862), .A(n23231), .ZN(n24651) );
  OAI211_X1 U1555 ( .C1(n23695), .C2(n5482), .A(n5481), .B(n5480), .ZN(n24809)
         );
  NOR2_X1 U4283 ( .A1(n22948), .A2(n22947), .ZN(n24542) );
  INV_X1 U174 ( .A(n24378), .ZN(n1828) );
  MUX2_X1 U12517 ( .A(n23133), .B(n23132), .S(n23678), .Z(n24532) );
  AND2_X2 U12955 ( .A1(n24544), .A2(n2054), .ZN(n24547) );
  OAI211_X1 U25549 ( .C1(n24237), .C2(n24236), .A(n24235), .B(n24234), .ZN(
        n25745) );
  MUX2_X1 U437 ( .A(n24156), .B(n24649), .S(n3061), .Z(n25261) );
  AOI21_X1 U1544 ( .B1(n23027), .B2(n24310), .A(n23026), .ZN(n25910) );
  NAND2_X1 U4492 ( .A1(n24080), .A2(n1128), .ZN(n25251) );
  BUF_X1 U438 ( .A(n25844), .Z(n363) );
  OAI21_X1 U22309 ( .B1(n1777), .B2(n1828), .A(n23094), .ZN(n28628) );
  NAND3_X1 U5081 ( .A1(n1495), .A2(n1653), .A3(n1652), .ZN(n25262) );
  XNOR2_X1 U25089 ( .A(n23414), .B(n23413), .ZN(n26793) );
  XNOR2_X1 U2266 ( .A(n25078), .B(n25077), .ZN(n26920) );
  XNOR2_X1 U15484 ( .A(n25765), .B(n25766), .ZN(n26989) );
  INV_X1 U7456 ( .A(n26911), .ZN(n5625) );
  AND2_X1 U6338 ( .A1(n3589), .A2(n3590), .ZN(n27819) );
  OR2_X1 U2193 ( .A1(n27725), .A2(n27724), .ZN(n26889) );
  AND2_X1 U2206 ( .A1(n1944), .A2(n5373), .ZN(n27382) );
  BUF_X1 U22972 ( .A(n27997), .Z(n28636) );
  CLKBUF_X1 U12488 ( .A(n27913), .Z(n1843) );
  CLKBUF_X1 U2097 ( .A(Key[30]), .Z(n3423) );
  CLKBUF_X1 U1603 ( .A(Key[144]), .Z(n28327) );
  NAND2_X1 U11983 ( .A1(n10687), .A2(n10963), .ZN(n10966) );
  OR2_X1 U3138 ( .A1(n10168), .A2(n10167), .ZN(n12125) );
  OR2_X1 U1558 ( .A1(n11877), .A2(n10868), .ZN(n1630) );
  NAND2_X1 U1455 ( .A1(n6645), .A2(n11361), .ZN(n6647) );
  CLKBUF_X1 U13059 ( .A(n17541), .Z(n28454) );
  INV_X1 U11129 ( .A(n17478), .ZN(n3883) );
  INV_X1 U20340 ( .A(n16904), .ZN(n17710) );
  OAI21_X1 U21390 ( .B1(n17736), .B2(n17735), .A(n17734), .ZN(n17965) );
  INV_X1 U2608 ( .A(n20324), .ZN(n502) );
  OR2_X1 U2588 ( .A1(n20020), .A2(n19795), .ZN(n19796) );
  AOI21_X1 U1508 ( .B1(n3973), .B2(n3974), .A(n20586), .ZN(n21134) );
  NAND2_X2 U8285 ( .A1(n21611), .A2(n21610), .ZN(n21326) );
  INV_X1 U2353 ( .A(n24367), .ZN(n23897) );
  NOR2_X1 U10287 ( .A1(n24650), .A2(n24155), .ZN(n24524) );
  BUF_X1 U5925 ( .A(n26850), .Z(n26849) );
  NOR2_X1 U4002 ( .A1(n27898), .A2(n26510), .ZN(n27904) );
  NOR2_X1 U143 ( .A1(n28403), .A2(n27818), .ZN(n27812) );
  NOR2_X1 U26338 ( .A1(n27433), .A2(n27439), .ZN(n27432) );
  AND3_X2 U870 ( .A1(n2626), .A2(n2625), .A3(n2629), .ZN(n8504) );
  OR2_X2 U27190 ( .A1(n5640), .A2(n5643), .ZN(n16498) );
  AND3_X2 U453 ( .A1(n782), .A2(n778), .A3(n781), .ZN(n18242) );
  OR2_X2 U8286 ( .A1(n7409), .A2(n2491), .ZN(n9133) );
  NAND2_X2 U8399 ( .A1(n2772), .A2(n7894), .ZN(n8658) );
  BUF_X2 U1400 ( .A(n17474), .Z(n16725) );
  AND2_X2 U21643 ( .A1(n18207), .A2(n18208), .ZN(n19491) );
  BUF_X1 U4311 ( .A(n19855), .Z(n20552) );
  BUF_X2 U3012 ( .A(n13744), .Z(n14254) );
  OAI211_X2 U409 ( .C1(n13769), .C2(n15199), .A(n13741), .B(n13740), .ZN(
        n15379) );
  AND2_X2 U11685 ( .A1(n4390), .A2(n10744), .ZN(n11671) );
  OAI21_X2 U3282 ( .B1(n9002), .B2(n9200), .A(n4302), .ZN(n10426) );
  NAND4_X2 U1160 ( .A1(n7735), .A2(n7031), .A3(n7032), .A4(n3115), .ZN(n8874)
         );
  AND2_X2 U5074 ( .A1(n1490), .A2(n1489), .ZN(n13380) );
  OAI211_X2 U9006 ( .C1(n21544), .C2(n21543), .A(n2725), .B(n2724), .ZN(n21980) );
  AND4_X2 U45 ( .A1(n2857), .A2(n2856), .A3(n17507), .A4(n2858), .ZN(n520) );
  AOI21_X2 U1252 ( .B1(n8791), .B2(n8787), .A(n8723), .ZN(n9877) );
  BUF_X2 U1084 ( .A(n23867), .Z(n24716) );
  BUF_X2 U1520 ( .A(n11037), .Z(n279) );
  OAI211_X2 U1063 ( .C1(n12162), .C2(n10897), .A(n10896), .B(n11843), .ZN(
        n13556) );
  OR2_X2 U25717 ( .A1(n28689), .A2(n7757), .ZN(n10022) );
  OR2_X2 U5069 ( .A1(n19884), .A2(n19885), .ZN(n4193) );
  AND3_X2 U466 ( .A1(n1307), .A2(n1306), .A3(n2234), .ZN(n18017) );
  NAND3_X2 U8411 ( .A1(n11342), .A2(n11343), .A3(n2580), .ZN(n12281) );
  XNOR2_X2 U1615 ( .A(n18004), .B(n18005), .ZN(n20200) );
  AND2_X2 U24300 ( .A1(n22217), .A2(n22216), .ZN(n24735) );
  BUF_X2 U17451 ( .A(n13017), .Z(n12894) );
  NAND2_X2 U1125 ( .A1(n17874), .A2(n1034), .ZN(n19643) );
  AND2_X2 U4436 ( .A1(n1102), .A2(n1101), .ZN(n13260) );
  OAI211_X2 U3278 ( .C1(n9105), .C2(n9104), .A(n4969), .B(n9121), .ZN(n4714)
         );
  NOR2_X1 U112 ( .A1(n3127), .A2(n3128), .ZN(n9430) );
  AND2_X2 U10250 ( .A1(n3392), .A2(n3391), .ZN(n24383) );
  AND4_X2 U5852 ( .A1(n17189), .A2(n4168), .A3(n4480), .A4(n4241), .ZN(n18410)
         );
  XNOR2_X2 U9677 ( .A(n18363), .B(n18362), .ZN(n20546) );
  BUF_X2 U7358 ( .A(n7192), .Z(n7985) );
  AND2_X2 U10892 ( .A1(n6076), .A2(n6078), .ZN(n19225) );
  NOR2_X2 U3879 ( .A1(n5626), .A2(n5627), .ZN(n2209) );
  XNOR2_X2 U1989 ( .A(n13409), .B(n13408), .ZN(n1368) );
  XNOR2_X2 U9136 ( .A(n13605), .B(n13604), .ZN(n17425) );
  OR2_X2 U14976 ( .A1(n7392), .A2(n7391), .ZN(n9132) );
  AND2_X2 U1278 ( .A1(n2947), .A2(n10109), .ZN(n11990) );
  NAND3_X2 U912 ( .A1(n15442), .A2(n5681), .A3(n15443), .ZN(n16303) );
  NOR2_X2 U1301 ( .A1(n27900), .A2(n27899), .ZN(n27919) );
  OAI21_X2 U1043 ( .B1(n7961), .B2(n7960), .A(n3368), .ZN(n8666) );
  OAI211_X2 U9858 ( .C1(n8496), .C2(n8495), .A(n8494), .B(n8493), .ZN(n9771)
         );
  BUF_X2 U571 ( .A(n7040), .Z(n7982) );
  NAND3_X2 U4367 ( .A1(n1107), .A2(n11916), .A3(n11917), .ZN(n13482) );
  AND2_X2 U14504 ( .A1(n7014), .A2(n7013), .ZN(n8881) );
  AOI21_X2 U7409 ( .B1(n16754), .B2(n16753), .A(n16752), .ZN(n18179) );
  AND3_X2 U564 ( .A1(n2162), .A2(n2073), .A3(n2160), .ZN(n15780) );
  NAND3_X2 U3268 ( .A1(n8190), .A2(n8189), .A3(n8188), .ZN(n9295) );
  XNOR2_X2 U3462 ( .A(Key[116]), .B(Plaintext[116]), .ZN(n7935) );
  NAND3_X2 U897 ( .A1(n1020), .A2(n13304), .A3(n13303), .ZN(n15690) );
  OAI21_X2 U10092 ( .B1(n19746), .B2(n4362), .A(n19745), .ZN(n22141) );
  AND2_X2 U946 ( .A1(n169), .A2(n168), .ZN(n16579) );
  AND2_X2 U2662 ( .A1(n17776), .A2(n17777), .ZN(n19481) );
  AND2_X2 U1329 ( .A1(n6743), .A2(n4733), .ZN(n4298) );
  OAI21_X2 U2891 ( .B1(n15180), .B2(n15181), .A(n15179), .ZN(n15850) );
  XNOR2_X2 U424 ( .A(n21206), .B(n21205), .ZN(n23131) );
  XNOR2_X2 U1716 ( .A(n15455), .B(n15454), .ZN(n17415) );
  OAI21_X2 U21723 ( .B1(n18394), .B2(n18393), .A(n18392), .ZN(n18863) );
  XNOR2_X2 U14473 ( .A(n6997), .B(Key[122]), .ZN(n7909) );
  NAND3_X1 U1413 ( .A1(n4584), .A2(n7442), .A3(n7443), .ZN(n9754) );
  NAND3_X1 U12843 ( .A1(n9061), .A2(n9062), .A3(n9060), .ZN(n5537) );
  OAI211_X1 U16942 ( .C1(n11322), .C2(n11181), .A(n10475), .B(n10474), .ZN(
        n12338) );
  AND2_X1 U3114 ( .A1(n11428), .A2(n11426), .ZN(n11487) );
  NAND3_X1 U1072 ( .A1(n10885), .A2(n11028), .A3(n10886), .ZN(n12164) );
  AND2_X1 U8134 ( .A1(n2295), .A2(n2294), .ZN(n15423) );
  OAI21_X1 U5546 ( .B1(n15232), .B2(n15231), .A(n15230), .ZN(n16271) );
  NAND4_X1 U19506 ( .A1(n14649), .A2(n14648), .A3(n14647), .A4(n14646), .ZN(
        n15817) );
  AND3_X1 U109 ( .A1(n16672), .A2(n16671), .A3(n16670), .ZN(n17947) );
  OAI21_X1 U3609 ( .B1(n19811), .B2(n20285), .A(n19813), .ZN(n20864) );
  NAND3_X1 U13021 ( .A1(n24571), .A2(n24570), .A3(n24569), .ZN(n25696) );
  OAI21_X2 U1664 ( .B1(n26444), .B2(n26950), .A(n26443), .ZN(n27300) );
  AOI21_X1 U10 ( .B1(n21225), .B2(n21224), .A(n21223), .ZN(n28517) );
  AND2_X1 U11 ( .A1(n17060), .A2(n18337), .ZN(n29204) );
  BUF_X1 U28 ( .A(n10816), .Z(n28157) );
  BUF_X1 U151 ( .A(n10472), .Z(n11183) );
  AND4_X2 U203 ( .A1(n20731), .A2(n20732), .A3(n20730), .A4(n4776), .ZN(n21990) );
  INV_X2 U236 ( .A(n15400), .ZN(n28196) );
  OAI211_X2 U238 ( .C1(n5956), .C2(n5285), .A(n5284), .B(n5283), .ZN(n15183)
         );
  AND2_X2 U240 ( .A1(n16848), .A2(n16849), .ZN(n18423) );
  MUX2_X2 U265 ( .A(n23869), .B(n23868), .S(n24720), .Z(n26040) );
  AOI21_X2 U266 ( .B1(n14711), .B2(n14598), .A(n14710), .ZN(n16568) );
  AND3_X2 U283 ( .A1(n3245), .A2(n23616), .A3(n23617), .ZN(n24791) );
  OAI211_X1 U330 ( .C1(n14006), .C2(n14007), .A(n6106), .B(n6105), .ZN(n15431)
         );
  XNOR2_X1 U345 ( .A(n16449), .B(n16305), .ZN(n16154) );
  BUF_X1 U349 ( .A(n22953), .Z(n23846) );
  BUF_X1 U356 ( .A(n20207), .Z(n21674) );
  OAI211_X1 U357 ( .C1(n17905), .C2(n18456), .A(n3865), .B(n3864), .ZN(n19346)
         );
  BUF_X1 U358 ( .A(n26452), .Z(n29105) );
  NOR2_X1 U363 ( .A1(n15334), .A2(n15338), .ZN(n28766) );
  NOR2_X1 U376 ( .A1(n14569), .A2(n15071), .ZN(n28767) );
  XOR2_X1 U382 ( .A(n15330), .B(n15329), .Z(n28768) );
  OAI21_X2 U387 ( .B1(n19876), .B2(n19985), .A(n19875), .ZN(n21159) );
  NOR2_X2 U389 ( .A1(n24774), .A2(n24773), .ZN(n29046) );
  XNOR2_X2 U407 ( .A(n25524), .B(n25523), .ZN(n29058) );
  OAI21_X2 U415 ( .B1(n5546), .B2(n26771), .A(n6769), .ZN(n27497) );
  OAI21_X2 U416 ( .B1(n27116), .B2(n27115), .A(n27114), .ZN(n29049) );
  OAI211_X2 U422 ( .C1(n17523), .C2(n18220), .A(n17533), .B(n1943), .ZN(n19377) );
  OAI211_X2 U427 ( .C1(n8771), .C2(n8770), .A(n8769), .B(n8768), .ZN(n9908) );
  XNOR2_X2 U434 ( .A(n13508), .B(n13507), .ZN(n14036) );
  OAI211_X1 U441 ( .C1(n23072), .C2(n24712), .A(n29249), .B(n29248), .ZN(
        n25908) );
  NAND3_X2 U458 ( .A1(n3857), .A2(n3858), .A3(n21189), .ZN(n22068) );
  NOR2_X2 U465 ( .A1(n21238), .A2(n952), .ZN(n22278) );
  NAND3_X2 U481 ( .A1(n28274), .A2(n1654), .A3(n1424), .ZN(n26070) );
  XNOR2_X1 U495 ( .A(Plaintext[137]), .B(Key[137]), .ZN(n8300) );
  NAND2_X2 U508 ( .A1(n3647), .A2(n3646), .ZN(n13338) );
  BUF_X1 U528 ( .A(n17175), .Z(n28775) );
  CLKBUF_X1 U530 ( .A(n17175), .Z(n28776) );
  XNOR2_X1 U531 ( .A(n16357), .B(n16356), .ZN(n17175) );
  AND2_X1 U573 ( .A1(n572), .A2(n11754), .ZN(n28878) );
  AND2_X2 U578 ( .A1(n6084), .A2(n6082), .ZN(n21448) );
  OAI211_X2 U597 ( .C1(n9167), .C2(n9163), .A(n8317), .B(n8316), .ZN(n28488)
         );
  NAND2_X2 U604 ( .A1(n828), .A2(n829), .ZN(n15515) );
  AND2_X1 U620 ( .A1(n25418), .A2(n26576), .ZN(n26574) );
  XNOR2_X1 U622 ( .A(n9576), .B(n9577), .ZN(n9933) );
  XNOR2_X2 U628 ( .A(n18971), .B(n18970), .ZN(n20219) );
  NAND2_X2 U637 ( .A1(n6557), .A2(n6558), .ZN(n23126) );
  XNOR2_X2 U639 ( .A(n9483), .B(n9482), .ZN(n2690) );
  NAND3_X2 U696 ( .A1(n2312), .A2(n1962), .A3(n3492), .ZN(n22628) );
  NOR2_X2 U719 ( .A1(n18352), .A2(n5920), .ZN(n18900) );
  XNOR2_X2 U725 ( .A(n10400), .B(n10399), .ZN(n10431) );
  INV_X2 U747 ( .A(n852), .ZN(n27357) );
  XNOR2_X2 U750 ( .A(n22367), .B(n22366), .ZN(n23621) );
  XNOR2_X1 U787 ( .A(n17684), .B(n19336), .ZN(n28140) );
  XNOR2_X2 U790 ( .A(n7007), .B(Key[69]), .ZN(n7846) );
  XNOR2_X1 U811 ( .A(n9022), .B(n9021), .ZN(n5595) );
  NOR2_X2 U820 ( .A1(n21434), .A2(n4311), .ZN(n22333) );
  AOI21_X2 U829 ( .B1(n10600), .B2(n10601), .A(n10599), .ZN(n11740) );
  BUF_X2 U891 ( .A(n24650), .Z(n28785) );
  OAI211_X1 U906 ( .C1(n23749), .C2(n23215), .A(n5041), .B(n3631), .ZN(n24650)
         );
  NAND3_X2 U929 ( .A1(n5609), .A2(n5610), .A3(n15646), .ZN(n18489) );
  XNOR2_X2 U934 ( .A(n6968), .B(Key[103]), .ZN(n7619) );
  OAI211_X2 U950 ( .C1(n13128), .C2(n15082), .A(n13127), .B(n4169), .ZN(n16476) );
  NAND3_X2 U951 ( .A1(n28938), .A2(n8997), .A3(n3056), .ZN(n9639) );
  NOR2_X2 U963 ( .A1(n24495), .A2(n24494), .ZN(n25849) );
  XNOR2_X2 U977 ( .A(n19581), .B(n19580), .ZN(n20323) );
  XNOR2_X2 U995 ( .A(n15570), .B(n15569), .ZN(n17336) );
  XNOR2_X2 U1018 ( .A(n9182), .B(n9181), .ZN(n11347) );
  OAI21_X2 U1035 ( .B1(n19781), .B2(n19754), .A(n19753), .ZN(n22145) );
  NOR2_X2 U1036 ( .A1(n21247), .A2(n21246), .ZN(n22204) );
  XNOR2_X2 U1087 ( .A(n7043), .B(Key[151]), .ZN(n7981) );
  OAI211_X2 U1112 ( .C1(n8209), .C2(n7842), .A(n1612), .B(n28365), .ZN(n8908)
         );
  INV_X1 U1128 ( .A(n24668), .ZN(n4195) );
  NAND3_X1 U1131 ( .A1(n21641), .A2(n21640), .A3(n3313), .ZN(n22180) );
  INV_X1 U1138 ( .A(n22023), .ZN(n28790) );
  INV_X1 U1147 ( .A(n21327), .ZN(n28791) );
  OR2_X2 U1164 ( .A1(n20741), .A2(n20736), .ZN(n20858) );
  NAND3_X1 U1168 ( .A1(n2135), .A2(n2136), .A3(n18191), .ZN(n19486) );
  INV_X2 U1170 ( .A(n17798), .ZN(n18456) );
  INV_X1 U1175 ( .A(n5891), .ZN(n28792) );
  INV_X1 U1177 ( .A(n17354), .ZN(n28793) );
  INV_X1 U1192 ( .A(n12354), .ZN(n29209) );
  INV_X1 U1201 ( .A(n10875), .ZN(n11220) );
  NAND2_X1 U1211 ( .A1(n8562), .A2(n9144), .ZN(n8937) );
  CLKBUF_X1 U1217 ( .A(Key[171]), .Z(n2986) );
  CLKBUF_X1 U1219 ( .A(Key[89]), .Z(n2477) );
  CLKBUF_X1 U1229 ( .A(Key[185]), .Z(n2465) );
  CLKBUF_X1 U1234 ( .A(Key[189]), .Z(n3554) );
  CLKBUF_X1 U1236 ( .A(Key[59]), .Z(n3223) );
  AND2_X1 U1263 ( .A1(n4485), .A2(n27047), .ZN(n27092) );
  AND2_X1 U1268 ( .A1(n29029), .A2(n29030), .ZN(n27944) );
  OAI21_X1 U1279 ( .B1(n26253), .B2(n26735), .A(n26252), .ZN(n28066) );
  BUF_X1 U1315 ( .A(n25465), .Z(n25782) );
  OAI21_X1 U1316 ( .B1(n23144), .B2(n24229), .A(n24895), .ZN(n25134) );
  NAND3_X1 U1339 ( .A1(n5293), .A2(n5292), .A3(n22499), .ZN(n29109) );
  INV_X1 U1340 ( .A(n5763), .ZN(n23284) );
  OR2_X1 U1344 ( .A1(n22877), .A2(n23810), .ZN(n5763) );
  INV_X1 U1372 ( .A(n23317), .ZN(n28963) );
  BUF_X1 U1388 ( .A(n23250), .Z(n28796) );
  AND2_X1 U1390 ( .A1(n22174), .A2(n23587), .ZN(n28824) );
  XNOR2_X1 U1398 ( .A(n21916), .B(n21915), .ZN(n23795) );
  OAI21_X1 U1409 ( .B1(n21153), .B2(n21152), .A(n21151), .ZN(n22419) );
  OR2_X1 U1424 ( .A1(n21462), .A2(n21457), .ZN(n28941) );
  OAI21_X1 U1426 ( .B1(n20998), .B2(n21217), .A(n28979), .ZN(n18788) );
  AND2_X1 U1427 ( .A1(n4344), .A2(n28937), .ZN(n21321) );
  NOR2_X1 U1434 ( .A1(n22025), .A2(n22026), .ZN(n22028) );
  NAND4_X1 U1435 ( .A1(n21217), .A2(n21218), .A3(n19914), .A4(n28980), .ZN(
        n28979) );
  AND2_X1 U1462 ( .A1(n21135), .A2(n21134), .ZN(n28937) );
  INV_X1 U1463 ( .A(n21394), .ZN(n28797) );
  AND3_X1 U1466 ( .A1(n28812), .A2(n29182), .A3(n29180), .ZN(n21749) );
  OAI21_X1 U1498 ( .B1(n28133), .B2(n20517), .A(n28992), .ZN(n19457) );
  XNOR2_X1 U1522 ( .A(n19121), .B(n19120), .ZN(n20498) );
  XNOR2_X1 U1527 ( .A(n19346), .B(n19486), .ZN(n19141) );
  AND2_X1 U1534 ( .A1(n1708), .A2(n18177), .ZN(n28981) );
  NAND3_X1 U1537 ( .A1(n28827), .A2(n28826), .A3(n17999), .ZN(n19428) );
  NAND2_X1 U1541 ( .A1(n17785), .A2(n28978), .ZN(n19378) );
  NAND3_X1 U1567 ( .A1(n18080), .A2(n18079), .A3(n46), .ZN(n19448) );
  OAI211_X1 U1588 ( .C1(n15939), .C2(n15938), .A(n15936), .B(n29007), .ZN(
        n19403) );
  AND2_X1 U1591 ( .A1(n18423), .A2(n17802), .ZN(n29274) );
  OR2_X1 U1600 ( .A1(n16985), .A2(n18188), .ZN(n29199) );
  OR2_X1 U1601 ( .A1(n18170), .A2(n4044), .ZN(n5203) );
  NAND2_X1 U1605 ( .A1(n29203), .A2(n4583), .ZN(n18338) );
  INV_X1 U1616 ( .A(n18135), .ZN(n526) );
  NAND2_X1 U1618 ( .A1(n16708), .A2(n1129), .ZN(n18198) );
  AND2_X1 U1620 ( .A1(n28831), .A2(n2600), .ZN(n17132) );
  NAND2_X1 U1630 ( .A1(n1088), .A2(n16818), .ZN(n18172) );
  OR2_X1 U1631 ( .A1(n2600), .A2(n17129), .ZN(n5733) );
  INV_X1 U1653 ( .A(n17455), .ZN(n28801) );
  NAND3_X1 U1670 ( .A1(n28816), .A2(n1164), .A3(n28818), .ZN(n16160) );
  AND3_X1 U1694 ( .A1(n29012), .A2(n29011), .A3(n29010), .ZN(n16395) );
  NAND2_X1 U1696 ( .A1(n14951), .A2(n28896), .ZN(n15999) );
  NOR2_X1 U1720 ( .A1(n14682), .A2(n14681), .ZN(n15802) );
  NOR2_X1 U1721 ( .A1(n14952), .A2(n15082), .ZN(n28897) );
  OR2_X1 U1735 ( .A1(n14990), .A2(n14989), .ZN(n3208) );
  AND3_X1 U1745 ( .A1(n734), .A2(n735), .A3(n12936), .ZN(n15082) );
  INV_X1 U1747 ( .A(n15333), .ZN(n28802) );
  BUF_X2 U1748 ( .A(n14981), .Z(n28803) );
  OR2_X1 U1750 ( .A1(n13699), .A2(n13306), .ZN(n28950) );
  AND2_X1 U1762 ( .A1(n13826), .A2(n14354), .ZN(n28899) );
  INV_X1 U1809 ( .A(n14401), .ZN(n28804) );
  INV_X1 U1842 ( .A(n14455), .ZN(n28806) );
  NAND2_X1 U1859 ( .A1(n2319), .A2(n11850), .ZN(n12872) );
  NAND3_X1 U1890 ( .A1(n29264), .A2(n11841), .A3(n4447), .ZN(n12787) );
  OR2_X1 U1926 ( .A1(n12030), .A2(n12031), .ZN(n1192) );
  OAI22_X1 U1939 ( .A1(n12299), .A2(n12300), .B1(n11769), .B2(n4197), .ZN(
        n5020) );
  OR2_X1 U1956 ( .A1(n11553), .A2(n11785), .ZN(n29291) );
  AND3_X1 U1974 ( .A1(n28811), .A2(n3449), .A3(n6361), .ZN(n11751) );
  INV_X1 U1983 ( .A(n569), .ZN(n28807) );
  NAND3_X1 U2108 ( .A1(n2868), .A2(n2867), .A3(n6242), .ZN(n11921) );
  AND2_X1 U2207 ( .A1(n8109), .A2(n9245), .ZN(n28911) );
  NAND2_X1 U2216 ( .A1(n2310), .A2(n7346), .ZN(n8185) );
  AND2_X1 U2219 ( .A1(n2695), .A2(n28814), .ZN(n8490) );
  INV_X1 U2262 ( .A(n8810), .ZN(n28808) );
  NAND2_X1 U2265 ( .A1(n29214), .A2(n7790), .ZN(n8353) );
  NAND4_X1 U2301 ( .A1(n7668), .A2(n901), .A3(n7667), .A4(n7666), .ZN(n8777)
         );
  MUX2_X1 U2306 ( .A(n7143), .B(n7142), .S(n7523), .Z(n28913) );
  OR2_X1 U2329 ( .A1(n7775), .A2(n7891), .ZN(n5494) );
  XNOR2_X1 U2331 ( .A(n6971), .B(Key[106]), .ZN(n7358) );
  INV_X1 U2374 ( .A(n9113), .ZN(n28810) );
  OR2_X1 U2377 ( .A1(n7017), .A2(n7690), .ZN(n7502) );
  CLKBUF_X1 U2435 ( .A(n7851), .Z(n371) );
  OR2_X1 U2445 ( .A1(n8034), .A2(n7508), .ZN(n8039) );
  AOI21_X1 U2458 ( .B1(n9436), .B2(n8998), .A(n9438), .ZN(n28989) );
  OR2_X1 U2459 ( .A1(n8868), .A2(n2006), .ZN(n3788) );
  INV_X1 U2463 ( .A(n8490), .ZN(n9099) );
  OAI211_X1 U2477 ( .C1(n8036), .C2(n7514), .A(n7513), .B(n7512), .ZN(n8817)
         );
  OAI211_X1 U2496 ( .C1(n8808), .C2(n28808), .A(n29242), .B(n29241), .ZN(n2899) );
  AND2_X1 U2510 ( .A1(n9213), .A2(n9212), .ZN(n28858) );
  XNOR2_X1 U2540 ( .A(n10037), .B(n9383), .ZN(n10421) );
  AND2_X1 U2558 ( .A1(n10808), .A2(n11149), .ZN(n29263) );
  XNOR2_X1 U2578 ( .A(n10142), .B(n10141), .ZN(n11084) );
  INV_X1 U2580 ( .A(n12313), .ZN(n12051) );
  NAND2_X1 U2617 ( .A1(n10270), .A2(n28929), .ZN(n28928) );
  OR2_X1 U2654 ( .A1(n11486), .A2(n6482), .ZN(n11793) );
  OR2_X1 U2669 ( .A1(n12356), .A2(n11739), .ZN(n919) );
  AND2_X1 U2693 ( .A1(n11656), .A2(n28828), .ZN(n11844) );
  MUX2_X1 U2749 ( .A(n10607), .B(n10606), .S(n10605), .Z(n10608) );
  OR2_X1 U2765 ( .A1(n11853), .A2(n10905), .ZN(n10906) );
  AND2_X1 U2766 ( .A1(n11658), .A2(n11657), .ZN(n28828) );
  OR2_X1 U2794 ( .A1(n11911), .A2(n12363), .ZN(n28961) );
  OAI21_X1 U2800 ( .B1(n11639), .B2(n11672), .A(n11671), .ZN(n11518) );
  OR2_X1 U2806 ( .A1(n11394), .A2(n11852), .ZN(n28886) );
  OR2_X1 U2815 ( .A1(n11686), .A2(n12000), .ZN(n29175) );
  AND2_X1 U2817 ( .A1(n11380), .A2(n11379), .ZN(n28917) );
  INV_X1 U2819 ( .A(n29244), .ZN(n29243) );
  NAND3_X1 U2850 ( .A1(n11160), .A2(n11161), .A3(n1140), .ZN(n13249) );
  BUF_X1 U2920 ( .A(n14171), .Z(n29097) );
  AOI21_X1 U2944 ( .B1(n6032), .B2(n13587), .A(n58), .ZN(n14041) );
  OR2_X1 U2985 ( .A1(n12744), .A2(n14465), .ZN(n28936) );
  OR2_X1 U2987 ( .A1(n14380), .A2(n14004), .ZN(n14005) );
  OR2_X1 U3063 ( .A1(n13824), .A2(n14126), .ZN(n14357) );
  OR2_X1 U3070 ( .A1(n14075), .A2(n14359), .ZN(n28952) );
  OAI21_X1 U3074 ( .B1(n14459), .B2(n13864), .A(n13863), .ZN(n15166) );
  NAND2_X1 U3076 ( .A1(n14490), .A2(n14489), .ZN(n15489) );
  INV_X1 U3088 ( .A(n15694), .ZN(n29011) );
  OR2_X1 U3100 ( .A1(n14837), .A2(n15290), .ZN(n14521) );
  NOR2_X1 U3121 ( .A1(n14601), .A2(n15284), .ZN(n28842) );
  NOR2_X1 U3134 ( .A1(n5596), .A2(n15172), .ZN(n28406) );
  OAI21_X1 U3151 ( .B1(n17160), .B2(n28497), .A(n17162), .ZN(n28852) );
  AND2_X1 U3175 ( .A1(n17282), .A2(n17283), .ZN(n29000) );
  INV_X1 U3185 ( .A(n17175), .ZN(n16874) );
  OR2_X1 U3242 ( .A1(n16614), .A2(n17496), .ZN(n28993) );
  AND2_X1 U3255 ( .A1(n4367), .A2(n4368), .ZN(n17126) );
  AND2_X1 U3261 ( .A1(n1880), .A2(n17249), .ZN(n968) );
  INV_X1 U3270 ( .A(n16837), .ZN(n17316) );
  OAI21_X1 U3280 ( .B1(n1090), .B2(n29000), .A(n29086), .ZN(n28999) );
  OR2_X1 U3309 ( .A1(n18710), .A2(n5023), .ZN(n3766) );
  AND4_X2 U3334 ( .A1(n16742), .A2(n16743), .A3(n16741), .A4(n16740), .ZN(
        n18277) );
  BUF_X1 U3361 ( .A(n18057), .Z(n1861) );
  OR2_X1 U3372 ( .A1(n17403), .A2(n16904), .ZN(n15934) );
  AOI22_X1 U3408 ( .A1(n1963), .A2(n17996), .B1(n18382), .B2(n17997), .ZN(
        n28826) );
  OR2_X1 U3449 ( .A1(n18349), .A2(n18000), .ZN(n28827) );
  NAND3_X1 U3476 ( .A1(n4120), .A2(n4119), .A3(n5992), .ZN(n18653) );
  XNOR2_X1 U3478 ( .A(n19603), .B(n18767), .ZN(n18768) );
  AND2_X1 U3548 ( .A1(n20148), .A2(n20146), .ZN(n28849) );
  OR2_X1 U3555 ( .A1(n21090), .A2(n5817), .ZN(n21931) );
  INV_X1 U3558 ( .A(n20286), .ZN(n29166) );
  XNOR2_X1 U3566 ( .A(n18917), .B(n18916), .ZN(n29134) );
  XNOR2_X1 U3573 ( .A(n19169), .B(n19168), .ZN(n20495) );
  OAI21_X1 U3596 ( .B1(n20307), .B2(n20305), .A(n19948), .ZN(n5194) );
  INV_X1 U3600 ( .A(n18919), .ZN(n4877) );
  OR2_X1 U3617 ( .A1(n29235), .A2(n20398), .ZN(n20402) );
  INV_X1 U3619 ( .A(n1875), .ZN(n28891) );
  OR2_X1 U3631 ( .A1(n21539), .A2(n21503), .ZN(n28991) );
  NAND2_X1 U3637 ( .A1(n19930), .A2(n29183), .ZN(n29182) );
  OR2_X1 U3638 ( .A1(n20459), .A2(n20273), .ZN(n29184) );
  CLKBUF_X1 U3639 ( .A(n28555), .Z(n20117) );
  OR2_X1 U3646 ( .A1(n20338), .A2(n29601), .ZN(n28982) );
  NOR3_X1 U3652 ( .A1(n20767), .A2(n29531), .A3(n20766), .ZN(n21153) );
  INV_X1 U3709 ( .A(n21376), .ZN(n29228) );
  OAI211_X1 U3786 ( .C1(n21553), .C2(n21547), .A(n1621), .B(n28890), .ZN(
        n21556) );
  INV_X1 U3817 ( .A(n21990), .ZN(n22763) );
  AND2_X1 U3826 ( .A1(n20712), .A2(n21269), .ZN(n29256) );
  OR2_X1 U3847 ( .A1(n23767), .A2(n23765), .ZN(n23333) );
  INV_X1 U3883 ( .A(n22078), .ZN(n28914) );
  OR2_X1 U3897 ( .A1(n23267), .A2(n28581), .ZN(n23217) );
  INV_X1 U3898 ( .A(n23353), .ZN(n4232) );
  BUF_X1 U3909 ( .A(n22877), .Z(n23808) );
  OR2_X1 U3910 ( .A1(n23493), .A2(n23795), .ZN(n23196) );
  MUX2_X1 U3920 ( .A(n23230), .B(n23229), .S(n22949), .Z(n23231) );
  INV_X1 U3966 ( .A(n24243), .ZN(n24239) );
  OR2_X1 U3990 ( .A1(n24246), .A2(n3061), .ZN(n29002) );
  OR2_X1 U3993 ( .A1(n24466), .A2(n24578), .ZN(n29013) );
  OR2_X1 U4017 ( .A1(n24612), .A2(n23922), .ZN(n4639) );
  OR2_X1 U4049 ( .A1(n462), .A2(n21303), .ZN(n29015) );
  MUX2_X1 U4086 ( .A(n24048), .B(n24047), .S(n469), .Z(n24049) );
  INV_X1 U4136 ( .A(n24532), .ZN(n24894) );
  AND3_X1 U4137 ( .A1(n24411), .A2(n24413), .A3(n24410), .ZN(n2261) );
  OAI21_X1 U4139 ( .B1(n4573), .B2(n4575), .A(n4572), .ZN(n24797) );
  AND2_X1 U4147 ( .A1(n26868), .A2(n26865), .ZN(n26870) );
  XNOR2_X1 U4152 ( .A(n25448), .B(n25447), .ZN(n26748) );
  BUF_X1 U4171 ( .A(n25365), .Z(n26489) );
  INV_X1 U4174 ( .A(n27382), .ZN(n29218) );
  OR2_X1 U4176 ( .A1(n27591), .A2(n27594), .ZN(n28967) );
  AND3_X1 U4204 ( .A1(n25048), .A2(n25047), .A3(n25050), .ZN(n28834) );
  CLKBUF_X1 U4221 ( .A(Key[71]), .Z(n3422) );
  XOR2_X1 U4274 ( .A(n10182), .B(n10181), .Z(n1851) );
  OR2_X1 U4285 ( .A1(n10740), .A2(n10806), .ZN(n28811) );
  OR2_X1 U4293 ( .A1(n19931), .A2(n5783), .ZN(n28812) );
  OR2_X1 U4307 ( .A1(n20395), .A2(n20400), .ZN(n28813) );
  AND2_X1 U4312 ( .A1(n4834), .A2(n4833), .ZN(n28814) );
  OR2_X1 U4330 ( .A1(n24978), .A2(n24976), .ZN(n28815) );
  OR2_X1 U4347 ( .A1(n15395), .A2(n14633), .ZN(n28816) );
  AND2_X1 U4357 ( .A1(n15233), .A2(n15234), .ZN(n28817) );
  INV_X1 U4368 ( .A(n7192), .ZN(n7644) );
  INV_X1 U4381 ( .A(n2238), .ZN(n29241) );
  NAND2_X1 U4382 ( .A1(n7622), .A2(n7623), .ZN(n9206) );
  INV_X1 U4397 ( .A(n14429), .ZN(n28986) );
  OR2_X1 U4405 ( .A1(n15391), .A2(n15390), .ZN(n28818) );
  XNOR2_X1 U4406 ( .A(n16049), .B(n16048), .ZN(n16860) );
  OR2_X1 U4415 ( .A1(n18170), .A2(n18168), .ZN(n28819) );
  XOR2_X1 U4419 ( .A(n18748), .B(n18747), .Z(n28820) );
  XNOR2_X1 U4426 ( .A(n19531), .B(n19530), .ZN(n20265) );
  INV_X1 U4427 ( .A(n20702), .ZN(n28980) );
  INV_X1 U4446 ( .A(n20619), .ZN(n28894) );
  INV_X1 U4451 ( .A(n21932), .ZN(n28916) );
  OR2_X1 U4455 ( .A1(n23209), .A2(n22984), .ZN(n28821) );
  OR2_X1 U4466 ( .A1(n26374), .A2(n26440), .ZN(n28822) );
  OR2_X1 U4476 ( .A1(n29330), .A2(n26800), .ZN(n28823) );
  NAND3_X1 U4481 ( .A1(n21157), .A2(n21156), .A3(n20744), .ZN(n19877) );
  NAND2_X1 U4488 ( .A1(n23715), .A2(n28824), .ZN(n23263) );
  NAND2_X1 U4494 ( .A1(n9057), .A2(n9058), .ZN(n9258) );
  NAND2_X1 U4498 ( .A1(n1174), .A2(n28825), .ZN(n11505) );
  OR2_X1 U4517 ( .A1(n11320), .A2(n4650), .ZN(n28825) );
  NAND2_X1 U4518 ( .A1(n15222), .A2(n15223), .ZN(n15351) );
  NAND3_X1 U4525 ( .A1(n21597), .A2(n21598), .A3(n5720), .ZN(n5719) );
  NAND3_X1 U4548 ( .A1(n10959), .A2(n10958), .A3(n10778), .ZN(n10603) );
  NAND3_X1 U4567 ( .A1(n11820), .A2(n4028), .A3(n11816), .ZN(n11823) );
  NAND2_X1 U4569 ( .A1(n8234), .A2(n7358), .ZN(n8239) );
  NAND2_X1 U4578 ( .A1(n23969), .A2(n24479), .ZN(n23553) );
  NAND2_X1 U4585 ( .A1(n24046), .A2(n23968), .ZN(n23969) );
  INV_X1 U4618 ( .A(n17070), .ZN(n17072) );
  NAND2_X1 U4661 ( .A1(n17829), .A2(n4270), .ZN(n17070) );
  NOR2_X1 U4678 ( .A1(n23311), .A2(n28829), .ZN(n28358) );
  INV_X1 U4688 ( .A(n23556), .ZN(n28829) );
  NAND2_X1 U4701 ( .A1(n23628), .A2(n23309), .ZN(n23556) );
  OAI21_X1 U4720 ( .B1(n17616), .B2(n17615), .A(n17613), .ZN(n17306) );
  NAND3_X1 U4754 ( .A1(n17305), .A2(n29152), .A3(n17421), .ZN(n17613) );
  MUX2_X1 U4759 ( .A(n27425), .B(n27429), .S(n27424), .Z(n27431) );
  NAND2_X1 U4774 ( .A1(n28491), .A2(n501), .ZN(n20021) );
  OAI21_X2 U4779 ( .B1(n20465), .B2(n21534), .A(n20464), .ZN(n22302) );
  OAI211_X1 U4789 ( .C1(n20218), .C2(n20496), .A(n6834), .B(n20217), .ZN(n2798) );
  NAND2_X1 U4792 ( .A1(n20496), .A2(n20493), .ZN(n20217) );
  XNOR2_X1 U4816 ( .A(n5809), .B(n28830), .ZN(n21353) );
  XNOR2_X1 U4841 ( .A(n19424), .B(n19425), .ZN(n28830) );
  NAND3_X1 U4857 ( .A1(n459), .A2(n5168), .A3(n24017), .ZN(n5218) );
  NAND2_X1 U4865 ( .A1(n6423), .A2(n6424), .ZN(n3459) );
  NAND2_X1 U4881 ( .A1(n24142), .A2(n24144), .ZN(n23931) );
  AND3_X2 U4902 ( .A1(n3538), .A2(n17905), .A3(n3539), .ZN(n19626) );
  NAND2_X1 U4905 ( .A1(n1337), .A2(n4801), .ZN(n10527) );
  NAND2_X1 U4917 ( .A1(n28801), .A2(n16797), .ZN(n2600) );
  NAND2_X1 U4918 ( .A1(n17128), .A2(n17451), .ZN(n28831) );
  NAND3_X2 U4934 ( .A1(n28832), .A2(n7419), .A3(n7417), .ZN(n9996) );
  NAND2_X1 U4957 ( .A1(n7416), .A2(n714), .ZN(n28832) );
  NAND3_X1 U4964 ( .A1(n2464), .A2(n4907), .A3(n11205), .ZN(n28875) );
  NAND2_X1 U4984 ( .A1(n25052), .A2(n28833), .ZN(Ciphertext[100]) );
  NAND2_X1 U5006 ( .A1(n25049), .A2(n28834), .ZN(n28833) );
  NAND2_X1 U5040 ( .A1(n9070), .A2(n8857), .ZN(n9069) );
  NAND3_X1 U5076 ( .A1(n5544), .A2(n21565), .A3(n20862), .ZN(n2918) );
  NAND3_X1 U5106 ( .A1(n18032), .A2(n18160), .A3(n18156), .ZN(n28973) );
  NAND2_X1 U5158 ( .A1(n17866), .A2(n28836), .ZN(n17870) );
  NAND3_X1 U5160 ( .A1(n511), .A2(n5690), .A3(n18216), .ZN(n28836) );
  NAND2_X1 U5171 ( .A1(n17485), .A2(n5737), .ZN(n5736) );
  NAND2_X1 U5172 ( .A1(n21198), .A2(n21509), .ZN(n21535) );
  NAND2_X1 U5174 ( .A1(n15237), .A2(n694), .ZN(n28837) );
  NAND2_X1 U5176 ( .A1(n5266), .A2(n10681), .ZN(n28838) );
  NAND2_X1 U5178 ( .A1(n5264), .A2(n10970), .ZN(n28839) );
  OAI21_X1 U5185 ( .B1(n8971), .B2(n8970), .A(n28840), .ZN(n9540) );
  NAND2_X1 U5210 ( .A1(n8969), .A2(n8968), .ZN(n28840) );
  NAND3_X2 U5218 ( .A1(n15287), .A2(n5930), .A3(n28841), .ZN(n16575) );
  NAND2_X1 U5224 ( .A1(n14696), .A2(n28842), .ZN(n28841) );
  NAND2_X1 U5235 ( .A1(n7814), .A2(n2273), .ZN(n8064) );
  NAND2_X1 U5294 ( .A1(n136), .A2(n23514), .ZN(n28844) );
  NOR2_X1 U5307 ( .A1(n8540), .A2(n6901), .ZN(n28845) );
  AND2_X2 U5327 ( .A1(n28847), .A2(n6394), .ZN(n22363) );
  NAND3_X1 U5353 ( .A1(n6396), .A2(n21272), .A3(n6397), .ZN(n28847) );
  NAND2_X1 U5355 ( .A1(n830), .A2(n14273), .ZN(n828) );
  NAND2_X1 U5363 ( .A1(n827), .A2(n14361), .ZN(n830) );
  NAND2_X1 U5365 ( .A1(n7248), .A2(n8052), .ZN(n1010) );
  OR2_X1 U5409 ( .A1(n8381), .A2(n8735), .ZN(n7575) );
  AND3_X2 U5460 ( .A1(n9816), .A2(n9814), .A3(n9815), .ZN(n11819) );
  AND2_X1 U5461 ( .A1(n9438), .A2(n8995), .ZN(n29221) );
  NAND2_X1 U5526 ( .A1(n6894), .A2(n28848), .ZN(n19012) );
  NAND2_X1 U5529 ( .A1(n20145), .A2(n28849), .ZN(n28848) );
  NAND2_X1 U5535 ( .A1(n20985), .A2(n20913), .ZN(n20921) );
  NAND2_X1 U5536 ( .A1(n27480), .A2(n27492), .ZN(n27475) );
  OAI21_X1 U5545 ( .B1(n24977), .B2(n24258), .A(n28815), .ZN(n24981) );
  INV_X1 U5554 ( .A(n8794), .ZN(n4839) );
  NAND2_X1 U5580 ( .A1(n9037), .A2(n9034), .ZN(n8794) );
  INV_X1 U5583 ( .A(n28852), .ZN(n28851) );
  NAND2_X1 U5602 ( .A1(n28853), .A2(n11261), .ZN(n3326) );
  NAND2_X1 U5633 ( .A1(n2754), .A2(n2755), .ZN(n28853) );
  NAND2_X1 U5634 ( .A1(n28855), .A2(n28854), .ZN(n23133) );
  NAND2_X1 U5668 ( .A1(n23366), .A2(n23364), .ZN(n28854) );
  NAND2_X1 U5675 ( .A1(n2921), .A2(n28604), .ZN(n28855) );
  NAND2_X1 U5700 ( .A1(n986), .A2(n988), .ZN(n5445) );
  NOR2_X2 U5710 ( .A1(n6198), .A2(n24298), .ZN(n25760) );
  NAND2_X1 U5718 ( .A1(n11274), .A2(n11034), .ZN(n11035) );
  NAND2_X1 U5726 ( .A1(n14569), .A2(n14570), .ZN(n6320) );
  NAND2_X1 U5742 ( .A1(n14967), .A2(n14964), .ZN(n28856) );
  NAND2_X1 U5747 ( .A1(n7658), .A2(n7659), .ZN(n28857) );
  NAND2_X1 U5763 ( .A1(n3325), .A2(n3326), .ZN(n11887) );
  INV_X1 U5897 ( .A(n1096), .ZN(n1356) );
  NAND3_X1 U5914 ( .A1(n28950), .A2(n13309), .A3(n13697), .ZN(n1096) );
  OR2_X1 U5941 ( .A1(n14349), .A2(n14354), .ZN(n6511) );
  NAND2_X1 U5953 ( .A1(n3911), .A2(n20049), .ZN(n20050) );
  OAI21_X2 U5980 ( .B1(n9215), .B2(n9214), .A(n28858), .ZN(n10356) );
  NAND3_X1 U5996 ( .A1(n22996), .A2(n23643), .A3(n23641), .ZN(n22258) );
  NAND2_X1 U6046 ( .A1(n9201), .A2(n9206), .ZN(n28860) );
  INV_X1 U6089 ( .A(n9206), .ZN(n28862) );
  NAND2_X1 U6146 ( .A1(n16602), .A2(n17518), .ZN(n3811) );
  NAND3_X1 U6188 ( .A1(n5333), .A2(n6509), .A3(n6508), .ZN(n21483) );
  NAND2_X1 U6231 ( .A1(n18128), .A2(n18124), .ZN(n18127) );
  OAI211_X2 U6236 ( .C1(n12260), .C2(n12261), .A(n12258), .B(n28863), .ZN(
        n12762) );
  OAI211_X1 U6309 ( .C1(n13993), .C2(n14578), .A(n15098), .B(n28864), .ZN(
        n12629) );
  NAND2_X1 U6327 ( .A1(n14578), .A2(n15097), .ZN(n28864) );
  NAND2_X1 U6393 ( .A1(n13358), .A2(n13914), .ZN(n28866) );
  NAND2_X1 U6406 ( .A1(n24602), .A2(n24734), .ZN(n5454) );
  NAND2_X1 U6434 ( .A1(n1992), .A2(n6663), .ZN(n3239) );
  NAND2_X1 U6442 ( .A1(n4979), .A2(n17181), .ZN(n16707) );
  AOI21_X1 U6443 ( .B1(n2286), .B2(n23697), .A(n28867), .ZN(n6942) );
  NAND2_X1 U6444 ( .A1(n23532), .A2(n6903), .ZN(n28867) );
  NOR2_X2 U6556 ( .A1(n13743), .A2(n4026), .ZN(n15382) );
  XNOR2_X1 U6578 ( .A(n28869), .B(n19210), .ZN(n19213) );
  INV_X1 U6611 ( .A(n19212), .ZN(n28869) );
  INV_X1 U6683 ( .A(n694), .ZN(n28871) );
  NAND2_X1 U6689 ( .A1(n28766), .A2(n694), .ZN(n28872) );
  NAND2_X1 U6737 ( .A1(n26984), .A2(n28019), .ZN(n28005) );
  NAND2_X1 U6773 ( .A1(n24228), .A2(n24532), .ZN(n24895) );
  NAND2_X1 U6808 ( .A1(n5030), .A2(n484), .ZN(n5029) );
  AND2_X1 U6809 ( .A1(n18107), .A2(n18106), .ZN(n29156) );
  NAND3_X1 U6849 ( .A1(n28874), .A2(n12299), .A3(n11767), .ZN(n11366) );
  NAND2_X1 U6856 ( .A1(n11769), .A2(n12302), .ZN(n28874) );
  NAND3_X1 U6864 ( .A1(n1657), .A2(n17258), .A3(n1574), .ZN(n16670) );
  NAND2_X1 U6865 ( .A1(n28875), .A2(n11208), .ZN(n12053) );
  NAND3_X1 U6895 ( .A1(n28627), .A2(n10806), .A3(n28876), .ZN(n10543) );
  INV_X1 U6899 ( .A(n10808), .ZN(n28876) );
  NAND2_X1 U6919 ( .A1(n10726), .A2(n1879), .ZN(n10727) );
  NAND2_X1 U6942 ( .A1(n2194), .A2(n2748), .ZN(n2193) );
  NAND2_X1 U6944 ( .A1(n2649), .A2(n24390), .ZN(n24691) );
  NAND3_X1 U6959 ( .A1(n893), .A2(n14833), .A3(n15036), .ZN(n14097) );
  NAND2_X1 U7110 ( .A1(n3849), .A2(n28241), .ZN(n28877) );
  NAND2_X1 U7124 ( .A1(n11686), .A2(n28878), .ZN(n11687) );
  AOI21_X1 U7126 ( .B1(n28879), .B2(n15466), .A(n15464), .ZN(n15467) );
  NAND2_X1 U7178 ( .A1(n4515), .A2(n15463), .ZN(n28879) );
  NAND2_X1 U7349 ( .A1(n11954), .A2(n4018), .ZN(n4017) );
  OAI22_X1 U7372 ( .A1(n2137), .A2(n58), .B1(n13999), .B2(n5918), .ZN(n6446)
         );
  NAND2_X1 U7390 ( .A1(n14036), .A2(n29089), .ZN(n2137) );
  NAND2_X1 U7391 ( .A1(n20886), .A2(n21587), .ZN(n21589) );
  NAND2_X1 U7509 ( .A1(n2250), .A2(n8350), .ZN(n28882) );
  OAI22_X2 U7620 ( .A1(n17871), .A2(n18063), .B1(n18303), .B2(n18061), .ZN(
        n19727) );
  OAI211_X2 U7683 ( .C1(n8766), .C2(n8765), .A(n9564), .B(n2168), .ZN(n9710)
         );
  AOI22_X1 U7695 ( .A1(n15074), .A2(n15073), .B1(n15076), .B2(n15075), .ZN(
        n15080) );
  NAND2_X1 U7709 ( .A1(n24653), .A2(n3061), .ZN(n24245) );
  OR2_X2 U7722 ( .A1(n23225), .A2(n23224), .ZN(n3061) );
  NOR2_X2 U7732 ( .A1(n26626), .A2(n5685), .ZN(n27977) );
  NAND2_X1 U7744 ( .A1(n5686), .A2(n5687), .ZN(n5685) );
  INV_X1 U7747 ( .A(n15980), .ZN(n539) );
  XNOR2_X1 U7748 ( .A(n15979), .B(n6455), .ZN(n15980) );
  NAND2_X1 U7771 ( .A1(n13615), .A2(n3346), .ZN(n15001) );
  OAI21_X1 U7796 ( .B1(n16936), .B2(n16935), .A(n17155), .ZN(n28883) );
  NAND2_X1 U7898 ( .A1(n21656), .A2(n20833), .ZN(n2641) );
  NAND2_X1 U7939 ( .A1(n28005), .A2(n28885), .ZN(n26986) );
  NAND2_X1 U7985 ( .A1(n28017), .A2(n445), .ZN(n28885) );
  NOR2_X2 U8008 ( .A1(n10967), .A2(n10968), .ZN(n349) );
  NAND2_X1 U8016 ( .A1(n11393), .A2(n28886), .ZN(n13025) );
  NAND2_X1 U8042 ( .A1(n3509), .A2(n29150), .ZN(n28887) );
  NAND2_X1 U8055 ( .A1(n28888), .A2(n4951), .ZN(n22862) );
  NAND2_X1 U8082 ( .A1(n29175), .A2(n11478), .ZN(n12954) );
  OR2_X1 U8096 ( .A1(n10913), .A2(n10735), .ZN(n10607) );
  NAND3_X1 U8149 ( .A1(n11215), .A2(n11216), .A3(n11214), .ZN(n12313) );
  NAND2_X1 U8193 ( .A1(n37), .A2(n39), .ZN(n11326) );
  NAND2_X1 U8198 ( .A1(n8177), .A2(n8173), .ZN(n7290) );
  OAI21_X2 U8203 ( .B1(n16840), .B2(n16839), .A(n28889), .ZN(n18190) );
  NAND2_X1 U8229 ( .A1(n1405), .A2(n29550), .ZN(n28889) );
  NAND2_X1 U8239 ( .A1(n21547), .A2(n28891), .ZN(n28890) );
  NAND2_X1 U8262 ( .A1(n15207), .A2(n15202), .ZN(n5515) );
  NAND2_X1 U8269 ( .A1(n20346), .A2(n20347), .ZN(n20348) );
  NAND2_X1 U8289 ( .A1(n28489), .A2(n20511), .ZN(n20347) );
  NAND3_X2 U8350 ( .A1(n13634), .A2(n13635), .A3(n4689), .ZN(n4688) );
  NAND3_X2 U8353 ( .A1(n73), .A2(n20727), .A3(n3252), .ZN(n22845) );
  OR2_X1 U8381 ( .A1(n20430), .A2(n28894), .ZN(n20622) );
  OR2_X1 U8404 ( .A1(n4346), .A2(n1931), .ZN(n10896) );
  INV_X1 U8445 ( .A(n12593), .ZN(n5069) );
  NAND2_X1 U8451 ( .A1(n29009), .A2(n2587), .ZN(n12593) );
  NAND2_X1 U8470 ( .A1(n28895), .A2(n5674), .ZN(n5673) );
  OAI21_X1 U8471 ( .B1(n6147), .B2(n9016), .A(n5676), .ZN(n28895) );
  INV_X1 U8473 ( .A(n12346), .ZN(n10649) );
  NOR2_X1 U8488 ( .A1(n21273), .A2(n6934), .ZN(n21274) );
  AND2_X1 U8491 ( .A1(n21373), .A2(n21372), .ZN(n6934) );
  NAND2_X1 U8497 ( .A1(n3776), .A2(n10722), .ZN(n11486) );
  NOR2_X1 U8498 ( .A1(n28767), .A2(n28897), .ZN(n28896) );
  OAI21_X1 U8501 ( .B1(n20359), .B2(n20238), .A(n20243), .ZN(n28898) );
  NAND3_X1 U8529 ( .A1(n9039), .A2(n9243), .A3(n9248), .ZN(n8694) );
  NAND2_X1 U8578 ( .A1(n14355), .A2(n28899), .ZN(n6873) );
  NAND2_X1 U8587 ( .A1(n28902), .A2(n28900), .ZN(n18084) );
  INV_X1 U8613 ( .A(n374), .ZN(n28901) );
  NAND2_X1 U8617 ( .A1(n18082), .A2(n374), .ZN(n28902) );
  XNOR2_X1 U8626 ( .A(n28903), .B(n3662), .ZN(Ciphertext[18]) );
  AOI22_X1 U8628 ( .A1(n26961), .A2(n27410), .B1(n28607), .B2(n26962), .ZN(
        n28903) );
  NAND2_X1 U8643 ( .A1(n2518), .A2(n11085), .ZN(n10165) );
  NAND2_X1 U8648 ( .A1(n23929), .A2(n24588), .ZN(n1283) );
  OR2_X2 U8649 ( .A1(n28245), .A2(n14925), .ZN(n16323) );
  NOR2_X2 U8657 ( .A1(n23670), .A2(n23671), .ZN(n24812) );
  NAND3_X1 U8665 ( .A1(n13255), .A2(n13578), .A3(n13254), .ZN(n6812) );
  NAND3_X2 U8675 ( .A1(n3484), .A2(n29176), .A3(n28904), .ZN(n18034) );
  NAND2_X1 U8679 ( .A1(n28906), .A2(n28905), .ZN(n28904) );
  INV_X1 U8717 ( .A(n17301), .ZN(n28905) );
  INV_X1 U8719 ( .A(n17300), .ZN(n28906) );
  NAND3_X1 U8720 ( .A1(n29174), .A2(n980), .A3(n24076), .ZN(n25398) );
  NAND2_X1 U8732 ( .A1(n28909), .A2(n28907), .ZN(n25243) );
  OR2_X1 U8742 ( .A1(n27395), .A2(n28908), .ZN(n28907) );
  INV_X1 U8749 ( .A(n26191), .ZN(n28908) );
  NAND2_X1 U8765 ( .A1(n27395), .A2(n27393), .ZN(n28909) );
  NAND2_X1 U8778 ( .A1(n28910), .A2(n10448), .ZN(n2272) );
  NAND2_X1 U8793 ( .A1(n6542), .A2(n10110), .ZN(n28910) );
  XNOR2_X2 U8806 ( .A(n16599), .B(n180), .ZN(n17518) );
  NAND2_X1 U8840 ( .A1(n9039), .A2(n28911), .ZN(n8697) );
  NAND2_X1 U8849 ( .A1(n29177), .A2(n17434), .ZN(n28912) );
  XNOR2_X1 U8894 ( .A(n22079), .B(n28914), .ZN(n28622) );
  NAND3_X1 U8928 ( .A1(n6586), .A2(n6585), .A3(n6584), .ZN(n6741) );
  XNOR2_X1 U8934 ( .A(n10183), .B(n10232), .ZN(n9606) );
  NAND2_X1 U8940 ( .A1(n28915), .A2(n20951), .ZN(n20957) );
  NAND2_X1 U8969 ( .A1(n21931), .A2(n28916), .ZN(n28915) );
  OAI21_X2 U8983 ( .B1(n11382), .B2(n11381), .A(n28917), .ZN(n13297) );
  NAND2_X1 U9032 ( .A1(n24539), .A2(n24540), .ZN(n24548) );
  OAI21_X1 U9039 ( .B1(n26209), .B2(n283), .A(n25665), .ZN(n25632) );
  OAI211_X1 U9101 ( .C1(n24162), .C2(n24802), .A(n24503), .B(n28918), .ZN(
        n24165) );
  NAND2_X1 U9169 ( .A1(n24162), .A2(n28919), .ZN(n28918) );
  INV_X1 U9216 ( .A(n24806), .ZN(n28919) );
  NAND2_X1 U9218 ( .A1(n24681), .A2(n24391), .ZN(n28262) );
  OAI211_X2 U9261 ( .C1(n24381), .C2(n24380), .A(n2905), .B(n2906), .ZN(n25352) );
  AOI21_X1 U9265 ( .B1(n4826), .B2(n28920), .A(n7641), .ZN(n4825) );
  NAND2_X1 U9279 ( .A1(n7985), .A2(n7642), .ZN(n28920) );
  OR2_X2 U9294 ( .A1(n1056), .A2(n8461), .ZN(n9930) );
  AND2_X1 U9319 ( .A1(n13653), .A2(n14327), .ZN(n13799) );
  INV_X1 U9324 ( .A(n8767), .ZN(n28921) );
  NAND2_X1 U9327 ( .A1(n28921), .A2(n9425), .ZN(n8769) );
  AND3_X2 U9329 ( .A1(n28924), .A2(n28923), .A3(n28922), .ZN(n24484) );
  NAND2_X1 U9336 ( .A1(n6941), .A2(n23458), .ZN(n28922) );
  NAND2_X1 U9341 ( .A1(n23117), .A2(n23460), .ZN(n28923) );
  INV_X1 U9363 ( .A(n11220), .ZN(n28929) );
  NOR2_X1 U9390 ( .A1(n10280), .A2(n28931), .ZN(n28930) );
  AND2_X1 U9394 ( .A1(n10269), .A2(n11220), .ZN(n28931) );
  AND2_X2 U9398 ( .A1(n1316), .A2(n1317), .ZN(n12813) );
  OR2_X1 U9402 ( .A1(n422), .A2(n16809), .ZN(n29195) );
  NAND2_X1 U9420 ( .A1(n2922), .A2(n28252), .ZN(n20434) );
  NAND2_X1 U9447 ( .A1(n17688), .A2(n1708), .ZN(n853) );
  NAND2_X1 U9467 ( .A1(n21579), .A2(n21578), .ZN(n5139) );
  NAND2_X1 U9557 ( .A1(n8049), .A2(n8131), .ZN(n28933) );
  NAND2_X1 U9586 ( .A1(n7556), .A2(n7127), .ZN(n28934) );
  NAND3_X2 U9592 ( .A1(n28935), .A2(n3885), .A3(n3884), .ZN(n18215) );
  NAND2_X1 U9618 ( .A1(n2559), .A2(n2560), .ZN(n28935) );
  NAND2_X1 U9629 ( .A1(n21392), .A2(n21632), .ZN(n21634) );
  NAND3_X1 U9652 ( .A1(n4754), .A2(n23119), .A3(n24479), .ZN(n23120) );
  NAND3_X1 U9682 ( .A1(n14281), .A2(n14082), .A3(n14081), .ZN(n14088) );
  NAND3_X2 U9685 ( .A1(n17245), .A2(n17244), .A3(n17243), .ZN(n2855) );
  OAI22_X1 U9687 ( .A1(n15337), .A2(n15338), .B1(n15339), .B2(n5777), .ZN(
        n15340) );
  NAND2_X1 U9688 ( .A1(n15233), .A2(n15333), .ZN(n15337) );
  AND4_X2 U9731 ( .A1(n6528), .A2(n21045), .A3(n21044), .A4(n21043), .ZN(
        n22488) );
  NAND2_X1 U9732 ( .A1(n1715), .A2(n1714), .ZN(n1207) );
  NAND2_X1 U9734 ( .A1(n4304), .A2(n9208), .ZN(n28938) );
  NOR2_X1 U9754 ( .A1(n24699), .A2(n28939), .ZN(n711) );
  INV_X1 U9756 ( .A(n24771), .ZN(n28939) );
  NAND2_X1 U9793 ( .A1(n24768), .A2(n24697), .ZN(n24771) );
  NAND3_X1 U9828 ( .A1(n22255), .A2(n22256), .A3(n23645), .ZN(n22257) );
  NAND2_X1 U9851 ( .A1(n7640), .A2(n7980), .ZN(n7647) );
  NAND2_X1 U9857 ( .A1(n7644), .A2(n7981), .ZN(n7640) );
  NAND2_X1 U9878 ( .A1(n29005), .A2(n14338), .ZN(n14339) );
  NAND2_X1 U9912 ( .A1(n2948), .A2(n10730), .ZN(n2947) );
  NAND2_X1 U9943 ( .A1(n2929), .A2(n3033), .ZN(n26462) );
  NAND3_X1 U9944 ( .A1(n24655), .A2(n3061), .A3(n24651), .ZN(n6223) );
  NAND3_X2 U9947 ( .A1(n28940), .A2(n28941), .A3(n6213), .ZN(n21728) );
  NAND3_X1 U9953 ( .A1(n21571), .A2(n20754), .A3(n21457), .ZN(n28940) );
  XNOR2_X2 U9954 ( .A(n7049), .B(Key[159]), .ZN(n1938) );
  OAI211_X1 U9984 ( .C1(n5234), .C2(n18391), .A(n18390), .B(n18389), .ZN(
        n18392) );
  NAND2_X1 U10004 ( .A1(n17732), .A2(n5234), .ZN(n18390) );
  NAND2_X1 U10008 ( .A1(n3844), .A2(n3846), .ZN(n16192) );
  NAND2_X1 U10009 ( .A1(n3845), .A2(n13865), .ZN(n3844) );
  AOI21_X2 U10061 ( .B1(n711), .B2(n28942), .A(n24701), .ZN(n25927) );
  NAND2_X1 U10090 ( .A1(n3054), .A2(n24700), .ZN(n28942) );
  NAND2_X1 U10120 ( .A1(n20867), .A2(n21497), .ZN(n28943) );
  AOI21_X1 U10132 ( .B1(n3442), .B2(n3441), .A(n28944), .ZN(n11247) );
  OAI211_X1 U10164 ( .C1(n16337), .C2(n2158), .A(n2157), .B(n28945), .ZN(n2155) );
  NAND2_X1 U10178 ( .A1(n16337), .A2(n538), .ZN(n28945) );
  NAND2_X1 U10201 ( .A1(n28947), .A2(n28946), .ZN(n17011) );
  NAND3_X1 U10213 ( .A1(n29088), .A2(n5891), .A3(n17428), .ZN(n28946) );
  NAND2_X1 U10246 ( .A1(n17006), .A2(n28792), .ZN(n28947) );
  NOR2_X1 U10247 ( .A1(n17942), .A2(n17762), .ZN(n1442) );
  NAND2_X1 U10294 ( .A1(n23518), .A2(n23519), .ZN(n23520) );
  NAND2_X1 U10331 ( .A1(n26801), .A2(n28823), .ZN(n28948) );
  NAND3_X1 U10342 ( .A1(n10408), .A2(n2891), .A3(n2892), .ZN(n29273) );
  OR2_X1 U10407 ( .A1(n23360), .A2(n23676), .ZN(n2888) );
  NAND2_X1 U10418 ( .A1(n2909), .A2(n21672), .ZN(n3903) );
  XNOR2_X1 U10474 ( .A(n26073), .B(n2350), .ZN(n25367) );
  NOR2_X1 U10489 ( .A1(n7534), .A2(n8014), .ZN(n3031) );
  NAND2_X1 U10490 ( .A1(n8013), .A2(n7743), .ZN(n7534) );
  INV_X1 U10518 ( .A(n27101), .ZN(n3542) );
  AND2_X1 U10519 ( .A1(n28949), .A2(n27101), .ZN(n3236) );
  NOR2_X2 U10521 ( .A1(n26854), .A2(n27839), .ZN(n27101) );
  INV_X1 U10533 ( .A(n27100), .ZN(n28949) );
  NAND2_X1 U10541 ( .A1(n14295), .A2(n13306), .ZN(n13309) );
  OAI211_X1 U10542 ( .C1(n23431), .C2(n408), .A(n23430), .B(n28951), .ZN(n1073) );
  NAND2_X1 U10552 ( .A1(n4178), .A2(n23431), .ZN(n28951) );
  NAND3_X1 U10560 ( .A1(n13618), .A2(n13617), .A3(n13616), .ZN(n28953) );
  NAND2_X1 U10568 ( .A1(n10990), .A2(n10995), .ZN(n10693) );
  NAND2_X1 U10591 ( .A1(n24634), .A2(n24635), .ZN(n24243) );
  NOR2_X1 U10637 ( .A1(n23792), .A2(n23790), .ZN(n28954) );
  INV_X1 U10646 ( .A(n23495), .ZN(n28955) );
  NAND2_X1 U10662 ( .A1(n1121), .A2(n17027), .ZN(n1120) );
  NAND2_X1 U10670 ( .A1(n5219), .A2(n884), .ZN(n24612) );
  NAND2_X1 U10677 ( .A1(n17930), .A2(n1863), .ZN(n19508) );
  OR3_X1 U10685 ( .A1(n1910), .A2(n8077), .A3(n8058), .ZN(n7807) );
  XNOR2_X1 U10700 ( .A(n28956), .B(n22619), .ZN(n6017) );
  NAND3_X1 U10702 ( .A1(n2665), .A2(n6015), .A3(n2667), .ZN(n28956) );
  OAI211_X2 U10703 ( .C1(n23299), .C2(n23300), .A(n5712), .B(n5713), .ZN(
        n24404) );
  NOR2_X1 U10732 ( .A1(n5181), .A2(n20149), .ZN(n20741) );
  NAND3_X1 U10768 ( .A1(n21561), .A2(n21465), .A3(n21464), .ZN(n28958) );
  INV_X1 U10797 ( .A(n10345), .ZN(n9612) );
  NAND2_X1 U10800 ( .A1(n203), .A2(n6688), .ZN(n10345) );
  NAND2_X1 U10876 ( .A1(n28960), .A2(n16906), .ZN(n1721) );
  NAND2_X1 U10882 ( .A1(n17228), .A2(n1723), .ZN(n28960) );
  OAI211_X1 U10909 ( .C1(n11907), .C2(n12359), .A(n919), .B(n12363), .ZN(
        n28962) );
  NAND3_X1 U10954 ( .A1(n28963), .A2(n23640), .A3(n22996), .ZN(n2622) );
  OAI211_X1 U10966 ( .C1(n11262), .C2(n29122), .A(n11265), .B(n6631), .ZN(
        n12293) );
  XNOR2_X1 U10967 ( .A(n19254), .B(n28964), .ZN(n4307) );
  XNOR2_X1 U10979 ( .A(n19383), .B(n28965), .ZN(n28964) );
  INV_X1 U10982 ( .A(n18737), .ZN(n28965) );
  NOR2_X1 U11027 ( .A1(n28966), .A2(n29026), .ZN(n23965) );
  INV_X1 U11042 ( .A(n24583), .ZN(n28966) );
  OAI21_X2 U11043 ( .B1(n21978), .B2(n23607), .A(n21977), .ZN(n24583) );
  OAI22_X1 U11054 ( .A1(n27266), .A2(n27596), .B1(n26346), .B2(n28967), .ZN(
        n27269) );
  NAND2_X1 U11084 ( .A1(n26372), .A2(n28970), .ZN(n28969) );
  INV_X1 U11107 ( .A(n26266), .ZN(n28970) );
  INV_X1 U11121 ( .A(n463), .ZN(n28971) );
  NAND3_X1 U11161 ( .A1(n28971), .A2(n24775), .A3(n24779), .ZN(n3836) );
  NAND2_X1 U11204 ( .A1(n3564), .A2(n4778), .ZN(n15184) );
  NAND3_X1 U11214 ( .A1(n3432), .A2(n3502), .A3(n23734), .ZN(n2481) );
  AOI22_X2 U11232 ( .A1(n17521), .A2(n17520), .B1(n17519), .B2(n796), .ZN(
        n18227) );
  XNOR2_X2 U11253 ( .A(n2257), .B(n19690), .ZN(n20440) );
  OAI21_X2 U11262 ( .B1(n4586), .B2(n13464), .A(n28972), .ZN(n13789) );
  NAND2_X1 U11268 ( .A1(n14148), .A2(n14376), .ZN(n28972) );
  OAI21_X1 U11286 ( .B1(n4854), .B2(n18033), .A(n28973), .ZN(n17827) );
  NAND2_X1 U11300 ( .A1(n4959), .A2(n28974), .ZN(n20861) );
  NAND3_X1 U11376 ( .A1(n20858), .A2(n21157), .A3(n21156), .ZN(n28974) );
  NAND3_X1 U11454 ( .A1(n27664), .A2(n28347), .A3(n27661), .ZN(n28373) );
  OAI21_X1 U11462 ( .B1(n20572), .B2(n20571), .A(n20570), .ZN(n20715) );
  NAND3_X1 U11474 ( .A1(n29557), .A2(n28975), .A3(n27225), .ZN(n4526) );
  INV_X1 U11477 ( .A(n4528), .ZN(n28975) );
  NAND2_X1 U11516 ( .A1(n11168), .A2(n10820), .ZN(n4107) );
  XNOR2_X1 U11517 ( .A(n28977), .B(n25322), .ZN(n24608) );
  NAND2_X1 U11560 ( .A1(n947), .A2(n946), .ZN(n28977) );
  OR2_X1 U11561 ( .A1(n21092), .A2(n18919), .ZN(n19870) );
  NAND3_X1 U11579 ( .A1(n14), .A2(n21158), .A3(n21157), .ZN(n13) );
  NAND3_X1 U11583 ( .A1(n29238), .A2(n2330), .A3(n28819), .ZN(n28978) );
  NOR2_X2 U11601 ( .A1(n18176), .A2(n28981), .ZN(n18880) );
  AOI21_X1 U11634 ( .B1(n7650), .B2(n7651), .A(n7649), .ZN(n7654) );
  NAND2_X1 U11656 ( .A1(n437), .A2(n29082), .ZN(n7650) );
  NAND3_X1 U11767 ( .A1(n8299), .A2(n8298), .A3(n8297), .ZN(n2405) );
  NAND2_X1 U11783 ( .A1(n1018), .A2(n1017), .ZN(n4005) );
  NAND2_X1 U11820 ( .A1(n14254), .A2(n29312), .ZN(n4376) );
  NAND3_X1 U11876 ( .A1(n2450), .A2(n17358), .A3(n2449), .ZN(n1752) );
  NAND3_X1 U11963 ( .A1(n23546), .A2(n4773), .A3(n4772), .ZN(n28983) );
  NAND2_X1 U11966 ( .A1(n28985), .A2(n28984), .ZN(n14610) );
  NAND2_X1 U12008 ( .A1(n14306), .A2(n14429), .ZN(n28984) );
  NAND2_X1 U12037 ( .A1(n28987), .A2(n28986), .ZN(n28985) );
  NAND2_X1 U12053 ( .A1(n14305), .A2(n4837), .ZN(n28987) );
  NAND2_X1 U12060 ( .A1(n9437), .A2(n28988), .ZN(n10045) );
  NAND2_X1 U12111 ( .A1(n28990), .A2(n28989), .ZN(n28988) );
  NAND2_X1 U12113 ( .A1(n9435), .A2(n9434), .ZN(n28990) );
  NAND2_X1 U12121 ( .A1(n28185), .A2(n28991), .ZN(n21193) );
  NAND2_X1 U12123 ( .A1(n21356), .A2(n28126), .ZN(n28992) );
  XNOR2_X1 U12151 ( .A(n29519), .B(n3462), .ZN(n22412) );
  NAND3_X1 U12201 ( .A1(n28994), .A2(n3629), .A3(n28993), .ZN(n18312) );
  NAND2_X1 U12213 ( .A1(n5587), .A2(n29373), .ZN(n28994) );
  NAND2_X1 U12220 ( .A1(n28198), .A2(n28995), .ZN(n4181) );
  NOR2_X1 U12221 ( .A1(n14845), .A2(n28996), .ZN(n28995) );
  INV_X1 U12227 ( .A(n15285), .ZN(n28996) );
  OAI21_X1 U12231 ( .B1(n7709), .B2(n7737), .A(n28998), .ZN(n7713) );
  NAND2_X1 U12309 ( .A1(n16859), .A2(n28999), .ZN(n17802) );
  NAND2_X1 U12319 ( .A1(n569), .A2(n12305), .ZN(n1238) );
  MUX2_X1 U12349 ( .A(n9095), .B(n8665), .S(n8490), .Z(n8668) );
  AOI21_X1 U12366 ( .B1(n10920), .B2(n10718), .A(n29001), .ZN(n10050) );
  NAND2_X1 U12390 ( .A1(n10031), .A2(n3862), .ZN(n29001) );
  NAND2_X1 U12426 ( .A1(n24248), .A2(n24155), .ZN(n24246) );
  NAND2_X1 U12436 ( .A1(n24524), .A2(n3061), .ZN(n29003) );
  NAND3_X1 U12439 ( .A1(n29004), .A2(n23921), .A3(n4783), .ZN(n24858) );
  NAND2_X1 U12441 ( .A1(n3295), .A2(n24582), .ZN(n29004) );
  NAND3_X1 U12465 ( .A1(n5190), .A2(n5189), .A3(n15311), .ZN(n29005) );
  OAI211_X2 U12471 ( .C1(n21381), .C2(n21380), .A(n4265), .B(n29006), .ZN(
        n22625) );
  NAND2_X1 U12474 ( .A1(n21380), .A2(n21253), .ZN(n29006) );
  NAND2_X1 U12484 ( .A1(n15939), .A2(n18061), .ZN(n29007) );
  NAND2_X1 U12504 ( .A1(n29008), .A2(n16874), .ZN(n4291) );
  NAND2_X1 U12510 ( .A1(n1262), .A2(n29512), .ZN(n21726) );
  AND2_X2 U12512 ( .A1(n2396), .A2(n3619), .ZN(n22387) );
  AOI22_X1 U12514 ( .A1(n12429), .A2(n12428), .B1(n10586), .B2(n10587), .ZN(
        n29009) );
  NAND2_X1 U12524 ( .A1(n1886), .A2(n15084), .ZN(n29010) );
  NAND2_X1 U12546 ( .A1(n15693), .A2(n15692), .ZN(n29012) );
  NAND2_X1 U12599 ( .A1(n21019), .A2(n22023), .ZN(n22025) );
  OAI21_X1 U12618 ( .B1(n24055), .B2(n24054), .A(n29013), .ZN(n24056) );
  OAI21_X1 U12665 ( .B1(n29015), .B2(n29545), .A(n29014), .ZN(n24026) );
  NAND2_X1 U12705 ( .A1(n24022), .A2(n462), .ZN(n29014) );
  BUF_X1 U12762 ( .A(n26459), .Z(n28476) );
  AOI22_X2 U12793 ( .A1(n23191), .A2(n23757), .B1(n5741), .B2(n23190), .ZN(
        n24635) );
  XNOR2_X1 U12866 ( .A(n19326), .B(n19325), .ZN(n20625) );
  XNOR2_X1 U12902 ( .A(n25841), .B(n25842), .ZN(n27120) );
  INV_X1 U12921 ( .A(n27092), .ZN(n27920) );
  OAI211_X1 U12938 ( .C1(n28550), .C2(n24747), .A(n24267), .B(n24266), .ZN(
        n29017) );
  NOR2_X2 U12949 ( .A1(n20657), .A2(n20656), .ZN(n28550) );
  BUF_X1 U12960 ( .A(n23432), .Z(n29018) );
  XNOR2_X1 U12982 ( .A(n3983), .B(n22660), .ZN(n23432) );
  AND2_X1 U12998 ( .A1(n21415), .A2(n29019), .ZN(n21050) );
  NAND2_X1 U13011 ( .A1(n21413), .A2(n20663), .ZN(n29019) );
  MUX2_X1 U13013 ( .A(n23914), .B(n23913), .S(n24667), .Z(n23915) );
  XNOR2_X1 U13046 ( .A(n22530), .B(n22529), .ZN(n23297) );
  AND3_X1 U13069 ( .A1(n3177), .A2(n26618), .A3(n26619), .ZN(n29021) );
  NAND3_X1 U13086 ( .A1(n3177), .A2(n26618), .A3(n26619), .ZN(n27979) );
  OR2_X1 U13125 ( .A1(n29104), .A2(n20041), .ZN(n20089) );
  NAND2_X1 U13232 ( .A1(n6492), .A2(n6026), .ZN(n29022) );
  OR2_X1 U13233 ( .A1(n24496), .A2(n5004), .ZN(n24207) );
  OAI22_X1 U13237 ( .A1(n6857), .A2(n5221), .B1(n27054), .B2(n1971), .ZN(
        n28025) );
  INV_X1 U13252 ( .A(n5234), .ZN(n29023) );
  INV_X1 U13288 ( .A(n5234), .ZN(n29024) );
  BUF_X1 U13296 ( .A(n26746), .Z(n28563) );
  XNOR2_X2 U13317 ( .A(n26027), .B(n26026), .ZN(n26865) );
  OAI21_X1 U13322 ( .B1(n22129), .B2(n28474), .A(n22128), .ZN(n29025) );
  OR2_X1 U13395 ( .A1(n26308), .A2(n26307), .ZN(n29027) );
  OAI21_X1 U13396 ( .B1(n22129), .B2(n28474), .A(n22128), .ZN(n24577) );
  XOR2_X1 U13409 ( .A(n24276), .B(n24275), .Z(n29028) );
  OR2_X1 U13491 ( .A1(n29075), .A2(n29500), .ZN(n27066) );
  AND2_X1 U13507 ( .A1(n5114), .A2(n5112), .ZN(n29029) );
  OR3_X1 U13516 ( .A1(n27074), .A2(n26992), .A3(n27076), .ZN(n29030) );
  AND2_X1 U13538 ( .A1(n3254), .A2(n25556), .ZN(n29031) );
  MUX2_X1 U13543 ( .A(n25462), .B(n25461), .S(n5760), .Z(n25472) );
  AND3_X1 U13545 ( .A1(n26669), .A2(n26531), .A3(n27417), .ZN(n26535) );
  MUX2_X1 U13546 ( .A(n29560), .B(n28548), .S(n26210), .Z(n26719) );
  AND2_X1 U13577 ( .A1(n25600), .A2(n25599), .ZN(n29032) );
  AND2_X1 U13582 ( .A1(n25600), .A2(n25599), .ZN(n28038) );
  BUF_X1 U13583 ( .A(n26028), .Z(n28534) );
  OAI211_X1 U13599 ( .C1(n24894), .C2(n23984), .A(n29269), .B(n29268), .ZN(
        n26028) );
  OAI21_X2 U13678 ( .B1(n26219), .B2(n26716), .A(n26218), .ZN(n28063) );
  AOI21_X2 U13708 ( .B1(n26269), .B2(n26775), .A(n26268), .ZN(n27594) );
  BUF_X1 U13709 ( .A(n27052), .Z(n28446) );
  NAND2_X1 U13712 ( .A1(n23813), .A2(n1239), .ZN(n29033) );
  OR2_X1 U13740 ( .A1(n17257), .A2(n17256), .ZN(n29034) );
  AND2_X1 U13748 ( .A1(n17972), .A2(n17973), .ZN(n29035) );
  NOR2_X1 U13753 ( .A1(n18034), .A2(n18033), .ZN(n18164) );
  OR2_X1 U13756 ( .A1(n17743), .A2(n18034), .ZN(n29289) );
  XOR2_X1 U13764 ( .A(n21979), .B(n22880), .Z(n21986) );
  OAI211_X2 U13766 ( .C1(n20846), .C2(n20841), .A(n20845), .B(n3555), .ZN(
        n22703) );
  OAI211_X1 U13781 ( .C1(n220), .C2(n24464), .A(n24462), .B(n24463), .ZN(
        n29053) );
  OAI211_X1 U13796 ( .C1(n220), .C2(n24464), .A(n24462), .B(n24463), .ZN(
        n25889) );
  XNOR2_X1 U13810 ( .A(n12767), .B(n12766), .ZN(n29036) );
  XNOR2_X1 U13876 ( .A(n12767), .B(n12766), .ZN(n29037) );
  OAI211_X1 U13881 ( .C1(n18240), .C2(n17290), .A(n17289), .B(n17288), .ZN(
        n29038) );
  OAI211_X1 U13882 ( .C1(n18240), .C2(n17290), .A(n17289), .B(n17288), .ZN(
        n18935) );
  AOI22_X1 U13923 ( .A1(n24407), .A2(n3797), .B1(n24086), .B2(n24085), .ZN(
        n25913) );
  XNOR2_X1 U13965 ( .A(n19039), .B(n19381), .ZN(n6569) );
  INV_X1 U13976 ( .A(n500), .ZN(n29040) );
  XNOR2_X1 U14001 ( .A(n18637), .B(n18636), .ZN(n29041) );
  XOR2_X1 U14040 ( .A(n22907), .B(n22906), .Z(n29042) );
  OR2_X1 U14063 ( .A1(n20862), .A2(n29236), .ZN(n4543) );
  XNOR2_X1 U14090 ( .A(n21986), .B(n21985), .ZN(n23735) );
  OAI211_X1 U14100 ( .C1(n23035), .C2(n23034), .A(n4935), .B(n4934), .ZN(
        n24704) );
  BUF_X1 U14111 ( .A(n26466), .Z(n280) );
  NAND2_X1 U14113 ( .A1(n2484), .A2(n16832), .ZN(n29044) );
  NAND2_X1 U14120 ( .A1(n2484), .A2(n16832), .ZN(n19561) );
  XOR2_X1 U14124 ( .A(n18991), .B(n18992), .Z(n18997) );
  XOR2_X1 U14125 ( .A(n19245), .B(n19669), .Z(n17597) );
  XNOR2_X1 U14135 ( .A(n15598), .B(n15599), .ZN(n29045) );
  INV_X1 U14151 ( .A(n22053), .ZN(n22731) );
  NOR2_X2 U14181 ( .A1(n1008), .A2(n26324), .ZN(n27795) );
  NOR2_X1 U14262 ( .A1(n24774), .A2(n24773), .ZN(n29047) );
  AND2_X1 U14285 ( .A1(n446), .A2(n27377), .ZN(n29219) );
  XNOR2_X1 U14361 ( .A(n26064), .B(n26063), .ZN(n29048) );
  NOR2_X1 U14391 ( .A1(n27902), .A2(n26848), .ZN(n26852) );
  BUF_X1 U14417 ( .A(n26579), .Z(n28477) );
  AND2_X1 U14496 ( .A1(n26926), .A2(n26579), .ZN(n26929) );
  XOR2_X1 U14502 ( .A(n10368), .B(n9703), .Z(n9708) );
  AND2_X1 U14503 ( .A1(n24095), .A2(n4532), .ZN(n29051) );
  AND2_X1 U14522 ( .A1(n4532), .A2(n24095), .ZN(n23874) );
  AND2_X1 U14544 ( .A1(n28669), .A2(n5422), .ZN(n29052) );
  AND2_X1 U14581 ( .A1(n28669), .A2(n5422), .ZN(n27352) );
  XNOR2_X1 U14721 ( .A(n24787), .B(n24786), .ZN(n29054) );
  OR2_X1 U14741 ( .A1(n26200), .A2(n26235), .ZN(n29055) );
  BUF_X1 U14788 ( .A(n29052), .Z(n27351) );
  AND4_X1 U14810 ( .A1(n679), .A2(n16893), .A3(n16892), .A4(n16894), .ZN(
        n29057) );
  OR2_X1 U14862 ( .A1(n17113), .A2(n29539), .ZN(n3099) );
  XNOR2_X1 U14870 ( .A(n28311), .B(n1987), .ZN(n29059) );
  XNOR2_X1 U14881 ( .A(n28311), .B(n1987), .ZN(n14008) );
  XNOR2_X1 U14935 ( .A(n26037), .B(n26036), .ZN(n29060) );
  XNOR2_X1 U15010 ( .A(n22565), .B(n22564), .ZN(n22566) );
  AOI22_X1 U15060 ( .A1(n26611), .A2(n28394), .B1(n295), .B2(n26610), .ZN(
        n5651) );
  XNOR2_X1 U15074 ( .A(n25483), .B(n25482), .ZN(n29062) );
  OR2_X1 U15084 ( .A1(n26626), .A2(n5685), .ZN(n29063) );
  XNOR2_X1 U15100 ( .A(n25483), .B(n25482), .ZN(n27050) );
  OAI21_X1 U15101 ( .B1(n11359), .B2(n12401), .A(n11358), .ZN(n29064) );
  INV_X1 U15114 ( .A(n2656), .ZN(n29065) );
  OAI21_X1 U15150 ( .B1(n11359), .B2(n12401), .A(n11358), .ZN(n12746) );
  AOI21_X1 U15157 ( .B1(n16968), .B2(n6130), .A(n6126), .ZN(n17889) );
  XNOR2_X1 U15167 ( .A(n18866), .B(n18865), .ZN(n29066) );
  OAI21_X1 U15169 ( .B1(n24414), .B2(n4136), .A(n2261), .ZN(n29067) );
  XNOR2_X1 U15174 ( .A(n18866), .B(n18865), .ZN(n20161) );
  OAI21_X1 U15175 ( .B1(n24414), .B2(n4136), .A(n2261), .ZN(n25550) );
  NOR2_X1 U15191 ( .A1(n25797), .A2(n25800), .ZN(n29069) );
  NOR2_X1 U15216 ( .A1(n25797), .A2(n25800), .ZN(n25729) );
  XNOR2_X1 U15227 ( .A(n25163), .B(n25164), .ZN(n29071) );
  XNOR2_X1 U15380 ( .A(n25163), .B(n25164), .ZN(n26952) );
  BUF_X1 U15381 ( .A(n17296), .Z(n29072) );
  AOI21_X1 U15447 ( .B1(n24034), .B2(n24033), .A(n24032), .ZN(n29073) );
  AOI21_X1 U15458 ( .B1(n24034), .B2(n24033), .A(n24032), .ZN(n25886) );
  OAI21_X1 U15520 ( .B1(n3671), .B2(n24513), .A(n3618), .ZN(n29193) );
  XNOR2_X1 U15553 ( .A(n22237), .B(n22236), .ZN(n29074) );
  XNOR2_X1 U15554 ( .A(n22237), .B(n22236), .ZN(n23642) );
  XOR2_X1 U15693 ( .A(n25700), .B(n25699), .Z(n29075) );
  XOR2_X1 U15844 ( .A(n25700), .B(n25699), .Z(n29076) );
  CLKBUF_X1 U15907 ( .A(n25344), .Z(n26737) );
  XNOR2_X1 U15930 ( .A(n9346), .B(n9347), .ZN(n29077) );
  XNOR2_X1 U15938 ( .A(n9346), .B(n9347), .ZN(n29078) );
  BUF_X1 U16008 ( .A(n22783), .Z(n29079) );
  XNOR2_X1 U16039 ( .A(n7058), .B(Key[167]), .ZN(n29081) );
  XNOR2_X1 U16071 ( .A(n7058), .B(Key[167]), .ZN(n29082) );
  XNOR2_X1 U16216 ( .A(n1257), .B(n1258), .ZN(n29083) );
  XNOR2_X1 U16217 ( .A(n7058), .B(Key[167]), .ZN(n7876) );
  XNOR2_X1 U16250 ( .A(n1257), .B(n1258), .ZN(n16811) );
  NAND3_X1 U16251 ( .A1(n15034), .A2(n15035), .A3(n15033), .ZN(n29084) );
  NAND3_X1 U16340 ( .A1(n15034), .A2(n15035), .A3(n15033), .ZN(n15966) );
  NAND2_X1 U16360 ( .A1(n26395), .A2(n56), .ZN(n29085) );
  NAND2_X1 U16375 ( .A1(n26395), .A2(n56), .ZN(n27572) );
  XOR2_X1 U16437 ( .A(n16049), .B(n16048), .Z(n29086) );
  XOR2_X1 U16444 ( .A(n22053), .B(n22052), .Z(n29087) );
  INV_X1 U16445 ( .A(n6013), .ZN(n29088) );
  XOR2_X1 U16688 ( .A(n13477), .B(n13476), .Z(n29089) );
  NAND3_X2 U16689 ( .A1(n2051), .A2(n26233), .A3(n26232), .ZN(n28067) );
  NAND2_X1 U16785 ( .A1(n27164), .A2(n5993), .ZN(n29090) );
  NAND2_X1 U16824 ( .A1(n27164), .A2(n5993), .ZN(n29091) );
  NAND2_X1 U16832 ( .A1(n27164), .A2(n5993), .ZN(n27673) );
  OR2_X1 U16883 ( .A1(n26635), .A2(n26634), .ZN(n29092) );
  NOR2_X2 U16901 ( .A1(n26578), .A2(n26577), .ZN(n29093) );
  NOR2_X1 U16957 ( .A1(n26578), .A2(n26577), .ZN(n27494) );
  MUX2_X1 U16960 ( .A(n21027), .B(n21026), .S(n23016), .Z(n21060) );
  NOR2_X1 U17016 ( .A1(n146), .A2(n23904), .ZN(n29094) );
  NOR2_X1 U17032 ( .A1(n146), .A2(n23904), .ZN(n25246) );
  OAI21_X1 U17036 ( .B1(n28617), .B2(n8262), .A(n8261), .ZN(n29096) );
  OAI21_X1 U17070 ( .B1(n28617), .B2(n8262), .A(n8261), .ZN(n8954) );
  XNOR2_X1 U17072 ( .A(n11546), .B(n11545), .ZN(n14171) );
  XNOR2_X1 U17114 ( .A(n15883), .B(n15882), .ZN(n29098) );
  XNOR2_X1 U17127 ( .A(n25439), .B(n25438), .ZN(n29099) );
  XNOR2_X1 U17150 ( .A(n25439), .B(n25438), .ZN(n29100) );
  BUF_X1 U17222 ( .A(n21696), .Z(n29101) );
  XNOR2_X1 U17265 ( .A(n22622), .B(n22623), .ZN(n29102) );
  XNOR2_X1 U17270 ( .A(n22622), .B(n22623), .ZN(n23806) );
  NOR2_X1 U17318 ( .A1(n24733), .A2(n3725), .ZN(n29103) );
  NOR2_X1 U17376 ( .A1(n24733), .A2(n3725), .ZN(n25531) );
  XNOR2_X1 U17383 ( .A(n18747), .B(n18748), .ZN(n29104) );
  XNOR2_X1 U17384 ( .A(n13182), .B(n13183), .ZN(n29107) );
  XNOR2_X1 U17393 ( .A(n7008), .B(Key[71]), .ZN(n7011) );
  XNOR2_X1 U17406 ( .A(n13182), .B(n13183), .ZN(n13920) );
  XNOR2_X1 U17457 ( .A(n24937), .B(n25560), .ZN(n27703) );
  XNOR2_X1 U17472 ( .A(n21456), .B(n21455), .ZN(n23427) );
  NAND2_X1 U17479 ( .A1(n20035), .A2(n29186), .ZN(n22643) );
  NAND3_X1 U17498 ( .A1(n5293), .A2(n5292), .A3(n22499), .ZN(n24613) );
  BUF_X1 U17598 ( .A(n8237), .Z(n29110) );
  XNOR2_X1 U17604 ( .A(n6969), .B(Key[104]), .ZN(n8237) );
  BUF_X1 U17606 ( .A(n26089), .Z(n29111) );
  OAI22_X1 U17618 ( .A1(n23951), .A2(n23950), .B1(n5004), .B2(n24810), .ZN(
        n26089) );
  XNOR2_X1 U17715 ( .A(n22361), .B(n22360), .ZN(n960) );
  XNOR2_X1 U17716 ( .A(n7085), .B(Key[4]), .ZN(n29112) );
  XNOR2_X1 U17802 ( .A(n7085), .B(Key[4]), .ZN(n7891) );
  BUF_X1 U17959 ( .A(n23733), .Z(n1862) );
  BUF_X1 U18090 ( .A(n23562), .Z(n29115) );
  XNOR2_X1 U18120 ( .A(n18742), .B(n18741), .ZN(n20090) );
  BUF_X2 U18139 ( .A(n11288), .Z(n29116) );
  XNOR2_X1 U18354 ( .A(n10326), .B(n10325), .ZN(n11288) );
  NOR2_X1 U18470 ( .A1(n26293), .A2(n26294), .ZN(n29117) );
  NOR2_X1 U18476 ( .A1(n26293), .A2(n26294), .ZN(n29118) );
  NOR2_X1 U18735 ( .A1(n26293), .A2(n26294), .ZN(n27768) );
  XNOR2_X1 U18820 ( .A(Key[44]), .B(Plaintext[44]), .ZN(n29119) );
  OR2_X1 U18974 ( .A1(n23782), .A2(n23781), .ZN(n29120) );
  XNOR2_X1 U18981 ( .A(Key[44]), .B(Plaintext[44]), .ZN(n8136) );
  MUX2_X2 U18999 ( .A(n21102), .B(n21101), .S(n28916), .Z(n22768) );
  INV_X1 U19073 ( .A(n28091), .ZN(n29121) );
  AOI22_X1 U19094 ( .A1(n26732), .A2(n1623), .B1(n26730), .B2(n29579), .ZN(
        n28091) );
  INV_X1 U19113 ( .A(n20333), .ZN(n28186) );
  XNOR2_X1 U19118 ( .A(n1141), .B(n9628), .ZN(n29122) );
  XNOR2_X1 U19127 ( .A(n1141), .B(n9628), .ZN(n11260) );
  XOR2_X1 U19235 ( .A(n18863), .B(n18395), .Z(n29124) );
  BUF_X1 U19317 ( .A(n19562), .Z(n29125) );
  XOR2_X1 U19338 ( .A(n22385), .B(n22384), .Z(n29126) );
  OAI211_X1 U19351 ( .C1(n17224), .C2(n16908), .A(n16917), .B(n16835), .ZN(
        n19562) );
  XOR2_X1 U19389 ( .A(n16209), .B(n16210), .Z(n29127) );
  AOI22_X1 U19398 ( .A1(n22989), .A2(n22990), .B1(n23624), .B2(n22988), .ZN(
        n29128) );
  AOI22_X1 U19440 ( .A1(n22989), .A2(n22990), .B1(n23624), .B2(n22988), .ZN(
        n24436) );
  NAND3_X1 U19475 ( .A1(n28362), .A2(n3359), .A3(n28361), .ZN(n29129) );
  NAND3_X1 U19517 ( .A1(n28362), .A2(n3359), .A3(n28361), .ZN(n26073) );
  XNOR2_X1 U19543 ( .A(Key[68]), .B(Plaintext[68]), .ZN(n29130) );
  XNOR2_X1 U19548 ( .A(Key[68]), .B(Plaintext[68]), .ZN(n8023) );
  AND2_X1 U19687 ( .A1(n10884), .A2(n11282), .ZN(n29212) );
  XOR2_X1 U19695 ( .A(n22335), .B(n22336), .Z(n29131) );
  AOI22_X1 U19732 ( .A1(n1362), .A2(n17314), .B1(n1361), .B2(n29550), .ZN(
        n17826) );
  XNOR2_X1 U19733 ( .A(n24866), .B(n24865), .ZN(n29132) );
  XNOR2_X1 U19734 ( .A(n12412), .B(n12411), .ZN(n29133) );
  XNOR2_X1 U19835 ( .A(n18916), .B(n18917), .ZN(n21092) );
  NOR2_X2 U19840 ( .A1(n28103), .A2(n5037), .ZN(n28089) );
  XOR2_X1 U19856 ( .A(n10149), .B(n9619), .Z(n9906) );
  XNOR2_X1 U19911 ( .A(n21999), .B(n22812), .ZN(n29136) );
  XNOR2_X1 U19912 ( .A(Key[119]), .B(Plaintext[119]), .ZN(n9113) );
  OAI21_X1 U20079 ( .B1(n11143), .B2(n11142), .A(n1452), .ZN(n29137) );
  BUF_X1 U20140 ( .A(n17565), .Z(n29138) );
  XNOR2_X1 U20284 ( .A(n2790), .B(n16267), .ZN(n17565) );
  OR2_X1 U20316 ( .A1(n29330), .A2(n26280), .ZN(n26801) );
  OAI21_X1 U20341 ( .B1(n11644), .B2(n11643), .A(n11642), .ZN(n29140) );
  NOR2_X1 U20444 ( .A1(n11636), .A2(n11633), .ZN(n11673) );
  OAI21_X1 U20544 ( .B1(n11644), .B2(n11643), .A(n11642), .ZN(n13012) );
  CLKBUF_X3 U20743 ( .A(n27378), .Z(n295) );
  XNOR2_X1 U20822 ( .A(n15827), .B(n15826), .ZN(n29142) );
  INV_X1 U20831 ( .A(n19838), .ZN(n29143) );
  XNOR2_X1 U20839 ( .A(n15827), .B(n15826), .ZN(n17557) );
  XNOR2_X1 U20843 ( .A(n17813), .B(n17812), .ZN(n29144) );
  XNOR2_X1 U20879 ( .A(n18563), .B(n18564), .ZN(n29145) );
  XNOR2_X1 U20950 ( .A(n18564), .B(n18563), .ZN(n29146) );
  XNOR2_X1 U20959 ( .A(n9599), .B(n9600), .ZN(n29149) );
  AND2_X1 U20984 ( .A1(n11126), .A2(n10114), .ZN(n11403) );
  AND2_X1 U21031 ( .A1(n29618), .A2(n22452), .ZN(n29169) );
  OAI21_X1 U21051 ( .B1(n15298), .B2(n15297), .A(n15296), .ZN(n29151) );
  XNOR2_X1 U21079 ( .A(n15330), .B(n15329), .ZN(n29152) );
  OAI21_X1 U21099 ( .B1(n15298), .B2(n15297), .A(n15296), .ZN(n16580) );
  OAI211_X1 U21116 ( .C1(n13888), .C2(n14313), .A(n13887), .B(n3602), .ZN(
        n29153) );
  AOI21_X1 U21117 ( .B1(n3634), .B2(n24459), .A(n24458), .ZN(n29154) );
  AOI21_X1 U21174 ( .B1(n3634), .B2(n24459), .A(n24458), .ZN(n29155) );
  OAI211_X1 U21177 ( .C1(n13888), .C2(n14313), .A(n13887), .B(n3602), .ZN(
        n15160) );
  AOI21_X1 U21179 ( .B1(n3634), .B2(n24459), .A(n24458), .ZN(n25759) );
  NAND2_X1 U21180 ( .A1(n18456), .A2(n29156), .ZN(n3865) );
  OR3_X1 U21242 ( .A1(n27492), .A2(n27494), .A3(n27497), .ZN(n27500) );
  XOR2_X1 U21251 ( .A(n22115), .B(n22114), .Z(n29157) );
  INV_X1 U21272 ( .A(n2433), .ZN(n29158) );
  XNOR2_X1 U21348 ( .A(n25452), .B(n25451), .ZN(n29159) );
  NOR2_X1 U21367 ( .A1(n25472), .A2(n28670), .ZN(n29160) );
  NOR2_X1 U21384 ( .A1(n25472), .A2(n28670), .ZN(n29161) );
  NOR2_X1 U21386 ( .A1(n25472), .A2(n28670), .ZN(n28024) );
  NAND2_X1 U21422 ( .A1(n4305), .A2(n9211), .ZN(n9207) );
  XNOR2_X1 U21423 ( .A(n29163), .B(n22761), .ZN(n22767) );
  XNOR2_X1 U21447 ( .A(n22758), .B(n22757), .ZN(n29163) );
  NAND2_X1 U21487 ( .A1(n29165), .A2(n29164), .ZN(n20767) );
  NAND2_X1 U21565 ( .A1(n20287), .A2(n20286), .ZN(n29164) );
  NAND2_X1 U21591 ( .A1(n20288), .A2(n29166), .ZN(n29165) );
  NOR3_X1 U21621 ( .A1(n29168), .A2(n26536), .A3(n26535), .ZN(Ciphertext[25])
         );
  NAND2_X1 U21632 ( .A1(n28605), .A2(n8200), .ZN(n28246) );
  NAND2_X1 U21722 ( .A1(n7423), .A2(n3112), .ZN(n7370) );
  NAND3_X1 U21826 ( .A1(n3161), .A2(n11349), .A3(n11355), .ZN(n11354) );
  NAND2_X1 U21889 ( .A1(n10765), .A2(n10764), .ZN(n13109) );
  NAND2_X1 U22216 ( .A1(n13889), .A2(n29153), .ZN(n29171) );
  NAND2_X1 U22218 ( .A1(n13890), .A2(n545), .ZN(n29172) );
  NAND2_X1 U22347 ( .A1(n4835), .A2(n15464), .ZN(n29173) );
  NAND2_X1 U22363 ( .A1(n24073), .A2(n24072), .ZN(n29174) );
  NAND2_X1 U22390 ( .A1(n5856), .A2(n23418), .ZN(n23097) );
  NAND2_X1 U22437 ( .A1(n4274), .A2(n4275), .ZN(n10545) );
  NAND3_X1 U22474 ( .A1(n386), .A2(n4306), .A3(n28408), .ZN(n5358) );
  NAND2_X1 U22506 ( .A1(n17873), .A2(n17938), .ZN(n17874) );
  NAND3_X1 U22514 ( .A1(n17416), .A2(n5430), .A3(n17413), .ZN(n29176) );
  NAND3_X1 U22573 ( .A1(n21661), .A2(n21654), .A3(n21655), .ZN(n20835) );
  NAND2_X1 U22692 ( .A1(n529), .A2(n17439), .ZN(n29177) );
  NAND2_X1 U22799 ( .A1(n17846), .A2(n18137), .ZN(n17848) );
  NAND2_X1 U22807 ( .A1(n8590), .A2(n8973), .ZN(n8597) );
  NAND2_X1 U22818 ( .A1(n21449), .A2(n21448), .ZN(n29178) );
  NAND2_X1 U22819 ( .A1(n29179), .A2(n11873), .ZN(n12849) );
  NAND2_X1 U22829 ( .A1(n6305), .A2(n6304), .ZN(n29179) );
  NAND2_X1 U22837 ( .A1(n29181), .A2(n20265), .ZN(n29180) );
  NAND2_X1 U22840 ( .A1(n6202), .A2(n6204), .ZN(n29181) );
  INV_X1 U22848 ( .A(n20265), .ZN(n29183) );
  NAND3_X1 U22904 ( .A1(n28745), .A2(n18486), .A3(n18493), .ZN(n1997) );
  NAND2_X1 U22910 ( .A1(n20478), .A2(n20477), .ZN(n20232) );
  XNOR2_X2 U22915 ( .A(n15560), .B(n15559), .ZN(n17338) );
  NAND3_X1 U22987 ( .A1(n412), .A2(n21678), .A3(n21448), .ZN(n2909) );
  NAND2_X1 U22988 ( .A1(n29185), .A2(n585), .ZN(n2954) );
  NAND2_X1 U22996 ( .A1(n11026), .A2(n11027), .ZN(n29185) );
  OAI211_X1 U23024 ( .C1(n21633), .C2(n21631), .A(n21036), .B(n28797), .ZN(
        n29186) );
  NAND2_X1 U23054 ( .A1(n24155), .A2(n28785), .ZN(n24249) );
  NAND4_X1 U23086 ( .A1(n25671), .A2(n25672), .A3(n29188), .A4(n29187), .ZN(
        n25675) );
  NAND2_X1 U23087 ( .A1(n25658), .A2(n27350), .ZN(n29187) );
  NAND2_X1 U23120 ( .A1(n27351), .A2(n25657), .ZN(n29188) );
  NAND2_X1 U23288 ( .A1(n23535), .A2(n23531), .ZN(n5481) );
  OR2_X1 U23311 ( .A1(n24237), .A2(n29642), .ZN(n6238) );
  NAND2_X1 U23384 ( .A1(n29189), .A2(n28821), .ZN(n24155) );
  NAND2_X1 U23385 ( .A1(n23608), .A2(n23211), .ZN(n29189) );
  NAND2_X1 U23434 ( .A1(n3549), .A2(n17364), .ZN(n16760) );
  NAND2_X1 U23435 ( .A1(n17234), .A2(n17368), .ZN(n17364) );
  NAND2_X1 U23506 ( .A1(n1576), .A2(n512), .ZN(n29191) );
  NAND2_X1 U23535 ( .A1(n1577), .A2(n16862), .ZN(n29192) );
  NAND2_X2 U23543 ( .A1(n29193), .A2(n24519), .ZN(n25909) );
  NAND2_X1 U23563 ( .A1(n28284), .A2(n28285), .ZN(n26578) );
  NOR2_X2 U23587 ( .A1(n5194), .A2(n19962), .ZN(n21472) );
  NAND2_X1 U23683 ( .A1(n4914), .A2(n1574), .ZN(n29194) );
  AND3_X2 U23684 ( .A1(n19185), .A2(n29197), .A3(n29196), .ZN(n21372) );
  NAND2_X1 U23723 ( .A1(n19179), .A2(n19863), .ZN(n29196) );
  NAND2_X1 U23724 ( .A1(n1041), .A2(n19867), .ZN(n29197) );
  OAI211_X2 U23756 ( .C1(n1750), .C2(n9410), .A(n29198), .B(n6505), .ZN(n10271) );
  NAND2_X1 U23806 ( .A1(n9040), .A2(n9410), .ZN(n29198) );
  NAND3_X1 U23938 ( .A1(n2422), .A2(n10699), .A3(n2423), .ZN(n11491) );
  NAND3_X1 U23965 ( .A1(n16830), .A2(n2485), .A3(n16829), .ZN(n2484) );
  NAND3_X1 U24032 ( .A1(n10754), .A2(n11152), .A3(n10804), .ZN(n10755) );
  NAND3_X1 U24033 ( .A1(n12022), .A2(n29209), .A3(n12428), .ZN(n1369) );
  NAND3_X1 U24079 ( .A1(n6434), .A2(n6307), .A3(n14310), .ZN(n6433) );
  NAND2_X1 U24098 ( .A1(n5981), .A2(n14393), .ZN(n29201) );
  NOR2_X1 U24135 ( .A1(n29202), .A2(n11831), .ZN(n11832) );
  NOR3_X1 U24137 ( .A1(n6281), .A2(n12207), .A3(n12206), .ZN(n29202) );
  NAND2_X1 U24228 ( .A1(n465), .A2(n24633), .ZN(n24560) );
  NAND3_X1 U24268 ( .A1(n15322), .A2(n15327), .A3(n15013), .ZN(n1106) );
  NAND2_X1 U24326 ( .A1(n1068), .A2(n27955), .ZN(n29277) );
  NAND3_X1 U24334 ( .A1(n18158), .A2(n18160), .A3(n18159), .ZN(n18161) );
  NOR2_X1 U24392 ( .A1(n4214), .A2(n29204), .ZN(n17061) );
  NAND2_X1 U24431 ( .A1(n7750), .A2(n8161), .ZN(n7157) );
  NAND2_X1 U24623 ( .A1(n29206), .A2(n29205), .ZN(n16840) );
  NAND2_X1 U24624 ( .A1(n17312), .A2(n29550), .ZN(n29205) );
  NAND2_X1 U24713 ( .A1(n16836), .A2(n17560), .ZN(n29206) );
  NAND2_X1 U24747 ( .A1(n15514), .A2(n15515), .ZN(n15277) );
  NAND2_X1 U24807 ( .A1(n14886), .A2(n29207), .ZN(n6668) );
  OR2_X1 U24811 ( .A1(n14972), .A2(n14969), .ZN(n29207) );
  INV_X1 U24813 ( .A(n10816), .ZN(n28207) );
  XNOR2_X1 U24890 ( .A(n8479), .B(n8480), .ZN(n10816) );
  NAND3_X1 U24909 ( .A1(n512), .A2(n17802), .A3(n29507), .ZN(n227) );
  NAND3_X1 U24928 ( .A1(n28820), .A2(n20039), .A3(n20090), .ZN(n6410) );
  OR2_X1 U24964 ( .A1(n22991), .A2(n23563), .ZN(n22993) );
  NAND2_X1 U24972 ( .A1(n15436), .A2(n15300), .ZN(n14664) );
  NAND2_X1 U24976 ( .A1(n17508), .A2(n17829), .ZN(n28323) );
  OAI21_X1 U24977 ( .B1(n10568), .B2(n10623), .A(n11896), .ZN(n29208) );
  NAND2_X1 U24987 ( .A1(n29210), .A2(n29209), .ZN(n26) );
  NAND2_X1 U24994 ( .A1(n11467), .A2(n12428), .ZN(n29210) );
  OAI211_X2 U25003 ( .C1(n15268), .C2(n15494), .A(n14619), .B(n29211), .ZN(
        n16399) );
  NAND2_X1 U25023 ( .A1(n11283), .A2(n29212), .ZN(n10380) );
  NAND2_X1 U25047 ( .A1(n10779), .A2(n10966), .ZN(n10782) );
  NAND2_X1 U25127 ( .A1(n6556), .A2(n24538), .ZN(n24539) );
  NAND3_X1 U25140 ( .A1(n6692), .A2(n6691), .A3(n8979), .ZN(n203) );
  OAI21_X1 U25141 ( .B1(n7784), .B2(n2670), .A(n7783), .ZN(n29214) );
  NAND2_X1 U25193 ( .A1(n454), .A2(n4820), .ZN(n6435) );
  NAND2_X1 U25216 ( .A1(n27908), .A2(n27092), .ZN(n27883) );
  NAND3_X1 U25242 ( .A1(n11930), .A2(n568), .A3(n12267), .ZN(n1491) );
  MUX2_X1 U25243 ( .A(n17767), .B(n18387), .S(n18388), .Z(n17736) );
  NAND2_X1 U25269 ( .A1(n29215), .A2(n10488), .ZN(n10648) );
  NAND2_X1 U25294 ( .A1(n10485), .A2(n11057), .ZN(n29215) );
  OAI21_X1 U25305 ( .B1(n2425), .B2(n2029), .A(n8958), .ZN(n8624) );
  OR2_X1 U25345 ( .A1(n18414), .A2(n18121), .ZN(n3915) );
  NAND2_X1 U25360 ( .A1(n27381), .A2(n29217), .ZN(n27385) );
  OAI21_X1 U25400 ( .B1(n27376), .B2(n29219), .A(n29218), .ZN(n29217) );
  NAND2_X1 U25401 ( .A1(n29220), .A2(n22878), .ZN(n24278) );
  NAND4_X1 U25408 ( .A1(n1151), .A2(n1284), .A3(n2202), .A4(n1150), .ZN(n29220) );
  NAND2_X1 U25495 ( .A1(n28332), .A2(n28334), .ZN(n11180) );
  NAND2_X1 U25496 ( .A1(n9435), .A2(n29221), .ZN(n7683) );
  NAND3_X1 U25541 ( .A1(n15029), .A2(n15430), .A3(n15028), .ZN(n15035) );
  AOI22_X2 U25551 ( .A1(n9693), .A2(n28405), .B1(n9694), .B2(n592), .ZN(n12186) );
  NAND2_X1 U25589 ( .A1(n29222), .A2(n9060), .ZN(n8107) );
  OAI21_X1 U25607 ( .B1(n9059), .B2(n9064), .A(n8397), .ZN(n29222) );
  NAND2_X1 U25704 ( .A1(n29223), .A2(n17434), .ZN(n4428) );
  NAND2_X1 U25723 ( .A1(n17308), .A2(n16962), .ZN(n29223) );
  NAND2_X1 U25765 ( .A1(n21375), .A2(n21702), .ZN(n29224) );
  NAND2_X1 U25766 ( .A1(n29226), .A2(n29227), .ZN(n29225) );
  INV_X1 U25801 ( .A(n21378), .ZN(n29226) );
  INV_X2 U25920 ( .A(n21709), .ZN(n29227) );
  OAI21_X1 U25998 ( .B1(n7795), .B2(n7796), .A(n29229), .ZN(n7544) );
  NAND2_X1 U25999 ( .A1(n7796), .A2(n7542), .ZN(n29229) );
  NAND3_X1 U26068 ( .A1(n29230), .A2(n7685), .A3(n7520), .ZN(n7013) );
  NAND2_X1 U26069 ( .A1(n7684), .A2(n7517), .ZN(n29230) );
  AND3_X2 U26110 ( .A1(n2270), .A2(n26335), .A3(n2269), .ZN(n27818) );
  XNOR2_X2 U26172 ( .A(n6467), .B(n19163), .ZN(n5225) );
  OAI21_X1 U26240 ( .B1(n27819), .B2(n29232), .A(n29231), .ZN(n26679) );
  NAND2_X1 U26255 ( .A1(n27819), .A2(n27818), .ZN(n29231) );
  INV_X1 U26339 ( .A(n27795), .ZN(n29232) );
  NAND3_X1 U26385 ( .A1(n20056), .A2(n6114), .A3(n20171), .ZN(n29233) );
  NAND2_X1 U26397 ( .A1(n11242), .A2(n11069), .ZN(n10198) );
  NAND2_X1 U26523 ( .A1(n7980), .A2(n7985), .ZN(n7459) );
  OAI21_X1 U26555 ( .B1(n20400), .B2(n20401), .A(n20562), .ZN(n29235) );
  INV_X1 U26582 ( .A(n28580), .ZN(n29236) );
  NAND2_X1 U26596 ( .A1(n21560), .A2(n5953), .ZN(n20862) );
  NAND3_X1 U26618 ( .A1(n5126), .A2(n28658), .A3(n29315), .ZN(n4472) );
  NAND2_X1 U26649 ( .A1(n28542), .A2(n26948), .ZN(n6469) );
  NAND2_X1 U26716 ( .A1(n1333), .A2(n1332), .ZN(n29237) );
  NAND2_X1 U26769 ( .A1(n2329), .A2(n1708), .ZN(n29238) );
  AND3_X2 U26783 ( .A1(n29239), .A2(n11766), .A3(n6725), .ZN(n15108) );
  NAND2_X1 U26910 ( .A1(n11765), .A2(n293), .ZN(n29239) );
  NAND3_X1 U27074 ( .A1(n7074), .A2(n7884), .A3(n7882), .ZN(n7076) );
  NAND2_X1 U27089 ( .A1(n9083), .A2(n9082), .ZN(n7490) );
  NAND2_X1 U27141 ( .A1(n2099), .A2(n8270), .ZN(n9083) );
  XNOR2_X2 U27142 ( .A(n20471), .B(n20472), .ZN(n23531) );
  AOI21_X2 U27143 ( .B1(n17231), .B2(n871), .A(n17230), .ZN(n18148) );
  NAND2_X1 U27253 ( .A1(n2357), .A2(n12162), .ZN(n12171) );
  OR2_X1 U27269 ( .A1(n17383), .A2(n17384), .ZN(n29240) );
  NAND2_X1 U27271 ( .A1(n8808), .A2(n8809), .ZN(n29242) );
  NAND2_X1 U27272 ( .A1(n4195), .A2(n24669), .ZN(n4194) );
  OR3_X1 U27304 ( .A1(n18042), .A2(n18421), .A3(n29507), .ZN(n18425) );
  NAND2_X1 U27339 ( .A1(n29245), .A2(n29243), .ZN(n13191) );
  OAI21_X1 U27344 ( .B1(n12004), .B2(n11760), .A(n11758), .ZN(n29244) );
  OAI21_X1 U27354 ( .B1(n11757), .B2(n11756), .A(n12004), .ZN(n29245) );
  NAND2_X1 U27425 ( .A1(n14424), .A2(n14425), .ZN(n4523) );
  NAND2_X1 U27487 ( .A1(n29246), .A2(n28813), .ZN(n21676) );
  NAND2_X1 U27513 ( .A1(n20211), .A2(n20210), .ZN(n29246) );
  NAND2_X1 U27519 ( .A1(n24351), .A2(n24712), .ZN(n29248) );
  NAND2_X1 U27547 ( .A1(n23070), .A2(n28416), .ZN(n29249) );
  NAND3_X1 U27582 ( .A1(n2281), .A2(n23816), .A3(n28609), .ZN(n3990) );
  NOR2_X1 U27600 ( .A1(n29251), .A2(n23819), .ZN(n23822) );
  NAND2_X1 U27611 ( .A1(n407), .A2(n23290), .ZN(n29251) );
  NAND2_X1 U27727 ( .A1(n21669), .A2(n22401), .ZN(n2072) );
  XNOR2_X2 U27729 ( .A(Key[80]), .B(Plaintext[80]), .ZN(n7690) );
  NAND2_X1 U27751 ( .A1(n29253), .A2(n23100), .ZN(n23101) );
  OAI21_X1 U27776 ( .B1(n23098), .B2(n23097), .A(n23096), .ZN(n29253) );
  INV_X1 U27790 ( .A(n24813), .ZN(n220) );
  NAND3_X1 U27934 ( .A1(n29255), .A2(n5707), .A3(n5710), .ZN(n5704) );
  NAND2_X1 U28001 ( .A1(n5709), .A2(n11237), .ZN(n29255) );
  NOR2_X2 U28033 ( .A1(n29256), .A2(n1312), .ZN(n22913) );
  NAND2_X1 U28036 ( .A1(n7744), .A2(n7743), .ZN(n7524) );
  NAND2_X1 U28110 ( .A1(n29257), .A2(n11538), .ZN(n6146) );
  NAND2_X1 U28124 ( .A1(n11685), .A2(n11540), .ZN(n29257) );
  OAI21_X1 U28125 ( .B1(n6906), .B2(n2107), .A(n24195), .ZN(n24197) );
  NAND2_X1 U28153 ( .A1(n24644), .A2(n24642), .ZN(n24195) );
  NAND2_X1 U28154 ( .A1(n14613), .A2(n14612), .ZN(n14614) );
  NAND2_X1 U28160 ( .A1(n7685), .A2(n7844), .ZN(n7686) );
  OAI211_X2 U28164 ( .C1(n21321), .C2(n21137), .A(n21589), .B(n4962), .ZN(
        n22418) );
  NOR2_X1 U28166 ( .A1(n29258), .A2(n27432), .ZN(n25426) );
  OAI21_X1 U28176 ( .B1(n26829), .B2(n27434), .A(n26708), .ZN(n29258) );
  AOI21_X1 U28197 ( .B1(n6194), .B2(n6197), .A(n6196), .ZN(n29259) );
  XNOR2_X1 U28199 ( .A(n29261), .B(n29260), .ZN(Ciphertext[153]) );
  INV_X1 U28205 ( .A(n27894), .ZN(n29260) );
  OAI211_X1 U28213 ( .C1(n27892), .C2(n27893), .A(n27891), .B(n27890), .ZN(
        n29261) );
  NOR2_X2 U28216 ( .A1(n29262), .A2(n20442), .ZN(n21513) );
  AOI22_X1 U28217 ( .A1(n20439), .A2(n20438), .B1(n20436), .B2(n29508), .ZN(
        n29262) );
  NAND2_X1 U28218 ( .A1(n6864), .A2(n6865), .ZN(n4238) );
  NAND2_X1 U28219 ( .A1(n10742), .A2(n29263), .ZN(n4274) );
  NAND2_X1 U28220 ( .A1(n223), .A2(n14894), .ZN(n3360) );
  NOR2_X2 U28221 ( .A1(n21517), .A2(n21518), .ZN(n22615) );
  NAND2_X1 U28222 ( .A1(n71), .A2(n4448), .ZN(n29264) );
  NAND3_X1 U28223 ( .A1(n20189), .A2(n6261), .A3(n19959), .ZN(n6260) );
  XNOR2_X1 U28224 ( .A(n15849), .B(n2465), .ZN(n15851) );
  NAND2_X1 U28225 ( .A1(n3777), .A2(n14875), .ZN(n15849) );
  NAND2_X1 U28226 ( .A1(n27156), .A2(n28180), .ZN(n27158) );
  NAND2_X1 U28227 ( .A1(n17687), .A2(n20417), .ZN(n20418) );
  NAND2_X1 U28229 ( .A1(n21623), .A2(n22141), .ZN(n29265) );
  NAND2_X1 U28230 ( .A1(n27663), .A2(n27661), .ZN(n27652) );
  NOR2_X2 U28231 ( .A1(n23278), .A2(n23279), .ZN(n24083) );
  NAND2_X1 U28234 ( .A1(n21708), .A2(n496), .ZN(n6104) );
  NAND2_X1 U28235 ( .A1(n21703), .A2(n21277), .ZN(n21708) );
  NAND2_X1 U28236 ( .A1(n6086), .A2(n20406), .ZN(n6085) );
  AND2_X2 U28237 ( .A1(n3308), .A2(n7335), .ZN(n8562) );
  NAND2_X1 U28240 ( .A1(n5054), .A2(n5055), .ZN(n3648) );
  NAND2_X1 U28242 ( .A1(n14417), .A2(n14418), .ZN(n14449) );
  NAND2_X1 U28243 ( .A1(n19052), .A2(n29584), .ZN(n19057) );
  NAND2_X1 U28244 ( .A1(n24894), .A2(n23982), .ZN(n29268) );
  NAND2_X1 U28245 ( .A1(n24295), .A2(n24294), .ZN(n29269) );
  NAND3_X1 U28246 ( .A1(n1268), .A2(n1267), .A3(n1269), .ZN(n1266) );
  NAND4_X2 U28247 ( .A1(n6216), .A2(n6217), .A3(n29271), .A4(n29270), .ZN(
        n16185) );
  NAND2_X1 U28248 ( .A1(n15502), .A2(n14923), .ZN(n29270) );
  NAND2_X1 U28249 ( .A1(n14707), .A2(n15506), .ZN(n29271) );
  NAND2_X1 U28250 ( .A1(n1739), .A2(n25656), .ZN(n28669) );
  NOR2_X1 U28251 ( .A1(n26738), .A2(n26737), .ZN(n1739) );
  INV_X1 U28252 ( .A(n7847), .ZN(n7260) );
  NAND2_X1 U28253 ( .A1(n7846), .A2(n8024), .ZN(n7847) );
  NAND2_X1 U28254 ( .A1(n26686), .A2(n395), .ZN(n29288) );
  NAND2_X1 U28255 ( .A1(n27300), .A2(n26879), .ZN(n26686) );
  NAND2_X1 U28256 ( .A1(n29272), .A2(n18334), .ZN(n18336) );
  NAND2_X1 U28257 ( .A1(n18333), .A2(n817), .ZN(n29272) );
  XNOR2_X1 U28258 ( .A(n29273), .B(n10409), .ZN(n10414) );
  NAND3_X1 U28259 ( .A1(n3877), .A2(n18423), .A3(n1942), .ZN(n3876) );
  NAND2_X1 U28260 ( .A1(n29274), .A2(n16862), .ZN(n5495) );
  NAND3_X1 U28261 ( .A1(n2789), .A2(n7511), .A3(n2788), .ZN(n3683) );
  XNOR2_X1 U28262 ( .A(n29275), .B(n28097), .ZN(Ciphertext[189]) );
  NAND3_X1 U28263 ( .A1(n28095), .A2(n3470), .A3(n3469), .ZN(n29275) );
  NAND2_X1 U28264 ( .A1(n29276), .A2(n11140), .ZN(n1452) );
  NAND2_X1 U28265 ( .A1(n11138), .A2(n11139), .ZN(n29276) );
  OR2_X1 U28266 ( .A1(n11473), .A2(n10648), .ZN(n12345) );
  INV_X1 U28267 ( .A(n14570), .ZN(n15076) );
  NAND2_X1 U28268 ( .A1(n14874), .A2(n15071), .ZN(n14570) );
  NAND2_X1 U28269 ( .A1(n142), .A2(n602), .ZN(n8130) );
  XNOR2_X1 U28270 ( .A(n29277), .B(n27957), .ZN(Ciphertext[162]) );
  AOI22_X1 U28272 ( .A1(n1684), .A2(n27364), .B1(n26496), .B2(n27370), .ZN(
        n29278) );
  NAND2_X1 U28273 ( .A1(n7919), .A2(n7619), .ZN(n7430) );
  AOI21_X1 U28274 ( .B1(n19898), .B2(n3009), .A(n19897), .ZN(n21124) );
  AND3_X2 U28275 ( .A1(n26154), .A2(n26153), .A3(n29279), .ZN(n27465) );
  NAND3_X1 U28276 ( .A1(n28286), .A2(n25418), .A3(n6826), .ZN(n29279) );
  NAND2_X1 U28277 ( .A1(n29281), .A2(n29280), .ZN(n26744) );
  NAND2_X1 U28278 ( .A1(n26739), .A2(n26235), .ZN(n29280) );
  NAND2_X1 U28279 ( .A1(n26738), .A2(n26737), .ZN(n29281) );
  OAI211_X2 U28280 ( .C1(n20846), .C2(n6247), .A(n5175), .B(n29282), .ZN(
        n22279) );
  NAND3_X1 U28281 ( .A1(n19904), .A2(n21125), .A3(n21461), .ZN(n29282) );
  OAI211_X1 U28282 ( .C1(n26608), .C2(n27458), .A(n29284), .B(n29283), .ZN(
        n26609) );
  NAND2_X1 U28283 ( .A1(n26605), .A2(n27447), .ZN(n29283) );
  NAND2_X1 U28284 ( .A1(n27458), .A2(n26606), .ZN(n29284) );
  NAND2_X1 U28285 ( .A1(n29286), .A2(n29285), .ZN(n26630) );
  OR3_X1 U28286 ( .A1(n29481), .A2(n26733), .A3(n26995), .ZN(n29285) );
  NAND2_X1 U28287 ( .A1(n26628), .A2(n26995), .ZN(n29286) );
  AOI22_X1 U28289 ( .A1(n26887), .A2(n5425), .B1(n29288), .B2(n29287), .ZN(
        n26446) );
  INV_X1 U28290 ( .A(n444), .ZN(n29287) );
  OAI21_X1 U28291 ( .B1(n18157), .B2(n17744), .A(n29289), .ZN(n2501) );
  NOR2_X1 U28292 ( .A1(n17614), .A2(n17616), .ZN(n17307) );
  NAND2_X1 U28293 ( .A1(n6001), .A2(n17303), .ZN(n17614) );
  NAND2_X1 U28294 ( .A1(n29290), .A2(n15399), .ZN(n6262) );
  NAND2_X1 U28296 ( .A1(n3900), .A2(n29291), .ZN(n3166) );
  NOR2_X2 U28297 ( .A1(n2534), .A2(n29292), .ZN(n21268) );
  NAND2_X1 U28298 ( .A1(n28383), .A2(n28384), .ZN(n29292) );
  NAND2_X1 U28299 ( .A1(n1109), .A2(n1110), .ZN(n21013) );
  NAND3_X1 U28302 ( .A1(n29121), .A2(n29056), .A3(n28089), .ZN(n28080) );
  OAI22_X1 U28303 ( .A1(n27204), .A2(n27547), .B1(n27205), .B2(n28422), .ZN(
        n27206) );
  XNOR2_X1 U28305 ( .A(n15721), .B(n15722), .ZN(n17362) );
  INV_X1 U28307 ( .A(n20351), .ZN(n21553) );
  XOR2_X1 U28308 ( .A(n24868), .B(n24869), .Z(n29293) );
  AOI21_X2 U2951 ( .B1(n12673), .B2(n190), .A(n12672), .ZN(n15103) );
  OAI21_X2 U1024 ( .B1(n22975), .B2(n22974), .A(n22973), .ZN(n24434) );
  OR2_X2 U827 ( .A1(n15479), .A2(n15478), .ZN(n16319) );
  OAI211_X2 U9166 ( .C1(n8130), .C2(n8129), .A(n8128), .B(n8127), .ZN(n2845)
         );
  BUF_X2 U18281 ( .A(n12711), .Z(n14204) );
  NAND2_X2 U3585 ( .A1(n4111), .A2(n6874), .ZN(n8642) );
  NAND3_X2 U1493 ( .A1(n28982), .A2(n5865), .A3(n1132), .ZN(n21549) );
  BUF_X2 U270 ( .A(n26841), .Z(n27088) );
  INV_X2 U1724 ( .A(n20425), .ZN(n21823) );
  NAND2_X2 U28187 ( .A1(n28756), .A2(n15210), .ZN(n16404) );
  AND2_X2 U1359 ( .A1(n5462), .A2(n12243), .ZN(n13054) );
  AND3_X2 U3064 ( .A1(n2682), .A2(n6280), .A3(n2685), .ZN(n13523) );
  BUF_X1 U2375 ( .A(n7838), .Z(n7700) );
  NOR2_X2 U1126 ( .A1(n23597), .A2(n23467), .ZN(n24975) );
  NAND3_X2 U730 ( .A1(n20126), .A2(n20127), .A3(n20128), .ZN(n5827) );
  BUF_X1 U426 ( .A(n10318), .Z(n11076) );
  BUF_X1 U2606 ( .A(n19787), .Z(n20632) );
  XNOR2_X2 U1531 ( .A(n19177), .B(n19178), .ZN(n20496) );
  XNOR2_X2 U1343 ( .A(n13023), .B(n13022), .ZN(n14362) );
  XNOR2_X2 U5227 ( .A(n1619), .B(n18641), .ZN(n20209) );
  NAND3_X2 U10374 ( .A1(n28372), .A2(n8010), .A3(n8011), .ZN(n9504) );
  AOI22_X2 U9320 ( .A1(n5022), .A2(n18406), .B1(n18709), .B2(n18407), .ZN(
        n18948) );
  AND2_X2 U619 ( .A1(n10841), .A2(n10840), .ZN(n12244) );
  AND2_X2 U2538 ( .A1(n3855), .A2(n21435), .ZN(n21442) );
  OAI21_X2 U9076 ( .B1(n17180), .B2(n1801), .A(n17178), .ZN(n18411) );
  OAI21_X2 U659 ( .B1(n23219), .B2(n23610), .A(n23218), .ZN(n24248) );
  BUF_X2 U312 ( .A(n8608), .Z(n9532) );
  BUF_X2 U678 ( .A(n17679), .Z(n18478) );
  BUF_X1 U1274 ( .A(n21729), .Z(n1929) );
  AND3_X2 U2913 ( .A1(n4519), .A2(n4521), .A3(n14430), .ZN(n15506) );
  NOR2_X2 U789 ( .A1(n2201), .A2(n22744), .ZN(n24551) );
  AOI21_X2 U10018 ( .B1(n18347), .B2(n18346), .A(n18345), .ZN(n18680) );
  NAND3_X2 U1500 ( .A1(n17510), .A2(n5807), .A3(n17511), .ZN(n17592) );
  AND3_X2 U7022 ( .A1(n4795), .A2(n5399), .A3(n16763), .ZN(n18441) );
  AND2_X2 U2528 ( .A1(n19987), .A2(n19988), .ZN(n20663) );
  BUF_X1 U3572 ( .A(n19795), .Z(n20261) );
  OR2_X2 U3562 ( .A1(n674), .A2(n23274), .ZN(n25008) );
  NAND2_X2 U1648 ( .A1(n689), .A2(n23944), .ZN(n25708) );
  OR2_X2 U16940 ( .A1(n10471), .A2(n10470), .ZN(n12339) );
  XNOR2_X2 U5184 ( .A(n15367), .B(n15368), .ZN(n17298) );
  NAND2_X2 U1222 ( .A1(n5550), .A2(n3719), .ZN(n19617) );
  BUF_X2 U618 ( .A(n11385), .Z(n12991) );
  INV_X2 U1569 ( .A(n18408), .ZN(n28798) );
  NAND2_X1 U82 ( .A1(n20739), .A2(n20737), .ZN(n21156) );
  XNOR2_X2 U11124 ( .A(n4989), .B(n5566), .ZN(n3880) );
  INV_X1 U10641 ( .A(n3829), .ZN(n11137) );
  INV_X2 U5413 ( .A(n5023), .ZN(n18709) );
  NOR2_X2 U2539 ( .A1(n18890), .A2(n18889), .ZN(n20988) );
  INV_X1 U19671 ( .A(n14921), .ZN(n16038) );
  BUF_X2 U1224 ( .A(n20013), .Z(n20510) );
  BUF_X2 U1622 ( .A(n27408), .Z(n28177) );
  OAI211_X2 U1416 ( .C1(n29228), .C2(n29227), .A(n29225), .B(n29224), .ZN(
        n22464) );
  BUF_X1 U4094 ( .A(n26682), .Z(n27434) );
  BUF_X1 U809 ( .A(n12955), .Z(n13218) );
  NAND2_X2 U1744 ( .A1(n28953), .A2(n28952), .ZN(n15127) );
  NAND2_X2 U18138 ( .A1(n14907), .A2(n14905), .ZN(n15098) );
  NAND3_X2 U3141 ( .A1(n9055), .A2(n9054), .A3(n9056), .ZN(n12200) );
  AND3_X2 U1672 ( .A1(n5445), .A2(n5444), .A3(n14515), .ZN(n15828) );
  MUX2_X2 U340 ( .A(n20297), .B(n20296), .S(n20295), .Z(n21308) );
  OAI21_X2 U7244 ( .B1(n22277), .B2(n23636), .A(n5457), .ZN(n22356) );
  NOR2_X2 U1002 ( .A1(n1339), .A2(n22014), .ZN(n22923) );
  BUF_X1 U15066 ( .A(n23633), .Z(n29061) );
  OR2_X2 U1519 ( .A1(n21275), .A2(n21283), .ZN(n21709) );
  OAI211_X2 U26 ( .C1(n6933), .C2(n4633), .A(n4632), .B(n4631), .ZN(n22882) );
  NAND2_X2 U1480 ( .A1(n20715), .A2(n20713), .ZN(n21591) );
  BUF_X1 U11677 ( .A(n26350), .Z(n28410) );
  BUF_X1 U2352 ( .A(n10008), .Z(n28616) );
  NAND2_X2 U2163 ( .A1(n11792), .A2(n28701), .ZN(n13020) );
  INV_X2 U2641 ( .A(n2571), .ZN(n19198) );
  NAND4_X1 U2361 ( .A1(n8986), .A2(n8985), .A3(n8988), .A4(n8987), .ZN(n10258)
         );
  NAND2_X2 U3354 ( .A1(n4695), .A2(n4698), .ZN(n9531) );
  AND2_X2 U1647 ( .A1(n28256), .A2(n28255), .ZN(n25509) );
  NOR2_X2 U1114 ( .A1(n27062), .A2(n27061), .ZN(n27905) );
  NAND3_X2 U9848 ( .A1(n15424), .A2(n15418), .A3(n15419), .ZN(n16569) );
  NAND2_X2 U956 ( .A1(n10899), .A2(n172), .ZN(n13101) );
  INV_X2 U3649 ( .A(n21657), .ZN(n6275) );
  NAND2_X2 U11637 ( .A1(n25359), .A2(n25357), .ZN(n27366) );
  MUX2_X2 U13179 ( .A(n26760), .B(n25276), .S(n26755), .Z(n25359) );
  XNOR2_X2 U796 ( .A(n22834), .B(n22833), .ZN(n23290) );
  AND2_X2 U1322 ( .A1(n5885), .A2(n5884), .ZN(n24631) );
  OAI21_X2 U1560 ( .B1(n15736), .B2(n15737), .A(n15735), .ZN(n19103) );
  OAI21_X1 U866 ( .B1(n14412), .B2(n14411), .A(n4001), .ZN(n14922) );
  OR2_X1 U6631 ( .A1(n2382), .A2(n7084), .ZN(n4675) );
  OAI21_X2 U2938 ( .B1(n13259), .B2(n14312), .A(n2331), .ZN(n14563) );
  NAND3_X2 U3830 ( .A1(n908), .A2(n4473), .A3(n907), .ZN(n24388) );
  OAI211_X2 U25124 ( .C1(n23510), .C2(n24081), .A(n23509), .B(n23508), .ZN(
        n25324) );
  MUX2_X2 U1638 ( .A(n8332), .B(n8331), .S(n8763), .Z(n10137) );
  XNOR2_X2 U1540 ( .A(n9945), .B(n9944), .ZN(n10461) );
  NAND3_X2 U1907 ( .A1(n15080), .A2(n15079), .A3(n28221), .ZN(n15865) );
  BUF_X1 U617 ( .A(n10657), .Z(n10872) );
  BUF_X2 U1083 ( .A(n23422), .Z(n23344) );
  NAND3_X2 U9543 ( .A1(n3051), .A2(n8750), .A3(n3050), .ZN(n10149) );
  XNOR2_X2 U3594 ( .A(n18742), .B(n18741), .ZN(n29114) );
  AND3_X2 U13051 ( .A1(n5749), .A2(n5750), .A3(n5748), .ZN(n25819) );
  XNOR2_X2 U3000 ( .A(n10772), .B(n10773), .ZN(n14107) );
  NAND2_X2 U2879 ( .A1(n11425), .A2(n11424), .ZN(n12420) );
  XNOR2_X2 U14814 ( .A(n7203), .B(Key[134]), .ZN(n7400) );
  AND3_X2 U102 ( .A1(n1597), .A2(n15130), .A3(n15129), .ZN(n3661) );
  AOI21_X1 U1491 ( .B1(n14183), .B2(n14470), .A(n5598), .ZN(n15165) );
  XNOR2_X2 U13203 ( .A(n6707), .B(n13927), .ZN(n5891) );
  OAI21_X1 U5292 ( .B1(n12452), .B2(n12451), .A(n1671), .ZN(n15097) );
  NAND2_X2 U931 ( .A1(n11987), .A2(n163), .ZN(n13543) );
  NAND2_X2 U11329 ( .A1(n10521), .A2(n4068), .ZN(n11449) );
  INV_X1 U3465 ( .A(n2984), .ZN(n624) );
  XNOR2_X1 U4478 ( .A(n26099), .B(n26098), .ZN(n27137) );
  NOR3_X1 U4475 ( .A1(n27147), .A2(n27142), .A3(n26858), .ZN(n27687) );
  OAI211_X2 U2885 ( .C1(n14690), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        n16238) );
  MUX2_X2 U24 ( .A(n20111), .B(n20110), .S(n20323), .Z(n20898) );
  CLKBUF_X3 U4355 ( .A(n9313), .Z(n9997) );
  BUF_X1 U362 ( .A(n18492), .Z(n28632) );
  BUF_X2 U1732 ( .A(n25059), .Z(n365) );
  BUF_X1 U1984 ( .A(n13595), .Z(n14372) );
  AOI22_X2 U26381 ( .A1(n26178), .A2(n26455), .B1(n25416), .B2(n25415), .ZN(
        n26830) );
  XNOR2_X2 U22103 ( .A(n18873), .B(n18872), .ZN(n20157) );
  NAND2_X2 U27041 ( .A1(n28712), .A2(n4242), .ZN(n22888) );
  INV_X1 U22730 ( .A(n19787), .ZN(n20635) );
  BUF_X1 U1124 ( .A(n24739), .Z(n29050) );
  MUX2_X2 U3086 ( .A(n12040), .B(n12039), .S(n375), .Z(n13171) );
  AOI21_X2 U9491 ( .B1(n23079), .B2(n23080), .A(n6580), .ZN(n23994) );
  NAND2_X2 U11723 ( .A1(n2314), .A2(n17122), .ZN(n17846) );
  OAI21_X2 U1142 ( .B1(n18844), .B2(n18843), .A(n18842), .ZN(n20816) );
  BUF_X1 U2816 ( .A(n17098), .Z(n17101) );
  AND2_X2 U1407 ( .A1(n23719), .A2(n23718), .ZN(n24517) );
  XNOR2_X2 U10604 ( .A(n7572), .B(n7573), .ZN(n11146) );
  INV_X1 U22633 ( .A(n19938), .ZN(n20281) );
  NAND3_X2 U12822 ( .A1(n13676), .A2(n13675), .A3(n5519), .ZN(n15388) );
  OAI211_X2 U943 ( .C1(n6785), .C2(n7618), .A(n3490), .B(n3489), .ZN(n329) );
  INV_X1 U1869 ( .A(n6309), .ZN(n24729) );
  OR2_X1 U10708 ( .A1(n7707), .A2(n371), .ZN(n4160) );
  BUF_X2 U1456 ( .A(n26507), .Z(n27084) );
  BUF_X1 U12305 ( .A(n23700), .Z(n28428) );
  AND3_X2 U182 ( .A1(n2072), .A2(n3474), .A3(n3475), .ZN(n22542) );
  NAND2_X2 U7564 ( .A1(n2552), .A2(n26844), .ZN(n27827) );
  INV_X1 U14609 ( .A(n7072), .ZN(n7886) );
  AOI21_X1 U4305 ( .B1(n20707), .B2(n20706), .A(n20705), .ZN(n22798) );
  NAND3_X2 U6191 ( .A1(n23895), .A2(n2265), .A3(n2266), .ZN(n25532) );
  NOR2_X1 U14436 ( .A1(n4466), .A2(n4465), .ZN(n22661) );
  AND3_X2 U5145 ( .A1(n1553), .A2(n1554), .A3(n5428), .ZN(n18263) );
  AND4_X2 U2566 ( .A1(n2177), .A2(n2179), .A3(n2082), .A4(n2182), .ZN(n21311)
         );
  AOI22_X2 U2871 ( .A1(n14820), .A2(n14819), .B1(n15444), .B2(n14818), .ZN(
        n16605) );
  NAND2_X2 U676 ( .A1(n20037), .A2(n3136), .ZN(n22023) );
  INV_X2 U6988 ( .A(n20225), .ZN(n20500) );
  XNOR2_X2 U21720 ( .A(n18385), .B(n18386), .ZN(n20290) );
  BUF_X2 U1715 ( .A(n20375), .Z(n351) );
  NAND3_X2 U5161 ( .A1(n8783), .A2(n9006), .A3(n1566), .ZN(n9716) );
  MUX2_X1 U6164 ( .A(n23548), .B(n23547), .S(n24772), .Z(n23549) );
  CLKBUF_X1 U1833 ( .A(Key[5]), .Z(n3219) );
  CLKBUF_X1 U1226 ( .A(Key[100]), .Z(n29247) );
  CLKBUF_X1 U1814 ( .A(Key[143]), .Z(n3049) );
  CLKBUF_X1 U51 ( .A(Key[183]), .Z(n3722) );
  CLKBUF_X1 U2113 ( .A(Key[102]), .Z(n26665) );
  CLKBUF_X1 U1832 ( .A(Key[6]), .Z(n3087) );
  XNOR2_X1 U14531 ( .A(Key[55]), .B(Plaintext[55]), .ZN(n7507) );
  CLKBUF_X1 U1230 ( .A(Key[0]), .Z(n1215) );
  XNOR2_X1 U5760 ( .A(Key[54]), .B(Plaintext[54]), .ZN(n7514) );
  CLKBUF_X1 U1235 ( .A(Key[175]), .Z(n3062) );
  XNOR2_X1 U3446 ( .A(Key[174]), .B(Plaintext[174]), .ZN(n7071) );
  XNOR2_X1 U14670 ( .A(Key[9]), .B(Plaintext[9]), .ZN(n7320) );
  XNOR2_X1 U14450 ( .A(Key[98]), .B(Plaintext[98]), .ZN(n7363) );
  XNOR2_X1 U14418 ( .A(Key[112]), .B(Plaintext[112]), .ZN(n8213) );
  XNOR2_X1 U933 ( .A(Key[182]), .B(Plaintext[182]), .ZN(n7092) );
  XNOR2_X1 U675 ( .A(n7098), .B(Key[17]), .ZN(n7759) );
  INV_X1 U16341 ( .A(n1196), .ZN(n24906) );
  XNOR2_X1 U247 ( .A(n6972), .B(Key[102]), .ZN(n8232) );
  XNOR2_X1 U14590 ( .A(n7057), .B(Key[166]), .ZN(n7999) );
  XNOR2_X1 U14568 ( .A(n7045), .B(Key[157]), .ZN(n7965) );
  XNOR2_X1 U14598 ( .A(n7062), .B(Key[162]), .ZN(n7992) );
  XNOR2_X1 U14699 ( .A(n7128), .B(Key[46]), .ZN(n8131) );
  XNOR2_X1 U14469 ( .A(n6995), .B(Key[120]), .ZN(n7628) );
  BUF_X1 U132 ( .A(n7110), .Z(n7898) );
  XNOR2_X1 U14542 ( .A(n7028), .B(Key[64]), .ZN(n7521) );
  BUF_X1 U3414 ( .A(n8290), .Z(n7915) );
  XNOR2_X1 U2413 ( .A(n7016), .B(Key[88]), .ZN(n7837) );
  BUF_X1 U3403 ( .A(n7404), .Z(n7976) );
  OR2_X1 U781 ( .A1(n7324), .A2(n7325), .ZN(n8579) );
  NAND3_X1 U694 ( .A1(n7951), .A2(n7950), .A3(n117), .ZN(n9107) );
  OR2_X1 U4546 ( .A1(n8026), .A2(n8025), .ZN(n8899) );
  MUX2_X1 U2453 ( .A(n7762), .B(n7761), .S(n7760), .Z(n7765) );
  OR2_X1 U1377 ( .A1(n7944), .A2(n7945), .ZN(n8914) );
  NAND2_X1 U4183 ( .A1(n7772), .A2(n3183), .ZN(n8351) );
  OAI21_X1 U680 ( .B1(n7152), .B2(n8148), .A(n7151), .ZN(n9247) );
  OR2_X1 U3388 ( .A1(n7429), .A2(n7428), .ZN(n9075) );
  OAI21_X1 U14453 ( .B1(n6983), .B2(n6982), .A(n6981), .ZN(n9229) );
  NAND3_X1 U665 ( .A1(n3185), .A2(n2221), .A3(n2222), .ZN(n8502) );
  NAND3_X1 U4505 ( .A1(n6802), .A2(n6801), .A3(n7593), .ZN(n8414) );
  OAI211_X1 U15204 ( .C1(n7732), .C2(n7733), .A(n7731), .B(n7730), .ZN(n9186)
         );
  NAND2_X1 U3348 ( .A1(n8152), .A2(n1512), .ZN(n8983) );
  OR2_X1 U1167 ( .A1(n7599), .A2(n7598), .ZN(n8788) );
  OR2_X1 U1065 ( .A1(n7713), .A2(n7712), .ZN(n9029) );
  OAI211_X1 U1442 ( .C1(n7673), .C2(n8275), .A(n7672), .B(n7671), .ZN(n8996)
         );
  OR2_X1 U1349 ( .A1(n2506), .A2(n7131), .ZN(n9041) );
  NOR2_X1 U1586 ( .A1(n3445), .A2(n155), .ZN(n28606) );
  BUF_X1 U1549 ( .A(n7726), .Z(n9188) );
  OR2_X1 U861 ( .A1(n732), .A2(n7739), .ZN(n8782) );
  AND2_X1 U410 ( .A1(n7904), .A2(n7903), .ZN(n8635) );
  NAND2_X1 U3343 ( .A1(n7972), .A2(n7973), .ZN(n8665) );
  MUX2_X1 U159 ( .A(n7217), .B(n7214), .S(n29673), .Z(n9228) );
  NAND2_X1 U8448 ( .A1(n2424), .A2(n2059), .ZN(n8719) );
  NAND2_X1 U654 ( .A1(n6199), .A2(n7242), .ZN(n8608) );
  BUF_X1 U1098 ( .A(n7175), .Z(n8537) );
  AND2_X1 U3333 ( .A1(n1042), .A2(n7195), .ZN(n8685) );
  AND2_X1 U3366 ( .A1(n7558), .A2(n7559), .ZN(n8872) );
  OR2_X1 U8480 ( .A1(n8785), .A2(n8414), .ZN(n8438) );
  OR2_X1 U6238 ( .A1(n9063), .A2(n9062), .ZN(n5536) );
  OR2_X1 U86 ( .A1(n8943), .A2(n8944), .ZN(n2168) );
  NAND3_X1 U910 ( .A1(n8489), .A2(n6318), .A3(n6317), .ZN(n10386) );
  MUX2_X1 U8663 ( .A(n8437), .B(n8436), .S(n9210), .Z(n9735) );
  OR2_X1 U15739 ( .A1(n8646), .A2(n8762), .ZN(n10406) );
  OR2_X1 U834 ( .A1(n9011), .A2(n9010), .ZN(n9512) );
  OR2_X1 U533 ( .A1(n9341), .A2(n2229), .ZN(n9979) );
  OR2_X1 U868 ( .A1(n8895), .A2(n8894), .ZN(n9824) );
  AND3_X1 U136 ( .A1(n2247), .A2(n3755), .A3(n28882), .ZN(n9648) );
  OR2_X1 U5888 ( .A1(n127), .A2(n8713), .ZN(n9575) );
  NAND2_X1 U556 ( .A1(n9415), .A2(n9414), .ZN(n10392) );
  MUX2_X1 U5623 ( .A(n8442), .B(n8441), .S(n8440), .Z(n1920) );
  OR2_X1 U15283 ( .A1(n7956), .A2(n7955), .ZN(n10357) );
  NAND3_X1 U3276 ( .A1(n3182), .A2(n8841), .A3(n3181), .ZN(n10272) );
  NAND2_X1 U9258 ( .A1(n8618), .A2(n2907), .ZN(n10043) );
  OR2_X1 U3291 ( .A1(n5308), .A2(n8645), .ZN(n10184) );
  OAI21_X1 U2564 ( .B1(n8662), .B2(n5677), .A(n5673), .ZN(n10134) );
  OAI211_X1 U740 ( .C1(n9227), .C2(n9228), .A(n9225), .B(n9226), .ZN(n10335)
         );
  XNOR2_X1 U15807 ( .A(n9295), .B(n26656), .ZN(n8772) );
  OAI21_X1 U4121 ( .B1(n8356), .B2(n8431), .A(n971), .ZN(n10282) );
  XNOR2_X1 U5645 ( .A(n10321), .B(n2845), .ZN(n9770) );
  NAND2_X1 U3267 ( .A1(n2334), .A2(n2336), .ZN(n10294) );
  NAND3_X1 U3274 ( .A1(n8387), .A2(n8386), .A3(n8385), .ZN(n10074) );
  NAND2_X1 U10996 ( .A1(n3781), .A2(n3780), .ZN(n10208) );
  OAI21_X1 U1448 ( .B1(n29147), .B2(n8198), .A(n8197), .ZN(n10060) );
  XNOR2_X1 U2143 ( .A(n9908), .B(n10021), .ZN(n10319) );
  XNOR2_X1 U516 ( .A(n9916), .B(n9698), .ZN(n10342) );
  XNOR2_X1 U16058 ( .A(n9280), .B(n9279), .ZN(n10705) );
  XNOR2_X1 U2333 ( .A(n5401), .B(n5400), .ZN(n11135) );
  XNOR2_X1 U16011 ( .A(n9217), .B(n9216), .ZN(n11349) );
  XNOR2_X1 U1667 ( .A(n9651), .B(n9652), .ZN(n11267) );
  XNOR2_X1 U3220 ( .A(n9159), .B(n9158), .ZN(n10847) );
  XNOR2_X1 U451 ( .A(n9898), .B(n9897), .ZN(n11120) );
  XNOR2_X1 U3217 ( .A(n10378), .B(n10377), .ZN(n11281) );
  BUF_X1 U269 ( .A(n10096), .Z(n29150) );
  XNOR2_X1 U3189 ( .A(n3437), .B(n5860), .ZN(n10958) );
  XNOR2_X1 U217 ( .A(n9792), .B(n9791), .ZN(n10995) );
  XNOR2_X1 U1338 ( .A(n5562), .B(n10286), .ZN(n11290) );
  OR2_X1 U9884 ( .A1(n11237), .A2(n11010), .ZN(n11234) );
  XNOR2_X1 U669 ( .A(n4590), .B(n4589), .ZN(n11165) );
  XNOR2_X1 U3200 ( .A(n9361), .B(n9360), .ZN(n10962) );
  BUF_X2 U1000 ( .A(n11064), .Z(n11069) );
  XNOR2_X1 U198 ( .A(n9328), .B(n9327), .ZN(n10913) );
  BUF_X1 U7569 ( .A(n10097), .Z(n11114) );
  NOR2_X1 U2665 ( .A1(n11199), .A2(n28207), .ZN(n10749) );
  BUF_X1 U3201 ( .A(n10855), .Z(n11308) );
  OAI211_X1 U17250 ( .C1(n10989), .C2(n10988), .A(n10987), .B(n10986), .ZN(
        n12249) );
  MUX2_X1 U3164 ( .A(n10631), .B(n9848), .S(n10783), .Z(n9865) );
  OR2_X1 U17119 ( .A1(n10737), .A2(n10736), .ZN(n11426) );
  NAND2_X1 U860 ( .A1(n3165), .A2(n10092), .ZN(n10905) );
  NAND3_X1 U6206 ( .A1(n1080), .A2(n10633), .A3(n10634), .ZN(n12218) );
  AOI22_X1 U3158 ( .A1(n11224), .A2(n11223), .B1(n11222), .B2(n11221), .ZN(
        n12320) );
  OAI211_X1 U2006 ( .C1(n10822), .C2(n28208), .A(n10824), .B(n6885), .ZN(
        n12146) );
  NAND2_X1 U4145 ( .A1(n1214), .A2(n3018), .ZN(n12058) );
  AND3_X1 U1587 ( .A1(n10217), .A2(n10216), .A3(n10215), .ZN(n11824) );
  AND2_X1 U4024 ( .A1(n898), .A2(n1146), .ZN(n12271) );
  OR2_X1 U2140 ( .A1(n10762), .A2(n6918), .ZN(n11405) );
  OR2_X1 U838 ( .A1(n10654), .A2(n10653), .ZN(n1986) );
  NOR2_X1 U2875 ( .A1(n11636), .A2(n11633), .ZN(n29139) );
  OAI21_X1 U4349 ( .B1(n4815), .B2(n4325), .A(n4328), .ZN(n12156) );
  AND3_X1 U1487 ( .A1(n3815), .A2(n4800), .A3(n3814), .ZN(n12111) );
  OR2_X1 U745 ( .A1(n11660), .A2(n10895), .ZN(n11377) );
  NAND3_X1 U717 ( .A1(n4710), .A2(n10511), .A3(n6271), .ZN(n11500) );
  NAND2_X1 U229 ( .A1(n28282), .A2(n28283), .ZN(n6482) );
  NAND3_X1 U7444 ( .A1(n3373), .A2(n8623), .A3(n8622), .ZN(n12203) );
  INV_X1 U13632 ( .A(n11794), .ZN(n10717) );
  AND3_X1 U1797 ( .A1(n2943), .A2(n11102), .A3(n1945), .ZN(n12516) );
  BUF_X1 U3112 ( .A(n11390), .Z(n11851) );
  NAND2_X1 U5451 ( .A1(n1786), .A2(n1787), .ZN(n12251) );
  AND2_X1 U187 ( .A1(n11495), .A2(n11493), .ZN(n569) );
  BUF_X1 U55 ( .A(n11878), .Z(n287) );
  NAND2_X1 U17867 ( .A1(n12198), .A2(n12189), .ZN(n12131) );
  BUF_X1 U5971 ( .A(n11859), .Z(n11943) );
  BUF_X1 U7578 ( .A(n12307), .Z(n4197) );
  NAND2_X1 U4540 ( .A1(n10604), .A2(n3322), .ZN(n12356) );
  INV_X1 U6298 ( .A(n12307), .ZN(n12300) );
  OR2_X1 U11157 ( .A1(n3910), .A2(n3908), .ZN(n4341) );
  INV_X1 U7445 ( .A(n12203), .ZN(n4844) );
  INV_X1 U3125 ( .A(n11058), .ZN(n12267) );
  BUF_X1 U652 ( .A(n11505), .Z(n12400) );
  BUF_X1 U3127 ( .A(n11419), .Z(n11785) );
  BUF_X1 U16436 ( .A(n9692), .Z(n12109) );
  NAND2_X1 U5761 ( .A1(n11887), .A2(n11886), .ZN(n12327) );
  OR2_X1 U6287 ( .A1(n11622), .A2(n11194), .ZN(n11580) );
  MUX2_X1 U10185 ( .A(n10118), .B(n10117), .S(n12507), .Z(n13167) );
  NAND3_X1 U10906 ( .A1(n11909), .A2(n28962), .A3(n28961), .ZN(n13413) );
  NAND3_X1 U1095 ( .A1(n11573), .A2(n11572), .A3(n3745), .ZN(n13291) );
  AND2_X1 U1169 ( .A1(n3795), .A2(n3794), .ZN(n13493) );
  OAI211_X1 U5628 ( .C1(n11485), .C2(n11484), .A(n11483), .B(n11612), .ZN(
        n13244) );
  NOR2_X1 U20964 ( .A1(n12185), .A2(n12184), .ZN(n13261) );
  OAI211_X1 U1190 ( .C1(n11711), .C2(n5169), .A(n3688), .B(n11414), .ZN(n12723) );
  OAI21_X1 U590 ( .B1(n12225), .B2(n12224), .A(n12223), .ZN(n13285) );
  AND2_X1 U12374 ( .A1(n5096), .A2(n5095), .ZN(n13236) );
  NAND2_X1 U2954 ( .A1(n11475), .A2(n3592), .ZN(n13018) );
  OAI21_X1 U13713 ( .B1(n6481), .B2(n6478), .A(n11721), .ZN(n13067) );
  NAND2_X1 U1265 ( .A1(n3566), .A2(n233), .ZN(n13159) );
  XNOR2_X1 U3056 ( .A(n13166), .B(n13219), .ZN(n13522) );
  BUF_X1 U1307 ( .A(n12752), .Z(n12783) );
  OAI21_X1 U1100 ( .B1(n1401), .B2(n12431), .A(n12430), .ZN(n13369) );
  XNOR2_X1 U8956 ( .A(n13523), .B(n1885), .ZN(n12454) );
  NAND2_X1 U1846 ( .A1(n10651), .A2(n10650), .ZN(n12560) );
  XNOR2_X1 U759 ( .A(n12719), .B(n12720), .ZN(n13933) );
  XNOR2_X1 U3031 ( .A(n12970), .B(n12969), .ZN(n14091) );
  XNOR2_X1 U817 ( .A(n12476), .B(n12477), .ZN(n12480) );
  XNOR2_X1 U1288 ( .A(n12540), .B(n12539), .ZN(n14426) );
  XNOR2_X1 U18060 ( .A(n12463), .B(n12464), .ZN(n14217) );
  BUF_X1 U3034 ( .A(n13755), .Z(n14475) );
  XNOR2_X1 U3036 ( .A(n12139), .B(n12138), .ZN(n14166) );
  XNOR2_X1 U3001 ( .A(n2962), .B(n3110), .ZN(n14435) );
  BUF_X1 U91 ( .A(n13749), .Z(n14261) );
  XNOR2_X1 U3009 ( .A(n13065), .B(n13064), .ZN(n14351) );
  XNOR2_X1 U994 ( .A(n12984), .B(n12983), .ZN(n14358) );
  BUF_X1 U1308 ( .A(n13686), .Z(n14415) );
  XNOR2_X1 U758 ( .A(n2173), .B(n2171), .ZN(n14376) );
  OAI21_X1 U2978 ( .B1(n13696), .B2(n13656), .A(n13655), .ZN(n14743) );
  OR2_X1 U972 ( .A1(n14042), .A2(n14041), .ZN(n14600) );
  OAI21_X1 U18988 ( .B1(n13696), .B2(n14325), .A(n13695), .ZN(n14115) );
  MUX2_X1 U10527 ( .A(n13165), .B(n13164), .S(n14328), .Z(n15692) );
  NAND3_X1 U23940 ( .A1(n1345), .A2(n14329), .A3(n1344), .ZN(n15306) );
  NOR2_X1 U751 ( .A1(n13665), .A2(n2373), .ZN(n14514) );
  INV_X1 U2961 ( .A(n14115), .ZN(n15138) );
  AND2_X1 U1361 ( .A1(n13905), .A2(n13904), .ZN(n14807) );
  NAND3_X1 U28161 ( .A1(n28754), .A2(n1016), .A3(n28753), .ZN(n14773) );
  INV_X1 U3187 ( .A(n14600), .ZN(n14601) );
  AND2_X1 U2955 ( .A1(n4163), .A2(n14277), .ZN(n14763) );
  OR2_X1 U2973 ( .A1(n14378), .A2(n14377), .ZN(n15511) );
  AND3_X1 U1743 ( .A1(n12758), .A2(n14471), .A3(n28936), .ZN(n15101) );
  OR2_X1 U225 ( .A1(n6446), .A2(n13590), .ZN(n15400) );
  AOI22_X1 U2969 ( .A1(n13746), .A2(n13745), .B1(n14076), .B2(n4376), .ZN(
        n15383) );
  OAI211_X1 U1642 ( .C1(n14009), .C2(n5404), .A(n6614), .B(n6613), .ZN(n14826)
         );
  AND2_X1 U226 ( .A1(n14830), .A2(n14834), .ZN(n15292) );
  NAND2_X1 U5803 ( .A1(n13705), .A2(n3435), .ZN(n15250) );
  NAND2_X1 U9541 ( .A1(n1627), .A2(n14472), .ZN(n15491) );
  OR2_X1 U11705 ( .A1(n13979), .A2(n14743), .ZN(n14744) );
  NOR2_X1 U18975 ( .A1(n14990), .A2(n14989), .ZN(n15395) );
  AOI21_X1 U1162 ( .B1(n5823), .B2(n293), .A(n5820), .ZN(n14986) );
  OAI21_X1 U6391 ( .B1(n5834), .B2(n13336), .A(n28866), .ZN(n14882) );
  NOR2_X1 U3081 ( .A1(n13596), .A2(n13597), .ZN(n13638) );
  NAND2_X1 U876 ( .A1(n2562), .A2(n2561), .ZN(n15174) );
  INV_X2 U6901 ( .A(n15311), .ZN(n14851) );
  BUF_X1 U2915 ( .A(n14518), .Z(n15036) );
  INV_X1 U895 ( .A(n14518), .ZN(n3827) );
  INV_X1 U4766 ( .A(n14575), .ZN(n15105) );
  NOR2_X1 U3120 ( .A1(n3208), .A2(n15387), .ZN(n14994) );
  OAI211_X1 U15633 ( .C1(n14968), .C2(n14961), .A(n13787), .B(n13786), .ZN(
        n16284) );
  OR2_X1 U1492 ( .A1(n15495), .A2(n15491), .ZN(n264) );
  AND3_X1 U1710 ( .A1(n29173), .A2(n29172), .A3(n29171), .ZN(n16634) );
  NAND2_X1 U537 ( .A1(n88), .A2(n14794), .ZN(n16509) );
  AND4_X1 U892 ( .A1(n5052), .A2(n5051), .A3(n14919), .A4(n5050), .ZN(n15977)
         );
  NOR2_X1 U2881 ( .A1(n14828), .A2(n14829), .ZN(n16526) );
  NAND2_X1 U621 ( .A1(n3682), .A2(n15364), .ZN(n16230) );
  NAND2_X1 U9696 ( .A1(n15220), .A2(n15221), .ZN(n15642) );
  NAND2_X1 U4770 ( .A1(n15270), .A2(n1243), .ZN(n16242) );
  AOI21_X1 U3900 ( .B1(n13978), .B2(n15014), .A(n13977), .ZN(n16146) );
  OR2_X1 U2877 ( .A1(n4720), .A2(n4718), .ZN(n15618) );
  AND2_X1 U1688 ( .A1(n14626), .A2(n14627), .ZN(n16043) );
  OR2_X1 U1264 ( .A1(n15149), .A2(n15148), .ZN(n16051) );
  NAND3_X1 U1690 ( .A1(n28837), .A2(n15240), .A3(n2885), .ZN(n16105) );
  NAND3_X1 U10506 ( .A1(n4417), .A2(n3550), .A3(n14599), .ZN(n16233) );
  NAND2_X1 U509 ( .A1(n82), .A2(n1964), .ZN(n16589) );
  XNOR2_X1 U1683 ( .A(n15846), .B(n15845), .ZN(n16908) );
  XNOR2_X1 U1960 ( .A(n14720), .B(n14721), .ZN(n17393) );
  XNOR2_X1 U2823 ( .A(n16573), .B(n16572), .ZN(n17516) );
  BUF_X1 U67 ( .A(n15551), .Z(n17348) );
  XNOR2_X1 U1243 ( .A(n15684), .B(n15683), .ZN(n17548) );
  XNOR2_X1 U19897 ( .A(n15429), .B(n15428), .ZN(n17411) );
  XNOR2_X1 U2839 ( .A(n15913), .B(n15912), .ZN(n17572) );
  XNOR2_X1 U10567 ( .A(n16515), .B(n16516), .ZN(n17450) );
  XNOR2_X1 U595 ( .A(n15776), .B(n15775), .ZN(n17543) );
  XNOR2_X1 U713 ( .A(n16195), .B(n16194), .ZN(n16888) );
  BUF_X1 U1650 ( .A(n17466), .Z(n28800) );
  XNOR2_X1 U10409 ( .A(n6502), .B(n16380), .ZN(n17375) );
  INV_X1 U2810 ( .A(n4316), .ZN(n17229) );
  BUF_X1 U1273 ( .A(n16137), .Z(n17262) );
  BUF_X1 U3149 ( .A(n16837), .Z(n17562) );
  MUX2_X1 U10593 ( .A(n16905), .B(n17706), .S(n4156), .Z(n18268) );
  OAI21_X1 U3287 ( .B1(n17194), .B2(n5260), .A(n17193), .ZN(n18121) );
  AOI22_X1 U26675 ( .A1(n3169), .A2(n3172), .B1(n16725), .B2(n16660), .ZN(
        n16663) );
  MUX2_X1 U616 ( .A(n16886), .B(n16885), .S(n17158), .Z(n18516) );
  INV_X1 U2769 ( .A(n19562), .ZN(n527) );
  OR2_X1 U4223 ( .A1(n16688), .A2(n16689), .ZN(n18342) );
  NAND2_X1 U1844 ( .A1(n14507), .A2(n17009), .ZN(n18306) );
  AND3_X1 U2731 ( .A1(n16979), .A2(n6538), .A3(n16978), .ZN(n18081) );
  OAI21_X1 U1614 ( .B1(n17161), .B2(n17386), .A(n28851), .ZN(n18376) );
  NAND3_X1 U473 ( .A1(n4702), .A2(n4700), .A3(n4699), .ZN(n18276) );
  AND3_X1 U6121 ( .A1(n3811), .A2(n3812), .A3(n5620), .ZN(n18356) );
  OR2_X1 U1943 ( .A1(n17144), .A2(n17145), .ZN(n5383) );
  NAND2_X1 U4793 ( .A1(n1264), .A2(n16692), .ZN(n18344) );
  NAND2_X1 U457 ( .A1(n5250), .A2(n783), .ZN(n17969) );
  OR2_X1 U56 ( .A1(n17306), .A2(n17307), .ZN(n17620) );
  BUF_X1 U1242 ( .A(n17826), .Z(n18160) );
  NAND2_X1 U27347 ( .A1(n6175), .A2(n6176), .ZN(n18527) );
  NAND2_X1 U27746 ( .A1(n28728), .A2(n1367), .ZN(n16985) );
  AND2_X1 U2719 ( .A1(n2702), .A2(n4280), .ZN(n18260) );
  AND2_X1 U1619 ( .A1(n29240), .A2(n4040), .ZN(n18248) );
  BUF_X1 U1753 ( .A(n18522), .Z(n373) );
  AND2_X1 U9048 ( .A1(n5326), .A2(n5327), .ZN(n18286) );
  NOR2_X1 U6979 ( .A1(n18298), .A2(n18063), .ZN(n2791) );
  INV_X1 U78 ( .A(n17207), .ZN(n17835) );
  OR2_X1 U100 ( .A1(n18304), .A2(n17679), .ZN(n18012) );
  AOI21_X1 U21364 ( .B1(n16898), .B2(n18276), .A(n18279), .ZN(n18206) );
  NAND2_X1 U2677 ( .A1(n16901), .A2(n16900), .ZN(n19111) );
  OAI211_X1 U884 ( .C1(n18163), .C2(n18164), .A(n18162), .B(n18161), .ZN(
        n19678) );
  OAI21_X1 U2681 ( .B1(n6326), .B2(n18454), .A(n18453), .ZN(n19220) );
  NAND2_X1 U351 ( .A1(n40), .A2(n18287), .ZN(n19695) );
  NAND2_X1 U1220 ( .A1(n2214), .A2(n2212), .ZN(n18638) );
  NAND2_X1 U2643 ( .A1(n2566), .A2(n17841), .ZN(n19704) );
  NAND2_X1 U1760 ( .A1(n28733), .A2(n17648), .ZN(n19108) );
  OAI21_X1 U1713 ( .B1(n18359), .B2(n18360), .A(n18358), .ZN(n18798) );
  AND2_X1 U1051 ( .A1(n1784), .A2(n17981), .ZN(n18959) );
  XNOR2_X1 U21921 ( .A(n19111), .B(n2889), .ZN(n18671) );
  XNOR2_X1 U21441 ( .A(n28447), .B(n19706), .ZN(n19285) );
  INV_X1 U6079 ( .A(n18867), .ZN(n19087) );
  NAND2_X1 U4051 ( .A1(n916), .A2(n913), .ZN(n19697) );
  XNOR2_X1 U22429 ( .A(n19312), .B(n19311), .ZN(n20626) );
  XNOR2_X1 U9673 ( .A(n19264), .B(n3111), .ZN(n20601) );
  XNOR2_X1 U1341 ( .A(n19684), .B(n19683), .ZN(n20607) );
  XNOR2_X1 U468 ( .A(n19722), .B(n19721), .ZN(n20614) );
  XNOR2_X1 U303 ( .A(n19494), .B(n19493), .ZN(n20444) );
  XNOR2_X1 U9769 ( .A(n18771), .B(n19455), .ZN(n20063) );
  BUF_X1 U1922 ( .A(n19995), .Z(n20478) );
  BUF_X1 U773 ( .A(n28140), .Z(n28779) );
  BUF_X1 U273 ( .A(n20224), .Z(n297) );
  BUF_X1 U8041 ( .A(n17954), .Z(n20311) );
  BUF_X1 U4723 ( .A(n19928), .Z(n20449) );
  NOR3_X1 U3608 ( .A1(n20545), .A2(n20546), .A3(n20547), .ZN(n21585) );
  MUX2_X1 U690 ( .A(n20543), .B(n20542), .S(n20541), .Z(n21586) );
  AND2_X1 U3516 ( .A1(n5302), .A2(n5305), .ZN(n21047) );
  OAI21_X1 U534 ( .B1(n20411), .B2(n20410), .A(n20409), .ZN(n21503) );
  OAI21_X1 U25346 ( .B1(n18833), .B2(n20097), .A(n28326), .ZN(n20878) );
  BUF_X1 U7131 ( .A(n20722), .Z(n21598) );
  BUF_X2 U23326 ( .A(n20782), .Z(n21551) );
  OR2_X1 U252 ( .A1(n20254), .A2(n28295), .ZN(n21014) );
  AND2_X1 U2553 ( .A1(n2747), .A2(n5376), .ZN(n21534) );
  AND3_X1 U593 ( .A1(n20566), .A2(n20564), .A3(n20565), .ZN(n5684) );
  MUX2_X1 U1916 ( .A(n19742), .B(n19741), .S(n19740), .Z(n22140) );
  NAND3_X1 U4621 ( .A1(n19853), .A2(n19854), .A3(n19852), .ZN(n21574) );
  OR2_X1 U1910 ( .A1(n19998), .A2(n6028), .ZN(n21171) );
  NOR2_X1 U419 ( .A1(n1099), .A2(n1335), .ZN(n20783) );
  OR2_X1 U19739 ( .A1(n28662), .A2(n28661), .ZN(n28584) );
  NAND3_X1 U1913 ( .A1(n20004), .A2(n6137), .A3(n20003), .ZN(n21408) );
  OR2_X1 U2484 ( .A1(n1327), .A2(n21749), .ZN(n5975) );
  NOR2_X1 U22532 ( .A1(n19459), .A2(n19458), .ZN(n21717) );
  OR2_X1 U1773 ( .A1(n21645), .A2(n497), .ZN(n21237) );
  OAI21_X1 U2483 ( .B1(n21685), .B2(n21684), .A(n21683), .ZN(n22221) );
  AOI21_X1 U10007 ( .B1(n21405), .B2(n21404), .A(n21403), .ZN(n22411) );
  MUX2_X1 U7087 ( .A(n18549), .B(n18548), .S(n28440), .Z(n21825) );
  OAI21_X1 U588 ( .B1(n20364), .B2(n20365), .A(n20363), .ZN(n22472) );
  NAND2_X1 U10079 ( .A1(n21201), .A2(n3288), .ZN(n22854) );
  AND2_X1 U2474 ( .A1(n1084), .A2(n1083), .ZN(n22414) );
  AND3_X1 U2475 ( .A1(n6694), .A2(n6695), .A3(n6696), .ZN(n22437) );
  AND4_X1 U761 ( .A1(n21486), .A2(n21488), .A3(n6369), .A4(n21487), .ZN(n22337) );
  NAND3_X1 U927 ( .A1(n6350), .A2(n21444), .A3(n6349), .ZN(n22479) );
  AOI21_X1 U1423 ( .B1(n21214), .B2(n21213), .A(n872), .ZN(n22783) );
  NOR2_X1 U218 ( .A1(n18788), .A2(n18787), .ZN(n2805) );
  NAND2_X1 U1585 ( .A1(n21285), .A2(n21284), .ZN(n22501) );
  AND3_X1 U1538 ( .A1(n6041), .A2(n6040), .A3(n6039), .ZN(n22710) );
  OAI211_X1 U5415 ( .C1(n20530), .C2(n20531), .A(n20529), .B(n20528), .ZN(
        n22750) );
  NAND2_X1 U1901 ( .A1(n2991), .A2(n2988), .ZN(n22525) );
  XNOR2_X1 U145 ( .A(n21948), .B(n274), .ZN(n23606) );
  XNOR2_X1 U1178 ( .A(n4760), .B(n21803), .ZN(n23769) );
  XNOR2_X1 U3913 ( .A(n22385), .B(n22384), .ZN(n23566) );
  XNOR2_X1 U908 ( .A(n21968), .B(n21969), .ZN(n23607) );
  XNOR2_X1 U1706 ( .A(n22005), .B(n22004), .ZN(n2141) );
  XNOR2_X1 U13805 ( .A(n22795), .B(n22794), .ZN(n23416) );
  BUF_X1 U13034 ( .A(n23297), .Z(n29020) );
  BUF_X1 U1513 ( .A(n22946), .Z(n23741) );
  BUF_X1 U2400 ( .A(n23233), .Z(n23714) );
  BUF_X1 U224 ( .A(n23280), .Z(n28418) );
  OR2_X1 U1677 ( .A1(n23088), .A2(n23087), .ZN(n24378) );
  NAND2_X1 U901 ( .A1(n22176), .A2(n22175), .ZN(n24582) );
  OR2_X1 U777 ( .A1(n5346), .A2(n23208), .ZN(n138) );
  OAI21_X1 U13361 ( .B1(n22129), .B2(n28474), .A(n22128), .ZN(n29026) );
  NAND3_X1 U9865 ( .A1(n6764), .A2(n6763), .A3(n1965), .ZN(n24391) );
  OR2_X1 U2351 ( .A1(n2835), .A2(n2076), .ZN(n24800) );
  NAND2_X1 U271 ( .A1(n1446), .A2(n28695), .ZN(n24081) );
  OAI211_X1 U1334 ( .C1(n23035), .C2(n23034), .A(n4935), .B(n4934), .ZN(n29043) );
  NAND2_X1 U1662 ( .A1(n5456), .A2(n28224), .ZN(n24602) );
  AND2_X1 U9787 ( .A1(n2818), .A2(n2817), .ZN(n24420) );
  AND2_X1 U26111 ( .A1(n23730), .A2(n23731), .ZN(n24520) );
  BUF_X1 U14362 ( .A(n23932), .Z(n24597) );
  BUF_X1 U435 ( .A(n25908), .Z(n28769) );
  AOI21_X1 U14356 ( .B1(n23975), .B2(n23974), .A(n23973), .ZN(n25187) );
  AND2_X1 U1389 ( .A1(n964), .A2(n967), .ZN(n26100) );
  OAI211_X1 U207 ( .C1(n4749), .C2(n4748), .A(n24147), .B(n24148), .ZN(n26093)
         );
  XNOR2_X1 U1473 ( .A(n25111), .B(n25110), .ZN(n26800) );
  XNOR2_X1 U2260 ( .A(n25707), .B(n25706), .ZN(n27069) );
  AND2_X1 U6580 ( .A1(n26865), .A2(n27110), .ZN(n27152) );
  MUX2_X1 U27064 ( .A(n26351), .B(n26350), .S(n27701), .Z(n26355) );
  AND2_X1 U26887 ( .A1(n26128), .A2(n27161), .ZN(n27707) );
  OAI21_X1 U10327 ( .B1(n26365), .B2(n28948), .A(n26363), .ZN(n27632) );
  NAND2_X1 U1221 ( .A1(n2966), .A2(n26564), .ZN(n27496) );
  NAND2_X1 U16604 ( .A1(n26243), .A2(n26244), .ZN(n28543) );
  CLKBUF_X1 U1238 ( .A(Key[153]), .Z(n3537) );
  XNOR2_X1 U14692 ( .A(Key[43]), .B(Plaintext[43]), .ZN(n8048) );
  BUF_X1 U4207 ( .A(Key[161]), .Z(n3787) );
  BUF_X1 U2473 ( .A(Key[134]), .Z(n28693) );
  BUF_X1 U3497 ( .A(Key[70]), .Z(n3036) );
  BUF_X1 U2063 ( .A(Key[79]), .Z(n26214) );
  BUF_X1 U1829 ( .A(Key[131]), .Z(n3491) );
  BUF_X2 U1604 ( .A(Key[186]), .Z(n3015) );
  CLKBUF_X1 U4208 ( .A(Key[162]), .Z(n3196) );
  OR2_X1 U8405 ( .A1(n2406), .A2(n6999), .ZN(n9045) );
  OR2_X1 U1205 ( .A1(n7339), .A2(n7338), .ZN(n9144) );
  NOR2_X1 U2227 ( .A1(n7661), .A2(n28857), .ZN(n8995) );
  INV_X1 U3387 ( .A(n29303), .ZN(n610) );
  OR2_X1 U11936 ( .A1(n4671), .A2(n7319), .ZN(n8327) );
  NAND2_X1 U157 ( .A1(n3179), .A2(n7617), .ZN(n9196) );
  BUF_X1 U124 ( .A(n9363), .Z(n284) );
  INV_X1 U3325 ( .A(n8384), .ZN(n8739) );
  NAND2_X1 U2379 ( .A1(n28751), .A2(n2480), .ZN(n8741) );
  NAND2_X1 U14462 ( .A1(n7482), .A2(n7483), .ZN(n28500) );
  OAI211_X1 U5458 ( .C1(n1792), .C2(n1794), .A(n1789), .B(n2844), .ZN(n9696)
         );
  OAI211_X1 U1367 ( .C1(n9169), .C2(n8250), .A(n8249), .B(n8248), .ZN(n10178)
         );
  OAI21_X1 U517 ( .B1(n2713), .B2(n8339), .A(n2712), .ZN(n9698) );
  NAND2_X1 U643 ( .A1(n5867), .A2(n3678), .ZN(n9991) );
  NAND2_X1 U3254 ( .A1(n8255), .A2(n8254), .ZN(n10059) );
  XNOR2_X1 U3192 ( .A(n9912), .B(n9911), .ZN(n11124) );
  INV_X1 U1800 ( .A(n10993), .ZN(n3454) );
  BUF_X1 U1660 ( .A(n11226), .Z(n333) );
  INV_X1 U2018 ( .A(n11086), .ZN(n433) );
  BUF_X1 U2013 ( .A(n10528), .Z(n11261) );
  INV_X2 U1565 ( .A(n11140), .ZN(n3862) );
  BUF_X1 U688 ( .A(n9344), .Z(n10916) );
  OAI22_X1 U8343 ( .A1(n10881), .A2(n10880), .B1(n5063), .B2(n10641), .ZN(
        n12166) );
  MUX2_X1 U16995 ( .A(n10565), .B(n10564), .S(n11196), .Z(n10567) );
  NAND2_X1 U3545 ( .A1(n2351), .A2(n3807), .ZN(n11782) );
  AND2_X1 U9362 ( .A1(n28930), .A2(n28928), .ZN(n11730) );
  INV_X2 U1194 ( .A(n11500), .ZN(n390) );
  NOR2_X1 U1256 ( .A1(n11673), .A2(n11671), .ZN(n11677) );
  INV_X1 U3775 ( .A(n12233), .ZN(n776) );
  NAND3_X1 U3084 ( .A1(n6550), .A2(n6551), .A3(n6549), .ZN(n13461) );
  AND3_X1 U2183 ( .A1(n3200), .A2(n3202), .A3(n2074), .ZN(n12854) );
  NAND3_X1 U8733 ( .A1(n6561), .A2(n10770), .A3(n2538), .ZN(n13547) );
  BUF_X2 U5788 ( .A(n12954), .Z(n12763) );
  NAND4_X1 U1993 ( .A1(n12171), .A2(n12170), .A3(n12168), .A4(n12169), .ZN(
        n13113) );
  NAND2_X1 U1254 ( .A1(n2979), .A2(n12323), .ZN(n13272) );
  XNOR2_X1 U18116 ( .A(n12521), .B(n12919), .ZN(n13434) );
  XNOR2_X1 U5993 ( .A(n12975), .B(n12974), .ZN(n14365) );
  INV_X1 U1546 ( .A(n15194), .ZN(n28172) );
  INV_X1 U1810 ( .A(n13953), .ZN(n28805) );
  AOI22_X1 U1982 ( .A1(n14065), .A2(n14324), .B1(n14328), .B2(n14327), .ZN(
        n13696) );
  INV_X2 U1987 ( .A(n14200), .ZN(n427) );
  AOI21_X1 U5809 ( .B1(n5796), .B2(n308), .A(n14371), .ZN(n14697) );
  AOI22_X1 U19252 ( .A1(n14124), .A2(n14123), .B1(n308), .B2(n14121), .ZN(
        n14153) );
  AOI21_X1 U202 ( .B1(n13768), .B2(n13769), .A(n15193), .ZN(n14961) );
  MUX2_X1 U949 ( .A(n14595), .B(n14594), .S(n14593), .Z(n14762) );
  AND2_X1 U59 ( .A1(n912), .A2(n14096), .ZN(n14518) );
  NAND2_X1 U25597 ( .A1(n14203), .A2(n28684), .ZN(n15338) );
  NAND2_X1 U350 ( .A1(n15346), .A2(n15344), .ZN(n15222) );
  OR2_X1 U14278 ( .A1(n14903), .A2(n14902), .ZN(n15100) );
  BUF_X1 U2825 ( .A(n16691), .Z(n17476) );
  INV_X1 U2788 ( .A(n16944), .ZN(n5398) );
  AND2_X1 U10024 ( .A1(n6013), .A2(n17424), .ZN(n16846) );
  NAND3_X1 U1951 ( .A1(n16277), .A2(n4653), .A3(n4654), .ZN(n1384) );
  NAND2_X1 U11426 ( .A1(n4155), .A2(n4154), .ZN(n17771) );
  NAND2_X1 U2734 ( .A1(n5518), .A2(n5517), .ZN(n17977) );
  OR2_X1 U2757 ( .A1(n17042), .A2(n17041), .ZN(n18334) );
  INV_X1 U3485 ( .A(n15810), .ZN(n18298) );
  NAND3_X1 U1839 ( .A1(n2375), .A2(n6554), .A3(n6553), .ZN(n18020) );
  BUF_X1 U939 ( .A(n17695), .Z(n18279) );
  INV_X1 U386 ( .A(n18017), .ZN(n524) );
  CLKBUF_X1 U569 ( .A(n17207), .Z(n18126) );
  OAI21_X1 U9098 ( .B1(n2791), .B2(n18303), .A(n18302), .ZN(n19631) );
  NAND3_X1 U8367 ( .A1(n2457), .A2(n16189), .A3(n5417), .ZN(n5416) );
  AND2_X1 U1345 ( .A1(n6655), .A2(n6654), .ZN(n18735) );
  NAND2_X1 U5162 ( .A1(n16821), .A2(n28254), .ZN(n18395) );
  OAI211_X1 U21575 ( .C1(n18147), .C2(n18049), .A(n18048), .B(n18047), .ZN(
        n19421) );
  XNOR2_X1 U1737 ( .A(n19051), .B(n19050), .ZN(n20475) );
  NOR2_X1 U22712 ( .A1(n19985), .A2(n29066), .ZN(n20163) );
  INV_X2 U1027 ( .A(n20133), .ZN(n415) );
  NAND2_X1 U10214 ( .A1(n18847), .A2(n835), .ZN(n20875) );
  NAND3_X1 U3960 ( .A1(n2872), .A2(n3411), .A3(n5469), .ZN(n21221) );
  INV_X1 U1132 ( .A(n20864), .ZN(n28789) );
  INV_X1 U7106 ( .A(n21581), .ZN(n5142) );
  OAI211_X1 U22817 ( .C1(n21452), .C2(n21451), .A(n1445), .B(n29178), .ZN(
        n22334) );
  MUX2_X1 U27 ( .A(n20856), .B(n20855), .S(n21143), .Z(n22526) );
  OAI21_X1 U1033 ( .B1(n18851), .B2(n29553), .A(n18850), .ZN(n6520) );
  AND3_X1 U8276 ( .A1(n5634), .A2(n21107), .A3(n21108), .ZN(n22052) );
  NAND2_X1 U9514 ( .A1(n21050), .A2(n3039), .ZN(n22820) );
  NAND3_X1 U12935 ( .A1(n2299), .A2(n19803), .A3(n4225), .ZN(n28450) );
  INV_X1 U24256 ( .A(n23262), .ZN(n23716) );
  CLKBUF_X1 U2427 ( .A(n22954), .Z(n23845) );
  INV_X1 U2404 ( .A(n6227), .ZN(n4231) );
  BUF_X1 U1468 ( .A(n23745), .Z(n24516) );
  MUX2_X1 U20339 ( .A(n23866), .B(n23865), .S(n28531), .Z(n25790) );
  CLKBUF_X1 U13900 ( .A(n25913), .Z(n29039) );
  NAND2_X2 U1060 ( .A1(n6055), .A2(n24587), .ZN(n945) );
  NOR2_X1 U25579 ( .A1(n24286), .A2(n24285), .ZN(n25341) );
  AND4_X1 U1209 ( .A1(n5118), .A2(n5117), .A3(n5115), .A4(n2997), .ZN(n25820)
         );
  INV_X1 U26202 ( .A(n26440), .ZN(n26775) );
  OR2_X1 U5111 ( .A1(n26502), .A2(n3632), .ZN(n27852) );
  AND3_X1 U1612 ( .A1(n6627), .A2(n26759), .A3(n6626), .ZN(n28107) );
  CLKBUF_X1 U2186 ( .A(n27582), .Z(n27586) );
  AOI21_X2 U1001 ( .B1(n11738), .B2(n11737), .A(n11736), .ZN(n13511) );
  AND3_X2 U9975 ( .A1(n2547), .A2(n7929), .A3(n8214), .ZN(n8669) );
  XNOR2_X2 U14673 ( .A(Key[10]), .B(Plaintext[10]), .ZN(n7342) );
  MUX2_X2 U5636 ( .A(n17559), .B(n17558), .S(n29142), .Z(n18251) );
  AND3_X2 U1299 ( .A1(n5081), .A2(n16778), .A3(n16777), .ZN(n18106) );
  OAI21_X2 U10548 ( .B1(n4000), .B2(n11753), .A(n11752), .ZN(n12699) );
  AND2_X2 U1202 ( .A1(n4904), .A2(n4903), .ZN(n11622) );
  OAI211_X2 U9516 ( .C1(n3082), .C2(n6573), .A(n11579), .B(n6572), .ZN(n15415)
         );
  NAND2_X2 U885 ( .A1(n722), .A2(n11464), .ZN(n12817) );
  BUF_X2 U1189 ( .A(n6988), .Z(n7821) );
  OR2_X2 U10359 ( .A1(n5073), .A2(n14397), .ZN(n15265) );
  NAND2_X2 U9835 ( .A1(n18119), .A2(n268), .ZN(n21692) );
  XNOR2_X2 U8364 ( .A(n2387), .B(Key[164]), .ZN(n7997) );
  NAND3_X2 U5117 ( .A1(n6412), .A2(n14782), .A3(n2047), .ZN(n16321) );
  OR2_X2 U313 ( .A1(n17237), .A2(n17238), .ZN(n18433) );
  BUF_X2 U542 ( .A(n7285), .Z(n7796) );
  AND2_X2 U2160 ( .A1(n28720), .A2(n28719), .ZN(n12696) );
  NOR2_X2 U1275 ( .A1(n1929), .A2(n21736), .ZN(n21388) );
  XNOR2_X2 U183 ( .A(n7205), .B(Key[136]), .ZN(n7655) );
  AND2_X2 U1804 ( .A1(n8240), .A2(n8241), .ZN(n8963) );
  AND3_X2 U852 ( .A1(n3525), .A2(n3524), .A3(n3523), .ZN(n19615) );
  NOR2_X2 U483 ( .A1(n9730), .A2(n28269), .ZN(n12198) );
  NAND2_X2 U3921 ( .A1(n7005), .A2(n7006), .ZN(n8699) );
  AND3_X2 U61 ( .A1(n4614), .A2(n4612), .A3(n4613), .ZN(n17942) );
  NOR2_X2 U655 ( .A1(n23130), .A2(n23129), .ZN(n25738) );
  NAND3_X2 U9015 ( .A1(n3979), .A2(n2730), .A3(n3977), .ZN(n16305) );
  NAND2_X2 U565 ( .A1(n13764), .A2(n2408), .ZN(n15202) );
  BUF_X2 U687 ( .A(n14407), .Z(n14332) );
  OR2_X2 U200 ( .A1(n23032), .A2(n23151), .ZN(n24706) );
  INV_X2 U133 ( .A(n6958), .ZN(n7925) );
  NAND2_X2 U15740 ( .A1(n10407), .A2(n10406), .ZN(n10283) );
  AND2_X2 U3126 ( .A1(n2749), .A2(n11783), .ZN(n11550) );
  AND2_X2 U1928 ( .A1(n12368), .A2(n12369), .ZN(n14937) );
  BUF_X2 U23 ( .A(n21775), .Z(n23788) );
  NOR2_X2 U2343 ( .A1(n9239), .A2(n9240), .ZN(n9352) );
  BUF_X2 U2830 ( .A(n16730), .Z(n17497) );
  OAI21_X2 U832 ( .B1(n1237), .B2(n7287), .A(n7286), .ZN(n8891) );
  XNOR2_X2 U526 ( .A(n16220), .B(n16219), .ZN(n17139) );
  NAND2_X2 U31 ( .A1(n4813), .A2(n20073), .ZN(n22013) );
  MUX2_X2 U10898 ( .A(n24385), .B(n24384), .S(n4195), .Z(n26071) );
  BUF_X2 U1402 ( .A(n15018), .Z(n15022) );
  OAI211_X2 U21435 ( .C1(n17810), .C2(n18195), .A(n17809), .B(n17808), .ZN(
        n19679) );
  AND4_X2 U842 ( .A1(n4203), .A2(n4206), .A3(n4202), .A4(n4201), .ZN(n22245)
         );
  AND4_X2 U12983 ( .A1(n15267), .A2(n5721), .A3(n5722), .A4(n5723), .ZN(n16084) );
  XNOR2_X2 U3205 ( .A(n10084), .B(n10083), .ZN(n11152) );
  XNOR2_X2 U24938 ( .A(n18728), .B(n5586), .ZN(n20039) );
  OR2_X2 U2937 ( .A1(n13975), .A2(n13974), .ZN(n15321) );
  XNOR2_X2 U3240 ( .A(n9812), .B(n9510), .ZN(n11038) );
  AND3_X2 U1807 ( .A1(n5919), .A2(n5921), .A3(n2048), .ZN(n18383) );
  NAND2_X2 U1405 ( .A1(n9556), .A2(n9557), .ZN(n12206) );
  OR2_X2 U633 ( .A1(n8949), .A2(n8948), .ZN(n10371) );
  MUX2_X2 U19217 ( .A(n14035), .B(n14034), .S(n14033), .Z(n15284) );
  OAI211_X2 U28241 ( .C1(n14423), .C2(n14422), .A(n14449), .B(n14448), .ZN(
        n15503) );
  XNOR2_X2 U733 ( .A(n7009), .B(Key[66]), .ZN(n8024) );
  OR2_X2 U1200 ( .A1(n3280), .A2(n21936), .ZN(n22811) );
  MUX2_X2 U15590 ( .A(n8447), .B(n8446), .S(n9187), .Z(n10298) );
  BUF_X2 U635 ( .A(n10853), .Z(n1933) );
  OAI21_X2 U13431 ( .B1(n6143), .B2(n14170), .A(n6142), .ZN(n14666) );
  NAND2_X2 U1610 ( .A1(n29237), .A2(n4564), .ZN(n18173) );
  NAND3_X2 U430 ( .A1(n3076), .A2(n3077), .A3(n5668), .ZN(n21090) );
  NAND2_X2 U10767 ( .A1(n24670), .A2(n4603), .ZN(n25869) );
  BUF_X2 U18966 ( .A(n13674), .Z(n14498) );
  NAND2_X2 U8804 ( .A1(n4970), .A2(n10557), .ZN(n12000) );
  AND3_X2 U14887 ( .A1(n7264), .A2(n7263), .A3(n7262), .ZN(n8944) );
  AND2_X2 U3346 ( .A1(n1007), .A2(n7213), .ZN(n9221) );
  OAI21_X2 U114 ( .B1(n984), .B2(n23038), .A(n23037), .ZN(n24707) );
  NAND2_X2 U2888 ( .A1(n6456), .A2(n15317), .ZN(n16625) );
  OAI21_X2 U20139 ( .B1(n24038), .B2(n24039), .A(n24037), .ZN(n28592) );
  INV_X2 U3124 ( .A(n11195), .ZN(n6706) );
  BUF_X2 U262 ( .A(n12607), .Z(n13699) );
  NAND3_X2 U63 ( .A1(n18073), .A2(n4846), .A3(n4845), .ZN(n18508) );
  XNOR2_X2 U16244 ( .A(n9463), .B(n9464), .ZN(n10929) );
  NAND3_X2 U2294 ( .A1(n818), .A2(n23912), .A3(n812), .ZN(n25372) );
  AND3_X2 U1108 ( .A1(n6256), .A2(n18514), .A3(n6255), .ZN(n18652) );
  AND3_X2 U990 ( .A1(n17461), .A2(n17462), .A3(n17460), .ZN(n18213) );
  AND2_X2 U3075 ( .A1(n4276), .A2(n12074), .ZN(n12377) );
  BUF_X2 U1392 ( .A(n23049), .Z(n23193) );
  XNOR2_X2 U1712 ( .A(n20279), .B(n20280), .ZN(n23067) );
  XNOR2_X2 U18588 ( .A(n13100), .B(n6922), .ZN(n14346) );
  XNOR2_X2 U1892 ( .A(n21747), .B(n21746), .ZN(n23787) );
  NAND2_X2 U703 ( .A1(n3733), .A2(n13991), .ZN(n16295) );
  OR2_X2 U14667 ( .A1(n7113), .A2(n7112), .ZN(n8826) );
  NAND2_X2 U392 ( .A1(n21139), .A2(n3534), .ZN(n22822) );
  OAI211_X2 U23141 ( .C1(n29521), .C2(n20514), .A(n20513), .B(n20512), .ZN(
        n21612) );
  NAND2_X2 U869 ( .A1(n2227), .A2(n1163), .ZN(n12332) );
  OR2_X2 U1180 ( .A1(n7190), .A2(n7189), .ZN(n8687) );
  XNOR2_X2 U574 ( .A(n21846), .B(n21845), .ZN(n23776) );
  NAND2_X2 U139 ( .A1(n24418), .A2(n24419), .ZN(n25737) );
  XNOR2_X2 U11087 ( .A(n21169), .B(n21170), .ZN(n23672) );
  XNOR2_X2 U18174 ( .A(n12571), .B(n6923), .ZN(n14314) );
  BUF_X2 U3397 ( .A(n7106), .Z(n7895) );
  BUF_X2 U5534 ( .A(n12712), .Z(n14460) );
  MUX2_X2 U560 ( .A(n16751), .B(n16750), .S(n28454), .Z(n18096) );
  AND2_X2 U3186 ( .A1(n17143), .A2(n17138), .ZN(n17088) );
  AND3_X2 U8731 ( .A1(n2087), .A2(n4087), .A3(n2847), .ZN(n12042) );
  OR2_X2 U1104 ( .A1(n7505), .A2(n7504), .ZN(n8819) );
  AND3_X2 U1073 ( .A1(n5385), .A2(n20507), .A3(n20508), .ZN(n21327) );
  AND2_X2 U370 ( .A1(n1294), .A2(n8789), .ZN(n9934) );
  XNOR2_X2 U28134 ( .A(n15842), .B(n15841), .ZN(n17554) );
  XNOR2_X2 U11101 ( .A(n6051), .B(n13431), .ZN(n3860) );
  MUX2_X2 U8862 ( .A(n9077), .B(n9076), .S(n9075), .Z(n9695) );
  BUF_X2 U4700 ( .A(n16724), .Z(n17477) );
  XNOR2_X2 U11029 ( .A(n9835), .B(n9834), .ZN(n10989) );
  INV_X2 U3272 ( .A(n9785), .ZN(n9677) );
  INV_X2 U2292 ( .A(n24272), .ZN(n26095) );
  XNOR2_X2 U1470 ( .A(n25070), .B(n4810), .ZN(n26919) );
  AND2_X2 U2408 ( .A1(n23651), .A2(n23472), .ZN(n1740) );
  AND3_X2 U3136 ( .A1(n6778), .A2(n6780), .A3(n6777), .ZN(n12304) );
  OAI21_X2 U2744 ( .B1(n17085), .B2(n2609), .A(n17084), .ZN(n18595) );
  XNOR2_X2 U12795 ( .A(n21584), .B(n21583), .ZN(n23666) );
  XNOR2_X2 U2618 ( .A(n19091), .B(n19090), .ZN(n20483) );
  AND2_X2 U1543 ( .A1(n6313), .A2(n6312), .ZN(n22248) );
  MUX2_X2 U178 ( .A(n24154), .B(n24153), .S(n23597), .Z(n25366) );
  OAI21_X2 U23404 ( .B1(n20905), .B2(n20904), .A(n20903), .ZN(n22459) );
  NAND2_X2 U1535 ( .A1(n28727), .A2(n14946), .ZN(n15949) );
  NAND3_X2 U3933 ( .A1(n860), .A2(n4016), .A3(n11957), .ZN(n13488) );
  AND2_X2 U11168 ( .A1(n15349), .A2(n15345), .ZN(n15046) );
  AND3_X2 U1231 ( .A1(n24478), .A2(n24477), .A3(n24476), .ZN(n5146) );
  XNOR2_X2 U980 ( .A(n13492), .B(n13491), .ZN(n5918) );
  OR2_X2 U2878 ( .A1(n3925), .A2(n3923), .ZN(n1967) );
  AND3_X2 U2024 ( .A1(n8822), .A2(n1813), .A3(n8821), .ZN(n9505) );
  NAND2_X2 U7787 ( .A1(n28883), .A2(n16938), .ZN(n18529) );
  XNOR2_X2 U16435 ( .A(n9690), .B(n9691), .ZN(n11053) );
  NAND4_X2 U4855 ( .A1(n8640), .A2(n8641), .A3(n8842), .A4(n1311), .ZN(n9746)
         );
  OAI211_X2 U1163 ( .C1(n6640), .C2(n6639), .A(n13466), .B(n3613), .ZN(n14972)
         );
  XNOR2_X2 U5890 ( .A(n9299), .B(n9300), .ZN(n10976) );
  XNOR2_X2 U3216 ( .A(n16317), .B(n16316), .ZN(n17062) );
  NOR2_X2 U677 ( .A1(n8374), .A2(n8373), .ZN(n10330) );
  INV_X2 U23881 ( .A(n22618), .ZN(n22724) );
  AND3_X2 U1708 ( .A1(n28259), .A2(n20246), .A3(n28258), .ZN(n22618) );
  INV_X2 U6509 ( .A(n21649), .ZN(n22610) );
  OAI211_X2 U3154 ( .C1(n6021), .C2(n11130), .A(n11129), .B(n11128), .ZN(
        n11778) );
  AND2_X2 U2943 ( .A1(n1321), .A2(n14548), .ZN(n15171) );
  BUF_X2 U28304 ( .A(n13824), .Z(n13826) );
  AND2_X2 U2718 ( .A1(n17096), .A2(n17095), .ZN(n18144) );
  XNOR2_X2 U4429 ( .A(n19366), .B(n19365), .ZN(n20619) );
  BUF_X2 U1292 ( .A(n16289), .Z(n321) );
  OR2_X2 U2005 ( .A1(n10812), .A2(n10813), .ZN(n11715) );
  AOI21_X2 U297 ( .B1(n18036), .B2(n17745), .A(n17622), .ZN(n18738) );
  NAND2_X2 U12120 ( .A1(n26803), .A2(n3075), .ZN(n27277) );
  NOR2_X2 U9761 ( .A1(n20337), .A2(n3144), .ZN(n21177) );
  AND2_X2 U148 ( .A1(n15194), .A2(n14241), .ZN(n14172) );
  XNOR2_X2 U815 ( .A(n11481), .B(n11480), .ZN(n14241) );
  XNOR2_X2 U2373 ( .A(Key[119]), .B(Plaintext[119]), .ZN(n29135) );
  XNOR2_X2 U577 ( .A(n16490), .B(n16489), .ZN(n17484) );
  OAI21_X2 U985 ( .B1(n7908), .B2(n8651), .A(n7907), .ZN(n4479) );
  OR2_X2 U384 ( .A1(n839), .A2(n8344), .ZN(n10138) );
  AND3_X2 U272 ( .A1(n28292), .A2(n18227), .A3(n28672), .ZN(n5439) );
  BUF_X2 U3402 ( .A(n7072), .Z(n7580) );
  AND3_X2 U13726 ( .A1(n15277), .A2(n15278), .A3(n6493), .ZN(n15545) );
  AOI21_X2 U442 ( .B1(n19817), .B2(n19816), .A(n1970), .ZN(n21493) );
  MUX2_X2 U9471 ( .A(n23328), .B(n23327), .S(n23474), .Z(n24677) );
  NAND3_X2 U1934 ( .A1(n5843), .A2(n5842), .A3(n16664), .ZN(n1741) );
  NAND2_X2 U2293 ( .A1(n3206), .A2(n2473), .ZN(n26118) );
  NOR2_X2 U27119 ( .A1(n26417), .A2(n26416), .ZN(n27255) );
  OAI21_X2 U208 ( .B1(n23479), .B2(n23478), .A(n23477), .ZN(n24779) );
  XNOR2_X2 U3477 ( .A(Key[2]), .B(Plaintext[2]), .ZN(n7089) );
  XNOR2_X2 U11002 ( .A(n15610), .B(n15609), .ZN(n17385) );
  XNOR2_X2 U14687 ( .A(n7123), .B(Key[40]), .ZN(n8143) );
  OAI21_X2 U19888 ( .B1(n15416), .B2(n223), .A(n15414), .ZN(n16649) );
  OAI211_X2 U1655 ( .C1(n11062), .C2(n11061), .A(n11060), .B(n11059), .ZN(
        n12827) );
  XNOR2_X2 U3245 ( .A(n9497), .B(n9496), .ZN(n11315) );
  NAND2_X2 U1239 ( .A1(n1298), .A2(n1297), .ZN(n8760) );
  NOR2_X1 U3654 ( .A1(n3760), .A2(n3759), .ZN(n3758) );
  XNOR2_X2 U553 ( .A(n19068), .B(n19067), .ZN(n20481) );
  AND2_X2 U8225 ( .A1(n6093), .A2(n6094), .ZN(n9028) );
  INV_X1 U22984 ( .A(n20207), .ZN(n21678) );
  AND2_X2 U255 ( .A1(n17789), .A2(n17788), .ZN(n18181) );
  XNOR2_X2 U447 ( .A(n18631), .B(n18632), .ZN(n20401) );
  AND2_X2 U2667 ( .A1(n2775), .A2(n2774), .ZN(n19370) );
  NOR2_X2 U322 ( .A1(n10168), .A2(n10167), .ZN(n1890) );
  INV_X2 U640 ( .A(n18782), .ZN(n19592) );
  OR2_X2 U641 ( .A1(n18427), .A2(n18428), .ZN(n18782) );
  NAND4_X2 U657 ( .A1(n1791), .A2(n5957), .A3(n8333), .A4(n1790), .ZN(n10171)
         );
  OAI211_X2 U184 ( .C1(n11558), .C2(n3946), .A(n3944), .B(n11557), .ZN(n13364)
         );
  MUX2_X2 U10840 ( .A(n17311), .B(n17310), .S(n17440), .Z(n18156) );
  AND2_X2 U2740 ( .A1(n5107), .A2(n2030), .ZN(n17989) );
  AND2_X2 U1656 ( .A1(n2106), .A2(n2105), .ZN(n26004) );
  OAI211_X2 U5736 ( .C1(n14967), .C2(n14968), .A(n14966), .B(n28856), .ZN(
        n16534) );
  NAND2_X2 U1061 ( .A1(n195), .A2(n3578), .ZN(n22791) );
  INV_X2 U1210 ( .A(n11247), .ZN(n12049) );
  OR2_X2 U2365 ( .A1(n5626), .A2(n5627), .ZN(n24643) );
  NAND2_X2 U287 ( .A1(n12126), .A2(n13203), .ZN(n13406) );
  BUF_X2 U1383 ( .A(n19678), .Z(n19464) );
  NOR2_X2 U1970 ( .A1(n14733), .A2(n14115), .ZN(n14512) );
  BUF_X2 U5930 ( .A(n6958), .Z(n7625) );
  OR3_X2 U27246 ( .A1(n26596), .A2(n27875), .A3(n27865), .ZN(n26597) );
  BUF_X2 U2403 ( .A(n23245), .Z(n23577) );
  OR2_X2 U3379 ( .A1(n7833), .A2(n7834), .ZN(n8910) );
  BUF_X1 U3050 ( .A(n12388), .Z(n12684) );
  MUX2_X2 U2298 ( .A(n24399), .B(n24398), .S(n24676), .Z(n25900) );
  AOI21_X2 U16703 ( .B1(n10054), .B2(n10053), .A(n10052), .ZN(n11853) );
  OAI211_X2 U3266 ( .C1(n8761), .C2(n8569), .A(n7387), .B(n7386), .ZN(n10364)
         );
  NAND2_X2 U13669 ( .A1(n10533), .A2(n6430), .ZN(n6432) );
  NAND2_X2 U19744 ( .A1(n15064), .A2(n15063), .ZN(n16619) );
  XNOR2_X2 U14444 ( .A(n6978), .B(Key[97]), .ZN(n7634) );
  BUF_X2 U296 ( .A(n27081), .Z(n27085) );
  NAND3_X2 U4545 ( .A1(n1805), .A2(n23044), .A3(n23043), .ZN(n1808) );
  OAI21_X2 U13124 ( .B1(n20912), .B2(n21607), .A(n20911), .ZN(n22123) );
  OR2_X1 U3384 ( .A1(n8315), .A2(n8314), .ZN(n8802) );
  AND4_X1 U367 ( .A1(n7270), .A2(n7272), .A3(n7269), .A4(n7271), .ZN(n8762) );
  BUF_X1 U1590 ( .A(Key[167]), .Z(n27225) );
  BUF_X1 U501 ( .A(n9913), .Z(n11121) );
  BUF_X1 U580 ( .A(n13837), .Z(n14150) );
  NAND3_X1 U2929 ( .A1(n5641), .A2(n2969), .A3(n5642), .ZN(n14916) );
  OAI21_X1 U1972 ( .B1(n13736), .B2(n557), .A(n13735), .ZN(n15371) );
  BUF_X2 U1497 ( .A(n15085), .Z(n323) );
  AND2_X1 U8561 ( .A1(n14501), .A2(n6797), .ZN(n15494) );
  INV_X1 U6023 ( .A(n15108), .ZN(n15406) );
  BUF_X1 U2940 ( .A(n14621), .Z(n15502) );
  OAI21_X1 U12513 ( .B1(n13950), .B2(n14667), .A(n13949), .ZN(n16564) );
  MUX2_X1 U1965 ( .A(n14525), .B(n14524), .S(n550), .Z(n16405) );
  BUF_X1 U20056 ( .A(n15617), .Z(n16636) );
  AND2_X1 U1193 ( .A1(n3917), .A2(n3919), .ZN(n16556) );
  OAI21_X1 U46 ( .B1(n16705), .B2(n28574), .A(n16704), .ZN(n18449) );
  AND2_X1 U2721 ( .A1(n16441), .A2(n16440), .ZN(n18467) );
  AOI21_X2 U12232 ( .B1(n17503), .B2(n17504), .A(n4963), .ZN(n18393) );
  BUF_X2 U1503 ( .A(n17534), .Z(n17842) );
  AND2_X1 U3841 ( .A1(n16663), .A2(n824), .ZN(n18311) );
  BUF_X1 U755 ( .A(n19556), .Z(n28144) );
  AND2_X1 U189 ( .A1(n28898), .A2(n4793), .ZN(n21656) );
  BUF_X1 U1181 ( .A(n22765), .Z(n28162) );
  INV_X1 U7245 ( .A(n22356), .ZN(n24744) );
  BUF_X1 U4 ( .A(n25182), .Z(n25441) );
  NAND3_X1 U5 ( .A1(n29352), .A2(n153), .A3(n24126), .ZN(n26110) );
  NOR2_X1 U13 ( .A1(n1330), .A2(n1329), .ZN(n20814) );
  INV_X1 U15 ( .A(n17881), .ZN(n17883) );
  AND3_X1 U17 ( .A1(n5894), .A2(n5893), .A3(n13925), .ZN(n16090) );
  XNOR2_X1 U19 ( .A(n12703), .B(n12702), .ZN(n14459) );
  BUF_X1 U20 ( .A(n5595), .Z(n29316) );
  BUF_X2 U36 ( .A(n18613), .Z(n20383) );
  OR2_X2 U37 ( .A1(n26744), .A2(n26743), .ZN(n29056) );
  NOR2_X2 U38 ( .A1(n23346), .A2(n23345), .ZN(n24074) );
  OR2_X2 U71 ( .A1(n6181), .A2(n11869), .ZN(n11457) );
  AND3_X2 U80 ( .A1(n6260), .A2(n28215), .A3(n6259), .ZN(n21675) );
  NOR2_X1 U101 ( .A1(n20860), .A2(n20861), .ZN(n22670) );
  BUF_X2 U104 ( .A(n25267), .Z(n26757) );
  MUX2_X2 U107 ( .A(n12533), .B(n12532), .S(n13872), .Z(n14907) );
  NAND2_X2 U110 ( .A1(n15273), .A2(n15954), .ZN(n16387) );
  NAND2_X2 U116 ( .A1(n8467), .A2(n29439), .ZN(n9964) );
  AOI211_X2 U117 ( .C1(n11232), .C2(n9709), .A(n10621), .B(n28568), .ZN(n10626) );
  NAND2_X2 U125 ( .A1(n10608), .A2(n29710), .ZN(n12362) );
  NAND2_X2 U131 ( .A1(n3563), .A2(n3562), .ZN(n22891) );
  OAI22_X2 U134 ( .A1(n20697), .A2(n20983), .B1(n20698), .B2(n20699), .ZN(
        n22796) );
  XNOR2_X2 U138 ( .A(n13544), .B(n29798), .ZN(n13572) );
  BUF_X2 U141 ( .A(n16993), .Z(n29299) );
  NOR2_X2 U144 ( .A1(n19750), .A2(n20383), .ZN(n20571) );
  AOI21_X2 U152 ( .B1(n24004), .B2(n24547), .A(n24003), .ZN(n26109) );
  NAND4_X2 U156 ( .A1(n13680), .A2(n13681), .A3(n14187), .A4(n13679), .ZN(
        n15144) );
  OAI21_X2 U162 ( .B1(n3529), .B2(n29718), .A(n6335), .ZN(n17818) );
  OR2_X2 U163 ( .A1(n29794), .A2(n7526), .ZN(n8593) );
  OAI21_X2 U169 ( .B1(n15191), .B2(n15190), .A(n15189), .ZN(n16407) );
  XNOR2_X2 U170 ( .A(n15876), .B(n15875), .ZN(n17568) );
  AND2_X2 U180 ( .A1(n26431), .A2(n26382), .ZN(n26380) );
  BUF_X2 U230 ( .A(n12053), .Z(n285) );
  OAI211_X2 U251 ( .C1(n14804), .C2(n14803), .A(n14805), .B(n785), .ZN(n4504)
         );
  XNOR2_X2 U259 ( .A(n25023), .B(n25022), .ZN(n27181) );
  AND2_X2 U260 ( .A1(n20617), .A2(n20618), .ZN(n19890) );
  BUF_X2 U261 ( .A(n26728), .Z(n29501) );
  AND2_X2 U263 ( .A1(n4597), .A2(n4594), .ZN(n24758) );
  XNOR2_X2 U264 ( .A(n7073), .B(Key[179]), .ZN(n7887) );
  BUF_X2 U274 ( .A(n25998), .Z(n27368) );
  AOI21_X2 U281 ( .B1(n12090), .B2(n12089), .A(n430), .ZN(n12995) );
  INV_X2 U286 ( .A(n2155), .ZN(n18465) );
  AND3_X2 U288 ( .A1(n28983), .A2(n4768), .A3(n4770), .ZN(n24745) );
  INV_X2 U289 ( .A(n19843), .ZN(n29315) );
  AND2_X2 U290 ( .A1(n1832), .A2(n20864), .ZN(n21183) );
  AOI21_X2 U294 ( .B1(n21469), .B2(n28155), .A(n29435), .ZN(n22677) );
  NOR2_X2 U298 ( .A1(n12995), .A2(n12101), .ZN(n13331) );
  OAI211_X2 U304 ( .C1(n8882), .C2(n8881), .A(n8880), .B(n8879), .ZN(n1852) );
  AND2_X1 U309 ( .A1(n26434), .A2(n26433), .ZN(n29493) );
  AND3_X1 U321 ( .A1(n26453), .A2(n6736), .A3(n2043), .ZN(n29542) );
  INV_X1 U360 ( .A(n25633), .ZN(n27386) );
  AND2_X1 U379 ( .A1(n21655), .A2(n21656), .ZN(n29334) );
  OR2_X1 U385 ( .A1(n14702), .A2(n14916), .ZN(n15268) );
  AND2_X1 U390 ( .A1(n18471), .A2(n18467), .ZN(n18315) );
  BUF_X1 U401 ( .A(n26575), .Z(n29576) );
  OR2_X1 U412 ( .A1(n6578), .A2(n20219), .ZN(n2096) );
  BUF_X1 U413 ( .A(n24214), .Z(n29307) );
  BUF_X1 U431 ( .A(n24214), .Z(n29309) );
  OAI211_X1 U432 ( .C1(n8430), .C2(n7809), .A(n7808), .B(n7807), .ZN(n9550) );
  CLKBUF_X1 U436 ( .A(n11646), .Z(n11712) );
  CLKBUF_X1 U454 ( .A(n15167), .Z(n15474) );
  XOR2_X1 U456 ( .A(n16372), .B(n16371), .Z(n29294) );
  NOR2_X2 U472 ( .A1(n17870), .A2(n17869), .ZN(n18760) );
  OAI211_X2 U485 ( .C1(n19764), .C2(n29491), .A(n19763), .B(n1699), .ZN(n21118) );
  AOI22_X1 U487 ( .A1(n21480), .A2(n29314), .B1(n21478), .B2(n21479), .ZN(
        n21649) );
  NOR2_X2 U489 ( .A1(n22930), .A2(n22929), .ZN(n24593) );
  AOI21_X2 U494 ( .B1(n22454), .B2(n22453), .A(n29169), .ZN(n24614) );
  XNOR2_X2 U496 ( .A(n25073), .B(n26104), .ZN(n26782) );
  OAI21_X2 U498 ( .B1(n19063), .B2(n19062), .A(n19061), .ZN(n21703) );
  XNOR2_X2 U499 ( .A(n7202), .B(Key[133]), .ZN(n7657) );
  OAI21_X2 U502 ( .B1(n23105), .B2(n23301), .A(n23104), .ZN(n24209) );
  AOI21_X2 U523 ( .B1(n11292), .B2(n10663), .A(n10327), .ZN(n12177) );
  XNOR2_X2 U529 ( .A(n13326), .B(n13327), .ZN(n13730) );
  BUF_X1 U546 ( .A(n23450), .Z(n29295) );
  BUF_X1 U554 ( .A(n23450), .Z(n29296) );
  XNOR2_X1 U558 ( .A(n22695), .B(n22696), .ZN(n23450) );
  NOR2_X2 U570 ( .A1(n7044), .A2(n4825), .ZN(n8808) );
  AND3_X2 U579 ( .A1(n19911), .A2(n5938), .A3(n29265), .ZN(n22330) );
  AOI22_X2 U581 ( .A1(n7224), .A2(n7465), .B1(n7223), .B2(n7222), .ZN(n9220)
         );
  CLKBUF_X1 U596 ( .A(n16993), .Z(n29297) );
  CLKBUF_X1 U600 ( .A(n16993), .Z(n29298) );
  XNOR2_X1 U615 ( .A(n14592), .B(n14591), .ZN(n16993) );
  MUX2_X2 U629 ( .A(n14880), .B(n14879), .S(n15691), .Z(n15982) );
  XNOR2_X2 U630 ( .A(n19908), .B(n19909), .ZN(n23529) );
  NAND3_X2 U631 ( .A1(n5975), .A2(n19943), .A3(n5976), .ZN(n22265) );
  XNOR2_X2 U638 ( .A(n7029), .B(Key[61]), .ZN(n8032) );
  XNOR2_X2 U644 ( .A(n12845), .B(n12844), .ZN(n14193) );
  OR2_X2 U646 ( .A1(n7435), .A2(n7434), .ZN(n9070) );
  CLKBUF_X1 U647 ( .A(n359), .Z(n29300) );
  BUF_X1 U664 ( .A(n359), .Z(n29301) );
  BUF_X1 U666 ( .A(n359), .Z(n29302) );
  XNOR2_X1 U673 ( .A(Plaintext[158]), .B(Key[158]), .ZN(n359) );
  XNOR2_X2 U692 ( .A(n29451), .B(Key[169]), .ZN(n441) );
  XNOR2_X2 U693 ( .A(n10182), .B(n10181), .ZN(n11242) );
  INV_X1 U707 ( .A(n11192), .ZN(n11355) );
  CLKBUF_X1 U711 ( .A(n9123), .Z(n29303) );
  BUF_X2 U712 ( .A(n9123), .Z(n29304) );
  XNOR2_X2 U714 ( .A(n22505), .B(n22504), .ZN(n22531) );
  NAND3_X2 U716 ( .A1(n7848), .A2(n7847), .A3(n29771), .ZN(n9014) );
  CLKBUF_X1 U724 ( .A(n13946), .Z(n29305) );
  BUF_X2 U727 ( .A(n13946), .Z(n29306) );
  XNOR2_X1 U728 ( .A(n12048), .B(n12047), .ZN(n13946) );
  XNOR2_X2 U729 ( .A(n12825), .B(n6343), .ZN(n14194) );
  NOR2_X2 U742 ( .A1(n14839), .A2(n14840), .ZN(n15887) );
  BUF_X1 U748 ( .A(n24214), .Z(n29308) );
  AOI22_X1 U762 ( .A1(n23473), .A2(n23654), .B1(n28391), .B2(n23471), .ZN(
        n24214) );
  CLKBUF_X1 U764 ( .A(n28606), .Z(n29310) );
  BUF_X1 U770 ( .A(n28606), .Z(n29311) );
  XNOR2_X2 U774 ( .A(n6208), .B(Key[168]), .ZN(n7591) );
  BUF_X2 U788 ( .A(n22494), .Z(n23839) );
  OAI21_X2 U791 ( .B1(n8601), .B2(n9062), .A(n8600), .ZN(n9601) );
  NAND2_X2 U792 ( .A1(n5243), .A2(n5239), .ZN(n8828) );
  NAND2_X2 U795 ( .A1(n2895), .A2(n12372), .ZN(n16310) );
  OAI21_X2 U797 ( .B1(n11490), .B2(n11489), .A(n11488), .ZN(n13263) );
  NOR2_X2 U805 ( .A1(n5320), .A2(n23255), .ZN(n24368) );
  XNOR2_X2 U813 ( .A(n7026), .B(Key[62]), .ZN(n7265) );
  OAI211_X2 U816 ( .C1(n17664), .C2(n17665), .A(n5700), .B(n5701), .ZN(n19465)
         );
  XNOR2_X2 U818 ( .A(n12175), .B(n12174), .ZN(n14260) );
  XNOR2_X2 U823 ( .A(n10049), .B(n6107), .ZN(n10919) );
  AOI21_X2 U824 ( .B1(n13996), .B2(n13995), .A(n13994), .ZN(n16062) );
  BUF_X2 U825 ( .A(n28588), .Z(n29312) );
  XNOR2_X2 U826 ( .A(n7052), .B(Key[171]), .ZN(n7231) );
  XNOR2_X2 U828 ( .A(Key[118]), .B(Plaintext[118]), .ZN(n7933) );
  XNOR2_X2 U830 ( .A(n13344), .B(n13345), .ZN(n13912) );
  OAI21_X2 U835 ( .B1(n4022), .B2(n8274), .A(n8273), .ZN(n8958) );
  XNOR2_X2 U840 ( .A(Key[70]), .B(Plaintext[70]), .ZN(n7844) );
  XNOR2_X2 U841 ( .A(n6989), .B(Key[91]), .ZN(n7822) );
  NAND2_X2 U844 ( .A1(n938), .A2(n1171), .ZN(n10183) );
  NAND4_X2 U862 ( .A1(n14537), .A2(n14538), .A3(n14536), .A4(n14535), .ZN(
        n15927) );
  XNOR2_X2 U872 ( .A(n7061), .B(Key[163]), .ZN(n7995) );
  AOI21_X2 U874 ( .B1(n7344), .B2(n4051), .A(n7343), .ZN(n8563) );
  OAI22_X2 U879 ( .A1(n6811), .A2(n6429), .B1(n18254), .B2(n28370), .ZN(n28516) );
  XNOR2_X2 U880 ( .A(n21952), .B(n21953), .ZN(n23247) );
  OAI21_X2 U886 ( .B1(n6346), .B2(n20803), .A(n6345), .ZN(n22903) );
  BUF_X2 U888 ( .A(n21359), .Z(n28586) );
  XNOR2_X2 U917 ( .A(Key[142]), .B(Plaintext[142]), .ZN(n8280) );
  XNOR2_X2 U919 ( .A(n12656), .B(n12655), .ZN(n14452) );
  XNOR2_X2 U928 ( .A(n12552), .B(n12553), .ZN(n14317) );
  XNOR2_X2 U935 ( .A(Key[117]), .B(Plaintext[117]), .ZN(n7614) );
  OAI211_X2 U944 ( .C1(n6716), .C2(n6019), .A(n6243), .B(n2935), .ZN(n19632)
         );
  NAND2_X2 U945 ( .A1(n4192), .A2(n4905), .ZN(n6314) );
  OAI22_X2 U952 ( .A1(n8538), .A2(n28845), .B1(n8542), .B2(n8731), .ZN(n9626)
         );
  XNOR2_X2 U957 ( .A(n18257), .B(n18258), .ZN(n20547) );
  XNOR2_X2 U962 ( .A(n16474), .B(n16475), .ZN(n17505) );
  XNOR2_X2 U966 ( .A(n8125), .B(n8126), .ZN(n11330) );
  OAI21_X2 U967 ( .B1(n9192), .B2(n9191), .A(n9190), .ZN(n10072) );
  XNOR2_X2 U971 ( .A(n16413), .B(n16412), .ZN(n17181) );
  XNOR2_X2 U974 ( .A(n16098), .B(n15521), .ZN(n17414) );
  XNOR2_X2 U975 ( .A(Key[183]), .B(Plaintext[183]), .ZN(n7172) );
  OAI21_X2 U976 ( .B1(n21181), .B2(n21180), .A(n879), .ZN(n22514) );
  XNOR2_X2 U981 ( .A(n7046), .B(Key[156]), .ZN(n7675) );
  NOR2_X2 U982 ( .A1(n26462), .A2(n6221), .ZN(n27426) );
  MUX2_X2 U984 ( .A(n10095), .B(n10094), .S(n10905), .Z(n13219) );
  OAI211_X2 U996 ( .C1(n5040), .C2(n12134), .A(n5039), .B(n5038), .ZN(n13459)
         );
  NOR2_X2 U997 ( .A1(n29351), .A2(n21830), .ZN(n24726) );
  XNOR2_X2 U1017 ( .A(Key[127]), .B(Plaintext[127]), .ZN(n7618) );
  OAI211_X2 U1019 ( .C1(n8609), .C2(n7419), .A(n6405), .B(n6404), .ZN(n4713)
         );
  OAI211_X2 U1025 ( .C1(n8463), .C2(n7120), .A(n7119), .B(n2410), .ZN(n9799)
         );
  OAI211_X2 U1034 ( .C1(n4895), .C2(n4896), .A(n6873), .B(n4894), .ZN(n15456)
         );
  AND3_X2 U1037 ( .A1(n1676), .A2(n2451), .A3(n1675), .ZN(n24373) );
  AOI21_X2 U1044 ( .B1(n21529), .B2(n21528), .A(n1263), .ZN(n24751) );
  XNOR2_X2 U1046 ( .A(n19259), .B(n4307), .ZN(n4569) );
  XNOR2_X2 U1047 ( .A(n7008), .B(Key[71]), .ZN(n29106) );
  XNOR2_X2 U1054 ( .A(n9459), .B(n9458), .ZN(n10932) );
  XNOR2_X2 U1069 ( .A(n12446), .B(n12445), .ZN(n14402) );
  OAI22_X2 U1070 ( .A1(n3201), .A2(n11854), .B1(n3307), .B2(n3306), .ZN(n12978) );
  XNOR2_X2 U1081 ( .A(n14954), .B(n14955), .ZN(n17437) );
  XNOR2_X2 U1088 ( .A(Plaintext[32]), .B(Key[32]), .ZN(n7349) );
  NOR2_X2 U1109 ( .A1(n4343), .A2(n21324), .ZN(n22386) );
  OR2_X1 U1111 ( .A1(n442), .A2(n27625), .ZN(n29463) );
  INV_X1 U1115 ( .A(n4823), .ZN(n27458) );
  OAI211_X1 U1116 ( .C1(n2140), .C2(n1950), .A(n2139), .B(n2038), .ZN(n27628)
         );
  INV_X1 U1130 ( .A(n24433), .ZN(n29726) );
  INV_X1 U1150 ( .A(n23525), .ZN(n23663) );
  INV_X1 U1156 ( .A(n21291), .ZN(n29313) );
  INV_X1 U1159 ( .A(n21387), .ZN(n29314) );
  NAND2_X1 U1165 ( .A1(n29425), .A2(n18446), .ZN(n19219) );
  NAND2_X1 U1212 ( .A1(n3597), .A2(n17764), .ZN(n2759) );
  INV_X2 U1213 ( .A(n14894), .ZN(n3362) );
  AND3_X1 U1225 ( .A1(n13723), .A2(n13722), .A3(n2144), .ZN(n15372) );
  INV_X2 U1248 ( .A(n14317), .ZN(n14313) );
  NAND3_X1 U1255 ( .A1(n29466), .A2(n11966), .A3(n2976), .ZN(n13209) );
  NAND2_X1 U1271 ( .A1(n12154), .A2(n29705), .ZN(n13433) );
  INV_X2 U1276 ( .A(n12428), .ZN(n29735) );
  BUF_X1 U1284 ( .A(n12577), .Z(n28202) );
  OR2_X1 U1286 ( .A1(n7035), .A2(n7034), .ZN(n10297) );
  BUF_X1 U1290 ( .A(n7114), .Z(n8824) );
  OAI21_X1 U1291 ( .B1(n7999), .B2(n7881), .A(n5363), .ZN(n8500) );
  AND2_X1 U1298 ( .A1(n7844), .A2(n29321), .ZN(n29772) );
  BUF_X1 U1306 ( .A(Key[39]), .Z(n3083) );
  CLKBUF_X1 U1309 ( .A(Key[62]), .Z(n2350) );
  BUF_X1 U1310 ( .A(Key[53]), .Z(n27422) );
  BUF_X1 U1312 ( .A(Key[165]), .Z(n3565) );
  BUF_X1 U1313 ( .A(Key[45]), .Z(n3643) );
  BUF_X2 U1314 ( .A(n8300), .Z(n29317) );
  OR2_X1 U1320 ( .A1(n307), .A2(n26817), .ZN(n29389) );
  NAND2_X1 U1328 ( .A1(n26137), .A2(n26136), .ZN(n27711) );
  BUF_X2 U1330 ( .A(n28091), .Z(n28794) );
  NAND4_X1 U1331 ( .A1(n6302), .A2(n6300), .A3(n26327), .A4(n6301), .ZN(n27807) );
  AND3_X1 U1336 ( .A1(n768), .A2(n28100), .A3(n767), .ZN(n28111) );
  AND3_X1 U1337 ( .A1(n29454), .A2(n28822), .A3(n28969), .ZN(n27571) );
  OAI21_X1 U1346 ( .B1(n4739), .B2(n28410), .A(n28398), .ZN(n27650) );
  INV_X1 U1354 ( .A(n27551), .ZN(n29445) );
  AND2_X1 U1366 ( .A1(n29778), .A2(n5300), .ZN(n27859) );
  OAI21_X1 U1375 ( .B1(n6823), .B2(n26574), .A(n6825), .ZN(n6824) );
  BUF_X1 U1378 ( .A(n27120), .Z(n29016) );
  BUF_X1 U1397 ( .A(n27044), .Z(n28130) );
  XNOR2_X1 U1399 ( .A(n25539), .B(n25538), .ZN(n28783) );
  INV_X1 U1411 ( .A(n26079), .ZN(n29410) );
  AND2_X1 U1419 ( .A1(n5101), .A2(n5104), .ZN(n25921) );
  OR2_X1 U1420 ( .A1(n24128), .A2(n5752), .ZN(n29352) );
  INV_X1 U1431 ( .A(n28223), .ZN(n29677) );
  AND2_X1 U1432 ( .A1(n5647), .A2(n5646), .ZN(n24544) );
  AND3_X1 U1438 ( .A1(n6764), .A2(n6763), .A3(n1965), .ZN(n29471) );
  AND3_X1 U1452 ( .A1(n23653), .A2(n5555), .A3(n23652), .ZN(n24794) );
  AND3_X1 U1483 ( .A1(n23359), .A2(n23358), .A3(n6628), .ZN(n24666) );
  AOI22_X1 U1490 ( .A1(n23316), .A2(n28390), .B1(n23317), .B2(n23565), .ZN(
        n28635) );
  BUF_X1 U1499 ( .A(n22566), .Z(n29564) );
  OR2_X1 U1505 ( .A1(n22458), .A2(n28183), .ZN(n29729) );
  XNOR2_X1 U1510 ( .A(n22254), .B(n22253), .ZN(n23640) );
  BUF_X1 U1516 ( .A(n23773), .Z(n29641) );
  INV_X1 U1518 ( .A(n28582), .ZN(n29402) );
  XNOR2_X1 U1525 ( .A(n6520), .B(n22670), .ZN(n22828) );
  AOI22_X1 U1526 ( .A1(n21115), .A2(n1897), .B1(n21114), .B2(n21463), .ZN(
        n29519) );
  INV_X1 U1536 ( .A(n20857), .ZN(n21157) );
  INV_X1 U1547 ( .A(n20756), .ZN(n21463) );
  INV_X1 U1554 ( .A(n20786), .ZN(n29586) );
  NAND3_X1 U1556 ( .A1(n3972), .A2(n21134), .A3(n3971), .ZN(n20886) );
  NAND2_X1 U1562 ( .A1(n19866), .A2(n29348), .ZN(n21155) );
  OAI211_X1 U1571 ( .C1(n19972), .C2(n19973), .A(n29347), .B(n29346), .ZN(
        n21387) );
  AND2_X1 U1577 ( .A1(n20334), .A2(n20626), .ZN(n20006) );
  BUF_X2 U1581 ( .A(n19766), .Z(n21091) );
  BUF_X1 U1583 ( .A(n21353), .Z(n28491) );
  XNOR2_X1 U1592 ( .A(n5005), .B(n5006), .ZN(n20441) );
  AND3_X1 U1633 ( .A1(n29386), .A2(n6483), .A3(n29385), .ZN(n18778) );
  INV_X1 U1643 ( .A(n3444), .ZN(n29318) );
  OAI21_X1 U1668 ( .B1(n18297), .B2(n18296), .A(n18295), .ZN(n19482) );
  NAND2_X1 U1693 ( .A1(n2501), .A2(n2498), .ZN(n19332) );
  OR2_X1 U1704 ( .A1(n17014), .A2(n18600), .ZN(n4419) );
  OR2_X1 U1707 ( .A1(n1436), .A2(n17765), .ZN(n3597) );
  OR2_X1 U1714 ( .A1(n17976), .A2(n521), .ZN(n29715) );
  AND2_X1 U1722 ( .A1(n29191), .A2(n29192), .ZN(n16868) );
  OR2_X1 U1726 ( .A1(n17746), .A2(n29663), .ZN(n17809) );
  BUF_X2 U1728 ( .A(n18601), .Z(n28142) );
  OAI21_X1 U1741 ( .B1(n5287), .B2(n5288), .A(n29674), .ZN(n18304) );
  OR2_X1 U1749 ( .A1(n18507), .A2(n18508), .ZN(n29350) );
  NAND2_X1 U1756 ( .A1(n17499), .A2(n18226), .ZN(n18388) );
  INV_X1 U1757 ( .A(n18195), .ZN(n29663) );
  INV_X1 U1763 ( .A(n18530), .ZN(n29336) );
  OAI21_X1 U1778 ( .B1(n16748), .B2(n17350), .A(n17349), .ZN(n18090) );
  NOR2_X1 U1782 ( .A1(n16806), .A2(n16668), .ZN(n16850) );
  BUF_X1 U1783 ( .A(n17250), .Z(n29503) );
  XNOR2_X1 U1791 ( .A(n15832), .B(n15831), .ZN(n17553) );
  XNOR2_X1 U1806 ( .A(n14603), .B(n14602), .ZN(n14629) );
  XNOR2_X1 U1840 ( .A(n15995), .B(n15996), .ZN(n17248) );
  XNOR2_X1 U1847 ( .A(n16480), .B(n1967), .ZN(n15973) );
  AND3_X1 U1849 ( .A1(n29326), .A2(n1000), .A3(n1006), .ZN(n15971) );
  INV_X1 U1866 ( .A(n16322), .ZN(n29319) );
  NOR2_X1 U1871 ( .A1(n15022), .A2(n15303), .ZN(n14657) );
  OR2_X1 U1883 ( .A1(n15223), .A2(n15224), .ZN(n29355) );
  AND2_X1 U1888 ( .A1(n1111), .A2(n13584), .ZN(n14944) );
  AND3_X1 U1903 ( .A1(n3357), .A2(n3356), .A3(n29325), .ZN(n15132) );
  OR2_X1 U1906 ( .A1(n1660), .A2(n13900), .ZN(n29682) );
  AND2_X1 U1908 ( .A1(n14415), .A2(n14215), .ZN(n29760) );
  OR2_X1 U1935 ( .A1(n4893), .A2(n13826), .ZN(n14125) );
  OR2_X1 U1962 ( .A1(n14484), .A2(n29305), .ZN(n14167) );
  INV_X1 U1967 ( .A(n14480), .ZN(n29320) );
  NAND2_X1 U1976 ( .A1(n12029), .A2(n1192), .ZN(n12913) );
  OAI21_X1 U1996 ( .B1(n11588), .B2(n11589), .A(n29354), .ZN(n13061) );
  AND2_X1 U2029 ( .A1(n4997), .A2(n4996), .ZN(n12632) );
  OAI211_X1 U2045 ( .C1(n11521), .C2(n11836), .A(n11520), .B(n29670), .ZN(
        n13270) );
  AND2_X1 U2053 ( .A1(n11990), .A2(n12508), .ZN(n29671) );
  OR2_X1 U2091 ( .A1(n29462), .A2(n29460), .ZN(n12315) );
  NAND3_X1 U2096 ( .A1(n10583), .A2(n10581), .A3(n10582), .ZN(n12022) );
  AND2_X1 U2099 ( .A1(n5704), .A2(n5705), .ZN(n12150) );
  INV_X1 U2102 ( .A(n11896), .ZN(n29461) );
  NAND2_X1 U2138 ( .A1(n8577), .A2(n4440), .ZN(n9763) );
  NAND3_X1 U2152 ( .A1(n29393), .A2(n749), .A3(n8613), .ZN(n748) );
  NAND2_X1 U2157 ( .A1(n8854), .A2(n8853), .ZN(n9619) );
  AND3_X1 U2211 ( .A1(n9537), .A2(n29660), .A3(n29661), .ZN(n10033) );
  BUF_X2 U2212 ( .A(n10222), .Z(n301) );
  NAND2_X1 U2214 ( .A1(n6172), .A2(n29650), .ZN(n9794) );
  INV_X1 U2230 ( .A(n8500), .ZN(n29416) );
  AND3_X1 U2242 ( .A1(n8017), .A2(n6807), .A3(n8020), .ZN(n9122) );
  NAND2_X1 U2243 ( .A1(n7469), .A2(n29756), .ZN(n8726) );
  INV_X1 U2246 ( .A(n24166), .ZN(n5490) );
  XNOR2_X1 U2248 ( .A(n7153), .B(Key[31]), .ZN(n8165) );
  XNOR2_X1 U2257 ( .A(n7218), .B(Key[130]), .ZN(n6782) );
  OR2_X1 U2268 ( .A1(n7162), .A2(n7320), .ZN(n7769) );
  XNOR2_X1 U2275 ( .A(Key[59]), .B(Plaintext[59]), .ZN(n29629) );
  INV_X1 U2277 ( .A(n7850), .ZN(n29321) );
  AND2_X1 U2290 ( .A1(n7468), .A2(n7467), .ZN(n29756) );
  XNOR2_X1 U2291 ( .A(Key[50]), .B(Plaintext[50]), .ZN(n7141) );
  OR2_X1 U2299 ( .A1(n9196), .A2(n9206), .ZN(n28861) );
  INV_X1 U2346 ( .A(n8891), .ZN(n8887) );
  AOI22_X1 U2402 ( .A1(n6689), .A2(n8591), .B1(n8975), .B2(n607), .ZN(n6688)
         );
  OR2_X1 U2420 ( .A1(n9126), .A2(n284), .ZN(n29650) );
  OR2_X1 U2428 ( .A1(n8956), .A2(n8955), .ZN(n8625) );
  OAI21_X1 U2438 ( .B1(n604), .B2(n8770), .A(n8579), .ZN(n9582) );
  CLKBUF_X1 U2444 ( .A(n8586), .Z(n29147) );
  OAI21_X1 U2469 ( .B1(n9137), .B2(n8552), .A(n8551), .ZN(n9851) );
  OR2_X1 U2512 ( .A1(n11045), .A2(n11267), .ZN(n2754) );
  XNOR2_X1 U2513 ( .A(n10022), .B(n9550), .ZN(n10179) );
  XNOR2_X1 U2515 ( .A(n10043), .B(n27422), .ZN(n9750) );
  BUF_X1 U2522 ( .A(n9863), .Z(n10957) );
  XNOR2_X1 U2523 ( .A(n9960), .B(n9959), .ZN(n10497) );
  XNOR2_X1 U2536 ( .A(n9600), .B(n9599), .ZN(n29148) );
  AND3_X1 U2547 ( .A1(n3801), .A2(n3800), .A3(n3805), .ZN(n12097) );
  XNOR2_X1 U2554 ( .A(n9813), .B(n9812), .ZN(n10991) );
  BUF_X1 U2567 ( .A(n10747), .Z(n10563) );
  OR2_X1 U2571 ( .A1(n10696), .A2(n10980), .ZN(n2422) );
  OR2_X1 U2658 ( .A1(n11782), .A2(n11419), .ZN(n1493) );
  INV_X1 U2675 ( .A(n12111), .ZN(n6281) );
  BUF_X1 U2679 ( .A(n11730), .Z(n13206) );
  NAND3_X1 U2690 ( .A1(n29208), .A2(n3103), .A3(n11899), .ZN(n12352) );
  AND2_X1 U2703 ( .A1(n11947), .A2(n11945), .ZN(n11861) );
  OAI21_X1 U2732 ( .B1(n11008), .B2(n11009), .A(n3013), .ZN(n12070) );
  NOR2_X1 U2750 ( .A1(n11869), .A2(n11867), .ZN(n11501) );
  AND2_X1 U2775 ( .A1(n12207), .A2(n12211), .ZN(n12115) );
  AND2_X1 U2778 ( .A1(n11587), .A2(n11586), .ZN(n29354) );
  CLKBUF_X1 U2824 ( .A(n11058), .Z(n11435) );
  INV_X1 U2845 ( .A(n11878), .ZN(n567) );
  NAND2_X1 U2848 ( .A1(n2272), .A2(n2271), .ZN(n10453) );
  OAI21_X1 U2853 ( .B1(n12516), .B2(n11567), .A(n11566), .ZN(n3871) );
  NAND2_X1 U2856 ( .A1(n12293), .A2(n12290), .ZN(n12289) );
  XNOR2_X1 U2898 ( .A(n13413), .B(n11912), .ZN(n13274) );
  OAI21_X1 U2908 ( .B1(n14213), .B2(n14402), .A(n14212), .ZN(n15239) );
  XNOR2_X1 U2911 ( .A(n12897), .B(n12898), .ZN(n14082) );
  BUF_X1 U2965 ( .A(n14479), .Z(n293) );
  MUX2_X1 U2974 ( .A(n14154), .B(n14155), .S(n29037), .Z(n15346) );
  OAI211_X1 U3010 ( .C1(n14480), .C2(n293), .A(n14478), .B(n14477), .ZN(n15485) );
  OR2_X1 U3048 ( .A1(n15250), .A2(n15135), .ZN(n14729) );
  OR2_X1 U3062 ( .A1(n14639), .A2(n14874), .ZN(n15081) );
  BUF_X1 U3069 ( .A(n15001), .Z(n14998) );
  NAND2_X1 U3072 ( .A1(n3012), .A2(n3010), .ZN(n15224) );
  AOI21_X1 U3080 ( .B1(n15091), .B2(n15690), .A(n15694), .ZN(n15089) );
  OR2_X1 U3083 ( .A1(n15041), .A2(n15040), .ZN(n28306) );
  OR2_X1 U3140 ( .A1(n15245), .A2(n15244), .ZN(n29675) );
  OAI211_X1 U3143 ( .C1(n15168), .C2(n15473), .A(n14801), .B(n15472), .ZN(
        n3856) );
  AND4_X2 U3184 ( .A1(n6332), .A2(n6333), .A3(n15016), .A4(n15017), .ZN(n16283) );
  XNOR2_X1 U3226 ( .A(n16509), .B(n16585), .ZN(n16119) );
  XNOR2_X1 U3230 ( .A(n15865), .B(n15092), .ZN(n16598) );
  OR2_X1 U3248 ( .A1(n17293), .A2(n17401), .ZN(n5487) );
  OR2_X1 U3289 ( .A1(n17120), .A2(n16811), .ZN(n17116) );
  XNOR2_X1 U3304 ( .A(n16336), .B(n16335), .ZN(n17491) );
  INV_X1 U3389 ( .A(n17498), .ZN(n538) );
  XNOR2_X1 U3440 ( .A(n16021), .B(n16020), .ZN(n17018) );
  INV_X1 U3451 ( .A(n17275), .ZN(n29421) );
  XOR2_X1 U3466 ( .A(n15604), .B(n15603), .Z(n28497) );
  OR2_X1 U3486 ( .A1(n29373), .A2(n17491), .ZN(n17493) );
  INV_X1 U3488 ( .A(n17720), .ZN(n17431) );
  XNOR2_X1 U3512 ( .A(n15748), .B(n15749), .ZN(n29550) );
  BUF_X1 U3552 ( .A(n17433), .Z(n29566) );
  OR2_X1 U3569 ( .A1(n6927), .A2(n2656), .ZN(n2216) );
  OR2_X1 U3571 ( .A1(n16986), .A2(n18087), .ZN(n18186) );
  INV_X1 U3581 ( .A(n16611), .ZN(n518) );
  OR2_X1 U3589 ( .A1(n17842), .A2(n18241), .ZN(n17757) );
  OR2_X1 U3590 ( .A1(n18448), .A2(n18447), .ZN(n29425) );
  OR2_X1 U3601 ( .A1(n18143), .A2(n18144), .ZN(n2635) );
  OR2_X1 U3673 ( .A1(n5589), .A2(n6484), .ZN(n29385) );
  AOI22_X1 U3681 ( .A1(n18381), .A2(n18382), .B1(n5670), .B2(n17883), .ZN(
        n3207) );
  BUF_X1 U3685 ( .A(n17793), .Z(n18445) );
  NAND2_X1 U3687 ( .A1(n3874), .A2(n3876), .ZN(n19278) );
  BUF_X1 U3699 ( .A(n20017), .Z(n28489) );
  INV_X1 U3734 ( .A(n20568), .ZN(n97) );
  OR2_X1 U3744 ( .A1(n97), .A2(n19833), .ZN(n20570) );
  OAI21_X1 U3754 ( .B1(n19867), .B2(n499), .A(n20491), .ZN(n29349) );
  INV_X1 U3780 ( .A(n20227), .ZN(n29426) );
  BUF_X1 U3796 ( .A(n20484), .Z(n29527) );
  AND2_X1 U3802 ( .A1(n29315), .A2(n18838), .ZN(n19779) );
  BUF_X1 U3844 ( .A(n21355), .Z(n28126) );
  INV_X1 U3848 ( .A(n506), .ZN(n29707) );
  AND2_X1 U3878 ( .A1(n20488), .A2(n19093), .ZN(n20359) );
  AND2_X1 U3888 ( .A1(n28236), .A2(n28235), .ZN(n29659) );
  NAND2_X1 U3895 ( .A1(n3551), .A2(n20301), .ZN(n29531) );
  NOR2_X1 U3896 ( .A1(n21410), .A2(n20663), .ZN(n21230) );
  OAI211_X1 U3925 ( .C1(n20460), .C2(n28408), .A(n4568), .B(n29184), .ZN(
        n21509) );
  OR2_X1 U3939 ( .A1(n20728), .A2(n21292), .ZN(n3252) );
  OR2_X1 U3959 ( .A1(n21481), .A2(n21483), .ZN(n21579) );
  OR2_X1 U3968 ( .A1(n20979), .A2(n20978), .ZN(n29591) );
  NAND3_X1 U3981 ( .A1(n5139), .A2(n5141), .A3(n5140), .ZN(n21987) );
  XNOR2_X1 U4007 ( .A(n29763), .B(n22884), .ZN(n5862) );
  INV_X1 U4016 ( .A(n21798), .ZN(n29417) );
  XNOR2_X1 U4020 ( .A(n22121), .B(n22120), .ZN(n28484) );
  OR2_X1 U4033 ( .A1(n5883), .A2(n23517), .ZN(n29358) );
  BUF_X1 U4037 ( .A(n23156), .Z(n23779) );
  CLKBUF_X1 U4056 ( .A(n23525), .Z(n29123) );
  INV_X1 U4163 ( .A(n23386), .ZN(n22084) );
  XNOR2_X1 U4173 ( .A(n21799), .B(n29417), .ZN(n28554) );
  BUF_X1 U4213 ( .A(n23629), .Z(n23636) );
  CLKBUF_X1 U4214 ( .A(n22174), .Z(n23260) );
  BUF_X1 U4233 ( .A(n24409), .Z(n28524) );
  OR2_X1 U4238 ( .A1(n23803), .A2(n23541), .ZN(n6763) );
  OAI22_X1 U4255 ( .A1(n4686), .A2(n23660), .B1(n405), .B2(n23659), .ZN(n24813) );
  NAND2_X1 U4257 ( .A1(n29259), .A2(n6195), .ZN(n24629) );
  AOI21_X1 U4259 ( .B1(n23846), .B2(n22455), .A(n23843), .ZN(n22129) );
  INV_X1 U4260 ( .A(n22931), .ZN(n23819) );
  OR2_X1 U4272 ( .A1(n29128), .A2(n24347), .ZN(n29727) );
  BUF_X1 U4289 ( .A(n24813), .Z(n24810) );
  OAI211_X1 U4300 ( .C1(n23500), .C2(n5355), .A(n5353), .B(n5354), .ZN(n23945)
         );
  CLKBUF_X1 U4314 ( .A(Key[126]), .Z(n4029) );
  MUX2_X1 U4359 ( .A(n3671), .B(n23752), .S(n24420), .Z(n23753) );
  OR2_X1 U4363 ( .A1(n29028), .A2(n26466), .ZN(n25617) );
  XNOR2_X1 U4378 ( .A(n26043), .B(n26042), .ZN(n26050) );
  XNOR2_X1 U4390 ( .A(n26071), .B(n1459), .ZN(n25541) );
  OR2_X1 U4404 ( .A1(n29479), .A2(n26240), .ZN(n29388) );
  NOR2_X1 U4418 ( .A1(n1874), .A2(n26740), .ZN(n29459) );
  XNOR2_X1 U4457 ( .A(n23919), .B(n23920), .ZN(n26449) );
  OR2_X1 U4461 ( .A1(n26791), .A2(n23862), .ZN(n28709) );
  XOR2_X1 U4467 ( .A(n24989), .B(n24988), .Z(n28535) );
  CLKBUF_X1 U4504 ( .A(n1907), .Z(n29487) );
  INV_X1 U4543 ( .A(n27663), .ZN(n29449) );
  XNOR2_X1 U4555 ( .A(n26078), .B(n29410), .ZN(n29633) );
  OR2_X1 U4556 ( .A1(n29480), .A2(n29121), .ZN(n29681) );
  AND2_X1 U4566 ( .A1(n6492), .A2(n6026), .ZN(n29070) );
  OR3_X1 U4568 ( .A1(n27442), .A2(n27433), .A3(n26682), .ZN(n25423) );
  MUX2_X1 U4581 ( .A(n27180), .B(n27179), .S(n27178), .Z(n27661) );
  OAI211_X1 U4598 ( .C1(n5299), .C2(n26511), .A(n5297), .B(n29615), .ZN(n29778) );
  NAND2_X1 U4610 ( .A1(n26337), .A2(n5485), .ZN(n27817) );
  CLKBUF_X1 U4628 ( .A(Key[133]), .Z(n2389) );
  INV_X1 U4669 ( .A(n1193), .ZN(n26713) );
  CLKBUF_X1 U4677 ( .A(Key[84]), .Z(n1225) );
  CLKBUF_X1 U4683 ( .A(Key[31]), .Z(n3414) );
  CLKBUF_X1 U4684 ( .A(Key[7]), .Z(n1079) );
  CLKBUF_X1 U4690 ( .A(Key[36]), .Z(n3256) );
  CLKBUF_X1 U4691 ( .A(Key[124]), .Z(n2960) );
  AND3_X1 U4725 ( .A1(n17898), .A2(n18356), .A3(n18355), .ZN(n29322) );
  AND2_X1 U4732 ( .A1(n673), .A2(n28481), .ZN(n29323) );
  INV_X1 U4744 ( .A(n9530), .ZN(n29662) );
  INV_X1 U4753 ( .A(n8749), .ZN(n29395) );
  NAND2_X1 U4757 ( .A1(n28674), .A2(n28913), .ZN(n8693) );
  AND2_X1 U4761 ( .A1(n4095), .A2(n5717), .ZN(n29324) );
  OR2_X1 U4772 ( .A1(n14080), .A2(n561), .ZN(n29325) );
  INV_X1 U4776 ( .A(n14278), .ZN(n29691) );
  NAND2_X1 U4788 ( .A1(n15120), .A2(n1904), .ZN(n29326) );
  INV_X1 U4798 ( .A(n15144), .ZN(n29380) );
  INV_X1 U4830 ( .A(n17470), .ZN(n29406) );
  XNOR2_X1 U4861 ( .A(n16181), .B(n16180), .ZN(n17280) );
  INV_X1 U4869 ( .A(n17280), .ZN(n29737) );
  CLKBUF_X1 U4874 ( .A(n19054), .Z(n20177) );
  AND2_X1 U4878 ( .A1(n18529), .A2(n29335), .ZN(n29327) );
  AND2_X1 U4882 ( .A1(n3551), .A2(n20301), .ZN(n29328) );
  OR3_X1 U4886 ( .A1(n21709), .A2(n21372), .A3(n21277), .ZN(n29329) );
  INV_X1 U4895 ( .A(n21211), .ZN(n29364) );
  NOR2_X1 U4896 ( .A1(n1330), .A2(n1329), .ZN(n29488) );
  INV_X1 U4898 ( .A(n24373), .ZN(n29340) );
  INV_X1 U4987 ( .A(n24258), .ZN(n24976) );
  OAI211_X1 U4991 ( .C1(n23466), .C2(n23465), .A(n23464), .B(n23463), .ZN(
        n24258) );
  INV_X1 U5031 ( .A(n27364), .ZN(n29387) );
  XOR2_X1 U5042 ( .A(n25093), .B(n25092), .Z(n29330) );
  BUF_X1 U5055 ( .A(n27028), .Z(n306) );
  OR3_X1 U5061 ( .A1(n27417), .A2(n26531), .A3(n26530), .ZN(n29331) );
  NAND2_X1 U5070 ( .A1(n26195), .A2(n27393), .ZN(n29332) );
  NAND2_X1 U5073 ( .A1(n3967), .A2(n19798), .ZN(n20756) );
  NOR2_X2 U5114 ( .A1(n11581), .A2(n6848), .ZN(n12881) );
  NAND3_X2 U5148 ( .A1(n20836), .A2(n20835), .A3(n29333), .ZN(n6458) );
  NAND2_X1 U5175 ( .A1(n6275), .A2(n29334), .ZN(n29333) );
  NAND3_X1 U5177 ( .A1(n29336), .A2(n4280), .A3(n4281), .ZN(n29335) );
  NAND2_X1 U5193 ( .A1(n29337), .A2(n23399), .ZN(n751) );
  NAND2_X1 U5211 ( .A1(n754), .A2(n755), .ZN(n29337) );
  OR2_X1 U5234 ( .A1(n17030), .A2(n17357), .ZN(n4279) );
  OAI21_X1 U5239 ( .B1(n27025), .B2(n24364), .A(n29338), .ZN(n27033) );
  NAND2_X1 U5247 ( .A1(n27029), .A2(n27025), .ZN(n29338) );
  OAI21_X2 U5252 ( .B1(n2726), .B2(n14114), .A(n14113), .ZN(n16329) );
  OAI21_X1 U5304 ( .B1(n23995), .B2(n29340), .A(n29339), .ZN(n23905) );
  NAND2_X1 U5305 ( .A1(n23995), .A2(n24380), .ZN(n29339) );
  NAND2_X1 U5319 ( .A1(n29341), .A2(n23235), .ZN(n23236) );
  NAND2_X1 U5324 ( .A1(n23584), .A2(n23260), .ZN(n29341) );
  NAND3_X1 U5326 ( .A1(n1836), .A2(n11874), .A3(n11360), .ZN(n2355) );
  OR2_X1 U5335 ( .A1(n24577), .A2(n6741), .ZN(n1204) );
  OAI21_X1 U5369 ( .B1(n18429), .B2(n420), .A(n29342), .ZN(n29797) );
  NAND3_X1 U5403 ( .A1(n2853), .A2(n2855), .A3(n18431), .ZN(n29342) );
  NAND4_X2 U5489 ( .A1(n6547), .A2(n2816), .A3(n6548), .A4(n24424), .ZN(n25864) );
  OAI22_X1 U5490 ( .A1(n15146), .A2(n3208), .B1(n1326), .B2(n15145), .ZN(
        n15149) );
  NAND2_X1 U5495 ( .A1(n17557), .A2(n17553), .ZN(n17224) );
  NAND2_X2 U5530 ( .A1(n29343), .A2(n26144), .ZN(n27725) );
  NOR2_X1 U5532 ( .A1(n26141), .A2(n26142), .ZN(n29343) );
  NAND2_X1 U5542 ( .A1(n14833), .A2(n893), .ZN(n15291) );
  NAND2_X1 U5543 ( .A1(n14095), .A2(n6000), .ZN(n14833) );
  NAND2_X1 U5548 ( .A1(n17123), .A2(n29344), .ZN(n17125) );
  NAND3_X1 U5561 ( .A1(n17477), .A2(n1816), .A3(n3883), .ZN(n29344) );
  NAND2_X1 U5606 ( .A1(n7159), .A2(n29345), .ZN(n10346) );
  OR2_X1 U5714 ( .A1(n7160), .A2(n7161), .ZN(n29345) );
  MUX2_X1 U5716 ( .A(n24726), .B(n24596), .S(n24725), .Z(n21944) );
  NAND2_X1 U5729 ( .A1(n29733), .A2(n21864), .ZN(n24725) );
  NAND2_X1 U5798 ( .A1(n19973), .A2(n20295), .ZN(n29346) );
  NAND2_X1 U5826 ( .A1(n19970), .A2(n20290), .ZN(n29347) );
  NAND2_X1 U5883 ( .A1(n20857), .A2(n21155), .ZN(n3762) );
  INV_X1 U5901 ( .A(n29349), .ZN(n29348) );
  NAND2_X1 U5995 ( .A1(n27188), .A2(n26401), .ZN(n26360) );
  NAND3_X1 U6011 ( .A1(n3360), .A2(n15108), .A3(n3361), .ZN(n3919) );
  NAND2_X1 U6018 ( .A1(n16868), .A2(n16867), .ZN(n18761) );
  OAI211_X1 U6030 ( .C1(n18512), .C2(n418), .A(n29350), .B(n18516), .ZN(n6256)
         );
  NAND2_X1 U6038 ( .A1(n28353), .A2(n6461), .ZN(n29351) );
  NAND3_X2 U6053 ( .A1(n16786), .A2(n1226), .A3(n16785), .ZN(n18107) );
  XNOR2_X1 U6058 ( .A(n25891), .B(n5146), .ZN(n24487) );
  NOR2_X2 U6063 ( .A1(n6420), .A2(n6422), .ZN(n25891) );
  XNOR2_X2 U6091 ( .A(n29353), .B(n22850), .ZN(n28182) );
  INV_X1 U6125 ( .A(n22849), .ZN(n29353) );
  NAND3_X1 U6133 ( .A1(n24578), .A2(n24468), .A3(n24582), .ZN(n6421) );
  NAND2_X1 U6181 ( .A1(n1631), .A2(n24617), .ZN(n24024) );
  AND2_X2 U6204 ( .A1(n29658), .A2(n29659), .ZN(n21192) );
  OR2_X2 U6225 ( .A1(n28337), .A2(n1210), .ZN(n6095) );
  NAND3_X1 U6228 ( .A1(n5669), .A2(n273), .A3(n4235), .ZN(n5817) );
  INV_X1 U6261 ( .A(n25659), .ZN(n25660) );
  XNOR2_X1 U6263 ( .A(n25296), .B(n25297), .ZN(n25659) );
  NAND2_X1 U6290 ( .A1(n15226), .A2(n29355), .ZN(n15231) );
  XNOR2_X1 U6313 ( .A(n19687), .B(n19688), .ZN(n29769) );
  NAND4_X2 U6352 ( .A1(n5235), .A2(n5232), .A3(n5231), .A4(n17768), .ZN(n19687) );
  NAND2_X1 U6387 ( .A1(n18511), .A2(n18512), .ZN(n18513) );
  NAND2_X1 U6395 ( .A1(n24236), .A2(n24568), .ZN(n23176) );
  NAND2_X1 U6403 ( .A1(n24643), .A2(n24638), .ZN(n24236) );
  NAND2_X1 U6469 ( .A1(n29356), .A2(n6600), .ZN(n6597) );
  OAI21_X1 U6477 ( .B1(n24162), .B2(n28522), .A(n24802), .ZN(n29356) );
  OAI21_X1 U6501 ( .B1(n23211), .B2(n22985), .A(n29357), .ZN(n2621) );
  NAND3_X1 U6516 ( .A1(n23604), .A2(n23583), .A3(n23578), .ZN(n29357) );
  NAND2_X1 U6550 ( .A1(n21159), .A2(n20744), .ZN(n20746) );
  NAND2_X1 U6568 ( .A1(n5881), .A2(n29358), .ZN(n5885) );
  NAND3_X1 U6596 ( .A1(n29359), .A2(n19802), .A3(n20631), .ZN(n21464) );
  NAND2_X1 U6613 ( .A1(n6059), .A2(n20012), .ZN(n29359) );
  NAND2_X1 U6615 ( .A1(n14426), .A2(n4522), .ZN(n13704) );
  NOR2_X2 U6643 ( .A1(n23907), .A2(n3028), .ZN(n26055) );
  NAND3_X2 U6644 ( .A1(n29361), .A2(n3059), .A3(n29360), .ZN(n25577) );
  NAND2_X1 U6666 ( .A1(n29323), .A2(n24653), .ZN(n29360) );
  OR2_X1 U6676 ( .A1(n24006), .A2(n24653), .ZN(n29361) );
  AND2_X2 U6704 ( .A1(n3231), .A2(n3230), .ZN(n28456) );
  NAND2_X1 U6722 ( .A1(n14413), .A2(n14414), .ZN(n14446) );
  NAND2_X1 U6780 ( .A1(n12481), .A2(n14444), .ZN(n14413) );
  NAND2_X1 U6946 ( .A1(n14754), .A2(n29362), .ZN(n16495) );
  OAI21_X1 U6954 ( .B1(n14750), .B2(n14751), .A(n15243), .ZN(n29362) );
  NAND3_X1 U7025 ( .A1(n5927), .A2(n20141), .A3(n21088), .ZN(n1245) );
  OAI211_X2 U7058 ( .C1(n23542), .C2(n23541), .A(n2326), .B(n712), .ZN(n24768)
         );
  NAND2_X1 U7073 ( .A1(n29477), .A2(n2070), .ZN(n5618) );
  OR2_X1 U7095 ( .A1(n5023), .A2(n18708), .ZN(n863) );
  NAND2_X1 U7100 ( .A1(n15095), .A2(n15096), .ZN(n2497) );
  NOR2_X1 U7184 ( .A1(n17992), .A2(n17994), .ZN(n17881) );
  OAI22_X1 U7195 ( .A1(n241), .A2(n17339), .B1(n5226), .B2(n17342), .ZN(n17992) );
  NAND3_X2 U7201 ( .A1(n3648), .A2(n4409), .A3(n4410), .ZN(n22286) );
  INV_X1 U7224 ( .A(n22294), .ZN(n22027) );
  NAND2_X1 U7280 ( .A1(n29364), .A2(n29363), .ZN(n22294) );
  INV_X1 U7346 ( .A(n21208), .ZN(n29363) );
  NAND3_X1 U7398 ( .A1(n15293), .A2(n3827), .A3(n15291), .ZN(n14520) );
  NAND2_X1 U7405 ( .A1(n29366), .A2(n29365), .ZN(n26349) );
  NAND2_X1 U7423 ( .A1(n26347), .A2(n27585), .ZN(n29365) );
  NAND2_X1 U7424 ( .A1(n26348), .A2(n27591), .ZN(n29366) );
  AND2_X2 U7472 ( .A1(n3713), .A2(n29367), .ZN(n25826) );
  INV_X1 U7491 ( .A(n29368), .ZN(n29367) );
  OAI21_X1 U7492 ( .B1(n3715), .B2(n464), .A(n3714), .ZN(n29368) );
  OAI21_X1 U7518 ( .B1(n23628), .B2(n23632), .A(n23040), .ZN(n22277) );
  NAND3_X1 U7528 ( .A1(n122), .A2(n18087), .A3(n123), .ZN(n28892) );
  NOR2_X1 U7593 ( .A1(n20616), .A2(n19920), .ZN(n20430) );
  XNOR2_X2 U7604 ( .A(n19358), .B(n19357), .ZN(n20616) );
  NAND2_X1 U7631 ( .A1(n19825), .A2(n19826), .ZN(n1832) );
  NAND2_X1 U7679 ( .A1(n26567), .A2(n26912), .ZN(n4455) );
  AND3_X2 U7686 ( .A1(n3130), .A2(n3129), .A3(n2431), .ZN(n11640) );
  NAND2_X1 U7745 ( .A1(n18197), .A2(n18193), .ZN(n18194) );
  NAND2_X1 U7772 ( .A1(n29369), .A2(n6494), .ZN(n20749) );
  NAND2_X1 U7789 ( .A1(n4472), .A2(n19848), .ZN(n29369) );
  NAND3_X1 U7809 ( .A1(n16729), .A2(n2578), .A3(n2579), .ZN(n4705) );
  OAI22_X2 U7815 ( .A1(n21165), .A2(n21166), .B1(n21326), .B2(n159), .ZN(
        n22506) );
  MUX2_X1 U7828 ( .A(n29139), .B(n11671), .S(n11640), .Z(n11402) );
  NAND2_X1 U7878 ( .A1(n5868), .A2(n8523), .ZN(n5867) );
  OAI21_X1 U7896 ( .B1(n24579), .B2(n24578), .A(n24469), .ZN(n6422) );
  XNOR2_X1 U7963 ( .A(n29370), .B(n2389), .ZN(Ciphertext[8]) );
  NAND2_X1 U7982 ( .A1(n1681), .A2(n29278), .ZN(n29370) );
  NAND2_X1 U7983 ( .A1(n11239), .A2(n29371), .ZN(n28944) );
  NAND3_X1 U8005 ( .A1(n11235), .A2(n11237), .A3(n11236), .ZN(n29371) );
  AND2_X2 U8021 ( .A1(n29372), .A2(n7311), .ZN(n9425) );
  NAND3_X1 U8029 ( .A1(n7307), .A2(n4438), .A3(n4439), .ZN(n29372) );
  INV_X1 U8034 ( .A(n16612), .ZN(n29373) );
  OAI211_X2 U8047 ( .C1(n4539), .C2(n10693), .A(n4537), .B(n10692), .ZN(n12303) );
  NAND2_X1 U8048 ( .A1(n8163), .A2(n8164), .ZN(n8172) );
  NAND3_X1 U8064 ( .A1(n747), .A2(n746), .A3(n7895), .ZN(n997) );
  NAND3_X1 U8066 ( .A1(n28839), .A2(n29374), .A3(n28838), .ZN(n11739) );
  AOI22_X1 U8085 ( .A1(n10612), .A2(n10972), .B1(n10969), .B2(n5267), .ZN(
        n29374) );
  NAND2_X1 U8104 ( .A1(n29375), .A2(n196), .ZN(n27634) );
  NAND2_X1 U8141 ( .A1(n2414), .A2(n2415), .ZN(n29375) );
  NAND2_X1 U8144 ( .A1(n16739), .A2(n16738), .ZN(n18204) );
  NAND2_X1 U8151 ( .A1(n8167), .A2(n7298), .ZN(n8169) );
  NAND2_X1 U8177 ( .A1(n29376), .A2(n21463), .ZN(n2299) );
  NAND2_X1 U8180 ( .A1(n4224), .A2(n4223), .ZN(n29376) );
  NAND2_X1 U8196 ( .A1(n29377), .A2(n18260), .ZN(n2705) );
  OAI21_X1 U8204 ( .B1(n17699), .B2(n18535), .A(n18259), .ZN(n29377) );
  OAI21_X1 U8264 ( .B1(n16824), .B2(n17291), .A(n28729), .ZN(n28728) );
  NOR2_X1 U8284 ( .A1(n17395), .A2(n17397), .ZN(n17291) );
  AND2_X2 U8290 ( .A1(n1373), .A2(n1656), .ZN(n18241) );
  NAND2_X1 U8291 ( .A1(n29433), .A2(n6464), .ZN(n29432) );
  OR2_X2 U8293 ( .A1(n17608), .A2(n3847), .ZN(n18799) );
  NAND3_X1 U8295 ( .A1(n6020), .A2(n11702), .A3(n4844), .ZN(n11705) );
  NAND3_X1 U8314 ( .A1(n11952), .A2(n11944), .A3(n11943), .ZN(n2440) );
  NAND2_X1 U8323 ( .A1(n4455), .A2(n29378), .ZN(n1021) );
  NAND2_X1 U8371 ( .A1(n26786), .A2(n26565), .ZN(n29378) );
  INV_X1 U8375 ( .A(n14633), .ZN(n14722) );
  NAND2_X1 U8383 ( .A1(n29379), .A2(n15389), .ZN(n14634) );
  NAND2_X1 U8446 ( .A1(n14633), .A2(n29380), .ZN(n29379) );
  NAND2_X1 U8459 ( .A1(n14992), .A2(n15387), .ZN(n14633) );
  NAND2_X1 U8479 ( .A1(n28871), .A2(n28817), .ZN(n29787) );
  NOR2_X2 U8482 ( .A1(n29382), .A2(n29381), .ZN(n25386) );
  OAI22_X1 U8487 ( .A1(n24311), .A2(n24390), .B1(n24312), .B2(n2649), .ZN(
        n29381) );
  AND2_X1 U8513 ( .A1(n24314), .A2(n24682), .ZN(n29382) );
  NAND2_X1 U8528 ( .A1(n28901), .A2(n18083), .ZN(n28900) );
  OR2_X1 U8541 ( .A1(n19938), .A2(n19810), .ZN(n29706) );
  OAI211_X1 U8544 ( .C1(n4232), .C2(n23140), .A(n23012), .B(n29383), .ZN(
        n23014) );
  NAND3_X1 U8550 ( .A1(n23011), .A2(n4232), .A3(n23351), .ZN(n29383) );
  NOR2_X2 U8575 ( .A1(n3732), .A2(n5972), .ZN(n13262) );
  OR2_X1 U8597 ( .A1(n17155), .A2(n17336), .ZN(n6336) );
  OAI21_X1 U8603 ( .B1(n27443), .B2(n26833), .A(n26832), .ZN(n26834) );
  NAND3_X1 U8605 ( .A1(n20982), .A2(n21008), .A3(n21809), .ZN(n2259) );
  NAND2_X1 U8606 ( .A1(n3637), .A2(n29384), .ZN(n7693) );
  NAND3_X1 U8619 ( .A1(n7691), .A2(n7818), .A3(n7690), .ZN(n29384) );
  NOR2_X1 U8631 ( .A1(n17900), .A2(n29322), .ZN(n29386) );
  NAND3_X1 U8632 ( .A1(n29541), .A2(n28562), .A3(n29387), .ZN(n5359) );
  NAND4_X2 U8637 ( .A1(n6882), .A2(n6881), .A3(n20260), .A4(n6883), .ZN(n5151)
         );
  XNOR2_X1 U8640 ( .A(n16255), .B(n16126), .ZN(n16499) );
  NAND3_X2 U8642 ( .A1(n15325), .A2(n3626), .A3(n3627), .ZN(n16255) );
  NAND2_X1 U8647 ( .A1(n25649), .A2(n29388), .ZN(n25975) );
  OAI211_X2 U8661 ( .C1(n6341), .C2(n6113), .A(n29233), .B(n29739), .ZN(n20786) );
  NAND3_X1 U8668 ( .A1(n5084), .A2(n5083), .A3(n6484), .ZN(n5082) );
  NAND2_X1 U8669 ( .A1(n23426), .A2(n23339), .ZN(n6197) );
  NAND3_X1 U8697 ( .A1(n4133), .A2(n26816), .A3(n29389), .ZN(n4925) );
  NAND3_X1 U8726 ( .A1(n3440), .A2(n623), .A3(n3439), .ZN(n1729) );
  NAND2_X1 U8740 ( .A1(n4545), .A2(n521), .ZN(n3440) );
  NAND2_X1 U8741 ( .A1(n29390), .A2(n1202), .ZN(n23967) );
  NAND2_X1 U8762 ( .A1(n23965), .A2(n24582), .ZN(n29390) );
  NAND2_X1 U8772 ( .A1(n28133), .A2(n28610), .ZN(n20328) );
  NAND2_X1 U8773 ( .A1(n29391), .A2(n21163), .ZN(n20731) );
  INV_X1 U8784 ( .A(n21162), .ZN(n29391) );
  NAND2_X1 U8826 ( .A1(n21334), .A2(n21612), .ZN(n21162) );
  AND3_X2 U8833 ( .A1(n29392), .A2(n26383), .A3(n1029), .ZN(n27551) );
  NAND2_X1 U8851 ( .A1(n26379), .A2(n26425), .ZN(n29392) );
  NAND2_X1 U8856 ( .A1(n28860), .A2(n28861), .ZN(n7639) );
  NAND2_X1 U8858 ( .A1(n8611), .A2(n29394), .ZN(n29393) );
  NAND2_X1 U8885 ( .A1(n9532), .A2(n29395), .ZN(n29394) );
  OR2_X1 U8905 ( .A1(n9037), .A2(n8792), .ZN(n3353) );
  XNOR2_X1 U8906 ( .A(n19462), .B(n19299), .ZN(n19077) );
  NAND2_X2 U8916 ( .A1(n6036), .A2(n28877), .ZN(n19462) );
  NOR2_X2 U8920 ( .A1(n16988), .A2(n29396), .ZN(n19408) );
  NAND2_X1 U8932 ( .A1(n28892), .A2(n2444), .ZN(n29396) );
  AND3_X2 U8938 ( .A1(n1299), .A2(n6597), .A3(n6595), .ZN(n25928) );
  AND2_X2 U8944 ( .A1(n1462), .A2(n1460), .ZN(n21410) );
  NAND2_X1 U8955 ( .A1(n12990), .A2(n12150), .ZN(n12994) );
  INV_X1 U8984 ( .A(n10793), .ZN(n12990) );
  NAND3_X2 U8986 ( .A1(n29397), .A2(n23451), .A3(n23452), .ZN(n24972) );
  OAI21_X1 U8987 ( .B1(n23444), .B2(n23443), .A(n4794), .ZN(n29397) );
  NAND2_X1 U9007 ( .A1(n1249), .A2(n1250), .ZN(n24153) );
  NAND3_X1 U9035 ( .A1(n29398), .A2(n26210), .A3(n26209), .ZN(n29657) );
  NAND2_X1 U9049 ( .A1(n26723), .A2(n26208), .ZN(n29398) );
  OAI21_X1 U9085 ( .B1(n24248), .B2(n24523), .A(n24030), .ZN(n24006) );
  NAND2_X1 U9088 ( .A1(n28785), .A2(n24248), .ZN(n24030) );
  NAND2_X1 U9147 ( .A1(n3145), .A2(n1078), .ZN(n22681) );
  NAND2_X1 U9180 ( .A1(n3701), .A2(n18505), .ZN(n18517) );
  OAI21_X1 U9194 ( .B1(n26772), .B2(n26771), .A(n29399), .ZN(n26773) );
  NAND3_X1 U9202 ( .A1(n28421), .A2(n26768), .A3(n26935), .ZN(n29399) );
  NAND2_X1 U9227 ( .A1(n26940), .A2(n26941), .ZN(n26772) );
  XNOR2_X1 U9244 ( .A(n25134), .B(n25133), .ZN(n25136) );
  AND2_X2 U9247 ( .A1(n29401), .A2(n29400), .ZN(n25133) );
  NAND2_X1 U9255 ( .A1(n24149), .A2(n29050), .ZN(n29400) );
  NAND2_X1 U9274 ( .A1(n23935), .A2(n24744), .ZN(n29401) );
  NAND3_X1 U9291 ( .A1(n29403), .A2(n760), .A3(n29402), .ZN(n23616) );
  INV_X1 U9307 ( .A(n476), .ZN(n29403) );
  NAND2_X1 U9321 ( .A1(n29404), .A2(n19931), .ZN(n4268) );
  NAND2_X1 U9322 ( .A1(n19573), .A2(n6205), .ZN(n29404) );
  NAND2_X1 U9323 ( .A1(n23363), .A2(n23673), .ZN(n23361) );
  NAND2_X1 U9328 ( .A1(n29407), .A2(n29405), .ZN(n16602) );
  NAND2_X1 U9345 ( .A1(n17106), .A2(n29406), .ZN(n29405) );
  NAND2_X1 U9356 ( .A1(n17083), .A2(n17470), .ZN(n29407) );
  NAND3_X1 U9357 ( .A1(n29408), .A2(n28208), .A3(n4107), .ZN(n248) );
  NAND2_X1 U9359 ( .A1(n11331), .A2(n11169), .ZN(n29408) );
  XNOR2_X1 U9367 ( .A(n29409), .B(Key[13]), .ZN(Ciphertext[128]) );
  NAND2_X1 U9378 ( .A1(n96), .A2(n26341), .ZN(n29409) );
  NAND2_X1 U9384 ( .A1(n29411), .A2(n8500), .ZN(n8115) );
  INV_X1 U9482 ( .A(n8116), .ZN(n29411) );
  OAI211_X2 U9490 ( .C1(n11894), .C2(n10794), .A(n10798), .B(n29412), .ZN(
        n12088) );
  NAND2_X1 U9492 ( .A1(n10796), .A2(n11893), .ZN(n29412) );
  XNOR2_X1 U9497 ( .A(n29413), .B(n27534), .ZN(Ciphertext[58]) );
  NAND2_X1 U9499 ( .A1(n27532), .A2(n27533), .ZN(n29413) );
  NAND2_X1 U9504 ( .A1(n29415), .A2(n29414), .ZN(n7908) );
  NAND2_X1 U9528 ( .A1(n8652), .A2(n8500), .ZN(n29414) );
  NAND2_X1 U9533 ( .A1(n8655), .A2(n29416), .ZN(n29415) );
  NAND3_X1 U9535 ( .A1(n28912), .A2(n16926), .A3(n15069), .ZN(n29674) );
  NAND3_X1 U9542 ( .A1(n23584), .A2(n23710), .A3(n380), .ZN(n6154) );
  NAND2_X1 U9549 ( .A1(n29418), .A2(n29332), .ZN(n27387) );
  NOR2_X1 U9585 ( .A1(n27392), .A2(n29419), .ZN(n29418) );
  NOR2_X1 U9632 ( .A1(n25621), .A2(n6685), .ZN(n29419) );
  OAI211_X1 U9638 ( .C1(n4681), .C2(n6465), .A(n29421), .B(n29420), .ZN(n5107)
         );
  NAND2_X1 U9644 ( .A1(n4681), .A2(n17277), .ZN(n29420) );
  XNOR2_X2 U9678 ( .A(n5433), .B(n5434), .ZN(n26935) );
  NAND3_X1 U9719 ( .A1(n11705), .A2(n6073), .A3(n29422), .ZN(n3438) );
  NAND2_X1 U9729 ( .A1(n12205), .A2(n11703), .ZN(n29422) );
  NAND2_X1 U9737 ( .A1(n16791), .A2(n16792), .ZN(n17798) );
  NAND2_X1 U9774 ( .A1(n20025), .A2(n20026), .ZN(n21632) );
  OR2_X1 U9781 ( .A1(n10544), .A2(n11149), .ZN(n1064) );
  NAND2_X1 U9794 ( .A1(n24113), .A2(n24111), .ZN(n23870) );
  NOR2_X1 U9840 ( .A1(n19656), .A2(n19659), .ZN(n19606) );
  NAND3_X1 U9842 ( .A1(n7580), .A2(n7887), .A3(n7581), .ZN(n7083) );
  OAI21_X1 U9874 ( .B1(n9211), .B2(n8995), .A(n8994), .ZN(n8436) );
  NAND2_X1 U9883 ( .A1(n9211), .A2(n8996), .ZN(n8994) );
  NAND3_X1 U9888 ( .A1(n29424), .A2(n29423), .A3(n11112), .ZN(n2351) );
  NAND2_X1 U9907 ( .A1(n5109), .A2(n11111), .ZN(n29423) );
  NAND2_X1 U9909 ( .A1(n243), .A2(n242), .ZN(n29424) );
  NAND2_X1 U9917 ( .A1(n16715), .A2(n16716), .ZN(n18197) );
  OAI211_X1 U9961 ( .C1(n17196), .C2(n29546), .A(n16714), .B(n4283), .ZN(
        n16715) );
  AOI21_X1 U10012 ( .B1(n29427), .B2(n29426), .A(n20008), .ZN(n20010) );
  NAND2_X1 U10030 ( .A1(n4991), .A2(n6156), .ZN(n29427) );
  AND2_X1 U10032 ( .A1(n6309), .A2(n24726), .ZN(n4749) );
  NAND3_X1 U10059 ( .A1(n17339), .A2(n17340), .A3(n17338), .ZN(n17341) );
  OAI21_X1 U10063 ( .B1(n26532), .B2(n26528), .A(n29331), .ZN(n29168) );
  NAND2_X1 U10068 ( .A1(n29429), .A2(n29428), .ZN(n19801) );
  NAND2_X1 U10070 ( .A1(n19800), .A2(n29601), .ZN(n29428) );
  NAND2_X1 U10077 ( .A1(n19799), .A2(n1624), .ZN(n29429) );
  NAND2_X1 U10110 ( .A1(n29431), .A2(n29430), .ZN(n15767) );
  NAND2_X1 U10121 ( .A1(n532), .A2(n17316), .ZN(n29430) );
  NAND2_X1 U10139 ( .A1(n790), .A2(n17562), .ZN(n29431) );
  NOR2_X2 U10157 ( .A1(n6635), .A2(n19801), .ZN(n21465) );
  XNOR2_X1 U10159 ( .A(n29432), .B(n26287), .ZN(Ciphertext[84]) );
  OR2_X1 U10187 ( .A1(n26286), .A2(n26346), .ZN(n29433) );
  OAI21_X1 U10195 ( .B1(n325), .B2(n27711), .A(n29434), .ZN(n27713) );
  NAND2_X1 U10200 ( .A1(n325), .A2(n27716), .ZN(n29434) );
  NAND2_X1 U10207 ( .A1(n28958), .A2(n21467), .ZN(n29435) );
  OAI21_X1 U10208 ( .B1(n29437), .B2(n1931), .A(n29436), .ZN(n12106) );
  NAND2_X1 U10212 ( .A1(n12104), .A2(n1931), .ZN(n29436) );
  NOR2_X1 U10225 ( .A1(n11656), .A2(n12162), .ZN(n29437) );
  NAND3_X1 U10263 ( .A1(n23296), .A2(n29020), .A3(n22864), .ZN(n5712) );
  NAND2_X1 U10283 ( .A1(n23837), .A2(n23391), .ZN(n23281) );
  NAND3_X1 U10291 ( .A1(n8027), .A2(n8029), .A3(n8028), .ZN(n29464) );
  NAND2_X1 U10325 ( .A1(n29438), .A2(n724), .ZN(n22393) );
  NAND2_X1 U10385 ( .A1(n726), .A2(n22392), .ZN(n29438) );
  NOR2_X1 U10452 ( .A1(n27286), .A2(n27287), .ZN(n26811) );
  NOR2_X2 U10455 ( .A1(n26795), .A2(n26796), .ZN(n27287) );
  NAND3_X1 U10472 ( .A1(n8465), .A2(n8464), .A3(n8826), .ZN(n29439) );
  MUX2_X1 U10477 ( .A(n18398), .B(n18231), .S(n18233), .Z(n18235) );
  NAND4_X2 U10540 ( .A1(n4987), .A2(n4988), .A3(n5459), .A4(n5458), .ZN(n18233) );
  OR2_X2 U10546 ( .A1(n29440), .A2(n17922), .ZN(n19413) );
  AOI21_X1 U10580 ( .B1(n17919), .B2(n17920), .A(n18357), .ZN(n29440) );
  NAND3_X2 U10616 ( .A1(n29441), .A2(n5979), .A3(n5977), .ZN(n15447) );
  NAND3_X1 U10623 ( .A1(n29201), .A2(n28805), .A3(n5980), .ZN(n29441) );
  NAND2_X1 U10632 ( .A1(n26404), .A2(n29442), .ZN(n26406) );
  NAND3_X1 U10633 ( .A1(n2433), .A2(n29444), .A3(n29443), .ZN(n29442) );
  NAND2_X1 U10645 ( .A1(n27553), .A2(n27551), .ZN(n29443) );
  NAND2_X1 U10649 ( .A1(n27552), .A2(n29445), .ZN(n29444) );
  NAND2_X1 U10650 ( .A1(n1120), .A2(n1122), .ZN(n29203) );
  NAND2_X1 U10653 ( .A1(n29446), .A2(n7235), .ZN(n6382) );
  OAI21_X1 U10661 ( .B1(n7232), .B2(n6384), .A(n2833), .ZN(n29446) );
  INV_X1 U10664 ( .A(n25617), .ZN(n27394) );
  OAI211_X2 U10688 ( .C1(n19982), .C2(n18886), .A(n18884), .B(n18885), .ZN(
        n21288) );
  NAND2_X1 U10697 ( .A1(n29448), .A2(n29447), .ZN(n27666) );
  NAND2_X1 U10705 ( .A1(n27664), .A2(n27663), .ZN(n29447) );
  NAND2_X1 U10718 ( .A1(n29450), .A2(n29449), .ZN(n29448) );
  NAND2_X1 U10751 ( .A1(n27674), .A2(n28655), .ZN(n29450) );
  INV_X1 U10753 ( .A(Plaintext[169]), .ZN(n29451) );
  INV_X1 U10761 ( .A(n21971), .ZN(n22555) );
  XNOR2_X1 U10763 ( .A(n21801), .B(n20798), .ZN(n21971) );
  AND2_X2 U10764 ( .A1(n29453), .A2(n29452), .ZN(n21364) );
  NAND2_X1 U10773 ( .A1(n19240), .A2(n28489), .ZN(n29452) );
  NAND2_X1 U10785 ( .A1(n19241), .A2(n20511), .ZN(n29453) );
  NAND2_X1 U10789 ( .A1(n26373), .A2(n26266), .ZN(n29454) );
  NAND2_X1 U10818 ( .A1(n14101), .A2(n14105), .ZN(n6563) );
  NAND2_X1 U10821 ( .A1(n29455), .A2(n113), .ZN(n4803) );
  NAND2_X1 U10864 ( .A1(n112), .A2(n111), .ZN(n29455) );
  NAND2_X1 U10885 ( .A1(n21184), .A2(n21497), .ZN(n21186) );
  XNOR2_X2 U10888 ( .A(n21891), .B(n21892), .ZN(n23800) );
  NAND2_X1 U10893 ( .A1(n27386), .A2(n27410), .ZN(n27388) );
  NOR2_X2 U10927 ( .A1(n25626), .A2(n4013), .ZN(n27410) );
  OAI21_X1 U10933 ( .B1(n23342), .B2(n23428), .A(n29456), .ZN(n23346) );
  NAND3_X1 U10938 ( .A1(n23341), .A2(n23340), .A3(n28570), .ZN(n29456) );
  OAI21_X1 U10959 ( .B1(n530), .B2(n29636), .A(n29457), .ZN(n17164) );
  NAND2_X1 U10997 ( .A1(n17374), .A2(n29635), .ZN(n29457) );
  AND2_X1 U11012 ( .A1(n20158), .A2(n20157), .ZN(n19769) );
  NAND2_X1 U11013 ( .A1(n4433), .A2(n4434), .ZN(n4432) );
  NAND2_X1 U11038 ( .A1(n2777), .A2(n739), .ZN(n2774) );
  NAND2_X1 U11052 ( .A1(n19772), .A2(n19771), .ZN(n21144) );
  NAND2_X1 U11060 ( .A1(n22963), .A2(n22964), .ZN(n4672) );
  NAND3_X1 U11070 ( .A1(n23696), .A2(n23693), .A3(n4086), .ZN(n5480) );
  INV_X1 U11083 ( .A(n20814), .ZN(n21266) );
  MUX2_X1 U11114 ( .A(n20878), .B(n21269), .S(n20814), .Z(n18851) );
  NAND2_X1 U11176 ( .A1(n29459), .A2(n29458), .ZN(n798) );
  NAND2_X1 U11215 ( .A1(n26204), .A2(n26235), .ZN(n29458) );
  OR3_X1 U11224 ( .A1(n17439), .A2(n17437), .A3(n17433), .ZN(n1387) );
  OAI22_X1 U11238 ( .A1(n11228), .A2(n29461), .B1(n11232), .B2(n11231), .ZN(
        n29460) );
  NOR2_X1 U11248 ( .A1(n11229), .A2(n11896), .ZN(n29462) );
  NAND3_X1 U11296 ( .A1(n3367), .A2(n3366), .A3(n29463), .ZN(n196) );
  NAND3_X1 U11301 ( .A1(n3153), .A2(n18063), .A3(n17672), .ZN(n4347) );
  XNOR2_X1 U11334 ( .A(n26102), .B(n3256), .ZN(n26103) );
  AOI22_X2 U11352 ( .A1(n24197), .A2(n6238), .B1(n24196), .B2(n6239), .ZN(
        n26102) );
  NAND3_X2 U11361 ( .A1(n29464), .A2(n8031), .A3(n4061), .ZN(n9124) );
  OAI211_X2 U11436 ( .C1(n5382), .C2(n15105), .A(n5379), .B(n29465), .ZN(
        n16229) );
  NAND2_X1 U11506 ( .A1(n5381), .A2(n15105), .ZN(n29465) );
  NAND2_X1 U11566 ( .A1(n28725), .A2(n11964), .ZN(n29466) );
  NAND2_X1 U11595 ( .A1(n11998), .A2(n11536), .ZN(n11685) );
  AOI22_X2 U11602 ( .A1(n10552), .A2(n10551), .B1(n10550), .B2(n10461), .ZN(
        n11998) );
  AOI22_X2 U11691 ( .A1(n18973), .A2(n2096), .B1(n18974), .B2(n19060), .ZN(
        n21290) );
  BUF_X1 U11726 ( .A(n14416), .Z(n29638) );
  XOR2_X1 U11728 ( .A(n23919), .B(n23920), .Z(n29467) );
  NAND2_X1 U11731 ( .A1(n29696), .A2(n26164), .ZN(n29468) );
  OR2_X1 U11736 ( .A1(n26519), .A2(n29633), .ZN(n27690) );
  NOR2_X1 U11749 ( .A1(n26312), .A2(n6669), .ZN(n27777) );
  NAND2_X1 U11766 ( .A1(n29696), .A2(n26164), .ZN(n27463) );
  INV_X1 U11768 ( .A(n26177), .ZN(n29697) );
  XNOR2_X1 U11797 ( .A(n9856), .B(n9855), .ZN(n10983) );
  AND2_X1 U11811 ( .A1(n26337), .A2(n5485), .ZN(n29469) );
  BUF_X2 U11838 ( .A(n24078), .Z(n29470) );
  MUX2_X1 U11900 ( .A(n23900), .B(n23899), .S(n24688), .Z(n23904) );
  OAI21_X1 U11975 ( .B1(n26160), .B2(n26161), .A(n29697), .ZN(n29696) );
  XNOR2_X1 U12001 ( .A(n24910), .B(n24909), .ZN(n27191) );
  AND2_X1 U12042 ( .A1(n2263), .A2(n29472), .ZN(n28590) );
  AND2_X1 U12043 ( .A1(n2262), .A2(n29473), .ZN(n29472) );
  INV_X1 U12083 ( .A(n26724), .ZN(n29473) );
  XNOR2_X1 U12148 ( .A(n26049), .B(n26050), .ZN(n29474) );
  OR2_X1 U12155 ( .A1(n27780), .A2(n29070), .ZN(n29475) );
  XNOR2_X1 U12163 ( .A(n26049), .B(n26050), .ZN(n27110) );
  OR2_X1 U12164 ( .A1(n29649), .A2(n14278), .ZN(n4163) );
  OR2_X1 U12182 ( .A1(n15420), .A2(n15103), .ZN(n15419) );
  AND2_X1 U12228 ( .A1(n16952), .A2(n17354), .ZN(n29476) );
  XNOR2_X1 U12258 ( .A(n15638), .B(n15637), .ZN(n17354) );
  AOI22_X1 U12260 ( .A1(n6610), .A2(n23390), .B1(n6279), .B2(n23837), .ZN(
        n29477) );
  OR2_X1 U12296 ( .A1(n27310), .A2(n29478), .ZN(n29701) );
  OR2_X1 U12303 ( .A1(n29493), .A2(n27308), .ZN(n29478) );
  NAND2_X1 U12327 ( .A1(n29748), .A2(n10865), .ZN(n13552) );
  XOR2_X1 U12363 ( .A(n25258), .B(n25259), .Z(n29479) );
  NAND3_X1 U12389 ( .A1(n6627), .A2(n26759), .A3(n6626), .ZN(n29480) );
  XNOR2_X1 U12417 ( .A(n25594), .B(n25593), .ZN(n29481) );
  XOR2_X1 U12419 ( .A(n25594), .B(n25593), .Z(n29482) );
  AND2_X1 U12427 ( .A1(n23097), .A2(n2452), .ZN(n3612) );
  BUF_X2 U12429 ( .A(n27128), .Z(n397) );
  XOR2_X1 U12435 ( .A(n15665), .B(n15664), .Z(n29483) );
  AND4_X1 U12437 ( .A1(n17578), .A2(n3086), .A3(n3085), .A4(n3084), .ZN(n29484) );
  INV_X1 U12449 ( .A(n17534), .ZN(n18243) );
  OAI21_X1 U12463 ( .B1(n24607), .B2(n24606), .A(n24605), .ZN(n29485) );
  OAI21_X1 U12479 ( .B1(n24607), .B2(n24606), .A(n24605), .ZN(n25754) );
  INV_X1 U12501 ( .A(n11955), .ZN(n571) );
  OR2_X1 U12505 ( .A1(n26997), .A2(n26998), .ZN(n29486) );
  XNOR2_X2 U12506 ( .A(n25568), .B(n25567), .ZN(n26998) );
  XNOR2_X1 U12562 ( .A(n24971), .B(n24970), .ZN(n1907) );
  AND2_X1 U12568 ( .A1(n2263), .A2(n29472), .ZN(n28115) );
  BUF_X1 U12580 ( .A(n25597), .Z(n26229) );
  XNOR2_X1 U12585 ( .A(n24915), .B(n24914), .ZN(n27124) );
  INV_X1 U12625 ( .A(n24666), .ZN(n29754) );
  OAI21_X1 U12656 ( .B1(n1391), .B2(n1642), .A(n1390), .ZN(n24237) );
  OAI211_X1 U12673 ( .C1(n20641), .C2(n1908), .A(n19790), .B(n19789), .ZN(
        n21113) );
  AOI21_X1 U12675 ( .B1(n21197), .B2(n21196), .A(n21195), .ZN(n29489) );
  AOI21_X1 U12678 ( .B1(n21197), .B2(n21196), .A(n21195), .ZN(n29490) );
  AOI21_X1 U12697 ( .B1(n21197), .B2(n21196), .A(n21195), .ZN(n22428) );
  INV_X1 U12726 ( .A(n3911), .ZN(n29491) );
  BUF_X1 U12737 ( .A(n18845), .Z(n19765) );
  OR2_X1 U12782 ( .A1(n22286), .A2(n21213), .ZN(n20666) );
  MUX2_X1 U12849 ( .A(n19989), .B(n20165), .S(n19993), .Z(n19862) );
  BUF_X1 U12890 ( .A(n26717), .Z(n283) );
  NAND3_X1 U12892 ( .A1(n4516), .A2(n28), .A3(n27), .ZN(n29492) );
  NAND3_X1 U12893 ( .A1(n4516), .A2(n28), .A3(n27), .ZN(n18756) );
  OR2_X1 U12905 ( .A1(n4118), .A2(n17569), .ZN(n17228) );
  OAI211_X1 U12929 ( .C1(n11375), .C2(n11831), .A(n3685), .B(n3684), .ZN(
        n29494) );
  OAI211_X1 U12947 ( .C1(n11375), .C2(n11831), .A(n3685), .B(n3684), .ZN(
        n29495) );
  OAI211_X1 U12964 ( .C1(n11375), .C2(n11831), .A(n3685), .B(n3684), .ZN(
        n13401) );
  NAND2_X1 U12993 ( .A1(n18071), .A2(n18070), .ZN(n29496) );
  XNOR2_X1 U13016 ( .A(n25907), .B(n25906), .ZN(n29497) );
  NAND2_X1 U13017 ( .A1(n4095), .A2(n5717), .ZN(n29498) );
  NAND2_X1 U13033 ( .A1(n4095), .A2(n5717), .ZN(n29499) );
  XNOR2_X1 U13039 ( .A(n3168), .B(n25712), .ZN(n29500) );
  XNOR2_X1 U13057 ( .A(n25236), .B(n25235), .ZN(n26728) );
  AND2_X1 U13068 ( .A1(n16716), .A2(n16715), .ZN(n29502) );
  XNOR2_X1 U13089 ( .A(n25681), .B(n25396), .ZN(n25807) );
  CLKBUF_X1 U13094 ( .A(n27871), .Z(n29504) );
  BUF_X1 U13112 ( .A(n23874), .Z(n24470) );
  OAI21_X1 U13116 ( .B1(n29227), .B2(n21378), .A(n29329), .ZN(n29652) );
  XOR2_X1 U13130 ( .A(n16171), .B(n15920), .Z(n15924) );
  NAND4_X1 U13153 ( .A1(n4076), .A2(n4077), .A3(n4075), .A4(n16694), .ZN(
        n29505) );
  NAND4_X1 U13174 ( .A1(n4076), .A2(n4077), .A3(n4075), .A4(n16694), .ZN(
        n29506) );
  NAND4_X1 U13175 ( .A1(n4076), .A2(n4077), .A3(n4075), .A4(n16694), .ZN(
        n19707) );
  OAI211_X1 U13180 ( .C1(n4865), .C2(n4866), .A(n4864), .B(n29738), .ZN(n29507) );
  XNOR2_X1 U13196 ( .A(n6804), .B(n19730), .ZN(n29508) );
  OAI211_X1 U13259 ( .C1(n4865), .C2(n4866), .A(n4864), .B(n29738), .ZN(n18422) );
  XNOR2_X1 U13378 ( .A(n6804), .B(n19730), .ZN(n20437) );
  INV_X1 U13379 ( .A(n10383), .ZN(n29509) );
  CLKBUF_X1 U13386 ( .A(n28174), .Z(n29510) );
  AND2_X1 U13392 ( .A1(n1907), .A2(n26387), .ZN(n27167) );
  CLKBUF_X1 U13397 ( .A(n16449), .Z(n29511) );
  OR2_X1 U13419 ( .A1(n21303), .A2(n24745), .ZN(n29512) );
  CLKBUF_X1 U13421 ( .A(n17571), .Z(n29513) );
  OAI21_X1 U13441 ( .B1(n21336), .B2(n21337), .A(n21335), .ZN(n29514) );
  OAI21_X1 U13453 ( .B1(n21336), .B2(n21337), .A(n21335), .ZN(n22668) );
  CLKBUF_X1 U13486 ( .A(n27418), .Z(n29515) );
  XOR2_X1 U13513 ( .A(n26972), .B(n24166), .Z(Ciphertext[27]) );
  NAND2_X1 U13524 ( .A1(n856), .A2(n18274), .ZN(n19320) );
  OR2_X1 U13539 ( .A1(n5540), .A2(n6268), .ZN(n25203) );
  OAI21_X1 U13584 ( .B1(n4955), .B2(n4957), .A(n14110), .ZN(n29516) );
  MUX2_X2 U13601 ( .A(n26226), .B(n26225), .S(n25453), .Z(n28069) );
  CLKBUF_X1 U13649 ( .A(n27629), .Z(n27626) );
  AOI21_X1 U13663 ( .B1(n25241), .B2(n25240), .A(n26464), .ZN(n25242) );
  INV_X1 U13664 ( .A(n25065), .ZN(n26114) );
  BUF_X1 U13667 ( .A(n23261), .Z(n23715) );
  AND2_X2 U13668 ( .A1(n5365), .A2(n16923), .ZN(n18324) );
  XNOR2_X1 U13695 ( .A(n10430), .B(n10429), .ZN(n29517) );
  XNOR2_X1 U13699 ( .A(n10430), .B(n10429), .ZN(n11206) );
  OAI211_X2 U13700 ( .C1(n23143), .C2(n4772), .A(n3886), .B(n2058), .ZN(n24891) );
  OAI211_X1 U13780 ( .C1(n20615), .C2(n20614), .A(n20613), .B(n20612), .ZN(
        n21600) );
  XNOR2_X1 U13789 ( .A(n29485), .B(n25714), .ZN(n29518) );
  INV_X1 U13819 ( .A(n26614), .ZN(n29520) );
  AOI22_X1 U13840 ( .A1(n21115), .A2(n1897), .B1(n21114), .B2(n21463), .ZN(
        n22410) );
  CLKBUF_X1 U13871 ( .A(n19785), .Z(n29521) );
  NAND2_X1 U13888 ( .A1(n26571), .A2(n26570), .ZN(n29522) );
  NAND2_X1 U13931 ( .A1(n26571), .A2(n26570), .ZN(n29523) );
  NAND2_X1 U13952 ( .A1(n26571), .A2(n26570), .ZN(n27498) );
  XNOR2_X1 U13971 ( .A(n10282), .B(n9648), .ZN(n9748) );
  XOR2_X1 U13981 ( .A(n25518), .B(n25519), .Z(n29524) );
  AND2_X1 U13990 ( .A1(n26227), .A2(n28063), .ZN(n28055) );
  AOI21_X1 U13992 ( .B1(n20298), .B2(n19903), .A(n19902), .ZN(n21459) );
  OAI211_X1 U14000 ( .C1(n1809), .C2(n15170), .A(n14553), .B(n14552), .ZN(
        n29525) );
  OAI211_X1 U14073 ( .C1(n19058), .C2(n20056), .A(n19056), .B(n19057), .ZN(
        n29526) );
  OAI211_X1 U14123 ( .C1(n19058), .C2(n20056), .A(n19056), .B(n19057), .ZN(
        n21277) );
  XNOR2_X1 U14129 ( .A(n19100), .B(n19099), .ZN(n20484) );
  XNOR2_X1 U14131 ( .A(n24130), .B(n24131), .ZN(n29528) );
  OR2_X1 U14147 ( .A1(n26479), .A2(n26478), .ZN(n29529) );
  XNOR2_X1 U14169 ( .A(n21456), .B(n21455), .ZN(n29108) );
  NAND2_X1 U14257 ( .A1(n3551), .A2(n20301), .ZN(n29530) );
  OAI21_X2 U14276 ( .B1(n24993), .B2(n29487), .A(n24992), .ZN(n29532) );
  OAI21_X1 U14294 ( .B1(n24993), .B2(n29487), .A(n24992), .ZN(n26671) );
  AOI21_X1 U14370 ( .B1(n23204), .B2(n28596), .A(n23203), .ZN(n29533) );
  AOI21_X1 U14381 ( .B1(n23204), .B2(n28596), .A(n23203), .ZN(n29534) );
  OR2_X1 U14406 ( .A1(n28403), .A2(n27818), .ZN(n29535) );
  XNOR2_X2 U14412 ( .A(n18797), .B(n18796), .ZN(n20155) );
  BUF_X1 U14499 ( .A(n26299), .Z(n29536) );
  OAI22_X1 U14529 ( .A1(n26300), .A2(n29497), .B1(n26301), .B2(n27060), .ZN(
        n29537) );
  OAI22_X1 U14594 ( .A1(n26300), .A2(n29497), .B1(n26301), .B2(n27060), .ZN(
        n27773) );
  OR2_X1 U14652 ( .A1(n25238), .A2(n25237), .ZN(n29538) );
  OR2_X1 U14684 ( .A1(n25238), .A2(n25237), .ZN(n25998) );
  XNOR2_X1 U14689 ( .A(n16074), .B(n16073), .ZN(n29539) );
  OAI211_X1 U14734 ( .C1(n19751), .C2(n28637), .A(n4361), .B(n3443), .ZN(
        n29540) );
  XNOR2_X1 U14798 ( .A(n16074), .B(n16073), .ZN(n16541) );
  OAI211_X1 U14835 ( .C1(n19751), .C2(n28637), .A(n4361), .B(n3443), .ZN(
        n21625) );
  NAND2_X2 U14864 ( .A1(n28680), .A2(n28217), .ZN(n28015) );
  NOR2_X2 U14882 ( .A1(n25243), .A2(n25242), .ZN(n29541) );
  NOR2_X1 U14902 ( .A1(n25243), .A2(n25242), .ZN(n27371) );
  AND3_X1 U14919 ( .A1(n26453), .A2(n6736), .A3(n2043), .ZN(n27424) );
  BUF_X1 U14953 ( .A(n26119), .Z(n29543) );
  AOI22_X1 U14954 ( .A1(n23924), .A2(n24017), .B1(n459), .B2(n23923), .ZN(
        n26119) );
  OR2_X1 U15041 ( .A1(n20017), .A2(n20349), .ZN(n20513) );
  XNOR2_X1 U15049 ( .A(n20960), .B(n20959), .ZN(n29544) );
  OR2_X1 U15051 ( .A1(n21060), .A2(n21059), .ZN(n29545) );
  XNOR2_X1 U15080 ( .A(n20960), .B(n20959), .ZN(n23683) );
  INV_X1 U15085 ( .A(n7404), .ZN(n742) );
  XNOR2_X1 U15176 ( .A(n2567), .B(n15641), .ZN(n29546) );
  AND2_X1 U15220 ( .A1(n3914), .A2(n17197), .ZN(n29547) );
  AND3_X1 U15228 ( .A1(n24), .A2(n5565), .A3(n5564), .ZN(n29548) );
  AND3_X1 U15323 ( .A1(n24), .A2(n5565), .A3(n5564), .ZN(n29549) );
  AND3_X1 U15401 ( .A1(n24), .A2(n5565), .A3(n5564), .ZN(n22705) );
  XNOR2_X1 U15417 ( .A(n15748), .B(n15749), .ZN(n17313) );
  XNOR2_X1 U15419 ( .A(n18572), .B(n19649), .ZN(n29551) );
  INV_X1 U15440 ( .A(n25421), .ZN(n29552) );
  XNOR2_X1 U15468 ( .A(n18572), .B(n19649), .ZN(n28526) );
  XNOR2_X1 U15470 ( .A(n22943), .B(n22942), .ZN(n26576) );
  OR2_X1 U15471 ( .A1(n2534), .A2(n29292), .ZN(n29553) );
  NAND3_X1 U15487 ( .A1(n17325), .A2(n3248), .A3(n17326), .ZN(n29554) );
  NAND3_X1 U15490 ( .A1(n17325), .A2(n3248), .A3(n17326), .ZN(n19670) );
  OR2_X1 U15585 ( .A1(n17234), .A2(n17361), .ZN(n17044) );
  XNOR2_X2 U15658 ( .A(n18559), .B(n18560), .ZN(n20081) );
  OR3_X1 U15708 ( .A1(n11195), .A2(n4341), .A3(n12257), .ZN(n5661) );
  NOR2_X1 U15717 ( .A1(n28358), .A2(n878), .ZN(n29555) );
  NOR2_X1 U15811 ( .A1(n28358), .A2(n878), .ZN(n24395) );
  INV_X1 U15812 ( .A(n4809), .ZN(n29556) );
  OR2_X1 U15813 ( .A1(n27502), .A2(n4808), .ZN(n29557) );
  CLKBUF_X1 U15845 ( .A(n13874), .Z(n29558) );
  XNOR2_X1 U15878 ( .A(n16030), .B(n16029), .ZN(n29559) );
  XNOR2_X1 U15926 ( .A(n16030), .B(n16029), .ZN(n17102) );
  XNOR2_X1 U16094 ( .A(n25314), .B(n25313), .ZN(n29560) );
  XNOR2_X1 U16368 ( .A(n25314), .B(n25313), .ZN(n26721) );
  NOR2_X1 U16414 ( .A1(n15848), .A2(n1241), .ZN(n29561) );
  NOR2_X1 U16415 ( .A1(n20820), .A2(n20819), .ZN(n29562) );
  NOR2_X1 U16480 ( .A1(n15848), .A2(n1241), .ZN(n18060) );
  NOR2_X1 U16534 ( .A1(n20820), .A2(n20819), .ZN(n22426) );
  OAI211_X1 U16646 ( .C1(n24743), .C2(n24744), .A(n24742), .B(n24741), .ZN(
        n29563) );
  XNOR2_X1 U16912 ( .A(n12119), .B(n12118), .ZN(n29565) );
  XNOR2_X1 U16945 ( .A(n12119), .B(n12118), .ZN(n14165) );
  XNOR2_X1 U16959 ( .A(n14932), .B(n1233), .ZN(n17433) );
  OR3_X1 U17012 ( .A1(n20589), .A2(n20314), .A3(n20585), .ZN(n6931) );
  INV_X1 U17018 ( .A(n19827), .ZN(n20589) );
  NOR2_X1 U17035 ( .A1(n23009), .A2(n23008), .ZN(n29567) );
  NOR2_X1 U17047 ( .A1(n23009), .A2(n23008), .ZN(n24390) );
  XNOR2_X2 U17068 ( .A(n12502), .B(n12501), .ZN(n12534) );
  XNOR2_X1 U17100 ( .A(n6998), .B(Key[123]), .ZN(n29568) );
  INV_X1 U17152 ( .A(n28584), .ZN(n29569) );
  NOR2_X1 U17153 ( .A1(n28662), .A2(n28661), .ZN(n21587) );
  AND2_X1 U17202 ( .A1(n18060), .A2(n17671), .ZN(n18301) );
  INV_X1 U17329 ( .A(n28009), .ZN(n26984) );
  XNOR2_X1 U17330 ( .A(n25529), .B(n25530), .ZN(n29570) );
  OAI211_X1 U17339 ( .C1(n15247), .C2(n14733), .A(n14732), .B(n14731), .ZN(
        n29571) );
  XNOR2_X1 U17340 ( .A(n14749), .B(n14748), .ZN(n29572) );
  OAI211_X1 U17341 ( .C1(n15247), .C2(n14733), .A(n14732), .B(n14731), .ZN(
        n16172) );
  XNOR2_X1 U17379 ( .A(n14749), .B(n14748), .ZN(n17401) );
  XNOR2_X1 U17380 ( .A(n25093), .B(n25092), .ZN(n29573) );
  XNOR2_X1 U17428 ( .A(n3677), .B(n5828), .ZN(n29574) );
  XOR2_X1 U17465 ( .A(n25926), .B(n25925), .Z(n29575) );
  XNOR2_X1 U17542 ( .A(n9317), .B(n9316), .ZN(n29577) );
  BUF_X1 U17558 ( .A(n27573), .Z(n29578) );
  XNOR2_X1 U17671 ( .A(n9317), .B(n9316), .ZN(n10971) );
  NOR2_X1 U17739 ( .A1(n26377), .A2(n6723), .ZN(n27573) );
  XNOR2_X1 U17747 ( .A(n25502), .B(n25208), .ZN(n29579) );
  XNOR2_X1 U17750 ( .A(n25502), .B(n25208), .ZN(n26731) );
  NAND3_X2 U17751 ( .A1(n4587), .A2(n19936), .A3(n19937), .ZN(n21645) );
  OAI21_X1 U17790 ( .B1(n4954), .B2(n671), .A(n4785), .ZN(n29580) );
  AND2_X1 U17846 ( .A1(n19771), .A2(n19772), .ZN(n29581) );
  OAI21_X1 U17853 ( .B1(n4954), .B2(n671), .A(n4785), .ZN(n19463) );
  INV_X1 U18127 ( .A(n29315), .ZN(n29582) );
  XNOR2_X1 U18347 ( .A(n20839), .B(n20838), .ZN(n29583) );
  XNOR2_X2 U18717 ( .A(n25468), .B(n25469), .ZN(n26747) );
  BUF_X1 U18749 ( .A(n20053), .Z(n29584) );
  XNOR2_X1 U18761 ( .A(n6122), .B(n24900), .ZN(n29585) );
  XNOR2_X1 U18918 ( .A(n6122), .B(n24900), .ZN(n2108) );
  XOR2_X1 U18919 ( .A(n18941), .B(n18940), .Z(n29587) );
  BUF_X1 U18976 ( .A(n27026), .Z(n29588) );
  XNOR2_X1 U18980 ( .A(n13376), .B(n13377), .ZN(n29589) );
  XNOR2_X1 U18997 ( .A(n13376), .B(n13377), .ZN(n14016) );
  XOR2_X1 U19128 ( .A(n7218), .B(Key[130]), .Z(n29590) );
  OR2_X1 U19148 ( .A1(n2719), .A2(n18144), .ZN(n2720) );
  BUF_X1 U19157 ( .A(n24215), .Z(n29592) );
  AOI22_X1 U19189 ( .A1(n23646), .A2(n6378), .B1(n23565), .B2(n23564), .ZN(
        n24215) );
  BUF_X1 U19214 ( .A(n10875), .Z(n29593) );
  OAI211_X1 U19254 ( .C1(n4005), .C2(n17001), .A(n4004), .B(n6638), .ZN(n29594) );
  OAI211_X1 U19291 ( .C1(n4005), .C2(n17001), .A(n4004), .B(n6638), .ZN(n29595) );
  OAI211_X1 U19312 ( .C1(n4005), .C2(n17001), .A(n4004), .B(n6638), .ZN(n18040) );
  OR2_X1 U19353 ( .A1(n26186), .A2(n26182), .ZN(n29596) );
  INV_X1 U19372 ( .A(n469), .ZN(n29597) );
  XOR2_X1 U19444 ( .A(n16108), .B(n16109), .Z(n29598) );
  OAI21_X1 U19458 ( .B1(n24623), .B2(n28223), .A(n24621), .ZN(n29599) );
  XNOR2_X1 U19465 ( .A(n14629), .B(n14628), .ZN(n29600) );
  BUF_X1 U19489 ( .A(n20506), .Z(n29601) );
  XNOR2_X1 U19490 ( .A(n14629), .B(n14628), .ZN(n16992) );
  XNOR2_X2 U19572 ( .A(n22540), .B(n22539), .ZN(n29602) );
  XNOR2_X1 U19574 ( .A(n22540), .B(n22539), .ZN(n23831) );
  AOI21_X1 U19735 ( .B1(n16928), .B2(n29566), .A(n16927), .ZN(n29603) );
  AOI21_X1 U19755 ( .B1(n16928), .B2(n29566), .A(n16927), .ZN(n18325) );
  XNOR2_X1 U19765 ( .A(n12811), .B(n12812), .ZN(n29604) );
  XNOR2_X1 U19792 ( .A(n12811), .B(n12812), .ZN(n2728) );
  XNOR2_X1 U19800 ( .A(n15924), .B(n15923), .ZN(n29605) );
  OAI22_X1 U19812 ( .A1(n24548), .A2(n24547), .B1(n24545), .B2(n24546), .ZN(
        n29606) );
  OAI22_X1 U19913 ( .A1(n24548), .A2(n24547), .B1(n24545), .B2(n24546), .ZN(
        n25534) );
  XNOR2_X1 U19983 ( .A(n12381), .B(n12382), .ZN(n29607) );
  AND2_X2 U20011 ( .A1(n29608), .A2(n29609), .ZN(n19215) );
  AND2_X1 U20051 ( .A1(n2901), .A2(n2031), .ZN(n29608) );
  OR2_X1 U20055 ( .A1(n17632), .A2(n17834), .ZN(n29609) );
  XNOR2_X1 U20063 ( .A(n12381), .B(n12382), .ZN(n14331) );
  XNOR2_X1 U20114 ( .A(n19456), .B(n19455), .ZN(n21359) );
  XNOR2_X2 U20209 ( .A(n3649), .B(n25371), .ZN(n29610) );
  XNOR2_X1 U20261 ( .A(n3649), .B(n25371), .ZN(n26912) );
  XNOR2_X1 U20297 ( .A(n13289), .B(n13288), .ZN(n29611) );
  NOR2_X1 U20342 ( .A1(n23753), .A2(n23754), .ZN(n29612) );
  NOR2_X1 U20344 ( .A1(n23753), .A2(n23754), .ZN(n29613) );
  XNOR2_X1 U20429 ( .A(n13289), .B(n13288), .ZN(n14301) );
  NOR2_X1 U20643 ( .A1(n23753), .A2(n23754), .ZN(n26056) );
  BUF_X1 U20744 ( .A(n25913), .Z(n29614) );
  OR2_X1 U20766 ( .A1(n27898), .A2(n26510), .ZN(n29615) );
  XNOR2_X1 U20855 ( .A(n19158), .B(n19157), .ZN(n29616) );
  CLKBUF_X1 U20856 ( .A(n26194), .Z(n29617) );
  XNOR2_X1 U20857 ( .A(n19158), .B(n19157), .ZN(n20493) );
  XNOR2_X1 U20867 ( .A(n22083), .B(n22082), .ZN(n29618) );
  INV_X1 U20886 ( .A(n6150), .ZN(n29619) );
  XNOR2_X1 U20936 ( .A(n22316), .B(n22317), .ZN(n29620) );
  XNOR2_X1 U20958 ( .A(n26124), .B(n26123), .ZN(n29621) );
  XNOR2_X1 U20968 ( .A(n26124), .B(n26123), .ZN(n27140) );
  XNOR2_X1 U21035 ( .A(n25726), .B(n25725), .ZN(n29622) );
  AOI21_X1 U21194 ( .B1(n26991), .B2(n25770), .A(n25769), .ZN(n29623) );
  AND2_X1 U21198 ( .A1(n7291), .A2(n7292), .ZN(n7784) );
  OAI21_X1 U21257 ( .B1(n23535), .B2(n23534), .A(n6942), .ZN(n29624) );
  XOR2_X1 U21288 ( .A(n19684), .B(n19683), .Z(n29625) );
  XOR2_X1 U21307 ( .A(n13135), .B(n3097), .Z(n29626) );
  XNOR2_X1 U21308 ( .A(n9952), .B(n9951), .ZN(n29627) );
  CLKBUF_X1 U21322 ( .A(n14401), .Z(n29628) );
  XNOR2_X1 U21394 ( .A(Key[59]), .B(Plaintext[59]), .ZN(n8034) );
  XOR2_X1 U21431 ( .A(n16495), .B(n14760), .Z(n29630) );
  XOR2_X1 U21462 ( .A(n25171), .B(n25170), .Z(n29631) );
  BUF_X1 U21478 ( .A(n24111), .Z(n24422) );
  XNOR2_X1 U21497 ( .A(n15556), .B(n15555), .ZN(n29632) );
  XNOR2_X1 U21610 ( .A(n15556), .B(n15555), .ZN(n17344) );
  OAI22_X1 U21630 ( .A1(n23951), .A2(n23950), .B1(n5004), .B2(n24810), .ZN(
        n29634) );
  XNOR2_X1 U21634 ( .A(n16372), .B(n16371), .ZN(n29635) );
  XNOR2_X1 U21651 ( .A(n16372), .B(n16371), .ZN(n29636) );
  BUF_X1 U21689 ( .A(n11056), .Z(n29637) );
  XNOR2_X1 U21700 ( .A(n4592), .B(n9659), .ZN(n11056) );
  MUX2_X2 U21769 ( .A(n27126), .B(n27127), .S(n4109), .Z(n27759) );
  MUX2_X1 U21770 ( .A(n7800), .B(n7898), .S(n7801), .Z(n7314) );
  XNOR2_X1 U21777 ( .A(n7103), .B(Key[187]), .ZN(n7801) );
  XNOR2_X1 U21778 ( .A(n10363), .B(n9401), .ZN(n10425) );
  XNOR2_X2 U21797 ( .A(n14985), .B(n14984), .ZN(n17439) );
  XNOR2_X2 U21845 ( .A(n21942), .B(n21941), .ZN(n23789) );
  NAND4_X2 U21994 ( .A1(n17377), .A2(n16875), .A3(n16877), .A4(n16876), .ZN(
        n18507) );
  XOR2_X1 U22057 ( .A(Key[148]), .B(Plaintext[148]), .Z(n29639) );
  CLKBUF_X1 U22060 ( .A(n12554), .Z(n29640) );
  OAI211_X1 U22078 ( .C1(n23161), .C2(n23489), .A(n28844), .B(n3026), .ZN(
        n29642) );
  OAI211_X1 U22080 ( .C1(n23161), .C2(n23489), .A(n28844), .B(n3026), .ZN(
        n29643) );
  OAI211_X1 U22093 ( .C1(n23161), .C2(n23489), .A(n28844), .B(n3026), .ZN(
        n24645) );
  XOR2_X1 U22175 ( .A(n18166), .B(n18167), .Z(n29644) );
  CLKBUF_X1 U22188 ( .A(n24644), .Z(n29645) );
  OAI21_X1 U22227 ( .B1(n23175), .B2(n23174), .A(n23173), .ZN(n24644) );
  XNOR2_X1 U22228 ( .A(n2638), .B(Key[47]), .ZN(n29646) );
  NAND2_X1 U22349 ( .A1(n29774), .A2(n29741), .ZN(n29647) );
  XNOR2_X1 U22350 ( .A(n2638), .B(Key[47]), .ZN(n7129) );
  XOR2_X1 U22364 ( .A(n9753), .B(n9752), .Z(n29648) );
  AOI21_X1 U22382 ( .B1(n14358), .B2(n14273), .A(n14271), .ZN(n29649) );
  NAND2_X1 U22457 ( .A1(n24686), .A2(n24687), .ZN(n2649) );
  NAND3_X1 U22530 ( .A1(n9031), .A2(n9029), .A3(n9030), .ZN(n9032) );
  NAND2_X1 U22657 ( .A1(n149), .A2(n23901), .ZN(n148) );
  NOR2_X2 U22714 ( .A1(n29652), .A2(n29651), .ZN(n22698) );
  INV_X1 U22721 ( .A(n19188), .ZN(n29651) );
  NAND3_X1 U22733 ( .A1(n7709), .A2(n8032), .A3(n7734), .ZN(n28998) );
  NAND2_X1 U22743 ( .A1(n29653), .A2(n15372), .ZN(n15378) );
  NAND2_X1 U22788 ( .A1(n683), .A2(n15369), .ZN(n29653) );
  OR2_X1 U22791 ( .A1(n14147), .A2(n14148), .ZN(n6254) );
  NAND2_X1 U22822 ( .A1(n2302), .A2(n2303), .ZN(n13179) );
  OAI21_X1 U22876 ( .B1(n17980), .B2(n18709), .A(n29654), .ZN(n18249) );
  NAND2_X1 U22892 ( .A1(n18709), .A2(n18248), .ZN(n29654) );
  NOR2_X2 U22894 ( .A1(n13033), .A2(n29655), .ZN(n14948) );
  NAND2_X1 U22911 ( .A1(n5351), .A2(n13024), .ZN(n29655) );
  NOR2_X1 U22918 ( .A1(n1725), .A2(n14657), .ZN(n14669) );
  NAND3_X1 U23006 ( .A1(n21484), .A2(n21575), .A3(n21485), .ZN(n21486) );
  NAND3_X1 U23047 ( .A1(n3454), .A2(n10991), .A3(n10992), .ZN(n9814) );
  NAND3_X2 U23049 ( .A1(n17049), .A2(n29709), .A3(n29708), .ZN(n18333) );
  NAND2_X1 U23083 ( .A1(n17263), .A2(n16995), .ZN(n17266) );
  XNOR2_X2 U23152 ( .A(n14656), .B(n14655), .ZN(n17263) );
  NAND2_X1 U23176 ( .A1(n10702), .A2(n28310), .ZN(n10710) );
  NAND3_X1 U23177 ( .A1(n21481), .A2(n21483), .A3(n21574), .ZN(n21488) );
  NAND2_X1 U23208 ( .A1(n29316), .A2(n11321), .ZN(n11188) );
  XNOR2_X2 U23209 ( .A(n9053), .B(n9052), .ZN(n11321) );
  NAND3_X1 U23216 ( .A1(n6706), .A2(n4341), .A3(n6687), .ZN(n28863) );
  NAND3_X1 U23217 ( .A1(n14901), .A2(n14906), .A3(n14904), .ZN(n14679) );
  NAND2_X1 U23219 ( .A1(n5733), .A2(n5734), .ZN(n5732) );
  XNOR2_X1 U23284 ( .A(n29656), .B(n21946), .ZN(n21104) );
  XNOR2_X1 U23285 ( .A(n21083), .B(n6520), .ZN(n29656) );
  XNOR2_X2 U23286 ( .A(n22329), .B(n1772), .ZN(n23474) );
  OR2_X1 U23369 ( .A1(n10484), .A2(n11258), .ZN(n29722) );
  AND3_X2 U23370 ( .A1(n29657), .A2(n26213), .A3(n26212), .ZN(n27213) );
  NOR2_X1 U23439 ( .A1(n21501), .A2(n21192), .ZN(n21504) );
  NAND2_X1 U23440 ( .A1(n20380), .A2(n20379), .ZN(n29658) );
  NAND3_X1 U23453 ( .A1(n20023), .A2(n28126), .A3(n19795), .ZN(n3969) );
  NAND3_X2 U23489 ( .A1(n29194), .A2(n16807), .A3(n29195), .ZN(n18170) );
  OR2_X1 U23504 ( .A1(n5200), .A2(n5222), .ZN(n4943) );
  NAND2_X1 U23514 ( .A1(n8321), .A2(n9530), .ZN(n29660) );
  NAND2_X1 U23583 ( .A1(n8322), .A2(n29662), .ZN(n29661) );
  NAND2_X1 U23590 ( .A1(n18449), .A2(n18198), .ZN(n17746) );
  NAND3_X1 U23638 ( .A1(n13935), .A2(n293), .A3(n29320), .ZN(n642) );
  NAND2_X1 U23731 ( .A1(n14614), .A2(n14615), .ZN(n1310) );
  NAND2_X1 U23732 ( .A1(n4799), .A2(n4837), .ZN(n13705) );
  NAND2_X1 U23733 ( .A1(n4627), .A2(n13704), .ZN(n4799) );
  NAND2_X1 U23738 ( .A1(n29664), .A2(n2554), .ZN(n10591) );
  NAND2_X1 U23741 ( .A1(n11005), .A2(n5573), .ZN(n29664) );
  XNOR2_X1 U23966 ( .A(n29665), .B(n2960), .ZN(Ciphertext[137]) );
  AOI22_X1 U24053 ( .A1(n27250), .A2(n27828), .B1(n27826), .B2(n27249), .ZN(
        n29665) );
  NAND2_X1 U24062 ( .A1(n29667), .A2(n29666), .ZN(n29749) );
  INV_X1 U24080 ( .A(n3817), .ZN(n29666) );
  NAND2_X1 U24134 ( .A1(n29669), .A2(n29668), .ZN(n29667) );
  NAND2_X1 U24145 ( .A1(n3820), .A2(n10833), .ZN(n29668) );
  NAND2_X1 U24184 ( .A1(n29148), .A2(n1338), .ZN(n29669) );
  NAND2_X1 U24207 ( .A1(n28349), .A2(n29671), .ZN(n29670) );
  NAND2_X1 U24303 ( .A1(n26728), .A2(n26481), .ZN(n26726) );
  NAND2_X1 U24331 ( .A1(n189), .A2(n192), .ZN(n15349) );
  NAND2_X1 U24351 ( .A1(n7478), .A2(n29672), .ZN(n7483) );
  NAND2_X1 U24399 ( .A1(n29673), .A2(n7477), .ZN(n29672) );
  NAND2_X1 U24481 ( .A1(n7975), .A2(n8275), .ZN(n7477) );
  INV_X1 U24495 ( .A(n7976), .ZN(n29673) );
  NAND3_X1 U24620 ( .A1(n6003), .A2(n6004), .A3(n29675), .ZN(n16360) );
  NAND2_X2 U24679 ( .A1(n29676), .A2(n23927), .ZN(n25328) );
  NAND2_X1 U24751 ( .A1(n29678), .A2(n29677), .ZN(n29676) );
  NAND2_X1 U24764 ( .A1(n29512), .A2(n24751), .ZN(n29678) );
  NAND2_X2 U24828 ( .A1(n29679), .A2(n1304), .ZN(n19702) );
  OAI21_X1 U24829 ( .B1(n18448), .B2(n18097), .A(n668), .ZN(n29679) );
  OAI21_X1 U24907 ( .B1(n28086), .B2(n28087), .A(n29680), .ZN(n3517) );
  NAND3_X1 U24960 ( .A1(n91), .A2(n2021), .A3(n29681), .ZN(n29680) );
  NAND2_X1 U24961 ( .A1(n1659), .A2(n29682), .ZN(n15009) );
  XNOR2_X1 U24978 ( .A(n14921), .B(n15575), .ZN(n16320) );
  AND2_X2 U25001 ( .A1(n29684), .A2(n29683), .ZN(n15575) );
  NAND2_X1 U25002 ( .A1(n6320), .A2(n14574), .ZN(n29683) );
  NAND2_X1 U25013 ( .A1(n14573), .A2(n14572), .ZN(n29684) );
  NOR2_X1 U25017 ( .A1(n20173), .A2(n20178), .ZN(n19002) );
  NAND3_X2 U25018 ( .A1(n3282), .A2(n7294), .A3(n28696), .ZN(n8336) );
  NAND2_X1 U25037 ( .A1(n29685), .A2(n715), .ZN(n19086) );
  NAND2_X1 U25040 ( .A1(n17861), .A2(n2292), .ZN(n29685) );
  NAND2_X1 U25051 ( .A1(n29687), .A2(n29686), .ZN(n8860) );
  NAND2_X1 U25058 ( .A1(n9075), .A2(n9069), .ZN(n29686) );
  NAND2_X1 U25068 ( .A1(n8859), .A2(n28212), .ZN(n29687) );
  NAND3_X1 U25104 ( .A1(n15460), .A2(n15457), .A3(n15459), .ZN(n2745) );
  NAND3_X1 U25129 ( .A1(n13831), .A2(n13830), .A3(n29688), .ZN(n14534) );
  NAND2_X1 U25134 ( .A1(n29690), .A2(n29689), .ZN(n29688) );
  AOI21_X1 U25137 ( .B1(n14359), .B2(n14278), .A(n13832), .ZN(n29689) );
  NAND2_X1 U25225 ( .A1(n28507), .A2(n29691), .ZN(n29690) );
  NAND3_X1 U25235 ( .A1(n2684), .A2(n2683), .A3(n6281), .ZN(n2682) );
  OAI21_X1 U25264 ( .B1(n29693), .B2(n22290), .A(n29692), .ZN(n20668) );
  NAND2_X1 U25268 ( .A1(n22290), .A2(n20666), .ZN(n29692) );
  INV_X1 U25312 ( .A(n20667), .ZN(n29693) );
  NAND3_X1 U25323 ( .A1(n7711), .A2(n8029), .A3(n618), .ZN(n1032) );
  NAND2_X1 U25336 ( .A1(n7734), .A2(n7265), .ZN(n7711) );
  NOR2_X1 U25354 ( .A1(n1019), .A2(n29694), .ZN(n1389) );
  NOR2_X1 U25382 ( .A1(n28257), .A2(n60), .ZN(n29694) );
  NAND2_X1 U25383 ( .A1(n29695), .A2(n24725), .ZN(n24148) );
  INV_X1 U25430 ( .A(n6309), .ZN(n29695) );
  NAND3_X2 U25494 ( .A1(n29698), .A2(n12994), .A3(n3008), .ZN(n13386) );
  NAND2_X1 U25584 ( .A1(n10801), .A2(n12149), .ZN(n29698) );
  NAND3_X1 U25594 ( .A1(n28076), .A2(n29700), .A3(n29699), .ZN(n28079) );
  INV_X1 U25618 ( .A(n28110), .ZN(n29699) );
  NAND2_X1 U25619 ( .A1(n28109), .A2(n28794), .ZN(n29700) );
  NAND2_X1 U25626 ( .A1(n1626), .A2(n1624), .ZN(n21435) );
  NAND3_X1 U25634 ( .A1(n17105), .A2(n17104), .A3(n17103), .ZN(n18135) );
  NAND4_X1 U25638 ( .A1(n29701), .A2(n1411), .A3(n1407), .A4(n27307), .ZN(
        n1410) );
  NAND2_X1 U25706 ( .A1(n2782), .A2(n14428), .ZN(n13875) );
  AND2_X2 U25724 ( .A1(n16022), .A2(n3729), .ZN(n17762) );
  NAND2_X1 U25727 ( .A1(n4871), .A2(n29702), .ZN(n24533) );
  NAND3_X1 U25866 ( .A1(n4892), .A2(n23146), .A3(n23457), .ZN(n29702) );
  NAND3_X1 U25913 ( .A1(n29703), .A2(n1949), .A3(n4096), .ZN(n21642) );
  NAND2_X1 U25959 ( .A1(n2487), .A2(n4278), .ZN(n29703) );
  NAND2_X1 U26011 ( .A1(n29704), .A2(n20221), .ZN(n1413) );
  NAND2_X1 U26039 ( .A1(n296), .A2(n20219), .ZN(n29704) );
  NAND3_X1 U26104 ( .A1(n15087), .A2(n13989), .A3(n15083), .ZN(n13990) );
  NAND3_X1 U26105 ( .A1(n14617), .A2(n14916), .A3(n14618), .ZN(n29211) );
  OAI211_X2 U26142 ( .C1(n12010), .C2(n14250), .A(n12009), .B(n5790), .ZN(
        n14894) );
  NOR3_X1 U26177 ( .A1(n15691), .A2(n15690), .A3(n14563), .ZN(n15694) );
  NAND3_X1 U26242 ( .A1(n28677), .A2(n28676), .A3(n12990), .ZN(n29705) );
  OAI21_X1 U26243 ( .B1(n20281), .B2(n29707), .A(n29706), .ZN(n19898) );
  OR2_X1 U26287 ( .A1(n17236), .A2(n15731), .ZN(n29708) );
  NAND2_X1 U26324 ( .A1(n7410), .A2(n8925), .ZN(n8926) );
  NAND2_X1 U26328 ( .A1(n17047), .A2(n17365), .ZN(n29709) );
  NAND2_X1 U26337 ( .A1(n29712), .A2(n29711), .ZN(n29710) );
  AOI21_X1 U26373 ( .B1(n10912), .B2(n9348), .A(n10609), .ZN(n29711) );
  NAND2_X1 U26374 ( .A1(n10915), .A2(n29078), .ZN(n29712) );
  NAND2_X1 U26414 ( .A1(n10898), .A2(n12361), .ZN(n870) );
  NAND3_X1 U26432 ( .A1(n3519), .A2(n4950), .A3(n28609), .ZN(n28888) );
  OR2_X1 U26475 ( .A1(n17428), .A2(n6013), .ZN(n14226) );
  NAND3_X1 U26487 ( .A1(n6097), .A2(n6098), .A3(n24489), .ZN(n24102) );
  OAI21_X1 U26496 ( .B1(n2018), .B2(n4586), .A(n29713), .ZN(n13596) );
  NAND3_X1 U26544 ( .A1(n4586), .A2(n14376), .A3(n2849), .ZN(n29713) );
  NAND2_X1 U26546 ( .A1(n29714), .A2(n2594), .ZN(n20675) );
  NAND2_X1 U26547 ( .A1(n20007), .A2(n20623), .ZN(n29714) );
  NAND2_X1 U26572 ( .A1(n11580), .A2(n11954), .ZN(n12260) );
  NAND4_X2 U26583 ( .A1(n29715), .A2(n17443), .A3(n17445), .A4(n17444), .ZN(
        n19468) );
  NAND2_X1 U26840 ( .A1(n15466), .A2(n15463), .ZN(n4734) );
  NAND4_X2 U26853 ( .A1(n3228), .A2(n4500), .A3(n13870), .A4(n13869), .ZN(
        n15466) );
  NAND3_X1 U26854 ( .A1(n3934), .A2(n11162), .A3(n3935), .ZN(n4037) );
  NOR2_X2 U26855 ( .A1(n20675), .A2(n20670), .ZN(n21394) );
  NAND3_X1 U26873 ( .A1(n10523), .A2(n11269), .A3(n11275), .ZN(n11270) );
  NAND2_X1 U26884 ( .A1(n29717), .A2(n29716), .ZN(n15590) );
  NAND2_X1 U26903 ( .A1(n15581), .A2(n17339), .ZN(n29716) );
  NAND2_X1 U26904 ( .A1(n15582), .A2(n29718), .ZN(n29717) );
  INV_X1 U26905 ( .A(n17339), .ZN(n29718) );
  OR2_X2 U26908 ( .A1(n4887), .A2(n19869), .ZN(n20857) );
  NAND2_X1 U26909 ( .A1(n9000), .A2(n9001), .ZN(n4303) );
  NAND2_X1 U26918 ( .A1(n9200), .A2(n329), .ZN(n9001) );
  NAND2_X1 U26935 ( .A1(n29719), .A2(n2232), .ZN(n12019) );
  NAND2_X1 U26958 ( .A1(n12018), .A2(n12017), .ZN(n29719) );
  NAND2_X1 U27024 ( .A1(n15), .A2(n1416), .ZN(n9786) );
  NAND2_X1 U27030 ( .A1(n8044), .A2(n8139), .ZN(n8045) );
  NAND3_X1 U27040 ( .A1(n16915), .A2(n186), .A3(n16914), .ZN(n18326) );
  BUF_X2 U27050 ( .A(n25908), .Z(n28771) );
  NAND2_X1 U27062 ( .A1(n29721), .A2(n29720), .ZN(n8801) );
  NAND2_X1 U27068 ( .A1(n8288), .A2(n8289), .ZN(n29720) );
  NAND2_X1 U27079 ( .A1(n8293), .A2(n8292), .ZN(n29721) );
  NAND2_X1 U27094 ( .A1(n23758), .A2(n29131), .ZN(n23475) );
  NAND2_X1 U27108 ( .A1(n2437), .A2(n2439), .ZN(n27253) );
  AOI21_X1 U27166 ( .B1(n8214), .B2(n8215), .A(n8213), .ZN(n8220) );
  NAND2_X1 U27167 ( .A1(n7625), .A2(n8216), .ZN(n8214) );
  NAND2_X1 U27177 ( .A1(n6855), .A2(n15398), .ZN(n29290) );
  NAND2_X1 U27199 ( .A1(n29723), .A2(n29722), .ZN(n12026) );
  OAI21_X1 U27200 ( .B1(n4650), .B2(n3882), .A(n4649), .ZN(n29723) );
  XNOR2_X1 U27225 ( .A(n29724), .B(n4607), .ZN(Ciphertext[112]) );
  NAND3_X1 U27252 ( .A1(n26147), .A2(n26148), .A3(n6952), .ZN(n29724) );
  AOI22_X2 U27273 ( .A1(n7874), .A2(n5360), .B1(n7875), .B2(n7959), .ZN(n8116)
         );
  NAND3_X1 U27331 ( .A1(n403), .A2(n29727), .A3(n29725), .ZN(n24349) );
  NAND2_X1 U27361 ( .A1(n29128), .A2(n29726), .ZN(n29725) );
  NAND2_X1 U27362 ( .A1(n14922), .A2(n14621), .ZN(n14706) );
  NAND2_X1 U27378 ( .A1(n29728), .A2(n28934), .ZN(n7558) );
  NAND2_X1 U27380 ( .A1(n28933), .A2(n29119), .ZN(n29728) );
  NAND3_X1 U27381 ( .A1(n29150), .A2(n11113), .A3(n10461), .ZN(n2868) );
  NAND3_X1 U27387 ( .A1(n382), .A2(n383), .A3(n19997), .ZN(n6452) );
  NAND3_X1 U27404 ( .A1(n7947), .A2(n8257), .A3(n8258), .ZN(n7467) );
  NAND2_X1 U27411 ( .A1(n22457), .A2(n29729), .ZN(n24610) );
  AND2_X2 U27495 ( .A1(n5342), .A2(n29730), .ZN(n15311) );
  NAND2_X1 U27499 ( .A1(n28273), .A2(n28351), .ZN(n29730) );
  AND3_X2 U27514 ( .A1(n14387), .A2(n14388), .A3(n14389), .ZN(n16443) );
  NAND2_X2 U27622 ( .A1(n29731), .A2(n5280), .ZN(n12181) );
  NAND2_X1 U27635 ( .A1(n5278), .A2(n5277), .ZN(n29731) );
  OAI211_X2 U27650 ( .C1(n24292), .C2(n24291), .A(n24290), .B(n24289), .ZN(
        n25890) );
  OAI21_X1 U27651 ( .B1(n13720), .B2(n13587), .A(n29732), .ZN(n13898) );
  NAND2_X1 U27747 ( .A1(n13587), .A2(n28569), .ZN(n29732) );
  AOI22_X1 U27808 ( .A1(n21861), .A2(n23779), .B1(n23514), .B2(n21862), .ZN(
        n29733) );
  NAND3_X1 U27809 ( .A1(n11905), .A2(n12430), .A3(n29734), .ZN(n11912) );
  NAND2_X1 U27846 ( .A1(n12429), .A2(n29735), .ZN(n29734) );
  NAND2_X1 U27874 ( .A1(n8351), .A2(n8077), .ZN(n8078) );
  OR2_X2 U27875 ( .A1(n7799), .A2(n7798), .ZN(n8077) );
  NAND3_X1 U27904 ( .A1(n20330), .A2(n1881), .A3(n20623), .ZN(n20331) );
  OAI22_X1 U27910 ( .A1(n26616), .A2(n28228), .B1(n29736), .B2(n922), .ZN(
        n26502) );
  NAND2_X1 U27945 ( .A1(n28452), .A2(n26614), .ZN(n29736) );
  NAND3_X1 U28102 ( .A1(n28800), .A2(n17467), .A3(n29737), .ZN(n3981) );
  NAND2_X1 U28105 ( .A1(n968), .A2(n17018), .ZN(n29738) );
  OR2_X1 U28108 ( .A1(n23010), .A2(n29583), .ZN(n23012) );
  NOR2_X2 U28132 ( .A1(n10590), .A2(n10591), .ZN(n12363) );
  NAND2_X1 U28136 ( .A1(n23020), .A2(n24691), .ZN(n23027) );
  NAND2_X1 U28137 ( .A1(n20175), .A2(n20174), .ZN(n29739) );
  NAND2_X1 U28169 ( .A1(n29740), .A2(n18441), .ZN(n17739) );
  NAND2_X1 U28173 ( .A1(n18181), .A2(n18178), .ZN(n29740) );
  NAND2_X1 U28177 ( .A1(n29774), .A2(n29741), .ZN(n18512) );
  NAND2_X1 U28180 ( .A1(n4089), .A2(n17492), .ZN(n29741) );
  NAND3_X1 U28189 ( .A1(n596), .A2(n8984), .A3(n8983), .ZN(n8985) );
  NAND2_X1 U28190 ( .A1(n26129), .A2(n27178), .ZN(n26264) );
  AND2_X2 U28193 ( .A1(n29743), .A2(n29742), .ZN(n22374) );
  NAND2_X1 U28211 ( .A1(n21505), .A2(n21506), .ZN(n29742) );
  NAND2_X1 U28214 ( .A1(n21508), .A2(n29744), .ZN(n29743) );
  NAND2_X1 U28228 ( .A1(n21504), .A2(n28611), .ZN(n29744) );
  OAI211_X1 U28232 ( .C1(n24597), .C2(n24595), .A(n24730), .B(n29745), .ZN(
        n5654) );
  NAND2_X1 U28233 ( .A1(n29746), .A2(n24595), .ZN(n29745) );
  INV_X1 U28238 ( .A(n24596), .ZN(n29746) );
  NAND3_X2 U28239 ( .A1(n28887), .A2(n10462), .A3(n4630), .ZN(n11877) );
  NAND3_X1 U28271 ( .A1(n14729), .A2(n14733), .A3(n14730), .ZN(n14732) );
  XNOR2_X1 U28288 ( .A(n19575), .B(n19016), .ZN(n18855) );
  XNOR2_X1 U28295 ( .A(n19075), .B(n19463), .ZN(n19016) );
  NAND2_X1 U28300 ( .A1(n29747), .A2(n530), .ZN(n16877) );
  AND2_X1 U28301 ( .A1(n29636), .A2(n28775), .ZN(n29747) );
  NAND2_X1 U28306 ( .A1(n491), .A2(n20933), .ZN(n20762) );
  OAI21_X1 U28309 ( .B1(n11617), .B2(n12507), .A(n10864), .ZN(n29748) );
  NAND3_X1 U28310 ( .A1(n7309), .A2(n7601), .A3(n5149), .ZN(n5361) );
  NAND2_X1 U28311 ( .A1(n1697), .A2(n4294), .ZN(n29008) );
  INV_X1 U28312 ( .A(n10723), .ZN(n10612) );
  NAND2_X1 U28313 ( .A1(n10976), .A2(n10948), .ZN(n10723) );
  NAND2_X1 U28314 ( .A1(n10648), .A2(n12337), .ZN(n12346) );
  NAND2_X2 U28315 ( .A1(n29749), .A2(n10480), .ZN(n12337) );
  NAND2_X1 U28316 ( .A1(n29752), .A2(n29750), .ZN(n7125) );
  NAND2_X1 U28317 ( .A1(n8139), .A2(n29751), .ZN(n29750) );
  INV_X1 U28318 ( .A(n7560), .ZN(n29751) );
  NAND2_X1 U28319 ( .A1(n8041), .A2(n7560), .ZN(n29752) );
  OAI21_X1 U28320 ( .B1(n24667), .B2(n29754), .A(n29753), .ZN(n24384) );
  NAND2_X1 U28321 ( .A1(n24667), .A2(n24383), .ZN(n29753) );
  AND2_X1 U28322 ( .A1(n23006), .A2(n23162), .ZN(n23523) );
  NAND3_X1 U28323 ( .A1(n18186), .A2(n18187), .A3(n29199), .ZN(n2136) );
  NOR2_X1 U28324 ( .A1(n29755), .A2(n26066), .ZN(n26067) );
  INV_X1 U28325 ( .A(n26309), .ZN(n29755) );
  NAND2_X1 U28326 ( .A1(n26865), .A2(n29048), .ZN(n26309) );
  OAI211_X2 U28327 ( .C1(n8871), .C2(n8872), .A(n8869), .B(n8870), .ZN(n10251)
         );
  NAND3_X1 U28328 ( .A1(n28808), .A2(n8812), .A3(n8808), .ZN(n8253) );
  OAI21_X1 U28329 ( .B1(n11956), .B2(n571), .A(n29757), .ZN(n11200) );
  NAND2_X1 U28330 ( .A1(n571), .A2(n12261), .ZN(n29757) );
  NAND2_X1 U28331 ( .A1(n11175), .A2(n11174), .ZN(n11178) );
  NAND2_X1 U28332 ( .A1(n3218), .A2(n29758), .ZN(n15617) );
  NAND2_X1 U28333 ( .A1(n2497), .A2(n2495), .ZN(n29758) );
  NAND2_X1 U28334 ( .A1(n29759), .A2(n17013), .ZN(n6130) );
  NAND2_X1 U28335 ( .A1(n16790), .A2(n5714), .ZN(n29759) );
  NAND2_X1 U28336 ( .A1(n13954), .A2(n29760), .ZN(n13894) );
  NAND2_X1 U28337 ( .A1(n14216), .A2(n14217), .ZN(n13954) );
  OAI211_X2 U28338 ( .C1(n4104), .C2(n20869), .A(n28943), .B(n29761), .ZN(
        n22523) );
  NAND2_X1 U28339 ( .A1(n20866), .A2(n4104), .ZN(n29761) );
  NAND2_X1 U28340 ( .A1(n514), .A2(n18343), .ZN(n1480) );
  XNOR2_X1 U28341 ( .A(n29762), .B(n1184), .ZN(Ciphertext[116]) );
  NAND3_X1 U28342 ( .A1(n2792), .A2(n1216), .A3(n2793), .ZN(n29762) );
  NAND2_X1 U28343 ( .A1(n4035), .A2(n4036), .ZN(n4034) );
  XNOR2_X1 U28344 ( .A(n22883), .B(n22882), .ZN(n29763) );
  XNOR2_X1 U28345 ( .A(n29764), .B(n17697), .ZN(n17726) );
  XNOR2_X1 U28346 ( .A(n17690), .B(n18114), .ZN(n29764) );
  NAND2_X1 U28347 ( .A1(n5917), .A2(n10749), .ZN(n3129) );
  XNOR2_X2 U28348 ( .A(n5002), .B(n5003), .ZN(n14414) );
  OAI211_X2 U28349 ( .C1(n24807), .C2(n4335), .A(n4334), .B(n4333), .ZN(n25515) );
  OAI21_X1 U28350 ( .B1(n400), .B2(n27702), .A(n29765), .ZN(n28667) );
  INV_X1 U28351 ( .A(n2011), .ZN(n29765) );
  OR3_X1 U28352 ( .A1(n23357), .A2(n23355), .A3(n1837), .ZN(n28924) );
  NAND3_X1 U28353 ( .A1(n4306), .A2(n20603), .A3(n1915), .ZN(n5252) );
  NAND2_X1 U28354 ( .A1(n4914), .A2(n29766), .ZN(n16855) );
  INV_X1 U28355 ( .A(n16850), .ZN(n29766) );
  NAND2_X2 U28356 ( .A1(n29768), .A2(n29767), .ZN(n15464) );
  NAND3_X1 U28357 ( .A1(n2344), .A2(n28804), .A3(n2346), .ZN(n29767) );
  NAND2_X1 U28358 ( .A1(n2607), .A2(n4012), .ZN(n29768) );
  XNOR2_X1 U28359 ( .A(n29769), .B(n19686), .ZN(n4042) );
  AND2_X2 U28360 ( .A1(n5163), .A2(n5162), .ZN(n19484) );
  INV_X1 U28361 ( .A(n16574), .ZN(n16009) );
  XNOR2_X1 U28362 ( .A(n16574), .B(n16039), .ZN(n16453) );
  NOR2_X2 U28363 ( .A1(n15468), .A2(n15467), .ZN(n16574) );
  NAND2_X1 U28364 ( .A1(n29770), .A2(n7619), .ZN(n7360) );
  OAI22_X1 U28365 ( .A1(n8236), .A2(n7920), .B1(n8231), .B2(n7919), .ZN(n29770) );
  NAND3_X1 U28366 ( .A1(n19976), .A2(n6114), .A3(n504), .ZN(n4889) );
  NAND2_X1 U28367 ( .A1(n29002), .A2(n29003), .ZN(n23240) );
  AND3_X2 U28368 ( .A1(n24535), .A2(n132), .A3(n24537), .ZN(n26080) );
  NAND2_X1 U28369 ( .A1(n16866), .A2(n17824), .ZN(n16867) );
  NAND2_X1 U28370 ( .A1(n27666), .A2(n28373), .ZN(n27670) );
  NAND2_X1 U28371 ( .A1(n14285), .A2(n14084), .ZN(n4451) );
  NAND2_X1 U28372 ( .A1(n7843), .A2(n29772), .ZN(n29771) );
  OR2_X1 U28373 ( .A1(n10929), .A2(n10932), .ZN(n9467) );
  OR2_X2 U28374 ( .A1(n29773), .A2(n16545), .ZN(n16611) );
  NAND2_X1 U28375 ( .A1(n16542), .A2(n16543), .ZN(n29773) );
  OR2_X2 U28376 ( .A1(n10495), .A2(n10496), .ZN(n11869) );
  OAI21_X1 U28377 ( .B1(n16881), .B2(n17495), .A(n17062), .ZN(n29774) );
  NAND2_X1 U28378 ( .A1(n29775), .A2(n23200), .ZN(n24634) );
  OAI21_X1 U28379 ( .B1(n28955), .B2(n28954), .A(n23795), .ZN(n29775) );
  INV_X1 U28380 ( .A(n23705), .ZN(n3616) );
  NOR2_X1 U28381 ( .A1(n23707), .A2(n29776), .ZN(n23708) );
  NAND2_X1 U28382 ( .A1(n29777), .A2(n23705), .ZN(n29776) );
  NAND2_X1 U28383 ( .A1(n23706), .A2(n29618), .ZN(n23705) );
  INV_X1 U28384 ( .A(n22451), .ZN(n29777) );
  INV_X1 U28385 ( .A(n22863), .ZN(n5541) );
  NAND2_X1 U28386 ( .A1(n23297), .A2(n23831), .ZN(n22863) );
  NAND3_X2 U28387 ( .A1(n1177), .A2(n1176), .A3(n6049), .ZN(n24817) );
  NAND2_X1 U28388 ( .A1(n29781), .A2(n29779), .ZN(n1078) );
  NAND2_X1 U28389 ( .A1(n29780), .A2(n21603), .ZN(n29779) );
  NAND2_X1 U28390 ( .A1(n21605), .A2(n20721), .ZN(n29780) );
  NAND2_X1 U28391 ( .A1(n29782), .A2(n20649), .ZN(n29781) );
  INV_X1 U28392 ( .A(n21603), .ZN(n29782) );
  NAND2_X1 U28393 ( .A1(n24376), .A2(n1883), .ZN(n23093) );
  NAND2_X2 U28394 ( .A1(n23120), .A2(n23121), .ZN(n25845) );
  OR2_X1 U28395 ( .A1(n11490), .A2(n11431), .ZN(n2302) );
  AOI22_X1 U28396 ( .A1(n11429), .A2(n11428), .B1(n6482), .B2(n11794), .ZN(
        n11490) );
  XNOR2_X1 U28397 ( .A(n16252), .B(n16414), .ZN(n15625) );
  OAI211_X2 U28398 ( .C1(n15461), .C2(n15460), .A(n1702), .B(n1701), .ZN(
        n16252) );
  AND2_X2 U28399 ( .A1(n28363), .A2(n28364), .ZN(n12232) );
  XNOR2_X1 U28400 ( .A(n29784), .B(n29783), .ZN(Ciphertext[35]) );
  INV_X1 U28401 ( .A(n3516), .ZN(n29783) );
  NAND2_X1 U28402 ( .A1(n29786), .A2(n29785), .ZN(n29784) );
  NAND2_X1 U28403 ( .A1(n26706), .A2(n28592), .ZN(n29785) );
  NAND2_X1 U28404 ( .A1(n26705), .A2(n393), .ZN(n29786) );
  NAND3_X1 U28405 ( .A1(n23529), .A2(n23531), .A3(n28164), .ZN(n23532) );
  XNOR2_X2 U28406 ( .A(n20061), .B(n20062), .ZN(n28164) );
  OAI211_X2 U28407 ( .C1(n15051), .C2(n15052), .A(n29787), .B(n28872), .ZN(
        n16480) );
  XNOR2_X1 U28408 ( .A(n15870), .B(n28585), .ZN(n15871) );
  OAI21_X2 U28409 ( .B1(n15461), .B2(n14980), .A(n14798), .ZN(n28585) );
  NAND2_X1 U28410 ( .A1(n29791), .A2(n29788), .ZN(n26803) );
  NAND2_X1 U28411 ( .A1(n29790), .A2(n29789), .ZN(n29788) );
  NOR2_X1 U28412 ( .A1(n26797), .A2(n26800), .ZN(n29789) );
  NAND2_X1 U28413 ( .A1(n26798), .A2(n26799), .ZN(n29790) );
  NAND2_X1 U28414 ( .A1(n26801), .A2(n26800), .ZN(n29791) );
  NAND2_X1 U28415 ( .A1(n5961), .A2(n8527), .ZN(n5960) );
  NAND2_X1 U28416 ( .A1(n906), .A2(n29328), .ZN(n6602) );
  NAND2_X1 U28417 ( .A1(n5639), .A2(n17436), .ZN(n237) );
  OAI21_X1 U28418 ( .B1(n1930), .B2(n29793), .A(n29792), .ZN(n20662) );
  NAND2_X1 U28419 ( .A1(n1929), .A2(n29314), .ZN(n29792) );
  INV_X1 U28420 ( .A(n21472), .ZN(n29793) );
  AOI21_X1 U28421 ( .B1(n7524), .B2(n7748), .A(n7533), .ZN(n29794) );
  NAND3_X1 U28422 ( .A1(n29795), .A2(n10842), .A3(n10843), .ZN(n10845) );
  NAND2_X1 U28423 ( .A1(n1812), .A2(n11038), .ZN(n29795) );
  OAI21_X2 U28424 ( .B1(n8094), .B2(n9037), .A(n29796), .ZN(n9878) );
  NAND2_X1 U28425 ( .A1(n6092), .A2(n8792), .ZN(n29796) );
  NAND2_X1 U28426 ( .A1(n23427), .A2(n28122), .ZN(n23340) );
  NOR2_X1 U28427 ( .A1(n17611), .A2(n29797), .ZN(n18408) );
  XNOR2_X1 U28428 ( .A(n6270), .B(n13542), .ZN(n29798) );
  NAND2_X1 U28429 ( .A1(n12511), .A2(n3653), .ZN(n11994) );
  NOR2_X1 U28430 ( .A1(n1746), .A2(n12507), .ZN(n12511) );
  XNOR2_X1 U28431 ( .A(n29799), .B(n2523), .ZN(Ciphertext[164]) );
  NAND2_X1 U28432 ( .A1(n3064), .A2(n3063), .ZN(n29799) );
  AOI21_X2 U28433 ( .B1(n14219), .B2(n29800), .A(n6231), .ZN(n15333) );
  NAND2_X1 U28434 ( .A1(n3045), .A2(n6466), .ZN(n29800) );
  NAND3_X2 U28435 ( .A1(n11525), .A2(n11526), .A3(n11523), .ZN(n11982) );
  XNOR2_X1 U28436 ( .A(n29801), .B(n10346), .ZN(n9663) );
  XNOR2_X1 U28437 ( .A(n1891), .B(n3501), .ZN(n29801) );
  NOR2_X1 U28438 ( .A1(n29570), .A2(n28783), .ZN(n26633) );
  AOI22_X1 U28439 ( .A1(n19990), .A2(n20166), .B1(n385), .B2(n19991), .ZN(
        n1460) );
  NOR3_X1 U28440 ( .A1(n18372), .A2(n18337), .A3(n18370), .ZN(n17888) );
  XNOR2_X2 U28441 ( .A(n15157), .B(n15158), .ZN(n17421) );
  XNOR2_X2 U28442 ( .A(n15549), .B(n15550), .ZN(n17347) );
  NOR2_X2 U28443 ( .A1(n26638), .A2(n26639), .ZN(n29095) );
endmodule


module SPEEDY_Top ( clk, Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFF_X1 \reg_in_reg[191]  ( .D(Plaintext[191]), .CK(clk), .Q(reg_in[191]) );
  DFF_X1 \reg_in_reg[190]  ( .D(Plaintext[190]), .CK(clk), .Q(reg_in[190]) );
  DFF_X1 \reg_in_reg[189]  ( .D(Plaintext[189]), .CK(clk), .Q(reg_in[189]) );
  DFF_X1 \reg_in_reg[188]  ( .D(Plaintext[188]), .CK(clk), .Q(reg_in[188]) );
  DFF_X1 \reg_in_reg[187]  ( .D(Plaintext[187]), .CK(clk), .Q(reg_in[187]) );
  DFF_X1 \reg_in_reg[186]  ( .D(Plaintext[186]), .CK(clk), .Q(reg_in[186]) );
  DFF_X1 \reg_in_reg[185]  ( .D(Plaintext[185]), .CK(clk), .Q(reg_in[185]) );
  DFF_X1 \reg_in_reg[184]  ( .D(Plaintext[184]), .CK(clk), .Q(reg_in[184]) );
  DFF_X1 \reg_in_reg[183]  ( .D(Plaintext[183]), .CK(clk), .Q(reg_in[183]) );
  DFF_X1 \reg_in_reg[182]  ( .D(Plaintext[182]), .CK(clk), .Q(reg_in[182]) );
  DFF_X1 \reg_in_reg[181]  ( .D(Plaintext[181]), .CK(clk), .Q(reg_in[181]) );
  DFF_X1 \reg_in_reg[180]  ( .D(Plaintext[180]), .CK(clk), .Q(reg_in[180]) );
  DFF_X1 \reg_in_reg[179]  ( .D(Plaintext[179]), .CK(clk), .Q(reg_in[179]) );
  DFF_X1 \reg_in_reg[178]  ( .D(Plaintext[178]), .CK(clk), .Q(reg_in[178]) );
  DFF_X1 \reg_in_reg[177]  ( .D(Plaintext[177]), .CK(clk), .Q(reg_in[177]) );
  DFF_X1 \reg_in_reg[176]  ( .D(Plaintext[176]), .CK(clk), .Q(reg_in[176]) );
  DFF_X1 \reg_in_reg[175]  ( .D(Plaintext[175]), .CK(clk), .Q(reg_in[175]) );
  DFF_X1 \reg_in_reg[174]  ( .D(Plaintext[174]), .CK(clk), .Q(reg_in[174]) );
  DFF_X1 \reg_in_reg[173]  ( .D(Plaintext[173]), .CK(clk), .Q(reg_in[173]) );
  DFF_X1 \reg_in_reg[172]  ( .D(Plaintext[172]), .CK(clk), .Q(reg_in[172]) );
  DFF_X1 \reg_in_reg[171]  ( .D(Plaintext[171]), .CK(clk), .Q(reg_in[171]) );
  DFF_X1 \reg_in_reg[170]  ( .D(Plaintext[170]), .CK(clk), .Q(reg_in[170]) );
  DFF_X1 \reg_in_reg[169]  ( .D(Plaintext[169]), .CK(clk), .Q(reg_in[169]) );
  DFF_X1 \reg_in_reg[168]  ( .D(Plaintext[168]), .CK(clk), .Q(reg_in[168]) );
  DFF_X1 \reg_in_reg[167]  ( .D(Plaintext[167]), .CK(clk), .Q(reg_in[167]) );
  DFF_X1 \reg_in_reg[166]  ( .D(Plaintext[166]), .CK(clk), .Q(reg_in[166]) );
  DFF_X1 \reg_in_reg[165]  ( .D(Plaintext[165]), .CK(clk), .Q(reg_in[165]) );
  DFF_X1 \reg_in_reg[164]  ( .D(Plaintext[164]), .CK(clk), .Q(reg_in[164]) );
  DFF_X1 \reg_in_reg[163]  ( .D(Plaintext[163]), .CK(clk), .Q(reg_in[163]) );
  DFF_X1 \reg_in_reg[162]  ( .D(Plaintext[162]), .CK(clk), .Q(reg_in[162]) );
  DFF_X1 \reg_in_reg[161]  ( .D(Plaintext[161]), .CK(clk), .Q(reg_in[161]) );
  DFF_X1 \reg_in_reg[160]  ( .D(Plaintext[160]), .CK(clk), .Q(reg_in[160]) );
  DFF_X1 \reg_in_reg[159]  ( .D(Plaintext[159]), .CK(clk), .Q(reg_in[159]) );
  DFF_X1 \reg_in_reg[158]  ( .D(Plaintext[158]), .CK(clk), .Q(reg_in[158]) );
  DFF_X1 \reg_in_reg[157]  ( .D(Plaintext[157]), .CK(clk), .Q(reg_in[157]) );
  DFF_X1 \reg_in_reg[156]  ( .D(Plaintext[156]), .CK(clk), .Q(reg_in[156]) );
  DFF_X1 \reg_in_reg[155]  ( .D(Plaintext[155]), .CK(clk), .Q(reg_in[155]) );
  DFF_X1 \reg_in_reg[154]  ( .D(Plaintext[154]), .CK(clk), .Q(reg_in[154]) );
  DFF_X1 \reg_in_reg[153]  ( .D(Plaintext[153]), .CK(clk), .Q(reg_in[153]) );
  DFF_X1 \reg_in_reg[152]  ( .D(Plaintext[152]), .CK(clk), .Q(reg_in[152]) );
  DFF_X1 \reg_in_reg[151]  ( .D(Plaintext[151]), .CK(clk), .Q(reg_in[151]) );
  DFF_X1 \reg_in_reg[150]  ( .D(Plaintext[150]), .CK(clk), .Q(reg_in[150]) );
  DFF_X1 \reg_in_reg[149]  ( .D(Plaintext[149]), .CK(clk), .Q(reg_in[149]) );
  DFF_X1 \reg_in_reg[148]  ( .D(Plaintext[148]), .CK(clk), .Q(reg_in[148]) );
  DFF_X1 \reg_in_reg[147]  ( .D(Plaintext[147]), .CK(clk), .Q(reg_in[147]) );
  DFF_X1 \reg_in_reg[146]  ( .D(Plaintext[146]), .CK(clk), .Q(reg_in[146]) );
  DFF_X1 \reg_in_reg[145]  ( .D(Plaintext[145]), .CK(clk), .Q(reg_in[145]) );
  DFF_X1 \reg_in_reg[144]  ( .D(Plaintext[144]), .CK(clk), .Q(reg_in[144]) );
  DFF_X1 \reg_in_reg[143]  ( .D(Plaintext[143]), .CK(clk), .Q(reg_in[143]) );
  DFF_X1 \reg_in_reg[142]  ( .D(Plaintext[142]), .CK(clk), .Q(reg_in[142]) );
  DFF_X1 \reg_in_reg[141]  ( .D(Plaintext[141]), .CK(clk), .Q(reg_in[141]) );
  DFF_X1 \reg_in_reg[140]  ( .D(Plaintext[140]), .CK(clk), .Q(reg_in[140]) );
  DFF_X1 \reg_in_reg[139]  ( .D(Plaintext[139]), .CK(clk), .Q(reg_in[139]) );
  DFF_X1 \reg_in_reg[138]  ( .D(Plaintext[138]), .CK(clk), .Q(reg_in[138]) );
  DFF_X1 \reg_in_reg[137]  ( .D(Plaintext[137]), .CK(clk), .Q(reg_in[137]) );
  DFF_X1 \reg_in_reg[136]  ( .D(Plaintext[136]), .CK(clk), .Q(reg_in[136]) );
  DFF_X1 \reg_in_reg[135]  ( .D(Plaintext[135]), .CK(clk), .Q(reg_in[135]) );
  DFF_X1 \reg_in_reg[134]  ( .D(Plaintext[134]), .CK(clk), .Q(reg_in[134]) );
  DFF_X1 \reg_in_reg[133]  ( .D(Plaintext[133]), .CK(clk), .Q(reg_in[133]) );
  DFF_X1 \reg_in_reg[132]  ( .D(Plaintext[132]), .CK(clk), .Q(reg_in[132]) );
  DFF_X1 \reg_in_reg[131]  ( .D(Plaintext[131]), .CK(clk), .Q(reg_in[131]) );
  DFF_X1 \reg_in_reg[130]  ( .D(Plaintext[130]), .CK(clk), .Q(reg_in[130]) );
  DFF_X1 \reg_in_reg[129]  ( .D(Plaintext[129]), .CK(clk), .Q(reg_in[129]) );
  DFF_X1 \reg_in_reg[128]  ( .D(Plaintext[128]), .CK(clk), .Q(reg_in[128]) );
  DFF_X1 \reg_in_reg[127]  ( .D(Plaintext[127]), .CK(clk), .Q(reg_in[127]) );
  DFF_X1 \reg_in_reg[126]  ( .D(Plaintext[126]), .CK(clk), .Q(reg_in[126]) );
  DFF_X1 \reg_in_reg[125]  ( .D(Plaintext[125]), .CK(clk), .Q(reg_in[125]) );
  DFF_X1 \reg_in_reg[124]  ( .D(Plaintext[124]), .CK(clk), .Q(reg_in[124]) );
  DFF_X1 \reg_in_reg[123]  ( .D(Plaintext[123]), .CK(clk), .Q(reg_in[123]) );
  DFF_X1 \reg_in_reg[122]  ( .D(Plaintext[122]), .CK(clk), .Q(reg_in[122]) );
  DFF_X1 \reg_in_reg[121]  ( .D(Plaintext[121]), .CK(clk), .Q(reg_in[121]) );
  DFF_X1 \reg_in_reg[120]  ( .D(Plaintext[120]), .CK(clk), .Q(reg_in[120]) );
  DFF_X1 \reg_in_reg[119]  ( .D(Plaintext[119]), .CK(clk), .Q(reg_in[119]) );
  DFF_X1 \reg_in_reg[118]  ( .D(Plaintext[118]), .CK(clk), .Q(reg_in[118]) );
  DFF_X1 \reg_in_reg[117]  ( .D(Plaintext[117]), .CK(clk), .Q(reg_in[117]) );
  DFF_X1 \reg_in_reg[116]  ( .D(Plaintext[116]), .CK(clk), .Q(reg_in[116]) );
  DFF_X1 \reg_in_reg[115]  ( .D(Plaintext[115]), .CK(clk), .Q(reg_in[115]) );
  DFF_X1 \reg_in_reg[114]  ( .D(Plaintext[114]), .CK(clk), .Q(reg_in[114]) );
  DFF_X1 \reg_in_reg[113]  ( .D(Plaintext[113]), .CK(clk), .Q(reg_in[113]) );
  DFF_X1 \reg_in_reg[112]  ( .D(Plaintext[112]), .CK(clk), .Q(reg_in[112]) );
  DFF_X1 \reg_in_reg[111]  ( .D(Plaintext[111]), .CK(clk), .Q(reg_in[111]) );
  DFF_X1 \reg_in_reg[110]  ( .D(Plaintext[110]), .CK(clk), .Q(reg_in[110]) );
  DFF_X1 \reg_in_reg[109]  ( .D(Plaintext[109]), .CK(clk), .Q(reg_in[109]) );
  DFF_X1 \reg_in_reg[108]  ( .D(Plaintext[108]), .CK(clk), .Q(reg_in[108]) );
  DFF_X1 \reg_in_reg[107]  ( .D(Plaintext[107]), .CK(clk), .Q(reg_in[107]) );
  DFF_X1 \reg_in_reg[106]  ( .D(Plaintext[106]), .CK(clk), .Q(reg_in[106]) );
  DFF_X1 \reg_in_reg[105]  ( .D(Plaintext[105]), .CK(clk), .Q(reg_in[105]) );
  DFF_X1 \reg_in_reg[104]  ( .D(Plaintext[104]), .CK(clk), .Q(reg_in[104]) );
  DFF_X1 \reg_in_reg[103]  ( .D(Plaintext[103]), .CK(clk), .Q(reg_in[103]) );
  DFF_X1 \reg_in_reg[102]  ( .D(Plaintext[102]), .CK(clk), .Q(reg_in[102]) );
  DFF_X1 \reg_in_reg[101]  ( .D(Plaintext[101]), .CK(clk), .Q(reg_in[101]) );
  DFF_X1 \reg_in_reg[100]  ( .D(Plaintext[100]), .CK(clk), .Q(reg_in[100]) );
  DFF_X1 \reg_in_reg[99]  ( .D(Plaintext[99]), .CK(clk), .Q(reg_in[99]) );
  DFF_X1 \reg_in_reg[98]  ( .D(Plaintext[98]), .CK(clk), .Q(reg_in[98]) );
  DFF_X1 \reg_in_reg[97]  ( .D(Plaintext[97]), .CK(clk), .Q(reg_in[97]) );
  DFF_X1 \reg_in_reg[96]  ( .D(Plaintext[96]), .CK(clk), .Q(reg_in[96]) );
  DFF_X1 \reg_in_reg[95]  ( .D(Plaintext[95]), .CK(clk), .Q(reg_in[95]) );
  DFF_X1 \reg_in_reg[94]  ( .D(Plaintext[94]), .CK(clk), .Q(reg_in[94]) );
  DFF_X1 \reg_in_reg[93]  ( .D(Plaintext[93]), .CK(clk), .Q(reg_in[93]) );
  DFF_X1 \reg_in_reg[92]  ( .D(Plaintext[92]), .CK(clk), .Q(reg_in[92]) );
  DFF_X1 \reg_in_reg[91]  ( .D(Plaintext[91]), .CK(clk), .Q(reg_in[91]) );
  DFF_X1 \reg_in_reg[90]  ( .D(Plaintext[90]), .CK(clk), .Q(reg_in[90]) );
  DFF_X1 \reg_in_reg[89]  ( .D(Plaintext[89]), .CK(clk), .Q(reg_in[89]) );
  DFF_X1 \reg_in_reg[88]  ( .D(Plaintext[88]), .CK(clk), .Q(reg_in[88]) );
  DFF_X1 \reg_in_reg[87]  ( .D(Plaintext[87]), .CK(clk), .Q(reg_in[87]) );
  DFF_X1 \reg_in_reg[86]  ( .D(Plaintext[86]), .CK(clk), .Q(reg_in[86]) );
  DFF_X1 \reg_in_reg[85]  ( .D(Plaintext[85]), .CK(clk), .Q(reg_in[85]) );
  DFF_X1 \reg_in_reg[84]  ( .D(Plaintext[84]), .CK(clk), .Q(reg_in[84]) );
  DFF_X1 \reg_in_reg[83]  ( .D(Plaintext[83]), .CK(clk), .Q(reg_in[83]) );
  DFF_X1 \reg_in_reg[82]  ( .D(Plaintext[82]), .CK(clk), .Q(reg_in[82]) );
  DFF_X1 \reg_in_reg[81]  ( .D(Plaintext[81]), .CK(clk), .Q(reg_in[81]) );
  DFF_X1 \reg_in_reg[80]  ( .D(Plaintext[80]), .CK(clk), .Q(reg_in[80]) );
  DFF_X1 \reg_in_reg[79]  ( .D(Plaintext[79]), .CK(clk), .Q(reg_in[79]) );
  DFF_X1 \reg_in_reg[78]  ( .D(Plaintext[78]), .CK(clk), .Q(reg_in[78]) );
  DFF_X1 \reg_in_reg[77]  ( .D(Plaintext[77]), .CK(clk), .Q(reg_in[77]) );
  DFF_X1 \reg_in_reg[76]  ( .D(Plaintext[76]), .CK(clk), .Q(reg_in[76]) );
  DFF_X1 \reg_in_reg[75]  ( .D(Plaintext[75]), .CK(clk), .Q(reg_in[75]) );
  DFF_X1 \reg_in_reg[74]  ( .D(Plaintext[74]), .CK(clk), .Q(reg_in[74]) );
  DFF_X1 \reg_in_reg[73]  ( .D(Plaintext[73]), .CK(clk), .Q(reg_in[73]) );
  DFF_X1 \reg_in_reg[72]  ( .D(Plaintext[72]), .CK(clk), .Q(reg_in[72]) );
  DFF_X1 \reg_in_reg[71]  ( .D(Plaintext[71]), .CK(clk), .Q(reg_in[71]) );
  DFF_X1 \reg_in_reg[70]  ( .D(Plaintext[70]), .CK(clk), .Q(reg_in[70]) );
  DFF_X1 \reg_in_reg[69]  ( .D(Plaintext[69]), .CK(clk), .Q(reg_in[69]) );
  DFF_X1 \reg_in_reg[68]  ( .D(Plaintext[68]), .CK(clk), .Q(reg_in[68]) );
  DFF_X1 \reg_in_reg[67]  ( .D(Plaintext[67]), .CK(clk), .Q(reg_in[67]) );
  DFF_X1 \reg_in_reg[66]  ( .D(Plaintext[66]), .CK(clk), .Q(reg_in[66]) );
  DFF_X1 \reg_in_reg[65]  ( .D(Plaintext[65]), .CK(clk), .Q(reg_in[65]) );
  DFF_X1 \reg_in_reg[64]  ( .D(Plaintext[64]), .CK(clk), .Q(reg_in[64]) );
  DFF_X1 \reg_in_reg[63]  ( .D(Plaintext[63]), .CK(clk), .Q(reg_in[63]) );
  DFF_X1 \reg_in_reg[62]  ( .D(Plaintext[62]), .CK(clk), .Q(reg_in[62]) );
  DFF_X1 \reg_in_reg[61]  ( .D(Plaintext[61]), .CK(clk), .Q(reg_in[61]) );
  DFF_X1 \reg_in_reg[60]  ( .D(Plaintext[60]), .CK(clk), .Q(reg_in[60]) );
  DFF_X1 \reg_in_reg[59]  ( .D(Plaintext[59]), .CK(clk), .Q(reg_in[59]) );
  DFF_X1 \reg_in_reg[58]  ( .D(Plaintext[58]), .CK(clk), .Q(reg_in[58]) );
  DFF_X1 \reg_in_reg[57]  ( .D(Plaintext[57]), .CK(clk), .Q(reg_in[57]) );
  DFF_X1 \reg_in_reg[56]  ( .D(Plaintext[56]), .CK(clk), .Q(reg_in[56]) );
  DFF_X1 \reg_in_reg[55]  ( .D(Plaintext[55]), .CK(clk), .Q(reg_in[55]) );
  DFF_X1 \reg_in_reg[54]  ( .D(Plaintext[54]), .CK(clk), .Q(reg_in[54]) );
  DFF_X1 \reg_in_reg[53]  ( .D(Plaintext[53]), .CK(clk), .Q(reg_in[53]) );
  DFF_X1 \reg_in_reg[52]  ( .D(Plaintext[52]), .CK(clk), .Q(reg_in[52]) );
  DFF_X1 \reg_in_reg[51]  ( .D(Plaintext[51]), .CK(clk), .Q(reg_in[51]) );
  DFF_X1 \reg_in_reg[50]  ( .D(Plaintext[50]), .CK(clk), .Q(reg_in[50]) );
  DFF_X1 \reg_in_reg[49]  ( .D(Plaintext[49]), .CK(clk), .Q(reg_in[49]) );
  DFF_X1 \reg_in_reg[48]  ( .D(Plaintext[48]), .CK(clk), .Q(reg_in[48]) );
  DFF_X1 \reg_in_reg[47]  ( .D(Plaintext[47]), .CK(clk), .Q(reg_in[47]) );
  DFF_X1 \reg_in_reg[46]  ( .D(Plaintext[46]), .CK(clk), .Q(reg_in[46]) );
  DFF_X1 \reg_in_reg[45]  ( .D(Plaintext[45]), .CK(clk), .Q(reg_in[45]) );
  DFF_X1 \reg_in_reg[44]  ( .D(Plaintext[44]), .CK(clk), .Q(reg_in[44]) );
  DFF_X1 \reg_in_reg[43]  ( .D(Plaintext[43]), .CK(clk), .Q(reg_in[43]) );
  DFF_X1 \reg_in_reg[42]  ( .D(Plaintext[42]), .CK(clk), .Q(reg_in[42]) );
  DFF_X1 \reg_in_reg[41]  ( .D(Plaintext[41]), .CK(clk), .Q(reg_in[41]) );
  DFF_X1 \reg_in_reg[40]  ( .D(Plaintext[40]), .CK(clk), .Q(reg_in[40]) );
  DFF_X1 \reg_in_reg[39]  ( .D(Plaintext[39]), .CK(clk), .Q(reg_in[39]) );
  DFF_X1 \reg_in_reg[38]  ( .D(Plaintext[38]), .CK(clk), .Q(reg_in[38]) );
  DFF_X1 \reg_in_reg[37]  ( .D(Plaintext[37]), .CK(clk), .Q(reg_in[37]) );
  DFF_X1 \reg_in_reg[36]  ( .D(Plaintext[36]), .CK(clk), .Q(reg_in[36]) );
  DFF_X1 \reg_in_reg[35]  ( .D(Plaintext[35]), .CK(clk), .Q(reg_in[35]) );
  DFF_X1 \reg_in_reg[34]  ( .D(Plaintext[34]), .CK(clk), .Q(reg_in[34]) );
  DFF_X1 \reg_in_reg[33]  ( .D(Plaintext[33]), .CK(clk), .Q(reg_in[33]) );
  DFF_X1 \reg_in_reg[32]  ( .D(Plaintext[32]), .CK(clk), .Q(reg_in[32]) );
  DFF_X1 \reg_in_reg[31]  ( .D(Plaintext[31]), .CK(clk), .Q(reg_in[31]) );
  DFF_X1 \reg_in_reg[30]  ( .D(Plaintext[30]), .CK(clk), .Q(reg_in[30]) );
  DFF_X1 \reg_in_reg[29]  ( .D(Plaintext[29]), .CK(clk), .Q(reg_in[29]) );
  DFF_X1 \reg_in_reg[28]  ( .D(Plaintext[28]), .CK(clk), .Q(reg_in[28]) );
  DFF_X1 \reg_in_reg[27]  ( .D(Plaintext[27]), .CK(clk), .Q(reg_in[27]) );
  DFF_X1 \reg_in_reg[26]  ( .D(Plaintext[26]), .CK(clk), .Q(reg_in[26]) );
  DFF_X1 \reg_in_reg[25]  ( .D(Plaintext[25]), .CK(clk), .Q(reg_in[25]) );
  DFF_X1 \reg_in_reg[24]  ( .D(Plaintext[24]), .CK(clk), .Q(reg_in[24]) );
  DFF_X1 \reg_in_reg[23]  ( .D(Plaintext[23]), .CK(clk), .Q(reg_in[23]) );
  DFF_X1 \reg_in_reg[22]  ( .D(Plaintext[22]), .CK(clk), .Q(reg_in[22]) );
  DFF_X1 \reg_in_reg[21]  ( .D(Plaintext[21]), .CK(clk), .Q(reg_in[21]) );
  DFF_X1 \reg_in_reg[20]  ( .D(Plaintext[20]), .CK(clk), .Q(reg_in[20]) );
  DFF_X1 \reg_in_reg[19]  ( .D(Plaintext[19]), .CK(clk), .Q(reg_in[19]) );
  DFF_X1 \reg_in_reg[18]  ( .D(Plaintext[18]), .CK(clk), .Q(reg_in[18]) );
  DFF_X1 \reg_in_reg[17]  ( .D(Plaintext[17]), .CK(clk), .Q(reg_in[17]) );
  DFF_X1 \reg_in_reg[16]  ( .D(Plaintext[16]), .CK(clk), .Q(reg_in[16]) );
  DFF_X1 \reg_in_reg[15]  ( .D(Plaintext[15]), .CK(clk), .Q(reg_in[15]) );
  DFF_X1 \reg_in_reg[14]  ( .D(Plaintext[14]), .CK(clk), .Q(reg_in[14]) );
  DFF_X1 \reg_in_reg[13]  ( .D(Plaintext[13]), .CK(clk), .Q(reg_in[13]) );
  DFF_X1 \reg_in_reg[12]  ( .D(Plaintext[12]), .CK(clk), .Q(reg_in[12]) );
  DFF_X1 \reg_in_reg[11]  ( .D(Plaintext[11]), .CK(clk), .Q(reg_in[11]) );
  DFF_X1 \reg_in_reg[10]  ( .D(Plaintext[10]), .CK(clk), .Q(reg_in[10]) );
  DFF_X1 \reg_in_reg[9]  ( .D(Plaintext[9]), .CK(clk), .Q(reg_in[9]) );
  DFF_X1 \reg_in_reg[8]  ( .D(Plaintext[8]), .CK(clk), .Q(reg_in[8]) );
  DFF_X1 \reg_in_reg[7]  ( .D(Plaintext[7]), .CK(clk), .Q(reg_in[7]) );
  DFF_X1 \reg_in_reg[6]  ( .D(Plaintext[6]), .CK(clk), .Q(reg_in[6]) );
  DFF_X1 \reg_in_reg[5]  ( .D(Plaintext[5]), .CK(clk), .Q(reg_in[5]) );
  DFF_X1 \reg_in_reg[4]  ( .D(Plaintext[4]), .CK(clk), .Q(reg_in[4]) );
  DFF_X1 \reg_in_reg[3]  ( .D(Plaintext[3]), .CK(clk), .Q(reg_in[3]) );
  DFF_X1 \reg_in_reg[2]  ( .D(Plaintext[2]), .CK(clk), .Q(reg_in[2]) );
  DFF_X1 \reg_in_reg[1]  ( .D(Plaintext[1]), .CK(clk), .Q(reg_in[1]) );
  DFF_X1 \reg_in_reg[0]  ( .D(Plaintext[0]), .CK(clk), .Q(reg_in[0]) );
  DFF_X1 \reg_key_reg[190]  ( .D(Key[190]), .CK(clk), .Q(reg_key[190]) );
  DFF_X1 \reg_key_reg[187]  ( .D(Key[187]), .CK(clk), .Q(reg_key[187]) );
  DFF_X1 \reg_key_reg[179]  ( .D(Key[179]), .CK(clk), .Q(reg_key[179]) );
  DFF_X1 \reg_key_reg[173]  ( .D(Key[173]), .CK(clk), .Q(reg_key[173]) );
  DFF_X1 \reg_key_reg[168]  ( .D(Key[168]), .CK(clk), .Q(reg_key[168]) );
  DFF_X1 \reg_key_reg[151]  ( .D(Key[151]), .CK(clk), .Q(reg_key[151]) );
  DFF_X1 \reg_key_reg[148]  ( .D(Key[148]), .CK(clk), .Q(reg_key[148]) );
  DFF_X1 \reg_key_reg[122]  ( .D(Key[122]), .CK(clk), .Q(reg_key[122]) );
  DFF_X1 \reg_key_reg[104]  ( .D(Key[104]), .CK(clk), .Q(reg_key[104]) );
  DFF_X1 \reg_key_reg[91]  ( .D(Key[91]), .CK(clk), .Q(reg_key[91]) );
  DFF_X1 \reg_key_reg[83]  ( .D(Key[83]), .CK(clk), .Q(reg_key[83]) );
  DFF_X1 \reg_key_reg[79]  ( .D(Key[79]), .CK(clk), .Q(reg_key[79]) );
  DFF_X1 \reg_key_reg[74]  ( .D(Key[74]), .CK(clk), .Q(reg_key[74]) );
  DFF_X1 \reg_key_reg[68]  ( .D(Key[68]), .CK(clk), .Q(reg_key[68]) );
  DFF_X1 \reg_key_reg[66]  ( .D(Key[66]), .CK(clk), .Q(reg_key[66]) );
  DFF_X1 \reg_key_reg[56]  ( .D(Key[56]), .CK(clk), .Q(reg_key[56]) );
  DFF_X1 \reg_key_reg[53]  ( .D(Key[53]), .CK(clk), .Q(reg_key[53]) );
  DFF_X1 \reg_key_reg[51]  ( .D(Key[51]), .CK(clk), .Q(reg_key[51]) );
  DFF_X1 \reg_key_reg[40]  ( .D(Key[40]), .CK(clk), .Q(reg_key[40]) );
  DFF_X1 \reg_key_reg[35]  ( .D(Key[35]), .CK(clk), .Q(reg_key[35]) );
  DFF_X1 \reg_key_reg[19]  ( .D(Key[19]), .CK(clk), .Q(reg_key[19]) );
  DFF_X1 \reg_key_reg[11]  ( .D(Key[11]), .CK(clk), .Q(reg_key[11]) );
  DFF_X1 \reg_key_reg[9]  ( .D(Key[9]), .CK(clk), .Q(reg_key[9]) );
  DFF_X1 \reg_key_reg[8]  ( .D(Key[8]), .CK(clk), .Q(reg_key[8]) );
  DFF_X1 \Ciphertext_reg[191]  ( .D(reg_out[191]), .CK(clk), .Q(
        Ciphertext[191]) );
  DFF_X1 \Ciphertext_reg[190]  ( .D(reg_out[190]), .CK(clk), .Q(
        Ciphertext[190]) );
  DFF_X1 \Ciphertext_reg[189]  ( .D(reg_out[189]), .CK(clk), .Q(
        Ciphertext[189]) );
  DFF_X1 \Ciphertext_reg[187]  ( .D(reg_out[187]), .CK(clk), .Q(
        Ciphertext[187]) );
  DFF_X1 \Ciphertext_reg[186]  ( .D(reg_out[186]), .CK(clk), .Q(
        Ciphertext[186]) );
  DFF_X1 \Ciphertext_reg[185]  ( .D(reg_out[185]), .CK(clk), .Q(
        Ciphertext[185]) );
  DFF_X1 \Ciphertext_reg[184]  ( .D(reg_out[184]), .CK(clk), .Q(
        Ciphertext[184]) );
  DFF_X1 \Ciphertext_reg[183]  ( .D(reg_out[183]), .CK(clk), .Q(
        Ciphertext[183]) );
  DFF_X1 \Ciphertext_reg[182]  ( .D(reg_out[182]), .CK(clk), .Q(
        Ciphertext[182]) );
  DFF_X1 \Ciphertext_reg[181]  ( .D(reg_out[181]), .CK(clk), .Q(
        Ciphertext[181]) );
  DFF_X1 \Ciphertext_reg[180]  ( .D(reg_out[180]), .CK(clk), .Q(
        Ciphertext[180]) );
  DFF_X1 \Ciphertext_reg[179]  ( .D(reg_out[179]), .CK(clk), .Q(
        Ciphertext[179]) );
  DFF_X1 \Ciphertext_reg[178]  ( .D(reg_out[178]), .CK(clk), .Q(
        Ciphertext[178]) );
  DFF_X1 \Ciphertext_reg[177]  ( .D(reg_out[177]), .CK(clk), .Q(
        Ciphertext[177]) );
  DFF_X1 \Ciphertext_reg[176]  ( .D(reg_out[176]), .CK(clk), .Q(
        Ciphertext[176]) );
  DFF_X1 \Ciphertext_reg[175]  ( .D(reg_out[175]), .CK(clk), .Q(
        Ciphertext[175]) );
  DFF_X1 \Ciphertext_reg[174]  ( .D(reg_out[174]), .CK(clk), .Q(
        Ciphertext[174]) );
  DFF_X1 \Ciphertext_reg[173]  ( .D(reg_out[173]), .CK(clk), .Q(
        Ciphertext[173]) );
  DFF_X1 \Ciphertext_reg[172]  ( .D(reg_out[172]), .CK(clk), .Q(
        Ciphertext[172]) );
  DFF_X1 \Ciphertext_reg[171]  ( .D(reg_out[171]), .CK(clk), .Q(
        Ciphertext[171]) );
  DFF_X1 \Ciphertext_reg[170]  ( .D(reg_out[170]), .CK(clk), .Q(
        Ciphertext[170]) );
  DFF_X1 \Ciphertext_reg[169]  ( .D(reg_out[169]), .CK(clk), .Q(
        Ciphertext[169]) );
  DFF_X1 \Ciphertext_reg[167]  ( .D(reg_out[167]), .CK(clk), .Q(
        Ciphertext[167]) );
  DFF_X1 \Ciphertext_reg[166]  ( .D(reg_out[166]), .CK(clk), .Q(
        Ciphertext[166]) );
  DFF_X1 \Ciphertext_reg[165]  ( .D(reg_out[165]), .CK(clk), .Q(
        Ciphertext[165]) );
  DFF_X1 \Ciphertext_reg[164]  ( .D(reg_out[164]), .CK(clk), .Q(
        Ciphertext[164]) );
  DFF_X1 \Ciphertext_reg[163]  ( .D(reg_out[163]), .CK(clk), .Q(
        Ciphertext[163]) );
  DFF_X1 \Ciphertext_reg[162]  ( .D(reg_out[162]), .CK(clk), .Q(
        Ciphertext[162]) );
  DFF_X1 \Ciphertext_reg[161]  ( .D(reg_out[161]), .CK(clk), .Q(
        Ciphertext[161]) );
  DFF_X1 \Ciphertext_reg[160]  ( .D(reg_out[160]), .CK(clk), .Q(
        Ciphertext[160]) );
  DFF_X1 \Ciphertext_reg[159]  ( .D(reg_out[159]), .CK(clk), .Q(
        Ciphertext[159]) );
  DFF_X1 \Ciphertext_reg[158]  ( .D(reg_out[158]), .CK(clk), .Q(
        Ciphertext[158]) );
  DFF_X1 \Ciphertext_reg[157]  ( .D(reg_out[157]), .CK(clk), .Q(
        Ciphertext[157]) );
  DFF_X1 \Ciphertext_reg[156]  ( .D(reg_out[156]), .CK(clk), .Q(
        Ciphertext[156]) );
  DFF_X1 \Ciphertext_reg[155]  ( .D(reg_out[155]), .CK(clk), .Q(
        Ciphertext[155]) );
  DFF_X1 \Ciphertext_reg[154]  ( .D(reg_out[154]), .CK(clk), .Q(
        Ciphertext[154]) );
  DFF_X1 \Ciphertext_reg[153]  ( .D(reg_out[153]), .CK(clk), .Q(
        Ciphertext[153]) );
  DFF_X1 \Ciphertext_reg[152]  ( .D(reg_out[152]), .CK(clk), .Q(
        Ciphertext[152]) );
  DFF_X1 \Ciphertext_reg[150]  ( .D(reg_out[150]), .CK(clk), .Q(
        Ciphertext[150]) );
  DFF_X1 \Ciphertext_reg[149]  ( .D(reg_out[149]), .CK(clk), .Q(
        Ciphertext[149]) );
  DFF_X1 \Ciphertext_reg[147]  ( .D(reg_out[147]), .CK(clk), .Q(
        Ciphertext[147]) );
  DFF_X1 \Ciphertext_reg[146]  ( .D(reg_out[146]), .CK(clk), .Q(
        Ciphertext[146]) );
  DFF_X1 \Ciphertext_reg[145]  ( .D(reg_out[145]), .CK(clk), .Q(
        Ciphertext[145]) );
  DFF_X1 \Ciphertext_reg[144]  ( .D(reg_out[144]), .CK(clk), .Q(
        Ciphertext[144]) );
  DFF_X1 \Ciphertext_reg[143]  ( .D(reg_out[143]), .CK(clk), .Q(
        Ciphertext[143]) );
  DFF_X1 \Ciphertext_reg[142]  ( .D(reg_out[142]), .CK(clk), .Q(
        Ciphertext[142]) );
  DFF_X1 \Ciphertext_reg[141]  ( .D(reg_out[141]), .CK(clk), .Q(
        Ciphertext[141]) );
  DFF_X1 \Ciphertext_reg[139]  ( .D(reg_out[139]), .CK(clk), .Q(
        Ciphertext[139]) );
  DFF_X1 \Ciphertext_reg[138]  ( .D(reg_out[138]), .CK(clk), .Q(
        Ciphertext[138]) );
  DFF_X1 \Ciphertext_reg[137]  ( .D(reg_out[137]), .CK(clk), .Q(
        Ciphertext[137]) );
  DFF_X1 \Ciphertext_reg[136]  ( .D(reg_out[136]), .CK(clk), .Q(
        Ciphertext[136]) );
  DFF_X1 \Ciphertext_reg[135]  ( .D(reg_out[135]), .CK(clk), .Q(
        Ciphertext[135]) );
  DFF_X1 \Ciphertext_reg[134]  ( .D(reg_out[134]), .CK(clk), .Q(
        Ciphertext[134]) );
  DFF_X1 \Ciphertext_reg[133]  ( .D(reg_out[133]), .CK(clk), .Q(
        Ciphertext[133]) );
  DFF_X1 \Ciphertext_reg[132]  ( .D(reg_out[132]), .CK(clk), .Q(
        Ciphertext[132]) );
  DFF_X1 \Ciphertext_reg[131]  ( .D(reg_out[131]), .CK(clk), .Q(
        Ciphertext[131]) );
  DFF_X1 \Ciphertext_reg[130]  ( .D(reg_out[130]), .CK(clk), .Q(
        Ciphertext[130]) );
  DFF_X1 \Ciphertext_reg[129]  ( .D(reg_out[129]), .CK(clk), .Q(
        Ciphertext[129]) );
  DFF_X1 \Ciphertext_reg[128]  ( .D(reg_out[128]), .CK(clk), .Q(
        Ciphertext[128]) );
  DFF_X1 \Ciphertext_reg[127]  ( .D(reg_out[127]), .CK(clk), .Q(
        Ciphertext[127]) );
  DFF_X1 \Ciphertext_reg[126]  ( .D(reg_out[126]), .CK(clk), .Q(
        Ciphertext[126]) );
  DFF_X1 \Ciphertext_reg[125]  ( .D(reg_out[125]), .CK(clk), .Q(
        Ciphertext[125]) );
  DFF_X1 \Ciphertext_reg[124]  ( .D(reg_out[124]), .CK(clk), .Q(
        Ciphertext[124]) );
  DFF_X1 \Ciphertext_reg[123]  ( .D(reg_out[123]), .CK(clk), .Q(
        Ciphertext[123]) );
  DFF_X1 \Ciphertext_reg[122]  ( .D(reg_out[122]), .CK(clk), .Q(
        Ciphertext[122]) );
  DFF_X1 \Ciphertext_reg[120]  ( .D(reg_out[120]), .CK(clk), .Q(
        Ciphertext[120]) );
  DFF_X1 \Ciphertext_reg[119]  ( .D(reg_out[119]), .CK(clk), .Q(
        Ciphertext[119]) );
  DFF_X1 \Ciphertext_reg[118]  ( .D(reg_out[118]), .CK(clk), .Q(
        Ciphertext[118]) );
  DFF_X1 \Ciphertext_reg[117]  ( .D(reg_out[117]), .CK(clk), .Q(
        Ciphertext[117]) );
  DFF_X1 \Ciphertext_reg[116]  ( .D(reg_out[116]), .CK(clk), .Q(
        Ciphertext[116]) );
  DFF_X1 \Ciphertext_reg[115]  ( .D(reg_out[115]), .CK(clk), .Q(
        Ciphertext[115]) );
  DFF_X1 \Ciphertext_reg[114]  ( .D(reg_out[114]), .CK(clk), .Q(
        Ciphertext[114]) );
  DFF_X1 \Ciphertext_reg[113]  ( .D(reg_out[113]), .CK(clk), .Q(
        Ciphertext[113]) );
  DFF_X1 \Ciphertext_reg[112]  ( .D(reg_out[112]), .CK(clk), .Q(
        Ciphertext[112]) );
  DFF_X1 \Ciphertext_reg[110]  ( .D(reg_out[110]), .CK(clk), .Q(
        Ciphertext[110]) );
  DFF_X1 \Ciphertext_reg[109]  ( .D(reg_out[109]), .CK(clk), .Q(
        Ciphertext[109]) );
  DFF_X1 \Ciphertext_reg[107]  ( .D(reg_out[107]), .CK(clk), .Q(
        Ciphertext[107]) );
  DFF_X1 \Ciphertext_reg[106]  ( .D(reg_out[106]), .CK(clk), .Q(
        Ciphertext[106]) );
  DFF_X1 \Ciphertext_reg[104]  ( .D(reg_out[104]), .CK(clk), .Q(
        Ciphertext[104]) );
  DFF_X1 \Ciphertext_reg[103]  ( .D(reg_out[103]), .CK(clk), .Q(
        Ciphertext[103]) );
  DFF_X1 \Ciphertext_reg[101]  ( .D(reg_out[101]), .CK(clk), .Q(
        Ciphertext[101]) );
  DFF_X1 \Ciphertext_reg[100]  ( .D(reg_out[100]), .CK(clk), .Q(
        Ciphertext[100]) );
  DFF_X1 \Ciphertext_reg[99]  ( .D(reg_out[99]), .CK(clk), .Q(Ciphertext[99])
         );
  DFF_X1 \Ciphertext_reg[98]  ( .D(reg_out[98]), .CK(clk), .Q(Ciphertext[98])
         );
  DFF_X1 \Ciphertext_reg[97]  ( .D(reg_out[97]), .CK(clk), .Q(Ciphertext[97])
         );
  DFF_X1 \Ciphertext_reg[96]  ( .D(reg_out[96]), .CK(clk), .Q(Ciphertext[96])
         );
  DFF_X1 \Ciphertext_reg[95]  ( .D(reg_out[95]), .CK(clk), .Q(Ciphertext[95])
         );
  DFF_X1 \Ciphertext_reg[94]  ( .D(reg_out[94]), .CK(clk), .Q(Ciphertext[94])
         );
  DFF_X1 \Ciphertext_reg[93]  ( .D(reg_out[93]), .CK(clk), .Q(Ciphertext[93])
         );
  DFF_X1 \Ciphertext_reg[92]  ( .D(reg_out[92]), .CK(clk), .Q(Ciphertext[92])
         );
  DFF_X1 \Ciphertext_reg[91]  ( .D(reg_out[91]), .CK(clk), .Q(Ciphertext[91])
         );
  DFF_X1 \Ciphertext_reg[90]  ( .D(reg_out[90]), .CK(clk), .Q(Ciphertext[90])
         );
  DFF_X1 \Ciphertext_reg[89]  ( .D(reg_out[89]), .CK(clk), .Q(Ciphertext[89])
         );
  DFF_X1 \Ciphertext_reg[88]  ( .D(reg_out[88]), .CK(clk), .Q(Ciphertext[88])
         );
  DFF_X1 \Ciphertext_reg[87]  ( .D(reg_out[87]), .CK(clk), .Q(Ciphertext[87])
         );
  DFF_X1 \Ciphertext_reg[86]  ( .D(reg_out[86]), .CK(clk), .Q(Ciphertext[86])
         );
  DFF_X1 \Ciphertext_reg[85]  ( .D(reg_out[85]), .CK(clk), .Q(Ciphertext[85])
         );
  DFF_X1 \Ciphertext_reg[83]  ( .D(reg_out[83]), .CK(clk), .Q(Ciphertext[83])
         );
  DFF_X1 \Ciphertext_reg[82]  ( .D(reg_out[82]), .CK(clk), .Q(Ciphertext[82])
         );
  DFF_X1 \Ciphertext_reg[81]  ( .D(reg_out[81]), .CK(clk), .Q(Ciphertext[81])
         );
  DFF_X1 \Ciphertext_reg[80]  ( .D(reg_out[80]), .CK(clk), .Q(Ciphertext[80])
         );
  DFF_X1 \Ciphertext_reg[79]  ( .D(reg_out[79]), .CK(clk), .Q(Ciphertext[79])
         );
  DFF_X1 \Ciphertext_reg[78]  ( .D(reg_out[78]), .CK(clk), .Q(Ciphertext[78])
         );
  DFF_X1 \Ciphertext_reg[77]  ( .D(reg_out[77]), .CK(clk), .Q(Ciphertext[77])
         );
  DFF_X1 \Ciphertext_reg[76]  ( .D(reg_out[76]), .CK(clk), .Q(Ciphertext[76])
         );
  DFF_X1 \Ciphertext_reg[75]  ( .D(reg_out[75]), .CK(clk), .Q(Ciphertext[75])
         );
  DFF_X1 \Ciphertext_reg[74]  ( .D(reg_out[74]), .CK(clk), .Q(Ciphertext[74])
         );
  DFF_X1 \Ciphertext_reg[72]  ( .D(reg_out[72]), .CK(clk), .Q(Ciphertext[72])
         );
  DFF_X1 \Ciphertext_reg[71]  ( .D(reg_out[71]), .CK(clk), .Q(Ciphertext[71])
         );
  DFF_X1 \Ciphertext_reg[70]  ( .D(reg_out[70]), .CK(clk), .Q(Ciphertext[70])
         );
  DFF_X1 \Ciphertext_reg[69]  ( .D(reg_out[69]), .CK(clk), .Q(Ciphertext[69])
         );
  DFF_X1 \Ciphertext_reg[68]  ( .D(reg_out[68]), .CK(clk), .Q(Ciphertext[68])
         );
  DFF_X1 \Ciphertext_reg[67]  ( .D(reg_out[67]), .CK(clk), .Q(Ciphertext[67])
         );
  DFF_X1 \Ciphertext_reg[66]  ( .D(reg_out[66]), .CK(clk), .Q(Ciphertext[66])
         );
  DFF_X1 \Ciphertext_reg[65]  ( .D(reg_out[65]), .CK(clk), .Q(Ciphertext[65])
         );
  DFF_X1 \Ciphertext_reg[64]  ( .D(reg_out[64]), .CK(clk), .Q(Ciphertext[64])
         );
  DFF_X1 \Ciphertext_reg[63]  ( .D(reg_out[63]), .CK(clk), .Q(Ciphertext[63])
         );
  DFF_X1 \Ciphertext_reg[62]  ( .D(reg_out[62]), .CK(clk), .Q(Ciphertext[62])
         );
  DFF_X1 \Ciphertext_reg[61]  ( .D(reg_out[61]), .CK(clk), .Q(Ciphertext[61])
         );
  DFF_X1 \Ciphertext_reg[60]  ( .D(reg_out[60]), .CK(clk), .Q(Ciphertext[60])
         );
  DFF_X1 \Ciphertext_reg[59]  ( .D(reg_out[59]), .CK(clk), .Q(Ciphertext[59])
         );
  DFF_X1 \Ciphertext_reg[58]  ( .D(reg_out[58]), .CK(clk), .Q(Ciphertext[58])
         );
  DFF_X1 \Ciphertext_reg[57]  ( .D(reg_out[57]), .CK(clk), .Q(Ciphertext[57])
         );
  DFF_X1 \Ciphertext_reg[56]  ( .D(reg_out[56]), .CK(clk), .Q(Ciphertext[56])
         );
  DFF_X1 \Ciphertext_reg[55]  ( .D(reg_out[55]), .CK(clk), .Q(Ciphertext[55])
         );
  DFF_X1 \Ciphertext_reg[54]  ( .D(reg_out[54]), .CK(clk), .Q(Ciphertext[54])
         );
  DFF_X1 \Ciphertext_reg[53]  ( .D(reg_out[53]), .CK(clk), .Q(Ciphertext[53])
         );
  DFF_X1 \Ciphertext_reg[52]  ( .D(reg_out[52]), .CK(clk), .Q(Ciphertext[52])
         );
  DFF_X1 \Ciphertext_reg[49]  ( .D(reg_out[49]), .CK(clk), .Q(Ciphertext[49])
         );
  DFF_X1 \Ciphertext_reg[48]  ( .D(reg_out[48]), .CK(clk), .Q(Ciphertext[48])
         );
  DFF_X1 \Ciphertext_reg[47]  ( .D(reg_out[47]), .CK(clk), .Q(Ciphertext[47])
         );
  DFF_X1 \Ciphertext_reg[46]  ( .D(reg_out[46]), .CK(clk), .Q(Ciphertext[46])
         );
  DFF_X1 \Ciphertext_reg[45]  ( .D(reg_out[45]), .CK(clk), .Q(Ciphertext[45])
         );
  DFF_X1 \Ciphertext_reg[43]  ( .D(reg_out[43]), .CK(clk), .Q(Ciphertext[43])
         );
  DFF_X1 \Ciphertext_reg[42]  ( .D(reg_out[42]), .CK(clk), .Q(Ciphertext[42])
         );
  DFF_X1 \Ciphertext_reg[41]  ( .D(reg_out[41]), .CK(clk), .Q(Ciphertext[41])
         );
  DFF_X1 \Ciphertext_reg[39]  ( .D(reg_out[39]), .CK(clk), .Q(Ciphertext[39])
         );
  DFF_X1 \Ciphertext_reg[38]  ( .D(reg_out[38]), .CK(clk), .Q(Ciphertext[38])
         );
  DFF_X1 \Ciphertext_reg[37]  ( .D(reg_out[37]), .CK(clk), .Q(Ciphertext[37])
         );
  DFF_X1 \Ciphertext_reg[36]  ( .D(reg_out[36]), .CK(clk), .Q(Ciphertext[36])
         );
  DFF_X1 \Ciphertext_reg[35]  ( .D(reg_out[35]), .CK(clk), .Q(Ciphertext[35])
         );
  DFF_X1 \Ciphertext_reg[34]  ( .D(reg_out[34]), .CK(clk), .Q(Ciphertext[34])
         );
  DFF_X1 \Ciphertext_reg[33]  ( .D(reg_out[33]), .CK(clk), .Q(Ciphertext[33])
         );
  DFF_X1 \Ciphertext_reg[32]  ( .D(reg_out[32]), .CK(clk), .Q(Ciphertext[32])
         );
  DFF_X1 \Ciphertext_reg[31]  ( .D(reg_out[31]), .CK(clk), .Q(Ciphertext[31])
         );
  DFF_X1 \Ciphertext_reg[30]  ( .D(reg_out[30]), .CK(clk), .Q(Ciphertext[30])
         );
  DFF_X1 \Ciphertext_reg[29]  ( .D(reg_out[29]), .CK(clk), .Q(Ciphertext[29])
         );
  DFF_X1 \Ciphertext_reg[27]  ( .D(reg_out[27]), .CK(clk), .Q(Ciphertext[27])
         );
  DFF_X1 \Ciphertext_reg[26]  ( .D(reg_out[26]), .CK(clk), .Q(Ciphertext[26])
         );
  DFF_X1 \Ciphertext_reg[25]  ( .D(reg_out[25]), .CK(clk), .Q(Ciphertext[25])
         );
  DFF_X1 \Ciphertext_reg[24]  ( .D(reg_out[24]), .CK(clk), .Q(Ciphertext[24])
         );
  DFF_X1 \Ciphertext_reg[23]  ( .D(reg_out[23]), .CK(clk), .Q(Ciphertext[23])
         );
  DFF_X1 \Ciphertext_reg[22]  ( .D(reg_out[22]), .CK(clk), .Q(Ciphertext[22])
         );
  DFF_X1 \Ciphertext_reg[21]  ( .D(reg_out[21]), .CK(clk), .Q(Ciphertext[21])
         );
  DFF_X1 \Ciphertext_reg[20]  ( .D(reg_out[20]), .CK(clk), .Q(Ciphertext[20])
         );
  DFF_X1 \Ciphertext_reg[19]  ( .D(reg_out[19]), .CK(clk), .Q(Ciphertext[19])
         );
  DFF_X1 \Ciphertext_reg[18]  ( .D(reg_out[18]), .CK(clk), .Q(Ciphertext[18])
         );
  DFF_X1 \Ciphertext_reg[17]  ( .D(reg_out[17]), .CK(clk), .Q(Ciphertext[17])
         );
  DFF_X1 \Ciphertext_reg[16]  ( .D(reg_out[16]), .CK(clk), .Q(Ciphertext[16])
         );
  DFF_X1 \Ciphertext_reg[15]  ( .D(reg_out[15]), .CK(clk), .Q(Ciphertext[15])
         );
  DFF_X1 \Ciphertext_reg[14]  ( .D(reg_out[14]), .CK(clk), .Q(Ciphertext[14])
         );
  DFF_X1 \Ciphertext_reg[13]  ( .D(reg_out[13]), .CK(clk), .Q(Ciphertext[13])
         );
  DFF_X1 \Ciphertext_reg[12]  ( .D(reg_out[12]), .CK(clk), .Q(Ciphertext[12])
         );
  DFF_X1 \Ciphertext_reg[11]  ( .D(reg_out[11]), .CK(clk), .Q(Ciphertext[11])
         );
  DFF_X1 \Ciphertext_reg[10]  ( .D(reg_out[10]), .CK(clk), .Q(Ciphertext[10])
         );
  DFF_X1 \Ciphertext_reg[9]  ( .D(reg_out[9]), .CK(clk), .Q(Ciphertext[9]) );
  DFF_X1 \Ciphertext_reg[8]  ( .D(reg_out[8]), .CK(clk), .Q(Ciphertext[8]) );
  DFF_X1 \Ciphertext_reg[7]  ( .D(reg_out[7]), .CK(clk), .Q(Ciphertext[7]) );
  DFF_X1 \Ciphertext_reg[6]  ( .D(reg_out[6]), .CK(clk), .Q(Ciphertext[6]) );
  DFF_X1 \Ciphertext_reg[5]  ( .D(reg_out[5]), .CK(clk), .Q(Ciphertext[5]) );
  DFF_X1 \Ciphertext_reg[4]  ( .D(reg_out[4]), .CK(clk), .Q(Ciphertext[4]) );
  DFF_X1 \Ciphertext_reg[3]  ( .D(reg_out[3]), .CK(clk), .Q(Ciphertext[3]) );
  DFF_X1 \Ciphertext_reg[2]  ( .D(reg_out[2]), .CK(clk), .Q(Ciphertext[2]) );
  DFF_X1 \Ciphertext_reg[1]  ( .D(reg_out[1]), .CK(clk), .Q(Ciphertext[1]) );
  DFF_X1 \Ciphertext_reg[40]  ( .D(reg_out[40]), .CK(clk), .Q(Ciphertext[40])
         );
  DFF_X1 \reg_key_reg[49]  ( .D(Key[49]), .CK(clk), .Q(reg_key[49]) );
  DFF_X1 \reg_key_reg[147]  ( .D(Key[147]), .CK(clk), .Q(reg_key[147]) );
  DFF_X1 \Ciphertext_reg[151]  ( .D(reg_out[151]), .CK(clk), .Q(
        Ciphertext[151]) );
  DFF_X1 \reg_key_reg[1]  ( .D(Key[1]), .CK(clk), .Q(reg_key[1]) );
  DFF_X1 \reg_key_reg[176]  ( .D(Key[176]), .CK(clk), .Q(reg_key[176]) );
  DFF_X1 \reg_key_reg[159]  ( .D(Key[159]), .CK(clk), .Q(reg_key[159]) );
  DFF_X1 \reg_key_reg[155]  ( .D(Key[155]), .CK(clk), .Q(reg_key[155]) );
  DFF_X1 \Ciphertext_reg[51]  ( .D(reg_out[51]), .CK(clk), .Q(Ciphertext[51])
         );
  DFF_X1 \reg_key_reg[119]  ( .D(Key[119]), .CK(clk), .Q(reg_key[119]) );
  DFF_X1 \reg_key_reg[44]  ( .D(Key[44]), .CK(clk), .Q(reg_key[44]) );
  DFF_X1 \reg_key_reg[116]  ( .D(Key[116]), .CK(clk), .Q(reg_key[116]) );
  DFF_X1 \reg_key_reg[137]  ( .D(Key[137]), .CK(clk), .Q(reg_key[137]) );
  DFF_X1 \reg_key_reg[167]  ( .D(Key[167]), .CK(clk), .Q(reg_key[167]) );
  DFF_X1 \reg_key_reg[50]  ( .D(Key[50]), .CK(clk), .Q(reg_key[50]) );
  DFF_X1 \reg_key_reg[129]  ( .D(Key[129]), .CK(clk), .Q(reg_key[129]) );
  DFF_X1 \reg_key_reg[111]  ( .D(Key[111]), .CK(clk), .Q(reg_key[111]) );
  DFF_X1 \reg_key_reg[20]  ( .D(Key[20]), .CK(clk), .Q(reg_key[20]) );
  DFF_X1 \reg_key_reg[33]  ( .D(Key[33]), .CK(clk), .Q(reg_key[33]) );
  DFF_X1 \reg_key_reg[178]  ( .D(Key[178]), .CK(clk), .Q(reg_key[178]) );
  DFF_X1 \reg_key_reg[135]  ( .D(Key[135]), .CK(clk), .Q(reg_key[135]) );
  DFF_X1 \reg_key_reg[2]  ( .D(Key[2]), .CK(clk), .Q(reg_key[2]) );
  DFF_X1 \reg_key_reg[77]  ( .D(Key[77]), .CK(clk), .Q(reg_key[77]) );
  DFF_X1 \reg_key_reg[101]  ( .D(Key[101]), .CK(clk), .Q(reg_key[101]) );
  DFF_X1 \reg_key_reg[125]  ( .D(Key[125]), .CK(clk), .Q(reg_key[125]) );
  DFF_X1 \reg_key_reg[191]  ( .D(Key[191]), .CK(clk), .Q(reg_key[191]) );
  DFF_X1 \reg_key_reg[175]  ( .D(Key[175]), .CK(clk), .Q(reg_key[175]) );
  DFF_X1 \reg_key_reg[3]  ( .D(Key[3]), .CK(clk), .Q(reg_key[3]) );
  DFF_X1 \reg_key_reg[153]  ( .D(Key[153]), .CK(clk), .Q(reg_key[153]) );
  DFF_X1 \reg_key_reg[32]  ( .D(Key[32]), .CK(clk), .Q(reg_key[32]) );
  DFF_X1 \reg_key_reg[112]  ( .D(Key[112]), .CK(clk), .Q(reg_key[112]) );
  DFF_X1 \reg_key_reg[80]  ( .D(Key[80]), .CK(clk), .Q(reg_key[80]) );
  DFF_X1 \reg_key_reg[150]  ( .D(Key[150]), .CK(clk), .Q(reg_key[150]) );
  DFF_X1 \reg_key_reg[107]  ( .D(Key[107]), .CK(clk), .Q(reg_key[107]) );
  DFF_X1 \reg_key_reg[98]  ( .D(Key[98]), .CK(clk), .Q(reg_key[98]) );
  DFF_X1 \reg_key_reg[87]  ( .D(Key[87]), .CK(clk), .Q(reg_key[87]) );
  DFF_X1 \reg_key_reg[189]  ( .D(Key[189]), .CK(clk), .Q(reg_key[189]) );
  DFF_X1 \reg_key_reg[174]  ( .D(Key[174]), .CK(clk), .Q(reg_key[174]) );
  DFF_X1 \reg_key_reg[28]  ( .D(Key[28]), .CK(clk), .Q(reg_key[28]) );
  DFF_X1 \reg_key_reg[26]  ( .D(Key[26]), .CK(clk), .Q(reg_key[26]) );
  DFF_X1 \reg_key_reg[134]  ( .D(Key[134]), .CK(clk), .Q(reg_key[134]) );
  DFF_X1 \reg_key_reg[70]  ( .D(Key[70]), .CK(clk), .Q(reg_key[70]) );
  DFF_X1 \reg_key_reg[177]  ( .D(Key[177]), .CK(clk), .Q(reg_key[177]) );
  DFF_X1 \reg_key_reg[82]  ( .D(Key[82]), .CK(clk), .Q(reg_key[82]) );
  DFF_X1 \reg_key_reg[92]  ( .D(Key[92]), .CK(clk), .Q(reg_key[92]) );
  DFF_X1 \reg_key_reg[140]  ( .D(Key[140]), .CK(clk), .Q(reg_key[140]) );
  DFF_X1 \reg_key_reg[57]  ( .D(Key[57]), .CK(clk), .Q(reg_key[57]) );
  DFF_X1 \reg_key_reg[183]  ( .D(Key[183]), .CK(clk), .Q(reg_key[183]) );
  DFF_X1 \reg_key_reg[171]  ( .D(Key[171]), .CK(clk), .Q(reg_key[171]) );
  DFF_X1 \reg_key_reg[152]  ( .D(Key[152]), .CK(clk), .Q(reg_key[152]) );
  DFF_X1 \reg_key_reg[108]  ( .D(Key[108]), .CK(clk), .Q(reg_key[108]) );
  DFF_X1 \reg_key_reg[41]  ( .D(Key[41]), .CK(clk), .Q(reg_key[41]) );
  DFF_X1 \reg_key_reg[130]  ( .D(Key[130]), .CK(clk), .Q(reg_key[130]) );
  DFF_X1 \reg_key_reg[27]  ( .D(Key[27]), .CK(clk), .Q(reg_key[27]) );
  DFF_X1 \reg_key_reg[23]  ( .D(Key[23]), .CK(clk), .Q(reg_key[23]) );
  DFF_X1 \reg_key_reg[43]  ( .D(Key[43]), .CK(clk), .Q(reg_key[43]) );
  DFF_X1 \reg_key_reg[169]  ( .D(Key[169]), .CK(clk), .Q(reg_key[169]) );
  DFF_X1 \reg_key_reg[131]  ( .D(Key[131]), .CK(clk), .Q(reg_key[131]) );
  DFF_X1 \reg_key_reg[185]  ( .D(Key[185]), .CK(clk), .Q(reg_key[185]) );
  DFF_X1 \reg_key_reg[36]  ( .D(Key[36]), .CK(clk), .Q(reg_key[36]) );
  DFF_X1 \reg_key_reg[86]  ( .D(Key[86]), .CK(clk), .Q(reg_key[86]) );
  DFF_X1 \reg_key_reg[161]  ( .D(Key[161]), .CK(clk), .Q(reg_key[161]) );
  DFF_X1 \reg_key_reg[71]  ( .D(Key[71]), .CK(clk), .Q(reg_key[71]) );
  DFF_X1 \reg_key_reg[123]  ( .D(Key[123]), .CK(clk), .Q(reg_key[123]) );
  DFF_X1 \reg_key_reg[157]  ( .D(Key[157]), .CK(clk), .Q(reg_key[157]) );
  DFF_X1 \reg_key_reg[170]  ( .D(Key[170]), .CK(clk), .Q(reg_key[170]) );
  DFF_X1 \Ciphertext_reg[44]  ( .D(reg_out[44]), .CK(clk), .Q(Ciphertext[44])
         );
  DFF_X1 \Ciphertext_reg[73]  ( .D(reg_out[73]), .CK(clk), .Q(Ciphertext[73])
         );
  DFF_X1 \reg_key_reg[22]  ( .D(Key[22]), .CK(clk), .Q(reg_key[22]) );
  DFF_X1 \reg_key_reg[186]  ( .D(Key[186]), .CK(clk), .Q(reg_key[186]) );
  DFF_X1 \reg_key_reg[76]  ( .D(Key[76]), .CK(clk), .Q(reg_key[76]) );
  DFF_X1 \reg_key_reg[103]  ( .D(Key[103]), .CK(clk), .Q(reg_key[103]) );
  DFF_X1 \reg_key_reg[48]  ( .D(Key[48]), .CK(clk), .Q(reg_key[48]) );
  DFF_X1 \reg_key_reg[47]  ( .D(Key[47]), .CK(clk), .Q(reg_key[47]) );
  DFF_X1 \reg_key_reg[184]  ( .D(Key[184]), .CK(clk), .Q(reg_key[184]) );
  DFF_X1 \reg_key_reg[156]  ( .D(Key[156]), .CK(clk), .Q(reg_key[156]) );
  DFF_X1 \reg_key_reg[46]  ( .D(Key[46]), .CK(clk), .Q(reg_key[46]) );
  DFF_X1 \reg_key_reg[128]  ( .D(Key[128]), .CK(clk), .Q(reg_key[128]) );
  DFF_X1 \reg_key_reg[73]  ( .D(Key[73]), .CK(clk), .Q(reg_key[73]) );
  DFF_X1 \reg_key_reg[45]  ( .D(Key[45]), .CK(clk), .Q(reg_key[45]) );
  DFF_X1 \reg_key_reg[17]  ( .D(Key[17]), .CK(clk), .Q(reg_key[17]) );
  DFF_X1 \reg_key_reg[154]  ( .D(Key[154]), .CK(clk), .Q(reg_key[154]) );
  DFF_X1 \reg_key_reg[180]  ( .D(Key[180]), .CK(clk), .Q(reg_key[180]) );
  DFF_X1 \reg_key_reg[124]  ( .D(Key[124]), .CK(clk), .Q(reg_key[124]) );
  DFF_X1 \reg_key_reg[96]  ( .D(Key[96]), .CK(clk), .Q(reg_key[96]) );
  DFF_X1 \reg_key_reg[67]  ( .D(Key[67]), .CK(clk), .Q(reg_key[67]) );
  DFF_X1 \reg_key_reg[149]  ( .D(Key[149]), .CK(clk), .Q(reg_key[149]) );
  DFF_X1 \reg_key_reg[39]  ( .D(Key[39]), .CK(clk), .Q(reg_key[39]) );
  DFF_X1 \reg_key_reg[146]  ( .D(Key[146]), .CK(clk), .Q(reg_key[146]) );
  DFF_X1 \reg_key_reg[118]  ( .D(Key[118]), .CK(clk), .Q(reg_key[118]) );
  DFF_X1 \reg_key_reg[63]  ( .D(Key[63]), .CK(clk), .Q(reg_key[63]) );
  DFF_X1 \reg_key_reg[145]  ( .D(Key[145]), .CK(clk), .Q(reg_key[145]) );
  DFF_X1 \reg_key_reg[90]  ( .D(Key[90]), .CK(clk), .Q(reg_key[90]) );
  DFF_X1 \reg_key_reg[117]  ( .D(Key[117]), .CK(clk), .Q(reg_key[117]) );
  DFF_X1 \reg_key_reg[62]  ( .D(Key[62]), .CK(clk), .Q(reg_key[62]) );
  DFF_X1 \reg_key_reg[34]  ( .D(Key[34]), .CK(clk), .Q(reg_key[34]) );
  DFF_X1 \reg_key_reg[143]  ( .D(Key[143]), .CK(clk), .Q(reg_key[143]) );
  DFF_X1 \reg_key_reg[88]  ( .D(Key[88]), .CK(clk), .Q(reg_key[88]) );
  DFF_X1 \reg_key_reg[115]  ( .D(Key[115]), .CK(clk), .Q(reg_key[115]) );
  DFF_X1 \reg_key_reg[5]  ( .D(Key[5]), .CK(clk), .Q(reg_key[5]) );
  DFF_X1 \reg_key_reg[142]  ( .D(Key[142]), .CK(clk), .Q(reg_key[142]) );
  DFF_X1 \reg_key_reg[31]  ( .D(Key[31]), .CK(clk), .Q(reg_key[31]) );
  DFF_X1 \reg_key_reg[113]  ( .D(Key[113]), .CK(clk), .Q(reg_key[113]) );
  DFF_X1 \reg_key_reg[58]  ( .D(Key[58]), .CK(clk), .Q(reg_key[58]) );
  DFF_X1 \reg_key_reg[30]  ( .D(Key[30]), .CK(clk), .Q(reg_key[30]) );
  DFF_X1 \reg_key_reg[29]  ( .D(Key[29]), .CK(clk), .Q(reg_key[29]) );
  DFF_X1 \reg_key_reg[138]  ( .D(Key[138]), .CK(clk), .Q(reg_key[138]) );
  DFF_X1 \reg_key_reg[110]  ( .D(Key[110]), .CK(clk), .Q(reg_key[110]) );
  DFF_X1 \reg_key_reg[55]  ( .D(Key[55]), .CK(clk), .Q(reg_key[55]) );
  DFF_X1 \reg_key_reg[164]  ( .D(Key[164]), .CK(clk), .Q(reg_key[164]) );
  DFF_X1 \reg_key_reg[109]  ( .D(Key[109]), .CK(clk), .Q(reg_key[109]) );
  DFF_X1 \reg_key_reg[136]  ( .D(Key[136]), .CK(clk), .Q(reg_key[136]) );
  DFF_X1 \reg_key_reg[81]  ( .D(Key[81]), .CK(clk), .Q(reg_key[81]) );
  DFF_X1 \reg_key_reg[163]  ( .D(Key[163]), .CK(clk), .Q(reg_key[163]) );
  DFF_X1 \reg_key_reg[162]  ( .D(Key[162]), .CK(clk), .Q(reg_key[162]) );
  DFF_X1 \reg_key_reg[106]  ( .D(Key[106]), .CK(clk), .Q(reg_key[106]) );
  DFF_X1 \reg_key_reg[133]  ( .D(Key[133]), .CK(clk), .Q(reg_key[133]) );
  DFF_X1 \reg_key_reg[105]  ( .D(Key[105]), .CK(clk), .Q(reg_key[105]) );
  DFF_X1 \reg_key_reg[165]  ( .D(Key[165]), .CK(clk), .Q(reg_key[165]) );
  DFF_X1 \reg_key_reg[97]  ( .D(Key[97]), .CK(clk), .Q(reg_key[97]) );
  DFF_X1 \reg_key_reg[158]  ( .D(Key[158]), .CK(clk), .Q(reg_key[158]) );
  DFF_X1 \reg_key_reg[102]  ( .D(Key[102]), .CK(clk), .Q(reg_key[102]) );
  DFF_X1 \reg_key_reg[18]  ( .D(Key[18]), .CK(clk), .Q(reg_key[18]) );
  DFF_X1 \reg_key_reg[182]  ( .D(Key[182]), .CK(clk), .Q(reg_key[182]) );
  DFF_X1 \reg_key_reg[72]  ( .D(Key[72]), .CK(clk), .Q(reg_key[72]) );
  DFF_X1 \reg_key_reg[99]  ( .D(Key[99]), .CK(clk), .Q(reg_key[99]) );
  DFF_X1 \reg_key_reg[181]  ( .D(Key[181]), .CK(clk), .Q(reg_key[181]) );
  DFF_X1 \reg_key_reg[42]  ( .D(Key[42]), .CK(clk), .Q(reg_key[42]) );
  DFF_X1 \reg_key_reg[14]  ( .D(Key[14]), .CK(clk), .Q(reg_key[14]) );
  DFF_X1 \reg_key_reg[12]  ( .D(Key[12]), .CK(clk), .Q(reg_key[12]) );
  DFF_X1 \reg_key_reg[38]  ( .D(Key[38]), .CK(clk), .Q(reg_key[38]) );
  DFF_X1 \reg_key_reg[120]  ( .D(Key[120]), .CK(clk), .Q(reg_key[120]) );
  DFF_X1 \reg_key_reg[10]  ( .D(Key[10]), .CK(clk), .Q(reg_key[10]) );
  DFF_X1 \reg_key_reg[89]  ( .D(Key[89]), .CK(clk), .Q(reg_key[89]) );
  DFF_X1 \reg_key_reg[59]  ( .D(Key[59]), .CK(clk), .Q(reg_key[59]) );
  DFF_X1 \reg_key_reg[85]  ( .D(Key[85]), .CK(clk), .Q(reg_key[85]) );
  DFF_X1 \reg_key_reg[139]  ( .D(Key[139]), .CK(clk), .Q(reg_key[139]) );
  DFF_X1 \reg_key_reg[52]  ( .D(Key[52]), .CK(clk), .Q(reg_key[52]) );
  DFF_X1 \reg_key_reg[132]  ( .D(Key[132]), .CK(clk), .Q(reg_key[132]) );
  DFF_X1 \reg_key_reg[126]  ( .D(Key[126]), .CK(clk), .Q(reg_key[126]) );
  DFF_X1 \reg_key_reg[75]  ( .D(Key[75]), .CK(clk), .Q(reg_key[75]) );
  DFF_X1 \reg_key_reg[127]  ( .D(Key[127]), .CK(clk), .Q(reg_key[127]) );
  DFF_X1 \reg_key_reg[69]  ( .D(Key[69]), .CK(clk), .Q(reg_key[69]) );
  DFF_X1 \reg_key_reg[114]  ( .D(Key[114]), .CK(clk), .Q(reg_key[114]) );
  DFF_X1 \reg_key_reg[141]  ( .D(Key[141]), .CK(clk), .Q(reg_key[141]) );
  DFF_X1 \reg_key_reg[188]  ( .D(Key[188]), .CK(clk), .Q(reg_key[188]) );
  DFF_X1 \reg_key_reg[60]  ( .D(Key[60]), .CK(clk), .Q(reg_key[60]) );
  DFF_X1 \reg_key_reg[6]  ( .D(Key[6]), .CK(clk), .Q(reg_key[6]) );
  DFF_X1 \reg_key_reg[4]  ( .D(Key[4]), .CK(clk), .Q(reg_key[4]) );
  DFF_X1 \reg_key_reg[15]  ( .D(Key[15]), .CK(clk), .Q(reg_key[15]) );
  DFF_X1 \reg_key_reg[24]  ( .D(Key[24]), .CK(clk), .Q(reg_key[24]) );
  DFF_X1 \reg_key_reg[65]  ( .D(Key[65]), .CK(clk), .Q(reg_key[65]) );
  DFF_X1 \reg_key_reg[16]  ( .D(Key[16]), .CK(clk), .Q(reg_key[16]) );
  DFF_X1 \reg_key_reg[0]  ( .D(Key[0]), .CK(clk), .Q(reg_key[0]) );
  DFF_X1 \reg_key_reg[13]  ( .D(Key[13]), .CK(clk), .Q(reg_key[13]) );
  DFF_X1 \reg_key_reg[37]  ( .D(Key[37]), .CK(clk), .Q(reg_key[37]) );
  DFF_X1 \reg_key_reg[93]  ( .D(Key[93]), .CK(clk), .Q(reg_key[93]) );
  DFF_X1 \reg_key_reg[94]  ( .D(Key[94]), .CK(clk), .Q(reg_key[94]) );
  DFF_X1 \reg_key_reg[21]  ( .D(Key[21]), .CK(clk), .Q(reg_key[21]) );
  DFF_X1 \reg_key_reg[7]  ( .D(Key[7]), .CK(clk), .Q(reg_key[7]) );
  DFF_X1 \reg_key_reg[95]  ( .D(Key[95]), .CK(clk), .Q(reg_key[95]) );
  DFF_X1 \reg_key_reg[61]  ( .D(Key[61]), .CK(clk), .Q(reg_key[61]) );
  DFF_X1 \reg_key_reg[121]  ( .D(Key[121]), .CK(clk), .Q(reg_key[121]) );
  DFF_X1 \reg_key_reg[64]  ( .D(Key[64]), .CK(clk), .Q(reg_key[64]) );
  DFF_X1 \reg_key_reg[166]  ( .D(Key[166]), .CK(clk), .Q(reg_key[166]) );
  DFF_X1 \reg_key_reg[84]  ( .D(Key[84]), .CK(clk), .Q(reg_key[84]) );
  DFF_X1 \reg_key_reg[54]  ( .D(Key[54]), .CK(clk), .Q(reg_key[54]) );
  DFF_X1 \reg_key_reg[160]  ( .D(Key[160]), .CK(clk), .Q(reg_key[160]) );
  DFF_X1 \reg_key_reg[25]  ( .D(Key[25]), .CK(clk), .Q(reg_key[25]) );
  DFF_X1 \reg_key_reg[78]  ( .D(Key[78]), .CK(clk), .Q(reg_key[78]) );
  DFF_X2 \Ciphertext_reg[105]  ( .D(reg_out[105]), .CK(clk), .Q(
        Ciphertext[105]) );
  DFF_X1 \Ciphertext_reg[102]  ( .D(reg_out[102]), .CK(clk), .Q(
        Ciphertext[102]) );
  DFF_X2 \Ciphertext_reg[28]  ( .D(reg_out[28]), .CK(clk), .Q(Ciphertext[28])
         );
  DFF_X1 \reg_key_reg[144]  ( .D(Key[144]), .CK(clk), .Q(reg_key[144]) );
  DFF_X1 \reg_key_reg[172]  ( .D(Key[172]), .CK(clk), .Q(reg_key[172]) );
  DFFRS_X1 \Ciphertext_reg[50]  ( .D(reg_out[50]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Ciphertext[50]) );
  DFF_X1 \Ciphertext_reg[168]  ( .D(reg_out[168]), .CK(clk), .Q(
        Ciphertext[168]) );
  DFF_X1 \Ciphertext_reg[140]  ( .D(reg_out[140]), .CK(clk), .Q(
        Ciphertext[140]) );
  DFF_X1 \reg_key_reg[100]  ( .D(Key[100]), .CK(clk), .Q(reg_key[100]) );
  SPEEDY_Rounds7_0 SPEEDY_instance ( .Plaintext(reg_in), .Key(reg_key), 
        .Ciphertext(reg_out) );
  DFF_X2 \Ciphertext_reg[111]  ( .D(reg_out[111]), .CK(clk), .Q(
        Ciphertext[111]) );
  DFF_X2 \Ciphertext_reg[108]  ( .D(reg_out[108]), .CK(clk), .Q(
        Ciphertext[108]) );
  DFFRS_X1 \Ciphertext_reg[121]  ( .D(reg_out[121]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Ciphertext[121]) );
  DFF_X2 \Ciphertext_reg[84]  ( .D(reg_out[84]), .CK(clk), .Q(Ciphertext[84])
         );
  DFF_X2 \Ciphertext_reg[188]  ( .D(reg_out[188]), .CK(clk), .Q(
        Ciphertext[188]) );
  DFF_X1 \Ciphertext_reg[0]  ( .D(reg_out[0]), .CK(clk), .Q(Ciphertext[0]) );
  DFF_X1 \Ciphertext_reg[148]  ( .D(reg_out[148]), .CK(clk), .Q(
        Ciphertext[148]) );
endmodule

