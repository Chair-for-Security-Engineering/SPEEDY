
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_SPEEDY_Top is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_SPEEDY_Top;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Rounds5_0 is

   port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : out
         std_logic_vector (191 downto 0));

end SPEEDY_Rounds5_0;

architecture SYN_Behavioral of SPEEDY_Rounds5_0 is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n7, n8, n9, n11, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n40, n41, n44, n45, n46, n48, n49, n50, n52, n53, n55, n57, n60, 
      n61, n63, n64, n65, n66, n67, n68, n70, n71, n73, n74, n75, n76, n78, n79
      , n80, n81, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n95, 
      n98, n99, n100, n102, n103, n104, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n117, n118, n119, n121, n122, n123, n125, n126, n128, 
      n129, n130, n131, n132, n133, n134, n135, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n160, n163, n164, n169, n170, n176, n177, n178, n179, n180, n182, n190, 
      n191, n192, n193, n195, n196, n197, n198, n199, n200, n201, n202, n204, 
      n205, n207, n208, n209, n210, n212, n213, n214, n215, n216, n219, n220, 
      n221, n222, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n273, n274, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n298, n299, n300, n301, n302, n303, n304, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n328, n329, n331, n332, n333, n334, n335, n336, n338, 
      n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
      n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
      n363, n364, n365, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n382, n383, n385, n386, n387, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n409, n410, n411, n412, n415, n416, n417, n419, n420, n421, 
      n422, n423, n424, n425, n427, n428, n429, n430, n431, n432, n434, n435, 
      n436, n437, n439, n440, n443, n444, n445, n446, n447, n448, n449, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n469, n470, n471, n472, n473, n474, n475, n477, 
      n478, n479, n480, n481, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n499, n502, n504, n505, n506, n507, 
      n508, n509, n510, n512, n513, n515, n516, n517, n518, n519, n520, n521, 
      n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, 
      n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, 
      n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, 
      n558, n559, n560, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n581, n582, n583, 
      n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, 
      n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, 
      n609, n610, n611, n612, n613, n614, n615, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n637, n638, n639, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n654, n655, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n667, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
      n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, 
      n786, n787, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n841, n842, n843, n844, n845, n846, n847, n848, 
      n850, n851, n852, n854, n855, n856, n857, n859, n860, n861, n862, n864, 
      n865, n868, n870, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n888, n889, n890, n891, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
      n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n933, 
      n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n946, n947, 
      n948, n951, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, 
      n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, 
      n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, 
      n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
      n1072, n1073, n1074, n1075, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1122, n1123, 
      n1124, n1126, n1127, n1128, n1129, n1131, n1132, n1133, n1136, n1137, 
      n1139, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, 
      n1162, n1163, n1164, n1165, n1166, n1167, n1170, n1173, n1174, n1175, 
      n1176, n1177, n1178, n1179, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1192, n1193, n1194, n1195, n1196, n1197, 
      n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
      n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
      n1218, n1219, n1220, n1221, n1223, n1224, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1270, n1271, 
      n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, 
      n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, 
      n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
      n1302, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, 
      n1324, n1325, n1326, n1327, n1329, n1330, n1331, n1332, n1333, n1334, 
      n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1343, n1344, n1345, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1356, n1357, 
      n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, 
      n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1376, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, 
      n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
      n1431, n1432, n1433, n1435, n1436, n1437, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1452, n1453, 
      n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, 
      n1464, n1465, n1466, n1468, n1469, n1470, n1471, n1472, n1473, n1474, 
      n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1546, n1547, 
      n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
      n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, 
      n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, 
      n1578, n1579, n1580, n1581, n1584, n1585, n1586, n1587, n1588, n1589, 
      n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
      n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
      n1610, n1611, n1613, n1614, n1615, n1616, n1618, n1619, n1620, n1621, 
      n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, 
      n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, 
      n1642, n1643, n1644, n1645, n1646, n1647, n1649, n1650, n1651, n1652, 
      n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, 
      n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, 
      n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
      n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
      n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1710, n1711, n1712, n1714, n1715, n1716, n1717, 
      n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, 
      n1728, n1729, n1730, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1761, n1762, n1763, n1764, n1765, n1766, n1768, n1769, n1770, 
      n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, 
      n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, 
      n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
      n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
      n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, 
      n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, 
      n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, 
      n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, 
      n1885, n1886, n1887, n1888, n1890, n1891, n1892, n1893, n1894, n1895, 
      n1896, n1897, n1898, n1899, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1914, n1915, n1916, n1917, 
      n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n1950, n1951, n1952, n1954, n1955, n1956, n1957, n1958, n1959, n1960, 
      n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
      n1971, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, 
      n1982, n1983, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, 
      n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, 
      n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, 
      n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, 
      n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, 
      n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2065, 
      n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
      n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2108, 
      n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2118, n2120, 
      n2121, n2122, n2123, n2125, n2126, n2127, n2129, n2130, n2132, n2133, 
      n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, 
      n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, 
      n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, 
      n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, 
      n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, 
      n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, 
      n2195, n2196, n2197, n2199, n2200, n2201, n2202, n2203, n2204, n2205, 
      n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, 
      n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, 
      n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, 
      n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2246, n2247, 
      n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, 
      n2289, n2290, n2291, n2292, n2293, n2294, n2296, n2297, n2298, n2299, 
      n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, 
      n2310, n2311, n2312, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
      n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2372, n2373, 
      n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, 
      n2384, n2385, n2386, n2387, n2389, n2390, n2391, n2392, n2393, n2394, 
      n2395, n2396, n2397, n2399, n2400, n2401, n2402, n2403, n2404, n2405, 
      n2406, n2407, n2408, n2410, n2411, n2412, n2413, n2414, n2415, n2417, 
      n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
      n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2437, n2438, 
      n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2448, n2449, 
      n2450, n2451, n2452, n2454, n2455, n2456, n2457, n2458, n2460, n2461, 
      n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, 
      n2472, n2473, n2474, n2475, n2476, n2478, n2479, n2480, n2481, n2482, 
      n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
      n2493, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, 
      n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, 
      n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
      n2524, n2525, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2535, n2536, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, 
      n2546, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2570, n2571, n2572, n2573, n2576, n2577, n2578, n2579, 
      n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2590, n2591, 
      n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2600, n2601, n2602, 
      n2603, n2604, n2605, n2606, n2607, n2608, n2610, n2611, n2612, n2613, 
      n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
      n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
      n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, 
      n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, 
      n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2664, 
      n2665, n2666, n2668, n2669, n2670, n2671, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2684, n2685, n2686, n2687, 
      n2688, n2689, n2690, n2691, n2692, n2693, n2695, n2696, n2697, n2698, 
      n2699, n2701, n2702, n2703, n2704, n2705, n2707, n2709, n2711, n2712, 
      n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
      n2723, n2724, n2725, n2726, n2727, n2729, n2730, n2731, n2732, n2733, 
      n2734, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, 
      n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, 
      n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, 
      n2766, n2767, n2768, n2769, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2781, n2782, n2783, n2784, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2828, n2829, n2830, 
      n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, 
      n2842, n2843, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, 
      n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
      n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
      n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
      n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
      n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
      n2905, n2906, n2907, n2908, n2910, n2911, n2912, n2913, n2914, n2915, 
      n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
      n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, 
      n2936, n2937, n2938, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2964, n2965, n2966, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, 
      n2979, n2980, n2981, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
      n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
      n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, 
      n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
      n3020, n3021, n3022, n3023, n3024, n3025, n3027, n3028, n3030, n3031, 
      n3034, n3035, n3036, n3038, n3039, n3040, n3041, n3042, n3043, n3044, 
      n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, 
      n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3064, n3065, 
      n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, 
      n3076, n3078, n3079, n3080, n3081, n3082, n3085, n3086, n3087, n3088, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
      n3099, n3100, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, 
      n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, 
      n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, 
      n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, 
      n3141, n3142, n3143, n3146, n3147, n3148, n3149, n3150, n3151, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3164, 
      n3165, n3166, n3167, n3168, n3169, n3171, n3172, n3173, n3174, n3175, 
      n3176, n3177, n3178, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3203, n3204, n3205, n3206, n3207, 
      n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3234, n3235, n3236, n3237, n3238, n3239, 
      n3240, n3241, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, 
      n3251, n3252, n3253, n3254, n3256, n3257, n3258, n3259, n3260, n3261, 
      n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, 
      n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
      n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, 
      n3293, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
      n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
      n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, 
      n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, 
      n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3343, n3344, 
      n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, 
      n3355, n3356, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, 
      n3366, n3367, n3368, n3369, n3370, n3371, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3436, n3437, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3453, n3454, n3455, n3456, n3457, n3458, n3459, 
      n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, 
      n3470, n3471, n3472, n3473, n3475, n3476, n3477, n3478, n3479, n3480, 
      n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, 
      n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, 
      n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, 
      n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, 
      n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, 
      n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, 
      n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, 
      n3552, n3553, n3554, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3572, n3573, 
      n3574, n3575, n3576, n3578, n3579, n3580, n3581, n3583, n3584, n3585, 
      n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, 
      n3596, n3597, n3598, n3599, n3601, n3602, n3603, n3604, n3605, n3606, 
      n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, 
      n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, 
      n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, 
      n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, 
      n3647, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, 
      n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, 
      n3669, n3670, n3671, n3672, n3674, n3675, n3676, n3677, n3678, n3679, 
      n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, 
      n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, 
      n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3709, n3710, 
      n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, 
      n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, 
      n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, 
      n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, 
      n3752, n3753, n3754, n3755, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3774, 
      n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, 
      n3785, n3787, n3788, n3789, n3791, n3793, n3794, n3795, n3796, n3797, 
      n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, 
      n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, 
      n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, 
      n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3838, 
      n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, 
      n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, 
      n3859, n3860, n3861, n3862, n3864, n3865, n3866, n3867, n3868, n3869, 
      n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, 
      n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, 
      n3890, n3891, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, 
      n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, 
      n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, 
      n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, 
      n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3941, 
      n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, 
      n3952, n3953, n3954, n3955, n3956, n3957, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3986, n3987, n3988, n3989, n3991, n3992, n3993, n3994, 
      n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, 
      n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, 
      n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, 
      n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, 
      n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, 
      n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, 
      n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, 
      n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, 
      n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, 
      n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, 
      n4095, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, 
      n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, 
      n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, 
      n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, 
      n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4146, 
      n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, 
      n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, 
      n4167, n4168, n4169, n4170, n4171, n4172, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4206, n4207, n4208, 
      n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
      n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, 
      n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, 
      n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, 
      n4250, n4251, n4253, n4254, n4255, n4256, n4257, n4259, n4260, n4261, 
      n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, 
      n4272, n4273, n4274, n4275, n4276, n4277, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4290, n4291, n4292, n4293, 
      n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
      n4304, n4305, n4306, n4307, n4308, n4309, n4311, n4312, n4313, n4314, 
      n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, 
      n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, 
      n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, 
      n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, 
      n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, 
      n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, 
      n4376, n4377, n4378, n4379, n4380, n4381, n4383, n4384, n4385, n4386, 
      n4387, n4388, n4389, n4390, n4391, n4392, n4395, n4396, n4397, n4398, 
      n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, 
      n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, 
      n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4428, n4430, 
      n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, 
      n4441, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, 
      n4452, n4453, n4454, n4455, n4456, n4457, n4459, n4460, n4461, n4462, 
      n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
      n4473, n4474, n4475, n4476, n4477, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4527, n4528, n4529, n4532, n4533, n4534, n4535, n4536, 
      n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, 
      n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, 
      n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, 
      n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, 
      n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, 
      n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, 
      n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, 
      n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, 
      n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, 
      n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, 
      n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, 
      n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, 
      n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, 
      n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, 
      n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, 
      n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, 
      n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, 
      n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, 
      n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, 
      n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, 
      n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, 
      n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, 
      n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, 
      n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, 
      n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, 
      n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, 
      n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, 
      n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, 
      n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, 
      n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, 
      n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, 
      n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, 
      n4857, n4858, n4859, n4860, n4862, n4863, n4864, n4865, n4866, n4867, 
      n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, 
      n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, 
      n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4896, n4897, n4898, 
      n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, 
      n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, 
      n4919, n4920, n4921, n4922, n4923, n4924, n4926, n4927, n4928, n4929, 
      n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, 
      n4940, n4941, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, 
      n4951, n4952, n4953, n4954, n4955, n4958, n4959, n4960, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, 
      n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
      n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, 
      n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5083, n5085, 
      n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, 
      n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, 
      n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, 
      n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, 
      n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, 
      n5136, n5137, n5138, n5139, n5141, n5142, n5143, n5144, n5145, n5146, 
      n5147, n5148, n5150, n5151, n5152, n5153, n5155, n5156, n5157, n5158, 
      n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, 
      n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, 
      n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, 
      n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, 
      n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, 
      n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, 
      n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, 
      n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, 
      n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5249, 
      n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, 
      n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, 
      n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, 
      n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, 
      n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, 
      n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, 
      n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, 
      n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, 
      n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, 
      n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, 
      n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, 
      n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, 
      n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, 
      n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, 
      n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, 
      n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, 
      n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, 
      n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, 
      n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, 
      n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, 
      n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, 
      n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, 
      n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, 
      n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, 
      n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, 
      n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, 
      n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, 
      n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, 
      n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, 
      n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, 
      n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, 
      n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, 
      n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, 
      n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, 
      n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, 
      n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, 
      n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, 
      n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, 
      n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, 
      n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, 
      n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, 
      n5662, n5663, n5664, n5665, n5666, n5668, n5669, n5670, n5671, n5672, 
      n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, 
      n5693, n5694, n5695, n5697, n5698, n5699, n5700, n5701, n5702, n5703, 
      n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, 
      n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, 
      n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, 
      n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, 
      n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, 
      n5754, n5756, n5757, n5758, n5759, n5760, n5762, n5763, n5764, n5765, 
      n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, 
      n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, 
      n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, 
      n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, 
      n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, 
      n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, 
      n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5837, 
      n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, 
      n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, 
      n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, 
      n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, 
      n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, 
      n5888, n5889, n5890, n5891, n5893, n5895, n5896, n5897, n5898, n5899, 
      n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, 
      n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, 
      n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, 
      n5930, n5931, n5932, n5934, n5935, n5936, n5937, n5938, n5939, n5940, 
      n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, 
      n5951, n5952, n5953, n5955, n5956, n5957, n5958, n5959, n5960, n5961, 
      n5962, n5963, n5965, n5967, n5968, n5969, n5970, n5971, n5972, n5973, 
      n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, 
      n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6010, n6011, n6012, n6013, n6014, n6015, 
      n6016, n6017, n6018, n6020, n6021, n6022, n6023, n6024, n6025, n6026, 
      n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, 
      n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, 
      n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, 
      n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, 
      n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, 
      n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, 
      n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, 
      n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, 
      n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, 
      n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, 
      n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, 
      n6137, n6138, n6139, n6140, n6141, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
      n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, 
      n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, 
      n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, 
      n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, 
      n6198, n6199, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, 
      n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, 
      n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, 
      n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, 
      n6240, n6241, n6242, n6243, n6244, n6246, n6247, n6248, n6249, n6250, 
      n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, 
      n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, 
      n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, 
      n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, 
      n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, 
      n6301, n6302, n6303, n6304, n6305, n6307, n6308, n6309, n6310, n6311, 
      n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, 
      n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, 
      n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
      n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, 
      n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, 
      n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
      n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
      n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, 
      n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, 
      n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, 
      n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
      n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, 
      n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, 
      n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, 
      n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, 
      n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, 
      n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, 
      n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, 
      n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, 
      n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, 
      n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, 
      n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, 
      n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, 
      n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, 
      n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, 
      n6562, n6563, n6564, n6565, n6566, n6567, n6569, n6570, n6571, n6572, 
      n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, 
      n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, 
      n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, 
      n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, 
      n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, 
      n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, 
      n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, 
      n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, 
      n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, 
      n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, 
      n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, 
      n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, 
      n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, 
      n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6792, n6793, n6794, 
      n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, 
      n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, 
      n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, 
      n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, 
      n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, 
      n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, 
      n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, 
      n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
      n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
      n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, 
      n6896, n6897, n6898, n6900, n6901, n6902, n6903, n6904, n6905, n6906, 
      n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, 
      n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, 
      n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, 
      n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, 
      n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, 
      n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, 
      n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, 
      n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, 
      n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, 
      n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, 
      n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, 
      n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, 
      n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, 
      n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, 
      n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7057, 
      n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, 
      n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, 
      n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, 
      n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, 
      n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, 
      n7108, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, 
      n7119, n7121, n7122, n7123, n7125, n7126, n7127, n7128, n7129, n7130, 
      n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, 
      n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, 
      n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, 
      n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, 
      n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, 
      n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, 
      n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, 
      n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, 
      n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, 
      n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, 
      n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, 
      n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, 
      n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, 
      n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, 
      n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, 
      n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, 
      n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, 
      n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, 
      n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, 
      n7321, n7322, n7323, n7324, n7325, n7326, n7328, n7329, n7330, n7331, 
      n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, 
      n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, 
      n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, 
      n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, 
      n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, 
      n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, 
      n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, 
      n7402, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, 
      n7413, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7440, n7441, n7442, n7443, n7444, 
      n7445, n7446, n7447, n7448, n7449, n7452, n7453, n7454, n7455, n7456, 
      n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, 
      n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, 
      n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, 
      n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, 
      n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, 
      n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, 
      n7517, n7519, n7520, n7521, n7523, n7524, n7525, n7526, n7527, n7528, 
      n7529, n7530, n7531, n7533, n7534, n7535, n7536, n7537, n7538, n7539, 
      n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, 
      n7551, n7552, n7553, n7554, n7555, n7556, n7558, n7559, n7560, n7561, 
      n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, 
      n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, 
      n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7590, n7591, n7592, 
      n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, 
      n7603, n7604, n7605, n7606, n7607, n7608, n7610, n7611, n7612, n7613, 
      n7615, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, 
      n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7636, 
      n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, 
      n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, 
      n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, 
      n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, 
      n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, 
      n7687, n7688, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, 
      n7698, n7701, n7702, n7703, n7704, n7705, n7706, n7708, n7709, n7710, 
      n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, 
      n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, 
      n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, 
      n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, 
      n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, 
      n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, 
      n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, 
      n7781, n7782, n7783, n7784, n7786, n7787, n7788, n7789, n7790, n7791, 
      n7792, n7793, n7794, n7795, n7796, n7797, n7799, n7800, n7801, n7802, 
      n7803, n7804, n7805, n7806, n7807, n7808, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, 
      n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, 
      n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, 
      n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, 
      n7855, n7856, n7857, n7858, n7859, n7861, n7862, n7863, n7864, n7865, 
      n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, 
      n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, 
      n7886, n7887, n7888, n7889, n7890, n7892, n7893, n7894, n7895, n7896, 
      n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7908, 
      n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, 
      n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, 
      n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7938, n7939, 
      n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, 
      n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, 
      n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, 
      n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, 
      n7980, n7981, n7982, n7984, n7985, n7986, n7987, n7988, n7989, n7990, 
      n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n8000, n8001, 
      n8002, n8003, n8004, n8006, n8007, n8008, n8009, n8010, n8011, n8012, 
      n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8059, n8060, n8061, n8062, n8063, n8064, 
      n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, 
      n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, 
      n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8093, n8094, n8095, 
      n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, 
      n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8116, 
      n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, 
      n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, 
      n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, 
      n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, 
      n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, 
      n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, 
      n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, 
      n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, 
      n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, 
      n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, 
      n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, 
      n8227, n8228, n8230, n8232, n8234, n8235, n8236, n8237, n8238, n8239, 
      n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, 
      n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, 
      n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8268, n8269, n8270, 
      n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, 
      n8281, n8282, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, 
      n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, 
      n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8312, n8313, n8314, 
      n8315, n8316, n8317, n8318, n8319, n8320, n8322, n8323, n8324, n8325, 
      n8326, n8327, n8328, n8330, n8331, n8332, n8333, n8334, n8335, n8336, 
      n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, 
      n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, 
      n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, 
      n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8375, n8376, n8377, 
      n8378, n8379, n8380, n8381, n8382, n8384, n8385, n8386, n8387, n8388, 
      n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, 
      n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, 
      n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, 
      n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, 
      n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, 
      n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, 
      n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, 
      n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, 
      n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, 
      n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8489, 
      n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, 
      n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, 
      n8510, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, 
      n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, 
      n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, 
      n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8550, n8551, n8552, 
      n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, 
      n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, 
      n8573, n8574, n8575, n8577, n8578, n8579, n8580, n8581, n8583, n8584, 
      n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, 
      n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, 
      n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, 
      n8615, n8616, n8617, n8618, n8619, n8622, n8623, n8624, n8625, n8626, 
      n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8638, 
      n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, 
      n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, 
      n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8668, n8669, 
      n8670, n8671, n8672, n8673, n8674, n8676, n8677, n8678, n8679, n8680, 
      n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, 
      n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, 
      n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8710, n8711, n8712, 
      n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, 
      n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, 
      n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, 
      n8743, n8744, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8754, 
      n8755, n8756, n8757, n8759, n8760, n8761, n8762, n8763, n8764, n8765, 
      n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, 
      n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, 
      n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, 
      n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, 
      n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, 
      n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, 
      n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, 
      n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, 
      n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, 
      n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, 
      n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, 
      n8876, n8877, n8878, n8879, n8881, n8882, n8883, n8884, n8885, n8886, 
      n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, 
      n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, 
      n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, 
      n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, 
      n8927, n8928, n8929, n8931, n8932, n8933, n8934, n8935, n8936, n8937, 
      n8939, n8940, n8941, n8942, n8944, n8945, n8946, n8947, n8948, n8949, 
      n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, 
      n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, 
      n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8979, n8980, 
      n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, 
      n8991, n8993, n8994, n8995, n8997, n8998, n8999, n9000, n9001, n9002, 
      n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, 
      n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, 
      n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, 
      n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, 
      n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, 
      n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, 
      n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, 
      n9073, n9074, n9075, n9076, n9078, n9079, n9080, n9081, n9082, n9083, 
      n9084, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, 
      n9096, n9097, n9098, n9099, n9100, n9103, n9104, n9105, n9106, n9107, 
      n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, 
      n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, 
      n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, 
      n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9147, n9148, 
      n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, 
      n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, 
      n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, 
      n9179, n9180, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, 
      n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, 
      n9200, n9201, n9202, n9204, n9206, n9207, n9208, n9209, n9210, n9211, 
      n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, 
      n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, 
      n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, 
      n9242, n9243, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, 
      n9253, n9255, n9256, n9257, n9258, n9260, n9261, n9262, n9264, n9265, 
      n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, 
      n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, 
      n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, 
      n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, 
      n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, 
      n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, 
      n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, 
      n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, 
      n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, 
      n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, 
      n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, 
      n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, 
      n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, 
      n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, 
      n9406, n9407, n9408, n9409, n9410, n9411, n9413, n9414, n9415, n9416, 
      n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, 
      n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, 
      n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, 
      n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, 
      n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, 
      n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, 
      n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, 
      n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, 
      n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, 
      n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, 
      n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, 
      n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, 
      n9537, n9538, n9539, n9540, n9541, n9543, n9544, n9545, n9546, n9547, 
      n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, 
      n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9566, n9567, n9568, 
      n9569, n9570, n9571, n9572, n9573, n9575, n9576, n9577, n9578, n9579, 
      n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, 
      n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, 
      n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, 
      n9610, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, 
      n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, 
      n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, 
      n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, 
      n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, 
      n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, 
      n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, 
      n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, 
      n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, 
      n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, 
      n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, 
      n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, 
      n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, 
      n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, 
      n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9760, n9761, 
      n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, 
      n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, 
      n9782, n9783, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, 
      n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, 
      n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, 
      n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, 
      n9824, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9834, n9836, 
      n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, 
      n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, 
      n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9867, n9868, 
      n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, 
      n9879, n9880, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9891, 
      n9892, n9893, n9894, n9895, n9898, n9899, n9900, n9901, n9902, n9904, 
      n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, 
      n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, 
      n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, 
      n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, 
      n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, 
      n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, 
      n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, 
      n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, 
      n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, 
      n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004
      , n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
      n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, 
      n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, 
      n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, 
      n10042, n10043, n10044, n10046, n10047, n10048, n10049, n10050, n10051, 
      n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, 
      n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, 
      n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, 
      n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, 
      n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, 
      n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, 
      n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, 
      n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, 
      n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, 
      n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, 
      n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, 
      n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, 
      n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, 
      n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, 
      n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, 
      n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, 
      n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, 
      n10205, n10206, n10207, n10208, n10209, n10210, n10213, n10214, n10215, 
      n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, 
      n10225, n10226, n10227, n10229, n10230, n10231, n10232, n10233, n10234, 
      n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, 
      n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, 
      n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, 
      n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, 
      n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, 
      n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, 
      n10289, n10290, n10291, n10292, n10293, n10295, n10296, n10297, n10298, 
      n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, 
      n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, 
      n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, 
      n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, 
      n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, 
      n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, 
      n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, 
      n10362, n10363, n10364, n10365, n10366, n10367, n10369, n10370, n10371, 
      n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, 
      n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, 
      n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, 
      n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, 
      n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, 
      n10417, n10418, n10419, n10420, n10421, n10422, n10424, n10425, n10426, 
      n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, 
      n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, 
      n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, 
      n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, 
      n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, 
      n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, 
      n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, 
      n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, 
      n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, 
      n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, 
      n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, 
      n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, 
      n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, 
      n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, 
      n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, 
      n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, 
      n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, 
      n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, 
      n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, 
      n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, 
      n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10615, n10616, 
      n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10625, n10626, 
      n10627, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, 
      n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, 
      n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, 
      n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, 
      n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, 
      n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, 
      n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, 
      n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, 
      n10701, n10702, n10703, n10704, n10705, n10707, n10708, n10709, n10710, 
      n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, 
      n10720, n10721, n10722, n10724, n10725, n10726, n10727, n10728, n10729, 
      n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, 
      n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, 
      n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, 
      n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, 
      n10766, n10767, n10768, n10769, n10770, n10772, n10773, n10774, n10775, 
      n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, 
      n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, 
      n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, 
      n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, 
      n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, 
      n10821, n10822, n10824, n10825, n10826, n10827, n10828, n10829, n10830, 
      n10831, n10832, n10833, n10835, n10836, n10837, n10838, n10839, n10840, 
      n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, 
      n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, 
      n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, 
      n10868, n10869, n10870, n10871, n10873, n10874, n10875, n10876, n10877, 
      n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, 
      n10887, n10888, n10889, n10890, n10892, n10893, n10894, n10895, n10896, 
      n10897, n10898, n10899, n10900, n10901, n10903, n10904, n10905, n10906, 
      n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, 
      n10916, n10917, n10918, n10919, n10921, n10922, n10923, n10924, n10925, 
      n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, 
      n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10944, 
      n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, 
      n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, 
      n10964, n10965, n10966, n10967, n10968, n10970, n10971, n10972, n10973, 
      n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, 
      n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, 
      n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, 
      n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, 
      n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, 
      n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, 
      n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, 
      n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, 
      n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, 
      n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, 
      n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, 
      n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, 
      n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, 
      n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, 
      n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11109, 
      n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11119, 
      n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, 
      n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, 
      n11138, n11139, n11140, n11142, n11143, n11144, n11145, n11146, n11147, 
      n11148, n11149, n11151, n11152, n11153, n11154, n11155, n11156, n11157, 
      n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, 
      n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, 
      n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, 
      n11185, n11186, n11187, n11188, n11189, n11191, n11192, n11193, n11194, 
      n11195, n11196, n11198, n11199, n11200, n11201, n11202, n11203, n11204, 
      n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, 
      n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, 
      n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, 
      n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, 
      n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, 
      n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, 
      n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, 
      n11268, n11269, n11270, n11271, n11274, n11275, n11276, n11277, n11278, 
      n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, 
      n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, 
      n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, 
      n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, 
      n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, 
      n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, 
      n11334, n11335, n11336, n11337, n11339, n11340, n11341, n11342, n11343, 
      n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, 
      n11353, n11354, n11355, n11356, n11358, n11359, n11360, n11361, n11362, 
      n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, 
      n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, 
      n11381, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, 
      n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, 
      n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, 
      n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, 
      n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11427, n11428, 
      n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, 
      n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, 
      n11447, n11448, n11450, n11451, n11452, n11453, n11454, n11455, n11456, 
      n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, 
      n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, 
      n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, 
      n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11493, 
      n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, 
      n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11512, 
      n11513, n11514, n11515, n11517, n11518, n11519, n11520, n11521, n11522, 
      n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, 
      n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, 
      n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, 
      n11550, n11551, n11553, n11554, n11555, n11556, n11557, n11559, n11560, 
      n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, 
      n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, 
      n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, 
      n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, 
      n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, 
      n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, 
      n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, 
      n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, 
      n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, 
      n11643, n11644, n11645, n11646, n11647, n11648, n11650, n11651, n11652, 
      n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, 
      n11662, n11663, n11664, n11666, n11667, n11668, n11669, n11670, n11671, 
      n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, 
      n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11690, 
      n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, 
      n11700, n11701, n11702, n11703, n11705, n11706, n11707, n11708, n11709, 
      n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, 
      n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, 
      n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, 
      n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, 
      n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, 
      n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, 
      n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, 
      n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, 
      n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11791, 
      n11792, n11793, n11794, n11795, n11796, n11798, n11799, n11800, n11801, 
      n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, 
      n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, 
      n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, 
      n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, 
      n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, 
      n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, 
      n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, 
      n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, 
      n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11883, 
      n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, 
      n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, 
      n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, 
      n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, 
      n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, 
      n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, 
      n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, 
      n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, 
      n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, 
      n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, 
      n11975, n11976, n11977, n11978, n11979, n11981, n11982, n11983, n11984, 
      n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, 
      n11994, n11995, n11996, n11997, n11999, n12000, n12001, n12002, n12003, 
      n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, 
      n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, 
      n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, 
      n12031, n12032, n12033, n12035, n12036, n12037, n12038, n12039, n12040, 
      n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, 
      n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, 
      n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, 
      n12068, n12069, n12070, n12071, n12072, n12073, n12075, n12076, n12077, 
      n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, 
      n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, 
      n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, 
      n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, 
      n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, 
      n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, 
      n12132, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, 
      n12142, n12143, n12144, n12145, n12147, n12148, n12149, n12151, n12152, 
      n12153, n12154, n12155, n12156, n12157, n12159, n12160, n12161, n12162, 
      n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, 
      n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, 
      n12181, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12192, 
      n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, 
      n12202, n12203, n12205, n12206, n12207, n12208, n12209, n12210, n12211, 
      n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, 
      n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, 
      n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, 
      n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, 
      n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, 
      n12257, n12258, n12260, n12261, n12262, n12263, n12264, n12265, n12266, 
      n12267, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, 
      n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12286, 
      n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12295, n12296, 
      n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, 
      n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, 
      n12315, n12316, n12317, n12318, n12319, n12321, n12322, n12323, n12324, 
      n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, 
      n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, 
      n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, 
      n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, 
      n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, 
      n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, 
      n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, 
      n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, 
      n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, 
      n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, 
      n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, 
      n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, 
      n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, 
      n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, 
      n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, 
      n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, 
      n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, 
      n12478, n12479, n12480, n12482, n12483, n12484, n12485, n12486, n12487, 
      n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, 
      n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, 
      n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, 
      n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, 
      n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, 
      n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, 
      n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, 
      n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, 
      n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, 
      n12569, n12570, n12571, n12572, n12573, n12574, n12576, n12577, n12578, 
      n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, 
      n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, 
      n12597, n12598, n12599, n12600, n12601, n12603, n12604, n12605, n12606, 
      n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, 
      n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, 
      n12625, n12626, n12627, n12629, n12630, n12631, n12632, n12633, n12634, 
      n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, 
      n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, 
      n12653, n12654, n12655, n12657, n12658, n12659, n12660, n12661, n12662, 
      n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, 
      n12672, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, 
      n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, 
      n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, 
      n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, 
      n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, 
      n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, 
      n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, 
      n12739, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, 
      n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, 
      n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, 
      n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, 
      n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, 
      n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, 
      n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, 
      n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, 
      n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, 
      n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, 
      n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, 
      n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, 
      n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, 
      n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, 
      n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, 
      n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, 
      n12884, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, 
      n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, 
      n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, 
      n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, 
      n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, 
      n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, 
      n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, 
      n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, 
      n12957, n12958, n12959, n12960, n12961, n12962, n12964, n12965, n12966, 
      n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, 
      n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, 
      n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, 
      n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, 
      n13004, n13005, n13006, n13007, n13008, n13010, n13011, n13012, n13013, 
      n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, 
      n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, 
      n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, 
      n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, 
      n13050, n13051, n13052, n13053, n13055, n13056, n13057, n13058, n13059, 
      n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, 
      n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, 
      n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, 
      n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, 
      n13096, n13097, n13099, n13100, n13101, n13102, n13103, n13104, n13105, 
      n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, 
      n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, 
      n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, 
      n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, 
      n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, 
      n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, 
      n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, 
      n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, 
      n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, 
      n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, 
      n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13204, n13205, 
      n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, 
      n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, 
      n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, 
      n13233, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, 
      n13243, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, 
      n13253, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, 
      n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, 
      n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, 
      n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, 
      n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, 
      n13299, n13300, n13302, n13303, n13304, n13305, n13306, n13307, n13308, 
      n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, 
      n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, 
      n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, 
      n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, 
      n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, 
      n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, 
      n13363, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, 
      n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13382, 
      n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, 
      n13392, n13393, n13396, n13397, n13398, n13399, n13400, n13401, n13402, 
      n13403, n13404, n13405, n13406, n13407, n13409, n13410, n13411, n13412, 
      n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, 
      n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, 
      n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, 
      n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, 
      n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, 
      n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13467, 
      n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, 
      n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, 
      n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, 
      n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, 
      n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, 
      n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, 
      n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, 
      n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, 
      n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, 
      n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, 
      n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, 
      n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, 
      n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, 
      n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, 
      n13595, n13596, n13597, n13598, n13600, n13601, n13602, n13603, n13604, 
      n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, 
      n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, 
      n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, 
      n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, 
      n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, 
      n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, 
      n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, 
      n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, 
      n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, 
      n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, 
      n13695, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, 
      n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, 
      n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, 
      n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, 
      n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, 
      n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, 
      n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, 
      n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, 
      n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, 
      n13778, n13779, n13780, n13781, n13783, n13784, n13785, n13786, n13787, 
      n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13797, 
      n13798, n13799, n13800, n13801, n13802, n13804, n13805, n13806, n13807, 
      n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, 
      n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, 
      n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, 
      n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, 
      n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, 
      n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, 
      n13863, n13864, n13865, n13866, n13867, n13868, n13870, n13871, n13872, 
      n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, 
      n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, 
      n13891, n13892, n13893, n13895, n13896, n13897, n13898, n13899, n13900, 
      n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, 
      n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, 
      n13919, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, 
      n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, 
      n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, 
      n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, 
      n13956, n13957, n13958, n13959, n13960, n13961, n13963, n13964, n13965, 
      n13966, n13967, n13968, n13969, n13970, n13971, n13973, n13974, n13975, 
      n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, 
      n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, 
      n13994, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, 
      n14004, n14005, n14006, n14007, n14008, n14010, n14011, n14012, n14013, 
      n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, 
      n14023, n14024, n14025, n14027, n14028, n14029, n14030, n14031, n14032, 
      n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, 
      n14042, n14043, n14044, n14045, n14047, n14049, n14050, n14051, n14052, 
      n14053, n14054, n14056, n14057, n14058, n14059, n14060, n14061, n14062, 
      n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14072, 
      n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, 
      n14082, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, 
      n14092, n14093, n14094, n14095, n14096, n14098, n14099, n14100, n14101, 
      n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, 
      n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, 
      n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, 
      n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, 
      n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, 
      n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, 
      n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, 
      n14165, n14166, n14167, n14168, n14171, n14172, n14173, n14174, n14176, 
      n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, 
      n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, 
      n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14203, n14204, 
      n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, 
      n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, 
      n14225, n14226, n14227, n14228, n14229, n14230, n14232, n14233, n14234, 
      n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, 
      n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, 
      n14253, n14254, n14255, n14257, n14258, n14259, n14260, n14261, n14262, 
      n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, 
      n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, 
      n14281, n14282, n14283, n14284, n14285, n14287, n14288, n14289, n14290, 
      n14291, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, 
      n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, 
      n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, 
      n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, 
      n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, 
      n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, 
      n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, 
      n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, 
      n14365, n14367, n14368, n14369, n14371, n14372, n14373, n14374, n14375, 
      n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, 
      n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, 
      n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14403, 
      n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, 
      n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, 
      n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, 
      n14431, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, 
      n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, 
      n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, 
      n14459, n14460, n14461, n14462, n14464, n14465, n14466, n14467, n14468, 
      n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, 
      n14478, n14479, n14480, n14481, n14482, n14483, n14485, n14486, n14487, 
      n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, 
      n14497, n14498, n14499, n14501, n14502, n14504, n14505, n14506, n14507, 
      n14508, n14509, n14511, n14512, n14513, n14514, n14515, n14516, n14518, 
      n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, 
      n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, 
      n14537, n14538, n14539, n14542, n14543, n14544, n14545, n14546, n14547, 
      n14548, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, 
      n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, 
      n14567, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, 
      n14577, n14578, n14580, n14581, n14582, n14583, n14584, n14585, n14586, 
      n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14596, 
      n14597, n14598, n14599, n14600, n14601, n14603, n14604, n14606, n14607, 
      n14608, n14609, n14611, n14612, n14613, n14614, n14615, n14616, n14617, 
      n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, 
      n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, 
      n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, 
      n14645, n14646, n14648, n14649, n14651, n14652, n14653, n14654, n14655, 
      n14656, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, 
      n14666, n14667, n14668, n14669, n14670, n14671, n14673, n14674, n14675, 
      n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, 
      n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, 
      n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, 
      n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, 
      n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, 
      n14722, n14723, n14724, n14726, n14727, n14728, n14729, n14730, n14731, 
      n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, 
      n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, 
      n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, 
      n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, 
      n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14778, 
      n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, 
      n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14796, n14797, 
      n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, 
      n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, 
      n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14826, 
      n14827, n14828, n14829, n14831, n14832, n14833, n14834, n14835, n14836, 
      n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, 
      n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, 
      n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, 
      n14864, n14865, n14866, n14868, n14869, n14870, n14871, n14872, n14873, 
      n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, 
      n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, 
      n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, 
      n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, 
      n14911, n14913, n14914, n14915, n14916, n14917, n14918, n14920, n14921, 
      n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, 
      n14931, n14932, n14933, n14935, n14936, n14937, n14938, n14939, n14940, 
      n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, 
      n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, 
      n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, 
      n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, 
      n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14986, n14987, 
      n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14997, 
      n14998, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, 
      n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, 
      n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, 
      n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, 
      n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, 
      n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, 
      n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, 
      n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, 
      n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, 
      n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, 
      n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, 
      n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, 
      n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, 
      n15117, n15118, n15119, n15120, n15121, n15123, n15124, n15125, n15126, 
      n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, 
      n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, 
      n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, 
      n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, 
      n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, 
      n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, 
      n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, 
      n15190, n15191, n15192, n15193, n15195, n15196, n15197, n15198, n15199, 
      n15200, n15201, n15203, n15204, n15205, n15206, n15207, n15208, n15209, 
      n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, 
      n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, 
      n15228, n15229, n15230, n15231, n15233, n15234, n15235, n15236, n15237, 
      n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, 
      n15247, n15248, n15249, n15250, n15252, n15253, n15254, n15255, n15256, 
      n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, 
      n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15274, n15275, 
      n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, 
      n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, 
      n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, 
      n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, 
      n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, 
      n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, 
      n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, 
      n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, 
      n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, 
      n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, 
      n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, 
      n15375, n15376, n15377, n15378, n15379, n15380, n15382, n15383, n15384, 
      n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, 
      n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, 
      n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, 
      n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, 
      n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, 
      n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, 
      n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, 
      n15449, n15450, n15451, n15453, n15454, n15456, n15457, n15458, n15459, 
      n15460, n15461, n15462, n15463, n15465, n15466, n15467, n15468, n15469, 
      n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, 
      n15479, n15480, n15481, n15482, n15483, n15485, n15487, n15488, n15489, 
      n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, 
      n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, 
      n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, 
      n15517, n15518, n15519, n15521, n15522, n15523, n15524, n15525, n15526, 
      n15527, n15528, n15529, n15530, n15531, n15532, n15534, n15535, n15536, 
      n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, 
      n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, 
      n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, 
      n15564, n15565, n15566, n15567, n15568, n15570, n15571, n15572, n15573, 
      n15574, n15575, n15576, n15577, n15578, n15579, n15581, n15582, n15583, 
      n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, 
      n15593, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, 
      n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, 
      n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, 
      n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, 
      n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, 
      n15640, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, 
      n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, 
      n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, 
      n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, 
      n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, 
      n15686, n15687, n15689, n15690, n15691, n15692, n15693, n15694, n15695, 
      n15696, n15697, n15698, n15700, n15701, n15702, n15703, n15704, n15705, 
      n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, 
      n15715, n15716, n15718, n15719, n15720, n15721, n15722, n15723, n15724, 
      n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15733, n15734, 
      n15735, n15736, n15737, n15739, n15740, n15741, n15742, n15743, n15744, 
      n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, 
      n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, 
      n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, 
      n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15782, 
      n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, 
      n15793, n15794, n15796, n15797, n15798, n15800, n15801, n15802, n15803, 
      n15804, n15805, n15807, n15808, n15809, n15810, n15811, n15812, n15813, 
      n15814, n15815, n15816, n15817, n15819, n15820, n15821, n15822, n15823, 
      n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, 
      n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, 
      n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, 
      n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, 
      n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15869, 
      n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, 
      n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, 
      n15888, n15889, n15890, n15891, n15892, n15895, n15896, n15897, n15898, 
      n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, 
      n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, 
      n15917, n15919, n15920, n15921, n15923, n15924, n15925, n15926, n15927, 
      n15928, n15929, n15930, n15932, n15933, n15934, n15935, n15936, n15937, 
      n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, 
      n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, 
      n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, 
      n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, 
      n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, 
      n15983, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, 
      n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, 
      n16002, n16003, n16004, n16005, n16006, n16007, n16009, n16010, n16011, 
      n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, 
      n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, 
      n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, 
      n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, 
      n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, 
      n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, 
      n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, 
      n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, 
      n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, 
      n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, 
      n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, 
      n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, 
      n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, 
      n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, 
      n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, 
      n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, 
      n16159, n16160, n16161, n16163, n16164, n16165, n16166, n16167, n16168, 
      n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, 
      n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, 
      n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, 
      n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, 
      n16206, n16207, n16208, n16209, n16210, n16211, n16213, n16214, n16215, 
      n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, 
      n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, 
      n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, 
      n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16251, n16253, 
      n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, 
      n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, 
      n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, 
      n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, 
      n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, 
      n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, 
      n16308, n16309, n16310, n16311, n16312, n16314, n16315, n16316, n16317, 
      n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, 
      n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, 
      n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, 
      n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, 
      n16354, n16355, n16356, n16357, n16359, n16360, n16361, n16362, n16363, 
      n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16373, 
      n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, 
      n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, 
      n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, 
      n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, 
      n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, 
      n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, 
      n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, 
      n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, 
      n16449, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, 
      n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, 
      n16468, n16469, n16470, n16471, n16472, n16473, n16476, n16477, n16478, 
      n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, 
      n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, 
      n16497, n16498, n16499, n16500, n16501, n16503, n16504, n16505, n16506, 
      n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, 
      n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, 
      n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, 
      n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, 
      n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, 
      n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, 
      n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, 
      n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16579, 
      n16580, n16581, n16583, n16584, n16585, n16586, n16587, n16588, n16589, 
      n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, 
      n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, 
      n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, 
      n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, 
      n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, 
      n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, 
      n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, 
      n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, 
      n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, 
      n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, 
      n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, 
      n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, 
      n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, 
      n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, 
      n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, 
      n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, 
      n16735, n16736, n16737, n16738, n16739, n16741, n16742, n16743, n16744, 
      n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, 
      n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, 
      n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, 
      n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, 
      n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, 
      n16790, n16791, n16792, n16794, n16795, n16796, n16797, n16798, n16799, 
      n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, 
      n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, 
      n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, 
      n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, 
      n16836, n16837, n16838, n16839, n16840, n16842, n16843, n16844, n16845, 
      n16846, n16847, n16848, n16849, n16851, n16852, n16853, n16854, n16855, 
      n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, 
      n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, 
      n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, 
      n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, 
      n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, 
      n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, 
      n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, 
      n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, 
      n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, 
      n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, 
      n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, 
      n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, 
      n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, 
      n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, 
      n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, 
      n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, 
      n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, 
      n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, 
      n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, 
      n17028, n17029, n17030, n17031, n17032, n17034, n17035, n17036, n17037, 
      n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, 
      n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, 
      n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, 
      n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, 
      n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17082, n17083, 
      n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, 
      n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, 
      n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, 
      n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, 
      n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, 
      n17129, n17130, n17131, n17132, n17133, n17135, n17136, n17138, n17139, 
      n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, 
      n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, 
      n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, 
      n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, 
      n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, 
      n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, 
      n17194, n17195, n17196, n17197, n17198, n17200, n17201, n17202, n17203, 
      n17204, n17205, n17206, n17208, n17209, n17210, n17211, n17212, n17213, 
      n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, 
      n17223, n17224, n17225, n17227, n17228, n17229, n17230, n17231, n17232, 
      n17233, n17234, n17235, n17236, n17238, n17240, n17241, n17242, n17243, 
      n17244, n17245, n17246, n17247, n17249, n17250, n17251, n17252, n17253, 
      n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17263, 
      n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, 
      n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, 
      n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, 
      n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, 
      n17300, n17301, n17302, n17303, n17307, n17308, n17309, n17310, n17311, 
      n17312, n17313, n17315, n17316, n17317, n17318, n17319, n17320, n17321, 
      n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, 
      n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, 
      n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, 
      n17349, n17350, n17351, n17352, n17353, n17355, n17356, n17357, n17358, 
      n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, 
      n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, 
      n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, 
      n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, 
      n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, 
      n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, 
      n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, 
      n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, 
      n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, 
      n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, 
      n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, 
      n17458, n17459, n17460, n17461, n17463, n17464, n17465, n17466, n17467, 
      n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, 
      n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, 
      n17486, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, 
      n17496, n17497, n17498, n17499, n17501, n17502, n17503, n17504, n17505, 
      n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, 
      n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, 
      n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, 
      n17533, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, 
      n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, 
      n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, 
      n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, 
      n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, 
      n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, 
      n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, 
      n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, 
      n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, 
      n17615, n17616, n17617, n17618, n17620, n17621, n17622, n17623, n17624, 
      n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, 
      n17634, n17635, n17637, n17638, n17639, n17640, n17641, n17642, n17643, 
      n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, 
      n17653, n17654, n17656, n17658, n17659, n17661, n17662, n17663, n17664, 
      n17665, n17666, n17667, n17668, n17669, n17670, n17672, n17673, n17674, 
      n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, 
      n17684, n17685, n17686, n17687, n17688, n17690, n17691, n17692, n17693, 
      n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, 
      n17703, n17705, n17706, n17707, n17708, n17709, n17710, n17712, n17713, 
      n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, 
      n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17731, n17732, 
      n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, 
      n17742, n17743, n17745, n17746, n17747, n17748, n17749, n17750, n17751, 
      n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, 
      n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, 
      n17770, n17771, n17772, n17773, n17774, n17776, n17777, n17778, n17779, 
      n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, 
      n17789, n17790, n17791, n17793, n17794, n17795, n17796, n17797, n17799, 
      n17800, n17802, n17803, n17804, n17805, n17807, n17808, n17809, n17810, 
      n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, 
      n17820, n17822, n17823, n17824, n17825, n17826, n17828, n17829, n17830, 
      n17831, n17832, n17833, n17834, n17835, n17836, n17838, n17839, n17840, 
      n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, 
      n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, 
      n17860, n17861, n17863, n17864, n17865, n17866, n17867, n17868, n17869, 
      n17872, n17873, n17874, n17875, n17876, n17878, n17879, n17881, n17882, 
      n17883, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, 
      n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, 
      n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, 
      n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, 
      n17921, n17922, n17923, n17925, n17927, n17928, n17929, n17930, n17931, 
      n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, 
      n17941, n17943, n17944, n17945, n17946, n17950, n17951, n17952, n17953, 
      n17954, n17955, n17956, n17957, n17958, n17959, n17961, n17962, n17963, 
      n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, 
      n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, 
      n17982, n17983, n17985, n17986, n17987, n17988, n17989, n17991, n17992, 
      n17993, n17994, n17996, n17997, n17998, n17999, n18000, n18001, n18002, 
      n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, 
      n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, 
      n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18032, 
      n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18042, 
      n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, 
      n18052, n18054, n18055, n18057, n18058, n18059, n18060, n18061, n18062, 
      n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, 
      n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18080, n18081, 
      n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, 
      n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, 
      n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18109, 
      n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18119, 
      n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, 
      n18129, n18130, n18131, n18133, n18134, n18135, n18136, n18137, n18138, 
      n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, 
      n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, 
      n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, 
      n18166, n18168, n18169, n18170, n18171, n18172, n18174, n18175, n18176, 
      n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, 
      n18186, n18187, n18188, n18190, n18191, n18192, n18193, n18194, n18195, 
      n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, 
      n18205, n18206, n18207, n18208, n18209, n18211, n18212, n18213, n18214, 
      n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18223, n18224, 
      n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, 
      n18234, n18235, n18236, n18237, n18238, n18240, n18241, n18245, n18246, 
      n18247, n18248, n18249, n18250, n18251, n18254, n18255, n18256, n18257, 
      n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, 
      n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, 
      n18276, n18277, n18278, n18279, n18281, n18282, n18283, n18284, n18285, 
      n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, 
      n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, 
      n18304, n18305, n18306, n18307, n18308, n18309, n18311, n18313, n18314, 
      n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, 
      n18324, n18325, n18326, n18327, n18328, n18329, n18331, n18332, n18333, 
      n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, 
      n18343, n18344, n18345, n18346, n18348, n18349, n18350, n18351, n18352, 
      n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, 
      n18362, n18364, n18365, n18366, n18367, n18368, n18369, n18371, n18372, 
      n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18381, n18382, 
      n18383, n18384, n18385, n18386, n18387, n18389, n18392, n18393, n18394, 
      n18395, n18396, n18397, n18398, n18399, n18400, n18402, n18403, n18404, 
      n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, 
      n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, 
      n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18433, 
      n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, 
      n18443, n18444, n18445, n18446, n18448, n18449, n18450, n18451, n18453, 
      n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18463, 
      n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, 
      n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, 
      n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18491, 
      n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, 
      n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18509, n18510, 
      n18511, n18512, n18513, n18514, n18515, n18517, n18518, n18519, n18520, 
      n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, 
      n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, 
      n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, 
      n18548, n18549, n18551, n18552, n18553, n18554, n18555, n18556, n18557, 
      n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, 
      n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18575, n18576, 
      n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, 
      n18587, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, 
      n18597, n18598, n18599, n18600, n18601, n18603, n18604, n18605, n18606, 
      n18607, n18608, n18609, n18610, n18612, n18613, n18614, n18615, n18616, 
      n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, 
      n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, 
      n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18644, 
      n18645, n18646, n18647, n18648, n18650, n18651, n18652, n18653, n18654, 
      n18655, n18656, n18658, n18659, n18660, n18661, n18662, n18663, n18664, 
      n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, 
      n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18682, n18683, 
      n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18693, 
      n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, 
      n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18711, n18712, 
      n18713, n18714, n18715, n18716, n18717, n18719, n18720, n18721, n18722, 
      n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, 
      n18732, n18733, n18735, n18736, n18737, n18741, n18742, n18743, n18744, 
      n18745, n18746, n18747, n18749, n18750, n18751, n18752, n18753, n18754, 
      n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, 
      n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, 
      n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, 
      n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, 
      n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, 
      n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, 
      n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, 
      n18819, n18820, n18822, n18823, n18825, n18826, n18827, n18829, n18830, 
      n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, 
      n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, 
      n18849, n18850, n18852, n18853, n18854, n18855, n18856, n18857, n18858, 
      n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18868, 
      n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, 
      n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, 
      n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, 
      n18896, n18897, n18898, n18899, n18901, n18902, n18903, n18904, n18905, 
      n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, 
      n18916, n18917, n18918, n18919, n18920, n18921, n18923, n18924, n18925, 
      n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, 
      n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, 
      n18944, n18946, n18948, n18949, n18950, n18951, n18952, n18953, n18954, 
      n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, 
      n18964, n18965, n18966, n18967, n18968, n18970, n18971, n18972, n18973, 
      n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18983, 
      n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, 
      n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19001, n19002, 
      n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, 
      n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, 
      n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, 
      n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, 
      n19040, n19041, n19042, n19043, n19045, n19046, n19047, n19048, n19049, 
      n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, 
      n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, 
      n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, 
      n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, 
      n19086, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, 
      n19096, n19097, n19098, n19100, n19101, n19102, n19103, n19105, n19106, 
      n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19115, n19116, 
      n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, 
      n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, 
      n19135, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, 
      n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, 
      n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, 
      n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, 
      n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, 
      n19181, n19182, n19183, n19185, n19186, n19187, n19188, n19189, n19190, 
      n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, 
      n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, 
      n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, 
      n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19227, 
      n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, 
      n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, 
      n19246, n19247, n19248, n19249, n19250, n19251, n19253, n19254, n19255, 
      n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, 
      n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, 
      n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, 
      n19283, n19284, n19285, n19286, n19288, n19290, n19291, n19292, n19293, 
      n19294, n19295, n19296, n19297, n19298, n19299, n19301, n19302, n19303, 
      n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, 
      n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, 
      n19322, n19324, n19325, n19326, n19327, n19329, n19330, n19331, n19332, 
      n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, 
      n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19351, 
      n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, 
      n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, 
      n19370, n19371, n19372, n19373, n19374, n19375, n19377, n19378, n19379, 
      n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, 
      n19389, n19390, n19391, n19392, n19393, n19395, n19396, n19397, n19398, 
      n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, 
      n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, 
      n19418, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, 
      n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, 
      n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, 
      n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19456, 
      n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, 
      n19466, n19467, n19468, n19472, n19474, n19475, n19476, n19485, n19488, 
      n19490, n19492, n19496, n19501, n19502, n19503, n19504, n19505, n19506, 
      n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, 
      n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, 
      n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, 
      n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, 
      n19543, n19544, n19546, n19547, n19548, n19549, n19550, n19551, n19552, 
      n19553, n19554, n19555, n19557, n19558, n19559, n19561, n19562, n19563, 
      n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19573, 
      n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, 
      n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, 
      n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, 
      n19601, n19602, n19603, n19604, n19606, n19607, n19608, n19609, n19610, 
      n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, 
      n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19629, 
      n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, 
      n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, 
      n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, 
      n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, 
      n19666, n19667, n19668, n19669, n19670, n19672, n19673, n19674, n19675, 
      n19676, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, 
      n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, 
      n19695, n19697, n19698, n19699, n19700, n19702, n19703, n19704, n19705, 
      n19706, n19707, n19708, n19709, n19710, n19711, n19713, n19715, n19716, 
      n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, 
      n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, 
      n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, 
      n19744, n19745, n19746, n19748, n19749, n19750, n19751, n19752, n19753, 
      n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19763, 
      n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19773, 
      n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, 
      n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, 
      n19792, n19794, n19796, n19797, n19798, n19799, n19802, n19803, n19804, 
      n19805, n19806, n19807, n19809, n19811, n19812, n19813, n19814, n19815, 
      n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, 
      n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, 
      n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, 
      n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, 
      n19854, n19855, n19856, n19857, n19859, n19860, n19861, n19862, n19863, 
      n19864, n19865, n19866, n19867, n19868, n19869, n19871, n19872, n19874, 
      n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, 
      n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, 
      n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, 
      n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, 
      n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, 
      n19921, n19922, n19923, n19924, n19925, n19927, n19928, n19929, n19930, 
      n19931, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, 
      n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, 
      n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, 
      n19962, n19963, n19964, n19966, n19967, n19968, n19969, n19970, n19971, 
      n19972, n19973, n19974, n19975, n19977, n19978, n19979, n19980, n19983, 
      n19984, n19985, n19986, n19988, n19989, n19990, n19992, n19993, n19997, 
      n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, 
      n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, 
      n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, 
      n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, 
      n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, 
      n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, 
      n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, 
      n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, 
      n20070, n20071, n20072, n20073, n20074, n20076, n20077, n20079, n20080, 
      n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, 
      n20091, n20092, n20093, n20094, n20095, n20097, n20098, n20099, n20100, 
      n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, 
      n20110, n20111, n20112, n20113, n20114, n20115, n20117, n20119, n20120, 
      n20121, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, 
      n20131, n20132, n20133, n20134, n20135, n20138, n20139, n20140, n20141, 
      n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, 
      n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, 
      n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, 
      n20169, n20170, n20171, n20172, n20173, n20174, n20176, n20177, n20178, 
      n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, 
      n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, 
      n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, 
      n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, 
      n20216, n20217, n20218, n20219, n20221, n20222, n20223, n20224, n20225, 
      n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, 
      n20235, n20236, n20237, n20239, n20240, n20241, n20242, n20243, n20244, 
      n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20256, 
      n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, 
      n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, 
      n20275, n20276, n20277, n20278, n20279, n20281, n20282, n20283, n20284, 
      n20285, n20286, n20288, n20290, n20291, n20292, n20293, n20294, n20295, 
      n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, 
      n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, 
      n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, 
      n20324, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, 
      n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, 
      n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, 
      n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, 
      n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, 
      n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, 
      n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, 
      n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, 
      n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, 
      n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, 
      n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, 
      n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, 
      n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, 
      n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, 
      n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, 
      n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, 
      n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, 
      n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, 
      n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, 
      n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, 
      n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, 
      n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, 
      n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, 
      n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, 
      n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, 
      n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, 
      n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, 
      n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, 
      n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, 
      n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, 
      n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, 
      n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, 
      n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, 
      n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, 
      n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, 
      n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, 
      n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, 
      n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, 
      n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, 
      n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, 
      n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, 
      n20694, n20695, n20696, n20697 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n19081, A2 => n19082, ZN => n1);
   U2 : OR2_X1 port map( A1 => n17858, A2 => n15, ZN => n14);
   U8 : AND2_X1 port map( A1 => n18948, A2 => n17812, ZN => n20);
   U9 : AND3_X1 port map( A1 => n3414, A2 => n3413, A3 => n15736, ZN => n16988)
                           ;
   U11 : NAND2_X1 port map( A1 => n14372, A2 => n2720, ZN => n16406);
   U12 : OAI21_X1 port map( B1 => n15862, B2 => n15864, A => n9, ZN => n15173);
   U13 : AND2_X1 port map( A1 => n15720, A2 => n15861, ZN => n15328);
   U20 : OR2_X1 port map( A1 => n13909, A2 => n14611, ZN => n133);
   U21 : OR2_X1 port map( A1 => n15121, A2 => n14520, ZN => n14320);
   U22 : BUF_X1 port map( A => n12911, Z => n14439);
   U28 : OR2_X1 port map( A1 => n12606, A2 => n12237, ZN => n12604);
   U29 : OR2_X1 port map( A1 => n19833, A2 => n12479, ZN => n6);
   U30 : AND2_X1 port map( A1 => n12207, A2 => n12208, ZN => n4);
   U32 : BUF_X1 port map( A => n10625, Z => n11820);
   U33 : INV_X1 port map( A => n11598, ZN => n11828);
   U34 : AND2_X1 port map( A1 => n3630, A2 => n3629, ZN => n122);
   U36 : OR2_X1 port map( A1 => n10960, A2 => n20366, ZN => n142);
   U37 : INV_X1 port map( A => n20366, ZN => n143);
   U39 : OR2_X1 port map( A1 => n11365, A2 => n10677, ZN => n2765);
   U41 : NOR2_X1 port map( A1 => n9570, A2 => n9569, ZN => n9843);
   U43 : OR2_X1 port map( A1 => n8547, A2 => n8546, ZN => n10339);
   U45 : OR2_X1 port map( A1 => n8946, A2 => n111, ZN => n109);
   U47 : AND3_X1 port map( A1 => n6957, A2 => n6956, A3 => n6955, ZN => n9163);
   U49 : INV_X1 port map( A => n8127, ZN => n9088);
   U53 : OR2_X1 port map( A1 => n7507, A2 => n7508, ZN => n1540);
   U54 : XNOR2_X1 port map( A => n6040, B => n6732, ZN => n8193);
   U55 : XNOR2_X1 port map( A => n7070, B => n6947, ZN => n6770);
   U57 : CLKBUF_X1 port map( A => Key(108), Z => n19027);
   U59 : OAI21_X1 port map( B1 => n19790, B2 => n5929, A => n41, ZN => n5597);
   U60 : OAI21_X1 port map( B1 => n6060, B2 => n6061, A => n6059, ZN => n6062);
   U61 : OR2_X1 port map( A1 => n5349, A2 => n6150, ZN => n6154);
   U63 : INV_X1 port map( A => n6042, ZN => n135);
   U64 : INV_X1 port map( A => n5632, ZN => n31);
   U65 : INV_X1 port map( A => n5215, ZN => n32);
   U66 : OR2_X1 port map( A1 => n4174, A2 => n4175, ZN => n117);
   U69 : AND2_X1 port map( A1 => n4819, A2 => n4820, ZN => n5953);
   U70 : NAND2_X1 port map( A1 => n2215, A2 => n2214, ZN => n6017);
   U71 : OR2_X1 port map( A1 => n5038, A2 => n303, ZN => n1320);
   U72 : AND2_X1 port map( A1 => n4524, A2 => n4342, ZN => n87);
   U74 : OR2_X1 port map( A1 => n176, A2 => n4685, ZN => n4487);
   U76 : AND2_X1 port map( A1 => n4313, A2 => n4601, ZN => n29);
   U78 : NAND2_X2 port map( A1 => n1186, A2 => n8561, ZN => n10171);
   U80 : OAI211_X1 port map( C1 => n11791, C2 => n14588, A => n108, B => n107, 
                           ZN => n12658);
   U83 : OAI21_X1 port map( B1 => n16679, B2 => n132, A => n131, ZN => n17675);
   U85 : AND2_X1 port map( A1 => n19056, A2 => n19071, ZN => n70);
   U88 : OR2_X1 port map( A1 => n18935, A2 => n18936, ZN => n7);
   U90 : INV_X1 port map( A => n19400, ZN => n2);
   U92 : OR2_X1 port map( A1 => n14010, A2 => n14406, ZN => n35);
   U93 : NOR3_X1 port map( A1 => n19292, A2 => n19283, A3 => n19282, ZN => 
                           n19294);
   U94 : OR2_X1 port map( A1 => n19290, A2 => n19304, ZN => n138);
   U95 : XNOR2_X1 port map( A => n13834, B => n13079, ZN => n13389);
   U96 : OAI22_X2 port map( A1 => n15472, A2 => n15471, B1 => n15470, B2 => 
                           n20503, ZN => n17298);
   U102 : INV_X1 port map( A => n3516, ZN => n139);
   U103 : INV_X1 port map( A => n701, ZN => n14443);
   U106 : XNOR2_X1 port map( A => n6915, B => n6916, ZN => n8342);
   U107 : AND2_X1 port map( A1 => n14601, A2 => n14250, ZN => n14248);
   U110 : OR2_X1 port map( A1 => n19402, A2 => n17650, ZN => n81);
   U118 : AND2_X1 port map( A1 => n19021, A2 => n19009, ZN => n19004);
   U123 : AND2_X1 port map( A1 => n6064, A2 => n5304, ZN => n6061);
   U125 : AOI21_X1 port map( B1 => n16638, B2 => n19353, A => n16637, ZN => 
                           n17935);
   U128 : AND2_X1 port map( A1 => n17656, A2 => n19396, ZN => n3);
   U130 : INV_X1 port map( A => n16306, ZN => n17);
   U131 : OR2_X1 port map( A1 => n19360, A2 => n17861, ZN => n132);
   U132 : NOR2_X1 port map( A1 => n15896, A2 => n15538, ZN => n15890);
   U133 : BUF_X1 port map( A => n15896, Z => n15402);
   U134 : INV_X1 port map( A => n14792, ZN => n12627);
   U138 : OR2_X1 port map( A1 => n15266, A2 => n15845, ZN => n717);
   U139 : NAND2_X2 port map( A1 => n14745, A2 => n14744, ZN => n17294);
   U143 : OAI21_X2 port map( B1 => n15231, B2 => n15449, A => n15230, ZN => 
                           n16861);
   U144 : OR2_X1 port map( A1 => n8542, A2 => n9066, ZN => n8860);
   U146 : NAND2_X1 port map( A1 => n19080, A2 => n1, ZN => n19084);
   U147 : OAI21_X1 port map( B1 => n19511, B2 => n3, A => n2, ZN => n17658);
   U149 : INV_X1 port map( A => n17856, ZN => n18);
   U150 : OAI21_X1 port map( B1 => n1690, B2 => n8179, A => n1851, ZN => n8796)
                           ;
   U152 : NAND2_X1 port map( A1 => n12211, A2 => n4, ZN => n12218);
   U156 : OR2_X2 port map( A1 => n5538, A2 => n5537, ZN => n5736);
   U158 : AND2_X2 port map( A1 => n2750, A2 => n1002, ZN => n2749);
   U160 : NAND2_X1 port map( A1 => n11223, A2 => n6, ZN => n12784);
   U162 : NAND2_X1 port map( A1 => n3607, A2 => n3752, ZN => n3658);
   U163 : OR2_X1 port map( A1 => n352, A2 => n9563, ZN => n2170);
   U169 : NAND3_X1 port map( A1 => n18933, A2 => n18934, A3 => n7, ZN => n2062)
                           ;
   U170 : NAND2_X1 port map( A1 => n8, A2 => n1912, ZN => n8330);
   U172 : NAND2_X1 port map( A1 => n4825, A2 => n4826, ZN => n4831);
   U174 : NAND2_X1 port map( A1 => n15862, A2 => n15327, ZN => n9);
   U176 : NAND2_X1 port map( A1 => n18923, A2 => n11, ZN => n18925);
   U177 : NAND2_X1 port map( A1 => n18920, A2 => n18921, ZN => n11);
   U178 : XNOR2_X2 port map( A => n16910, B => n16909, ZN => n18221);
   U182 : NAND2_X1 port map( A1 => n9527, A2 => n9530, ZN => n9754);
   U186 : NAND4_X2 port map( A1 => n5127, A2 => n5126, A3 => n5125, A4 => n1096
                           , ZN => n7179);
   U188 : AND3_X2 port map( A1 => n1251, A2 => n1249, A3 => n1447, ZN => n13577
                           );
   U190 : XNOR2_X2 port map( A => n16100, B => n16099, ZN => n17891);
   U194 : NAND2_X1 port map( A1 => n1487, A2 => n8832, ZN => n2150);
   U195 : INV_X1 port map( A => n14285, ZN => n15066);
   U199 : OR2_X1 port map( A1 => n11664, A2 => n121, ZN => n11666);
   U200 : NOR2_X2 port map( A1 => n16, A2 => n14, ZN => n19242);
   U202 : NOR2_X1 port map( A1 => n18, A2 => n17, ZN => n16);
   U205 : NAND3_X1 port map( A1 => n5928, A2 => n6027, A3 => n5929, ZN => n19);
   U206 : INV_X2 port map( A => n8129, ZN => n9451);
   U208 : MUX2_X2 port map( A => n12086, B => n12085, S => n12416, Z => n12906)
                           ;
   U209 : NAND2_X1 port map( A1 => n18047, A2 => n20, ZN => n3544);
   U210 : NAND2_X1 port map( A1 => n24, A2 => n21, ZN => n7523);
   U211 : NAND2_X1 port map( A1 => n23, A2 => n22, ZN => n21);
   U212 : INV_X1 port map( A => n7922, ZN => n22);
   U213 : NAND2_X1 port map( A1 => n2176, A2 => n776, ZN => n23);
   U214 : NAND2_X1 port map( A1 => n7521, A2 => n7922, ZN => n24);
   U219 : NAND2_X1 port map( A1 => n15740, A2 => n26, ZN => n25);
   U220 : INV_X1 port map( A => n15751, ZN => n26);
   U222 : NAND3_X1 port map( A1 => n12068, A2 => n12069, A3 => n1878, ZN => 
                           n13710);
   U227 : NAND2_X1 port map( A1 => n1938, A2 => n13892, ZN => n1352);
   U228 : INV_X1 port map( A => n6117, ZN => n6122);
   U229 : NAND2_X1 port map( A1 => n5868, A2 => n6118, ZN => n6117);
   U230 : NAND2_X1 port map( A1 => n4354, A2 => n29, ZN => n4314);
   U233 : NAND2_X1 port map( A1 => n32, A2 => n31, ZN => n30);
   U235 : OAI21_X1 port map( B1 => n12032, B2 => n12033, A => n12272, ZN => n33
                           );
   U237 : NAND2_X1 port map( A1 => n703, A2 => n12185, ZN => n1981);
   U239 : AOI21_X1 port map( B1 => n11374, B2 => n11375, A => n11373, ZN => 
                           n12552);
   U241 : OR2_X1 port map( A1 => n7965, A2 => n20490, ZN => n8019);
   U242 : AOI21_X1 port map( B1 => n34, B2 => n5530, A => n5529, ZN => n5536);
   U243 : NAND2_X1 port map( A1 => n2940, A2 => n5569, ZN => n34);
   U248 : NAND2_X1 port map( A1 => n14007, A2 => n14236, ZN => n36);
   U250 : OR2_X1 port map( A1 => n11995, A2 => n11820, ZN => n12327);
   U251 : NAND3_X1 port map( A1 => n261, A2 => n9151, A3 => n2499, ZN => n391);
   U254 : OAI21_X1 port map( B1 => n3028, B2 => n19989, A => n679, ZN => n18862
                           );
   U258 : NAND3_X1 port map( A1 => n15794, A2 => n15791, A3 => n859, ZN => 
                           n2309);
   U265 : NAND2_X1 port map( A1 => n14211, A2 => n14213, ZN => n14084);
   U267 : OR2_X1 port map( A1 => n11921, A2 => n11920, ZN => n40);
   U269 : NAND2_X1 port map( A1 => n19790, A2 => n6025, ZN => n41);
   U270 : OAI21_X1 port map( B1 => n8814, B2 => n8812, A => n8810, ZN => n44);
   U271 : INV_X1 port map( A => n9119, ZN => n45);
   U272 : NOR2_X1 port map( A1 => n14441, A2 => n20262, ZN => n140);
   U273 : OAI22_X1 port map( A1 => n11126, A2 => n19949, B1 => n10814, B2 => 
                           n2729, ZN => n11128);
   U274 : OAI21_X1 port map( B1 => n48, B2 => n15150, A => n46, ZN => n14922);
   U275 : NAND2_X1 port map( A1 => n15713, A2 => n19514, ZN => n46);
   U277 : NAND2_X1 port map( A1 => n49, A2 => n20178, ZN => n48);
   U278 : INV_X1 port map( A => n15712, ZN => n49);
   U286 : NAND2_X1 port map( A1 => n1764, A2 => n5114, ZN => n4068);
   U288 : AOI22_X1 port map( A1 => n3703, A2 => n2749, B1 => n19606, B2 => 
                           n8544, ZN => n88);
   U290 : NAND2_X1 port map( A1 => n52, A2 => n50, ZN => n18071);
   U291 : NAND2_X1 port map( A1 => n18069, A2 => n17091, ZN => n50);
   U292 : NAND2_X1 port map( A1 => n18068, A2 => n2516, ZN => n52);
   U294 : NAND3_X2 port map( A1 => n11123, A2 => n11122, A3 => n2033, ZN => 
                           n12463);
   U295 : XNOR2_X1 port map( A => n13222, B => n13724, ZN => n13761);
   U298 : AOI21_X1 port map( B1 => n53, B2 => n19891, A => n15256, ZN => n15000
                           );
   U299 : NAND2_X1 port map( A1 => n2223, A2 => n19931, ZN => n53);
   U302 : NAND2_X1 port map( A1 => n15201, A2 => n3431, ZN => n55);
   U304 : NAND2_X1 port map( A1 => n15200, A2 => n15495, ZN => n57);
   U307 : NAND2_X1 port map( A1 => n1300, A2 => n1299, ZN => n1298);
   U311 : NAND2_X1 port map( A1 => n14101, A2 => n14102, ZN => n14106);
   U312 : INV_X1 port map( A => n7462, ZN => n7461);
   U313 : NAND2_X1 port map( A1 => n8061, A2 => n8060, ZN => n7462);
   U314 : NAND2_X1 port map( A1 => n16662, A2 => n1173, ZN => n60);
   U316 : AOI21_X1 port map( B1 => n4345, B2 => n4344, A => n4516, ZN => n61);
   U318 : AND2_X1 port map( A1 => n19998, A2 => n11500, ZN => n11082);
   U319 : XNOR2_X2 port map( A => n10556, B => n10555, ZN => n11500);
   U321 : NAND2_X1 port map( A1 => n12126, A2 => n1508, ZN => n11703);
   U323 : NAND2_X1 port map( A1 => n2241, A2 => n2242, ZN => n63);
   U324 : AND2_X1 port map( A1 => n11256, A2 => n11253, ZN => n10774);
   U326 : NAND2_X1 port map( A1 => n81, A2 => n16291, ZN => n16497);
   U328 : AND2_X2 port map( A1 => n65, A2 => n64, ZN => n13791);
   U329 : NAND2_X1 port map( A1 => n1439, A2 => n1440, ZN => n64);
   U330 : NAND2_X1 port map( A1 => n12292, A2 => n12291, ZN => n65);
   U334 : NAND2_X1 port map( A1 => n19294, A2 => n20515, ZN => n18166);
   U337 : OAI21_X1 port map( B1 => n18269, B2 => n17766, A => n100, ZN => 
                           n16869);
   U345 : NAND3_X2 port map( A1 => n2543, A2 => n8199, A3 => n1361, ZN => n9217
                           );
   U347 : NAND3_X1 port map( A1 => n15782, A2 => n15686, A3 => n15687, ZN => 
                           n93);
   U351 : NAND2_X1 port map( A1 => n13802, A2 => n14148, ZN => n67);
   U352 : NAND2_X1 port map( A1 => n6035, A2 => n6037, ZN => n86);
   U354 : NAND3_X1 port map( A1 => n2311, A2 => n2005, A3 => n15678, ZN => 
                           n2003);
   U355 : OR2_X2 port map( A1 => n4973, A2 => n4972, ZN => n6036);
   U356 : XNOR2_X1 port map( A => n15218, B => n15219, ZN => n17245);
   U358 : XNOR2_X1 port map( A => n68, B => n7303, ZN => n5759);
   U359 : XNOR2_X1 port map( A => n6942, B => n5754, ZN => n68);
   U360 : XNOR2_X1 port map( A => n6872, B => n106, ZN => n6874);
   U361 : NAND2_X1 port map( A1 => n495, A2 => n497, ZN => n6872);
   U362 : NAND2_X1 port map( A1 => n71, A2 => n70, ZN => n2362);
   U367 : NAND2_X1 port map( A1 => n153, A2 => n4706, ZN => n4453);
   U369 : XNOR2_X1 port map( A => n12681, B => n12682, ZN => n13937);
   U370 : NAND2_X1 port map( A1 => n10688, A2 => n11411, ZN => n11006);
   U375 : OR2_X1 port map( A1 => n8733, A2 => n8736, ZN => n8333);
   U377 : NAND3_X1 port map( A1 => n15507, A2 => n1758, A3 => n15188, ZN => 
                           n14937);
   U383 : NAND2_X1 port map( A1 => n4846, A2 => n4839, ZN => n4661);
   U384 : NAND2_X1 port map( A1 => n164, A2 => n4657, ZN => n4846);
   U386 : AND2_X1 port map( A1 => n11952, A2 => n11598, ZN => n9613);
   U389 : NAND2_X1 port map( A1 => n3873, A2 => n1920, ZN => n5798);
   U390 : NAND3_X1 port map( A1 => n3896, A2 => n74, A3 => n4467, ZN => n3895);
   U391 : NAND2_X1 port map( A1 => n4117, A2 => n4114, ZN => n74);
   U393 : NAND2_X1 port map( A1 => n4916, A2 => n76, ZN => n75);
   U394 : NAND2_X1 port map( A1 => n4952, A2 => n4953, ZN => n76);
   U396 : NAND2_X1 port map( A1 => n4955, A2 => n4954, ZN => n78);
   U401 : AND2_X2 port map( A1 => n10666, A2 => n10665, ZN => n12110);
   U403 : AND2_X2 port map( A1 => n80, A2 => n79, ZN => n10570);
   U404 : NAND2_X1 port map( A1 => n8452, A2 => n19880, ZN => n79);
   U405 : NAND2_X1 port map( A1 => n8453, A2 => n8454, ZN => n80);
   U406 : OR2_X1 port map( A1 => n3948, A2 => n4541, ZN => n4538);
   U407 : BUF_X1 port map( A => n4220, Z => n4845);
   U417 : NAND3_X1 port map( A1 => n626, A2 => n2003, A3 => n625, ZN => n17444)
                           ;
   U419 : AND3_X2 port map( A1 => n1291, A2 => n2715, A3 => n1287, ZN => n16973
                           );
   U424 : NAND3_X1 port map( A1 => n8916, A2 => n19518, A3 => n8917, ZN => 
                           n8918);
   U432 : XNOR2_X2 port map( A => n5854, B => n5853, ZN => n8040);
   U434 : NAND2_X1 port map( A1 => n11469, A2 => n927, ZN => n10884);
   U437 : NAND3_X1 port map( A1 => n3431, A2 => n15607, A3 => n16128, ZN => 
                           n417);
   U443 : NAND2_X1 port map( A1 => n2626, A2 => n19748, ZN => n2439);
   U444 : NAND2_X1 port map( A1 => n1034, A2 => n1033, ZN => n2626);
   U446 : AND2_X2 port map( A1 => n16018, A2 => n16017, ZN => n17347);
   U448 : NAND3_X1 port map( A1 => n8259, A2 => n8159, A3 => n6831, ZN => n6847
                           );
   U452 : NAND2_X1 port map( A1 => n9309, A2 => n1751, ZN => n9229);
   U454 : NAND3_X2 port map( A1 => n8207, A2 => n2885, A3 => n8206, ZN => n9114
                           );
   U457 : NAND2_X1 port map( A1 => n595, A2 => n596, ZN => n594);
   U458 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => n10787);
   U459 : NAND2_X1 port map( A1 => n11879, A2 => n10259, ZN => n83);
   U460 : NAND2_X1 port map( A1 => n10786, A2 => n85, ZN => n84);
   U461 : INV_X1 port map( A => n10259, ZN => n85);
   U462 : NAND2_X1 port map( A1 => n10808, A2 => n11884, ZN => n10786);
   U464 : NAND3_X1 port map( A1 => n15685, A2 => n15779, A3 => n20362, ZN => 
                           n15689);
   U465 : NAND2_X1 port map( A1 => n9338, A2 => n9070, ZN => n8699);
   U469 : BUF_X1 port map( A => n4233, Z => n4499);
   U473 : NAND2_X1 port map( A1 => n86, A2 => n5531, ZN => n1708);
   U474 : XNOR2_X1 port map( A => n13808, B => n12614, ZN => n12626);
   U475 : XNOR2_X1 port map( A => n13376, B => n13518, ZN => n13808);
   U478 : OR2_X2 port map( A1 => n12039, A2 => n11172, ZN => n12282);
   U481 : NAND2_X1 port map( A1 => n3925, A2 => n87, ZN => n4189);
   U483 : NAND2_X1 port map( A1 => n4595, A2 => n4596, ZN => n6477);
   U487 : INV_X1 port map( A => n7961, ZN => n90);
   U488 : INV_X1 port map( A => n7773, ZN => n91);
   U489 : NAND3_X1 port map( A1 => n7961, A2 => n7917, A3 => n1231, ZN => n92);
   U493 : XNOR2_X2 port map( A => Key(145), B => Plaintext(145), ZN => n5010);
   U494 : AOI22_X2 port map( A1 => n9274, A2 => n3618, B1 => n8649, B2 => n8449
                           , ZN => n10114);
   U496 : NAND3_X1 port map( A1 => n94, A2 => n14433, A3 => n2811, ZN => n14488
                           );
   U497 : NAND3_X1 port map( A1 => n14485, A2 => n14486, A3 => n14487, ZN => 
                           n94);
   U498 : NAND2_X1 port map( A1 => n5425, A2 => n5668, ZN => n5674);
   U500 : NOR2_X2 port map( A1 => n14805, A2 => n14804, ZN => n15812);
   U502 : NAND2_X1 port map( A1 => n95, A2 => n11114, ZN => n1813);
   U503 : NOR2_X1 port map( A1 => n1812, A2 => n11452, ZN => n95);
   U511 : NAND2_X1 port map( A1 => n9363, A2 => n8958, ZN => n8965);
   U515 : BUF_X1 port map( A => n10685, Z => n11271);
   U517 : NAND2_X1 port map( A1 => n98, A2 => n8083, ZN => n7558);
   U518 : OAI21_X1 port map( B1 => n8230, B2 => n20107, A => n8085, ZN => n98);
   U519 : NAND2_X1 port map( A1 => n10677, A2 => n11231, ZN => n11235);
   U525 : NAND2_X1 port map( A1 => n18269, A2 => n18275, ZN => n100);
   U528 : NAND2_X1 port map( A1 => n8592, A2 => n9358, ZN => n9530);
   U529 : NAND3_X1 port map( A1 => n647, A2 => n11547, A3 => n258, ZN => n10764
                           );
   U532 : NAND3_X1 port map( A1 => n15831, A2 => n15642, A3 => n2223, ZN => 
                           n15646);
   U534 : NAND2_X1 port map( A1 => n8565, A2 => n8884, ZN => n8471);
   U536 : NAND2_X1 port map( A1 => n443, A2 => n444, ZN => n102);
   U537 : NAND3_X1 port map( A1 => n2600, A2 => n2598, A3 => n12543, ZN => 
                           n11798);
   U551 : OAI211_X1 port map( C1 => n1714, C2 => n1729, A => n103, B => n1727, 
                           ZN => Ciphertext(10));
   U552 : NAND2_X1 port map( A1 => n1714, A2 => n1728, ZN => n103);
   U553 : OR2_X1 port map( A1 => n11717, A2 => n12279, ZN => n12278);
   U558 : NAND2_X1 port map( A1 => n15600, A2 => n15275, ZN => n15277);
   U560 : AOI21_X1 port map( B1 => n11447, B2 => n11448, A => n11446, ZN => 
                           n104);
   U565 : NAND2_X1 port map( A1 => n19375, A2 => n19380, ZN => n17236);
   U566 : NAND2_X2 port map( A1 => n435, A2 => n15570, ZN => n17014);
   U569 : NAND2_X1 port map( A1 => n14809, A2 => n14813, ZN => n107);
   U570 : NAND2_X1 port map( A1 => n474, A2 => n239, ZN => n108);
   U571 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => n8491);
   U572 : NAND2_X1 port map( A1 => n8940, A2 => n8644, ZN => n8946);
   U573 : NAND2_X1 port map( A1 => n8489, A2 => n111, ZN => n110);
   U574 : INV_X1 port map( A => n8947, ZN => n111);
   U575 : BUF_X1 port map( A => n16639, Z => n17219);
   U577 : OAI21_X2 port map( B1 => n11301, B2 => n11398, A => n11300, ZN => 
                           n12399);
   U578 : OAI211_X2 port map( C1 => n17450, C2 => n17946, A => n2290, B => 
                           n2289, ZN => n18697);
   U581 : NAND3_X1 port map( A1 => n12335, A2 => n12339, A3 => n11992, ZN => 
                           n11971);
   U582 : XNOR2_X1 port map( A => n13600, B => n112, ZN => n13257);
   U583 : INV_X1 port map( A => n13255, ZN => n112);
   U587 : NAND2_X1 port map( A1 => n5630, A2 => n5631, ZN => n5634);
   U588 : INV_X1 port map( A => n17882, ZN => n113);
   U589 : NOR2_X1 port map( A1 => n5635, A2 => n5636, ZN => n6301);
   U593 : NAND2_X1 port map( A1 => n20258, A2 => n18238, ZN => n114);
   U594 : OR3_X1 port map( A1 => n15081, A2 => n15422, A3 => n15531, ZN => 
                           n14257);
   U595 : XNOR2_X1 port map( A => n6667, B => n6666, ZN => n6671);
   U597 : INV_X1 port map( A => n5752, ZN => n5750);
   U598 : NAND2_X1 port map( A1 => n5744, A2 => n5743, ZN => n5752);
   U603 : NAND2_X1 port map( A1 => n12488, A2 => n12811, ZN => n11693);
   U606 : OR2_X1 port map( A1 => n11283, A2 => n10693, ZN => n11286);
   U607 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => n5649);
   U608 : NAND2_X1 port map( A1 => n4172, A2 => n4171, ZN => n118);
   U612 : NAND3_X1 port map( A1 => n11185, A2 => n2948, A3 => n2949, ZN => 
                           n12141);
   U613 : NAND2_X1 port map( A1 => n8126, A2 => n9453, ZN => n8127);
   U616 : NAND2_X1 port map( A1 => n8597, A2 => n8928, ZN => n8598);
   U618 : OAI22_X1 port map( A1 => n17396, A2 => n18264, B1 => n17762, B2 => 
                           n18750, ZN => n17397);
   U619 : AOI22_X2 port map( A1 => n1223, A2 => n228, B1 => n15815, B2 => 
                           n15036, ZN => n17358);
   U620 : OAI211_X1 port map( C1 => n11439, C2 => n11116, A => n11034, B => 
                           n119, ZN => n3160);
   U621 : OR2_X1 port map( A1 => n11115, A2 => n11440, ZN => n119);
   U631 : NAND2_X1 port map( A1 => n122, A2 => n11990, ZN => n121);
   U632 : OR2_X2 port map( A1 => n775, A2 => n3901, ZN => n5428);
   U634 : NAND2_X2 port map( A1 => n3998, A2 => n3997, ZN => n6067);
   U635 : NAND2_X1 port map( A1 => n201, A2 => n12500, ZN => n2016);
   U636 : AND2_X2 port map( A1 => n3981, A2 => n3320, ZN => n3319);
   U638 : OR2_X1 port map( A1 => n14796, A2 => n13891, ZN => n14213);
   U642 : MUX2_X2 port map( A => n14383, B => n14382, S => n14381, Z => n15838)
                           ;
   U643 : NAND2_X1 port map( A1 => n8768, A2 => n8477, ZN => n1470);
   U644 : NAND2_X1 port map( A1 => n1672, A2 => n1671, ZN => n8768);
   U646 : XNOR2_X2 port map( A => n12496, B => n12495, ZN => n14789);
   U648 : NAND2_X1 port map( A1 => n12759, A2 => n123, ZN => n1828);
   U649 : NOR2_X1 port map( A1 => n2523, A2 => n12754, ZN => n123);
   U651 : NAND2_X1 port map( A1 => n4555, A2 => n20229, ZN => n4731);
   U654 : NAND2_X1 port map( A1 => n2056, A2 => n12595, ZN => n125);
   U655 : XNOR2_X2 port map( A => n2264, B => n11682, ZN => n14813);
   U659 : OAI21_X1 port map( B1 => n12008, B2 => n12009, A => n126, ZN => 
                           n11662);
   U664 : AND2_X1 port map( A1 => n11539, A2 => n11168, ZN => n11537);
   U666 : OR2_X1 port map( A1 => n18697, A2 => n18702, ZN => n18706);
   U667 : NAND2_X1 port map( A1 => n12412, A2 => n12390, ZN => n3082);
   U668 : NAND2_X1 port map( A1 => n128, A2 => n4206, ZN => n4209);
   U669 : NAND2_X1 port map( A1 => n5003, A2 => n4750, ZN => n128);
   U670 : NAND2_X1 port map( A1 => n20168, A2 => n17501, ZN => n17503);
   U671 : BUF_X2 port map( A => n5250, Z => n5323);
   U673 : NAND2_X1 port map( A1 => n1976, A2 => n1977, ZN => n129);
   U678 : NAND2_X1 port map( A1 => n3734, A2 => n12261, ZN => n1045);
   U686 : AND3_X2 port map( A1 => n7555, A2 => n7554, A3 => n7553, ZN => n8961)
                           ;
   U695 : OAI211_X2 port map( C1 => n10944, C2 => n12048, A => n10942, B => 
                           n130, ZN => n13058);
   U696 : NAND3_X1 port map( A1 => n10944, A2 => n10934, A3 => n11647, ZN => 
                           n130);
   U697 : NAND3_X1 port map( A1 => n1213, A2 => n12337, A3 => n12338, ZN => 
                           n12342);
   U698 : NAND2_X1 port map( A1 => n4108, A2 => n567, ZN => n3290);
   U703 : AND2_X2 port map( A1 => n14391, A2 => n1021, ZN => n1288);
   U704 : NAND3_X1 port map( A1 => n8892, A2 => n8893, A3 => n9010, ZN => n8894
                           );
   U706 : OR2_X2 port map( A1 => n13926, A2 => n13925, ZN => n14935);
   U709 : NAND2_X1 port map( A1 => n11926, A2 => n11683, ZN => n12579);
   U710 : NAND3_X2 port map( A1 => n11004, A2 => n411, A3 => n11003, ZN => 
                           n11926);
   U712 : NAND3_X1 port map( A1 => n1266, A2 => n1265, A3 => n15314, ZN => 
                           n1129);
   U713 : OAI21_X2 port map( B1 => n15383, B2 => n3621, A => n2862, ZN => 
                           n16840);
   U714 : MUX2_X2 port map( A => n14030, B => n14029, S => n20120, Z => n15491)
                           ;
   U715 : NOR2_X1 port map( A1 => n5251, A2 => n5323, ZN => n5392);
   U719 : NAND2_X2 port map( A1 => n10470, A2 => n10471, ZN => n11995);
   U726 : XNOR2_X2 port map( A => n4040, B => Key(120), ZN => n4708);
   U729 : NAND2_X1 port map( A1 => n17670, A2 => n19360, ZN => n131);
   U732 : NAND3_X2 port map( A1 => n14144, A2 => n14145, A3 => n133, ZN => 
                           n15509);
   U733 : OR2_X2 port map( A1 => n14774, A2 => n14773, ZN => n16964);
   U735 : OAI21_X1 port map( B1 => n6041, B2 => n135, A => n134, ZN => n5889);
   U736 : NAND2_X1 port map( A1 => n6041, A2 => n1214, ZN => n134);
   U741 : XNOR2_X1 port map( A => n137, B => n1259, ZN => Ciphertext(171));
   U744 : NAND2_X2 port map( A1 => n9270, A2 => n1157, ZN => n10360);
   U752 : NAND2_X1 port map( A1 => n2596, A2 => n4137, ZN => n4139);
   U755 : NAND3_X1 port map( A1 => n2773, A2 => n140, A3 => n139, ZN => n564);
   U759 : OAI211_X1 port map( C1 => n19090, C2 => n19089, A => n141, B => 
                           n19088, ZN => n19091);
   U760 : NAND2_X1 port map( A1 => n19086, A2 => n19109, ZN => n141);
   U766 : BUF_X1 port map( A => n14952, Z => n15803);
   U767 : OAI211_X1 port map( C1 => n143, C2 => n3515, A => n142, B => n11142, 
                           ZN => n1669);
   U768 : NAND2_X1 port map( A1 => n273, A2 => n8014, ZN => n7992);
   U769 : AOI21_X2 port map( B1 => n144, B2 => n307, A => n1000, ZN => n16961);
   U770 : NOR2_X1 port map( A1 => n14983, A2 => n15522, ZN => n144);
   U774 : NOR2_X1 port map( A1 => n8879, A2 => n9249, ZN => n1618);
   U779 : OR2_X1 port map( A1 => n6090, A2 => n5176, ZN => n806);
   U780 : OR2_X1 port map( A1 => n6090, A2 => n6087, ZN => n1468);
   U782 : OR3_X1 port map( A1 => n5997, A2 => n5434, A3 => n5704, ZN => n5814);
   U783 : OR2_X1 port map( A1 => n19980, A2 => n6007, ZN => n6014);
   U784 : INV_X1 port map( A => n7421, ZN => n585);
   U786 : OR2_X1 port map( A1 => n20257, A2 => n5941, ZN => n1834);
   U787 : AND2_X1 port map( A1 => n8542, A2 => n9065, ZN => n8544);
   U789 : INV_X1 port map( A => n2749, ZN => n545);
   U790 : XNOR2_X1 port map( A => n694, B => n10027, ZN => n10319);
   U792 : NOR2_X1 port map( A1 => n15495, A2 => n747, ZN => n3425);
   U793 : OAI21_X1 port map( B1 => n15574, B2 => n15365, A => n15796, ZN => 
                           n15366);
   U794 : OAI21_X1 port map( B1 => n18094, B2 => n19774, A => n424, ZN => 
                           n17166);
   U795 : AND2_X1 port map( A1 => n19935, A2 => n18650, ZN => n18645);
   U796 : OR2_X1 port map( A1 => n19456, A2 => n19459, ZN => n810);
   U797 : AND2_X1 port map( A1 => n5955, A2 => n6107, ZN => n145);
   U798 : AND2_X1 port map( A1 => n5780, A2 => n5778, ZN => n146);
   U799 : AND2_X2 port map( A1 => n7636, A2 => n1404, ZN => n8602);
   U800 : NAND4_X2 port map( A1 => n7107, A2 => n7104, A3 => n7105, A4 => n7106
                           , ZN => n8851);
   U803 : AND2_X1 port map( A1 => n951, A2 => n20443, ZN => n147);
   U805 : NAND2_X2 port map( A1 => n2152, A2 => n2153, ZN => n15573);
   U806 : OR2_X1 port map( A1 => n14916, A2 => n15863, ZN => n148);
   U807 : NAND2_X2 port map( A1 => n12933, A2 => n2535, ZN => n15380);
   U808 : OR2_X1 port map( A1 => n15093, A2 => n15636, ZN => n149);
   U810 : OR2_X1 port map( A1 => n19708, A2 => n19163, ZN => n150);
   U812 : OR2_X1 port map( A1 => n19031, A2 => n20074, ZN => n151);
   U813 : AND3_X1 port map( A1 => n19775, A2 => n16453, A3 => n16452, ZN => 
                           n152);
   U821 : XNOR2_X1 port map( A => Key(122), B => Plaintext(122), ZN => n5031);
   U830 : XNOR2_X1 port map( A => Key(177), B => Plaintext(177), ZN => n4638);
   U842 : MUX2_X2 port map( A => n8346, B => n8345, S => n8344, Z => n9135);
   U846 : XNOR2_X2 port map( A => n6893, B => n6892, ZN => n8347);
   U856 : XNOR2_X1 port map( A => Key(69), B => Plaintext(69), ZN => n4656);
   U858 : XNOR2_X2 port map( A => Key(162), B => Plaintext(162), ZN => n4539);
   U867 : OAI21_X2 port map( B1 => n5210, B2 => n861, A => n5209, ZN => n6854);
   U872 : INV_X2 port map( A => n5106, ZN => n5102);
   U874 : AND2_X2 port map( A1 => n1131, A2 => n1393, ZN => n7345);
   U879 : AND2_X2 port map( A1 => n1445, A2 => n4900, ZN => n5682);
   U888 : XNOR2_X2 port map( A => n13140, B => n13471, ZN => n14667);
   U894 : XNOR2_X2 port map( A => Key(87), B => Plaintext(87), ZN => n5073);
   U901 : XNOR2_X2 port map( A => n13170, B => n13171, ZN => n14666);
   U905 : OAI21_X2 port map( B1 => n3193, B2 => n12878, A => n12881, ZN => 
                           n15167);
   U911 : AOI22_X1 port map( A1 => n4655, A2 => n4654, B1 => n4863, B2 => n4653
                           , ZN => n6167);
   U932 : XNOR2_X1 port map( A => n6885, B => n6884, ZN => n8349);
   U934 : BUF_X1 port map( A => n4686, Z => n177);
   U935 : BUF_X1 port map( A => n4686, Z => n178);
   U936 : XNOR2_X1 port map( A => Key(57), B => Plaintext(57), ZN => n4686);
   U937 : OAI21_X2 port map( B1 => n5708, B2 => n4113, A => n622, ZN => n7390);
   U950 : OR2_X1 port map( A1 => n7967, A2 => n278, ZN => n7976);
   U951 : XNOR2_X2 port map( A => n3953, B => Key(187), ZN => n4614);
   U952 : NAND2_X2 port map( A1 => n6197, A2 => n6198, ZN => n7031);
   U954 : NAND2_X2 port map( A1 => n1983, A2 => n1982, ZN => n7134);
   U956 : AOI22_X2 port map( A1 => n17980, A2 => n18752, B1 => n17979, B2 => 
                           n17978, ZN => n18682);
   U960 : OAI21_X2 port map( B1 => n8575, B2 => n9059, A => n8574, ZN => n10186
                           );
   U962 : AOI21_X2 port map( B1 => n8643, B2 => n8642, A => n8641, ZN => n10240
                           );
   U963 : XNOR2_X2 port map( A => n3880, B => Key(0), ZN => n4169);
   U975 : XNOR2_X2 port map( A => n2745, B => n2744, ZN => n10677);
   U977 : OAI22_X2 port map( A1 => n11969, A2 => n11631, B1 => n11629, B2 => 
                           n11630, ZN => n12986);
   U978 : OAI21_X2 port map( B1 => n6074, B2 => n6075, A => n6073, ZN => n7391)
                           ;
   U984 : BUF_X1 port map( A => n11325, Z => n190);
   U987 : NOR2_X1 port map( A1 => n18454, A2 => n20139, ZN => n18469);
   U989 : OAI21_X1 port map( B1 => n17679, B2 => n20514, A => n17678, ZN => 
                           n1205);
   U991 : OAI21_X1 port map( B1 => n222, B2 => n17876, A => n600, ZN => n19248)
                           ;
   U993 : OR2_X1 port map( A1 => n14838, A2 => n15018, ZN => n322);
   U994 : INV_X1 port map( A => n16011, ZN => n192);
   U1002 : INV_X1 port map( A => n12589, ZN => n193);
   U1005 : CLKBUF_X1 port map( A => n10684, Z => n12104);
   U1006 : NAND2_X1 port map( A1 => n7284, A2 => n3210, ZN => n8932);
   U1009 : NAND3_X1 port map( A1 => n8151, A2 => n7864, A3 => n8261, ZN => 
                           n7572);
   U1010 : NAND2_X1 port map( A1 => n8175, A2 => n8179, ZN => n7887);
   U1012 : CLKBUF_X1 port map( A => n7508, Z => n7910);
   U1014 : NAND4_X1 port map( A1 => n5353, A2 => n5352, A3 => n5351, A4 => 
                           n5350, ZN => n7146);
   U1017 : CLKBUF_X1 port map( A => n4176, Z => n4613);
   U1019 : CLKBUF_X1 port map( A => Key(14), Z => n16035);
   U1020 : CLKBUF_X1 port map( A => Key(118), Z => n2329);
   U1021 : CLKBUF_X1 port map( A => Key(104), Z => n2454);
   U1022 : CLKBUF_X1 port map( A => Key(147), Z => n2344);
   U1023 : CLKBUF_X1 port map( A => Key(141), Z => n2446);
   U1024 : CLKBUF_X1 port map( A => Key(128), Z => n2096);
   U1025 : CLKBUF_X1 port map( A => Key(45), Z => n17365);
   U1027 : CLKBUF_X1 port map( A => Key(32), Z => n1857);
   U1028 : CLKBUF_X1 port map( A => Key(68), Z => n18478);
   U1029 : CLKBUF_X1 port map( A => Key(29), Z => n18801);
   U1031 : CLKBUF_X1 port map( A => Key(157), Z => n1969);
   U1032 : CLKBUF_X1 port map( A => Key(145), Z => n2082);
   U1033 : CLKBUF_X1 port map( A => Key(101), Z => n18420);
   U1034 : CLKBUF_X1 port map( A => Key(67), Z => n18170);
   U1035 : CLKBUF_X1 port map( A => Key(171), Z => n17733);
   U1036 : AOI21_X1 port map( B1 => n19267, B2 => n19276, A => n658, ZN => 
                           n19279);
   U1038 : NAND2_X1 port map( A1 => n1557, A2 => n1556, ZN => n19146);
   U1043 : MUX2_X1 port map( A => n16043, B => n16042, S => n19707, Z => n19168
                           );
   U1044 : INV_X1 port map( A => n19164, ZN => n195);
   U1045 : AND2_X1 port map( A1 => n3039, A2 => n17906, ZN => n18358);
   U1046 : OAI211_X1 port map( C1 => n220, C2 => n20127, A => n17193, B => n326
                           , ZN => n17820);
   U1047 : CLKBUF_X1 port map( A => n17225, Z => n17510);
   U1048 : CLKBUF_X1 port map( A => n16251, Z => n16629);
   U1049 : CLKBUF_X1 port map( A => n17394, Z => n18754);
   U1050 : INV_X1 port map( A => n17676, ZN => n1112);
   U1051 : XNOR2_X1 port map( A => n16935, B => n16934, ZN => n18948);
   U1055 : BUF_X1 port map( A => n16171, Z => n17507);
   U1057 : XNOR2_X1 port map( A => n16433, B => n16432, ZN => n18092);
   U1058 : INV_X1 port map( A => n17876, ZN => n196);
   U1061 : XNOR2_X1 port map( A => n15979, B => n17143, ZN => n16553);
   U1065 : INV_X1 port map( A => n15310, ZN => n197);
   U1066 : INV_X1 port map( A => n15714, ZN => n198);
   U1067 : INV_X1 port map( A => n14707, ZN => n14273);
   U1068 : INV_X1 port map( A => n14547, ZN => n199);
   U1069 : AND2_X1 port map( A1 => n14562, A2 => n14566, ZN => n14708);
   U1072 : INV_X1 port map( A => n14692, ZN => n200);
   U1074 : XNOR2_X1 port map( A => n11789, B => n11788, ZN => n14199);
   U1076 : XNOR2_X1 port map( A => n12173, B => n294, ZN => n13636);
   U1077 : XNOR2_X1 port map( A => n12173, B => n299, ZN => n12850);
   U1078 : XNOR2_X1 port map( A => n12173, B => n304, ZN => n13049);
   U1082 : AND3_X1 port map( A1 => n12164, A2 => n3476, A3 => n12163, ZN => 
                           n12173);
   U1084 : OR2_X1 port map( A1 => n1252, A2 => n193, ZN => n1251);
   U1085 : INV_X1 port map( A => n248, ZN => n685);
   U1086 : CLKBUF_X1 port map( A => n12275, Z => n920);
   U1093 : NAND3_X1 port map( A1 => n10847, A2 => n11202, A3 => n19920, ZN => 
                           n10848);
   U1094 : AND3_X1 port map( A1 => n11177, A2 => n11174, A3 => n9486, ZN => 
                           n3219);
   U1095 : INV_X1 port map( A => n11330, ZN => n202);
   U1096 : CLKBUF_X1 port map( A => n9548, Z => n10952);
   U1098 : CLKBUF_X1 port map( A => n9351, Z => n9486);
   U1099 : INV_X1 port map( A => n11216, ZN => n204);
   U1100 : XNOR2_X1 port map( A => n9409, B => n9410, ZN => n10947);
   U1101 : INV_X1 port map( A => n11129, ZN => n205);
   U1102 : XNOR2_X1 port map( A => n10030, B => n298, ZN => n9404);
   U1103 : XNOR2_X1 port map( A => n9646, B => n296, ZN => n8716);
   U1104 : XNOR2_X1 port map( A => n260, B => n9646, ZN => n9910);
   U1105 : XNOR2_X1 port map( A => n10030, B => n300, ZN => n9417);
   U1107 : NOR2_X1 port map( A1 => n8847, A2 => n3201, ZN => n9623);
   U1113 : INV_X1 port map( A => n8959, ZN => n207);
   U1115 : OR2_X1 port map( A1 => n1231, A2 => n277, ZN => n377);
   U1117 : CLKBUF_X1 port map( A => n6734, Z => n8373);
   U1119 : INV_X1 port map( A => n8016, ZN => n208);
   U1120 : XNOR2_X1 port map( A => n1369, B => n6630, ZN => n8068);
   U1121 : XNOR2_X1 port map( A => n3570, B => n3572, ZN => n7479);
   U1122 : XNOR2_X1 port map( A => n5249, B => n295, ZN => n6386);
   U1123 : XNOR2_X1 port map( A => n5249, B => n293, ZN => n6620);
   U1125 : OR2_X1 port map( A1 => n5947, A2 => n5946, ZN => n7127);
   U1126 : NAND3_X1 port map( A1 => n5187, A2 => n2978, A3 => n5186, ZN => 
                           n7178);
   U1127 : AND2_X1 port map( A1 => n355, A2 => n5848, ZN => n354);
   U1129 : OAI211_X1 port map( C1 => n5943, C2 => n6172, A => n6175, B => n5221
                           , ZN => n6873);
   U1131 : OR2_X1 port map( A1 => n5816, A2 => n285, ZN => n5820);
   U1132 : NAND2_X1 port map( A1 => n827, A2 => n830, ZN => n5435);
   U1133 : NOR3_X1 port map( A1 => n6166, A2 => n170, A3 => n6171, ZN => n569);
   U1135 : AND2_X1 port map( A1 => n762, A2 => n3714, ZN => n5747);
   U1137 : INV_X1 port map( A => n6067, ZN => n209);
   U1139 : OR2_X1 port map( A1 => n5079, A2 => n20002, ZN => n4809);
   U1141 : INV_X1 port map( A => n4899, ZN => n210);
   U1142 : CLKBUF_X1 port map( A => Key(85), Z => n18848);
   U1143 : CLKBUF_X1 port map( A => Key(46), Z => n632);
   U1144 : CLKBUF_X1 port map( A => Key(83), Z => n19336);
   U1146 : CLKBUF_X1 port map( A => Key(163), Z => n2347);
   U1147 : CLKBUF_X1 port map( A => Key(34), Z => n2376);
   U1148 : CLKBUF_X1 port map( A => Key(133), Z => n17170);
   U1150 : CLKBUF_X1 port map( A => Key(25), Z => n2218);
   U1151 : CLKBUF_X1 port map( A => Key(21), Z => n2375);
   U1152 : CLKBUF_X1 port map( A => Key(8), Z => n2298);
   U1153 : CLKBUF_X1 port map( A => Key(191), Z => n2123);
   U1154 : CLKBUF_X1 port map( A => Key(170), Z => n2284);
   U1155 : CLKBUF_X1 port map( A => Key(44), Z => n484);
   U1156 : CLKBUF_X1 port map( A => Key(18), Z => n19216);
   U1157 : CLKBUF_X1 port map( A => Key(96), Z => n2369);
   U1158 : CLKBUF_X1 port map( A => Key(58), Z => n1148);
   U1159 : CLKBUF_X1 port map( A => Key(182), Z => n1904);
   U1160 : CLKBUF_X1 port map( A => Key(90), Z => n18779);
   U1161 : CLKBUF_X1 port map( A => Key(11), Z => n2087);
   U1162 : CLKBUF_X1 port map( A => Key(111), Z => n16030);
   U1163 : CLKBUF_X1 port map( A => Key(168), Z => n2257);
   U1164 : CLKBUF_X1 port map( A => Key(15), Z => n16424);
   U1165 : CLKBUF_X1 port map( A => Key(161), Z => n2392);
   U1166 : CLKBUF_X1 port map( A => Key(125), Z => n19436);
   U1167 : CLKBUF_X1 port map( A => Key(89), Z => n1386);
   U1168 : CLKBUF_X1 port map( A => Key(86), Z => n2248);
   U1169 : CLKBUF_X1 port map( A => Key(0), Z => n2341);
   U1170 : CLKBUF_X1 port map( A => Key(64), Z => n457);
   U1171 : CLKBUF_X1 port map( A => Key(4), Z => n1996);
   U1172 : CLKBUF_X1 port map( A => Key(91), Z => n18006);
   U1173 : CLKBUF_X1 port map( A => Key(72), Z => n2122);
   U1174 : CLKBUF_X1 port map( A => Key(87), Z => n311);
   U1175 : CLKBUF_X1 port map( A => Key(116), Z => n16366);
   U1176 : CLKBUF_X1 port map( A => Key(150), Z => n642);
   U1177 : CLKBUF_X1 port map( A => Key(143), Z => n2448);
   U1178 : CLKBUF_X1 port map( A => Key(172), Z => n2323);
   U1179 : CLKBUF_X1 port map( A => Key(106), Z => n621);
   U1180 : CLKBUF_X1 port map( A => Key(37), Z => n2368);
   U1181 : CLKBUF_X1 port map( A => Key(130), Z => n573);
   U1182 : CLKBUF_X1 port map( A => Key(140), Z => n18090);
   U1183 : CLKBUF_X1 port map( A => Key(23), Z => n2410);
   U1184 : CLKBUF_X1 port map( A => Key(153), Z => n18070);
   U1185 : CLKBUF_X1 port map( A => Key(27), Z => n2395);
   U1186 : CLKBUF_X1 port map( A => Key(5), Z => n19018);
   U1187 : CLKBUF_X1 port map( A => Key(26), Z => n18433);
   U1188 : CLKBUF_X1 port map( A => Key(126), Z => n875);
   U1190 : CLKBUF_X1 port map( A => Key(71), Z => n18830);
   U1191 : CLKBUF_X1 port map( A => Key(92), Z => n15479);
   U1193 : CLKBUF_X1 port map( A => Key(40), Z => n347);
   U1194 : CLKBUF_X1 port map( A => Key(19), Z => n18208);
   U1195 : CLKBUF_X1 port map( A => Key(70), Z => n2067);
   U1197 : CLKBUF_X1 port map( A => Key(112), Z => n18304);
   U1198 : CLKBUF_X1 port map( A => Key(149), Z => n19243);
   U1200 : CLKBUF_X1 port map( A => Key(49), Z => n17587);
   U1201 : CLKBUF_X1 port map( A => Key(178), Z => n1869);
   U1202 : CLKBUF_X1 port map( A => Key(151), Z => n18716);
   U1203 : CLKBUF_X1 port map( A => Key(12), Z => n2280);
   U1204 : CLKBUF_X1 port map( A => Key(154), Z => n2424);
   U1205 : CLKBUF_X1 port map( A => Key(20), Z => n2222);
   U1206 : CLKBUF_X1 port map( A => Key(158), Z => n19321);
   U1207 : CLKBUF_X1 port map( A => Key(109), Z => n17466);
   U1208 : CLKBUF_X1 port map( A => Key(74), Z => n2356);
   U1209 : CLKBUF_X1 port map( A => Key(80), Z => n18988);
   U1210 : CLKBUF_X1 port map( A => Key(2), Z => n18203);
   U1211 : CLKBUF_X1 port map( A => Key(131), Z => n2385);
   U1212 : CLKBUF_X1 port map( A => Key(105), Z => n2208);
   U1213 : CLKBUF_X1 port map( A => Key(138), Z => n538);
   U1214 : CLKBUF_X1 port map( A => Key(152), Z => n2233);
   U1216 : CLKBUF_X1 port map( A => Key(166), Z => n2337);
   U1217 : CLKBUF_X1 port map( A => Key(134), Z => n641);
   U1218 : CLKBUF_X1 port map( A => Key(107), Z => n19205);
   U1219 : CLKBUF_X1 port map( A => Key(61), Z => n610);
   U1220 : CLKBUF_X1 port map( A => Key(115), Z => n16487);
   U1221 : CLKBUF_X1 port map( A => Key(135), Z => n19222);
   U1222 : CLKBUF_X1 port map( A => Key(77), Z => n17932);
   U1225 : CLKBUF_X1 port map( A => Key(122), Z => n18065);
   U1226 : CLKBUF_X1 port map( A => Key(16), Z => n404);
   U1227 : CLKBUF_X1 port map( A => Key(102), Z => n16242);
   U1228 : CLKBUF_X1 port map( A => Key(9), Z => n17089);
   U1229 : CLKBUF_X1 port map( A => Key(55), Z => n2310);
   U1230 : CLKBUF_X1 port map( A => Key(56), Z => n18338);
   U1231 : CLKBUF_X1 port map( A => Key(113), Z => n18863);
   U1232 : CLKBUF_X1 port map( A => Key(78), Z => n19467);
   U1233 : CLKBUF_X1 port map( A => Key(129), Z => n18439);
   U1235 : CLKBUF_X1 port map( A => Key(48), Z => n17804);
   U1236 : CLKBUF_X1 port map( A => Key(121), Z => n2296);
   U1237 : CLKBUF_X1 port map( A => Key(187), Z => n19158);
   U1238 : CLKBUF_X1 port map( A => Key(24), Z => n2164);
   U1239 : CLKBUF_X1 port map( A => Key(110), Z => n2307);
   U1240 : CLKBUF_X1 port map( A => Key(38), Z => n18887);
   U1241 : CLKBUF_X1 port map( A => Key(52), Z => n2203);
   U1242 : CLKBUF_X1 port map( A => Key(84), Z => n649);
   U1243 : CLKBUF_X1 port map( A => Key(76), Z => n18768);
   U1244 : CLKBUF_X1 port map( A => Key(169), Z => n18984);
   U1245 : CLKBUF_X1 port map( A => Key(148), Z => n2305);
   U1246 : CLKBUF_X1 port map( A => Key(114), Z => n2221);
   U1248 : CLKBUF_X1 port map( A => Key(47), Z => n19052);
   U1249 : CLKBUF_X1 port map( A => Key(73), Z => n2394);
   U1250 : CLKBUF_X1 port map( A => Key(17), Z => n18366);
   U1251 : CLKBUF_X1 port map( A => Key(62), Z => n18726);
   U1252 : CLKBUF_X1 port map( A => Key(127), Z => n2151);
   U1253 : CLKBUF_X1 port map( A => Key(188), Z => n18854);
   U1254 : CLKBUF_X1 port map( A => Key(146), Z => n17993);
   U1255 : CLKBUF_X1 port map( A => Key(155), Z => n17060);
   U1256 : CLKBUF_X1 port map( A => Key(10), Z => n18055);
   U1257 : CLKBUF_X1 port map( A => Key(181), Z => n2032);
   U1258 : CLKBUF_X1 port map( A => Key(162), Z => n18396);
   U1259 : CLKBUF_X1 port map( A => Key(120), Z => n16651);
   U1261 : CLKBUF_X1 port map( A => Key(43), Z => n2055);
   U1262 : CLKBUF_X1 port map( A => Key(66), Z => n2442);
   U1263 : CLKBUF_X1 port map( A => Key(31), Z => n2413);
   U1264 : CLKBUF_X1 port map( A => Key(35), Z => n18011);
   U1265 : CLKBUF_X1 port map( A => Key(3), Z => n2192);
   U1267 : INV_X1 port map( A => n19125, ZN => n833);
   U1269 : MUX2_X1 port map( A => n17088, B => n17087, S => n19683, Z => n17090
                           );
   U1270 : OAI21_X1 port map( B1 => n18201, B2 => n16446, A => n2208, ZN => 
                           n628);
   U1271 : OR2_X1 port map( A1 => n17997, A2 => n18555, ZN => n16459);
   U1272 : AND2_X1 port map( A1 => n18646, A2 => n299, ZN => n842);
   U1274 : OAI22_X1 port map( A1 => n19692, A2 => n19163, B1 => n19948, B2 => 
                           n18306, ZN => n19166);
   U1275 : CLKBUF_X1 port map( A => n18311, Z => n19334);
   U1277 : NOR2_X1 port map( A1 => n18465, A2 => n20110, ZN => n18441);
   U1278 : OR2_X1 port map( A1 => n18638, A2 => n18637, ZN => n583);
   U1283 : AND2_X1 port map( A1 => n930, A2 => n931, ZN => n19460);
   U1284 : INV_X1 port map( A => n18009, ZN => n18504);
   U1285 : AND2_X1 port map( A1 => n19009, A2 => n19002, ZN => n310);
   U1287 : AND3_X1 port map( A1 => n16405, A2 => n1147, A3 => n1146, ZN => 
                           n18559);
   U1288 : INV_X1 port map( A => n19190, ZN => n19197);
   U1292 : INV_X1 port map( A => n19452, ZN => n212);
   U1293 : INV_X1 port map( A => n18795, ZN => n213);
   U1297 : AND3_X1 port map( A1 => n1906, A2 => n1905, A3 => n982, ZN => n19233
                           );
   U1298 : INV_X1 port map( A => n18511, ZN => n214);
   U1306 : OAI21_X1 port map( B1 => n18268, B2 => n16869, A => n16868, ZN => 
                           n17054);
   U1308 : MUX2_X1 port map( A => n17151, B => n17150, S => n17957, Z => n17152
                           );
   U1309 : OAI21_X1 port map( B1 => n612, B2 => n18262, A => n611, ZN => n17398
                           );
   U1311 : INV_X1 port map( A => n1205, ZN => n215);
   U1312 : NOR2_X1 port map( A1 => n17164, A2 => n759, ZN => n17165);
   U1313 : OR2_X1 port map( A1 => n17864, A2 => n17595, ZN => n601);
   U1314 : OR2_X1 port map( A1 => n17762, A2 => n18264, ZN => n18140);
   U1316 : OAI211_X1 port map( C1 => n17161, C2 => n16792, A => n16791, B => 
                           n18542, ZN => n17584);
   U1317 : INV_X1 port map( A => n18869, ZN => n216);
   U1318 : OR2_X1 port map( A1 => n196, A2 => n17879, ZN => n17610);
   U1319 : NOR2_X1 port map( A1 => n17495, A2 => n17492, ZN => n17490);
   U1320 : INV_X1 port map( A => n17492, ZN => n16801);
   U1321 : CLKBUF_X1 port map( A => n17458, Z => n17559);
   U1322 : OR2_X1 port map( A1 => n19846, A2 => n18948, ZN => n17315);
   U1324 : MUX2_X1 port map( A => n17830, B => n17829, S => n20221, Z => n17834
                           );
   U1332 : AND2_X1 port map( A1 => n18221, A2 => n18977, ZN => n18224);
   U1334 : INV_X1 port map( A => n18956, ZN => n219);
   U1335 : OR2_X1 port map( A1 => n18273, A2 => n18033, ZN => n17764);
   U1337 : INV_X1 port map( A => n19380, ZN => n635);
   U1338 : XNOR2_X1 port map( A => n16060, B => n16061, ZN => n17879);
   U1339 : AOI21_X1 port map( B1 => n18221, B2 => n20499, A => n18976, ZN => 
                           n320);
   U1340 : BUF_X1 port map( A => n17187, Z => n18935);
   U1341 : INV_X1 port map( A => n17245, ZN => n812);
   U1342 : XNOR2_X1 port map( A => n16520, B => n16519, ZN => n17861);
   U1344 : BUF_X1 port map( A => n16540, Z => n19348);
   U1345 : INV_X1 port map( A => n18968, ZN => n220);
   U1348 : INV_X1 port map( A => n18273, ZN => n221);
   U1350 : XNOR2_X1 port map( A => n15949, B => n15950, ZN => n17825);
   U1351 : INV_X1 port map( A => n19823, ZN => n815);
   U1354 : INV_X1 port map( A => n17881, ZN => n222);
   U1356 : XNOR2_X1 port map( A => n16904, B => n16903, ZN => n18976);
   U1359 : INV_X1 port map( A => n18221, ZN => n224);
   U1360 : INV_X1 port map( A => n20499, ZN => n225);
   U1362 : XNOR2_X1 port map( A => n16585, B => n16586, ZN => n19396);
   U1363 : INV_X1 port map( A => n18092, ZN => n226);
   U1364 : XNOR2_X1 port map( A => n15557, B => n15556, ZN => n16666);
   U1365 : INV_X1 port map( A => n17818, ZN => n227);
   U1366 : XNOR2_X1 port map( A => n17102, B => n334, ZN => n16132);
   U1367 : INV_X1 port map( A => n15979, ZN => n17005);
   U1369 : AND3_X1 port map( A1 => n15035, A2 => n3314, A3 => n1898, ZN => 
                           n16969);
   U1374 : AND3_X1 port map( A1 => n1079, A2 => n1077, A3 => n1075, ZN => 
                           n16240);
   U1375 : INV_X1 port map( A => n16045, ZN => n335);
   U1378 : NAND2_X1 port map( A1 => n565, A2 => n1154, ZN => n16292);
   U1379 : NAND3_X1 port map( A1 => n1645, A2 => n1644, A3 => n1650, ZN => 
                           n16507);
   U1381 : NAND2_X1 port map( A1 => n15796, A2 => n691, ZN => n690);
   U1382 : OR2_X1 port map( A1 => n15771, A2 => n15665, ZN => n1443);
   U1383 : MUX2_X1 port map( A => n15058, B => n15057, S => n15409, Z => n16269
                           );
   U1385 : OR2_X1 port map( A1 => n717, A2 => n15846, ZN => n714);
   U1386 : OR2_X1 port map( A1 => n15227, A2 => n15451, ZN => n349);
   U1387 : OAI21_X1 port map( B1 => n15307, B2 => n15306, A => n361, ZN => 
                           n2969);
   U1388 : MUX2_X1 port map( A => n15364, B => n15045, S => n1520, Z => n14951)
                           ;
   U1389 : INV_X1 port map( A => n717, ZN => n15640);
   U1390 : AND2_X1 port map( A1 => n13181, A2 => n2023, ZN => n783);
   U1391 : NOR2_X1 port map( A1 => n15857, A2 => n15720, ZN => n15171);
   U1392 : NAND2_X1 port map( A1 => n3496, A2 => n14586, ZN => n15270);
   U1395 : AND2_X1 port map( A1 => n16128, A2 => n15734, ZN => n387);
   U1398 : INV_X1 port map( A => n14954, ZN => n15808);
   U1399 : OR2_X1 port map( A1 => n546, A2 => n15474, ZN => n2113);
   U1400 : INV_X1 port map( A => n15060, ZN => n15307);
   U1401 : NAND2_X1 port map( A1 => n15812, A2 => n15813, ZN => n3313);
   U1403 : CLKBUF_X1 port map( A => n14312, Z => n15056);
   U1405 : AND2_X1 port map( A1 => n15070, A2 => n15405, ZN => n15617);
   U1406 : OR2_X1 port map( A1 => n14754, A2 => n14757, ZN => n15822);
   U1407 : AND2_X1 port map( A1 => n2889, A2 => n14702, ZN => n942);
   U1408 : INV_X1 port map( A => n15796, ZN => n15364);
   U1409 : OAI21_X1 port map( B1 => n914, B2 => n14489, A => n14488, ZN => 
                           n15132);
   U1411 : INV_X1 port map( A => n15311, ZN => n361);
   U1412 : INV_X1 port map( A => n15028, ZN => n3621);
   U1413 : INV_X1 port map( A => n15671, ZN => n15666);
   U1414 : INV_X1 port map( A => n15812, ZN => n228);
   U1415 : AND3_X1 port map( A1 => n1743, A2 => n1741, A3 => n1739, ZN => 
                           n15673);
   U1417 : AOI21_X1 port map( B1 => n14538, B2 => n2676, A => n14537, ZN => 
                           n14997);
   U1420 : NOR2_X1 port map( A1 => n14670, A2 => n14671, ZN => n859);
   U1421 : INV_X1 port map( A => n15657, ZN => n229);
   U1422 : INV_X1 port map( A => n15846, ZN => n230);
   U1429 : INV_X1 port map( A => n15491, ZN => n15755);
   U1431 : OAI22_X1 port map( A1 => n13953, A2 => n13952, B1 => n2642, B2 => 
                           n14134, ZN => n16011);
   U1432 : INV_X1 port map( A => n15490, ZN => n15588);
   U1433 : INV_X1 port map( A => n20183, ZN => n232);
   U1435 : OR2_X1 port map( A1 => n15815, A2 => n15813, ZN => n15035);
   U1436 : INV_X1 port map( A => n15813, ZN => n233);
   U1437 : OR3_X1 port map( A1 => n14198, A2 => n14197, A3 => n14590, ZN => 
                           n2789);
   U1438 : INV_X1 port map( A => n15667, ZN => n234);
   U1439 : OR2_X1 port map( A1 => n13957, A2 => n14705, ZN => n402);
   U1441 : MUX2_X1 port map( A => n14669, B => n14668, S => n14667, Z => n14670
                           );
   U1442 : XNOR2_X1 port map( A => n13680, B => n13681, ZN => n14718);
   U1443 : MUX2_X1 port map( A => n13948, B => n13947, S => n200, Z => n13949);
   U1445 : BUF_X1 port map( A => n13901, Z => n14782);
   U1446 : BUF_X1 port map( A => n14727, Z => n14408);
   U1447 : INV_X1 port map( A => n14548, ZN => n14654);
   U1448 : INV_X1 port map( A => n13940, ZN => n2039);
   U1450 : XNOR2_X1 port map( A => n3236, B => n12015, ZN => n14203);
   U1452 : AND2_X1 port map( A1 => n13865, A2 => n14441, ZN => n2983);
   U1457 : XNOR2_X1 port map( A => n13187, B => n13188, ZN => n14548);
   U1459 : INV_X1 port map( A => n14818, ZN => n3444);
   U1460 : INV_X1 port map( A => n14820, ZN => n235);
   U1462 : CLKBUF_X1 port map( A => n13872, Z => n14524);
   U1463 : INV_X1 port map( A => n14724, ZN => n236);
   U1464 : AND2_X1 port map( A1 => n951, A2 => n14648, ZN => n779);
   U1465 : XNOR2_X1 port map( A => n13034, B => n2240, ZN => n13868);
   U1467 : INV_X1 port map( A => n14522, ZN => n237);
   U1469 : INV_X1 port map( A => n14442, ZN => n238);
   U1471 : INV_X1 port map( A => n14199, ZN => n239);
   U1472 : XNOR2_X1 port map( A => n13669, B => n13670, ZN => n14714);
   U1473 : XNOR2_X1 port map( A => n13286, B => n13285, ZN => n14563);
   U1475 : XNOR2_X1 port map( A => n13801, B => n13800, ZN => n14239);
   U1476 : INV_X1 port map( A => n14228, ZN => n240);
   U1477 : INV_X1 port map( A => n20266, ZN => n241);
   U1478 : XNOR2_X1 port map( A => n13242, B => n627, ZN => n13246);
   U1479 : XNOR2_X1 port map( A => n13028, B => n979, ZN => n1089);
   U1480 : INV_X1 port map( A => n12977, ZN => n13757);
   U1481 : INV_X1 port map( A => n13231, ZN => n13706);
   U1482 : XNOR2_X1 port map( A => n13136, B => n13088, ZN => n13382);
   U1483 : XNOR2_X1 port map( A => n13193, B => n18478, ZN => n12999);
   U1485 : XNOR2_X1 port map( A => n13755, B => n13687, ZN => n627);
   U1490 : XNOR2_X1 port map( A => n12173, B => n357, ZN => n13086);
   U1493 : XNOR2_X1 port map( A => n13703, B => n13059, ZN => n12826);
   U1494 : AND4_X1 port map( A1 => n3530, A2 => n11139, A3 => n11137, A4 => 
                           n11138, ZN => n13330);
   U1496 : INV_X1 port map( A => n12709, ZN => n13827);
   U1497 : AND2_X1 port map( A1 => n553, A2 => n552, ZN => n551);
   U1501 : OR2_X1 port map( A1 => n12557, A2 => n12558, ZN => n13017);
   U1505 : OAI21_X1 port map( B1 => n12815, B2 => n12814, A => n12813, ZN => 
                           n13287);
   U1506 : NAND3_X1 port map( A1 => n2432, A2 => n12140, A3 => n2431, ZN => 
                           n13446);
   U1507 : XNOR2_X1 port map( A => n13511, B => n19205, ZN => n3365);
   U1509 : INV_X1 port map( A => n12770, ZN => n13745);
   U1511 : OAI211_X1 port map( C1 => n12359, C2 => n12506, A => n12012, B => 
                           n12011, ZN => n13673);
   U1513 : OAI211_X1 port map( C1 => n741, C2 => n11730, A => n3816, B => n740,
                           ZN => n12770);
   U1514 : OR2_X1 port map( A1 => n1366, A2 => n685, ZN => n684);
   U1515 : AOI22_X1 port map( A1 => n10822, A2 => n12206, B1 => n2713, B2 => 
                           n12211, ZN => n2711);
   U1516 : OAI21_X1 port map( B1 => n11983, B2 => n12619, A => n11982, ZN => 
                           n13634);
   U1519 : OR2_X1 port map( A1 => n11832, A2 => n11833, ZN => n1471);
   U1520 : INV_X1 port map( A => n11793, ZN => n850);
   U1523 : OR2_X1 port map( A1 => n20457, A2 => n12642, ZN => n491);
   U1524 : AND2_X1 port map( A1 => n13145, A2 => n13147, ZN => n356);
   U1526 : AND2_X1 port map( A1 => n12589, A2 => n12202, ZN => n563);
   U1527 : OR2_X1 port map( A1 => n11658, A2 => n11951, ZN => n488);
   U1528 : NOR2_X1 port map( A1 => n12639, A2 => n12455, ZN => n12637);
   U1529 : OAI21_X1 port map( B1 => n698, B2 => n12131, A => n12130, ZN => n697
                           );
   U1531 : NOR2_X1 port map( A1 => n12084, A2 => n12416, ZN => n369);
   U1532 : INV_X1 port map( A => n12174, ZN => n415);
   U1534 : OR2_X1 port map( A1 => n11670, A2 => n12180, ZN => n11672);
   U1535 : OR2_X1 port map( A1 => n12514, A2 => n11997, ZN => n521);
   U1536 : AND3_X1 port map( A1 => n10848, A2 => n2060, A3 => n2061, ZN => 
                           n12201);
   U1537 : INV_X1 port map( A => n12250, ZN => n242);
   U1538 : OAI211_X1 port map( C1 => n12437, C2 => n12442, A => n11942, B => 
                           n12443, ZN => n10686);
   U1539 : OR2_X1 port map( A1 => n11845, A2 => n20427, ZN => n588);
   U1543 : OR2_X1 port map( A1 => n11478, A2 => n3481, ZN => n313);
   U1544 : INV_X1 port map( A => n12532, ZN => n243);
   U1545 : OR2_X1 port map( A1 => n12636, A2 => n12449, ZN => n11948);
   U1546 : OR3_X1 port map( A1 => n12576, A2 => n11683, A3 => n11926, ZN => 
                           n3816);
   U1549 : INV_X1 port map( A => n953, ZN => n3586);
   U1551 : AND2_X1 port map( A1 => n3639, A2 => n3638, ZN => n12257);
   U1552 : INV_X1 port map( A => n12255, ZN => n244);
   U1553 : INV_X1 port map( A => n12759, ZN => n245);
   U1554 : INV_X1 port map( A => n11618, ZN => n246);
   U1556 : INV_X1 port map( A => n948, ZN => n247);
   U1558 : OR2_X1 port map( A1 => n10930, A2 => n10926, ZN => n1892);
   U1560 : CLKBUF_X1 port map( A => n11061, Z => n12016);
   U1561 : INV_X1 port map( A => n12417, ZN => n12084);
   U1562 : INV_X1 port map( A => n12263, ZN => n248);
   U1564 : NAND3_X1 port map( A1 => n11576, A2 => n11575, A3 => n3151, ZN => 
                           n12273);
   U1566 : INV_X1 port map( A => n12349, ZN => n249);
   U1569 : OAI21_X1 port map( B1 => n11407, B2 => n19506, A => n2810, ZN => 
                           n12544);
   U1570 : INV_X1 port map( A => n12554, ZN => n250);
   U1571 : INV_X1 port map( A => n12442, ZN => n251);
   U1575 : INV_X1 port map( A => n12180, ZN => n252);
   U1576 : INV_X1 port map( A => n12399, ZN => n253);
   U1577 : INV_X1 port map( A => n12408, ZN => n254);
   U1579 : OR2_X1 port map( A1 => n1279, A2 => n1280, ZN => n766);
   U1580 : AND2_X1 port map( A1 => n2043, A2 => n10861, ZN => n874);
   U1582 : AND2_X1 port map( A1 => n727, A2 => n725, ZN => n724);
   U1583 : INV_X1 port map( A => n12126, ZN => n255);
   U1585 : NOR2_X1 port map( A1 => n9413, A2 => n11281, ZN => n606);
   U1586 : INV_X1 port map( A => n11673, ZN => n256);
   U1587 : INV_X1 port map( A => n12415, ZN => n257);
   U1589 : OAI21_X1 port map( B1 => n11340, B2 => n10198, A => n10197, ZN => 
                           n11992);
   U1590 : OAI211_X1 port map( C1 => n11458, C2 => n1814, A => n11457, B => 
                           n1813, ZN => n12290);
   U1592 : CLKBUF_X1 port map( A => n10785, Z => n10814);
   U1593 : OR2_X1 port map( A1 => n11200, A2 => n11493, ZN => n798);
   U1594 : MUX2_X1 port map( A => n11525, B => n11524, S => n11523, Z => n11741
                           );
   U1595 : OR2_X1 port map( A1 => n10845, A2 => n10726, ZN => n11203);
   U1597 : INV_X1 port map( A => n12107, ZN => n765);
   U1598 : OR2_X1 port map( A1 => n11264, A2 => n11339, ZN => n753);
   U1599 : INV_X1 port map( A => n11574, ZN => n723);
   U1601 : OR2_X1 port map( A1 => n11006, A2 => n11005, ZN => n411);
   U1602 : OR2_X1 port map( A1 => n11079, A2 => n3482, ZN => n11080);
   U1603 : OAI21_X1 port map( B1 => n732, B2 => n11539, A => n731, ZN => n10738
                           );
   U1604 : NOR2_X1 port map( A1 => n11168, A2 => n11538, ZN => n732);
   U1605 : AND2_X1 port map( A1 => n12103, A2 => n11381, ZN => n12107);
   U1607 : INV_X1 port map( A => n11538, ZN => n11171);
   U1608 : MUX2_X1 port map( A => n10758, B => n10757, S => n10756, Z => n10759
                           );
   U1609 : INV_X1 port map( A => n11275, ZN => n764);
   U1610 : OR2_X1 port map( A1 => n20517, A2 => n11866, ZN => n1403);
   U1611 : BUF_X1 port map( A => n9616, Z => n10701);
   U1612 : INV_X1 port map( A => n11087, ZN => n11114);
   U1613 : OR2_X1 port map( A1 => n11538, A2 => n10640, ZN => n11540);
   U1614 : OR2_X1 port map( A1 => n9830, A2 => n10673, ZN => n756);
   U1615 : NAND2_X1 port map( A1 => n11133, A2 => n19959, ZN => n3295);
   U1616 : OR2_X1 port map( A1 => n11476, A2 => n11475, ZN => n10893);
   U1617 : NOR2_X1 port map( A1 => n3588, A2 => n11294, ZN => n11405);
   U1620 : OR2_X1 port map( A1 => n11489, A2 => n11493, ZN => n11198);
   U1622 : OR2_X1 port map( A1 => n11437, A2 => n11440, ZN => n11916);
   U1625 : XNOR2_X1 port map( A => n9428, B => n9944, ZN => n11277);
   U1627 : CLKBUF_X1 port map( A => n10726, Z => n11201);
   U1628 : XNOR2_X1 port map( A => n10269, B => n10268, ZN => n11325);
   U1631 : INV_X1 port map( A => n11535, ZN => n731);
   U1632 : OR2_X1 port map( A1 => n11302, A2 => n19750, ZN => n11387);
   U1634 : INV_X1 port map( A => n11550, ZN => n258);
   U1635 : XNOR2_X1 port map( A => n9816, B => n9815, ZN => n9830);
   U1636 : XNOR2_X1 port map( A => n2938, B => n9997, ZN => n11513);
   U1637 : INV_X1 port map( A => n11510, ZN => n259);
   U1638 : CLKBUF_X1 port map( A => n11113, Z => n11456);
   U1640 : CLKBUF_X1 port map( A => n9551, Z => n11010);
   U1643 : XNOR2_X1 port map( A => n8900, B => n8899, ZN => n11539);
   U1644 : XNOR2_X1 port map( A => n10162, B => n10161, ZN => n11428);
   U1646 : XNOR2_X1 port map( A => n9829, B => n9828, ZN => n11339);
   U1647 : XNOR2_X1 port map( A => n10408, B => n10407, ZN => n10829);
   U1653 : XNOR2_X1 port map( A => n802, B => n801, ZN => n9603);
   U1655 : INV_X1 port map( A => n9462, ZN => n790);
   U1656 : XNOR2_X1 port map( A => n9602, B => n9983, ZN => n802);
   U1657 : CLKBUF_X1 port map( A => n9537, Z => n10483);
   U1658 : XNOR2_X1 port map( A => n9646, B => n768, ZN => n10238);
   U1659 : XNOR2_X1 port map( A => n10281, B => n9862, ZN => n10563);
   U1660 : INV_X1 port map( A => n10185, ZN => n10441);
   U1661 : XNOR2_X1 port map( A => n9623, B => n9624, ZN => n10343);
   U1662 : XNOR2_X1 port map( A => n9646, B => n767, ZN => n9388);
   U1665 : INV_X1 port map( A => n9414, ZN => n10143);
   U1666 : BUF_X1 port map( A => n9856, Z => n10205);
   U1667 : XNOR2_X1 port map( A => n10237, B => n1228, ZN => n1227);
   U1670 : NAND4_X1 port map( A1 => n3200, A2 => n8935, A3 => n3199, A4 => 
                           n3799, ZN => n9624);
   U1672 : NAND3_X1 port map( A1 => n7900, A2 => n7901, A3 => n7899, ZN => 
                           n10528);
   U1674 : OAI211_X1 port map( C1 => n9218, C2 => n8670, A => n8669, B => n8668
                           , ZN => n10332);
   U1675 : XNOR2_X1 port map( A => n9414, B => n17024, ZN => n801);
   U1676 : OAI211_X1 port map( C1 => n6215, C2 => n9238, A => n6214, B => n6213
                           , ZN => n9819);
   U1681 : NAND2_X1 port map( A1 => n7658, A2 => n2336, ZN => n9430);
   U1682 : AND3_X1 port map( A1 => n8851, A2 => n590, A3 => n589, ZN => n7175);
   U1683 : AND2_X1 port map( A1 => n9160, A2 => n436, ZN => n1257);
   U1685 : OAI211_X1 port map( C1 => n9152, C2 => n1544, A => n1543, B => n1542
                           , ZN => n10061);
   U1688 : AND2_X1 port map( A1 => n8475, A2 => n8976, ZN => n577);
   U1692 : OR2_X1 port map( A1 => n9566, A2 => n9346, ZN => n2171);
   U1693 : INV_X1 port map( A => n10157, ZN => n260);
   U1694 : OR2_X1 port map( A1 => n9059, A2 => n9031, ZN => n3072);
   U1695 : OR2_X1 port map( A1 => n9298, A2 => n7424, ZN => n7440);
   U1696 : NOR2_X1 port map( A1 => n8987, A2 => n9172, ZN => n8763);
   U1697 : OR2_X1 port map( A1 => n1765, A2 => n9031, ZN => n1766);
   U1698 : OR2_X1 port map( A1 => n8498, A2 => n8499, ZN => n704);
   U1699 : OR2_X1 port map( A1 => n8965, A2 => n207, ZN => n838);
   U1702 : OR2_X1 port map( A1 => n8960, A2 => n8959, ZN => n7559);
   U1703 : OR2_X1 port map( A1 => n8338, A2 => n8790, ZN => n8439);
   U1706 : INV_X1 port map( A => n9300, ZN => n9297);
   U1707 : OR2_X1 port map( A1 => n978, A2 => n19490, ZN => n464);
   U1709 : INV_X1 port map( A => n2097, ZN => n9238);
   U1711 : AND2_X1 port map( A1 => n778, A2 => n777, ZN => n7996);
   U1712 : AND2_X1 port map( A1 => n8499, A2 => n8733, ZN => n7665);
   U1714 : INV_X1 port map( A => n8923, ZN => n3645);
   U1715 : INV_X1 port map( A => n8786, ZN => n261);
   U1716 : NOR2_X1 port map( A1 => n8125, A2 => n8124, ZN => n8995);
   U1719 : NAND2_X1 port map( A1 => n737, A2 => n7509, ZN => n9049);
   U1720 : OAI211_X1 port map( C1 => n7505, C2 => n7931, A => n7506, B => n1402
                           , ZN => n9287);
   U1721 : AND2_X1 port map( A1 => n9114, A2 => n9113, ZN => n9219);
   U1722 : INV_X1 port map( A => n9333, ZN => n262);
   U1723 : OR2_X1 port map( A1 => n9168, A2 => n8569, ZN => n777);
   U1726 : INV_X1 port map( A => n9210, ZN => n263);
   U1727 : NAND3_X1 port map( A1 => n2156, A2 => n2155, A3 => n6894, ZN => 
                           n9228);
   U1728 : INV_X1 port map( A => n655, ZN => n9233);
   U1729 : INV_X1 port map( A => n8569, ZN => n264);
   U1730 : OAI21_X1 port map( B1 => n8137, B2 => n8138, A => n8136, ZN => n352)
                           ;
   U1732 : OAI21_X1 port map( B1 => n6701, B2 => n8261, A => n6700, ZN => n9305
                           );
   U1733 : INV_X1 port map( A => n8985, ZN => n265);
   U1736 : INV_X1 port map( A => n9162, ZN => n437);
   U1741 : INV_X1 port map( A => n9189, ZN => n266);
   U1742 : INV_X1 port map( A => n6587, ZN => n267);
   U1745 : INV_X1 port map( A => n9242, ZN => n268);
   U1747 : INV_X1 port map( A => n8568, ZN => n269);
   U1748 : INV_X1 port map( A => n9018, ZN => n270);
   U1751 : INV_X1 port map( A => n770, ZN => n8434);
   U1753 : INV_X1 port map( A => n9166, ZN => n8705);
   U1756 : AND3_X1 port map( A1 => n493, A2 => n6284, A3 => n6283, ZN => n8470)
                           ;
   U1757 : OR2_X1 port map( A1 => n7807, A2 => n462, ZN => n461);
   U1758 : OR2_X1 port map( A1 => n8236, A2 => n6539, ZN => n770);
   U1760 : OR2_X1 port map( A1 => n7499, A2 => n163, ZN => n3377);
   U1761 : CLKBUF_X1 port map( A => n7717, Z => n7723);
   U1764 : AND3_X1 port map( A1 => n7760, A2 => n6903, A3 => n3089, ZN => n9162
                           );
   U1767 : AOI21_X1 port map( B1 => n1198, B2 => n7541, A => n1197, ZN => n8823
                           );
   U1769 : AND3_X1 port map( A1 => n2934, A2 => n8368, A3 => n8367, ZN => n8420
                           );
   U1770 : AND2_X1 port map( A1 => n7513, A2 => n7514, ZN => n738);
   U1771 : AOI211_X1 port map( C1 => n7912, C2 => n7745, A => n6908, B => n7911
                           , ZN => n6909);
   U1772 : INV_X1 port map( A => n7602, ZN => n7793);
   U1773 : OR2_X1 port map( A1 => n7417, A2 => n8068, ZN => n428);
   U1774 : INV_X1 port map( A => n8091, ZN => n718);
   U1775 : OR2_X1 port map( A1 => n6539, A2 => n19826, ZN => n358);
   U1776 : NAND3_X1 port map( A1 => n8183, A2 => n7464, A3 => n7463, ZN => 
                           n9023);
   U1777 : BUF_X1 port map( A => n7389, Z => n7807);
   U1778 : AND2_X1 port map( A1 => n20195, A2 => n7936, ZN => n6244);
   U1779 : AND2_X1 port map( A1 => n8010, A2 => n1560, ZN => n427);
   U1780 : INV_X1 port map( A => n1726, ZN => n505);
   U1783 : INV_X1 port map( A => n8003, ZN => n324);
   U1785 : OR2_X1 port map( A1 => n7903, A2 => n7530, ZN => n494);
   U1786 : OR2_X1 port map( A1 => n7918, A2 => n7917, ZN => n376);
   U1787 : AND2_X1 port map( A1 => n8212, A2 => n8095, ZN => n8091);
   U1788 : NOR2_X1 port map( A1 => n7801, A2 => n208, ZN => n629);
   U1789 : AND2_X1 port map( A1 => n8300, A2 => n5941, ZN => n7787);
   U1790 : INV_X1 port map( A => n7967, ZN => n776);
   U1794 : XNOR2_X1 port map( A => n1074, B => n1073, ZN => n8251);
   U1796 : XNOR2_X1 port map( A => n6823, B => n6822, ZN => n8159);
   U1799 : BUF_X1 port map( A => n6312, Z => n7982);
   U1800 : OR2_X1 port map( A1 => n7833, A2 => n8910, ZN => n7773);
   U1801 : INV_X1 port map( A => n7991, ZN => n273);
   U1802 : INV_X1 port map( A => n7908, ZN => n274);
   U1806 : XNOR2_X1 port map( A => n639, B => n6691, ZN => n895);
   U1807 : INV_X1 port map( A => n8325, ZN => n276);
   U1808 : XNOR2_X1 port map( A => n6372, B => n6371, ZN => n7709);
   U1809 : XNOR2_X1 port map( A => n6583, B => n6582, ZN => n8111);
   U1810 : XNOR2_X1 port map( A => n6291, B => n6292, ZN => n7978);
   U1811 : INV_X1 port map( A => n7631, ZN => n2703);
   U1812 : INV_X1 port map( A => n2977, ZN => n277);
   U1813 : XNOR2_X1 port map( A => n2622, B => n5898, ZN => n5941);
   U1814 : INV_X1 port map( A => n7971, ZN => n278);
   U1815 : XNOR2_X1 port map( A => n7075, B => n7076, ZN => n1560);
   U1817 : INV_X1 port map( A => n7855, ZN => n279);
   U1819 : INV_X1 port map( A => n7754, ZN => n280);
   U1820 : INV_X1 port map( A => n7475, ZN => n281);
   U1821 : XNOR2_X1 port map( A => n7236, B => n7235, ZN => n8016);
   U1823 : INV_X1 port map( A => n6830, ZN => n282);
   U1826 : AND2_X1 port map( A1 => n6217, A2 => n6221, ZN => n7360);
   U1827 : INV_X1 port map( A => n6690, ZN => n639);
   U1828 : XNOR2_X1 port map( A => n459, B => n6032, ZN => n6040);
   U1829 : XNOR2_X1 port map( A => n7178, B => n7273, ZN => n6838);
   U1830 : XNOR2_X1 port map( A => n6024, B => n7333, ZN => n459);
   U1833 : INV_X1 port map( A => n3068, ZN => n7305);
   U1834 : INV_X1 port map( A => n7143, ZN => n353);
   U1836 : OAI21_X1 port map( B1 => n6148, B2 => n6147, A => n6146, ZN => n7206
                           );
   U1838 : XNOR2_X1 port map( A => n354, B => n7274, ZN => n6593);
   U1840 : OAI211_X1 port map( C1 => n5620, C2 => n6143, A => n5619, B => n5618
                           , ZN => n6713);
   U1844 : AND2_X1 port map( A1 => n6207, A2 => n6208, ZN => n6221);
   U1846 : INV_X1 port map( A => n354, ZN => n6793);
   U1847 : XNOR2_X1 port map( A => n3663, B => n7146, ZN => n6506);
   U1853 : NAND2_X1 port map( A1 => n2524, A2 => n480, ZN => n6719);
   U1854 : OR2_X1 port map( A1 => n5359, A2 => n5358, ZN => n7142);
   U1859 : OAI21_X1 port map( B1 => n6192, B2 => n5234, A => n5233, ZN => n6919
                           );
   U1862 : INV_X1 port map( A => n6220, ZN => n3674);
   U1864 : AOI22_X1 port map( A1 => n5348, A2 => n5720, B1 => n3664, B2 => 
                           n5347, ZN => n5984);
   U1865 : MUX2_X1 port map( A => n4689, B => n4688, S => n6172, Z => n4690);
   U1869 : MUX2_X1 port map( A => n5446, B => n5445, S => n5645, Z => n7257);
   U1870 : OR2_X1 port map( A1 => n6003, A2 => n6000, ZN => n3602);
   U1873 : NOR2_X1 port map( A1 => n6173, A2 => n5842, ZN => n568);
   U1875 : OR2_X1 port map( A1 => n5868, A2 => n6119, ZN => n2092);
   U1877 : AOI21_X1 port map( B1 => n2407, B2 => n5790, A => n5428, ZN => n2879
                           );
   U1878 : OR2_X1 port map( A1 => n6379, A2 => n5847, ZN => n5848);
   U1879 : INV_X1 port map( A => n5953, ZN => n283);
   U1880 : OR2_X1 port map( A1 => n5622, A2 => n5623, ZN => n6134);
   U1881 : OR2_X1 port map( A1 => n5745, A2 => n5742, ZN => n1883);
   U1883 : OAI21_X1 port map( B1 => n5322, B2 => n5395, A => n1838, ZN => n533)
                           ;
   U1884 : AND2_X1 port map( A1 => n5930, A2 => n6027, ZN => n5596);
   U1885 : AND2_X1 port map( A1 => n5201, A2 => n5745, ZN => n455);
   U1886 : OR3_X1 port map( A1 => n5823, A2 => n6017, A3 => n6016, ZN => n5829)
                           ;
   U1888 : AND2_X1 port map( A1 => n618, A2 => n617, ZN => n5742);
   U1890 : NOR2_X1 port map( A1 => n1685, A2 => n3606, ZN => n5718);
   U1891 : OR2_X1 port map( A1 => n5393, A2 => n5395, ZN => n5369);
   U1892 : BUF_X1 port map( A => n5483, Z => n5716);
   U1893 : INV_X1 port map( A => n3701, ZN => n5748);
   U1894 : OR2_X1 port map( A1 => n5328, A2 => n6049, ZN => n3919);
   U1895 : INV_X1 port map( A => n6124, ZN => n6120);
   U1896 : AND2_X1 port map( A1 => n4282, A2 => n4281, ZN => n508);
   U1898 : INV_X1 port map( A => n5952, ZN => n284);
   U1902 : INV_X1 port map( A => n733, ZN => n5571);
   U1905 : INV_X1 port map( A => n5985, ZN => n285);
   U1906 : NAND4_X1 port map( A1 => n760, A2 => n761, A3 => n3714, A4 => n762, 
                           ZN => n3701);
   U1907 : NAND2_X1 port map( A1 => n2572, A2 => n2573, ZN => n5611);
   U1908 : INV_X1 port map( A => n5802, ZN => n5378);
   U1909 : INV_X1 port map( A => n6068, ZN => n473);
   U1910 : NAND2_X1 port map( A1 => n4301, A2 => n4300, ZN => n5363);
   U1911 : NAND2_X1 port map( A1 => n4120, A2 => n4121, ZN => n5971);
   U1912 : OAI21_X1 port map( B1 => n4124, B2 => n4985, A => n4123, ZN => n5699
                           );
   U1917 : INV_X1 port map( A => n5251, ZN => n5398);
   U1918 : INV_X1 port map( A => n5172, ZN => n5957);
   U1919 : NOR2_X1 port map( A1 => n5531, A2 => n6036, ZN => n5566);
   U1921 : INV_X1 port map( A => n5747, ZN => n286);
   U1926 : OAI21_X1 port map( B1 => n4364, B2 => n604, A => n603, ZN => n4375);
   U1927 : OR2_X1 port map( A1 => n4034, A2 => n4033, ZN => n1214);
   U1930 : OAI211_X1 port map( C1 => n4980, C2 => n4979, A => n4978, B => n3517
                           , ZN => n5563);
   U1931 : OAI211_X1 port map( C1 => n4964, C2 => n210, A => n3232, B => n3229,
                           ZN => n5531);
   U1932 : MUX2_X1 port map( A => n4949, B => n4948, S => n4947, Z => n5532);
   U1933 : OAI21_X1 port map( B1 => n4506, B2 => n4567, A => n4505, ZN => n5766
                           );
   U1936 : OR2_X1 port map( A1 => n821, A2 => n4652, ZN => n4873);
   U1937 : OAI211_X1 port map( C1 => n4607, C2 => n4153, A => n1253, B => n680,
                           ZN => n733);
   U1938 : INV_X1 port map( A => n6205, ZN => n287);
   U1940 : OR2_X1 port map( A1 => n665, A2 => n4569, ZN => n643);
   U1941 : INV_X1 port map( A => n19475, ZN => n288);
   U1942 : INV_X1 port map( A => n5072, ZN => n828);
   U1943 : OR2_X1 port map( A1 => n4681, A2 => n4387, ZN => n523);
   U1944 : AND2_X1 port map( A1 => n4337, A2 => n20487, ZN => n4535);
   U1945 : OR2_X1 port map( A1 => n3624, A2 => n20487, ZN => n393);
   U1947 : OR2_X1 port map( A1 => n3854, A2 => n4674, ZN => n306);
   U1948 : OR2_X1 port map( A1 => n4732, A2 => n3683, ZN => n3682);
   U1949 : AND2_X1 port map( A1 => n4365, A2 => n4013, ZN => n1535);
   U1950 : BUF_X1 port map( A => n4021, Z => n4976);
   U1951 : OR2_X1 port map( A1 => n896, A2 => n20357, ZN => n453);
   U1953 : OR2_X1 port map( A1 => n5100, A2 => n5101, ZN => n4049);
   U1954 : OR2_X1 port map( A1 => n4652, A2 => n20357, ZN => n4863);
   U1955 : CLKBUF_X1 port map( A => n3995, Z => n4387);
   U1956 : OR2_X1 port map( A1 => n4548, A2 => n4152, ZN => n4153);
   U1957 : CLKBUF_X1 port map( A => n4232, Z => n4902);
   U1959 : CLKBUF_X1 port map( A => n4445, Z => n4585);
   U1961 : OR2_X1 port map( A1 => n4271, A2 => n4268, ZN => n556);
   U1962 : INV_X1 port map( A => n2233, ZN => n357);
   U1963 : INV_X1 port map( A => n20355, ZN => n289);
   U1964 : INV_X1 port map( A => n5079, ZN => n378);
   U1966 : AND2_X1 port map( A1 => n5022, A2 => n19788, ZN => n315);
   U1967 : INV_X1 port map( A => n4365, ZN => n290);
   U1968 : INV_X1 port map( A => n4663, ZN => n291);
   U1969 : CLKBUF_X1 port map( A => n4602, Z => n4361);
   U1970 : OR2_X1 port map( A1 => n4638, A2 => n4528, ZN => n4636);
   U1971 : BUF_X1 port map( A => n4439, Z => n5042);
   U1972 : CLKBUF_X1 port map( A => n4187, Z => n4522);
   U1973 : OR2_X1 port map( A1 => n4110, A2 => n4277, ZN => n672);
   U1974 : XNOR2_X1 port map( A => n1581, B => Key(76), ZN => n4214);
   U1975 : OR2_X1 port map( A1 => n20143, A2 => n4285, ZN => n4630);
   U1976 : CLKBUF_X1 port map( A => n4048, Z => n5105);
   U1977 : AND2_X1 port map( A1 => n4623, A2 => n4626, ZN => n531);
   U1979 : BUF_X1 port map( A => n4575, Z => n4372);
   U1980 : CLKBUF_X1 port map( A => Key(183), Z => n18997);
   U1982 : CLKBUF_X1 port map( A => Key(190), Z => n2035);
   U1983 : CLKBUF_X1 port map( A => Key(176), Z => n2382);
   U1984 : INV_X1 port map( A => n4894, ZN => n292);
   U1985 : CLKBUF_X1 port map( A => Key(136), Z => n2417);
   U1987 : INV_X1 port map( A => n2082, ZN => n293);
   U1988 : INV_X1 port map( A => n1857, ZN => n294);
   U1989 : INV_X1 port map( A => n2218, ZN => n295);
   U1990 : XNOR2_X1 port map( A => Key(81), B => Plaintext(81), ZN => n5117);
   U1991 : CLKBUF_X1 port map( A => Key(50), Z => n19457);
   U1992 : INV_X1 port map( A => n18801, ZN => n296);
   U1993 : CLKBUF_X1 port map( A => Key(1), Z => n17787);
   U1995 : CLKBUF_X1 port map( A => Key(22), Z => n2275);
   U1996 : CLKBUF_X1 port map( A => Key(165), Z => n2381);
   U2000 : CLKBUF_X1 port map( A => Key(95), Z => n17989);
   U2001 : CLKBUF_X1 port map( A => Key(81), Z => n17024);
   U2002 : CLKBUF_X1 port map( A => Key(53), Z => n18146);
   U2003 : CLKBUF_X1 port map( A => Key(99), Z => n18308);
   U2004 : CLKBUF_X1 port map( A => Key(97), Z => n19410);
   U2005 : CLKBUF_X1 port map( A => Key(177), Z => n17686);
   U2006 : INV_X1 port map( A => n17544, ZN => n298);
   U2007 : CLKBUF_X1 port map( A => Key(184), Z => n2401);
   U2008 : CLKBUF_X1 port map( A => Key(132), Z => n18809);
   U2009 : CLKBUF_X1 port map( A => Key(79), Z => n19180);
   U2010 : CLKBUF_X1 port map( A => Key(139), Z => n2383);
   U2011 : CLKBUF_X1 port map( A => Key(160), Z => n18819);
   U2012 : CLKBUF_X1 port map( A => Key(13), Z => n2455);
   U2013 : CLKBUF_X1 port map( A => Key(65), Z => n1840);
   U2015 : XNOR2_X1 port map( A => Key(72), B => Plaintext(72), ZN => n4829);
   U2016 : CLKBUF_X1 port map( A => Key(59), Z => n18078);
   U2017 : INV_X1 port map( A => n2096, ZN => n299);
   U2018 : CLKBUF_X1 port map( A => Key(174), Z => n2108);
   U2019 : CLKBUF_X1 port map( A => Key(180), Z => n17637);
   U2020 : INV_X1 port map( A => n17733, ZN => n300);
   U2022 : INV_X1 port map( A => n4541, ZN => n301);
   U2023 : CLKBUF_X1 port map( A => Key(164), Z => n2384);
   U2024 : INV_X1 port map( A => n1969, ZN => n302);
   U2025 : CLKBUF_X1 port map( A => Key(189), Z => n2420);
   U2026 : XNOR2_X1 port map( A => Key(166), B => Plaintext(166), ZN => n4349);
   U2031 : INV_X1 port map( A => n4107, ZN => n303);
   U2032 : CLKBUF_X1 port map( A => Key(42), Z => n2216);
   U2033 : INV_X1 port map( A => n16035, ZN => n304);
   U2034 : CLKBUF_X1 port map( A => Key(7), Z => n2423);
   U2035 : CLKBUF_X1 port map( A => Key(28), Z => n1911);
   U2036 : CLKBUF_X1 port map( A => Key(98), Z => n17791);
   U2038 : NAND2_X1 port map( A1 => n4828, A2 => n19688, ZN => n4674);
   U2039 : NOR2_X1 port map( A1 => n14984, A2 => n15180, ZN => n307);
   U2040 : NAND3_X1 port map( A1 => n1822, A2 => n262, A3 => n8121, ZN => n8122
                           );
   U2041 : NOR3_X1 port map( A1 => n12223, A2 => n308, A3 => n10925, ZN => 
                           n12225);
   U2042 : INV_X1 port map( A => n12220, ZN => n308);
   U2043 : AND2_X1 port map( A1 => n8937, A2 => n8729, ZN => n8942);
   U2044 : NAND2_X1 port map( A1 => n8097, A2 => n309, ZN => n8103);
   U2045 : OAI21_X1 port map( B1 => n8210, B2 => n8091, A => n7631, ZN => n309)
                           ;
   U2046 : NAND2_X1 port map( A1 => n19724, A2 => n310, ZN => n18992);
   U2049 : OAI21_X1 port map( B1 => n19751, B2 => n19753, A => n312, ZN => 
                           n17630);
   U2050 : NAND2_X1 port map( A1 => n18703, A2 => n18697, ZN => n312);
   U2052 : NAND3_X1 port map( A1 => n3711, A2 => n11218, A3 => n3482, ZN => 
                           n11220);
   U2053 : NAND2_X1 port map( A1 => n1142, A2 => n1144, ZN => n1236);
   U2054 : NAND2_X1 port map( A1 => n314, A2 => n1235, ZN => n11597);
   U2055 : NAND2_X1 port map( A1 => n1234, A2 => n245, ZN => n314);
   U2057 : NAND2_X1 port map( A1 => n4581, A2 => n315, ZN => n4583);
   U2060 : INV_X1 port map( A => n8941, ZN => n317);
   U2061 : NAND2_X1 port map( A1 => n8942, A2 => n8941, ZN => n318);
   U2063 : NAND2_X1 port map( A1 => n321, A2 => n320, ZN => n319);
   U2064 : NAND2_X1 port map( A1 => n20129, A2 => n225, ZN => n321);
   U2066 : OR2_X1 port map( A1 => n5444, A2 => n5641, ZN => n5640);
   U2067 : NAND3_X1 port map( A1 => n3109, A2 => n4610, A3 => n4615, ZN => 
                           n3108);
   U2068 : NAND3_X1 port map( A1 => n7601, A2 => n7602, A3 => n8286, ZN => 
                           n2315);
   U2069 : OAI21_X2 port map( B1 => n14840, B2 => n14839, A => n322, ZN => 
                           n16614);
   U2070 : OAI21_X1 port map( B1 => n8004, B2 => n324, A => n323, ZN => n8009);
   U2071 : NAND2_X1 port map( A1 => n281, A2 => n8004, ZN => n323);
   U2072 : NOR2_X1 port map( A1 => n325, A2 => n147, ZN => n2152);
   U2073 : NOR2_X1 port map( A1 => n14652, A2 => n14651, ZN => n325);
   U2074 : NAND2_X1 port map( A1 => n17818, A2 => n18962, ZN => n326);
   U2075 : NAND3_X1 port map( A1 => n4789, A2 => n5092, A3 => n4782, ZN => 
                           n4070);
   U2076 : NAND2_X1 port map( A1 => n2460, A2 => n4405, ZN => n4789);
   U2078 : NAND3_X1 port map( A1 => n4604, A2 => n4603, A3 => n4354, ZN => 
                           n4606);
   U2079 : NAND2_X1 port map( A1 => n329, A2 => n2281, ZN => n478);
   U2080 : NAND2_X1 port map( A1 => n13955, A2 => n14566, ZN => n329);
   U2081 : NAND2_X1 port map( A1 => n10995, A2 => n10996, ZN => n10997);
   U2082 : NAND2_X1 port map( A1 => n4495, A2 => n4496, ZN => n4500);
   U2083 : NAND3_X1 port map( A1 => n20368, A2 => n6013, A3 => n5921, ZN => 
                           n5516);
   U2084 : OAI211_X1 port map( C1 => n245, C2 => n12754, A => n331, B => n12389
                           , ZN => n609);
   U2085 : NAND2_X1 port map( A1 => n12410, A2 => n254, ZN => n331);
   U2086 : NAND2_X1 port map( A1 => n12399, A2 => n953, ZN => n11912);
   U2089 : NAND2_X1 port map( A1 => n11336, A2 => n11265, ZN => n332);
   U2090 : NAND2_X1 port map( A1 => n11335, A2 => n11337, ZN => n333);
   U2091 : OAI22_X1 port map( A1 => n252, A2 => n256, B1 => n11673, B2 => 
                           n20427, ZN => n703);
   U2092 : NAND2_X1 port map( A1 => n7600, A2 => n8033, ZN => n7602);
   U2094 : NAND2_X1 port map( A1 => n4696, A2 => n4795, ZN => n4029);
   U2096 : NAND2_X1 port map( A1 => n7864, A2 => n8153, ZN => n6698);
   U2097 : OAI211_X1 port map( C1 => n9314, C2 => n9313, A => n9312, B => n9311
                           , ZN => n9856);
   U2098 : XNOR2_X1 port map( A => n17406, B => n335, ZN => n334);
   U2101 : NAND3_X1 port map( A1 => n336, A2 => n15467, A3 => n15466, ZN => 
                           n15472);
   U2102 : NAND2_X1 port map( A1 => n20502, A2 => n15465, ZN => n336);
   U2103 : OAI21_X1 port map( B1 => n3725, B2 => n15257, A => n1349, ZN => 
                           n15261);
   U2105 : NAND3_X1 port map( A1 => n5465, A2 => n5464, A3 => n5633, ZN => 
                           n5469);
   U2106 : NAND2_X1 port map( A1 => n5632, A2 => n5364, ZN => n5465);
   U2111 : NAND2_X1 port map( A1 => n12662, A2 => n12661, ZN => n338);
   U2112 : INV_X1 port map( A => n339, ZN => n17499);
   U2114 : NOR2_X1 port map( A1 => n20648, A2 => n17504, ZN => n339);
   U2115 : NAND2_X1 port map( A1 => n7766, A2 => n7919, ZN => n7536);
   U2118 : NAND2_X1 port map( A1 => n358, A2 => n7425, ZN => n7427);
   U2120 : NAND2_X1 port map( A1 => n14045, A2 => n14826, ZN => n340);
   U2121 : NAND2_X1 port map( A1 => n14833, A2 => n19859, ZN => n341);
   U2122 : NAND2_X1 port map( A1 => n1955, A2 => n15339, ZN => n2069);
   U2124 : NAND2_X1 port map( A1 => n5435, A2 => n5704, ZN => n6003);
   U2125 : NAND3_X1 port map( A1 => n19916, A2 => n17687, A3 => n18042, ZN => 
                           n17813);
   U2126 : NAND3_X1 port map( A1 => n15895, A2 => n19838, A3 => n15896, ZN => 
                           n15897);
   U2127 : NAND2_X1 port map( A1 => n5037, A2 => n153, ZN => n713);
   U2128 : XNOR2_X1 port map( A => n9987, B => n9947, ZN => n10417);
   U2129 : OAI21_X1 port map( B1 => n18223, B2 => n18977, A => n342, ZN => 
                           n16911);
   U2130 : NAND2_X1 port map( A1 => n224, A2 => n18977, ZN => n342);
   U2131 : OAI21_X1 port map( B1 => n684, B2 => n11726, A => n683, ZN => n682);
   U2132 : NAND2_X1 port map( A1 => n1177, A2 => n14954, ZN => n14743);
   U2134 : NAND2_X1 port map( A1 => n12250, A2 => n12573, ZN => n541);
   U2137 : NAND2_X1 port map( A1 => n6100, A2 => n283, ZN => n343);
   U2138 : NAND2_X1 port map( A1 => n5663, A2 => n5952, ZN => n6100);
   U2141 : NAND2_X1 port map( A1 => n11364, A2 => n2765, ZN => n344);
   U2142 : OR2_X1 port map( A1 => n8386, A2 => n8132, ZN => n2441);
   U2143 : XNOR2_X1 port map( A => n10593, B => n10592, ZN => n3051);
   U2144 : INV_X1 port map( A => n5428, ZN => n5797);
   U2145 : NAND2_X1 port map( A1 => n5338, A2 => n6124, ZN => n1382);
   U2146 : AND2_X2 port map( A1 => n1051, A2 => n1050, ZN => n6124);
   U2147 : NAND2_X1 port map( A1 => n19476, A2 => n6379, ZN => n5844);
   U2149 : NAND3_X1 port map( A1 => n6056, A2 => n20670, A3 => n5785, ZN => 
                           n5305);
   U2151 : NAND2_X1 port map( A1 => n346, A2 => n2618, ZN => n2617);
   U2152 : NAND2_X1 port map( A1 => n9174, A2 => n9175, ZN => n346);
   U2153 : NAND3_X1 port map( A1 => n820, A2 => n8202, A3 => n8201, ZN => n8207
                           );
   U2154 : NAND3_X1 port map( A1 => n3532, A2 => n14600, A3 => n20181, ZN => 
                           n1824);
   U2155 : NAND3_X1 port map( A1 => n3410, A2 => n5931, A3 => n5930, ZN => 
                           n5932);
   U2157 : NAND2_X1 port map( A1 => n14866, A2 => n15684, ZN => n15226);
   U2159 : NAND2_X1 port map( A1 => n9874, A2 => n11230, ZN => n348);
   U2161 : NAND2_X1 port map( A1 => n1987, A2 => n1183, ZN => n350);
   U2163 : NAND3_X1 port map( A1 => n6844, A2 => n279, A3 => n7852, ZN => n6845
                           );
   U2164 : NOR2_X1 port map( A1 => n351, A2 => n18504, ZN => n1660);
   U2165 : AOI21_X1 port map( B1 => n18518, B2 => n18511, A => n18512, ZN => 
                           n351);
   U2166 : AOI22_X1 port map( A1 => n11835, A2 => n12506, B1 => n12507, B2 => 
                           n12505, ZN => n11840);
   U2167 : NOR2_X1 port map( A1 => n390, A2 => n12642, ZN => n389);
   U2168 : NAND2_X1 port map( A1 => n352, A2 => n9564, ZN => n9193);
   U2169 : NAND2_X1 port map( A1 => n9338, A2 => n352, ZN => n8155);
   U2171 : XNOR2_X1 port map( A => n353, B => n6793, ZN => n7089);
   U2172 : XNOR2_X1 port map( A => n354, B => n7088, ZN => n6722);
   U2173 : NAND2_X1 port map( A1 => n5850, A2 => n5849, ZN => n355);
   U2174 : NAND2_X1 port map( A1 => n356, A2 => n244, ZN => n12018);
   U2175 : NAND2_X1 port map( A1 => n242, A2 => n356, ZN => n542);
   U2176 : INV_X1 port map( A => n358, ZN => n7859);
   U2178 : NAND2_X1 port map( A1 => n359, A2 => n9559, ZN => n3489);
   U2179 : NAND2_X1 port map( A1 => n2734, A2 => n10996, ZN => n359);
   U2180 : INV_X1 port map( A => n1640, ZN => n360);
   U2181 : NAND2_X1 port map( A1 => n15397, A2 => n361, ZN => n15064);
   U2182 : AND3_X2 port map( A1 => n3267, A2 => n3266, A3 => n3268, ZN => 
                           n15311);
   U2183 : OAI21_X1 port map( B1 => n8439, B2 => n2499, A => n364, ZN => n362);
   U2184 : AOI21_X1 port map( B1 => n365, B2 => n8337, A => n9144, ZN => n363);
   U2185 : NAND2_X1 port map( A1 => n9145, A2 => n2499, ZN => n364);
   U2186 : NAND2_X1 port map( A1 => n8338, A2 => n8786, ZN => n365);
   U2187 : NAND2_X1 port map( A1 => n8338, A2 => n2499, ZN => n8337);
   U2188 : NAND2_X1 port map( A1 => n6105, A2 => n6109, ZN => n368);
   U2189 : NAND2_X1 port map( A1 => n1623, A2 => n368, ZN => n1620);
   U2193 : NOR2_X1 port map( A1 => n5957, A2 => n368, ZN => n367);
   U2195 : NAND2_X1 port map( A1 => n12502, A2 => n12004, ZN => n12345);
   U2197 : NAND2_X1 port map( A1 => n19999, A2 => n11521, ZN => n370);
   U2199 : NAND3_X1 port map( A1 => n372, A2 => n1446, A3 => n10930, ZN => n371
                           );
   U2200 : NAND2_X1 port map( A1 => n10889, A2 => n11550, ZN => n10930);
   U2201 : NAND2_X1 port map( A1 => n10068, A2 => n11544, ZN => n372);
   U2202 : NAND2_X1 port map( A1 => n374, A2 => n646, ZN => n373);
   U2203 : NAND2_X1 port map( A1 => n648, A2 => n647, ZN => n374);
   U2204 : INV_X1 port map( A => n4349, ZN => n4199);
   U2205 : NAND2_X1 port map( A1 => n4349, A2 => n4541, ZN => n4536);
   U2206 : XNOR2_X2 port map( A => Key(167), B => Plaintext(167), ZN => n4541);
   U2207 : NAND2_X1 port map( A1 => n15766, A2 => n15474, ZN => n12664);
   U2208 : NAND3_X1 port map( A1 => n15766, A2 => n15474, A3 => n15769, ZN => 
                           n375);
   U2209 : NAND3_X1 port map( A1 => n7916, A2 => n377, A3 => n376, ZN => n9143)
                           ;
   U2210 : NAND2_X1 port map( A1 => n8910, A2 => n7956, ZN => n1231);
   U2211 : NAND2_X1 port map( A1 => n20431, A2 => n378, ZN => n4083);
   U2212 : OAI21_X1 port map( B1 => n378, B2 => n5074, A => n4809, ZN => n4084)
                           ;
   U2213 : NAND2_X1 port map( A1 => n4810, A2 => n378, ZN => n1047);
   U2214 : NAND2_X2 port map( A1 => n379, A2 => n14033, ZN => n15760);
   U2215 : NAND2_X1 port map( A1 => n14301, A2 => n14512, ZN => n379);
   U2216 : NAND2_X1 port map( A1 => n13986, A2 => n2972, ZN => n14301);
   U2217 : NAND4_X2 port map( A1 => n5391, A2 => n5390, A3 => n5389, A4 => 
                           n5388, ZN => n7128);
   U2220 : NAND2_X1 port map( A1 => n10784, A2 => n11435, ZN => n382);
   U2221 : NAND2_X1 port map( A1 => n5664, A2 => n5949, ZN => n5458);
   U2222 : NOR3_X1 port map( A1 => n9296, A2 => n9300, A3 => n9295, ZN => n2225
                           );
   U2224 : OAI21_X1 port map( B1 => n8297, B2 => n20485, A => n383, ZN => n7582
                           );
   U2225 : NAND2_X1 port map( A1 => n7581, A2 => n8297, ZN => n383);
   U2227 : AOI22_X1 port map( A1 => n19166, A2 => n19165, B1 => n386, B2 => 
                           n19948, ZN => n19167);
   U2228 : NAND2_X1 port map( A1 => n19161, A2 => n150, ZN => n386);
   U2229 : OR2_X2 port map( A1 => n1967, A2 => n7423, ZN => n9018);
   U2230 : NAND2_X1 port map( A1 => n439, A2 => n387, ZN => n15735);
   U2233 : INV_X1 port map( A => n12639, ZN => n390);
   U2234 : NAND2_X1 port map( A1 => n8682, A2 => n9149, ZN => n392);
   U2237 : NAND2_X1 port map( A1 => n1525, A2 => n15148, ZN => n15149);
   U2238 : OAI21_X1 port map( B1 => n9211, B2 => n263, A => n394, ZN => n8448);
   U2239 : NAND2_X1 port map( A1 => n9211, A2 => n8444, ZN => n394);
   U2241 : XNOR2_X1 port map( A => n395, B => n9787, ZN => n9789);
   U2242 : XNOR2_X1 port map( A => n9788, B => n10387, ZN => n395);
   U2243 : AOI21_X1 port map( B1 => n17982, B2 => n18238, A => n396, ZN => 
                           n3208);
   U2244 : INV_X1 port map( A => n17981, ZN => n396);
   U2246 : OAI22_X1 port map( A1 => n19385, A2 => n17221, B1 => n17218, B2 => 
                           n19383, ZN => n19387);
   U2247 : NAND3_X1 port map( A1 => n4739, A2 => n5059, A3 => n5060, ZN => 
                           n4102);
   U2248 : OR2_X2 port map( A1 => n4103, A2 => n4104, ZN => n5985);
   U2250 : OR2_X1 port map( A1 => n8296, A2 => n8299, ZN => n397);
   U2251 : NOR2_X1 port map( A1 => n20000, A2 => n9107, ZN => n8555);
   U2252 : AOI21_X2 port map( B1 => n12506, B2 => n9887, A => n398, ZN => 
                           n13746);
   U2253 : OAI22_X1 port map( A1 => n9885, A2 => n12506, B1 => n9886, B2 => 
                           n12008, ZN => n398);
   U2254 : OAI21_X2 port map( B1 => n8130, B2 => n8129, A => n399, ZN => n9999)
                           ;
   U2255 : OAI211_X1 port map( C1 => n8127, C2 => n8128, A => n1651, B => n8889
                           , ZN => n399);
   U2256 : NOR2_X2 port map( A1 => n8724, A2 => n8725, ZN => n10273);
   U2257 : MUX2_X1 port map( A => n7724, B => n8161, S => n8160, Z => n8164);
   U2258 : NAND2_X1 port map( A1 => n7855, A2 => n8157, ZN => n8160);
   U2259 : NOR2_X1 port map( A1 => n5583, A2 => n5582, ZN => n5584);
   U2260 : NAND2_X1 port map( A1 => n3959, A2 => n3960, ZN => n5583);
   U2262 : NAND2_X1 port map( A1 => n15373, A2 => n548, ZN => n16996);
   U2263 : XNOR2_X1 port map( A => n400, B => n18985, ZN => Ciphertext(108));
   U2264 : NAND2_X1 port map( A1 => n2050, A2 => n18983, ZN => n400);
   U2265 : OAI211_X1 port map( C1 => n6439, C2 => n8128, A => n401, B => n9090,
                           ZN => n6440);
   U2268 : NAND3_X1 port map( A1 => n1118, A2 => n17913, A3 => n17914, ZN => 
                           n403);
   U2270 : OAI21_X1 port map( B1 => n650, B2 => n11423, A => n2440, ZN => 
                           n12524);
   U2271 : XNOR2_X1 port map( A => n403, B => n302, ZN => Ciphertext(24));
   U2272 : OR2_X1 port map( A1 => n4306, A2 => n4305, ZN => n4004);
   U2273 : XNOR2_X1 port map( A => n405, B => n17783, ZN => Ciphertext(87));
   U2274 : NAND3_X1 port map( A1 => n2219, A2 => n2177, A3 => n17782, ZN => 
                           n405);
   U2277 : NAND2_X1 port map( A1 => n3770, A2 => n410, ZN => n409);
   U2278 : OR2_X1 port map( A1 => n4233, A2 => n4856, ZN => n410);
   U2279 : NAND3_X1 port map( A1 => n412, A2 => n4153, A3 => n4607, ZN => n4154
                           );
   U2280 : NAND2_X1 port map( A1 => n4546, A2 => n4603, ZN => n412);
   U2281 : NOR2_X1 port map( A1 => n5581, A2 => n733, ZN => n5000);
   U2285 : OAI21_X1 port map( B1 => n415, B2 => n249, A => n12002, ZN => n2260)
                           ;
   U2287 : NAND3_X1 port map( A1 => n1687, A2 => n2465, A3 => n5145, ZN => 
                           n6674);
   U2288 : NAND2_X1 port map( A1 => n416, A2 => n7963, ZN => n7966);
   U2289 : NAND2_X1 port map( A1 => n208, A2 => n7801, ZN => n416);
   U2290 : OAI21_X1 port map( B1 => n14131, B2 => n15606, A => n417, ZN => 
                           n14139);
   U2293 : OR2_X1 port map( A1 => n10673, A2 => n10194, ZN => n11341);
   U2294 : NAND3_X2 port map( A1 => n419, A2 => n3107, A3 => n3106, ZN => 
                           n10229);
   U2296 : NAND3_X1 port map( A1 => n14728, A2 => n14731, A3 => n14224, ZN => 
                           n420);
   U2297 : OAI211_X1 port map( C1 => n12347, C2 => n201, A => n421, B => n12346
                           , ZN => n12348);
   U2298 : NAND2_X1 port map( A1 => n12345, A2 => n201, ZN => n421);
   U2299 : OR3_X1 port map( A1 => n3366, A2 => n14666, A3 => n14663, ZN => 
                           n14037);
   U2300 : NAND2_X1 port map( A1 => n806, A2 => n5495, ZN => n805);
   U2301 : AND3_X2 port map( A1 => n422, A2 => n1307, A3 => n1306, ZN => n13275
                           );
   U2302 : NAND2_X1 port map( A1 => n10366, A2 => n11451, ZN => n422);
   U2303 : NAND2_X1 port map( A1 => n9028, A2 => n9031, ZN => n9034);
   U2304 : NAND2_X1 port map( A1 => n2504, A2 => n8545, ZN => n544);
   U2305 : OAI21_X1 port map( B1 => n8263, B2 => n8262, A => n423, ZN => n8265)
                           ;
   U2306 : NAND2_X1 port map( A1 => n8263, A2 => n895, ZN => n423);
   U2307 : NAND3_X1 port map( A1 => n10705, A2 => n10708, A3 => n10953, ZN => 
                           n2045);
   U2308 : NAND2_X1 port map( A1 => n20470, A2 => n10952, ZN => n10705);
   U2309 : NAND2_X1 port map( A1 => n18101, A2 => n19774, ZN => n424);
   U2310 : NAND2_X1 port map( A1 => n14998, A2 => n15835, ZN => n15001);
   U2311 : OAI211_X2 port map( C1 => n12515, C2 => n1305, A => n2491, B => 
                           n1304, ZN => n13136);
   U2312 : XNOR2_X2 port map( A => n425, B => Key(93), ZN => n5093);
   U2313 : INV_X1 port map( A => Plaintext(93), ZN => n425);
   U2319 : NAND2_X1 port map( A1 => n7418, A2 => n19901, ZN => n429);
   U2320 : NAND2_X1 port map( A1 => n9243, A2 => n430, ZN => n8715);
   U2321 : NAND2_X1 port map( A1 => n431, A2 => n1777, ZN => n430);
   U2323 : OR2_X1 port map( A1 => n7584, A2 => n2548, ZN => n7588);
   U2324 : OR2_X1 port map( A1 => n4667, A2 => n19688, ZN => n4672);
   U2325 : AND2_X1 port map( A1 => n18094, A2 => n18096, ZN => n759);
   U2326 : NAND3_X1 port map( A1 => n4026, A2 => n4027, A3 => n20464, ZN => 
                           n432);
   U2327 : NAND2_X1 port map( A1 => n4029, A2 => n4698, ZN => n434);
   U2328 : NAND2_X1 port map( A1 => n15564, A2 => n232, ZN => n435);
   U2329 : AOI22_X1 port map( A1 => n14741, A2 => n14740, B1 => n14739, B2 => 
                           n14738, ZN => n14952);
   U2330 : NAND2_X1 port map( A1 => n9163, A2 => n437, ZN => n436);
   U2331 : INV_X1 port map( A => n12430, ZN => n3649);
   U2332 : XNOR2_X1 port map( A => n6415, B => n6414, ZN => n7750);
   U2333 : OR2_X1 port map( A1 => n8353, A2 => n8352, ZN => n823);
   U2335 : OAI211_X1 port map( C1 => n1334, C2 => n803, A => n1333, B => n3454,
                           ZN => n9748);
   U2336 : NAND2_X1 port map( A1 => n747, A2 => n16126, ZN => n439);
   U2337 : INV_X1 port map( A => n14410, ZN => n14132);
   U2338 : AND2_X1 port map( A1 => n236, A2 => n14410, ZN => n14223);
   U2340 : OAI211_X1 port map( C1 => n18472, C2 => n18471, A => n18470, B => 
                           n440, ZN => n18474);
   U2341 : NAND3_X1 port map( A1 => n18466, A2 => n20110, A3 => n20148, ZN => 
                           n440);
   U2342 : OR2_X1 port map( A1 => n20451, A2 => n14410, ZN => n14134);
   U2343 : NAND3_X1 port map( A1 => n11275, A2 => n10684, A3 => n11271, ZN => 
                           n11249);
   U2346 : AND2_X1 port map( A1 => n11428, A2 => n11106, ZN => n10769);
   U2347 : NAND2_X1 port map( A1 => n17817, A2 => n227, ZN => n443);
   U2348 : NAND2_X1 port map( A1 => n18966, A2 => n18968, ZN => n17817);
   U2349 : NAND2_X1 port map( A1 => n18965, A2 => n20127, ZN => n444);
   U2352 : NAND2_X1 port map( A1 => n5316, A2 => n3533, ZN => n446);
   U2353 : NAND2_X2 port map( A1 => n447, A2 => n7004, ZN => n9046);
   U2355 : NAND3_X1 port map( A1 => n16010, A2 => n15333, A3 => n13968, ZN => 
                           n527);
   U2356 : OAI21_X1 port map( B1 => n5078, B2 => n5077, A => n448, ZN => n5503)
                           ;
   U2357 : NAND2_X1 port map( A1 => n2162, A2 => n11418, ZN => n2161);
   U2358 : NAND3_X1 port map( A1 => n12685, A2 => n1091, A3 => n12686, ZN => 
                           n1092);
   U2359 : OR3_X1 port map( A1 => n7754, A2 => n7530, A3 => n7903, ZN => n644);
   U2360 : NAND2_X1 port map( A1 => n7998, A2 => n1425, ZN => n449);
   U2363 : NAND2_X1 port map( A1 => n8256, A2 => n8258, ZN => n7726);
   U2365 : NAND2_X1 port map( A1 => n3133, A2 => n3134, ZN => n2680);
   U2366 : INV_X1 port map( A => n15094, ZN => n451);
   U2367 : AND2_X2 port map( A1 => n451, A2 => n149, ZN => n17035);
   U2369 : NAND3_X1 port map( A1 => n4867, A2 => n2072, A3 => n453, ZN => n452)
                           ;
   U2370 : NAND2_X1 port map( A1 => n11712, A2 => n454, ZN => n13138);
   U2371 : OR2_X1 port map( A1 => n11713, A2 => n12155, ZN => n454);
   U2372 : OAI21_X1 port map( B1 => n10789, B2 => n10788, A => n10787, ZN => 
                           n12636);
   U2374 : NAND2_X1 port map( A1 => n4632, A2 => n455, ZN => n5179);
   U2375 : OR2_X1 port map( A1 => n8411, A2 => n655, ZN => n9183);
   U2376 : NOR2_X1 port map( A1 => n3468, A2 => n5985, ZN => n5438);
   U2377 : XNOR2_X1 port map( A => n10600, B => n9860, ZN => n550);
   U2378 : XNOR2_X2 port map( A => n7214, B => n7215, ZN => n8004);
   U2379 : NAND2_X1 port map( A1 => n4652, A2 => n4867, ZN => n3562);
   U2382 : NAND3_X1 port map( A1 => n11962, A2 => n2140, A3 => n2139, ZN => 
                           n458);
   U2385 : INV_X1 port map( A => n8289, ZN => n462);
   U2386 : NAND2_X1 port map( A1 => n7468, A2 => n7807, ZN => n463);
   U2387 : NAND2_X1 port map( A1 => n1658, A2 => n464, ZN => n9011);
   U2389 : OAI211_X2 port map( C1 => n7819, C2 => n7818, A => n7817, B => n465,
                           ZN => n8895);
   U2390 : NAND3_X1 port map( A1 => n466, A2 => n8379, A3 => n8378, ZN => n8445
                           );
   U2391 : NAND3_X1 port map( A1 => n8371, A2 => n8369, A3 => n8370, ZN => n466
                           );
   U2393 : NOR2_X2 port map( A1 => n7490, A2 => n467, ZN => n9122);
   U2394 : AOI21_X1 port map( B1 => n7489, B2 => n7488, A => n22, ZN => n467);
   U2395 : XNOR2_X1 port map( A => n20018, B => n13527, ZN => n12367);
   U2397 : OAI21_X1 port map( B1 => n5345, B2 => n6139, A => n469, ZN => n6724)
                           ;
   U2398 : NAND2_X1 port map( A1 => n5343, A2 => n5344, ZN => n469);
   U2399 : XNOR2_X1 port map( A => n470, B => n790, ZN => n8777);
   U2400 : XNOR2_X1 port map( A => n8776, B => n10030, ZN => n470);
   U2401 : NAND2_X1 port map( A1 => n5593, A2 => n5590, ZN => n5591);
   U2402 : NAND2_X1 port map( A1 => n8950, A2 => n8603, ZN => n9367);
   U2403 : NAND2_X1 port map( A1 => n2070, A2 => n1882, ZN => n3981);
   U2405 : NAND2_X1 port map( A1 => n472, A2 => n471, ZN => n4001);
   U2406 : NAND2_X1 port map( A1 => n3993, A2 => n6068, ZN => n471);
   U2407 : NAND2_X1 port map( A1 => n3992, A2 => n473, ZN => n472);
   U2408 : NAND2_X1 port map( A1 => n12473, A2 => n12142, ZN => n12393);
   U2409 : AOI21_X2 port map( B1 => n8351, B2 => n7549, A => n2778, ZN => n8960
                           );
   U2410 : AOI22_X1 port map( A1 => n9369, A2 => n904, B1 => n9370, B2 => n9371
                           , ZN => n9373);
   U2412 : NOR2_X1 port map( A1 => n14590, A2 => n19781, ZN => n474);
   U2414 : AOI22_X1 port map( A1 => n3250, A2 => n8141, B1 => n8270, B2 => 
                           n8350, ZN => n475);
   U2415 : NAND2_X1 port map( A1 => n12591, A2 => n12589, ZN => n12596);
   U2416 : NAND2_X1 port map( A1 => n15395, A2 => n14990, ZN => n3247);
   U2417 : OR2_X1 port map( A1 => n12658, A2 => n15657, ZN => n546);
   U2422 : NAND2_X1 port map( A1 => n7529, A2 => n274, ZN => n477);
   U2423 : NOR2_X1 port map( A1 => n13318, A2 => n478, ZN => n15672);
   U2426 : NOR2_X1 port map( A1 => n479, A2 => n17748, ZN => n780);
   U2427 : AND2_X1 port map( A1 => n18028, A2 => n17749, ZN => n479);
   U2428 : OAI22_X1 port map( A1 => n10688, A2 => n19851, B1 => n9547, B2 => 
                           n11277, ZN => n11276);
   U2429 : OAI211_X1 port map( C1 => n5745, C2 => n5741, A => n20509, B => n481
                           , ZN => n480);
   U2430 : NAND2_X1 port map( A1 => n5741, A2 => n286, ZN => n481);
   U2431 : XNOR2_X1 port map( A => n19844, B => n16429, ZN => n14163);
   U2435 : NAND2_X1 port map( A1 => n2541, A2 => n14277, ZN => n1409);
   U2441 : OAI21_X1 port map( B1 => n2320, B2 => n12147, A => n12149, ZN => 
                           n485);
   U2443 : NAND2_X1 port map( A1 => n486, A2 => n4334, ZN => n6165);
   U2444 : NAND2_X1 port map( A1 => n4333, A2 => n5632, ZN => n486);
   U2445 : NAND2_X1 port map( A1 => n15550, A2 => n15056, ZN => n14979);
   U2448 : NAND2_X1 port map( A1 => n11660, A2 => n11951, ZN => n487);
   U2449 : NAND2_X1 port map( A1 => n19248, A2 => n3345, ZN => n17667);
   U2450 : NOR2_X2 port map( A1 => n13998, A2 => n13999, ZN => n15701);
   U2451 : NAND2_X1 port map( A1 => n8263, A2 => n8262, ZN => n8106);
   U2453 : NAND2_X1 port map( A1 => n490, A2 => n489, ZN => n18861);
   U2454 : NAND2_X1 port map( A1 => n18860, A2 => n216, ZN => n489);
   U2455 : NAND2_X1 port map( A1 => n18859, A2 => n18869, ZN => n490);
   U2457 : NAND2_X1 port map( A1 => n492, A2 => n491, ZN => n11947);
   U2458 : NAND2_X1 port map( A1 => n11946, A2 => n20457, ZN => n492);
   U2459 : NAND2_X1 port map( A1 => n6272, A2 => n494, ZN => n493);
   U2461 : NAND3_X1 port map( A1 => n1812, A2 => n11452, A3 => n11455, ZN => 
                           n10733);
   U2462 : XNOR2_X2 port map( A => n16759, B => n16758, ZN => n18954);
   U2464 : NAND3_X1 port map( A1 => n14675, A2 => n13981, A3 => n14674, ZN => 
                           n687);
   U2465 : OAI22_X1 port map( A1 => n15475, A2 => n15244, B1 => n15656, B2 => 
                           n15243, ZN => n14859);
   U2466 : NAND2_X1 port map( A1 => n15658, A2 => n15474, ZN => n15244);
   U2467 : INV_X1 port map( A => n496, ZN => n495);
   U2468 : OAI21_X1 port map( B1 => n5713, B2 => n5985, A => n5712, ZN => n496)
                           ;
   U2469 : NAND2_X1 port map( A1 => n5710, A2 => n5986, ZN => n497);
   U2470 : NAND2_X1 port map( A1 => n12606, A2 => n3305, ZN => n11628);
   U2471 : NAND3_X2 port map( A1 => n1893, A2 => n1892, A3 => n10892, ZN => 
                           n12606);
   U2475 : INV_X1 port map( A => n8070, ZN => n8204);
   U2476 : NAND2_X1 port map( A1 => n4633, A2 => n20487, ZN => n4156);
   U2477 : NOR2_X1 port map( A1 => n12528, A2 => n12525, ZN => n12526);
   U2478 : NAND2_X1 port map( A1 => n182, A2 => n12523, ZN => n12525);
   U2479 : AND2_X1 port map( A1 => n1907, A2 => n17886, ZN => n17600);
   U2480 : XNOR2_X1 port map( A => n13711, B => n13659, ZN => n12079);
   U2483 : AND2_X1 port map( A1 => n11154, A2 => n1580, ZN => n532);
   U2486 : NOR3_X1 port map( A1 => n10979, A2 => n19506, A3 => n10982, ZN => 
                           n10984);
   U2487 : XNOR2_X1 port map( A => n16568, B => n17433, ZN => n17135);
   U2490 : INV_X1 port map( A => n11168, ZN => n11533);
   U2491 : NAND2_X1 port map( A1 => n11337, A2 => n11267, ZN => n755);
   U2492 : XNOR2_X1 port map( A => n657, B => n18177, ZN => n6832);
   U2493 : NAND2_X1 port map( A1 => n4405, A2 => n5093, ZN => n5096);
   U2494 : NAND2_X1 port map( A1 => n2234, A2 => n2235, ZN => n11922);
   U2497 : AND2_X1 port map( A1 => n9559, A2 => n19779, ZN => n11287);
   U2498 : NAND2_X1 port map( A1 => n4901, A2 => n4492, ZN => n4494);
   U2499 : NAND2_X1 port map( A1 => n504, A2 => n502, ZN => n1725);
   U2501 : NAND2_X1 port map( A1 => n7536, A2 => n505, ZN => n504);
   U2503 : NAND3_X1 port map( A1 => n9368, A2 => n8953, A3 => n8952, ZN => n506
                           );
   U2505 : OAI22_X1 port map( A1 => n3598, A2 => n3167, B1 => n5107, B2 => n507
                           , ZN => n3166);
   U2506 : NAND2_X1 port map( A1 => n5099, A2 => n4048, ZN => n507);
   U2507 : NAND2_X1 port map( A1 => n1338, A2 => n11574, ZN => n11576);
   U2508 : NAND2_X1 port map( A1 => n5326, A2 => n508, ZN => n4284);
   U2509 : NAND2_X1 port map( A1 => n510, A2 => n509, ZN => n12275);
   U2511 : NAND2_X1 port map( A1 => n11551, A2 => n11550, ZN => n510);
   U2512 : NAND2_X1 port map( A1 => n12030, A2 => n12304, ZN => n512);
   U2513 : NAND2_X1 port map( A1 => n12031, A2 => n11782, ZN => n513);
   U2516 : NAND2_X1 port map( A1 => n14506, A2 => n14305, ZN => n13507);
   U2518 : NAND2_X1 port map( A1 => n19113, A2 => n19112, ZN => n19120);
   U2520 : OAI21_X1 port map( B1 => n5951, B2 => n5950, A => n5949, ZN => n515)
                           ;
   U2522 : OR3_X1 port map( A1 => n5796, A2 => n5795, A3 => n5300, ZN => n5794)
                           ;
   U2523 : NAND2_X1 port map( A1 => n551, A2 => n516, ZN => n13231);
   U2524 : NAND2_X1 port map( A1 => n11624, A2 => n12441, ZN => n516);
   U2526 : NAND2_X1 port map( A1 => n5407, A2 => n517, ZN => n6404);
   U2527 : OR2_X1 port map( A1 => n5409, A2 => n5408, ZN => n517);
   U2528 : OAI21_X1 port map( B1 => n239, B2 => n19781, A => n518, ZN => n14200
                           );
   U2529 : NAND2_X1 port map( A1 => n19781, A2 => n14811, ZN => n518);
   U2531 : NAND3_X2 port map( A1 => n2452, A2 => n537, A3 => n536, ZN => n10247
                           );
   U2533 : NAND2_X1 port map( A1 => n2373, A2 => n921, ZN => n519);
   U2534 : NAND2_X1 port map( A1 => n520, A2 => n828, ZN => n827);
   U2535 : NAND2_X1 port map( A1 => n575, A2 => n829, ZN => n520);
   U2536 : NAND2_X1 port map( A1 => n522, A2 => n521, ZN => n10630);
   U2537 : NAND2_X1 port map( A1 => n12325, A2 => n12514, ZN => n522);
   U2539 : INV_X1 port map( A => n15333, ZN => n1817);
   U2540 : NAND2_X1 port map( A1 => n15879, A2 => n15153, ZN => n15333);
   U2542 : OR2_X2 port map( A1 => n9554, A2 => n9553, ZN => n11598);
   U2543 : NOR2_X1 port map( A1 => n12974, A2 => n3820, ZN => n12975);
   U2545 : NAND2_X1 port map( A1 => n7797, A2 => n7466, ZN => n7963);
   U2547 : NAND2_X1 port map( A1 => n1090, A2 => n14837, ZN => n14840);
   U2548 : OAI211_X2 port map( C1 => n10317, C2 => n10316, A => n525, B => n524
                           , ZN => n13352);
   U2549 : NAND2_X1 port map( A1 => n10313, A2 => n12336, ZN => n524);
   U2550 : NAND2_X1 port map( A1 => n10315, A2 => n10314, ZN => n525);
   U2551 : XNOR2_X1 port map( A => n526, B => n2145, ZN => n11113);
   U2552 : XNOR2_X1 port map( A => n10371, B => n10370, ZN => n526);
   U2553 : INV_X1 port map( A => n4714, ZN => n5097);
   U2554 : OAI22_X1 port map( A1 => n3804, A2 => n5891, B1 => n20670, B2 => 
                           n3249, ZN => n5893);
   U2555 : NAND2_X1 port map( A1 => n2217, A2 => n3662, ZN => n1989);
   U2558 : NAND2_X1 port map( A1 => n527, A2 => n15154, ZN => n15155);
   U2560 : XNOR2_X2 port map( A => n9736, B => n9737, ZN => n11395);
   U2561 : OR2_X1 port map( A1 => n5093, A2 => n4405, ZN => n4782);
   U2562 : NOR2_X1 port map( A1 => n12366, A2 => n12365, ZN => n915);
   U2564 : OAI22_X1 port map( A1 => n8944, A2 => n8945, B1 => n8947, B2 => 
                           n8946, ZN => n528);
   U2565 : NAND2_X1 port map( A1 => n5093, A2 => n5098, ZN => n4714);
   U2566 : AOI21_X2 port map( B1 => n15001, B2 => n15831, A => n15000, ZN => 
                           n16706);
   U2567 : INV_X1 port map( A => n14626, ZN => n14192);
   U2568 : XNOR2_X1 port map( A => n11901, B => n11900, ZN => n14626);
   U2569 : OAI21_X1 port map( B1 => n4349, B2 => n301, A => n4540, ZN => n3932)
                           ;
   U2570 : NAND2_X1 port map( A1 => n17977, A2 => n17758, ZN => n17762);
   U2572 : NAND3_X1 port map( A1 => n637, A2 => n9054, A3 => n9306, ZN => n529)
                           ;
   U2574 : AOI21_X1 port map( B1 => n3056, B2 => n13682, A => n13963, ZN => 
                           n530);
   U2575 : NAND2_X1 port map( A1 => n5394, A2 => n5395, ZN => n5326);
   U2576 : NAND2_X1 port map( A1 => n4167, A2 => n531, ZN => n4017);
   U2577 : OR3_X1 port map( A1 => n17480, A2 => n20354, A3 => n17479, ZN => 
                           n17485);
   U2578 : AOI21_X2 port map( B1 => n1971, B2 => n3382, A => n532, ZN => n12280
                           );
   U2579 : NAND2_X1 port map( A1 => n534, A2 => n533, ZN => n5253);
   U2580 : NAND2_X1 port map( A1 => n5252, A2 => n5323, ZN => n534);
   U2581 : NAND2_X1 port map( A1 => n3457, A2 => n15245, ZN => n12663);
   U2582 : NAND2_X1 port map( A1 => n8290, A2 => n20189, ZN => n7370);
   U2583 : OAI21_X1 port map( B1 => n5792, B2 => n1026, A => n535, ZN => n5157)
                           ;
   U2584 : NAND2_X1 port map( A1 => n5792, A2 => n5156, ZN => n535);
   U2585 : NAND2_X1 port map( A1 => n8800, A2 => n8799, ZN => n536);
   U2586 : NAND2_X1 port map( A1 => n908, A2 => n8798, ZN => n537);
   U2587 : NAND2_X1 port map( A1 => n539, A2 => n16364, ZN => n18556);
   U2588 : OAI21_X1 port map( B1 => n17966, B2 => n16363, A => n18112, ZN => 
                           n539);
   U2589 : NOR2_X1 port map( A1 => n8468, A2 => n8467, ZN => n9647);
   U2590 : OAI211_X1 port map( C1 => n3373, C2 => n20424, A => n2402, B => 
                           n14020, ZN => n688);
   U2591 : XNOR2_X1 port map( A => n540, B => n12679, ZN => n12681);
   U2592 : XNOR2_X1 port map( A => n12680, B => n13018, ZN => n540);
   U2593 : NAND2_X1 port map( A1 => n10896, A2 => n10745, ZN => n10059);
   U2596 : NAND2_X1 port map( A1 => n12534, A2 => n12162, ZN => n11804);
   U2597 : NOR2_X1 port map( A1 => n8547, A2 => n8546, ZN => n872);
   U2598 : NAND2_X1 port map( A1 => n544, A2 => n543, ZN => n8546);
   U2599 : NAND2_X1 port map( A1 => n8544, A2 => n2749, ZN => n543);
   U2600 : INV_X1 port map( A => n11133, ZN => n650);
   U2602 : NAND2_X1 port map( A1 => n4622, A2 => n4285, ZN => n4167);
   U2603 : NOR2_X2 port map( A1 => n14560, A2 => n14561, ZN => n15644);
   U2606 : AND2_X2 port map( A1 => n1132, A2 => n1133, ZN => n12359);
   U2607 : NAND3_X1 port map( A1 => n749, A2 => n748, A3 => n4610, ZN => n762);
   U2608 : NAND2_X1 port map( A1 => n20146, A2 => n9204, ZN => n771);
   U2610 : INV_X1 port map( A => Plaintext(188), ZN => n547);
   U2611 : NAND2_X1 port map( A1 => n549, A2 => n232, ZN => n548);
   U2612 : INV_X1 port map( A => n15374, ZN => n549);
   U2614 : NAND2_X1 port map( A1 => n11623, A2 => n12442, ZN => n552);
   U2615 : NAND2_X1 port map( A1 => n11622, A2 => n1522, ZN => n553);
   U2616 : AOI21_X1 port map( B1 => n11540, B2 => n11541, A => n11539, ZN => 
                           n11542);
   U2618 : NAND2_X1 port map( A1 => n5708, A2 => n5815, ZN => n5816);
   U2619 : NAND2_X1 port map( A1 => n557, A2 => n554, ZN => n4273);
   U2620 : NAND2_X1 port map( A1 => n555, A2 => n4765, ZN => n554);
   U2621 : NAND2_X1 port map( A1 => n4764, A2 => n556, ZN => n555);
   U2622 : NAND2_X1 port map( A1 => n4270, A2 => n19788, ZN => n557);
   U2623 : XOR2_X1 port map( A => n7087, B => n7316, Z => n826);
   U2625 : NOR2_X1 port map( A1 => n3247, A2 => n15306, ZN => n15062);
   U2626 : NAND2_X1 port map( A1 => n17882, A2 => n17881, ZN => n558);
   U2627 : NAND2_X1 port map( A1 => n17883, A2 => n222, ZN => n559);
   U2628 : NAND3_X1 port map( A1 => n593, A2 => n4437, A3 => n4438, ZN => n1919
                           );
   U2629 : NAND2_X1 port map( A1 => n562, A2 => n560, ZN => n17698);
   U2630 : NAND2_X1 port map( A1 => n17694, A2 => n17819, ZN => n560);
   U2631 : NAND2_X1 port map( A1 => n17693, A2 => n935, ZN => n562);
   U2633 : NAND3_X1 port map( A1 => n564, A2 => n773, A3 => n3087, ZN => n15059
                           );
   U2635 : OAI211_X1 port map( C1 => n15462, C2 => n1458, A => n15351, B => 
                           n15352, ZN => n565);
   U2637 : OR2_X1 port map( A1 => n2867, A2 => n2869, ZN => n566);
   U2638 : NAND2_X1 port map( A1 => n4707, A2 => n4706, ZN => n567);
   U2640 : NAND2_X1 port map( A1 => n1535, A2 => n619, ZN => n1534);
   U2641 : NOR2_X1 port map( A1 => n569, A2 => n568, ZN => n5843);
   U2642 : NAND2_X1 port map( A1 => n572, A2 => n570, ZN => n12597);
   U2643 : NAND2_X1 port map( A1 => n571, A2 => n12595, ZN => n570);
   U2644 : NAND2_X1 port map( A1 => n12593, A2 => n20430, ZN => n571);
   U2645 : NAND2_X1 port map( A1 => n12596, A2 => n11637, ZN => n572);
   U2646 : NAND2_X1 port map( A1 => n8851, A2 => n9038, ZN => n1979);
   U2648 : OAI211_X1 port map( C1 => n2600, C2 => n11977, A => n574, B => n250,
                           ZN => n11414);
   U2649 : NAND2_X1 port map( A1 => n2600, A2 => n12545, ZN => n574);
   U2650 : XNOR2_X1 port map( A => n638, B => n6732, ZN => n3484);
   U2651 : OR2_X1 port map( A1 => n291, A2 => n5073, ZN => n575);
   U2653 : NAND2_X1 port map( A1 => n9098, A2 => n10646, ZN => n576);
   U2654 : NAND2_X1 port map( A1 => n1959, A2 => n20149, ZN => n578);
   U2658 : XNOR2_X1 port map( A => n581, B => n295, ZN => Ciphertext(60));
   U2659 : NAND3_X1 port map( A1 => n582, A2 => n18641, A3 => n18640, ZN => 
                           n581);
   U2661 : NAND2_X1 port map( A1 => n19745, A2 => n583, ZN => n18639);
   U2663 : NAND2_X1 port map( A1 => n5760, A2 => n7421, ZN => n586);
   U2664 : NAND2_X1 port map( A1 => n18441, A2 => n18466, ZN => n18446);
   U2665 : XNOR2_X2 port map( A => n587, B => n13076, ZN => n14514);
   U2666 : XNOR2_X1 port map( A => n2200, B => n13077, ZN => n587);
   U2667 : NAND3_X1 port map( A1 => n243, A2 => n12537, A3 => n12534, ZN => 
                           n2328);
   U2669 : NAND2_X1 port map( A1 => n608, A2 => n20516, ZN => n607);
   U2670 : NAND2_X1 port map( A1 => n8852, A2 => n9038, ZN => n589);
   U2671 : NAND2_X1 port map( A1 => n8849, A2 => n591, ZN => n590);
   U2672 : INV_X1 port map( A => n9038, ZN => n591);
   U2673 : NAND2_X1 port map( A1 => n592, A2 => n8492, ZN => n7701);
   U2675 : NAND3_X1 port map( A1 => n5429, A2 => n1776, A3 => n5790, ZN => 
                           n2956);
   U2676 : NAND2_X1 port map( A1 => n9009, A2 => n9007, ZN => n1671);
   U2677 : OAI21_X1 port map( B1 => n4807, B2 => n4802, A => n4801, ZN => n593)
                           ;
   U2678 : XNOR2_X1 port map( A => n594, B => n17365, ZN => Ciphertext(8));
   U2680 : NAND2_X1 port map( A1 => n3455, A2 => n3456, ZN => n596);
   U2681 : NAND2_X1 port map( A1 => n1106, A2 => n3388, ZN => n18394);
   U2682 : OAI21_X2 port map( B1 => n11679, B2 => n12500, A => n1149, ZN => 
                           n12979);
   U2683 : AOI22_X1 port map( A1 => n20111, A2 => n18384, B1 => n20611, B2 => 
                           n18376, ZN => n18393);
   U2684 : NAND3_X1 port map( A1 => n4609, A2 => n4613, A3 => n4177, ZN => 
                           n3109);
   U2685 : NAND2_X1 port map( A1 => n14005, A2 => n2304, ZN => n14119);
   U2686 : AND2_X2 port map( A1 => n751, A2 => n752, ZN => n15696);
   U2687 : NAND2_X1 port map( A1 => n5444, A2 => n5641, ZN => n4179);
   U2688 : NAND3_X2 port map( A1 => n3110, A2 => n3108, A3 => n4178, ZN => 
                           n5444);
   U2689 : INV_X1 port map( A => n598, ZN => n597);
   U2691 : NAND2_X1 port map( A1 => n800, A2 => n9363, ZN => n599);
   U2692 : NOR2_X1 port map( A1 => n20005, A2 => n20133, ZN => n750);
   U2693 : NAND2_X1 port map( A1 => n17876, A2 => n16308, ZN => n600);
   U2694 : OR2_X1 port map( A1 => n10808, A2 => n10259, ZN => n10809);
   U2695 : NAND2_X1 port map( A1 => n4750, A2 => n4204, ZN => n4558);
   U2697 : AOI22_X1 port map( A1 => n11266, A2 => n11265, B1 => n11335, B2 => 
                           n11267, ZN => n602);
   U2698 : OAI211_X2 port map( C1 => n14521, C2 => n14520, A => n15126, B => 
                           n15125, ZN => n15018);
   U2699 : NAND2_X1 port map( A1 => n14518, A2 => n14519, ZN => n15126);
   U2701 : NAND2_X1 port map( A1 => n4366, A2 => n290, ZN => n603);
   U2702 : NAND2_X1 port map( A1 => n605, A2 => n4365, ZN => n604);
   U2703 : NAND2_X1 port map( A1 => n4011, A2 => n4614, ZN => n605);
   U2704 : NAND2_X1 port map( A1 => n11671, A2 => n11672, ZN => n11676);
   U2706 : NAND2_X1 port map( A1 => n8330, A2 => n8331, ZN => n9861);
   U2707 : NAND2_X1 port map( A1 => n2238, A2 => n7643, ZN => n8603);
   U2709 : NOR2_X1 port map( A1 => n15896, A2 => n15536, ZN => n15539);
   U2710 : AOI22_X1 port map( A1 => n11735, A2 => n242, B1 => n13149, B2 => 
                           n20153, ZN => n11736);
   U2711 : NAND2_X1 port map( A1 => n10803, A2 => n191, ZN => n10804);
   U2712 : NAND2_X1 port map( A1 => n18645, A2 => n18656, ZN => n18282);
   U2713 : INV_X1 port map( A => n4615, ZN => n748);
   U2715 : INV_X1 port map( A => n11159, ZN => n608);
   U2717 : INV_X1 port map( A => n4931, ZN => n4977);
   U2718 : OAI21_X1 port map( B1 => n3877, B2 => n3876, A => n4931, ZN => n3878
                           );
   U2719 : NAND2_X1 port map( A1 => n4979, A2 => n4297, ZN => n4931);
   U2721 : NAND2_X1 port map( A1 => n17395, A2 => n18257, ZN => n611);
   U2722 : OR2_X1 port map( A1 => n18260, A2 => n18257, ZN => n612);
   U2725 : NAND2_X1 port map( A1 => n613, A2 => n4010, ZN => n3955);
   U2726 : NAND2_X1 port map( A1 => n4364, A2 => n4614, ZN => n613);
   U2728 : NAND2_X1 port map( A1 => n2682, A2 => n14599, ZN => n3532);
   U2729 : INV_X1 port map( A => n9602, ZN => n10289);
   U2730 : NAND2_X1 port map( A1 => n7624, A2 => n7625, ZN => n8741);
   U2731 : NAND4_X1 port map( A1 => n4636, A2 => n4634, A3 => n4637, A4 => 
                           n4635, ZN => n614);
   U2732 : NAND2_X1 port map( A1 => n5319, A2 => n5406, ZN => n615);
   U2733 : NAND2_X1 port map( A1 => n13924, A2 => n3599, ZN => n3254);
   U2736 : NAND2_X1 port map( A1 => n6042, A2 => n1214, ZN => n5308);
   U2737 : AND2_X2 port map( A1 => n687, A2 => n688, ZN => n15796);
   U2738 : NAND2_X1 port map( A1 => n4616, A2 => n748, ZN => n617);
   U2739 : NAND2_X1 port map( A1 => n3715, A2 => n619, ZN => n618);
   U2740 : INV_X1 port map( A => n3717, ZN => n619);
   U2742 : MUX2_X1 port map( A => n4112, B => n5711, S => n5709, Z => n622);
   U2743 : AOI21_X1 port map( B1 => n1270, B2 => n3832, A => n20105, ZN => n623
                           );
   U2744 : NAND2_X1 port map( A1 => n624, A2 => n9346, ZN => n2168);
   U2745 : NAND2_X1 port map( A1 => n2170, A2 => n2169, ZN => n624);
   U2746 : NAND2_X1 port map( A1 => n4237, A2 => n4238, ZN => n2215);
   U2748 : NAND2_X1 port map( A1 => n15680, A2 => n15679, ZN => n625);
   U2749 : NAND2_X1 port map( A1 => n15681, A2 => n15682, ZN => n626);
   U2750 : NOR2_X1 port map( A1 => n152, A2 => n628, ZN => n16460);
   U2751 : NAND2_X1 port map( A1 => n630, A2 => n629, ZN => n3681);
   U2752 : INV_X1 port map( A => n8017, ZN => n630);
   U2753 : NAND2_X1 port map( A1 => n631, A2 => n14800, ZN => n14211);
   U2754 : XNOR2_X2 port map( A => n12249, B => n12248, ZN => n14800);
   U2755 : INV_X1 port map( A => n3440, ZN => n631);
   U2756 : NAND3_X1 port map( A1 => n252, A2 => n12179, A3 => n20427, ZN => 
                           n1980);
   U2757 : XNOR2_X1 port map( A => n735, B => n9478, ZN => n9551);
   U2758 : NAND3_X1 port map( A1 => n19742, A2 => n1089, A3 => n14501, ZN => 
                           n13053);
   U2759 : NAND2_X1 port map( A1 => n4807, A2 => n633, ZN => n4699);
   U2760 : AND2_X1 port map( A1 => n5087, A2 => n20202, ZN => n633);
   U2763 : NAND2_X1 port map( A1 => n16579, A2 => n635, ZN => n634);
   U2765 : NAND2_X1 port map( A1 => n1751, A2 => n9313, ZN => n637);
   U2766 : XNOR2_X1 port map( A => n6731, B => n6730, ZN => n638);
   U2767 : NAND2_X1 port map( A1 => n14731, A2 => n14729, ZN => n14137);
   U2768 : NAND2_X1 port map( A1 => n3086, A2 => n5602, ZN => n5485);
   U2773 : AND2_X2 port map( A1 => n5245, A2 => n5244, ZN => n5249);
   U2774 : NAND2_X1 port map( A1 => n7904, A2 => n7754, ZN => n3272);
   U2775 : NAND2_X1 port map( A1 => n7903, A2 => n20166, ZN => n7904);
   U2776 : OAI211_X2 port map( C1 => n7758, C2 => n7757, A => n7756, B => n644,
                           ZN => n8657);
   U2780 : NAND2_X1 port map( A1 => n10069, A2 => n11548, ZN => n646);
   U2781 : INV_X1 port map( A => n11548, ZN => n647);
   U2782 : NAND2_X1 port map( A1 => n11544, A2 => n10760, ZN => n648);
   U2783 : AND2_X1 port map( A1 => n205, A2 => n11133, ZN => n10830);
   U2784 : NAND2_X1 port map( A1 => n11052, A2 => n650, ZN => n11053);
   U2785 : NAND2_X1 port map( A1 => n11130, A2 => n650, ZN => n2106);
   U2788 : NAND2_X1 port map( A1 => n16685, A2 => n651, ZN => n654);
   U2792 : AOI22_X2 port map( A1 => n16686, A2 => n654, B1 => n19399, B2 => 
                           n16687, ZN => n19463);
   U2793 : NAND2_X1 port map( A1 => n654, A2 => n17654, ZN => n17659);
   U2794 : OR2_X2 port map( A1 => n5137, A2 => n5136, ZN => n655);
   U2795 : NOR2_X1 port map( A1 => n655, A2 => n9234, ZN => n8633);
   U2796 : NAND2_X1 port map( A1 => n19716, A2 => n655, ZN => n9236);
   U2797 : NAND3_X1 port map( A1 => n8411, A2 => n9234, A3 => n655, ZN => n6214
                           );
   U2798 : NAND2_X1 port map( A1 => n8630, A2 => n655, ZN => n8632);
   U2800 : NAND2_X1 port map( A1 => n656, A2 => n912, ZN => n2249);
   U2801 : MUX2_X1 port map( A => n14327, B => n14352, S => n14818, Z => n656);
   U2802 : XNOR2_X1 port map( A => n20224, B => n657, ZN => n6554);
   U2803 : XNOR2_X1 port map( A => n657, B => n18792, ZN => n6848);
   U2804 : XNOR2_X1 port map( A => n7206, B => n657, ZN => n6962);
   U2805 : XNOR2_X1 port map( A => n6743, B => n657, ZN => n7303);
   U2806 : INV_X1 port map( A => n2816, ZN => n660);
   U2807 : NOR2_X1 port map( A1 => n2816, A2 => n215, ZN => n658);
   U2808 : NAND3_X1 port map( A1 => n19278, A2 => n19269, A3 => n660, ZN => 
                           n19256);
   U2809 : MUX2_X1 port map( A => n19246, B => n19269, S => n2816, Z => n17682)
                           ;
   U2810 : NAND2_X1 port map( A1 => n19274, A2 => n2816, ZN => n659);
   U2811 : AOI21_X1 port map( B1 => n19275, B2 => n660, A => n20448, ZN => 
                           n19277);
   U2812 : OR2_X1 port map( A1 => n5021, A2 => n4277, ZN => n662);
   U2813 : NAND2_X1 port map( A1 => n4554, A2 => n663, ZN => n661);
   U2814 : NAND2_X1 port map( A1 => n5803, A2 => n5378, ZN => n5733);
   U2815 : AND2_X1 port map( A1 => n4734, A2 => n4555, ZN => n663);
   U2816 : MUX2_X1 port map( A => n666, B => n4568, S => n1391, Z => n664);
   U2817 : INV_X1 port map( A => n666, ZN => n665);
   U2818 : NAND2_X1 port map( A1 => n4563, A2 => n4754, ZN => n666);
   U2820 : NAND2_X1 port map( A1 => n7725, A2 => n7851, ZN => n667);
   U2822 : NAND2_X1 port map( A1 => n669, A2 => n8972, ZN => n3354);
   U2823 : OAI21_X1 port map( B1 => n8971, B2 => n9255, A => n8976, ZN => n669)
                           ;
   U2824 : NAND2_X1 port map( A1 => n671, A2 => n670, ZN => n8976);
   U2825 : INV_X1 port map( A => n9250, ZN => n671);
   U2826 : NAND2_X1 port map( A1 => n4731, A2 => n672, ZN => n4276);
   U2827 : NAND2_X1 port map( A1 => n4110, A2 => n5012, ZN => n5013);
   U2828 : NAND3_X1 port map( A1 => n5016, A2 => n4110, A3 => n4734, ZN => 
                           n4735);
   U2829 : NAND3_X1 port map( A1 => n5020, A2 => n5019, A3 => n673, ZN => n6027
                           );
   U2830 : OR2_X1 port map( A1 => n5021, A2 => n4110, ZN => n673);
   U2831 : XNOR2_X1 port map( A => n674, B => n18308, ZN => Ciphertext(98));
   U2832 : NAND2_X1 port map( A1 => n677, A2 => n675, ZN => n674);
   U2833 : NAND2_X1 port map( A1 => n676, A2 => n19988, ZN => n675);
   U2834 : MUX2_X1 port map( A => n20259, B => n18857, S => n20418, Z => n676);
   U2836 : NAND2_X1 port map( A1 => n678, A2 => n20535, ZN => n677);
   U2839 : OAI21_X1 port map( B1 => n5404, B2 => n5571, A => n5408, ZN => n5147
                           );
   U2840 : NAND3_X1 port map( A1 => n4607, A2 => n1908, A3 => n4312, ZN => n680
                           );
   U2842 : NAND2_X1 port map( A1 => n14658, A2 => n19748, ZN => n681);
   U2843 : XNOR2_X1 port map( A => n13185, B => n13248, ZN => n13186);
   U2844 : NAND2_X1 port map( A1 => n11725, A2 => n685, ZN => n683);
   U2845 : NAND2_X1 port map( A1 => n686, A2 => n924, ZN => n2143);
   U2846 : NAND2_X1 port map( A1 => n12537, A2 => n686, ZN => n11488);
   U2847 : INV_X1 port map( A => n12534, ZN => n686);
   U2849 : INV_X1 port map( A => n17315, ZN => n689);
   U2850 : NOR2_X1 port map( A1 => n690, A2 => n15573, ZN => n692);
   U2851 : INV_X1 port map( A => n15577, ZN => n691);
   U2852 : NAND2_X1 port map( A1 => n15791, A2 => n15796, ZN => n693);
   U2854 : XNOR2_X1 port map( A => n694, B => n17851, ZN => n10418);
   U2855 : XNOR2_X1 port map( A => n694, B => n9462, ZN => n9656);
   U2856 : XNOR2_X1 port map( A => n9799, B => n694, ZN => n8427);
   U2857 : XNOR2_X1 port map( A => n694, B => n9754, ZN => n9465);
   U2859 : NAND2_X1 port map( A1 => n699, A2 => n12126, ZN => n12134);
   U2860 : NAND2_X1 port map( A1 => n696, A2 => n699, ZN => n695);
   U2863 : NAND2_X1 port map( A1 => n2983, A2 => n238, ZN => n3172);
   U2864 : NAND2_X1 port map( A1 => n20262, A2 => n2983, ZN => n700);
   U2866 : NAND3_X1 port map( A1 => n9278, A2 => n9275, A3 => n8991, ZN => n702
                           );
   U2867 : INV_X1 port map( A => n11650, ZN => n11674);
   U2868 : OAI21_X1 port map( B1 => n3645, B2 => n8736, A => n19518, ZN => n708
                           );
   U2869 : INV_X1 port map( A => n8921, ZN => n705);
   U2870 : NAND2_X1 port map( A1 => n8497, A2 => n707, ZN => n706);
   U2871 : NOR2_X1 port map( A1 => n19518, A2 => n8923, ZN => n707);
   U2872 : NAND2_X1 port map( A1 => n8324, A2 => n276, ZN => n709);
   U2873 : NAND2_X1 port map( A1 => n711, A2 => n710, ZN => n9103);
   U2874 : NAND2_X1 port map( A1 => n8323, A2 => n1425, ZN => n710);
   U2875 : NAND2_X1 port map( A1 => n3611, A2 => n19856, ZN => n711);
   U2876 : NAND2_X1 port map( A1 => n3161, A2 => n3160, ZN => n712);
   U2878 : OAI22_X1 port map( A1 => n12383, A2 => n12138, B1 => n11917, B2 => 
                           n712, ZN => n11918);
   U2881 : NAND2_X1 port map( A1 => n2146, A2 => n15266, ZN => n716);
   U2882 : NAND3_X1 port map( A1 => n717, A2 => n15636, A3 => n716, ZN => n715)
                           ;
   U2883 : NAND3_X1 port map( A1 => n8214, A2 => n8213, A3 => n718, ZN => n9113
                           );
   U2884 : INV_X1 port map( A => n17886, ZN => n719);
   U2885 : NAND2_X1 port map( A1 => n719, A2 => n17887, ZN => n3214);
   U2886 : NAND2_X1 port map( A1 => n720, A2 => n12004, ZN => n1861);
   U2887 : NAND2_X1 port map( A1 => n12498, A2 => n12500, ZN => n720);
   U2890 : NAND2_X1 port map( A1 => n10007, A2 => n11575, ZN => n722);
   U2892 : NAND2_X1 port map( A1 => n10740, A2 => n11572, ZN => n727);
   U2894 : NAND2_X1 port map( A1 => n729, A2 => n3642, ZN => n728);
   U2895 : NAND2_X1 port map( A1 => n730, A2 => n14675, ZN => n729);
   U2896 : NAND2_X1 port map( A1 => n19530, A2 => n14542, ZN => n730);
   U2897 : XNOR2_X2 port map( A => n8757, B => n8756, ZN => n11538);
   U2898 : NAND2_X1 port map( A1 => n733, A2 => n5148, ZN => n3960);
   U2899 : AOI21_X1 port map( B1 => n5404, B2 => n733, A => n5582, ZN => n5409)
                           ;
   U2900 : MUX2_X1 port map( A => n5404, B => n733, S => n5148, Z => n3961);
   U2902 : XNOR2_X1 port map( A => n10494, B => n9477, ZN => n735);
   U2903 : XNOR2_X1 port map( A => n734, B => n10126, ZN => n10494);
   U2904 : INV_X1 port map( A => n9824, ZN => n734);
   U2906 : MUX2_X1 port map( A => n9576, B => n9291, S => n9049, Z => n736);
   U2907 : NAND2_X1 port map( A1 => n1541, A2 => n1538, ZN => n737);
   U2910 : NAND2_X1 port map( A1 => n11730, A2 => n11683, ZN => n740);
   U2911 : NAND2_X1 port map( A1 => n742, A2 => n11926, ZN => n741);
   U2912 : NAND2_X1 port map( A1 => n11923, A2 => n11922, ZN => n742);
   U2913 : OAI211_X1 port map( C1 => n9576, C2 => n9287, A => n743, B => n9291,
                           ZN => n744);
   U2914 : NAND2_X1 port map( A1 => n9576, A2 => n19715, ZN => n743);
   U2916 : NAND2_X1 port map( A1 => n9579, A2 => n746, ZN => n745);
   U2917 : OR2_X1 port map( A1 => n19519, A2 => n9576, ZN => n746);
   U2918 : NAND2_X1 port map( A1 => n747, A2 => n15607, ZN => n14975);
   U2919 : MUX2_X1 port map( A => n15608, B => n16126, S => n16129, Z => n14977
                           );
   U2920 : NAND2_X1 port map( A1 => n20007, A2 => n747, ZN => n15737);
   U2921 : NAND2_X1 port map( A1 => n15494, A2 => n747, ZN => n3432);
   U2922 : NAND2_X1 port map( A1 => n3415, A2 => n747, ZN => n3414);
   U2924 : NAND2_X1 port map( A1 => n749, A2 => n4610, ZN => n4616);
   U2925 : NAND2_X1 port map( A1 => n4365, A2 => n4013, ZN => n4610);
   U2926 : NAND2_X1 port map( A1 => n290, A2 => n4613, ZN => n749);
   U2927 : NAND2_X1 port map( A1 => n750, A2 => n20449, ZN => n1998);
   U2928 : NAND2_X1 port map( A1 => n14119, A2 => n19503, ZN => n751);
   U2929 : NAND2_X1 port map( A1 => n14006, A2 => n14232, ZN => n752);
   U2930 : NAND2_X1 port map( A1 => n754, A2 => n753, ZN => n11809);
   U2931 : NAND2_X1 port map( A1 => n1282, A2 => n9832, ZN => n754);
   U2933 : NAND2_X1 port map( A1 => n758, A2 => n757, ZN => n16441);
   U2934 : NAND2_X1 port map( A1 => n16434, A2 => n160, ZN => n757);
   U2935 : NAND2_X1 port map( A1 => n759, A2 => n226, ZN => n758);
   U2936 : NAND2_X1 port map( A1 => n4649, A2 => n4648, ZN => n760);
   U2937 : MUX2_X1 port map( A => n4644, B => n4643, S => n4642, Z => n761);
   U2938 : NAND2_X1 port map( A1 => n12107, A2 => n764, ZN => n974);
   U2939 : INV_X1 port map( A => n1840, ZN => n767);
   U2940 : INV_X1 port map( A => n2317, ZN => n768);
   U2942 : NAND2_X1 port map( A1 => n18953, A2 => n17831, ZN => n17830);
   U2943 : OR2_X1 port map( A1 => n7560, A2 => n8249, ZN => n769);
   U2944 : NAND2_X1 port map( A1 => n3540, A2 => n3541, ZN => n8435);
   U2945 : AND3_X2 port map( A1 => n3540, A2 => n3541, A3 => n770, ZN => n9780)
                           ;
   U2946 : NAND2_X1 port map( A1 => n3542, A2 => n9780, ZN => n772);
   U2947 : NAND2_X1 port map( A1 => n2983, A2 => n2773, ZN => n773);
   U2948 : NAND2_X1 port map( A1 => n15059, A2 => n15309, ZN => n15060);
   U2950 : NOR2_X1 port map( A1 => n14431, A2 => n14481, ZN => n774);
   U2951 : AOI21_X1 port map( B1 => n3900, B2 => n3899, A => n19822, ZN => n775
                           );
   U2952 : MUX2_X1 port map( A => n5791, B => n5300, S => n5428, Z => n5158);
   U2953 : NAND2_X1 port map( A1 => n776, A2 => n7922, ZN => n7923);
   U2956 : AOI21_X1 port map( B1 => n8705, B2 => n9168, A => n9167, ZN => n778)
                           ;
   U2957 : NAND2_X1 port map( A1 => n237, A2 => n779, ZN => n3244);
   U2958 : NAND2_X1 port map( A1 => n18332, A2 => n213, ZN => n18334);
   U2959 : INV_X1 port map( A => n781, ZN => n784);
   U2960 : AOI21_X1 port map( B1 => n13182, B2 => n13181, A => n2023, ZN => 
                           n781);
   U2962 : NAND2_X1 port map( A1 => n784, A2 => n782, ZN => n13183);
   U2963 : NAND2_X1 port map( A1 => n13182, A2 => n783, ZN => n782);
   U2964 : XNOR2_X1 port map( A => n785, B => n18587, ZN => n16573);
   U2965 : XNOR2_X1 port map( A => n785, B => n2376, ZN => n16046);
   U2966 : XNOR2_X1 port map( A => n785, B => n3162, ZN => n16386);
   U2967 : XNOR2_X1 port map( A => n16095, B => n785, ZN => n16828);
   U2968 : OR2_X1 port map( A1 => n7855, A2 => n282, ZN => n8259);
   U2969 : NAND2_X1 port map( A1 => n786, A2 => n8157, ZN => n7725);
   U2970 : NAND2_X1 port map( A1 => n7855, A2 => n282, ZN => n786);
   U2971 : NAND3_X1 port map( A1 => n279, A2 => n7724, A3 => n8157, ZN => n7554
                           );
   U2975 : NAND2_X1 port map( A1 => n15535, A2 => n15898, ZN => n789);
   U2976 : NAND2_X1 port map( A1 => n19838, A2 => n15401, ZN => n15535);
   U2977 : XNOR2_X1 port map( A => n10030, B => n791, ZN => n10383);
   U2978 : INV_X1 port map( A => Key(63), ZN => n791);
   U2979 : NAND3_X1 port map( A1 => n14023, A2 => n20266, A3 => n19748, ZN => 
                           n1977);
   U2982 : NAND2_X1 port map( A1 => n792, A2 => n20405, ZN => n2796);
   U2983 : XNOR2_X1 port map( A => n794, B => n793, ZN => Ciphertext(124));
   U2984 : INV_X1 port map( A => n1386, ZN => n793);
   U2985 : NAND2_X1 port map( A1 => n797, A2 => n795, ZN => n794);
   U2986 : AOI22_X1 port map( A1 => n796, A2 => n19069, B1 => n19653, B2 => 
                           n19070, ZN => n795);
   U2987 : INV_X1 port map( A => n19071, ZN => n796);
   U2988 : NAND2_X1 port map( A1 => n19072, A2 => n19071, ZN => n797);
   U2989 : NAND2_X1 port map( A1 => n19074, A2 => n19059, ZN => n19071);
   U2990 : NAND3_X2 port map( A1 => n11199, A2 => n799, A3 => n798, ZN => 
                           n12478);
   U2991 : NAND3_X1 port map( A1 => n19913, A2 => n19719, A3 => n11198, ZN => 
                           n799);
   U2992 : XNOR2_X2 port map( A => n10622, B => n3049, ZN => n11493);
   U2993 : INV_X1 port map( A => n7559, ZN => n800);
   U2994 : XNOR2_X1 port map( A => n5249, B => n302, ZN => n7027);
   U2996 : NAND2_X1 port map( A1 => n803, A2 => n9135, ZN => n2726);
   U2997 : NAND2_X1 port map( A1 => n9137, A2 => n803, ZN => n9215);
   U2998 : AOI22_X1 port map( A1 => n9135, A2 => n8446, B1 => n9134, B2 => n803
                           , ZN => n8447);
   U2999 : NOR2_X1 port map( A1 => n953, A2 => n12488, ZN => n11910);
   U3000 : NAND2_X1 port map( A1 => n5908, A2 => n890, ZN => n5495);
   U3001 : NAND2_X1 port map( A1 => n805, A2 => n5494, ZN => n804);
   U3003 : NAND2_X1 port map( A1 => n19462, A2 => n19463, ZN => n809);
   U3004 : XNOR2_X1 port map( A => n807, B => n16688, ZN => Ciphertext(189));
   U3005 : NAND3_X1 port map( A1 => n810, A2 => n808, A3 => n16682, ZN => n807)
                           ;
   U3006 : OAI211_X1 port map( C1 => n19463, C2 => n17091, A => n809, B => 
                           n20140, ZN => n808);
   U3007 : NAND2_X1 port map( A1 => n301, A2 => n4539, ZN => n4544);
   U3008 : NAND2_X1 port map( A1 => n4349, A2 => n301, ZN => n3760);
   U3009 : MUX2_X1 port map( A => n4347, B => n4348, S => n4541, Z => n4352);
   U3013 : NAND3_X1 port map( A1 => n17483, A2 => n17243, A3 => n812, ZN => 
                           n811);
   U3014 : NAND3_X1 port map( A1 => n815, A2 => n17479, A3 => n17480, ZN => 
                           n814);
   U3015 : NAND2_X1 port map( A1 => n817, A2 => n1718, ZN => n816);
   U3016 : OAI21_X1 port map( B1 => n17243, B2 => n17479, A => n818, ZN => n817
                           );
   U3017 : NAND2_X1 port map( A1 => n17479, A2 => n20353, ZN => n818);
   U3019 : NAND2_X1 port map( A1 => n2470, A2 => n10756, ZN => n11531);
   U3020 : NAND2_X1 port map( A1 => n819, A2 => n8200, ZN => n820);
   U3021 : INV_X1 port map( A => n8070, ZN => n819);
   U3022 : XNOR2_X2 port map( A => n5639, B => n5638, ZN => n8070);
   U3023 : NAND2_X1 port map( A1 => n289, A2 => n20459, ZN => n821);
   U3024 : NAND2_X1 port map( A1 => n1312, A2 => n1311, ZN => n822);
   U3025 : MUX2_X1 port map( A => n263, B => n9135, S => n9209, Z => n1334);
   U3026 : NAND2_X1 port map( A1 => n8351, A2 => n8350, ZN => n824);
   U3027 : XNOR2_X1 port map( A => n825, B => n6593, ZN => n5854);
   U3028 : INV_X1 port map( A => n3590, ZN => n825);
   U3029 : XNOR2_X1 port map( A => n3590, B => n826, ZN => n6638);
   U3030 : NAND2_X1 port map( A1 => n5073, A2 => n4664, ZN => n829);
   U3031 : NAND3_X1 port map( A1 => n4814, A2 => n5072, A3 => n4409, ZN => n830
                           );
   U3032 : NAND2_X1 port map( A1 => n4410, A2 => n5073, ZN => n4409);
   U3033 : XNOR2_X1 port map( A => n831, B => n18339, ZN => Ciphertext(133));
   U3034 : NAND2_X1 port map( A1 => n834, A2 => n832, ZN => n831);
   U3035 : NAND2_X1 port map( A1 => n835, A2 => n833, ZN => n832);
   U3036 : OAI22_X1 port map( A1 => n835, A2 => n19130, B1 => n20508, B2 => 
                           n19148, ZN => n834);
   U3037 : NAND2_X1 port map( A1 => n20508, A2 => n19135, ZN => n19130);
   U3038 : AND2_X1 port map( A1 => n18337, A2 => n19134, ZN => n835);
   U3039 : NAND2_X1 port map( A1 => n8322, A2 => n2548, ZN => n836);
   U3040 : AOI21_X1 port map( B1 => n7585, B2 => n8325, A => n8001, ZN => n837)
                           ;
   U3041 : NAND2_X1 port map( A1 => n8532, A2 => n8577, ZN => n839);
   U3042 : NAND3_X1 port map( A1 => n846, A2 => n843, A3 => n841, ZN => 
                           Ciphertext(61));
   U3043 : NAND2_X1 port map( A1 => n18647, A2 => n842, ZN => n841);
   U3044 : NAND2_X1 port map( A1 => n845, A2 => n844, ZN => n843);
   U3045 : AOI21_X1 port map( B1 => n18647, B2 => n18646, A => n299, ZN => n844
                           );
   U3046 : NAND2_X1 port map( A1 => n848, A2 => n18659, ZN => n845);
   U3047 : NAND2_X1 port map( A1 => n848, A2 => n847, ZN => n846);
   U3048 : AND2_X1 port map( A1 => n18659, A2 => n299, ZN => n847);
   U3049 : INV_X1 port map( A => n18645, ZN => n848);
   U3050 : OAI21_X1 port map( B1 => n850, B2 => n11794, A => n11792, ZN => n852
                           );
   U3053 : NAND3_X1 port map( A1 => n1511, A2 => n907, A3 => n12523, ZN => n851
                           );
   U3054 : INV_X1 port map( A => n12165, ZN => n1511);
   U3055 : INV_X1 port map( A => n16025, ZN => n854);
   U3056 : NAND2_X1 port map( A1 => n2732, A2 => n1339, ZN => n855);
   U3057 : OAI211_X1 port map( C1 => n8984, C2 => n8983, A => n8982, B => n3797
                           , ZN => n856);
   U3058 : OR2_X1 port map( A1 => n11128, A2 => n2029, ZN => n857);
   U3059 : OAI211_X1 port map( C1 => n1597, C2 => n2462, A => n1595, B => n1594
                           , ZN => n861);
   U3060 : OAI211_X1 port map( C1 => n1597, C2 => n2462, A => n1595, B => n1594
                           , ZN => n862);
   U3062 : OAI211_X1 port map( C1 => n1597, C2 => n2462, A => n1595, B => n1594
                           , ZN => n5920);
   U3065 : NAND2_X1 port map( A1 => n2300, A2 => n2299, ZN => n865);
   U3068 : OAI21_X1 port map( B1 => n14066, B2 => n14065, A => n14064, ZN => 
                           n15843);
   U3069 : XNOR2_X1 port map( A => n5690, B => n6534, ZN => n5727);
   U3070 : AOI21_X1 port map( B1 => n16726, B2 => n20127, A => n16725, ZN => 
                           n19143);
   U3072 : XNOR2_X1 port map( A => Key(126), B => Plaintext(126), ZN => n873);
   U3073 : INV_X1 port map( A => n12041, ZN => n876);
   U3074 : OAI211_X1 port map( C1 => n9260, C2 => n19516, A => n9258, B => 
                           n9257, ZN => n878);
   U3075 : OAI211_X1 port map( C1 => n15850, C2 => n15851, A => n15849, B => 
                           n15848, ZN => n879);
   U3076 : OAI211_X1 port map( C1 => n15850, C2 => n15851, A => n15849, B => 
                           n15848, ZN => n880);
   U3077 : XNOR2_X1 port map( A => n11593, B => n11592, ZN => n14779);
   U3078 : OAI211_X1 port map( C1 => n9260, C2 => n19516, A => n9258, B => 
                           n9257, ZN => n9878);
   U3080 : OR2_X1 port map( A1 => n18382, A2 => n18384, ZN => n881);
   U3081 : NAND2_X1 port map( A1 => n881, A2 => n18394, ZN => n2274);
   U3082 : OAI21_X1 port map( B1 => n11016, B2 => n1579, A => n10956, ZN => 
                           n882);
   U3083 : OAI211_X1 port map( C1 => n5242, C2 => n5714, A => n4376, B => n2207
                           , ZN => n883);
   U3084 : OAI21_X1 port map( B1 => n11016, B2 => n1579, A => n10956, ZN => 
                           n12127);
   U3085 : OAI211_X1 port map( C1 => n5242, C2 => n5714, A => n4376, B => n2207
                           , ZN => n7325);
   U3086 : OAI211_X2 port map( C1 => n14576, C2 => n14570, A => n14272, B => 
                           n14271, ZN => n15400);
   U3087 : INV_X1 port map( A => n7457, ZN => n8053);
   U3088 : OR2_X1 port map( A1 => n8361, A2 => n7709, ZN => n884);
   U3089 : NAND2_X1 port map( A1 => n884, A2 => n1994, ZN => n7512);
   U3090 : NAND2_X1 port map( A1 => n7875, A2 => n7874, ZN => n885);
   U3092 : XNOR2_X1 port map( A => n10609, B => n10610, ZN => n888);
   U3093 : XOR2_X1 port map( A => n17031, B => n17030, Z => n889);
   U3095 : XOR2_X1 port map( A => n6856, B => n6857, Z => n6862);
   U3096 : NAND2_X1 port map( A1 => n4838, A2 => n4837, ZN => n890);
   U3097 : INV_X1 port map( A => n9018, ZN => n891);
   U3098 : INV_X1 port map( A => n17729, ZN => n893);
   U3099 : AND2_X1 port map( A1 => n19755, A2 => n10873, ZN => n894);
   U3100 : XNOR2_X1 port map( A => Key(63), B => Plaintext(63), ZN => n896);
   U3103 : XNOR2_X1 port map( A => Key(63), B => Plaintext(63), ZN => n4866);
   U3105 : NAND2_X1 port map( A1 => n14877, A2 => n14878, ZN => n897);
   U3106 : XNOR2_X1 port map( A => n9964, B => n9963, ZN => n898);
   U3107 : NAND2_X1 port map( A1 => n14877, A2 => n14878, ZN => n16336);
   U3108 : XNOR2_X1 port map( A => n9964, B => n9963, ZN => n11182);
   U3110 : BUF_X1 port map( A => n15957, Z => n902);
   U3111 : OAI22_X1 port map( A1 => n15707, A2 => n15706, B1 => n2625, B2 => 
                           n16009, ZN => n15957);
   U3112 : NAND2_X1 port map( A1 => n5976, A2 => n5977, ZN => n903);
   U3113 : INV_X1 port map( A => n905, ZN => n904);
   U3114 : NAND2_X1 port map( A1 => n5976, A2 => n5977, ZN => n7372);
   U3115 : NAND2_X1 port map( A1 => n3850, A2 => n3849, ZN => n906);
   U3116 : INV_X1 port map( A => n11493, ZN => n3521);
   U3118 : OAI21_X1 port map( B1 => n11463, B2 => n11886, A => n11462, ZN => 
                           n907);
   U3119 : INV_X1 port map( A => n8795, ZN => n908);
   U3120 : XNOR2_X1 port map( A => n16347, B => n17411, ZN => n16921);
   U3121 : INV_X1 port map( A => n9748, ZN => n9977);
   U3123 : NOR2_X1 port map( A1 => n15819, A2 => n2114, ZN => n911);
   U3124 : XNOR2_X1 port map( A => n10602, B => n10601, ZN => n913);
   U3126 : XNOR2_X1 port map( A => n12830, B => n12829, ZN => n14820);
   U3129 : XNOR2_X1 port map( A => n12071, B => n12070, ZN => n13206);
   U3130 : XNOR2_X1 port map( A => n13720, B => n13719, ZN => n14228);
   U3131 : AND2_X1 port map( A1 => n20263, A2 => n14482, ZN => n914);
   U3132 : OR2_X1 port map( A1 => n12359, A2 => n12509, ZN => n916);
   U3133 : NOR2_X1 port map( A1 => n12366, A2 => n12365, ZN => n13781);
   U3134 : NAND3_X1 port map( A1 => n8170, A2 => n8169, A3 => n8168, ZN => n917
                           );
   U3135 : NAND3_X1 port map( A1 => n8170, A2 => n8169, A3 => n8168, ZN => n918
                           );
   U3136 : XOR2_X1 port map( A => n13286, B => n13285, Z => n919);
   U3138 : INV_X1 port map( A => n14159, ZN => n921);
   U3139 : XNOR2_X1 port map( A => n6638, B => n6637, ZN => n923);
   U3140 : XNOR2_X1 port map( A => n6638, B => n6637, ZN => n8066);
   U3141 : OR2_X1 port map( A1 => n17937, A2 => n18349, ZN => n925);
   U3142 : NAND2_X1 port map( A1 => n925, A2 => n17908, ZN => n17910);
   U3143 : XNOR2_X1 port map( A => n9440, B => n9439, ZN => n926);
   U3144 : XNOR2_X1 port map( A => n9956, B => n926, ZN => n927);
   U3145 : OAI211_X1 port map( C1 => n9142, C2 => n9213, A => n9141, B => n9140
                           , ZN => n928);
   U3147 : XNOR2_X1 port map( A => n9956, B => n926, ZN => n11566);
   U3148 : OAI211_X1 port map( C1 => n9142, C2 => n9213, A => n9141, B => n9140
                           , ZN => n10358);
   U3149 : AOI21_X1 port map( B1 => n19387, B2 => n15731, A => n15730, ZN => 
                           n18412);
   U3150 : XNOR2_X1 port map( A => n10621, B => n10321, ZN => n9951);
   U3151 : XNOR2_X2 port map( A => n6807, B => n6806, ZN => n7855);
   U3152 : XNOR2_X1 port map( A => n10247, B => n10008, ZN => n929);
   U3153 : NAND2_X1 port map( A1 => n17863, A2 => n16681, ZN => n930);
   U3154 : NAND2_X1 port map( A1 => n16680, A2 => n16679, ZN => n931);
   U3155 : XNOR2_X1 port map( A => n13453, B => n13369, ZN => n933);
   U3156 : XNOR2_X1 port map( A => n7378, B => n7379, ZN => n934);
   U3158 : INV_X1 port map( A => n17729, ZN => n18485);
   U3159 : OAI211_X2 port map( C1 => n2781, C2 => n8614, A => n8613, B => n8612
                           , ZN => n9879);
   U3160 : XNOR2_X1 port map( A => n16700, B => n16699, ZN => n935);
   U3161 : XNOR2_X1 port map( A => n16084, B => n16335, ZN => n936);
   U3162 : OR2_X1 port map( A1 => n17698, A2 => n17697, ZN => n938);
   U3163 : OR2_X1 port map( A1 => n14818, A2 => n14091, ZN => n939);
   U3165 : OAI21_X1 port map( B1 => n11618, B2 => n11897, A => n11896, ZN => 
                           n940);
   U3167 : OAI211_X1 port map( C1 => n5874, C2 => n5873, A => n5872, B => n5871
                           , ZN => n943);
   U3171 : OAI211_X1 port map( C1 => n5874, C2 => n5873, A => n5872, B => n5871
                           , ZN => n6249);
   U3172 : OAI21_X2 port map( B1 => n4416, B2 => n4415, A => n4414, ZN => n6123
                           );
   U3174 : AND2_X1 port map( A1 => n5573, A2 => n5574, ZN => n946);
   U3176 : OAI211_X2 port map( C1 => n14137, C2 => n14408, A => n14136, B => 
                           n14135, ZN => n16129);
   U3179 : INV_X1 port map( A => Plaintext(142), ZN => n2990);
   U3181 : XNOR2_X1 port map( A => n5727, B => n5726, ZN => n8200);
   U3182 : XNOR2_X1 port map( A => n6512, B => n6811, ZN => n7334);
   U3183 : XNOR2_X1 port map( A => n5759, B => n1863, ZN => n2886);
   U3184 : XNOR2_X1 port map( A => n6509, B => n3321, ZN => n8247);
   U3185 : OR2_X1 port map( A1 => n6904, A2 => n7753, ZN => n3271);
   U3187 : INV_X1 port map( A => n2886, ZN => n7421);
   U3188 : AND2_X1 port map( A1 => n8178, A2 => n8179, ZN => n7416);
   U3189 : INV_X1 port map( A => n8247, ZN => n8245);
   U3190 : INV_X1 port map( A => n8113, ZN => n7844);
   U3191 : OR2_X1 port map( A1 => n7722, A2 => n8352, ZN => n2155);
   U3192 : AND2_X1 port map( A1 => n7833, A2 => n8910, ZN => n7918);
   U3193 : OR2_X1 port map( A1 => n7507, A2 => n7748, ZN => n1548);
   U3195 : XNOR2_X1 port map( A => n10461, B => n10061, ZN => n10356);
   U3196 : XNOR2_X1 port map( A => n1031, B => n1029, ZN => n9432);
   U3197 : XNOR2_X1 port map( A => n10621, B => n3050, ZN => n3049);
   U3198 : XNOR2_X1 port map( A => n10620, B => n1605, ZN => n3050);
   U3199 : INV_X1 port map( A => n10960, ZN => n11143);
   U3200 : OR2_X1 port map( A1 => n11124, A2 => n85, ZN => n2033);
   U3201 : OR2_X1 port map( A1 => n11540, A2 => n11168, ZN => n3279);
   U3202 : AND2_X1 port map( A1 => n12289, A2 => n12288, ZN => n1440);
   U3203 : INV_X1 port map( A => n13697, ZN => n12769);
   U3204 : INV_X1 port map( A => n11640, ZN => n13792);
   U3205 : OAI211_X1 port map( C1 => n11647, C2 => n11646, A => n12227, B => 
                           n11692, ZN => n11648);
   U3206 : XNOR2_X1 port map( A => n13503, B => n13502, ZN => n14490);
   U3207 : XNOR2_X1 port map( A => n13139, B => n3498, ZN => n13471);
   U3208 : XNOR2_X1 port map( A => n12872, B => n12871, ZN => n13927);
   U3209 : AND2_X1 port map( A1 => n13927, A2 => n14451, ZN => n13559);
   U3210 : INV_X1 port map( A => n14493, ZN => n1936);
   U3211 : NOR2_X1 port map( A1 => n15424, A2 => n14238, ZN => n14243);
   U3212 : XNOR2_X1 port map( A => n3543, B => Key(53), ZN => n4233);
   U3213 : INV_X1 port map( A => n4950, ZN => n3265);
   U3214 : XNOR2_X1 port map( A => Plaintext(45), B => Key(45), ZN => n4969);
   U3215 : AND2_X1 port map( A1 => n5055, A2 => n4100, ZN => n5053);
   U3216 : INV_X1 port map( A => n4887, ZN => n4947);
   U3217 : INV_X1 port map( A => Plaintext(64), ZN => n1088);
   U3218 : INV_X1 port map( A => n6410, ZN => n7025);
   U3219 : OR2_X1 port map( A1 => n5763, A2 => n5736, ZN => n2239);
   U3220 : OR2_X1 port map( A1 => n5805, A2 => n6192, ZN => n4593);
   U3221 : XNOR2_X1 port map( A => n7054, B => n7053, ZN => n2977);
   U3222 : NOR2_X1 port map( A1 => n4062, A2 => n956, ZN => n1131);
   U3223 : INV_X1 port map( A => n6510, ZN => n8248);
   U3224 : OR2_X1 port map( A1 => n7982, A2 => n7981, ZN => n7767);
   U3225 : INV_X1 port map( A => n1507, ZN => n1574);
   U3226 : AND2_X1 port map( A1 => n7312, A2 => n7311, ZN => n8323);
   U3227 : AND2_X1 port map( A1 => n3395, A2 => n3394, ZN => n1841);
   U3228 : INV_X1 port map( A => n7311, ZN => n7590);
   U3229 : AND2_X1 port map( A1 => n7958, A2 => n2977, ZN => n2976);
   U3230 : AOI21_X1 port map( B1 => n8013, B2 => n8012, A => n7826, ZN => n3625
                           );
   U3231 : OR2_X1 port map( A1 => n8035, A2 => n8286, ZN => n2165);
   U3233 : NOR2_X1 port map( A1 => n7909, A2 => n274, ZN => n1785);
   U3234 : XNOR2_X1 port map( A => n6717, B => n6720, ZN => n2824);
   U3235 : INV_X1 port map( A => n7675, ZN => n1994);
   U3236 : OR2_X1 port map( A1 => n7622, A2 => n8177, ZN => n3523);
   U3237 : OR2_X1 port map( A1 => n7003, A2 => n7755, ZN => n7004);
   U3238 : NOR2_X1 port map( A1 => n8002, A2 => n3076, ZN => n3075);
   U3242 : XNOR2_X1 port map( A => n10151, B => n10491, ZN => n10549);
   U3243 : INV_X1 port map( A => n10980, ZN => n11291);
   U3244 : AND2_X1 port map( A1 => n10980, A2 => n11294, ZN => n11406);
   U3245 : XNOR2_X1 port map( A => n1284, B => n1283, ZN => n1285);
   U3246 : INV_X1 port map( A => n10808, ZN => n11883);
   U3247 : INV_X1 port map( A => n1040, ZN => n1317);
   U3248 : OR2_X1 port map( A1 => n3789, A2 => n11177, ZN => n10966);
   U3249 : XNOR2_X1 port map( A => n2202, B => n7664, ZN => n10945);
   U3250 : XNOR2_X1 port map( A => n10510, B => n1479, ZN => n11302);
   U3251 : XNOR2_X1 port map( A => n9771, B => n18379, ZN => n9772);
   U3252 : INV_X1 port map( A => n12463, ZN => n11915);
   U3254 : OR2_X1 port map( A1 => n11217, A2 => n11475, ZN => n3768);
   U3255 : OR2_X1 port map( A1 => n11289, A2 => n10950, ZN => n3023);
   U3257 : INV_X1 port map( A => n12252, ZN => n3637);
   U3258 : OR2_X1 port map( A1 => n11078, A2 => n11474, ZN => n2464);
   U3260 : OR2_X1 port map( A1 => n11006, A2 => n19851, ZN => n3175);
   U3261 : NAND2_X1 port map( A1 => n1663, A2 => n1664, ZN => n12255);
   U3262 : INV_X1 port map( A => n11243, ZN => n1599);
   U3263 : OAI21_X1 port map( B1 => n1748, B2 => n11140, A => n1747, ZN => 
                           n11146);
   U3264 : INV_X1 port map( A => n12600, ZN => n12072);
   U3265 : INV_X1 port map( A => n14623, ZN => n14001);
   U3266 : XNOR2_X1 port map( A => n13204, B => n977, ZN => n12654);
   U3268 : XNOR2_X1 port map( A => n13481, B => n13081, ZN => n13199);
   U3269 : INV_X1 port map( A => n12479, ZN => n2553);
   U3270 : XNOR2_X1 port map( A => n13204, B => n13205, ZN => n13209);
   U3271 : OR2_X1 port map( A1 => n1208, A2 => n14020, ZN => n1207);
   U3272 : XNOR2_X1 port map( A => n13807, B => n13251, ZN => n2832);
   U3273 : XNOR2_X1 port map( A => n3742, B => n3743, ZN => n14120);
   U3274 : XNOR2_X1 port map( A => n13773, B => n13770, ZN => n2623);
   U3275 : INV_X1 port map( A => n15313, ZN => n14146);
   U3276 : BUF_X1 port map( A => n14103, Z => n14788);
   U3278 : OR2_X1 port map( A1 => n14127, A2 => n19921, ZN => n13950);
   U3279 : INV_X1 port map( A => n14599, ZN => n1264);
   U3280 : XNOR2_X1 port map( A => n12972, B => n12971, ZN => n14032);
   U3281 : OR2_X1 port map( A1 => n14442, A2 => n14168, ZN => n2773);
   U3284 : NAND2_X1 port map( A1 => n15488, A2 => n15487, ZN => n15758);
   U3285 : OR2_X1 port map( A1 => n2808, A2 => n14196, ZN => n3006);
   U3286 : INV_X1 port map( A => n15421, ZN => n2974);
   U3287 : AND2_X1 port map( A1 => n19752, A2 => n15921, ZN => n1119);
   U3288 : OR2_X1 port map( A1 => n3174, A2 => n12919, ZN => n2088);
   U3289 : OR2_X1 port map( A1 => n13866, A2 => n15121, ZN => n1789);
   U3290 : OR2_X1 port map( A1 => n1795, A2 => n13559, ZN => n1794);
   U3291 : AND2_X1 port map( A1 => n14172, A2 => n14171, ZN => n13883);
   U3292 : OR2_X1 port map( A1 => n14750, A2 => n14747, ZN => n3267);
   U3293 : OR2_X1 port map( A1 => n14981, A2 => n15553, ZN => n3042);
   U3294 : OR2_X1 port map( A1 => n4824, A2 => n5258, ZN => n4825);
   U3295 : XNOR2_X1 port map( A => n3874, B => Key(23), ZN => n4021);
   U3297 : OR2_X1 port map( A1 => n177, A2 => n3995, ZN => n4682);
   U3298 : OR2_X1 port map( A1 => n4391, A2 => n4685, ZN => n4854);
   U3299 : OR2_X1 port map( A1 => n5079, A2 => n4719, ZN => n1163);
   U3300 : OR2_X1 port map( A1 => n5080, A2 => n5075, ZN => n5078);
   U3302 : INV_X1 port map( A => n4532, ZN => n3551);
   U3303 : INV_X1 port map( A => n5226, ZN => n6202);
   U3304 : INV_X1 port map( A => n4793, ZN => n3167);
   U3305 : OR2_X1 port map( A1 => n4056, A2 => n4060, ZN => n4741);
   U3306 : INV_X1 port map( A => n4796, ZN => n2670);
   U3307 : OR2_X1 port map( A1 => n4088, A2 => n5046, ZN => n5044);
   U3308 : INV_X1 port map( A => n4198, ZN => n1391);
   U3309 : OR2_X1 port map( A1 => n4504, A2 => n4565, ZN => n4753);
   U3310 : XNOR2_X1 port map( A => n3204, B => Key(124), ZN => n4706);
   U3311 : OR2_X1 port map( A1 => n4618, A2 => n4982, ZN => n1803);
   U3312 : OR2_X1 port map( A1 => n4114, A2 => n4940, ZN => n2389);
   U3313 : INV_X1 port map( A => n4271, ZN => n5025);
   U3314 : INV_X1 port map( A => n4440, ZN => n5040);
   U3316 : INV_X1 port map( A => n6168, ZN => n1867);
   U3317 : INV_X1 port map( A => n292, ZN => n3231);
   U3318 : OR2_X1 port map( A1 => n4613, A2 => n4614, ZN => n3716);
   U3319 : OR2_X1 port map( A1 => n4674, A2 => n4673, ZN => n3191);
   U3320 : OR2_X1 port map( A1 => n4969, A2 => n4968, ZN => n4971);
   U3321 : OR2_X1 port map( A1 => n5054, A2 => n5055, ZN => n2266);
   U3322 : OR2_X1 port map( A1 => n6003, A2 => n6002, ZN => n1454);
   U3323 : OR2_X1 port map( A1 => n6138, A2 => n3188, ZN => n4461);
   U3324 : AND2_X1 port map( A1 => n5996, A2 => n5998, ZN => n3604);
   U3325 : OR2_X1 port map( A1 => n4114, A2 => n4118, ZN => n3896);
   U3326 : MUX2_X1 port map( A => n4481, B => n4480, S => n4479, Z => n3043);
   U3327 : OR2_X2 port map( A1 => n4666, A2 => n4665, ZN => n6172);
   U3329 : OR2_X1 port map( A1 => n7445, A2 => n19686, ZN => n3662);
   U3331 : OR2_X1 port map( A1 => n5733, A2 => n6194, ZN => n2866);
   U3332 : INV_X1 port map( A => n7500, ZN => n8358);
   U3333 : INV_X1 port map( A => n7739, ZN => n8357);
   U3335 : AND2_X1 port map( A1 => n8112, A2 => n8241, ZN => n1271);
   U3336 : OR2_X1 port map( A1 => n9021, A2 => n8672, ZN => n8838);
   U3337 : OR2_X1 port map( A1 => n9023, A2 => n8510, ZN => n1631);
   U3338 : INV_X1 port map( A => n2499, ZN => n2501);
   U3339 : AND2_X1 port map( A1 => n8947, A2 => n8945, ZN => n8731);
   U3340 : INV_X1 port map( A => n7748, ZN => n7911);
   U3341 : INV_X1 port map( A => n7749, ZN => n7745);
   U3343 : OAI211_X1 port map( C1 => n8011, C2 => n7830, A => n8013, B => n273,
                           ZN => n7831);
   U3344 : INV_X1 port map( A => n9121, ZN => n9124);
   U3345 : NOR2_X1 port map( A1 => n8815, A2 => n8813, ZN => n9123);
   U3346 : AND2_X1 port map( A1 => n7745, A2 => n7507, ZN => n7694);
   U3347 : AND2_X1 port map( A1 => n7749, A2 => n3446, ZN => n7691);
   U3348 : OAI21_X1 port map( B1 => n3445, B2 => n1308, A => n3368, ZN => n8125
                           );
   U3349 : AOI21_X1 port map( B1 => n7769, B2 => n3376, A => n3375, ZN => n8772
                           );
   U3350 : INV_X1 port map( A => n3271, ZN => n7758);
   U3351 : INV_X1 port map( A => n9113, ZN => n1602);
   U3352 : AND2_X1 port map( A1 => n6617, A2 => n1962, ZN => n1961);
   U3353 : OR2_X1 port map( A1 => n8786, A2 => n2499, ZN => n2498);
   U3354 : OR2_X1 port map( A1 => n9236, A2 => n9235, ZN => n9237);
   U3355 : OAI21_X1 port map( B1 => n8439, B2 => n261, A => n8789, ZN => n1737)
                           ;
   U3356 : AOI21_X1 port map( B1 => n8332, B2 => n7533, A => n8499, ZN => n2747
                           );
   U3357 : AOI21_X1 port map( B1 => n19518, B2 => n8920, A => n8923, ZN => 
                           n2746);
   U3359 : INV_X1 port map( A => n9067, ZN => n2503);
   U3360 : AOI21_X1 port map( B1 => n9134, B2 => n9213, A => n1324, ZN => n1323
                           );
   U3361 : XNOR2_X1 port map( A => n10280, B => n10087, ZN => n10397);
   U3362 : OR2_X1 port map( A1 => n9069, A2 => n2749, ZN => n8075);
   U3363 : OAI211_X1 port map( C1 => n9840, C2 => n2749, A => n9839, B => n9838
                           , ZN => n9841);
   U3364 : XNOR2_X1 port map( A => n3628, B => n10091, ZN => n1040);
   U3365 : OR2_X1 port map( A1 => n7661, A2 => n8596, ZN => n2478);
   U3366 : OR2_X1 port map( A1 => n8924, A2 => n8749, ZN => n2479);
   U3367 : AND2_X1 port map( A1 => n9167, A2 => n9171, ZN => n7989);
   U3368 : NAND2_X1 port map( A1 => n2300, A2 => n2299, ZN => n10542);
   U3369 : OR2_X1 port map( A1 => n9064, A2 => n8829, ZN => n2299);
   U3370 : NAND2_X1 port map( A1 => n8922, A2 => n2301, ZN => n10039);
   U3371 : AND2_X1 port map( A1 => n8411, A2 => n9233, ZN => n2650);
   U3372 : OAI21_X1 port map( B1 => n9238, B2 => n8411, A => n2653, ZN => n2651
                           );
   U3373 : AND2_X1 port map( A1 => n11883, A2 => n3441, ZN => n11887);
   U3374 : OR2_X1 port map( A1 => n8941, A2 => n8945, ZN => n2400);
   U3375 : OR2_X1 port map( A1 => n3400, A2 => n12634, ZN => n1387);
   U3376 : OR2_X1 port map( A1 => n9147, A2 => n9145, ZN => n1542);
   U3377 : INV_X1 port map( A => n10046, ZN => n2689);
   U3378 : OR2_X1 port map( A1 => n8701, A2 => n9070, ZN => n8169);
   U3379 : INV_X1 port map( A => n9919, ZN => n11476);
   U3381 : INV_X1 port map( A => n11359, ZN => n3458);
   U3382 : OR2_X1 port map( A1 => n12129, A2 => n1508, ZN => n1546);
   U3383 : INV_X1 port map( A => n10683, ZN => n3601);
   U3384 : INV_X1 port map( A => n11500, ZN => n3234);
   U3385 : AND2_X1 port map( A1 => n19897, A2 => n20233, ZN => n2536);
   U3386 : INV_X1 port map( A => n3260, ZN => n12147);
   U3387 : OR2_X1 port map( A1 => n11293, A2 => n11294, ZN => n3585);
   U3388 : MUX2_X1 port map( A => n11520, B => n11519, S => n12533, Z => n13293
                           );
   U3389 : NAND3_X1 port map( A1 => n12632, A2 => n1689, A3 => n1240, ZN => 
                           n13596);
   U3390 : INV_X1 port map( A => n12002, ZN => n12355);
   U3391 : AOI21_X1 port map( B1 => n1396, B2 => n1397, A => n12338, ZN => 
                           n11669);
   U3393 : NOR2_X1 port map( A1 => n3781, A2 => n11699, ZN => n3780);
   U3396 : NOR2_X1 port map( A1 => n11642, A2 => n11586, ZN => n11590);
   U3397 : XNOR2_X1 port map( A => n13293, B => n13344, ZN => n13569);
   U3398 : OR2_X1 port map( A1 => n11018, A2 => n12576, ZN => n2345);
   U3399 : INV_X1 port map( A => n11730, ZN => n11017);
   U3400 : AOI22_X1 port map( A1 => n11938, A2 => n12443, B1 => n11937, B2 => 
                           n1522, ZN => n11941);
   U3401 : OR2_X1 port map( A1 => n11943, A2 => n11942, ZN => n1400);
   U3402 : XNOR2_X1 port map( A => n1260, B => n13330, ZN => n13332);
   U3403 : OAI21_X1 port map( B1 => n1578, B2 => n11953, A => n11659, ZN => 
                           n3024);
   U3404 : AND3_X1 port map( A1 => n1633, A2 => n12002, A3 => n11032, ZN => 
                           n1634);
   U3405 : OR2_X1 port map( A1 => n1636, A2 => n9380, ZN => n1635);
   U3406 : AOI22_X1 port map( A1 => n11775, A2 => n12281, B1 => n11776, B2 => 
                           n12282, ZN => n11780);
   U3407 : XNOR2_X1 port map( A => n13201, B => n13202, ZN => n14021);
   U3408 : AND2_X1 port map( A1 => n12684, A2 => n12429, ZN => n3647);
   U3409 : AND2_X1 port map( A1 => n12525, A2 => n12528, ZN => n12172);
   U3410 : OR2_X1 port map( A1 => n12231, A2 => n11646, ZN => n12233);
   U3411 : AND2_X1 port map( A1 => n11033, A2 => n11032, ZN => n3536);
   U3412 : XNOR2_X1 port map( A => n13319, B => n13596, ZN => n13842);
   U3414 : OR2_X1 port map( A1 => n3156, A2 => n19728, ZN => n3154);
   U3415 : OR2_X1 port map( A1 => n14032, A2 => n14642, ZN => n2972);
   U3416 : INV_X1 port map( A => n15120, ZN => n1802);
   U3417 : NOR2_X1 port map( A1 => n14487, A2 => n14172, ZN => n14481);
   U3418 : INV_X1 port map( A => n13872, ZN => n14651);
   U3419 : NOR2_X1 port map( A1 => n14516, A2 => n14321, ZN => n14519);
   U3421 : XNOR2_X1 port map( A => n13061, B => n13062, ZN => n15119);
   U3423 : XNOR2_X1 port map( A => n2947, B => n13549, ZN => n13553);
   U3424 : OR2_X1 port map( A1 => n13908, A2 => n14203, ZN => n13909);
   U3425 : INV_X1 port map( A => n13927, ZN => n14447);
   U3426 : NOR2_X1 port map( A1 => n192, A2 => n19740, ZN => n15335);
   U3427 : AND2_X1 port map( A1 => n15445, A2 => n15678, ZN => n2437);
   U3428 : OAI21_X1 port map( B1 => n15076, B2 => n15077, A => n15906, ZN => 
                           n1412);
   U3429 : OR2_X1 port map( A1 => n3019, A2 => n3778, ZN => n3576);
   U3430 : NOR2_X1 port map( A1 => n15081, A2 => n15430, ZN => n15433);
   U3431 : AND2_X1 port map( A1 => n14371, A2 => n2721, ZN => n2720);
   U3432 : AND3_X1 port map( A1 => n1181, A2 => n1925, A3 => n20094, ZN => 
                           n15877);
   U3433 : NAND3_X1 port map( A1 => n15189, A2 => n14935, A3 => n13933, ZN => 
                           n1757);
   U3435 : OR2_X1 port map( A1 => n3688, A2 => n15768, ZN => n3686);
   U3436 : OR2_X1 port map( A1 => n14938, A2 => n20449, ZN => n3136);
   U3437 : NOR2_X1 port map( A1 => n18948, A2 => n18946, ZN => n3546);
   U3438 : OR2_X1 port map( A1 => n15703, A2 => n15702, ZN => n1877);
   U3439 : AND2_X1 port map( A1 => n2364, A2 => n2363, ZN => n2862);
   U3440 : AOI21_X1 port map( B1 => n15439, B2 => n15775, A => n1639, ZN => 
                           n15440);
   U3441 : XNOR2_X1 port map( A => n16335, B => n16084, ZN => n16696);
   U3444 : INV_X1 port map( A => n17098, ZN => n15970);
   U3445 : XNOR2_X1 port map( A => n16597, B => n16598, ZN => n19389);
   U3446 : AND2_X1 port map( A1 => n19501, A2 => n18382, ZN => n2794);
   U3447 : INV_X1 port map( A => n17221, ZN => n3389);
   U3448 : INV_X1 port map( A => n16251, ZN => n17211);
   U3449 : NOR2_X1 port map( A1 => n17211, A2 => n19975, ZN => n17214);
   U3450 : AND2_X1 port map( A1 => n17210, A2 => n17208, ZN => n2841);
   U3451 : XNOR2_X1 port map( A => n3736, B => n16240, ZN => n3735);
   U3452 : XNOR2_X1 port map( A => n16921, B => n17291, ZN => n3574);
   U3453 : XNOR2_X1 port map( A => n16361, B => n16362, ZN => n18112);
   U3454 : NOR2_X1 port map( A1 => n17080, A2 => n17824, ZN => n3293);
   U3455 : XNOR2_X1 port map( A => n16033, B => n17371, ZN => n17181);
   U3456 : XNOR2_X1 port map( A => n16040, B => n16041, ZN => n16781);
   U3457 : NOR2_X1 port map( A1 => n4011, A2 => n1537, ZN => n1536);
   U3458 : INV_X1 port map( A => n20002, ZN => n3451);
   U3459 : OR2_X1 port map( A1 => n4960, A2 => n292, ZN => n4898);
   U3461 : INV_X1 port map( A => n5075, ZN => n4457);
   U3462 : OR2_X1 port map( A1 => n4539, A2 => n4350, ZN => n4348);
   U3463 : AND2_X1 port map( A1 => n3607, A2 => n3752, ZN => n3606);
   U3465 : INV_X1 port map( A => n5088, ZN => n5090);
   U3466 : OAI211_X1 port map( C1 => n5069, C2 => n2971, A => n5073, B => n291,
                           ZN => n5505);
   U3467 : OR2_X1 port map( A1 => n4438, A2 => n4804, ZN => n2115);
   U3468 : INV_X1 port map( A => n5866, ZN => n2158);
   U3470 : OR2_X1 port map( A1 => n5674, A2 => n5424, ZN => n4212);
   U3471 : AND2_X1 port map( A1 => n6113, A2 => n6107, ZN => n5658);
   U3472 : OR2_X1 port map( A1 => n5104, A2 => n5102, ZN => n1420);
   U3473 : AOI22_X1 port map( A1 => n4885, A2 => n4946, B1 => n4467, B2 => 
                           n4002, ZN => n5250);
   U3474 : OR2_X1 port map( A1 => n3760, A2 => n4540, ZN => n3759);
   U3475 : INV_X1 port map( A => n287, ZN => n3071);
   U3476 : INV_X1 port map( A => n5401, ZN => n4282);
   U3477 : INV_X1 port map( A => n6183, ZN => n3196);
   U3478 : OR2_X1 port map( A1 => n5114, A2 => n1915, ZN => n3650);
   U3479 : OR2_X1 port map( A1 => n5798, A2 => n1776, ZN => n5156);
   U3480 : OR2_X1 port map( A1 => n4722, A2 => n5076, ZN => n1569);
   U3481 : INV_X1 port map( A => n5927, ZN => n6026);
   U3482 : OR2_X1 port map( A1 => n5200, A2 => n5492, ZN => n6092);
   U3483 : OR2_X1 port map( A1 => n5697, A2 => n5699, ZN => n5528);
   U3484 : OAI21_X1 port map( B1 => n5929, B2 => n5030, A => n3371, ZN => n5521
                           );
   U3485 : OAI211_X1 port map( C1 => n6206, C2 => n287, A => n3044, B => n6204,
                           ZN => n3672);
   U3486 : AND2_X1 port map( A1 => n6207, A2 => n6208, ZN => n1890);
   U3487 : OR2_X1 port map( A1 => n4449, A2 => n5107, ZN => n3453);
   U3488 : OR2_X1 port map( A1 => n5188, A2 => n5675, ZN => n2978);
   U3489 : AOI21_X1 port map( B1 => n5969, B2 => n5973, A => n971, ZN => n5977)
                           ;
   U3490 : OR2_X1 port map( A1 => n5044, A2 => n5045, ZN => n4444);
   U3491 : OR2_X1 port map( A1 => n4048, A2 => n5100, ZN => n4076);
   U3492 : NAND2_X1 port map( A1 => n2870, A2 => n2873, ZN => n5845);
   U3493 : XNOR2_X1 port map( A => n3513, B => n6786, ZN => n7098);
   U3494 : INV_X1 port map( A => n6687, ZN => n3513);
   U3495 : OR2_X1 port map( A1 => n5495, A2 => n5494, ZN => n2099);
   U3496 : OR2_X1 port map( A1 => n5683, A2 => n5682, ZN => n5477);
   U3497 : NAND2_X1 port map( A1 => n2640, A2 => n3351, ZN => n2639);
   U3498 : OR2_X1 port map( A1 => n5855, A2 => n6159, ZN => n4403);
   U3499 : NOR2_X1 port map( A1 => n6193, A2 => n6192, ZN => n2869);
   U3500 : INV_X1 port map( A => n6016, ZN => n5826);
   U3501 : OR2_X1 port map( A1 => n4239, A2 => n4383, ZN => n2214);
   U3502 : OAI21_X1 port map( B1 => n7622, B2 => n8068, A => n19901, ZN => 
                           n2386);
   U3503 : INV_X1 port map( A => n8184, ZN => n2649);
   U3504 : OR2_X1 port map( A1 => n5474, A2 => n5475, ZN => n1885);
   U3505 : INV_X1 port map( A => n6072, ZN => n3999);
   U3506 : OR2_X1 port map( A1 => n5216, A2 => n5360, ZN => n1947);
   U3508 : XNOR2_X1 port map( A => n1081, B => n6985, ZN => n7377);
   U3509 : XNOR2_X1 port map( A => n6776, B => n6641, ZN => n7238);
   U3510 : OAI211_X1 port map( C1 => n5993, C2 => n5818, A => n3469, B => n3467
                           , ZN => n6947);
   U3511 : OR2_X1 port map( A1 => n3319, A2 => n6068, ZN => n1982);
   U3512 : AND2_X1 port map( A1 => n1958, A2 => n1274, ZN => n1957);
   U3513 : AND2_X1 port map( A1 => n6206, A2 => n287, ZN => n5838);
   U3515 : OR2_X1 port map( A1 => n5752, A2 => n5753, ZN => n2294);
   U3516 : OR2_X1 port map( A1 => n5320, A2 => n3319, ZN => n6071);
   U3517 : INV_X1 port map( A => n8720, ZN => n2756);
   U3518 : AND2_X1 port map( A1 => n20154, A2 => n1560, ZN => n7408);
   U3519 : OR2_X1 port map( A1 => n7096, A2 => n20154, ZN => n7407);
   U3520 : AND3_X1 port map( A1 => n7642, A2 => n7641, A3 => n7640, ZN => n2238
                           );
   U3521 : INV_X1 port map( A => n8347, ZN => n8271);
   U3522 : OR2_X1 port map( A1 => n6618, A2 => n8095, ZN => n1962);
   U3523 : INV_X1 port map( A => n9623, ZN => n10231);
   U3525 : INV_X1 port map( A => n9006, ZN => n8622);
   U3526 : OR2_X1 port map( A1 => n9007, A2 => n9008, ZN => n1484);
   U3528 : OR2_X1 port map( A1 => n9346, A2 => n8156, ZN => n8700);
   U3529 : OR2_X1 port map( A1 => n2727, A2 => n9210, ZN => n1326);
   U3530 : OR2_X1 port map( A1 => n9252, A2 => n9251, ZN => n1616);
   U3531 : INV_X1 port map( A => n8748, ZN => n8747);
   U3533 : INV_X1 port map( A => n9287, ZN => n8577);
   U3534 : OR2_X1 port map( A1 => n8727, A2 => n8961, ZN => n2850);
   U3535 : INV_X1 port map( A => n7668, ZN => n8336);
   U3536 : AOI21_X1 port map( B1 => n8728, B2 => n2955, A => n8731, ZN => n9382
                           );
   U3537 : AND2_X1 port map( A1 => n9121, A2 => n1233, ZN => n8553);
   U3539 : AND2_X1 port map( A1 => n9333, A2 => n9331, ZN => n9075);
   U3540 : OR2_X1 port map( A1 => n9122, A2 => n8552, ZN => n9127);
   U3541 : OR2_X1 port map( A1 => n9173, A2 => n9176, ZN => n2618);
   U3542 : OAI211_X1 port map( C1 => n9451, C2 => n6442, A => n6441, B => n6440
                           , ZN => n9957);
   U3543 : NAND2_X1 port map( A1 => n2690, A2 => n8651, ZN => n10351);
   U3544 : OR2_X1 port map( A1 => n8660, A2 => n8995, ZN => n3552);
   U3545 : XNOR2_X1 port map( A => n10171, B => n19853, ZN => n1283);
   U3546 : XNOR2_X1 port map( A => n9977, B => n9596, ZN => n1284);
   U3547 : XNOR2_X1 port map( A => n10472, B => n875, ZN => n9596);
   U3548 : XNOR2_X1 port map( A => n9646, B => n9991, ZN => n10348);
   U3549 : XNOR2_X1 port map( A => n9940, B => n9939, ZN => n10882);
   U3550 : INV_X1 port map( A => n9054, ZN => n1761);
   U3551 : NAND2_X1 port map( A1 => n8888, A2 => n1030, ZN => n9429);
   U3552 : OR2_X1 port map( A1 => n8889, A2 => n9451, ZN => n1030);
   U3553 : INV_X1 port map( A => n11378, ZN => n2611);
   U3554 : BUF_X1 port map( A => n10856, Z => n11331);
   U3555 : OR2_X1 port map( A1 => n8795, A2 => n9217, ZN => n8670);
   U3556 : AOI21_X1 port map( B1 => n1830, B2 => n8995, A => n1829, ZN => n8442
                           );
   U3557 : AND2_X1 port map( A1 => n8998, A2 => n8997, ZN => n1829);
   U3559 : OR2_X1 port map( A1 => n8420, A2 => n8445, ZN => n8444);
   U3560 : OR2_X1 port map( A1 => n9264, A2 => n9271, ZN => n1321);
   U3561 : INV_X1 port map( A => n9583, ZN => n9582);
   U3562 : XNOR2_X1 port map( A => n10617, B => n3812, ZN => n11489);
   U3563 : OR2_X1 port map( A1 => n7897, A2 => n8649, ZN => n7900);
   U3564 : OR2_X1 port map( A1 => n8818, A2 => n8817, ZN => n1964);
   U3565 : OR2_X1 port map( A1 => n8785, A2 => n9149, ZN => n8788);
   U3566 : INV_X1 port map( A => n9600, ZN => n8769);
   U3567 : INV_X1 port map( A => n10163, ZN => n8450);
   U3568 : INV_X1 port map( A => n9697, ZN => n9587);
   U3569 : INV_X1 port map( A => n9430, ZN => n9967);
   U3570 : INV_X1 port map( A => n9429, ZN => n10304);
   U3571 : OAI211_X1 port map( C1 => n8814, C2 => n8815, A => n8813, B => n2752
                           , ZN => n8456);
   U3572 : NOR2_X1 port map( A1 => n9546, A2 => n11412, ZN => n3617);
   U3574 : OAI21_X1 port map( B1 => n2611, B2 => n11331, A => n11375, ZN => 
                           n2610);
   U3575 : XNOR2_X1 port map( A => n2570, B => n9608, ZN => n3588);
   U3576 : OR2_X1 port map( A1 => n11460, A2 => n11880, ZN => n10246);
   U3577 : NOR2_X1 port map( A1 => n11093, A2 => n11446, ZN => n11204);
   U3578 : AOI21_X1 port map( B1 => n11233, B2 => n11366, A => n1600, ZN => 
                           n11252);
   U3579 : INV_X1 port map( A => n3482, ZN => n3481);
   U3580 : AND2_X1 port map( A1 => n11489, A2 => n11493, ZN => n2135);
   U3581 : NOR2_X1 port map( A1 => n11952, A2 => n11598, ZN => n11658);
   U3582 : OR2_X1 port map( A1 => n10998, A2 => n10999, ZN => n2234);
   U3584 : INV_X1 port map( A => n12207, ZN => n3692);
   U3585 : OR2_X1 port map( A1 => n11401, A2 => n2724, ZN => n1460);
   U3586 : INV_X1 port map( A => n11683, ZN => n12577);
   U3590 : INV_X1 port map( A => n11942, ZN => n12439);
   U3591 : AND2_X1 port map( A1 => n11942, A2 => n12110, ZN => n11938);
   U3592 : INV_X1 port map( A => n12606, ZN => n12603);
   U3593 : OR2_X1 port map( A1 => n11323, A2 => n11324, ZN => n10806);
   U3595 : BUF_X1 port map( A => n13451, Z => n12859);
   U3596 : NOR2_X1 port map( A1 => n20363, A2 => n924, ZN => n3811);
   U3598 : OR2_X1 port map( A1 => n12416, A2 => n11602, ZN => n2760);
   U3599 : AND2_X1 port map( A1 => n246, A2 => n180, ZN => n3405);
   U3600 : INV_X1 port map( A => n12429, ZN => n12685);
   U3601 : OAI21_X1 port map( B1 => n1547, B2 => n11642, A => n1546, ZN => 
                           n11705);
   U3602 : XNOR2_X1 port map( A => n13596, B => n13715, ZN => n13204);
   U3603 : INV_X1 port map( A => n12041, ZN => n12283);
   U3605 : INV_X1 port map( A => n924, ZN => n3164);
   U3606 : XNOR2_X1 port map( A => n13103, B => n13383, ZN => n13631);
   U3607 : NOR2_X1 port map( A1 => n11194, A2 => n3234, ZN => n11195);
   U3608 : OAI21_X1 port map( B1 => n11618, B2 => n11897, A => n11896, ZN => 
                           n13686);
   U3609 : AND2_X1 port map( A1 => n248, A2 => n12568, ZN => n11893);
   U3610 : OR2_X1 port map( A1 => n11173, A2 => n10912, ZN => n3360);
   U3611 : AOI21_X1 port map( B1 => n11210, B2 => n11480, A => n2536, ZN => 
                           n11215);
   U3613 : XNOR2_X1 port map( A => n12745, B => n13634, ZN => n12996);
   U3614 : XNOR2_X1 port map( A => n13677, B => n13833, ZN => n13433);
   U3616 : XNOR2_X1 port map( A => n12713, B => n13330, ZN => n2947);
   U3617 : OR2_X1 port map( A1 => n14790, A2 => n14787, ZN => n14102);
   U3618 : OR2_X1 port map( A1 => n14775, A2 => n14781, ZN => n13905);
   U3619 : OR2_X1 port map( A1 => n13270, A2 => n13275, ZN => n1304);
   U3620 : OR2_X1 port map( A1 => n11627, A2 => n12237, ZN => n3754);
   U3621 : OR2_X1 port map( A1 => n11628, A2 => n12237, ZN => n2910);
   U3622 : INV_X1 port map( A => n13335, ZN => n2312);
   U3623 : OR2_X1 port map( A1 => n14556, A2 => n14554, ZN => n2125);
   U3624 : OAI211_X1 port map( C1 => n11030, C2 => n12355, A => n3278, B => 
                           n1637, ZN => n3276);
   U3625 : INV_X1 port map( A => n2748, ZN => n14275);
   U3626 : INV_X1 port map( A => n19781, ZN => n1295);
   U3627 : XNOR2_X1 port map( A => n2657, B => n12913, ZN => n3236);
   U3628 : AND2_X1 port map( A1 => n12321, A2 => n2838, ZN => n14850);
   U3629 : NOR2_X1 port map( A1 => n14623, A2 => n19875, ZN => n15316);
   U3630 : INV_X1 port map( A => n19906, ZN => n14612);
   U3631 : INV_X1 port map( A => n14268, ZN => n14740);
   U3632 : INV_X1 port map( A => n14693, ZN => n1104);
   U3633 : NOR2_X1 port map( A1 => n14935, A2 => n15504, ZN => n3778);
   U3634 : NOR2_X1 port map( A1 => n14641, A2 => n14637, ZN => n14635);
   U3635 : INV_X1 port map( A => n14148, ZN => n14237);
   U3636 : OR2_X1 port map( A1 => n14497, A2 => n1089, ZN => n1876);
   U3637 : AND2_X1 port map( A1 => n2748, A2 => n14566, ZN => n14276);
   U3638 : AND2_X1 port map( A1 => n14673, A2 => n13981, ZN => n14263);
   U3639 : INV_X1 port map( A => n14746, ZN => n3158);
   U3640 : AND2_X1 port map( A1 => n15906, A2 => n2723, ZN => n2722);
   U3641 : INV_X1 port map( A => n19986, ZN => n13913);
   U3642 : OR2_X1 port map( A1 => n14828, A2 => n14826, ZN => n13914);
   U3643 : AND2_X1 port map( A1 => n13904, A2 => n3697, ZN => n3696);
   U3645 : OR2_X1 port map( A1 => n14728, A2 => n986, ZN => n1642);
   U3646 : OR2_X1 port map( A1 => n14644, A2 => n12973, ZN => n13986);
   U3647 : NOR2_X1 port map( A1 => n15378, A2 => n14874, ZN => n14875);
   U3648 : XNOR2_X1 port map( A => n1809, B => n12672, ZN => n14420);
   U3649 : XNOR2_X1 port map( A => n12678, B => n12677, ZN => n14052);
   U3650 : OR2_X1 port map( A1 => n20147, A2 => n15409, ZN => n2129);
   U3651 : OR2_X1 port map( A1 => n15544, A2 => n15070, ZN => n2800);
   U3652 : INV_X1 port map( A => n15608, ZN => n3427);
   U3653 : OR2_X1 port map( A1 => n15615, A2 => n15071, ZN => n15407);
   U3654 : INV_X1 port map( A => n17128, ZN => n3273);
   U3655 : OAI211_X1 port map( C1 => n14691, C2 => n19895, A => n14693, B => 
                           n2094, ZN => n2186);
   U3656 : INV_X1 port map( A => n15625, ZN => n15836);
   U3657 : OR2_X1 port map( A1 => n15914, A2 => n15915, ZN => n1152);
   U3658 : INV_X1 port map( A => n15409, ZN => n15413);
   U3659 : AND2_X1 port map( A1 => n14514, A2 => n14323, ZN => n3149);
   U3660 : INV_X1 port map( A => n15353, ZN => n1155);
   U3661 : OR2_X1 port map( A1 => n198, A2 => n20178, ZN => n15715);
   U3662 : OR2_X1 port map( A1 => n15870, A2 => n15709, ZN => n15711);
   U3663 : OAI21_X1 port map( B1 => n2674, B2 => n2677, A => n2673, ZN => 
                           n15712);
   U3664 : INV_X1 port map( A => n2678, ZN => n2674);
   U3665 : NOR2_X1 port map( A1 => n18105, A2 => n17954, ZN => n2661);
   U3666 : OR2_X1 port map( A1 => n14016, A2 => n14015, ZN => n2110);
   U3667 : INV_X1 port map( A => n17946, ZN => n3475);
   U3668 : NOR2_X1 port map( A1 => n15030, A2 => n15380, ZN => n2988);
   U3669 : NOR2_X1 port map( A1 => n16373, A2 => n2385, ZN => n16051);
   U3670 : AND2_X1 port map( A1 => n16373, A2 => n2385, ZN => n16052);
   U3671 : INV_X1 port map( A => n2216, ZN => n3102);
   U3673 : OR2_X1 port map( A1 => n19891, A2 => n15828, ZN => n14581);
   U3675 : OR2_X1 port map( A1 => n17511, A2 => n16633, ZN => n2335);
   U3676 : OAI21_X1 port map( B1 => n20240, B2 => n19352, A => n2668, ZN => 
                           n16638);
   U3677 : AND2_X1 port map( A1 => n20436, A2 => n17238, ZN => n3485);
   U3678 : OR2_X1 port map( A1 => n19647, A2 => n20436, ZN => n3486);
   U3681 : OAI21_X1 port map( B1 => n17492, B2 => n17491, A => n17155, ZN => 
                           n17158);
   U3682 : INV_X1 port map( A => n18131, ZN => n17777);
   U3683 : AND2_X1 port map( A1 => n20101, A2 => n19744, ZN => n17449);
   U3684 : BUF_X1 port map( A => n18138, Z => n18264);
   U3685 : XNOR2_X1 port map( A => n1529, B => n1528, ZN => n17981);
   U3686 : XNOR2_X1 port map( A => n17297, B => n17301, ZN => n1528);
   U3687 : XNOR2_X1 port map( A => n1417, B => n17290, ZN => n3207);
   U3688 : NOR2_X1 port map( A1 => n225, A2 => n18016, ZN => n18979);
   U3689 : XNOR2_X1 port map( A => n16138, B => n16137, ZN => n16731);
   U3692 : INV_X1 port map( A => n3287, ZN => n3150);
   U3693 : XNOR2_X1 port map( A => n2994, B => n16825, ZN => n2991);
   U3694 : XNOR2_X1 port map( A => n17355, B => n3749, ZN => n2993);
   U3695 : AND2_X1 port map( A1 => n17069, A2 => n19707, ZN => n17184);
   U3696 : INV_X1 port map( A => n17887, ZN => n1907);
   U3697 : AND2_X1 port map( A1 => n17536, A2 => n17537, ZN => n3535);
   U3698 : INV_X1 port map( A => n16465, ZN => n1115);
   U3699 : OR2_X1 port map( A1 => n17211, A2 => n20092, ZN => n1395);
   U3700 : OR2_X1 port map( A1 => n20111, A2 => n18392, ZN => n3455);
   U3701 : NAND2_X1 port map( A1 => n20111, A2 => n2793, ZN => n1733);
   U3703 : INV_X1 port map( A => n18078, ZN => n1728);
   U3704 : INV_X1 port map( A => n19352, ZN => n2669);
   U3705 : NAND2_X1 port map( A1 => n16468, A2 => n17507, ZN => n3080);
   U3706 : OAI21_X1 port map( B1 => n17214, B2 => n2841, A => n20135, ZN => 
                           n1844);
   U3707 : NOR2_X1 port map( A1 => n16249, A2 => n16248, ZN => n18501);
   U3712 : AND2_X1 port map( A1 => n17789, A2 => n1668, ZN => n19157);
   U3713 : OAI21_X1 port map( B1 => n17596, B2 => n16657, A => n16656, ZN => 
                           n19452);
   U3714 : OR2_X1 port map( A1 => n3078, A2 => n4952, ZN => n4910);
   U3715 : NOR2_X1 port map( A1 => n5018, A2 => n4555, ZN => n3683);
   U3716 : INV_X1 port map( A => n5520, ZN => n3410);
   U3717 : AND2_X1 port map( A1 => n19789, A2 => n6027, ZN => n5030);
   U3718 : OR2_X1 port map( A1 => n4355, A2 => n4601, ZN => n3095);
   U3719 : INV_X1 port map( A => n6101, ZN => n5664);
   U3721 : OR2_X1 port map( A1 => n4482, A2 => n4965, ZN => n4481);
   U3724 : INV_X1 port map( A => n4960, ZN => n3657);
   U3725 : INV_X1 port map( A => n5023, ZN => n4765);
   U3726 : OR2_X1 port map( A1 => n1232, A2 => n5073, ZN => n3838);
   U3727 : NOR2_X1 port map( A1 => n6171, A2 => n6168, ZN => n2434);
   U3728 : AND2_X1 port map( A1 => n6172, A2 => n6171, ZN => n2435);
   U3729 : INV_X1 port map( A => n6172, ZN => n2629);
   U3730 : OR2_X1 port map( A1 => n4840, A2 => n4656, ZN => n3980);
   U3731 : AND2_X1 port map( A1 => n6202, A2 => n6201, ZN => n1891);
   U3732 : OR2_X1 port map( A1 => n5363, A2 => n5364, ZN => n5464);
   U3733 : INV_X1 port map( A => n5631, ZN => n5467);
   U3734 : INV_X1 port map( A => n6118, ZN => n3483);
   U3735 : OR2_X1 port map( A1 => n5387, A2 => n6124, ZN => n2093);
   U3736 : INV_X1 port map( A => n6050, ZN => n5138);
   U3737 : INV_X1 port map( A => n5471, ZN => n5475);
   U3738 : INV_X1 port map( A => n5569, ZN => n6033);
   U3739 : AND2_X1 port map( A1 => n5676, A2 => n5279, ZN => n3128);
   U3740 : INV_X1 port map( A => n5628, ZN => n5632);
   U3741 : INV_X1 port map( A => n5930, ZN => n3434);
   U3743 : INV_X1 port map( A => n5930, ZN => n5929);
   U3744 : OR2_X1 port map( A1 => n5899, A2 => n3098, ZN => n3096);
   U3745 : INV_X1 port map( A => n5201, ZN => n1695);
   U3746 : AND2_X1 port map( A1 => n3802, A2 => n5218, ZN => n1465);
   U3747 : OR2_X1 port map( A1 => n4745, A2 => n5005, ZN => n4748);
   U3748 : OAI21_X1 port map( B1 => n6166, B2 => n1867, A => n6172, ZN => n1866
                           );
   U3749 : OR2_X1 port map( A1 => n4737, A2 => n4736, ZN => n3008);
   U3750 : NOR2_X1 port map( A1 => n3606, A2 => n3605, ZN => n3608);
   U3751 : OR2_X1 port map( A1 => n5570, A2 => n5569, ZN => n2377);
   U3752 : INV_X1 port map( A => n3188, ZN => n6148);
   U3754 : NOR2_X1 port map( A1 => n6138, A2 => n5859, ZN => n5864);
   U3755 : OR2_X1 port map( A1 => n4507, A2 => n4370, ZN => n3907);
   U3757 : AND2_X1 port map( A1 => n4305, A2 => n2490, ZN => n4124);
   U3758 : OR2_X1 port map( A1 => n4087, A2 => n19562, ZN => n2136);
   U3759 : OR2_X1 port map( A1 => n5279, A2 => n2719, ZN => n2718);
   U3760 : INV_X1 port map( A => n5444, ZN => n5647);
   U3761 : INV_X1 port map( A => n2557, ZN => n6742);
   U3762 : AND2_X1 port map( A1 => n6067, A2 => n6068, ZN => n2286);
   U3763 : AND2_X1 port map( A1 => n5803, A2 => n6189, ZN => n1986);
   U3765 : INV_X1 port map( A => n6022, ZN => n5447);
   U3766 : AND2_X1 port map( A1 => n3418, A2 => n9300, ZN => n2985);
   U3767 : OR2_X1 port map( A1 => n7974, A2 => n7972, ZN => n2176);
   U3768 : OR2_X1 port map( A1 => n5397, A2 => n5251, ZN => n5399);
   U3770 : OR2_X1 port map( A1 => n5826, A2 => n1096, ZN => n1095);
   U3771 : OR2_X1 port map( A1 => n6175, A2 => n170, ZN => n6177);
   U3772 : INV_X1 port map( A => n8284, ZN => n3660);
   U3773 : OR2_X1 port map( A1 => n5235, A2 => n1746, ZN => n1745);
   U3774 : NOR2_X1 port map( A1 => n5793, A2 => n5429, ZN => n2880);
   U3775 : OR2_X1 port map( A1 => n7990, A2 => n7096, ZN => n8013);
   U3776 : OR2_X1 port map( A1 => n8014, A2 => n7096, ZN => n7828);
   U3777 : OR2_X1 port map( A1 => n8070, A2 => n7420, ZN => n2379);
   U3778 : OR2_X1 port map( A1 => n6023, A2 => n6022, ZN => n1483);
   U3779 : INV_X1 port map( A => n6046, ZN => n5777);
   U3780 : AND2_X1 port map( A1 => n8271, A2 => n8272, ZN => n1608);
   U3781 : NAND3_X1 port map( A1 => n1568, A2 => n5384, A3 => n1570, ZN => 
                           n7065);
   U3782 : OR2_X1 port map( A1 => n5385, A2 => n19475, ZN => n1570);
   U3784 : OR2_X1 port map( A1 => n5870, A2 => n6124, ZN => n2175);
   U3785 : OR2_X1 port map( A1 => n7930, A2 => n2030, ZN => n1402);
   U3786 : XNOR2_X1 port map( A => n5337, B => n6630, ZN => n7600);
   U3787 : INV_X1 port map( A => n8132, ZN => n7497);
   U3788 : INV_X1 port map( A => n8220, ZN => n3655);
   U3789 : XNOR2_X1 port map( A => n3068, B => n7304, ZN => n3067);
   U3792 : INV_X1 port map( A => n8114, ZN => n1143);
   U3793 : AND2_X1 port map( A1 => n8060, A2 => n8062, ZN => n4730);
   U3794 : AND2_X1 port map( A1 => n8344, A2 => n8341, ZN => n3122);
   U3795 : AND2_X1 port map( A1 => n8239, A2 => n8238, ZN => n2987);
   U3796 : OR2_X1 port map( A1 => n7432, A2 => n2687, ZN => n7433);
   U3797 : AND2_X1 port map( A1 => n7416, A2 => n8068, ZN => n8793);
   U3798 : INV_X1 port map( A => n8603, ZN => n8952);
   U3799 : INV_X1 port map( A => n7898, ZN => n1405);
   U3800 : OR2_X1 port map( A1 => n7618, A2 => n8204, ZN => n1410);
   U3801 : AOI21_X1 port map( B1 => n266, B2 => n9241, A => n6587, ZN => n2476)
                           ;
   U3802 : INV_X1 port map( A => n9129, ZN => n8805);
   U3803 : INV_X1 port map( A => n7445, ZN => n8281);
   U3804 : INV_X1 port map( A => n8068, ZN => n8181);
   U3806 : INV_X1 port map( A => n8354, ZN => n7695);
   U3807 : AND2_X1 port map( A1 => n6750, A2 => n8142, ZN => n1197);
   U3808 : OAI21_X1 port map( B1 => n8264, B2 => n8262, A => n3765, ZN => n6701
                           );
   U3809 : OAI21_X1 port map( B1 => n7556, B2 => n1791, A => n7558, ZN => n8500
                           );
   U3810 : OR2_X1 port map( A1 => n7678, A2 => n8363, ZN => n3491);
   U3811 : OAI21_X1 port map( B1 => n8264, B2 => n8261, A => n8263, ZN => n3597
                           );
   U3812 : AND2_X1 port map( A1 => n8420, A2 => n9210, ZN => n8803);
   U3813 : OR2_X1 port map( A1 => n8111, A2 => n8098, ZN => n7436);
   U3814 : INV_X1 port map( A => n8248, ZN => n3312);
   U3815 : OR2_X1 port map( A1 => n8250, A2 => n8248, ZN => n3311);
   U3816 : OAI22_X1 port map( A1 => n1810, A2 => n8294, B1 => n7469, B2 => 
                           n8031, ZN => n8811);
   U3817 : AND2_X1 port map( A1 => n7469, A2 => n7471, ZN => n1810);
   U3818 : INV_X1 port map( A => n1560, ZN => n8015);
   U3819 : AND2_X1 port map( A1 => n7466, A2 => n7811, ZN => n7467);
   U3820 : AND2_X1 port map( A1 => n9210, A2 => n9135, ZN => n1324);
   U3821 : INV_X1 port map( A => n1567, ZN => n8515);
   U3822 : AND2_X1 port map( A1 => n8140, A2 => n8347, ZN => n3250);
   U3823 : NOR2_X1 port map( A1 => n8140, A2 => n8352, ZN => n8270);
   U3824 : INV_X1 port map( A => n9357, ZN => n1204);
   U3825 : OR2_X1 port map( A1 => n9359, A2 => n9528, ZN => n1201);
   U3826 : OR2_X1 port map( A1 => n9215, A2 => n9214, ZN => n1333);
   U3827 : NOR2_X1 port map( A1 => n9176, A2 => n8761, ZN => n8693);
   U3828 : XNOR2_X1 port map( A => n9934, B => n6461, ZN => n9935);
   U3829 : INV_X1 port map( A => n9105, ZN => n8779);
   U3830 : NOR2_X1 port map( A1 => n8077, A2 => n3795, ZN => n3794);
   U3831 : INV_X1 port map( A => n9266, ZN => n1587);
   U3833 : OR2_X1 port map( A1 => n8998, A2 => n8772, ZN => n1831);
   U3834 : AND2_X1 port map( A1 => n7408, A2 => n7826, ZN => n2405);
   U3835 : AND2_X1 port map( A1 => n8272, A2 => n8349, ZN => n1607);
   U3836 : INV_X1 port map( A => n6656, ZN => n9190);
   U3838 : INV_X1 port map( A => n9453, ZN => n8565);
   U3839 : OR2_X1 port map( A1 => n7863, A2 => n1502, ZN => n1499);
   U3840 : OR2_X1 port map( A1 => n8146, A2 => n8145, ZN => n8147);
   U3841 : OR2_X1 port map( A1 => n8708, A2 => n1037, ZN => n9182);
   U3842 : INV_X1 port map( A => n1032, ZN => n10016);
   U3843 : BUF_X1 port map( A => n8550, Z => n8818);
   U3844 : AND2_X1 port map( A1 => n9262, A2 => n9266, ZN => n8771);
   U3847 : INV_X1 port map( A => n1037, ZN => n2653);
   U3848 : AND2_X1 port map( A1 => n8708, A2 => n1037, ZN => n8630);
   U3850 : INV_X1 port map( A => n7562, ZN => n7564);
   U3851 : OR2_X1 port map( A1 => n9300, A2 => n9018, ZN => n9019);
   U3852 : INV_X1 port map( A => n8846, ZN => n9298);
   U3853 : INV_X1 port map( A => n9624, ZN => n9978);
   U3854 : AND2_X1 port map( A1 => n9836, A2 => n2749, ZN => n8467);
   U3855 : AND2_X1 port map( A1 => n9305, A2 => n9228, ZN => n1752);
   U3856 : INV_X1 port map( A => n20011, ZN => n1754);
   U3857 : INV_X1 port map( A => n8500, ZN => n9363);
   U3858 : INV_X1 port map( A => n8961, ZN => n8726);
   U3859 : OR2_X1 port map( A1 => n7659, A2 => n9038, ZN => n2336);
   U3861 : INV_X1 port map( A => n8729, ZN => n8939);
   U3862 : AND2_X1 port map( A1 => n20146, A2 => n9129, ZN => n9202);
   U3863 : INV_X1 port map( A => n9201, ZN => n8665);
   U3864 : AND2_X1 port map( A1 => n9130, A2 => n9201, ZN => n9782);
   U3865 : INV_X1 port map( A => n8812, ZN => n8552);
   U3866 : OR2_X1 port map( A1 => n7477, A2 => n7476, ZN => n3609);
   U3867 : OR2_X1 port map( A1 => n8815, A2 => n8812, ZN => n2752);
   U3868 : OR2_X1 port map( A1 => n3518, A2 => n7752, ZN => n1401);
   U3869 : INV_X1 port map( A => n8124, ZN => n3520);
   U3872 : INV_X1 port map( A => n10805, ZN => n10802);
   U3873 : MUX2_X1 port map( A => n9455, B => n9454, S => n9453, Z => n9868);
   U3874 : AND2_X1 port map( A1 => n10649, A2 => n10945, ZN => n11156);
   U3875 : OR2_X1 port map( A1 => n10960, A2 => n10701, ZN => n9614);
   U3876 : XNOR2_X1 port map( A => n9429, B => n9430, ZN => n1029);
   U3877 : OR2_X1 port map( A1 => n10971, A2 => n11162, ZN => n3487);
   U3878 : NOR2_X1 port map( A1 => n2498, A2 => n9145, ZN => n7942);
   U3879 : OR2_X1 port map( A1 => n11430, A2 => n11428, ZN => n1970);
   U3880 : XNOR2_X1 port map( A => n10496, B => n10495, ZN => n10783);
   U3881 : INV_X1 port map( A => n11440, ZN => n2272);
   U3882 : INV_X1 port map( A => n9960, ZN => n2506);
   U3883 : XNOR2_X1 port map( A => n9778, B => n1032, ZN => n9860);
   U3884 : XNOR2_X1 port map( A => n9389, B => n9390, ZN => n10946);
   U3885 : OR2_X1 port map( A1 => n9381, A2 => n9382, ZN => n9383);
   U3886 : NOR2_X1 port map( A1 => n247, A2 => n12209, ZN => n2713);
   U3887 : OR2_X1 port map( A1 => n204, A2 => n3507, ZN => n3712);
   U3888 : INV_X1 port map( A => n11383, ZN => n1330);
   U3889 : INV_X1 port map( A => n12212, ZN => n12067);
   U3890 : AND2_X1 port map( A1 => n12208, A2 => n247, ZN => n1879);
   U3891 : OAI21_X1 port map( B1 => n11463, B2 => n11886, A => n11462, ZN => 
                           n12168);
   U3893 : OR2_X1 port map( A1 => n11460, A2 => n11120, ZN => n11124);
   U3894 : OR2_X1 port map( A1 => n11256, A2 => n191, ZN => n10805);
   U3895 : INV_X1 port map( A => n10783, ZN => n11438);
   U3896 : NOR2_X1 port map( A1 => n12084, A2 => n12422, ZN => n2761);
   U3897 : AND2_X1 port map( A1 => n12639, A2 => n12449, ZN => n12638);
   U3898 : XNOR2_X1 port map( A => n9850, B => n9849, ZN => n11365);
   U3899 : XNOR2_X1 port map( A => n9853, B => n9855, ZN => n2744);
   U3900 : INV_X1 port map( A => n11322, ZN => n1124);
   U3902 : INV_X1 port map( A => n12636, ZN => n2256);
   U3903 : NOR2_X1 port map( A1 => n11562, A2 => n11561, ZN => n11563);
   U3904 : OR2_X1 port map( A1 => n12274, A2 => n12273, ZN => n11748);
   U3905 : INV_X1 port map( A => n2605, ZN => n2604);
   U3906 : OAI21_X1 port map( B1 => n2606, B2 => n2610, A => n10858, ZN => 
                           n2605);
   U3907 : BUF_X1 port map( A => n11709, Z => n12153);
   U3908 : INV_X1 port map( A => n12211, ZN => n12206);
   U3909 : INV_X1 port map( A => n11011, ZN => n3382);
   U3910 : INV_X1 port map( A => n11513, ZN => n11509);
   U3912 : AND4_X1 port map( A1 => n3488, A2 => n3489, A3 => n10949, A4 => 
                           n3487, ZN => n11761);
   U3913 : INV_X1 port map( A => n11539, ZN => n11532);
   U3914 : INV_X1 port map( A => n12282, ZN => n11582);
   U3915 : XNOR2_X1 port map( A => n6657, B => n6658, ZN => n1523);
   U3917 : OR2_X1 port map( A1 => n2610, A2 => n2606, ZN => n2607);
   U3918 : OR2_X1 port map( A1 => n11889, A2 => n11890, ZN => n3732);
   U3919 : OR2_X1 port map( A1 => n11042, A2 => n11041, ZN => n10192);
   U3920 : OR2_X1 port map( A1 => n12041, A2 => n12280, ZN => n1299);
   U3921 : AND2_X1 port map( A1 => n1387, A2 => n3676, ZN => n1414);
   U3922 : INV_X1 port map( A => n3617, ZN => n3614);
   U3923 : INV_X1 port map( A => n10756, ZN => n11523);
   U3924 : INV_X1 port map( A => n10742, ZN => n11572);
   U3925 : AND2_X1 port map( A1 => n11365, A2 => n11230, ZN => n10679);
   U3926 : INV_X1 port map( A => n10677, ZN => n11366);
   U3927 : NOR2_X1 port map( A1 => n10851, A2 => n11231, ZN => n11364);
   U3928 : INV_X1 port map( A => n19878, ZN => n3361);
   U3929 : INV_X1 port map( A => n2598, ZN => n2160);
   U3930 : NAND2_X1 port map( A1 => n2043, A2 => n10861, ZN => n12240);
   U3931 : AND2_X1 port map( A1 => n12554, A2 => n12542, ZN => n11795);
   U3932 : INV_X1 port map( A => n12440, ZN => n11939);
   U3933 : AOI21_X1 port map( B1 => n10871, B2 => n20235, A => n10870, ZN => 
                           n12617);
   U3934 : INV_X1 port map( A => n12269, ZN => n12020);
   U3935 : OR2_X1 port map( A1 => n2707, A2 => n12002, ZN => n3241);
   U3936 : AND2_X1 port map( A1 => n12250, A2 => n11733, ZN => n1139);
   U3937 : INV_X1 port map( A => n11717, ZN => n11776);
   U3939 : AOI21_X1 port map( B1 => n10310, B2 => n11254, A => n11327, ZN => 
                           n10312);
   U3940 : AND2_X1 port map( A1 => n3733, A2 => n12261, ZN => n1366);
   U3941 : OR2_X1 port map( A1 => n12374, A2 => n12373, ZN => n12375);
   U3942 : OR2_X1 port map( A1 => n10737, A2 => n19915, ZN => n10739);
   U3943 : OR2_X1 port map( A1 => n11599, A2 => n1578, ZN => n3633);
   U3944 : INV_X1 port map( A => n12273, ZN => n12298);
   U3945 : INV_X1 port map( A => n12274, ZN => n11781);
   U3946 : AND2_X1 port map( A1 => n12648, A2 => n12686, ZN => n12646);
   U3947 : NOR2_X1 port map( A1 => n3601, A2 => n1330, ZN => n12105);
   U3948 : OR2_X1 port map( A1 => n10900, A2 => n11210, ZN => n2898);
   U3950 : OR2_X1 port map( A1 => n10961, A2 => n10960, ZN => n1673);
   U3951 : AND2_X1 port map( A1 => n11761, A2 => n11586, ZN => n1735);
   U3952 : OAI211_X1 port map( C1 => n10829, C2 => n11131, A => n11418, B => 
                           n11051, ZN => n10413);
   U3953 : OR2_X1 port map( A1 => n10372, A2 => n11456, ZN => n1307);
   U3954 : OR2_X1 port map( A1 => n12002, A2 => n12354, ZN => n3278);
   U3955 : AND2_X1 port map( A1 => n11399, A2 => n2724, ZN => n9747);
   U3958 : OR2_X1 port map( A1 => n10924, A2 => n11526, ZN => n2522);
   U3959 : INV_X1 port map( A => n1260, ZN => n13790);
   U3960 : INV_X1 port map( A => n11646, ZN => n1952);
   U3961 : OR2_X1 port map( A1 => n11603, A2 => n12417, ZN => n12083);
   U3962 : NOR2_X1 port map( A1 => n12103, A2 => n11380, ZN => n1280);
   U3963 : OAI21_X1 port map( B1 => n10674, B2 => n10673, A => n10672, ZN => 
                           n12437);
   U3964 : INV_X1 port map( A => n13199, ZN => n2657);
   U3965 : OR2_X1 port map( A1 => n631, A2 => n14800, ZN => n12321);
   U3966 : XNOR2_X1 port map( A => n20155, B => n6461, ZN => n2518);
   U3967 : INV_X1 port map( A => n14420, ZN => n1808);
   U3968 : AND2_X1 port map( A1 => n12295, A2 => n20363, ZN => n2220);
   U3969 : INV_X1 port map( A => n13735, ZN => n2764);
   U3970 : OR2_X1 port map( A1 => n1819, A2 => n14269, ZN => n14270);
   U3971 : INV_X1 port map( A => n18517, ZN => n2954);
   U3972 : XNOR2_X1 port map( A => n13795, B => n2323, ZN => n3237);
   U3973 : INV_X1 port map( A => n3405, ZN => n3396);
   U3974 : XNOR2_X1 port map( A => n1260, B => n2035, ZN => n11653);
   U3975 : OR2_X1 port map( A1 => n11803, A2 => n19626, ZN => n3168);
   U3976 : OR2_X1 port map( A1 => n11804, A2 => n20363, ZN => n11805);
   U3977 : OR2_X1 port map( A1 => n12145, A2 => n19833, ZN => n2147);
   U3978 : INV_X1 port map( A => n13344, ZN => n12937);
   U3979 : INV_X1 port map( A => n13330, ZN => n12955);
   U3980 : AND2_X1 port map( A1 => n13971, A2 => n20380, ZN => n2563);
   U3981 : AND2_X1 port map( A1 => n14326, A2 => n14327, ZN => n14353);
   U3982 : INV_X1 port map( A => n14449, ZN => n1364);
   U3983 : OAI21_X1 port map( B1 => n19907, B2 => n14148, A => n2979, ZN => 
                           n15424);
   U3984 : INV_X1 port map( A => n240, ZN => n2891);
   U3985 : NOR2_X1 port map( A1 => n14599, A2 => n1262, ZN => n1261);
   U3986 : NAND2_X1 port map( A1 => n2439, A2 => n13951, ZN => n15153);
   U3987 : OAI21_X1 port map( B1 => n1699, B2 => n1593, A => n14023, ZN => 
                           n13951);
   U3988 : BUF_X1 port map( A => n14153, Z => n14598);
   U3989 : OR2_X1 port map( A1 => n14656, A2 => n14021, ZN => n3280);
   U3990 : NOR2_X1 port map( A1 => n241, A2 => n1593, ZN => n1740);
   U3991 : INV_X1 port map( A => n14023, ZN => n1744);
   U3992 : OR2_X1 port map( A1 => n13118, A2 => n13980, ZN => n14674);
   U3994 : AND2_X1 port map( A1 => n15256, A2 => n15828, ZN => n3722);
   U3995 : OAI21_X1 port map( B1 => n14035, B2 => n2937, A => n13164, ZN => 
                           n14038);
   U3996 : INV_X1 port map( A => n14481, ZN => n2811);
   U3997 : INV_X1 port map( A => n15905, ZN => n15008);
   U3998 : AND2_X1 port map( A1 => n2696, A2 => n2695, ZN => n2167);
   U3999 : XNOR2_X1 port map( A => n12714, B => n2947, ZN => n1755);
   U4000 : INV_X1 port map( A => n3252, ZN => n3299);
   U4001 : OR2_X1 port map( A1 => n14554, A2 => n14679, ZN => n14283);
   U4002 : NAND2_X1 port map( A1 => n14235, A2 => n14596, ZN => n15430);
   U4003 : XNOR2_X1 port map( A => n13314, B => n13315, ZN => n2748);
   U4004 : AND2_X1 port map( A1 => n20471, A2 => n14021, ZN => n1699);
   U4005 : AND2_X1 port map( A1 => n20266, A2 => n14656, ZN => n1698);
   U4006 : INV_X1 port map( A => n15906, ZN => n15078);
   U4007 : OR2_X1 port map( A1 => n14217, A2 => n3697, ZN => n3538);
   U4008 : OR2_X1 port map( A1 => n14141, A2 => n14593, ZN => n2809);
   U4010 : OAI211_X1 port map( C1 => n20262, C2 => n14167, A => n3088, B => 
                           n238, ZN => n3087);
   U4011 : OAI21_X1 port map( B1 => n14447, B2 => n14455, A => n1363, ZN => 
                           n1362);
   U4012 : OR2_X1 port map( A1 => n12911, A2 => n1724, ZN => n1723);
   U4013 : OR2_X1 port map( A1 => n13979, A2 => n14678, ZN => n2353);
   U4014 : INV_X1 port map( A => n13868, ZN => n14498);
   U4015 : OR2_X1 port map( A1 => n14265, A2 => n13981, ZN => n1573);
   U4016 : NOR2_X1 port map( A1 => n15327, A2 => n2655, ZN => n15722);
   U4017 : INV_X1 port map( A => n2655, ZN => n15863);
   U4018 : INV_X1 port map( A => n15007, ZN => n2578);
   U4019 : INV_X1 port map( A => n2723, ZN => n15910);
   U4020 : INV_X1 port map( A => n15397, ZN => n2500);
   U4021 : OAI21_X1 port map( B1 => n14186, B2 => n14185, A => n14184, ZN => 
                           n15308);
   U4022 : INV_X1 port map( A => n1288, ZN => n1286);
   U4023 : INV_X1 port map( A => n14935, ZN => n15506);
   U4024 : AND2_X1 port map( A1 => n15845, A2 => n15266, ZN => n15091);
   U4025 : INV_X1 port map( A => n19007, ZN => n1782);
   U4026 : NOR2_X1 port map( A1 => n20480, A2 => n14381, ZN => n3705);
   U4027 : AOI22_X1 port map( A1 => n15007, A2 => n15906, B1 => n15907, B2 => 
                           n15905, ZN => n15419);
   U4030 : INV_X1 port map( A => n15628, ZN => n15839);
   U4031 : INV_X1 port map( A => n15573, ZN => n1520);
   U4032 : INV_X1 port map( A => n15697, ZN => n15386);
   U4033 : INV_X1 port map( A => n15702, ZN => n15385);
   U4034 : INV_X1 port map( A => n15243, ZN => n3689);
   U4035 : AND2_X1 port map( A1 => n15767, A2 => n15657, ZN => n3690);
   U4036 : INV_X1 port map( A => n15698, ZN => n3138);
   U4037 : AND2_X1 port map( A1 => n15495, A2 => n15606, ZN => n3430);
   U4038 : INV_X1 port map( A => n15442, ZN => n15446);
   U4039 : OAI21_X1 port map( B1 => n15316, B2 => n15315, A => n2731, ZN => 
                           n1226);
   U4040 : NAND2_X1 port map( A1 => n20506, A2 => n17078, ZN => n1166);
   U4041 : NOR2_X1 port map( A1 => n14224, A2 => n14729, ZN => n2642);
   U4042 : INV_X1 port map( A => n19739, ZN => n16010);
   U4043 : OR2_X1 port map( A1 => n12664, A2 => n15767, ZN => n1383);
   U4045 : OR2_X1 port map( A1 => n13950, A2 => n14693, ZN => n2952);
   U4046 : OR2_X1 port map( A1 => n14387, A2 => n14695, ZN => n2716);
   U4047 : AND2_X1 port map( A1 => n19884, A2 => n1638, ZN => n1639);
   U4048 : AND2_X1 port map( A1 => n15574, A2 => n15365, ZN => n15045);
   U4049 : INV_X1 port map( A => n19828, ZN => n15642);
   U4050 : INV_X1 port map( A => n14119, ZN => n14123);
   U4051 : OR2_X1 port map( A1 => n14312, A2 => n14903, ZN => n14978);
   U4052 : INV_X1 port map( A => n15682, ZN => n2005);
   U4054 : INV_X1 port map( A => n15587, ZN => n15990);
   U4055 : AND2_X1 port map( A1 => n15282, A2 => n15284, ZN => n1656);
   U4056 : AOI21_X1 port map( B1 => n12876, B2 => n14339, A => n19485, ZN => 
                           n3193);
   U4058 : OR2_X1 port map( A1 => n14866, A2 => n15684, ZN => n13180);
   U4059 : OR2_X1 port map( A1 => n13868, A2 => n1089, ZN => n2276);
   U4060 : NOR2_X1 port map( A1 => n15413, A2 => n15551, ZN => n15412);
   U4061 : OR2_X1 port map( A1 => n15864, A2 => n15861, ZN => n1974);
   U4062 : NOR2_X1 port map( A1 => n13906, A2 => n3696, ZN => n3695);
   U4064 : INV_X1 port map( A => n15308, ZN => n15306);
   U4065 : INV_X1 port map( A => n15110, ZN => n2644);
   U4067 : OR2_X1 port map( A1 => n17494, A2 => n17493, ZN => n2422);
   U4068 : OR2_X1 port map( A1 => n15407, A2 => n2803, ZN => n2802);
   U4069 : INV_X1 port map( A => n642, ZN => n3209);
   U4070 : XNOR2_X1 port map( A => n17289, B => n17291, ZN => n1417);
   U4071 : OR2_X1 port map( A1 => n18927, A2 => n18928, ZN => n1068);
   U4073 : OAI21_X1 port map( B1 => n196, B2 => n16308, A => n20162, ZN => 
                           n3343);
   U4075 : XNOR2_X1 port map( A => n16045, B => n16269, ZN => n16906);
   U4077 : OR2_X1 port map( A1 => n15052, A2 => n15237, ZN => n13566);
   U4078 : XNOR2_X1 port map( A => n16330, B => n880, ZN => n3448);
   U4079 : XNOR2_X1 port map( A => n16374, B => n16507, ZN => n15726);
   U4080 : XNOR2_X1 port map( A => n14376, B => n14375, ZN => n17511);
   U4081 : OR2_X1 port map( A1 => n17149, A2 => n17956, ZN => n2662);
   U4082 : OR2_X1 port map( A1 => n18092, A2 => n20109, ZN => n17569);
   U4083 : OR3_X1 port map( A1 => n17973, A2 => n19771, A3 => n2836, ZN => 
                           n2835);
   U4084 : INV_X1 port map( A => n18130, ZN => n18126);
   U4085 : OR2_X1 port map( A1 => n19787, A2 => n18753, ZN => n18263);
   U4087 : NAND4_X1 port map( A1 => n3548, A2 => n3544, A3 => n3545, A4 => 
                           n3547, ZN => n18890);
   U4088 : OR2_X1 port map( A1 => n17812, A2 => n16959, ZN => n3547);
   U4089 : NOR2_X1 port map( A1 => n16153, A2 => n17715, ZN => n16730);
   U4092 : OR2_X1 port map( A1 => n20221, A2 => n2907, ZN => n2906);
   U4093 : OR2_X1 port map( A1 => n17891, A2 => n16261, ZN => n3216);
   U4094 : OR2_X1 port map( A1 => n17898, A2 => n17896, ZN => n1924);
   U4095 : XNOR2_X1 port map( A => n1436, B => n16509, ZN => n19363);
   U4096 : OR2_X1 port map( A1 => n18335, A2 => n18332, ZN => n2219);
   U4097 : OR2_X1 port map( A1 => n18404, A2 => n18425, ZN => n1875);
   U4098 : NOR2_X1 port map( A1 => n18414, A2 => n15529, ZN => n2018);
   U4099 : AND2_X1 port map( A1 => n2544, A2 => n2545, ZN => n2546);
   U4100 : OR2_X1 port map( A1 => n18423, A2 => n18412, ZN => n2544);
   U4101 : AOI21_X1 port map( B1 => n3045, B2 => n18436, A => n18444, ZN => 
                           n18445);
   U4102 : AND2_X1 port map( A1 => n17642, A2 => n17641, ZN => n2852);
   U4103 : AND2_X1 port map( A1 => n18500, A2 => n18485, ZN => n17639);
   U4104 : AND2_X1 port map( A1 => n18497, A2 => n18498, ZN => n1174);
   U4106 : INV_X1 port map( A => n18546, ZN => n18552);
   U4107 : INV_X1 port map( A => n17584, ZN => n17923);
   U4108 : AND2_X1 port map( A1 => n18559, A2 => n18555, ZN => n1862);
   U4109 : AND2_X1 port map( A1 => n19509, A2 => n18600, ZN => n1080);
   U4110 : OR2_X1 port map( A1 => n19757, A2 => n18600, ZN => n18603);
   U4111 : AND2_X1 port map( A1 => n3436, A2 => n3437, ZN => n1799);
   U4112 : INV_X1 port map( A => n18688, ZN => n17985);
   U4113 : INV_X1 port map( A => n18671, ZN => n17964);
   U4114 : OR2_X1 port map( A1 => n18667, A2 => n18671, ZN => n1532);
   U4115 : AND2_X1 port map( A1 => n18698, A2 => n18701, ZN => n17631);
   U4116 : OR2_X1 port map( A1 => n19766, A2 => n18834, ZN => n18814);
   U4118 : NOR2_X1 port map( A1 => n18882, A2 => n18921, ZN => n18918);
   U4121 : NOR2_X1 port map( A1 => n19151, A2 => n20508, ZN => n17807);
   U4123 : INV_X1 port map( A => n18306, ZN => n2918);
   U4124 : OAI21_X1 port map( B1 => n2918, B2 => n19165, A => n17790, ZN => 
                           n17793);
   U4125 : OR2_X1 port map( A1 => n195, A2 => n18306, ZN => n17789);
   U4126 : NOR2_X1 port map( A1 => n20460, A2 => n19168, ZN => n19171);
   U4127 : OR2_X1 port map( A1 => n17201, A2 => n16153, ZN => n2236);
   U4128 : INV_X1 port map( A => n17184, ZN => n1248);
   U4129 : OR2_X1 port map( A1 => n19241, A2 => n19242, ZN => n3338);
   U4130 : INV_X1 port map( A => n17665, ZN => n2819);
   U4131 : INV_X1 port map( A => n1205, ZN => n19274);
   U4132 : OR2_X1 port map( A1 => n20515, A2 => n18164, ZN => n2227);
   U4133 : INV_X1 port map( A => n17542, ZN => n2996);
   U4134 : OR2_X1 port map( A1 => n19404, A2 => n16306, ZN => n2965);
   U4135 : OR2_X1 port map( A1 => n19463, A2 => n20152, ZN => n1145);
   U4136 : OR2_X1 port map( A1 => n19453, A2 => n19452, ZN => n19456);
   U4137 : NOR2_X1 port map( A1 => n212, A2 => n19459, ZN => n2515);
   U4138 : INV_X1 port map( A => n17091, ZN => n2516);
   U4139 : OR2_X1 port map( A1 => n2514, A2 => n17095, ZN => n2509);
   U4140 : OR2_X1 port map( A1 => n17907, A2 => n18365, ZN => n16649);
   U4142 : NAND4_X1 port map( A1 => n1732, A2 => n18376, A3 => n1733, A4 => 
                           n1728, ZN => n1727);
   U4143 : AND2_X1 port map( A1 => n18409, A2 => n18407, ZN => n16492);
   U4145 : OR2_X1 port map( A1 => n17739, A2 => n2084, ZN => n17740);
   U4146 : OR2_X1 port map( A1 => n18583, A2 => n18596, ZN => n3411);
   U4147 : OAI211_X1 port map( C1 => n19917, C2 => n19988, A => n3028, B => 
                           n18857, ZN => n18852);
   U4148 : INV_X1 port map( A => n610, ZN => n2361);
   U4149 : INV_X1 port map( A => n17535, ZN => n2193);
   U4151 : OR2_X1 port map( A1 => n18164, A2 => n19298, ZN => n1775);
   U4153 : INV_X1 port map( A => n13918, ZN => n3516);
   U4154 : INV_X1 port map( A => n14250, ZN => n2682);
   U4155 : INV_X1 port map( A => n8212, ZN => n8209);
   U4157 : INV_X1 port map( A => n8262, ZN => n3766);
   U4158 : XNOR2_X1 port map( A => n3062, B => n13583, ZN => n14396);
   U4159 : AND2_X1 port map( A1 => n4052, A2 => n135, ZN => n956);
   U4160 : INV_X1 port map( A => n5250, ZN => n1838);
   U4161 : XNOR2_X1 port map( A => n962, B => n7252, ZN => n7801);
   U4163 : AND2_X1 port map( A1 => n5968, A2 => n5967, ZN => n957);
   U4164 : AND2_X1 port map( A1 => n11446, A2 => n11201, ZN => n958);
   U4165 : OR2_X1 port map( A1 => n19885, A2 => n17559, ZN => n959);
   U4166 : OR2_X1 port map( A1 => n16462, A2 => n17483, ZN => n960);
   U4167 : INV_X1 port map( A => n5684, ZN => n3529);
   U4168 : INV_X1 port map( A => n18600, ZN => n3693);
   U4169 : INV_X1 port map( A => n9047, ZN => n3395);
   U4170 : INV_X1 port map( A => n11244, ZN => n2861);
   U4171 : INV_X1 port map( A => n11297, ZN => n2724);
   U4172 : XOR2_X1 port map( A => n10252, B => n10249, Z => n961);
   U4173 : INV_X1 port map( A => n4013, ZN => n1537);
   U4174 : XNOR2_X1 port map( A => n10338, B => n10337, ZN => n11458);
   U4175 : INV_X1 port map( A => n14566, ZN => n2282);
   U4176 : INV_X1 port map( A => n14781, ZN => n3697);
   U4177 : XOR2_X1 port map( A => n7247, B => n7246, Z => n962);
   U4178 : XOR2_X1 port map( A => n17139, B => n17138, Z => n963);
   U4179 : XNOR2_X1 port map( A => n9631, B => n9630, ZN => n11381);
   U4181 : INV_X1 port map( A => n11990, ZN => n1213);
   U4184 : INV_X1 port map( A => n12004, ZN => n1859);
   U4185 : INV_X1 port map( A => n8179, ZN => n1850);
   U4186 : INV_X1 port map( A => n12262, ZN => n3734);
   U4187 : XNOR2_X1 port map( A => n1756, B => n1755, ZN => n14465);
   U4188 : INV_X1 port map( A => n3319, ZN => n6069);
   U4189 : INV_X1 port map( A => n15443, ZN => n1494);
   U4190 : OR2_X1 port map( A1 => n5003, A2 => n4745, ZN => n964);
   U4192 : OR2_X1 port map( A1 => n10814, A2 => n10113, ZN => n965);
   U4193 : OR2_X1 port map( A1 => n9209, A2 => n9135, ZN => n966);
   U4194 : OAI211_X1 port map( C1 => n11396, C2 => n11395, A => n1460, B => 
                           n11400, ZN => n12554);
   U4195 : OR2_X1 port map( A1 => n12282, A2 => n11721, ZN => n967);
   U4196 : INV_X1 port map( A => n11142, ZN => n1749);
   U4197 : OR2_X1 port map( A1 => n3373, A2 => n14020, ZN => n968);
   U4198 : OR3_X1 port map( A1 => n9178, A2 => n9177, A3 => n9176, ZN => n969);
   U4199 : INV_X1 port map( A => n15844, ZN => n2146);
   U4200 : OR2_X1 port map( A1 => n8309, A2 => n20057, ZN => n970);
   U4202 : INV_X1 port map( A => n4892, ZN => n4377);
   U4203 : INV_X1 port map( A => n12617, ZN => n1591);
   U4204 : AND2_X1 port map( A1 => n5968, A2 => n5971, ZN => n971);
   U4205 : XNOR2_X1 port map( A => n6437, B => n6436, ZN => n7507);
   U4206 : INV_X1 port map( A => n7750, ZN => n7912);
   U4207 : OR2_X1 port map( A1 => n9158, A2 => n8696, ZN => n972);
   U4208 : OR2_X1 port map( A1 => n4226, A2 => n4853, ZN => n973);
   U4209 : XNOR2_X1 port map( A => n9970, B => n9969, ZN => n11466);
   U4210 : INV_X1 port map( A => n5563, ZN => n2940);
   U4211 : INV_X1 port map( A => n8445, ZN => n2727);
   U4212 : NAND3_X1 port map( A1 => n17504, A2 => n19898, A3 => n19815, ZN => 
                           n975);
   U4213 : INV_X1 port map( A => n15627, ZN => n2472);
   U4215 : INV_X1 port map( A => n14584, ZN => n1351);
   U4216 : XNOR2_X1 port map( A => n12367, B => n12368, ZN => n14584);
   U4217 : OR3_X1 port map( A1 => n12016, A2 => n12262, A3 => n12264, ZN => 
                           n976);
   U4218 : INV_X1 port map( A => n5115, ZN => n1915);
   U4219 : INV_X1 port map( A => n17831, ZN => n2907);
   U4220 : INV_X1 port map( A => n12437, ZN => n1099);
   U4221 : INV_X1 port map( A => n9135, ZN => n9213);
   U4222 : INV_X1 port map( A => n14666, ZN => n2676);
   U4223 : XNOR2_X1 port map( A => n1524, B => n1523, ZN => n11158);
   U4224 : XNOR2_X1 port map( A => n13740, B => n13739, ZN => n14229);
   U4225 : XOR2_X1 port map( A => n13260, B => n17089, Z => n977);
   U4226 : INV_X1 port map( A => n5112, ZN => n2042);
   U4227 : AND2_X1 port map( A1 => n9008, A2 => n9007, ZN => n978);
   U4228 : OAI211_X1 port map( C1 => n18930, C2 => n18929, A => n1067, B => 
                           n1066, ZN => n19013);
   U4229 : INV_X1 port map( A => n19013, ZN => n2058);
   U4230 : XNOR2_X1 port map( A => n6601, B => n6600, ZN => n8211);
   U4231 : INV_X1 port map( A => n5328, ZN => n6054);
   U4232 : XNOR2_X1 port map( A => n9377, B => n9376, ZN => n10962);
   U4233 : XOR2_X1 port map( A => n13026, B => n13025, Z => n979);
   U4234 : OAI22_X1 port map( A1 => n11050, A2 => n11887, B1 => n11049, B2 => 
                           n11886, ZN => n12263);
   U4235 : XOR2_X1 port map( A => n6946, B => n2208, Z => n980);
   U4236 : AND2_X1 port map( A1 => n11659, A2 => n11829, ZN => n981);
   U4238 : OR3_X1 port map( A1 => n17891, A2 => n16261, A3 => n17890, ZN => 
                           n982);
   U4239 : XNOR2_X1 port map( A => n13575, B => n3823, ZN => n14154);
   U4240 : INV_X1 port map( A => n14154, ZN => n2926);
   U4241 : AND3_X1 port map( A1 => n4698, A2 => n5048, A3 => n4697, ZN => n983)
                           ;
   U4242 : INV_X1 port map( A => n12684, ZN => n2805);
   U4243 : AND2_X1 port map( A1 => n20513, A2 => n14601, ZN => n984);
   U4244 : INV_X1 port map( A => n14000, ZN => n14624);
   U4246 : XNOR2_X1 port map( A => n6298, B => n6297, ZN => n6312);
   U4247 : INV_X1 port map( A => n6312, ZN => n1726);
   U4248 : INV_X1 port map( A => n14535, ZN => n14664);
   U4249 : XNOR2_X1 port map( A => n13163, B => n13162, ZN => n14535);
   U4250 : AND2_X1 port map( A1 => n20261, A2 => n19985, ZN => n985);
   U4251 : OR2_X1 port map( A1 => n20451, A2 => n14724, ZN => n986);
   U4252 : XNOR2_X1 port map( A => n2046, B => n10025, ZN => n10746);
   U4253 : INV_X1 port map( A => n5941, ZN => n1835);
   U4254 : AND2_X1 port map( A1 => n6050, A2 => n6049, ZN => n987);
   U4255 : INV_X1 port map( A => n5971, ZN => n5700);
   U4256 : AND2_X1 port map( A1 => n18590, A2 => n19656, ZN => n988);
   U4257 : INV_X1 port map( A => n12658, ZN => n15659);
   U4258 : OR2_X1 port map( A1 => n5200, A2 => n5199, ZN => n989);
   U4259 : OR2_X1 port map( A1 => n11051, A2 => n11131, ZN => n990);
   U4260 : OR2_X1 port map( A1 => n11109, A2 => n11428, ZN => n991);
   U4261 : AND2_X1 port map( A1 => n19912, A2 => n5428, ZN => n992);
   U4263 : AND3_X1 port map( A1 => n18324, A2 => n18156, A3 => n2368, ZN => 
                           n993);
   U4264 : INV_X1 port map( A => n12110, ZN => n12441);
   U4265 : OR2_X2 port map( A1 => n4759, A2 => n4760, ZN => n6109);
   U4266 : AND2_X1 port map( A1 => n18522, A2 => n18512, ZN => n994);
   U4267 : OR2_X1 port map( A1 => n8241, A2 => n8100, ZN => n995);
   U4268 : AND2_X1 port map( A1 => n14447, A2 => n14448, ZN => n996);
   U4269 : AND2_X1 port map( A1 => n16128, A2 => n16129, ZN => n997);
   U4271 : INV_X1 port map( A => n15815, ZN => n3534);
   U4273 : AND2_X1 port map( A1 => n15742, A2 => n15521, ZN => n1000);
   U4274 : AND2_X1 port map( A1 => n1859, A2 => n12500, ZN => n1001);
   U4275 : INV_X1 port map( A => n3366, ZN => n2677);
   U4276 : INV_X1 port map( A => n14667, ZN => n3366);
   U4277 : OR2_X1 port map( A1 => n3055, A2 => n8194, ZN => n1002);
   U4278 : INV_X1 port map( A => n8657, ZN => n3518);
   U4279 : AND2_X1 port map( A1 => n12499, A2 => n201, ZN => n1003);
   U4280 : INV_X1 port map( A => n15607, ZN => n15606);
   U4281 : INV_X1 port map( A => n9666, ZN => n12103);
   U4282 : XOR2_X1 port map( A => n13843, B => n17544, Z => n1004);
   U4283 : OR2_X1 port map( A1 => n11639, A2 => n12214, ZN => n1005);
   U4284 : OR2_X1 port map( A1 => n7633, A2 => n20511, ZN => n1006);
   U4286 : INV_X1 port map( A => n9167, ZN => n9082);
   U4287 : AND2_X1 port map( A1 => n2928, A2 => n4057, ZN => n1007);
   U4288 : OR2_X1 port map( A1 => n11977, A2 => n250, ZN => n1008);
   U4289 : OR2_X1 port map( A1 => n12262, A2 => n3731, ZN => n1009);
   U4290 : AND2_X1 port map( A1 => n19922, A2 => n8203, ZN => n1010);
   U4291 : AND2_X1 port map( A1 => n284, A2 => n5953, ZN => n1011);
   U4292 : OR2_X1 port map( A1 => n9298, A2 => n891, ZN => n1012);
   U4293 : NAND2_X1 port map( A1 => n17097, A2 => n18111, ZN => n1013);
   U4294 : OR2_X1 port map( A1 => n13507, A2 => n14498, ZN => n1014);
   U4295 : NOR2_X2 port map( A1 => n11196, A2 => n11195, ZN => n12480);
   U4296 : INV_X1 port map( A => n12480, ZN => n2550);
   U4297 : AND2_X1 port map( A1 => n9021, A2 => n9023, ZN => n1015);
   U4298 : NAND2_X1 port map( A1 => n19033, A2 => n19992, ZN => n1016);
   U4299 : INV_X1 port map( A => n13939, ZN => n14422);
   U4300 : INV_X1 port map( A => n15822, ZN => n15507);
   U4301 : AND2_X1 port map( A1 => n19524, A2 => n4528, ZN => n1017);
   U4302 : INV_X1 port map( A => n7568, ZN => n8263);
   U4303 : OR2_X1 port map( A1 => n15674, A2 => n15673, ZN => n1018);
   U4304 : AND2_X1 port map( A1 => n14935, A2 => n15187, ZN => n1019);
   U4305 : INV_X1 port map( A => n9048, ZN => n3394);
   U4306 : INV_X1 port map( A => n9329, ZN => n2174);
   U4307 : OR2_X1 port map( A1 => n12647, A2 => n12684, ZN => n1020);
   U4308 : BUF_X1 port map( A => n15220, Z => n17479);
   U4309 : INV_X1 port map( A => n15187, ZN => n15504);
   U4310 : OR2_X1 port map( A1 => n14392, A2 => n14717, ZN => n1021);
   U4311 : OR2_X1 port map( A1 => n18072, A2 => n19753, ZN => n1022);
   U4312 : INV_X1 port map( A => n9159, ZN => n1230);
   U4313 : OR2_X1 port map( A1 => n8958, A2 => n8959, ZN => n1023);
   U4314 : OR2_X1 port map( A1 => n14266, A2 => n14265, ZN => n1024);
   U4315 : OR2_X1 port map( A1 => n6220, A2 => n5758, ZN => n1025);
   U4316 : INV_X1 port map( A => n4840, ZN => n4223);
   U4317 : INV_X1 port map( A => n19208, ZN => n2943);
   U4318 : INV_X1 port map( A => n8420, ZN => n9214);
   U4319 : AND2_X1 port map( A1 => n5300, A2 => n5428, ZN => n1026);
   U4321 : INV_X1 port map( A => n8708, ZN => n1041);
   U4322 : NAND2_X1 port map( A1 => n9082, A2 => n9166, ZN => n1027);
   U4323 : INV_X1 port map( A => n12549, ZN => n3615);
   U4324 : NAND3_X1 port map( A1 => n4841, A2 => n3978, A3 => n20105, ZN => 
                           n1028);
   U4325 : INV_X1 port map( A => n19410, ZN => n3749);
   U4327 : INV_X1 port map( A => n573, ZN => n1259);
   U4328 : INV_X1 port map( A => n2275, ZN => n2709);
   U4329 : INV_X1 port map( A => n1911, ZN => n1780);
   U4330 : INV_X1 port map( A => n18146, ZN => n1228);
   U4331 : INV_X1 port map( A => n2401, ZN => n1781);
   U4332 : INV_X1 port map( A => n18819, ZN => n1783);
   U4333 : XNOR2_X1 port map( A => n10163, B => n2329, ZN => n1031);
   U4334 : NAND2_X1 port map( A1 => n14547, A2 => n20266, ZN => n1033);
   U4336 : NAND2_X1 port map( A1 => n14656, A2 => n14021, ZN => n1034);
   U4337 : NOR2_X1 port map( A1 => n18319, A2 => n1035, ZN => n3776);
   U4339 : OAI21_X1 port map( B1 => n18317, B2 => n1035, A => n18157, ZN => 
                           n18059);
   U4341 : OAI211_X1 port map( C1 => n19174, C2 => n1035, A => n19168, B => 
                           n19169, ZN => n19173);
   U4343 : AND2_X1 port map( A1 => n1041, A2 => n1037, ZN => n3058);
   U4344 : OR2_X1 port map( A1 => n1041, A2 => n1037, ZN => n8711);
   U4345 : OAI21_X1 port map( B1 => n9233, B2 => n1037, A => n1036, ZN => n6215
                           );
   U4346 : NAND2_X1 port map( A1 => n8411, A2 => n1037, ZN => n1036);
   U4347 : OAI21_X1 port map( B1 => n11127, B2 => n1039, A => n1038, ZN => 
                           n10817);
   U4348 : NAND2_X1 port map( A1 => n11127, A2 => n1040, ZN => n1038);
   U4349 : NAND2_X1 port map( A1 => n20099, A2 => n1040, ZN => n2729);
   U4350 : NAND2_X1 port map( A1 => n1040, A2 => n19725, ZN => n11359);
   U4351 : NAND3_X1 port map( A1 => n9238, A2 => n8411, A3 => n2653, ZN => 
                           n8631);
   U4352 : AOI21_X1 port map( B1 => n9180, B2 => n9238, A => n2653, ZN => n9185
                           );
   U4353 : NOR2_X1 port map( A1 => n248, A2 => n1042, ZN => n1044);
   U4354 : NOR2_X1 port map( A1 => n11061, A2 => n12261, ZN => n1042);
   U4355 : NAND2_X1 port map( A1 => n1045, A2 => n1044, ZN => n1043);
   U4357 : NAND2_X1 port map( A1 => n248, A2 => n12262, ZN => n12565);
   U4358 : NAND2_X1 port map( A1 => n1048, A2 => n1046, ZN => n5304);
   U4359 : NAND2_X1 port map( A1 => n1047, A2 => n4457, ZN => n1046);
   U4361 : NAND2_X1 port map( A1 => n4720, A2 => n4081, ZN => n1048);
   U4362 : NAND2_X1 port map( A1 => n1049, A2 => n1163, ZN => n4720);
   U4363 : NAND2_X1 port map( A1 => n19868, A2 => n5075, ZN => n1049);
   U4364 : NAND2_X1 port map( A1 => n1472, A2 => n4667, ZN => n5255);
   U4365 : NAND3_X1 port map( A1 => n1472, A2 => n4667, A3 => n19688, ZN => 
                           n1050);
   U4366 : NAND2_X1 port map( A1 => n5257, A2 => n4668, ZN => n1051);
   U4367 : OR2_X1 port map( A1 => n12334, A2 => n11992, ZN => n11970);
   U4368 : INV_X1 port map( A => n11240, ZN => n11346);
   U4371 : INV_X1 port map( A => n11829, ZN => n1578);
   U4372 : OR2_X1 port map( A1 => n7855, A2 => n6830, ZN => n7857);
   U4373 : INV_X1 port map( A => n3959, ZN => n5580);
   U4374 : OAI21_X1 port map( B1 => n12416, B2 => n11312, A => n2758, ZN => 
                           n13031);
   U4375 : AND2_X1 port map( A1 => n4901, A2 => n4856, ZN => n3769);
   U4376 : INV_X1 port map( A => n5663, ZN => n6098);
   U4377 : OR2_X1 port map( A1 => n5663, A2 => n5953, ZN => n6099);
   U4378 : NOR2_X1 port map( A1 => n10513, A2 => n11034, ZN => n10836);
   U4379 : OR2_X1 port map( A1 => n10783, A2 => n11034, ZN => n2485);
   U4380 : INV_X1 port map( A => n11034, ZN => n11435);
   U4381 : INV_X1 port map( A => n8611, ZN => n2781);
   U4382 : OR2_X1 port map( A1 => n4197, A2 => n4755, ZN => n2034);
   U4383 : INV_X1 port map( A => n15756, ZN => n2103);
   U4384 : OR2_X1 port map( A1 => n3986, A2 => n20459, ZN => n1719);
   U4385 : AND2_X1 port map( A1 => n16810, A2 => n19655, ZN => n17927);
   U4386 : OR2_X1 port map( A1 => n19737, A2 => n19672, ZN => n17149);
   U4388 : AND2_X1 port map( A1 => n11193, A2 => n11186, ZN => n11083);
   U4389 : XNOR2_X1 port map( A => n2211, B => n6772, ZN => n7686);
   U4390 : NOR2_X1 port map( A1 => n10745, A2 => n20233, ZN => n1788);
   U4391 : INV_X1 port map( A => n8253, ZN => n6704);
   U4392 : OR2_X1 port map( A1 => n8253, A2 => n8251, ZN => n8250);
   U4393 : AND2_X1 port map( A1 => n1807, A2 => n4369, ZN => n2936);
   U4394 : INV_X1 port map( A => n1807, ZN => n1685);
   U4395 : INV_X1 port map( A => n17686, ZN => n1605);
   U4396 : INV_X1 port map( A => n14813, ZN => n14812);
   U4397 : OR2_X1 port map( A1 => n15582, A2 => n3315, ZN => n15811);
   U4398 : NOR2_X1 port map( A1 => n905, A2 => n8742, ZN => n2066);
   U4399 : OR2_X1 port map( A1 => n8482, A2 => n8743, ZN => n9370);
   U4400 : NAND2_X1 port map( A1 => n5568, A2 => n2377, ZN => n1052);
   U4401 : NAND2_X1 port map( A1 => n5568, A2 => n2377, ZN => n1053);
   U4402 : NAND2_X1 port map( A1 => n5568, A2 => n2377, ZN => n7287);
   U4403 : AND2_X1 port map( A1 => n8162, A2 => n7852, ZN => n8260);
   U4405 : AND2_X1 port map( A1 => n11158, A2 => n11160, ZN => n9555);
   U4406 : AND3_X1 port map( A1 => n14870, A2 => n14869, A3 => n14868, ZN => 
                           n1054);
   U4409 : OR2_X1 port map( A1 => n18350, A2 => n18287, ZN => n18354);
   U4410 : OR2_X1 port map( A1 => n15457, A2 => n15050, ZN => n15352);
   U4411 : MUX2_X1 port map( A => n15210, B => n15209, S => n3822, Z => n15215)
                           ;
   U4412 : NOR2_X1 port map( A1 => n15559, A2 => n3822, ZN => n15511);
   U4413 : OR2_X1 port map( A1 => n3822, A2 => n15558, ZN => n14964);
   U4414 : OR2_X1 port map( A1 => n14236, A2 => n14148, ZN => n14150);
   U4415 : INV_X1 port map( A => n11253, ZN => n10803);
   U4416 : NAND2_X1 port map( A1 => n3405, A2 => n10716, ZN => n3404);
   U4417 : OR2_X1 port map( A1 => n12003, A2 => n12001, ZN => n3240);
   U4418 : OR2_X1 port map( A1 => n3537, A2 => n12001, ZN => n2184);
   U4419 : OR2_X1 port map( A1 => n14150, A2 => n14239, ZN => n14008);
   U4420 : OR2_X1 port map( A1 => n14240, A2 => n14239, ZN => n14241);
   U4421 : NOR2_X1 port map( A1 => n9241, A2 => n9240, ZN => n1777);
   U4422 : AND2_X1 port map( A1 => n9189, A2 => n9240, ZN => n2444);
   U4423 : AND2_X1 port map( A1 => n9240, A2 => n8713, ZN => n6656);
   U4424 : OR2_X1 port map( A1 => n8569, A2 => n8568, ZN => n3227);
   U4425 : OAI21_X1 port map( B1 => n20490, B2 => n7466, A => n3680, ZN => 
                           n3679);
   U4426 : INV_X1 port map( A => n7797, ZN => n8017);
   U4427 : OR2_X1 port map( A1 => n5277, A2 => n5709, ZN => n3467);
   U4428 : AOI21_X1 port map( B1 => n5817, B2 => n5990, A => n5815, ZN => n3470
                           );
   U4429 : AND2_X1 port map( A1 => n12230, A2 => n12122, ZN => n12235);
   U4430 : INV_X1 port map( A => n12230, ZN => n12227);
   U4431 : AND2_X1 port map( A1 => n15510, A2 => n14159, ZN => n15210);
   U4432 : XNOR2_X1 port map( A => n9892, B => n9893, ZN => n3471);
   U4433 : INV_X1 port map( A => n3471, ZN => n11474);
   U4434 : NOR2_X1 port map( A1 => n11219, A2 => n3471, ZN => n11217);
   U4435 : XNOR2_X1 port map( A => n19746, B => n10425, ZN => n10340);
   U4436 : INV_X1 port map( A => n18697, ZN => n1055);
   U4437 : XNOR2_X1 port map( A => n13624, B => n641, ZN => n10793);
   U4438 : AND3_X1 port map( A1 => n8207, A2 => n8206, A3 => n2885, ZN => n1056
                           );
   U4439 : BUF_X1 port map( A => n10154, Z => n1057);
   U4440 : OR2_X1 port map( A1 => n8208, A2 => n2886, ZN => n2885);
   U4441 : OAI211_X1 port map( C1 => n9118, C2 => n9218, A => n9117, B => n9116
                           , ZN => n10154);
   U4442 : NOR2_X1 port map( A1 => n12609, A2 => n12601, ZN => n12607);
   U4444 : AOI21_X1 port map( B1 => n3898, B2 => n4005, A => n2490, ZN => n3901
                           );
   U4445 : OAI21_X1 port map( B1 => n1363, B2 => n1072, A => n1071, ZN => n1070
                           );
   U4446 : AND2_X1 port map( A1 => n11232, A2 => n10677, ZN => n1600);
   U4447 : XNOR2_X1 port map( A => n10596, B => n7663, ZN => n2202);
   U4448 : NAND2_X1 port map( A1 => n7427, A2 => n1791, ZN => n1058);
   U4449 : NAND2_X1 port map( A1 => n7426, A2 => n8232, ZN => n1059);
   U4450 : NAND2_X1 port map( A1 => n1058, A2 => n1059, ZN => n7429);
   U4451 : AND2_X1 port map( A1 => n20168, A2 => n19814, ZN => n1060);
   U4454 : INV_X1 port map( A => n5022, ZN => n4269);
   U4455 : INV_X1 port map( A => n14833, ZN => n2779);
   U4457 : OR2_X1 port map( A1 => n12100, A2 => n11381, ZN => n3325);
   U4458 : XNOR2_X1 port map( A => n6455, B => n6454, ZN => n8076);
   U4459 : INV_X1 port map( A => n14648, ZN => n3246);
   U4460 : AND2_X1 port map( A1 => n20181, A2 => n14249, ZN => n3685);
   U4461 : NOR2_X1 port map( A1 => n1960, A2 => n9106, ZN => n9104);
   U4462 : OR2_X1 port map( A1 => n4899, A2 => n4963, ZN => n3232);
   U4463 : OR2_X1 port map( A1 => n18559, A2 => n18556, ZN => n2960);
   U4464 : AND2_X1 port map( A1 => n9147, A2 => n8790, ZN => n8683);
   U4465 : OAI211_X1 port map( C1 => n5704, C2 => n19562, A => n5999, B => 
                           n2051, ZN => n5436);
   U4466 : NOR2_X1 port map( A1 => n19756, A2 => n12240, ZN => n12241);
   U4467 : NOR2_X1 port map( A1 => n20445, A2 => n18592, ZN => n18573);
   U4468 : AND2_X1 port map( A1 => n12524, A2 => n11464, ZN => n11768);
   U4470 : OAI21_X1 port map( B1 => n14597, B2 => n14598, A => n2926, ZN => 
                           n3758);
   U4471 : INV_X1 port map( A => n14396, ZN => n1527);
   U4472 : AND2_X1 port map( A1 => n14154, A2 => n14396, ZN => n13994);
   U4473 : INV_X1 port map( A => n11176, ZN => n11173);
   U4474 : OR2_X1 port map( A1 => n10657, A2 => n11176, ZN => n2231);
   U4475 : OR2_X1 port map( A1 => n11466, A2 => n11568, ZN => n10885);
   U4476 : XNOR2_X1 port map( A => n9414, B => n9854, ZN => n10321);
   U4478 : NOR2_X1 port map( A1 => n15459, A2 => n15350, ZN => n14860);
   U4479 : AND2_X1 port map( A1 => n190, A2 => n11321, ZN => n1123);
   U4480 : OR2_X1 port map( A1 => n11253, A2 => n19886, ZN => n10310);
   U4481 : XNOR2_X1 port map( A => n17377, B => n3209, ZN => n17263);
   U4482 : XNOR2_X1 port map( A => n17377, B => n3102, ZN => n16296);
   U4484 : OR2_X1 port map( A1 => n2984, A2 => n9304, ZN => n3788);
   U4485 : XNOR2_X1 port map( A => n9799, B => n9462, ZN => n10481);
   U4486 : AND2_X1 port map( A1 => n14662, A2 => n14663, ZN => n2937);
   U4487 : INV_X1 port map( A => n14663, ZN => n1552);
   U4488 : NAND2_X1 port map( A1 => n20263, A2 => n14483, ZN => n1062);
   U4489 : XOR2_X1 port map( A => n6252, B => n6251, Z => n1063);
   U4490 : XNOR2_X1 port map( A => n3744, B => n13709, ZN => n3743);
   U4491 : XNOR2_X1 port map( A => n13708, B => n13704, ZN => n3742);
   U4492 : XNOR2_X1 port map( A => n12861, B => n13020, ZN => n13708);
   U4493 : OR2_X1 port map( A1 => n11553, A2 => n9017, ZN => n10916);
   U4494 : INV_X1 port map( A => n20360, ZN => n1452);
   U4495 : OR2_X1 port map( A1 => n7519, A2 => n20359, ZN => n3089);
   U4496 : AND2_X1 port map( A1 => n9296, A2 => n9295, ZN => n8520);
   U4497 : INV_X1 port map( A => n9296, ZN => n3418);
   U4499 : NOR2_X1 port map( A1 => n17223, A2 => n3573, ZN => n16170);
   U4500 : AND2_X1 port map( A1 => n18233, A2 => n20179, ZN => n18120);
   U4501 : NOR2_X1 port map( A1 => n17545, A2 => n18233, ZN => n17973);
   U4502 : AND2_X1 port map( A1 => n18233, A2 => n18226, ZN => n2836);
   U4503 : INV_X1 port map( A => n19496, ZN => n2697);
   U4504 : AND2_X1 port map( A1 => n11292, A2 => n20235, ZN => n3587);
   U4505 : INV_X1 port map( A => n11292, ZN => n10978);
   U4506 : OR2_X1 port map( A1 => n8325, A2 => n19856, ZN => n7584);
   U4507 : INV_X1 port map( A => n3440, ZN => n3497);
   U4508 : NOR2_X1 port map( A1 => n244, A2 => n13147, ZN => n13149);
   U4509 : OR2_X1 port map( A1 => n7627, A2 => n20198, ZN => n6212);
   U4510 : AND2_X1 port map( A1 => n20198, A2 => n8192, ZN => n7878);
   U4511 : INV_X1 port map( A => n12095, ZN => n1091);
   U4512 : INV_X1 port map( A => n18311, ZN => n19324);
   U4513 : INV_X1 port map( A => n14269, ZN => n14574);
   U4514 : INV_X1 port map( A => n15167, ZN => n15378);
   U4515 : AND2_X1 port map( A1 => n13930, A2 => n12879, ZN => n14334);
   U4516 : BUF_X1 port map( A => n13930, Z => n14338);
   U4517 : XNOR2_X1 port map( A => n13341, B => n13342, ZN => n14692);
   U4519 : OR2_X1 port map( A1 => n15162, A2 => n15501, ZN => n2293);
   U4520 : OR2_X1 port map( A1 => n14434, A2 => n14487, ZN => n14433);
   U4521 : XNOR2_X1 port map( A => n13517, B => n2296, ZN => n2834);
   U4522 : OR2_X1 port map( A1 => n5405, A2 => n5408, ZN => n5146);
   U4525 : OAI211_X1 port map( C1 => n12502, C2 => n12004, A => n12500, B => 
                           n12499, ZN => n12006);
   U4527 : OR2_X1 port map( A1 => n8981, A2 => n9267, ZN => n3797);
   U4529 : INV_X1 port map( A => n17489, ZN => n3347);
   U4530 : OR2_X1 port map( A1 => n14529, A2 => n15018, ZN => n15281);
   U4531 : OR2_X1 port map( A1 => n5562, A2 => n6036, ZN => n5534);
   U4532 : INV_X1 port map( A => n12284, ZN => n13085);
   U4534 : AND2_X1 port map( A1 => n10829, A2 => n11133, ZN => n1165);
   U4535 : OR2_X1 port map( A1 => n8958, A2 => n8960, ZN => n1477);
   U4536 : AND2_X1 port map( A1 => n4816, A2 => n5073, ZN => n2022);
   U4537 : INV_X1 port map( A => n5073, ZN => n2287);
   U4539 : OR2_X1 port map( A1 => n15226, A2 => n15454, ZN => n1987);
   U4540 : OAI22_X1 port map( A1 => n19196, A2 => n19182, B1 => n19209, B2 => 
                           n19208, ZN => n19212);
   U4541 : INV_X1 port map( A => n14450, ZN => n1363);
   U4542 : AND2_X1 port map( A1 => n19986, A2 => n19859, ZN => n2316);
   U4543 : AOI21_X1 port map( B1 => n13928, B2 => n3025, A => n14448, ZN => 
                           n14756);
   U4544 : AOI21_X1 port map( B1 => n12407, B2 => n12408, A => n12754, ZN => 
                           n3012);
   U4545 : MUX2_X1 port map( A => n11595, B => n12755, S => n12754, Z => n11596
                           );
   U4546 : AND2_X1 port map( A1 => n12754, A2 => n12407, ZN => n1234);
   U4547 : NAND2_X1 port map( A1 => n1064, A2 => n5200, ZN => n3097);
   U4548 : OAI21_X1 port map( B1 => n6089, B2 => n5176, A => n4874, ZN => n1064
                           );
   U4549 : NAND2_X1 port map( A1 => n1064, A2 => n5495, ZN => n4875);
   U4550 : AOI21_X1 port map( B1 => n269, B2 => n1065, A => n9082, ZN => n9083)
                           ;
   U4551 : NAND2_X1 port map( A1 => n3227, A2 => n1065, ZN => n8403);
   U4552 : NAND2_X1 port map( A1 => n8569, A2 => n9168, ZN => n1065);
   U4553 : NOR2_X1 port map( A1 => n273, A2 => n1560, ZN => n7995);
   U4554 : AND2_X1 port map( A1 => n19001, A2 => n19013, ZN => n19023);
   U4555 : NAND3_X1 port map( A1 => n1068, A2 => n18929, A3 => n2120, ZN => 
                           n1066);
   U4556 : NAND2_X1 port map( A1 => n18928, A2 => n17749, ZN => n1067);
   U4557 : NAND2_X1 port map( A1 => n20009, A2 => n20146, ZN => n8278);
   U4558 : NAND2_X1 port map( A1 => n251, A2 => n12437, ZN => n11943);
   U4559 : NAND2_X1 port map( A1 => n20365, A2 => n18592, ZN => n17627);
   U4560 : NAND2_X1 port map( A1 => n17096, A2 => n18633, ZN => n1069);
   U4561 : NAND2_X1 port map( A1 => n14455, A2 => n14453, ZN => n1072);
   U4562 : INV_X1 port map( A => n1070, ZN => n1359);
   U4563 : NAND3_X1 port map( A1 => n13927, A2 => n14453, A3 => n14448, ZN => 
                           n1071);
   U4564 : XNOR2_X1 port map( A => n20208, B => n6514, ZN => n1073);
   U4565 : XNOR2_X1 port map( A => n6730, B => n6515, ZN => n1074);
   U4567 : NAND2_X1 port map( A1 => n1078, A2 => n15336, ZN => n1077);
   U4568 : NAND2_X1 port map( A1 => n15339, A2 => n15469, ZN => n15466);
   U4570 : INV_X1 port map( A => n15466, ZN => n1078);
   U4571 : NAND3_X1 port map( A1 => n14897, A2 => n19888, A3 => n15466, ZN => 
                           n1079);
   U4572 : NAND2_X1 port map( A1 => n1080, A2 => n18619, ZN => n18628);
   U4573 : NOR2_X1 port map( A1 => n1080, A2 => n18619, ZN => n18180);
   U4574 : XNOR2_X1 port map( A => n1081, B => n7143, ZN => n6374);
   U4575 : XNOR2_X1 port map( A => n1081, B => n6839, ZN => n6891);
   U4576 : XNOR2_X1 port map( A => n6307, B => n1081, ZN => n6309);
   U4577 : NAND2_X1 port map( A1 => n1083, A2 => n989, ZN => n1082);
   U4578 : INV_X1 port map( A => n5177, ZN => n1083);
   U4579 : NAND2_X1 port map( A1 => n1086, A2 => n1084, ZN => n9151);
   U4580 : NAND2_X1 port map( A1 => n1085, A2 => n7921, ZN => n1084);
   U4581 : MUX2_X1 port map( A => n7984, B => n7981, S => n6312, Z => n1085);
   U4582 : NAND3_X1 port map( A1 => n7920, A2 => n7768, A3 => n1087, ZN => 
                           n1086);
   U4583 : NAND2_X1 port map( A1 => n7919, A2 => n1726, ZN => n1087);
   U4584 : NAND2_X1 port map( A1 => n19812, A2 => n7978, ZN => n7920);
   U4585 : INV_X1 port map( A => n1089, ZN => n14304);
   U4586 : NAND2_X1 port map( A1 => n14506, A2 => n1089, ZN => n14502);
   U4588 : OAI21_X1 port map( B1 => n14498, B2 => n14506, A => n1089, ZN => 
                           n13974);
   U4589 : NAND2_X1 port map( A1 => n15020, A2 => n1090, ZN => n14960);
   U4590 : INV_X1 port map( A => n1656, ZN => n1090);
   U4591 : NAND2_X1 port map( A1 => n1091, A2 => n12686, ZN => n12428);
   U4592 : NOR2_X1 port map( A1 => n3649, A2 => n1094, ZN => n11944);
   U4593 : OAI21_X1 port map( B1 => n2805, B2 => n1094, A => n12428, ZN => 
                           n12434);
   U4594 : OAI21_X1 port map( B1 => n12687, B2 => n1094, A => n1092, ZN => 
                           n1550);
   U4595 : OAI211_X1 port map( C1 => n12651, C2 => n1094, A => n12650, B => 
                           n1093, ZN => n13543);
   U4596 : OAI21_X1 port map( B1 => n12646, B2 => n12685, A => n1094, ZN => 
                           n1093);
   U4597 : INV_X1 port map( A => n12095, ZN => n1094);
   U4598 : NAND2_X1 port map( A1 => n5823, A2 => n6017, ZN => n1096);
   U4599 : OAI21_X1 port map( B1 => n1098, B2 => n12442, A => n1097, ZN => 
                           n11067);
   U4600 : NAND2_X1 port map( A1 => n12442, A2 => n12443, ZN => n1097);
   U4601 : NAND2_X1 port map( A1 => n1099, A2 => n11942, ZN => n1098);
   U4602 : INV_X1 port map( A => n1101, ZN => n1100);
   U4603 : OAI22_X1 port map( A1 => n15614, A2 => n15546, B1 => n15619, B2 => 
                           n15547, ZN => n1101);
   U4604 : NAND2_X1 port map( A1 => n15071, A2 => n15615, ZN => n15614);
   U4605 : INV_X1 port map( A => n15615, ZN => n15619);
   U4606 : NAND2_X1 port map( A1 => n9071, A2 => n9346, ZN => n1102);
   U4607 : NAND2_X1 port map( A1 => n9072, A2 => n9339, ZN => n1103);
   U4608 : OAI21_X2 port map( B1 => n9243, B2 => n268, A => n2636, ZN => n9854)
                           ;
   U4609 : NAND2_X1 port map( A1 => n1486, A2 => n1104, ZN => n2717);
   U4610 : NAND3_X1 port map( A1 => n14125, A2 => n14126, A3 => n1104, ZN => 
                           n14129);
   U4611 : OR2_X1 port map( A1 => n19731, A2 => n14394, ZN => n2201);
   U4612 : AOI21_X1 port map( B1 => n1661, B2 => n214, A => n1660, ZN => n1659)
                           ;
   U4613 : OAI21_X1 port map( B1 => n15919, B2 => n15420, A => n3709, ZN => 
                           n14259);
   U4614 : NAND2_X1 port map( A1 => n1105, A2 => n8303, ZN => n1242);
   U4615 : NAND2_X1 port map( A1 => n1247, A2 => n7876, ZN => n1105);
   U4616 : NAND2_X1 port map( A1 => n1108, A2 => n1107, ZN => n1106);
   U4617 : INV_X1 port map( A => n3389, ZN => n1107);
   U4618 : NAND2_X1 port map( A1 => n3391, A2 => n3390, ZN => n1108);
   U4620 : NAND2_X1 port map( A1 => n1111, A2 => n1110, ZN => n1109);
   U4621 : AOI21_X1 port map( B1 => n17868, B2 => n17676, A => n17078, ZN => 
                           n1110);
   U4622 : NAND2_X1 port map( A1 => n17074, A2 => n1112, ZN => n1111);
   U4623 : NAND2_X1 port map( A1 => n1114, A2 => n1113, ZN => n16631);
   U4624 : NAND2_X1 port map( A1 => n16627, A2 => n16465, ZN => n1113);
   U4625 : NAND2_X1 port map( A1 => n16628, A2 => n1115, ZN => n1114);
   U4626 : NAND3_X1 port map( A1 => n9498, A2 => n11670, A3 => n11845, ZN => 
                           n1116);
   U4627 : NAND2_X1 port map( A1 => n9543, A2 => n12185, ZN => n1117);
   U4628 : XNOR2_X1 port map( A => n12286, B => n12287, ZN => n3440);
   U4629 : OAI21_X1 port map( B1 => n17911, B2 => n17912, A => n18501, ZN => 
                           n1118);
   U4630 : AOI21_X2 port map( B1 => n15924, B2 => n15923, A => n1119, ZN => 
                           n16224);
   U4631 : AND2_X1 port map( A1 => n7548, A2 => n7547, ZN => n2778);
   U4632 : INV_X1 port map( A => n14571, ZN => n14267);
   U4633 : NAND2_X1 port map( A1 => n12348, A2 => n1120, ZN => n13778);
   U4634 : NAND2_X1 port map( A1 => n1001, A2 => n12497, ZN => n1120);
   U4637 : NOR2_X1 port map( A1 => n1123, A2 => n11327, ZN => n1122);
   U4639 : NAND2_X1 port map( A1 => n11488, A2 => n12530, ZN => n11520);
   U4640 : NAND2_X1 port map( A1 => n11209, A2 => n11443, ZN => n10469);
   U4641 : NAND2_X1 port map( A1 => n4401, A2 => n4400, ZN => n6153);
   U4642 : NAND2_X1 port map( A1 => n14076, A2 => n14780, ZN => n14217);
   U4645 : OR2_X1 port map( A1 => n17812, A2 => n19846, ZN => n18949);
   U4647 : NAND2_X1 port map( A1 => n8571, A2 => n9062, ZN => n8572);
   U4648 : INV_X1 port map( A => n5845, ZN => n5847);
   U4649 : INV_X1 port map( A => n3507, ZN => n3711);
   U4650 : AND2_X1 port map( A1 => n1336, A2 => n920, ZN => n1872);
   U4651 : OAI211_X1 port map( C1 => n7227, C2 => n8313, A => n7226, B => n7225
                           , ZN => n8925);
   U4652 : INV_X1 port map( A => n9313, ZN => n9053);
   U4653 : AOI21_X1 port map( B1 => n3796, B2 => n20568, A => n2525, ZN => 
                           n2524);
   U4654 : INV_X1 port map( A => n8813, ZN => n8810);
   U4655 : AND3_X1 port map( A1 => n11094, A2 => n11443, A3 => n11445, ZN => 
                           n2656);
   U4656 : INV_X1 port map( A => n15422, ZN => n3710);
   U4657 : INV_X1 port map( A => n8602, ZN => n8956);
   U4659 : INV_X1 port map( A => n15521, ZN => n15593);
   U4660 : INV_X1 port map( A => n13041, ZN => n12697);
   U4661 : INV_X1 port map( A => n17494, ZN => n17488);
   U4662 : XNOR2_X1 port map( A => n6719, B => n6761, ZN => n7079);
   U4663 : XNOR2_X1 port map( A => n16980, B => n17109, ZN => n16892);
   U4664 : NOR2_X1 port map( A1 => n10919, A2 => n10755, ZN => n10923);
   U4666 : OR2_X1 port map( A1 => n9272, A2 => n9275, ZN => n9282);
   U4667 : XNOR2_X1 port map( A => n3162, B => n20064, ZN => n15087);
   U4668 : INV_X1 port map( A => n11769, ZN => n11792);
   U4669 : NAND2_X1 port map( A1 => n2271, A2 => n2270, ZN => n11769);
   U4670 : NAND2_X1 port map( A1 => n7694, A2 => n7911, ZN => n1679);
   U4671 : INV_X1 port map( A => n1770, ZN => n5624);
   U4674 : NAND2_X1 port map( A1 => n3429, A2 => n1126, ZN => n3428);
   U4675 : NAND2_X1 port map( A1 => n3431, A2 => n3427, ZN => n1126);
   U4678 : XNOR2_X2 port map( A => n12789, B => n12790, ZN => n14335);
   U4679 : NAND2_X1 port map( A1 => n1127, A2 => n2485, ZN => n2484);
   U4680 : NAND2_X1 port map( A1 => n11116, A2 => n11440, ZN => n1127);
   U4681 : NOR2_X1 port map( A1 => n3617, A2 => n12549, ZN => n3613);
   U4682 : NAND2_X1 port map( A1 => n1761, A2 => n1128, ZN => n1759);
   U4684 : NAND2_X1 port map( A1 => n5860, A2 => n6140, ZN => n5620);
   U4685 : OAI21_X2 port map( B1 => n4456, B2 => n153, A => n4455, ZN => n6140)
                           ;
   U4686 : NAND2_X1 port map( A1 => n15237, A2 => n15350, ZN => n15353);
   U4687 : OAI21_X2 port map( B1 => n13881, B2 => n13555, A => n13554, ZN => 
                           n15350);
   U4688 : NAND3_X2 port map( A1 => n1129, A2 => n2730, A3 => n14147, ZN => 
                           n15558);
   U4691 : NAND2_X1 port map( A1 => n12226, A2 => n12228, ZN => n11692);
   U4692 : NAND2_X1 port map( A1 => n10927, A2 => n10928, ZN => n10931);
   U4693 : NOR2_X1 port map( A1 => n11549, A2 => n11546, ZN => n10928);
   U4694 : NOR2_X1 port map( A1 => n11371, A2 => n11372, ZN => n13099);
   U4695 : XNOR2_X1 port map( A => n17005, B => n16873, ZN => n2994);
   U4697 : NOR2_X1 port map( A1 => n11834, A2 => n12359, ZN => n11835);
   U4699 : NAND2_X1 port map( A1 => n9831, A2 => n11343, ZN => n1133);
   U4700 : NAND2_X1 port map( A1 => n12631, A2 => n3401, ZN => n12632);
   U4702 : AND2_X1 port map( A1 => n5496, A2 => n5741, ZN => n2525);
   U4703 : AND2_X1 port map( A1 => n8017, A2 => n7965, ZN => n7811);
   U4704 : XNOR2_X1 port map( A => n7293, B => n7292, ZN => n7786);
   U4705 : AND2_X1 port map( A1 => n19434, A2 => n19433, ZN => n2450);
   U4706 : INV_X1 port map( A => n4021, ZN => n4131);
   U4707 : INV_X1 port map( A => n12523, ZN => n12288);
   U4708 : INV_X1 port map( A => n8890, ZN => n9005);
   U4712 : NAND2_X1 port map( A1 => n9331, A2 => n9330, ZN => n9076);
   U4713 : NAND2_X1 port map( A1 => n2924, A2 => n14394, ZN => n2923);
   U4714 : NAND2_X2 port map( A1 => n3412, A2 => n1136, ZN => n16128);
   U4715 : OR2_X1 port map( A1 => n14111, A2 => n20498, ZN => n1136);
   U4716 : NAND2_X1 port map( A1 => n2022, A2 => n5072, ZN => n1137);
   U4718 : NAND2_X1 port map( A1 => n874, A2 => n12616, ZN => n12243);
   U4720 : AOI22_X1 port map( A1 => n13865, A2 => n3516, B1 => n701, B2 => 
                           n14442, ZN => n3174);
   U4721 : NAND2_X1 port map( A1 => n11734, A2 => n1139, ZN => n11737);
   U4723 : NAND2_X1 port map( A1 => n7492, A2 => n7491, ZN => n10028);
   U4724 : NOR2_X1 port map( A1 => n17998, A2 => n1141, ZN => n18000);
   U4725 : OAI21_X1 port map( B1 => n2960, B2 => n18568, A => n2957, ZN => 
                           n1141);
   U4726 : NAND2_X1 port map( A1 => n6587, A2 => n9189, ZN => n9188);
   U4727 : NAND3_X1 port map( A1 => n1238, A2 => n1237, A3 => n1143, ZN => 
                           n1142);
   U4728 : NAND2_X1 port map( A1 => n7845, A2 => n8114, ZN => n1144);
   U4729 : NAND2_X1 port map( A1 => n13671, A2 => n14716, ZN => n14245);
   U4730 : NAND2_X1 port map( A1 => n19456, A2 => n1145, ZN => n18014);
   U4731 : NAND2_X1 port map( A1 => n16402, A2 => n16401, ZN => n1146);
   U4732 : NAND2_X1 port map( A1 => n16403, A2 => n16404, ZN => n1147);
   U4735 : XNOR2_X1 port map( A => n10370, B => n2900, ZN => n2046);
   U4738 : NAND2_X1 port map( A1 => n4848, A2 => n3996, ZN => n4849);
   U4739 : INV_X1 port map( A => n9616, ZN => n3515);
   U4740 : NAND2_X1 port map( A1 => n1858, A2 => n1861, ZN => n1149);
   U4743 : NAND2_X1 port map( A1 => n4899, A2 => n4962, ZN => n3974);
   U4744 : OR2_X1 port map( A1 => n9106, A2 => n9105, ZN => n8780);
   U4746 : OAI211_X1 port map( C1 => n19517, C2 => n8998, A => n8657, B => 
                           n3554, ZN => n3553);
   U4747 : OAI22_X1 port map( A1 => n15138, A2 => n15386, B1 => n15696, B2 => 
                           n15702, ZN => n15039);
   U4751 : NAND2_X1 port map( A1 => n5471, A2 => n6036, ZN => n5472);
   U4752 : NAND2_X1 port map( A1 => n5562, A2 => n5569, ZN => n5471);
   U4753 : XNOR2_X1 port map( A => n13588, B => n12770, ZN => n13490);
   U4754 : OR2_X1 port map( A1 => n17219, A2 => n19386, ZN => n3391);
   U4755 : XNOR2_X1 port map( A => n16225, B => n16134, ZN => n17119);
   U4756 : XNOR2_X1 port map( A => n1153, B => n13750, ZN => n13751);
   U4757 : XNOR2_X1 port map( A => n13748, B => n13749, ZN => n1153);
   U4758 : NAND2_X1 port map( A1 => n1155, A2 => n15049, ZN => n1154);
   U4759 : NAND2_X1 port map( A1 => n9190, A2 => n2443, ZN => n9700);
   U4761 : OAI21_X1 port map( B1 => n4131, B2 => n4293, A => n1156, ZN => n4135
                           );
   U4762 : NAND2_X1 port map( A1 => n4131, A2 => n4298, ZN => n1156);
   U4763 : NOR2_X1 port map( A1 => n11359, A2 => n20099, ZN => n3667);
   U4764 : NAND2_X1 port map( A1 => n19979, A2 => n5920, ZN => n6011);
   U4766 : NAND2_X1 port map( A1 => n1239, A2 => n4840, ZN => n4839);
   U4767 : NAND2_X1 port map( A1 => n11509, A2 => n20106, ZN => n10007);
   U4769 : INV_X1 port map( A => n1159, ZN => n1158);
   U4771 : NAND2_X1 port map( A1 => n7859, A2 => n8232, ZN => n1160);
   U4772 : OAI21_X1 port map( B1 => n12376, B2 => n19504, A => n12375, ZN => 
                           n2332);
   U4773 : NAND3_X1 port map( A1 => n5493, A2 => n5900, A3 => n6089, ZN => 
                           n2098);
   U4774 : OAI21_X1 port map( B1 => n1162, B2 => n1161, A => n20417, ZN => 
                           n17586);
   U4775 : NOR2_X1 port map( A1 => n19661, A2 => n19655, ZN => n1161);
   U4776 : INV_X1 port map( A => n18532, ZN => n1162);
   U4778 : NAND3_X1 port map( A1 => n8362, A2 => n8361, A3 => n8360, ZN => 
                           n2934);
   U4779 : NAND3_X1 port map( A1 => n14379, A2 => n2767, A3 => n20204, ZN => 
                           n2766);
   U4780 : NAND2_X1 port map( A1 => n14230, A2 => n14229, ZN => n14379);
   U4781 : AOI22_X2 port map( A1 => n15776, A2 => n15775, B1 => n15773, B2 => 
                           n15774, ZN => n16939);
   U4783 : INV_X1 port map( A => n12208, ZN => n12210);
   U4784 : AOI22_X1 port map( A1 => n10799, A2 => n11348, B1 => n10800, B2 => 
                           n11346, ZN => n1592);
   U4785 : OR2_X1 port map( A1 => n14228, A2 => n14229, ZN => n2304);
   U4788 : INV_X1 port map( A => n2627, ZN => n1164);
   U4789 : NAND2_X1 port map( A1 => n1680, A2 => n1165, ZN => n11134);
   U4790 : NAND2_X1 port map( A1 => n1167, A2 => n1166, ZN => n16728);
   U4791 : NAND2_X1 port map( A1 => n17677, A2 => n17074, ZN => n1167);
   U4793 : INV_X1 port map( A => n14451, ZN => n14180);
   U4794 : NOR2_X1 port map( A1 => n10639, A2 => n10932, ZN => n10737);
   U4795 : INV_X1 port map( A => n17214, ZN => n1173);
   U4796 : NAND2_X1 port map( A1 => n16466, A2 => n1395, ZN => n16662);
   U4797 : NOR2_X1 port map( A1 => n18496, A2 => n1174, ZN => n18499);
   U4798 : XNOR2_X1 port map( A => n17443, B => n16293, ZN => n14895);
   U4799 : OAI22_X2 port map( A1 => n14888, A2 => n14889, B1 => n15311, B2 => 
                           n14887, ZN => n17443);
   U4802 : AOI21_X1 port map( B1 => n9776, B2 => n10862, A => n11302, ZN => 
                           n1175);
   U4803 : NOR2_X1 port map( A1 => n996, A2 => n1362, ZN => n14459);
   U4804 : NAND2_X1 port map( A1 => n5085, A2 => n1596, ZN => n1360);
   U4805 : NAND2_X1 port map( A1 => n19980, A2 => n5917, ZN => n5588);
   U4806 : NOR2_X1 port map( A1 => n1176, A2 => n15336, ZN => n12874);
   U4807 : AND2_X1 port map( A1 => n12841, A2 => n12840, ZN => n1176);
   U4808 : NAND2_X1 port map( A1 => n7992, A2 => n8010, ZN => n7993);
   U4811 : NAND2_X1 port map( A1 => n1179, A2 => n1178, ZN => n14528);
   U4812 : NAND3_X1 port map( A1 => n14648, A2 => n14525, A3 => n14522, ZN => 
                           n1178);
   U4813 : NAND2_X1 port map( A1 => n14523, A2 => n19831, ZN => n1179);
   U4815 : NAND2_X1 port map( A1 => n15714, A2 => n15871, ZN => n1181);
   U4817 : NAND2_X1 port map( A1 => n14192, A2 => n14620, ZN => n1265);
   U4818 : OR2_X1 port map( A1 => n15813, A2 => n15581, ZN => n15816);
   U4820 : NAND3_X1 port map( A1 => n5316, A2 => n5572, A3 => n5583, ZN => 
                           n1182);
   U4821 : NAND2_X1 port map( A1 => n5605, A2 => n5714, ZN => n5243);
   U4822 : AOI21_X1 port map( B1 => n15782, B2 => n15783, A => n15686, ZN => 
                           n1183);
   U4823 : NOR2_X1 port map( A1 => n13912, A2 => n1184, ZN => n13917);
   U4824 : AND2_X1 port map( A1 => n15171, A2 => n15327, ZN => n1184);
   U4826 : INV_X1 port map( A => n12059, ZN => n2053);
   U4827 : XNOR2_X1 port map( A => n961, B => n1185, ZN => n1524);
   U4828 : INV_X1 port map( A => n8509, ZN => n1185);
   U4832 : XNOR2_X1 port map( A => n1187, B => n15225, ZN => n15250);
   U4833 : XNOR2_X1 port map( A => n16887, B => n16926, ZN => n1187);
   U4835 : NAND3_X1 port map( A1 => n1188, A2 => n15416, A3 => n15007, ZN => 
                           n14372);
   U4836 : NAND2_X1 port map( A1 => n15078, A2 => n15907, ZN => n1188);
   U4837 : NOR2_X2 port map( A1 => n3720, A2 => n11621, ZN => n13776);
   U4838 : OAI21_X1 port map( B1 => n8438, B2 => n9149, A => n1736, ZN => n1738
                           );
   U4839 : OAI21_X1 port map( B1 => n11160, B2 => n11159, A => n11161, ZN => 
                           n1903);
   U4840 : NAND2_X1 port map( A1 => n15443, A2 => n15442, ZN => n15312);
   U4841 : NAND3_X1 port map( A1 => n10801, A2 => n11060, A3 => n11057, ZN => 
                           n1189);
   U4842 : OR3_X1 port map( A1 => n19776, A2 => n5086, A3 => n20202, ZN => 
                           n4031);
   U4843 : NAND3_X1 port map( A1 => n17155, A2 => n19675, A3 => n17489, ZN => 
                           n2693);
   U4844 : AOI21_X1 port map( B1 => n12205, B2 => n12589, A => n1190, ZN => 
                           n12977);
   U4845 : AND2_X2 port map( A1 => n13862, A2 => n13863, ZN => n17288);
   U4846 : NOR2_X1 port map( A1 => n19509, A2 => n18600, ZN => n1195);
   U4847 : OAI21_X1 port map( B1 => n19509, B2 => n1192, A => n1193, ZN => 
                           n18219);
   U4848 : NAND2_X1 port map( A1 => n3693, A2 => n18215, ZN => n1192);
   U4849 : NAND2_X1 port map( A1 => n1195, A2 => n18625, ZN => n17576);
   U4851 : INV_X1 port map( A => n18215, ZN => n1194);
   U4852 : NAND2_X1 port map( A1 => n1196, A2 => n9006, ZN => n8767);
   U4853 : NAND2_X1 port map( A1 => n8890, A2 => n8895, ZN => n1196);
   U4854 : MUX2_X1 port map( A => n6182, B => n6181, S => n2865, Z => n6188);
   U4855 : MUX2_X2 port map( A => n6382, B => n6383, S => n6184, Z => n7355);
   U4856 : NAND2_X1 port map( A1 => n1198, A2 => n8372, ZN => n3490);
   U4857 : NAND2_X1 port map( A1 => n6733, A2 => n1199, ZN => n1198);
   U4858 : OR2_X1 port map( A1 => n6734, A2 => n8370, ZN => n1199);
   U4859 : NAND3_X1 port map( A1 => n20003, A2 => n15529, A3 => n18423, ZN => 
                           n16490);
   U4862 : INV_X1 port map( A => n1201, ZN => n9352);
   U4863 : INV_X1 port map( A => n9359, ZN => n9356);
   U4865 : NAND2_X1 port map( A1 => n9355, A2 => n1201, ZN => n1200);
   U4866 : OAI21_X1 port map( B1 => n1204, B2 => n9359, A => n1203, ZN => n1202
                           );
   U4867 : NAND2_X1 port map( A1 => n9358, A2 => n9359, ZN => n1203);
   U4868 : NAND2_X1 port map( A1 => n20447, A2 => n19269, ZN => n2533);
   U4869 : INV_X1 port map( A => n1206, ZN => n3558);
   U4870 : NAND2_X1 port map( A1 => n11513, A2 => n11510, ZN => n1206);
   U4871 : NAND2_X1 port map( A1 => n11575, A2 => n1206, ZN => n11512);
   U4872 : NAND2_X1 port map( A1 => n20424, A2 => n14542, ZN => n1208);
   U4873 : NAND2_X1 port map( A1 => n13982, A2 => n14542, ZN => n1209);
   U4874 : NAND2_X1 port map( A1 => n1918, A2 => n1210, ZN => n1917);
   U4875 : AOI21_X1 port map( B1 => n11397, B2 => n11297, A => n11399, ZN => 
                           n1210);
   U4876 : NAND2_X1 port map( A1 => n269, A2 => n8569, ZN => n1211);
   U4877 : AND2_X1 port map( A1 => n1212, A2 => n11990, ZN => n12340);
   U4878 : INV_X1 port map( A => n12334, ZN => n1212);
   U4880 : NOR2_X1 port map( A1 => n12337, A2 => n1213, ZN => n10315);
   U4881 : NAND2_X1 port map( A1 => n5309, A2 => n1214, ZN => n2466);
   U4882 : NOR2_X1 port map( A1 => n5144, A2 => n1214, ZN => n4052);
   U4884 : INV_X1 port map( A => n1215, ZN => n14587);
   U4885 : NAND2_X1 port map( A1 => n14811, A2 => n14593, ZN => n1215);
   U4886 : NAND2_X1 port map( A1 => n1215, A2 => n14812, ZN => n11791);
   U4887 : NAND2_X1 port map( A1 => n15271, A2 => n15274, ZN => n1218);
   U4888 : NAND3_X1 port map( A1 => n15604, A2 => n1221, A3 => n1216, ZN => 
                           n1219);
   U4889 : NAND2_X1 port map( A1 => n15271, A2 => n15601, ZN => n1216);
   U4891 : NAND2_X1 port map( A1 => n14986, A2 => n15274, ZN => n1220);
   U4892 : NAND2_X1 port map( A1 => n1217, A2 => n1220, ZN => n14987);
   U4893 : NAND2_X1 port map( A1 => n1218, A2 => n1219, ZN => n1217);
   U4894 : NAND2_X1 port map( A1 => n15270, A2 => n15600, ZN => n1221);
   U4895 : NAND2_X1 port map( A1 => n15275, A2 => n15276, ZN => n15604);
   U4896 : NAND2_X1 port map( A1 => n15035, A2 => n15034, ZN => n1223);
   U4897 : NAND2_X1 port map( A1 => n11843, A2 => n20201, ZN => n1224);
   U4899 : NOR2_X1 port map( A1 => n14620, A2 => n954, ZN => n15315);
   U4900 : INV_X1 port map( A => n14619, ZN => n15314);
   U4901 : NAND2_X1 port map( A1 => n13858, A2 => n1226, ZN => n15676);
   U4902 : XNOR2_X1 port map( A => n10563, B => n1227, ZN => n9526);
   U4903 : NAND2_X1 port map( A1 => n12083, A2 => n1229, ZN => n12085);
   U4904 : NAND2_X1 port map( A1 => n12415, A2 => n12417, ZN => n1229);
   U4905 : NAND2_X1 port map( A1 => n10637, A2 => n20279, ZN => n12415);
   U4906 : NAND2_X1 port map( A1 => n1230, A2 => n9158, ZN => n2782);
   U4907 : NAND2_X1 port map( A1 => n8247, A2 => n8253, ZN => n7562);
   U4908 : XNOR2_X2 port map( A => n6481, B => n6482, ZN => n8253);
   U4909 : NAND2_X1 port map( A1 => n291, A2 => n4410, ZN => n1232);
   U4910 : NAND2_X1 port map( A1 => n8334, A2 => n3645, ZN => n2301);
   U4911 : INV_X1 port map( A => n9123, ZN => n1233);
   U4912 : NAND2_X1 port map( A1 => n245, A2 => n1234, ZN => n3702);
   U4913 : NAND2_X1 port map( A1 => n12756, A2 => n12759, ZN => n1235);
   U4915 : NAND2_X1 port map( A1 => n8113, A2 => n8253, ZN => n1237);
   U4916 : NAND2_X1 port map( A1 => n6704, A2 => n3312, ZN => n1238);
   U4917 : INV_X1 port map( A => n4656, ZN => n1239);
   U4918 : NAND2_X1 port map( A1 => n4841, A2 => n1239, ZN => n4221);
   U4919 : NAND2_X1 port map( A1 => n19859, A2 => n985, ZN => n14831);
   U4920 : XNOR2_X1 port map( A => n12750, B => n12749, ZN => n2684);
   U4921 : NAND3_X1 port map( A1 => n1241, A2 => n1688, A3 => n246, ZN => n1240
                           );
   U4922 : NAND2_X1 port map( A1 => n10716, A2 => n12629, ZN => n1241);
   U4923 : NAND2_X1 port map( A1 => n8991, A2 => n8990, ZN => n8650);
   U4924 : NAND2_X1 port map( A1 => n1245, A2 => n20001, ZN => n1243);
   U4925 : NAND2_X1 port map( A1 => n8044, A2 => n8304, ZN => n1245);
   U4926 : INV_X1 port map( A => n8304, ZN => n8045);
   U4927 : NAND2_X1 port map( A1 => n8304, A2 => n8305, ZN => n1247);
   U4929 : NAND2_X1 port map( A1 => n1250, A2 => n1252, ZN => n1249);
   U4930 : NAND2_X1 port map( A1 => n12060, A2 => n11979, ZN => n1250);
   U4931 : INV_X1 port map( A => n4152, ZN => n4354);
   U4932 : NAND3_X1 port map( A1 => n4547, A2 => n4546, A3 => n4603, ZN => 
                           n1253);
   U4933 : NAND2_X1 port map( A1 => n2781, A2 => n9165, ZN => n1254);
   U4934 : NOR2_X1 port map( A1 => n9157, A2 => n1256, ZN => n1255);
   U4935 : NAND2_X1 port map( A1 => n9159, A2 => n9158, ZN => n1256);
   U4936 : NAND2_X1 port map( A1 => n11652, A2 => n11651, ZN => n1258);
   U4937 : XNOR2_X1 port map( A => n13790, B => n1259, ZN => n12786);
   U4938 : XNOR2_X1 port map( A => n1260, B => n13677, ZN => n12014);
   U4939 : XNOR2_X1 port map( A => n13734, B => n1260, ZN => n13486);
   U4940 : NAND2_X1 port map( A1 => n14251, A2 => n1261, ZN => n14254);
   U4943 : OAI211_X2 port map( C1 => n1264, C2 => n3329, A => n2681, B => n1263
                           , ZN => n15702);
   U4944 : NAND3_X1 port map( A1 => n1264, A2 => n20181, A3 => n19918, ZN => 
                           n1263);
   U4947 : NOR2_X1 port map( A1 => n7653, A2 => n8960, ZN => n1267);
   U4950 : NAND2_X1 port map( A1 => n2071, A2 => n4845, ZN => n1270);
   U4951 : OAI21_X1 port map( B1 => n4845, B2 => n4421, A => n1270, ZN => n4422
                           );
   U4952 : OR2_X1 port map( A1 => n1270, A2 => n4844, ZN => n5903);
   U4953 : NAND2_X1 port map( A1 => n1271, A2 => n3775, ZN => n2190);
   U4954 : NAND2_X1 port map( A1 => n1271, A2 => n1502, ZN => n1500);
   U4955 : NAND2_X1 port map( A1 => n1803, A2 => n1272, ZN => n4620);
   U4956 : OAI21_X1 port map( B1 => n4006, B2 => n4003, A => n1272, ZN => n4007
                           );
   U4957 : NAND3_X1 port map( A1 => n4308, A2 => n4307, A3 => n1272, ZN => 
                           n4309);
   U4958 : NAND2_X1 port map( A1 => n4302, A2 => n4306, ZN => n1272);
   U4959 : AND2_X2 port map( A1 => n12465, A2 => n991, ZN => n12138);
   U4960 : NAND2_X1 port map( A1 => n1273, A2 => n8046, ZN => n8050);
   U4961 : NAND3_X1 port map( A1 => n1273, A2 => n8046, A3 => n2597, ZN => 
                           n2635);
   U4962 : NAND2_X1 port map( A1 => n20001, A2 => n8303, ZN => n1273);
   U4963 : NOR2_X1 port map( A1 => n6105, A2 => n6109, ZN => n1275);
   U4964 : NOR2_X1 port map( A1 => n5957, A2 => n6105, ZN => n6111);
   U4965 : NAND2_X1 port map( A1 => n5172, A2 => n1275, ZN => n1274);
   U4966 : NAND2_X1 port map( A1 => n1276, A2 => n6155, ZN => n1347);
   U4967 : NAND2_X1 port map( A1 => n6153, A2 => n1277, ZN => n1276);
   U4968 : INV_X1 port map( A => n5349, ZN => n1277);
   U4969 : OAI21_X2 port map( B1 => n2585, B2 => n4380, A => n2584, ZN => n5349
                           );
   U4970 : NAND3_X1 port map( A1 => n12104, A2 => n11383, A3 => n20468, ZN => 
                           n1278);
   U4971 : NAND2_X1 port map( A1 => n10864, A2 => n11271, ZN => n1279);
   U4972 : NAND2_X1 port map( A1 => n1281, A2 => n10796, ZN => n11810);
   U4973 : INV_X1 port map( A => n9832, ZN => n1281);
   U4974 : INV_X1 port map( A => n10797, ZN => n1282);
   U4975 : NAND2_X1 port map( A1 => n15841, A2 => n1286, ZN => n15264);
   U4976 : MUX2_X1 port map( A => n15625, B => n15100, S => n1288, Z => n14417)
                           ;
   U4977 : NAND2_X1 port map( A1 => n2471, A2 => n1286, ZN => n15631);
   U4978 : NAND2_X1 port map( A1 => n1289, A2 => n1288, ZN => n1287);
   U4979 : NAND2_X1 port map( A1 => n15841, A2 => n1290, ZN => n1289);
   U4980 : NAND2_X1 port map( A1 => n15839, A2 => n15840, ZN => n1290);
   U4981 : NAND2_X1 port map( A1 => n15839, A2 => n15625, ZN => n15841);
   U4982 : NAND2_X1 port map( A1 => n15837, A2 => n15836, ZN => n1291);
   U4984 : NAND2_X1 port map( A1 => n3642, A2 => n14264, ZN => n1292);
   U4986 : MUX2_X1 port map( A => n15538, B => n15400, S => n15898, Z => n1293)
                           ;
   U4987 : NAND2_X1 port map( A1 => n14263, A2 => n14262, ZN => n1294);
   U4988 : NAND3_X1 port map( A1 => n1295, A2 => n14811, A3 => n14807, ZN => 
                           n14140);
   U4989 : NAND2_X1 port map( A1 => n1296, A2 => n18383, ZN => n18387);
   U4990 : OAI21_X1 port map( B1 => n1296, B2 => n18369, A => n18392, ZN => 
                           n18373);
   U4992 : NAND2_X2 port map( A1 => n1297, A2 => n1301, ZN => n13335);
   U4993 : NAND2_X1 port map( A1 => n1298, A2 => n11167, ZN => n1297);
   U4994 : NAND2_X1 port map( A1 => n12282, A2 => n12042, ZN => n1300);
   U4995 : NAND2_X1 port map( A1 => n1302, A2 => n12041, ZN => n1301);
   U4996 : OR2_X2 port map( A1 => n3017, A2 => n3016, ZN => n12041);
   U4997 : NAND2_X1 port map( A1 => n12278, A2 => n12282, ZN => n1302);
   U4999 : MUX2_X1 port map( A => n17391, B => n17392, S => n3066, Z => n17393)
                           ;
   U5000 : AOI22_X1 port map( A1 => n12514, A2 => n12513, B1 => n11995, B2 => 
                           n13275, ZN => n1305);
   U5001 : NAND2_X1 port map( A1 => n10365, A2 => n11110, ZN => n1306);
   U5002 : NAND2_X1 port map( A1 => n7912, A2 => n7910, ZN => n1308);
   U5003 : NAND2_X1 port map( A1 => n18772, A2 => n19803, ZN => n18713);
   U5004 : NAND3_X1 port map( A1 => n18277, A2 => n18276, A3 => n1309, ZN => 
                           n1310);
   U5005 : NAND3_X1 port map( A1 => n18772, A2 => n19803, A3 => n18781, ZN => 
                           n1309);
   U5006 : XNOR2_X1 port map( A => n1310, B => n18279, ZN => Ciphertext(82));
   U5007 : NAND2_X1 port map( A1 => n10980, A2 => n11290, ZN => n1311);
   U5008 : AOI21_X1 port map( B1 => n11292, B2 => n19506, A => n3588, ZN => 
                           n1312);
   U5009 : NAND3_X1 port map( A1 => n10813, A2 => n19949, A3 => n1039, ZN => 
                           n1314);
   U5010 : XNOR2_X1 port map( A => n10084, B => n10083, ZN => n10785);
   U5011 : OAI21_X1 port map( B1 => n1039, B2 => n1317, A => n1316, ZN => n1315
                           );
   U5012 : AOI21_X1 port map( B1 => n19725, B2 => n1039, A => n10813, ZN => 
                           n1316);
   U5013 : OR2_X1 port map( A1 => n11038, A2 => n19949, ZN => n1318);
   U5014 : NAND2_X1 port map( A1 => n10112, A2 => n11360, ZN => n11038);
   U5015 : NAND2_X1 port map( A1 => n1441, A2 => n1319, ZN => n5311);
   U5016 : AND2_X1 port map( A1 => n1320, A2 => n2468, ZN => n1319);
   U5017 : NAND3_X2 port map( A1 => n1501, A2 => n1503, A3 => n1321, ZN => 
                           n9462);
   U5018 : NAND2_X1 port map( A1 => n8979, A2 => n9265, ZN => n9264);
   U5020 : NAND2_X1 port map( A1 => n1325, A2 => n9214, ZN => n1322);
   U5021 : NAND2_X1 port map( A1 => n2726, A2 => n1326, ZN => n1325);
   U5022 : NAND3_X1 port map( A1 => n1332, A2 => n20496, A3 => n11384, ZN => 
                           n1327);
   U5023 : NAND2_X1 port map( A1 => n1331, A2 => n1330, ZN => n1329);
   U5024 : NAND2_X1 port map( A1 => n12101, A2 => n20468, ZN => n11384);
   U5025 : INV_X1 port map( A => n11384, ZN => n1331);
   U5026 : NAND2_X1 port map( A1 => n3601, A2 => n10684, ZN => n1332);
   U5028 : NAND2_X1 port map( A1 => n7879, A2 => n8053, ZN => n1335);
   U5030 : NAND2_X1 port map( A1 => n5797, A2 => n5796, ZN => n4182);
   U5031 : OAI21_X1 port map( B1 => n12298, B2 => n12299, A => n12274, ZN => 
                           n1336);
   U5032 : NAND3_X1 port map( A1 => n14576, A2 => n14574, A3 => n14575, ZN => 
                           n14577);
   U5033 : NAND2_X1 port map( A1 => n8070, A2 => n7420, ZN => n8208);
   U5034 : NAND2_X1 port map( A1 => n9317, A2 => n9065, ZN => n8466);
   U5037 : NAND2_X1 port map( A1 => n11572, A2 => n11573, ZN => n1338);
   U5039 : OAI22_X1 port map( A1 => n3458, A2 => n11125, B1 => n19949, B2 => 
                           n10813, ZN => n3459);
   U5041 : OAI21_X1 port map( B1 => n7671, B2 => n20252, A => n8377, ZN => 
                           n8145);
   U5042 : OR2_X1 port map( A1 => n14213, A2 => n3497, ZN => n3274);
   U5043 : NAND3_X1 port map( A1 => n16442, A2 => n16167, A3 => n17505, ZN => 
                           n2633);
   U5044 : NAND2_X1 port map( A1 => n2732, A2 => n1339, ZN => n2733);
   U5045 : AOI22_X1 port map( A1 => n12470, A2 => n12466, B1 => n12467, B2 => 
                           n12468, ZN => n1339);
   U5046 : NAND2_X1 port map( A1 => n5682, A2 => n5410, ZN => n5686);
   U5048 : NAND2_X1 port map( A1 => n4621, A2 => n20143, ZN => n4624);
   U5049 : NAND2_X1 port map( A1 => n18214, A2 => n18213, ZN => n17560);
   U5050 : NAND2_X1 port map( A1 => n2951, A2 => n2950, ZN => n18214);
   U5051 : NAND2_X1 port map( A1 => n3306, A2 => n1723, ZN => n1722);
   U5052 : NOR2_X1 port map( A1 => n9255, A2 => n8974, ZN => n8970);
   U5053 : INV_X1 port map( A => n11476, ZN => n3482);
   U5054 : NOR2_X1 port map( A1 => n15294, A2 => n14461, ZN => n15107);
   U5055 : INV_X1 port map( A => n8941, ZN => n8730);
   U5056 : OR2_X1 port map( A1 => n9320, A2 => n9836, ZN => n1855);
   U5057 : AND2_X1 port map( A1 => n6379, A2 => n5728, ZN => n5383);
   U5058 : OAI21_X1 port map( B1 => n5383, B2 => n19476, A => n5846, ZN => 
                           n1568);
   U5059 : INV_X1 port map( A => n13891, ZN => n14799);
   U5060 : INV_X1 port map( A => n1654, ZN => n11155);
   U5061 : XNOR2_X1 port map( A => n6794, B => n3590, ZN => n6684);
   U5062 : INV_X1 port map( A => n7932, ZN => n2031);
   U5063 : AOI21_X1 port map( B1 => n17080, B2 => n3114, A => n17825, ZN => 
                           n3115);
   U5064 : AOI22_X1 port map( A1 => n5433, A2 => n5432, B1 => n5996, B2 => 
                           n3627, ZN => n5437);
   U5065 : XNOR2_X1 port map( A => n2582, B => n13433, ZN => n1756);
   U5066 : NAND3_X1 port map( A1 => n5242, A2 => n3086, A3 => n5241, ZN => 
                           n5245);
   U5067 : OAI211_X2 port map( C1 => n5180, C2 => n4632, A => n5179, B => n5178
                           , ZN => n6985);
   U5068 : XNOR2_X1 port map( A => n13064, B => n19337, ZN => n13067);
   U5069 : OAI22_X1 port map( A1 => n8763, A2 => n8693, B1 => n2243, B2 => 
                           n9177, ZN => n8694);
   U5070 : OAI21_X2 port map( B1 => n8585, B2 => n9304, A => n1340, ZN => 
                           n10612);
   U5071 : NAND2_X1 port map( A1 => n2073, A2 => n2074, ZN => n1340);
   U5073 : NAND2_X1 port map( A1 => n19519, A2 => n9291, ZN => n9051);
   U5074 : AND2_X2 port map( A1 => n7896, A2 => n7895, ZN => n8649);
   U5075 : OAI21_X1 port map( B1 => n3711, B2 => n11216, A => n1341, ZN => 
                           n11477);
   U5076 : NAND2_X1 port map( A1 => n3711, A2 => n11076, ZN => n1341);
   U5077 : NAND3_X1 port map( A1 => n14937, A2 => n1344, A3 => n1343, ZN => 
                           n16045);
   U5078 : NAND2_X1 port map( A1 => n1019, A2 => n13933, ZN => n1343);
   U5079 : NAND2_X1 port map( A1 => n14936, A2 => n15506, ZN => n1344);
   U5080 : NAND2_X1 port map( A1 => n1347, A2 => n1345, ZN => n5247);
   U5081 : NAND2_X1 port map( A1 => n5246, A2 => n20405, ZN => n1345);
   U5083 : INV_X1 port map( A => n9188, ZN => n1778);
   U5084 : NAND3_X1 port map( A1 => n4222, A2 => n1028, A3 => n1348, ZN => 
                           n6022);
   U5085 : NAND2_X1 port map( A1 => n4840, A2 => n3977, ZN => n1348);
   U5086 : NAND2_X1 port map( A1 => n15257, A2 => n15256, ZN => n1349);
   U5087 : OR2_X1 port map( A1 => n11565, A2 => n11569, ZN => n2948);
   U5089 : NAND2_X1 port map( A1 => n13893, A2 => n1351, ZN => n1350);
   U5090 : NAND2_X1 port map( A1 => n14800, A2 => n14796, ZN => n13893);
   U5091 : INV_X1 port map( A => n12141, ZN => n11931);
   U5093 : NAND2_X1 port map( A1 => n12288, A2 => n11792, ZN => n1512);
   U5094 : NAND2_X1 port map( A1 => n4170, A2 => n4169, ZN => n4018);
   U5096 : NAND2_X1 port map( A1 => n2482, A2 => n1883, ZN => n1353);
   U5097 : INV_X1 port map( A => n2456, ZN => n1354);
   U5098 : NAND2_X1 port map( A1 => n19922, A2 => n7615, ZN => n2456);
   U5101 : INV_X1 port map( A => n4696, ZN => n2872);
   U5102 : NAND2_X1 port map( A1 => n4439, A2 => n4697, ZN => n4696);
   U5103 : NAND2_X1 port map( A1 => n10815, A2 => n10814, ZN => n1356);
   U5104 : NAND2_X1 port map( A1 => n10816, A2 => n19949, ZN => n1357);
   U5105 : OR2_X1 port map( A1 => n7801, A2 => n8016, ZN => n3211);
   U5106 : NAND2_X1 port map( A1 => n8079, A2 => n8219, ZN => n8077);
   U5107 : XNOR2_X2 port map( A => n6460, B => n6459, ZN => n8219);
   U5109 : NAND2_X1 port map( A1 => n4872, A2 => n4873, ZN => n5899);
   U5111 : NAND2_X1 port map( A1 => n1359, A2 => n1358, ZN => n15339);
   U5112 : OR2_X1 port map( A1 => n12873, A2 => n14448, ZN => n1358);
   U5113 : XNOR2_X2 port map( A => n5191, B => n5190, ZN => n8304);
   U5114 : OAI211_X1 port map( C1 => n12352, C2 => n12354, A => n3330, B => 
                           n12355, ZN => n12356);
   U5115 : XNOR2_X2 port map( A => n3944, B => Key(182), ZN => n4355);
   U5116 : INV_X1 port map( A => Plaintext(29), ZN => n2036);
   U5118 : NAND3_X1 port map( A1 => n8052, A2 => n8192, A3 => n8196, ZN => 
                           n1361);
   U5120 : NAND2_X1 port map( A1 => n2499, A2 => n8786, ZN => n9147);
   U5122 : OAI21_X1 port map( B1 => n11346, B2 => n11238, A => n1365, ZN => 
                           n10149);
   U5123 : NAND2_X1 port map( A1 => n11346, A2 => n11239, ZN => n1365);
   U5124 : NOR2_X1 port map( A1 => n3733, A2 => n12562, ZN => n11726);
   U5125 : OR2_X1 port map( A1 => n11990, A2 => n12334, ZN => n11667);
   U5126 : NAND2_X1 port map( A1 => n1367, A2 => n3589, ZN => n5665);
   U5127 : OAI21_X1 port map( B1 => n283, B2 => n5663, A => n5664, ZN => n1367)
                           ;
   U5128 : NAND2_X1 port map( A1 => n14660, A2 => n14659, ZN => n1368);
   U5129 : XNOR2_X1 port map( A => n6632, B => n6686, ZN => n1369);
   U5130 : XOR2_X1 port map( A => n13033, B => n13032, Z => n2240);
   U5131 : OAI21_X1 port map( B1 => n4913, B2 => n4911, A => n4477, ZN => n3871
                           );
   U5132 : AOI21_X1 port map( B1 => n14506, B2 => n14498, A => n14499, ZN => 
                           n1762);
   U5133 : NAND2_X1 port map( A1 => n1372, A2 => n1370, ZN => n11896);
   U5134 : NAND2_X1 port map( A1 => n11962, A2 => n1371, ZN => n1370);
   U5136 : NAND2_X1 port map( A1 => n1373, A2 => n180, ZN => n1372);
   U5137 : NAND2_X1 port map( A1 => n12629, A2 => n11618, ZN => n1373);
   U5138 : XNOR2_X1 port map( A => n1374, B => n18849, ZN => Ciphertext(96));
   U5140 : NAND2_X1 port map( A1 => n12283, A2 => n20215, ZN => n11580);
   U5142 : NAND2_X1 port map( A1 => n11107, A2 => n19830, ZN => n1376);
   U5144 : INV_X1 port map( A => n11431, ZN => n1378);
   U5145 : NOR2_X1 port map( A1 => n8957, A2 => n1379, ZN => n9670);
   U5146 : OAI22_X1 port map( A1 => n9370, A2 => n8602, B1 => n8951, B2 => 
                           n8950, ZN => n1379);
   U5148 : NAND2_X1 port map( A1 => n11708, A2 => n12479, ZN => n1380);
   U5149 : XNOR2_X1 port map( A => n13409, B => n13767, ZN => n11029);
   U5150 : NOR2_X2 port map( A1 => n11024, A2 => n11023, ZN => n13409);
   U5151 : NAND2_X1 port map( A1 => n1382, A2 => n1381, ZN => n5341);
   U5152 : NAND2_X1 port map( A1 => n6123, A2 => n5868, ZN => n1381);
   U5155 : NAND2_X1 port map( A1 => n1385, A2 => n1384, ZN => n19228);
   U5156 : NAND2_X1 port map( A1 => n19754, A2 => n19227, ZN => n1384);
   U5157 : NAND2_X1 port map( A1 => n20124, A2 => n19235, ZN => n1385);
   U5158 : OAI21_X2 port map( B1 => n4680, B2 => n169, A => n4679, ZN => n6166)
                           ;
   U5159 : OAI21_X1 port map( B1 => n11438, B2 => n11439, A => n11437, ZN => 
                           n11441);
   U5160 : NAND2_X1 port map( A1 => n8674, A2 => n8672, ZN => n7465);
   U5161 : NAND2_X1 port map( A1 => n8960, A2 => n8959, ZN => n8502);
   U5162 : NAND2_X1 port map( A1 => n15101, A2 => n15838, ZN => n15102);
   U5163 : NAND2_X1 port map( A1 => n4764, A2 => n19788, ZN => n5027);
   U5164 : NAND2_X1 port map( A1 => n13506, A2 => n1014, ZN => n13508);
   U5165 : NAND2_X1 port map( A1 => n12451, A2 => n12452, ZN => n12454);
   U5166 : OR2_X1 port map( A1 => n19474, A2 => n8193, ZN => n7881);
   U5168 : NAND2_X1 port map( A1 => n11143, A2 => n10957, ZN => n10702);
   U5169 : OR2_X1 port map( A1 => n11256, A2 => n11321, ZN => n10776);
   U5171 : NAND2_X2 port map( A1 => n7884, A2 => n7883, ZN => n9274);
   U5172 : OR2_X1 port map( A1 => n4440, A2 => n4439, ZN => n4795);
   U5174 : AOI22_X1 port map( A1 => n3468, A2 => n5985, B1 => n5989, B2 => 
                           n5711, ZN => n4113);
   U5175 : AOI21_X1 port map( B1 => n1388, B2 => n20472, A => n2225, ZN => 
                           n9303);
   U5176 : NOR2_X1 port map( A1 => n270, A2 => n9300, ZN => n1388);
   U5178 : NAND3_X1 port map( A1 => n3917, A2 => n3131, A3 => n4753, ZN => 
                           n1389);
   U5179 : NAND2_X1 port map( A1 => n3918, A2 => n1391, ZN => n1390);
   U5180 : NAND2_X1 port map( A1 => n2419, A2 => n9201, ZN => n2418);
   U5181 : NAND2_X1 port map( A1 => n20009, A2 => n9204, ZN => n2419);
   U5182 : NAND3_X1 port map( A1 => n5620, A2 => n6148, A3 => n6138, ZN => 
                           n5343);
   U5183 : NAND2_X1 port map( A1 => n2593, A2 => n2594, ZN => n2592);
   U5186 : NAND2_X1 port map( A1 => n1394, A2 => n6042, ZN => n1393);
   U5187 : OAI21_X1 port map( B1 => n6041, B2 => n5144, A => n2149, ZN => n1394
                           );
   U5188 : NAND2_X1 port map( A1 => n1213, A2 => n12334, ZN => n1396);
   U5189 : NAND2_X1 port map( A1 => n12335, A2 => n11990, ZN => n1397);
   U5190 : OAI21_X1 port map( B1 => n8424, B2 => n8423, A => n8781, ZN => n1398
                           );
   U5191 : OAI211_X2 port map( C1 => n8634, C2 => n8633, A => n8632, B => n8631
                           , ZN => n10359);
   U5192 : OAI21_X1 port map( B1 => n11989, B2 => n14623, A => n1399, ZN => 
                           n14849);
   U5193 : NAND2_X1 port map( A1 => n14195, A2 => n11988, ZN => n1399);
   U5194 : NAND2_X1 port map( A1 => n10995, A2 => n10946, ZN => n9560);
   U5195 : AOI21_X1 port map( B1 => n20165, B2 => n7770, A => n2976, ZN => 
                           n7772);
   U5196 : INV_X1 port map( A => n15503, ZN => n1758);
   U5197 : XNOR2_X1 port map( A => n13464, B => n2881, ZN => n2264);
   U5198 : NAND2_X1 port map( A1 => n1403, A2 => n11867, ZN => n2365);
   U5199 : XNOR2_X1 port map( A => n7289, B => n18170, ZN => n6932);
   U5201 : NAND2_X1 port map( A1 => n8602, A2 => n8482, ZN => n9372);
   U5202 : NAND2_X1 port map( A1 => n1405, A2 => n8093, ZN => n1404);
   U5203 : NAND2_X1 port map( A1 => n1407, A2 => n1406, ZN => n10470);
   U5204 : NAND2_X1 port map( A1 => n10468, A2 => n11201, ZN => n1406);
   U5205 : NAND2_X1 port map( A1 => n10469, A2 => n11093, ZN => n1407);
   U5206 : NAND2_X1 port map( A1 => n9931, A2 => n11523, ZN => n9932);
   U5207 : NAND2_X1 port map( A1 => n19270, A2 => n19271, ZN => n19272);
   U5209 : NAND2_X1 port map( A1 => n9328, A2 => n9330, ZN => n1408);
   U5211 : XNOR2_X1 port map( A => n10610, B => n10609, ZN => n10730);
   U5212 : OR2_X1 port map( A1 => n2527, A2 => n16306, ZN => n17648);
   U5213 : NOR2_X1 port map( A1 => n20000, A2 => n9105, ZN => n8423);
   U5214 : MUX2_X1 port map( A => n14525, B => n951, S => n14648, Z => n14310);
   U5216 : INV_X1 port map( A => n5046, ZN => n4796);
   U5217 : INV_X1 port map( A => n1508, ZN => n12130);
   U5218 : INV_X1 port map( A => n2005, ZN => n1491);
   U5219 : NOR2_X1 port map( A1 => n10911, A2 => n12606, ZN => n3764);
   U5220 : AOI22_X1 port map( A1 => n14944, A2 => n2645, B1 => n15107, B2 => 
                           n2644, ZN => n2643);
   U5221 : NAND2_X1 port map( A1 => n7618, A2 => n7420, ZN => n1411);
   U5223 : NAND3_X1 port map( A1 => n3404, A2 => n1414, A3 => n1413, ZN => 
                           n12284);
   U5224 : NAND2_X1 port map( A1 => n20184, A2 => n3402, ZN => n1413);
   U5225 : NAND2_X1 port map( A1 => n14509, A2 => n14644, ZN => n14508);
   U5226 : NAND2_X1 port map( A1 => n1415, A2 => n14354, ZN => n15909);
   U5227 : NAND2_X1 port map( A1 => n1572, A2 => n1571, ZN => n1415);
   U5229 : NOR2_X1 port map( A1 => n8315, A2 => n7475, ZN => n7594);
   U5230 : AOI21_X1 port map( B1 => n4543, B2 => n4544, A => n4542, ZN => n5538
                           );
   U5232 : NAND3_X1 port map( A1 => n8033, A2 => n20012, A3 => n8034, ZN => 
                           n1416);
   U5233 : NAND3_X2 port map( A1 => n2121, A2 => n11720, A3 => n967, ZN => 
                           n13491);
   U5234 : OR2_X1 port map( A1 => n11073, A2 => n10898, ZN => n1418);
   U5236 : NAND2_X1 port map( A1 => n2143, A2 => n11804, ZN => n1419);
   U5237 : OR2_X1 port map( A1 => n8200, A2 => n5762, ZN => n7872);
   U5238 : INV_X1 port map( A => n5102, ZN => n1421);
   U5239 : NAND2_X1 port map( A1 => n10923, A2 => n11523, ZN => n12222);
   U5240 : INV_X1 port map( A => n13017, ZN => n13576);
   U5241 : INV_X1 port map( A => n1640, ZN => n15395);
   U5243 : NAND2_X1 port map( A1 => n1423, A2 => n4413, ZN => n4414);
   U5244 : NAND2_X1 port map( A1 => n4412, A2 => n4411, ZN => n1423);
   U5245 : NAND2_X1 port map( A1 => n8324, A2 => n19856, ZN => n1424);
   U5246 : INV_X1 port map( A => n7786, ZN => n1425);
   U5247 : OR2_X1 port map( A1 => n12383, A2 => n12468, ZN => n3783);
   U5248 : OR2_X1 port map( A1 => n2628, A2 => n13891, ZN => n14797);
   U5249 : NAND2_X1 port map( A1 => n8619, A2 => n2243, ZN => n2242);
   U5250 : AND2_X1 port map( A1 => n2523, A2 => n12759, ZN => n12411);
   U5251 : NAND2_X1 port map( A1 => n1426, A2 => n6104, ZN => n5956);
   U5252 : OAI22_X1 port map( A1 => n5957, A2 => n6107, B1 => n6113, B2 => 
                           n6105, ZN => n1426);
   U5253 : OR2_X1 port map( A1 => n8650, A2 => n8649, ZN => n9281);
   U5254 : AOI22_X1 port map( A1 => n8252, A2 => n8251, B1 => n8253, B2 => 
                           n8254, ZN => n8255);
   U5256 : XNOR2_X1 port map( A => n1427, B => n12896, ZN => n12898);
   U5257 : XNOR2_X1 port map( A => n12897, B => n13126, ZN => n1427);
   U5259 : AND3_X1 port map( A1 => n14988, A2 => n14990, A3 => n14989, ZN => 
                           n14991);
   U5260 : OAI21_X1 port map( B1 => n12631, B2 => n12630, A => n11619, ZN => 
                           n11960);
   U5261 : INV_X1 port map( A => n15059, ZN => n15061);
   U5262 : XNOR2_X1 port map( A => n2285, B => n8508, ZN => n10755);
   U5263 : OAI21_X1 port map( B1 => n19657, B2 => n3522, A => n19819, ZN => 
                           n3253);
   U5265 : INV_X1 port map( A => n4233, ZN => n4860);
   U5266 : XNOR2_X1 port map( A => n10151, B => n10002, ZN => n9261);
   U5267 : INV_X1 port map( A => n1746, ZN => n6186);
   U5268 : INV_X1 port map( A => n1776, ZN => n2407);
   U5269 : INV_X1 port map( A => n15683, ZN => n15782);
   U5270 : INV_X1 port map( A => n12162, ZN => n12535);
   U5271 : NAND3_X1 port map( A1 => n19520, A2 => n7592, A3 => n8313, ZN => 
                           n7597);
   U5272 : INV_X1 port map( A => n15266, ZN => n15847);
   U5273 : INV_X1 port map( A => n8937, ZN => n8940);
   U5274 : OAI21_X1 port map( B1 => n19505, B2 => n19719, A => n11490, ZN => 
                           n2134);
   U5275 : XNOR2_X1 port map( A => n7303, B => n3067, ZN => n7310);
   U5276 : INV_X1 port map( A => n1603, ZN => n1428);
   U5277 : NAND2_X1 port map( A1 => n1430, A2 => n1429, ZN => n8724);
   U5278 : NAND3_X1 port map( A1 => n9358, A2 => n9359, A3 => n9528, ZN => 
                           n1429);
   U5279 : NAND2_X1 port map( A1 => n8723, A2 => n9356, ZN => n1430);
   U5280 : XNOR2_X1 port map( A => n6867, B => n6977, ZN => n7353);
   U5281 : NOR2_X2 port map( A1 => n8065, A2 => n1431, ZN => n9065);
   U5282 : NAND2_X1 port map( A1 => n1433, A2 => n1432, ZN => n1431);
   U5283 : NAND2_X1 port map( A1 => n8063, A2 => n8190, ZN => n1432);
   U5286 : AOI21_X1 port map( B1 => n4584, B2 => n4582, A => n4271, ZN => n2334
                           );
   U5287 : NAND2_X1 port map( A1 => n4269, A2 => n4095, ZN => n4584);
   U5289 : OAI21_X1 port map( B1 => n11145, B2 => n10642, A => n1749, ZN => 
                           n1670);
   U5290 : NAND2_X1 port map( A1 => n5698, A2 => n5973, ZN => n1435);
   U5291 : XNOR2_X1 port map( A => n17267, B => n16508, ZN => n1436);
   U5294 : NAND2_X1 port map( A1 => n7724, A2 => n8159, ZN => n8258);
   U5296 : NAND2_X1 port map( A1 => n12522, A2 => n182, ZN => n1439);
   U5297 : NAND2_X1 port map( A1 => n17665, A2 => n17662, ZN => n17086);
   U5298 : NAND3_X1 port map( A1 => n4360, A2 => n4359, A3 => n2370, ZN => 
                           n5483);
   U5299 : NOR2_X1 port map( A1 => n4363, A2 => n5719, ZN => n5240);
   U5301 : NOR2_X1 port map( A1 => n1442, A2 => n4033, ZN => n1441);
   U5303 : NAND2_X1 port map( A1 => n15438, A2 => n15775, ZN => n1444);
   U5305 : NAND2_X1 port map( A1 => n4896, A2 => n4897, ZN => n1445);
   U5306 : OAI22_X2 port map( A1 => n6047, A2 => n5313, B1 => n5312, B2 => 
                           n5781, ZN => n6728);
   U5307 : NAND2_X1 port map( A1 => n10889, A2 => n10926, ZN => n1446);
   U5308 : NAND2_X1 port map( A1 => n10844, A2 => n193, ZN => n1447);
   U5309 : NAND2_X1 port map( A1 => n1448, A2 => n709, ZN => n1485);
   U5310 : NOR2_X1 port map( A1 => n1449, A2 => n9103, ZN => n1448);
   U5311 : NAND2_X1 port map( A1 => n9100, A2 => n9099, ZN => n1449);
   U5312 : NOR2_X1 port map( A1 => n20007, A2 => n3430, ZN => n3429);
   U5314 : INV_X1 port map( A => n8917, ZN => n8734);
   U5315 : INV_X1 port map( A => n4337, ZN => n3753);
   U5316 : OR2_X1 port map( A1 => n3753, A2 => n1017, ZN => n3607);
   U5317 : NOR2_X1 port map( A1 => n14790, A2 => n14103, ZN => n2411);
   U5319 : NAND2_X1 port map( A1 => n17944, A2 => n19105, ZN => n1450);
   U5321 : NOR2_X2 port map( A1 => n14107, A2 => n14108, ZN => n16429);
   U5322 : NOR2_X1 port map( A1 => n11534, A2 => n19915, ZN => n11536);
   U5325 : NAND2_X1 port map( A1 => n9204, A2 => n9201, ZN => n8433);
   U5327 : NAND2_X1 port map( A1 => n14237, A2 => n14406, ZN => n14242);
   U5328 : NAND2_X1 port map( A1 => n12531, A2 => n924, ZN => n12530);
   U5330 : NAND2_X1 port map( A1 => n2048, A2 => n5997, ZN => n1455);
   U5331 : NAND2_X1 port map( A1 => n1457, A2 => n1456, ZN => n13568);
   U5332 : NAND2_X1 port map( A1 => n14860, A2 => n15237, ZN => n1456);
   U5333 : NAND2_X1 port map( A1 => n13561, A2 => n1458, ZN => n1457);
   U5334 : NAND2_X1 port map( A1 => n12154, A2 => n12152, ZN => n11711);
   U5335 : NAND2_X1 port map( A1 => n11169, A2 => n11170, ZN => n1459);
   U5336 : NAND2_X1 port map( A1 => n8840, A2 => n1461, ZN => n10422);
   U5337 : NAND3_X1 port map( A1 => n1631, A2 => n1630, A3 => n8676, ZN => 
                           n1461);
   U5338 : OAI21_X1 port map( B1 => n10667, B2 => n11399, A => n2044, ZN => 
                           n2043);
   U5339 : NAND3_X1 port map( A1 => n14430, A2 => n3154, A3 => n14494, ZN => 
                           n2138);
   U5340 : NAND2_X1 port map( A1 => n1462, A2 => n8205, ZN => n7874);
   U5341 : NAND2_X1 port map( A1 => n2378, A2 => n2379, ZN => n1462);
   U5342 : NAND2_X1 port map( A1 => n17891, A2 => n17890, ZN => n17662);
   U5343 : XNOR2_X2 port map( A => n16109, B => n16108, ZN => n17890);
   U5344 : INV_X1 port map( A => n12211, ZN => n2712);
   U5345 : NAND2_X1 port map( A1 => n1464, A2 => n1463, ZN => n9583);
   U5346 : NAND2_X1 port map( A1 => n9287, A2 => n9576, ZN => n1463);
   U5347 : NAND2_X1 port map( A1 => n9288, A2 => n9289, ZN => n1464);
   U5349 : INV_X1 port map( A => n1506, ZN => n3182);
   U5350 : NAND2_X1 port map( A1 => n8356, A2 => n1506, ZN => n1480);
   U5351 : NAND2_X1 port map( A1 => n3181, A2 => n7500, ZN => n1506);
   U5353 : NAND2_X1 port map( A1 => n9104, A2 => n8781, ZN => n9109);
   U5354 : NAND2_X1 port map( A1 => n1465, A2 => n4691, ZN => n4688);
   U5355 : NAND2_X1 port map( A1 => n1468, A2 => n1466, ZN => n2396);
   U5357 : NAND2_X1 port map( A1 => n1820, A2 => n14738, ZN => n1469);
   U5358 : NAND2_X1 port map( A1 => n1470, A2 => n8478, ZN => n10497);
   U5363 : XNOR2_X2 port map( A => Key(35), B => Plaintext(35), ZN => n4954);
   U5366 : OR2_X1 port map( A1 => n12579, A2 => n12576, ZN => n11924);
   U5367 : XNOR2_X1 port map( A => n7325, B => n2571, ZN => n6881);
   U5368 : INV_X1 port map( A => n4524, ZN => n4516);
   U5369 : INV_X1 port map( A => n8195, ZN => n8054);
   U5370 : INV_X1 port map( A => n2749, ZN => n2504);
   U5371 : NAND2_X1 port map( A1 => n4426, A2 => n4827, ZN => n1472);
   U5372 : OAI21_X1 port map( B1 => n1039, B2 => n1317, A => n1473, ZN => 
                           n11362);
   U5373 : NOR2_X1 port map( A1 => n11127, A2 => n19949, ZN => n1473);
   U5374 : INV_X1 port map( A => n1475, ZN => n1474);
   U5375 : OAI21_X1 port map( B1 => n5748, B2 => n2482, A => n5205, ZN => n1475
                           );
   U5376 : NAND2_X1 port map( A1 => n15295, A2 => n15297, ZN => n14770);
   U5378 : OAI22_X1 port map( A1 => n1806, A2 => n5730, B1 => n5847, B2 => 
                           n1805, ZN => n1476);
   U5379 : NAND2_X1 port map( A1 => n2461, A2 => n5098, ZN => n4712);
   U5380 : NAND2_X1 port map( A1 => n8722, A2 => n9359, ZN => n8721);
   U5381 : NAND2_X2 port map( A1 => n3490, A2 => n7672, ZN => n9359);
   U5382 : XNOR2_X1 port map( A => n6728, B => n456, ZN => n6729);
   U5383 : NAND2_X1 port map( A1 => n207, A2 => n8958, ZN => n1478);
   U5384 : INV_X1 port map( A => n12137, ZN => n12385);
   U5385 : NAND3_X1 port map( A1 => n12468, A2 => n12386, A3 => n12137, ZN => 
                           n1946);
   U5386 : XNOR2_X1 port map( A => n6960, B => n980, ZN => n6227);
   U5387 : XNOR2_X1 port map( A => n7348, B => n6226, ZN => n6960);
   U5388 : XNOR2_X1 port map( A => n9773, B => n9774, ZN => n1479);
   U5389 : INV_X1 port map( A => n6109, ZN => n5657);
   U5390 : NAND2_X1 port map( A1 => n1899, A2 => n1901, ZN => n14847);
   U5391 : NAND2_X1 port map( A1 => n11094, A2 => n11443, ZN => n11448);
   U5393 : NAND2_X1 port map( A1 => n14275, A2 => n20498, ZN => n13957);
   U5394 : NAND2_X1 port map( A1 => n8093, A2 => n8212, ZN => n7432);
   U5395 : NAND2_X1 port map( A1 => n4186, A2 => n4185, ZN => n3622);
   U5396 : NAND2_X1 port map( A1 => n4156, A2 => n3623, ZN => n4186);
   U5397 : NAND2_X1 port map( A1 => n1480, A2 => n1565, ZN => n2930);
   U5398 : OR2_X1 port map( A1 => n9251, A2 => n8974, ZN => n1481);
   U5399 : NOR2_X1 port map( A1 => n3403, A2 => n180, ZN => n3402);
   U5400 : OAI21_X1 port map( B1 => n11578, B2 => n11739, A => n11577, ZN => 
                           n2367);
   U5402 : NAND3_X2 port map( A1 => n1854, A2 => n11274, A3 => n974, ZN => 
                           n12807);
   U5403 : OAI211_X1 port map( C1 => n9004, C2 => n8890, A => n19490, B => 
                           n1484, ZN => n8626);
   U5404 : NAND2_X1 port map( A1 => n12545, A2 => n12542, ZN => n12306);
   U5405 : INV_X1 port map( A => n13989, ZN => n15302);
   U5406 : NAND2_X1 port map( A1 => n15714, A2 => n15874, ZN => n13989);
   U5407 : OAI21_X1 port map( B1 => n19515, B2 => n20000, A => n1485, ZN => 
                           n9110);
   U5409 : OAI21_X1 port map( B1 => n14688, B2 => n14690, A => n14385, ZN => 
                           n1486);
   U5410 : AOI21_X1 port map( B1 => n9028, B2 => n8829, A => n9029, ZN => n1487
                           );
   U5411 : NAND3_X1 port map( A1 => n885, A2 => n9274, A3 => n9275, ZN => n9280
                           );
   U5412 : XNOR2_X2 port map( A => Key(21), B => Plaintext(21), ZN => n4297);
   U5413 : XOR2_X1 port map( A => n13550, B => n13080, Z => n1809);
   U5414 : OAI211_X2 port map( C1 => n9069, C2 => n545, A => n2502, B => n2503,
                           ZN => n10220);
   U5415 : NAND2_X1 port map( A1 => n18427, A2 => n15529, ZN => n1701);
   U5416 : AND3_X2 port map( A1 => n2643, A2 => n2646, A3 => n3308, ZN => 
                           n17269);
   U5417 : OAI21_X1 port map( B1 => n17483, B2 => n19823, A => n1488, ZN => 
                           n15177);
   U5418 : NAND2_X1 port map( A1 => n1718, A2 => n17243, ZN => n1488);
   U5419 : NOR2_X1 port map( A1 => n15239, A2 => n3348, ZN => n1489);
   U5420 : INV_X1 port map( A => n9563, ZN => n9340);
   U5421 : NAND3_X1 port map( A1 => n1493, A2 => n1492, A3 => n1491, ZN => 
                           n1490);
   U5422 : NAND2_X1 port map( A1 => n15443, A2 => n15228, ZN => n1492);
   U5423 : NAND2_X1 port map( A1 => n15446, A2 => n1494, ZN => n1493);
   U5424 : NAND2_X1 port map( A1 => n1495, A2 => n9023, ZN => n2025);
   U5425 : OAI22_X1 port map( A1 => n8515, A2 => n9021, B1 => n8841, B2 => 
                           n8672, ZN => n1495);
   U5426 : AND3_X2 port map( A1 => n17567, A2 => n1496, A3 => n17561, ZN => 
                           n18600);
   U5427 : NAND2_X1 port map( A1 => n17563, A2 => n17562, ZN => n1496);
   U5428 : NAND2_X1 port map( A1 => n9411, A2 => n19817, ZN => n1497);
   U5430 : NAND3_X2 port map( A1 => n1500, A2 => n3771, A3 => n1499, ZN => 
                           n8979);
   U5431 : NAND2_X1 port map( A1 => n8771, A2 => n8979, ZN => n1501);
   U5432 : INV_X1 port map( A => n3775, ZN => n1502);
   U5433 : NAND2_X1 port map( A1 => n1504, A2 => n19880, ZN => n1503);
   U5434 : NAND2_X1 port map( A1 => n1505, A2 => n9266, ZN => n1504);
   U5435 : NAND2_X1 port map( A1 => n7866, A2 => n9262, ZN => n1505);
   U5436 : NAND2_X1 port map( A1 => n7742, A2 => n1506, ZN => n7698);
   U5440 : NAND2_X1 port map( A1 => n1507, A2 => n8126, ZN => n6439);
   U5441 : NOR2_X1 port map( A1 => n1507, A2 => n8470, ZN => n9087);
   U5442 : NOR2_X1 port map( A1 => n8565, A2 => n1507, ZN => n1575);
   U5443 : NAND3_X1 port map( A1 => n9091, A2 => n1507, A3 => n8884, ZN => 
                           n8887);
   U5444 : NAND2_X1 port map( A1 => n9090, A2 => n1507, ZN => n1577);
   U5445 : MUX2_X1 port map( A => n1507, B => n8565, S => n9091, Z => n8130);
   U5446 : NAND3_X1 port map( A1 => n8471, A2 => n1507, A3 => n8470, ZN => 
                           n8472);
   U5448 : OR2_X1 port map( A1 => n11586, A2 => n1508, ZN => n1547);
   U5449 : AND2_X1 port map( A1 => n12127, A2 => n1508, ZN => n1643);
   U5450 : NAND2_X1 port map( A1 => n10967, A2 => n1508, ZN => n10974);
   U5451 : OAI21_X1 port map( B1 => n11763, B2 => n12126, A => n1508, ZN => 
                           n11587);
   U5452 : AOI21_X1 port map( B1 => n10972, B2 => n1508, A => n1735, ZN => 
                           n10973);
   U5453 : NAND3_X1 port map( A1 => n1512, A2 => n1511, A3 => n1510, ZN => 
                           n1509);
   U5454 : NAND2_X1 port map( A1 => n12520, A2 => n12523, ZN => n1510);
   U5455 : NAND2_X1 port map( A1 => n11793, A2 => n12523, ZN => n1514);
   U5456 : OAI21_X1 port map( B1 => n9220, B2 => n1516, A => n1515, ZN => n2452
                           );
   U5457 : INV_X1 port map( A => n9218, ZN => n1515);
   U5458 : NOR2_X1 port map( A1 => n8797, A2 => n9113, ZN => n1516);
   U5459 : NOR2_X1 port map( A1 => n9112, A2 => n9114, ZN => n9220);
   U5460 : NAND2_X1 port map( A1 => n1517, A2 => n15364, ZN => n15367);
   U5461 : NAND2_X1 port map( A1 => n1520, A2 => n15577, ZN => n1517);
   U5462 : NAND2_X1 port map( A1 => n14643, A2 => n20473, ZN => n1518);
   U5463 : NAND2_X1 port map( A1 => n14646, A2 => n14645, ZN => n1519);
   U5464 : NAND2_X1 port map( A1 => n251, A2 => n12443, ZN => n1521);
   U5465 : OAI211_X1 port map( C1 => n12109, C2 => n1522, A => n1521, B => 
                           n12441, ZN => n12112);
   U5466 : INV_X1 port map( A => n12442, ZN => n1522);
   U5467 : OR2_X2 port map( A1 => n10682, A2 => n10681, ZN => n12442);
   U5468 : NAND2_X1 port map( A1 => n12441, A2 => n12442, ZN => n12444);
   U5469 : NAND2_X1 port map( A1 => n12438, A2 => n1522, ZN => n12113);
   U5470 : AOI22_X1 port map( A1 => n12438, A2 => n12437, B1 => n1522, B2 => 
                           n12436, ZN => n12447);
   U5471 : NAND2_X1 port map( A1 => n15711, A2 => n15871, ZN => n1525);
   U5475 : NOR2_X1 port map( A1 => n14154, A2 => n20171, ZN => n13996);
   U5476 : AND2_X1 port map( A1 => n1527, A2 => n14394, ZN => n14397);
   U5477 : NOR2_X1 port map( A1 => n5630, A2 => n5631, ZN => n1949);
   U5478 : OAI21_X2 port map( B1 => n4330, B2 => n4331, A => n4329, ZN => n5631
                           );
   U5479 : XNOR2_X1 port map( A => n17296, B => n17302, ZN => n1529);
   U5480 : XNOR2_X2 port map( A => n1530, B => Plaintext(191), ZN => n4615);
   U5481 : INV_X1 port map( A => Key(191), ZN => n1530);
   U5482 : NAND2_X1 port map( A1 => n1531, A2 => n18688, ZN => n17988);
   U5483 : NAND2_X1 port map( A1 => n17972, A2 => n1532, ZN => n1531);
   U5484 : INV_X1 port map( A => n18667, ZN => n18686);
   U5485 : NAND2_X1 port map( A1 => n5393, A2 => n5322, ZN => n5397);
   U5486 : NAND2_X1 port map( A1 => n1536, A2 => n4614, ZN => n1533);
   U5487 : NAND2_X1 port map( A1 => n1538, A2 => n7746, ZN => n2497);
   U5488 : NAND2_X1 port map( A1 => n1540, A2 => n1539, ZN => n1538);
   U5489 : NAND2_X1 port map( A1 => n7749, A2 => n7750, ZN => n1539);
   U5490 : INV_X1 port map( A => n7691, ZN => n1541);
   U5491 : NAND2_X1 port map( A1 => n9150, A2 => n9149, ZN => n1543);
   U5492 : OAI21_X1 port map( B1 => n8338, B2 => n2499, A => n9145, ZN => n1544
                           );
   U5493 : INV_X1 port map( A => n7507, ZN => n3445);
   U5495 : NAND3_X1 port map( A1 => n1549, A2 => n7912, A3 => n1548, ZN => 
                           n7913);
   U5496 : NAND2_X1 port map( A1 => n7910, A2 => n3445, ZN => n1549);
   U5500 : NOR2_X1 port map( A1 => n1552, A2 => n14666, ZN => n14669);
   U5501 : OAI21_X1 port map( B1 => n2676, B2 => n1552, A => n1551, ZN => n2675
                           );
   U5502 : NAND2_X1 port map( A1 => n1552, A2 => n14662, ZN => n1551);
   U5503 : AOI21_X1 port map( B1 => n14536, B2 => n13164, A => n1552, ZN => 
                           n14537);
   U5504 : NAND2_X1 port map( A1 => n15563, A2 => n3822, ZN => n1553);
   U5505 : NAND2_X1 port map( A1 => n15211, A2 => n15562, ZN => n1554);
   U5506 : NAND2_X1 port map( A1 => n921, A2 => n15510, ZN => n15211);
   U5507 : NAND2_X1 port map( A1 => n1555, A2 => n15866, ZN => n15859);
   U5508 : OAI21_X1 port map( B1 => n1555, B2 => n15866, A => n2655, ZN => 
                           n15172);
   U5509 : INV_X1 port map( A => n15857, ZN => n1555);
   U5510 : OR2_X1 port map( A1 => n16787, A2 => n16025, ZN => n1556);
   U5511 : NAND2_X1 port map( A1 => n1558, A2 => n16786, ZN => n1557);
   U5512 : NAND2_X1 port map( A1 => n1559, A2 => n16784, ZN => n1558);
   U5513 : NAND2_X1 port map( A1 => n1560, A2 => n8014, ZN => n7827);
   U5514 : NOR2_X1 port map( A1 => n1560, A2 => n20154, ZN => n7086);
   U5515 : NAND2_X1 port map( A1 => n7077, A2 => n1560, ZN => n7107);
   U5516 : NAND2_X1 port map( A1 => n5367, A2 => n1562, ZN => n1561);
   U5517 : NOR2_X1 port map( A1 => n5323, A2 => n5368, ZN => n1562);
   U5518 : NAND3_X1 port map( A1 => n4019, A2 => n5401, A3 => n1564, ZN => 
                           n1563);
   U5519 : NAND2_X1 port map( A1 => n5367, A2 => n5393, ZN => n1564);
   U5520 : NAND3_X1 port map( A1 => n15061, A2 => n15306, A3 => n1640, ZN => 
                           n14187);
   U5521 : NAND2_X1 port map( A1 => n8358, A2 => n1565, ZN => n7696);
   U5522 : NAND2_X1 port map( A1 => n8357, A2 => n1565, ZN => n2931);
   U5523 : INV_X1 port map( A => n7741, ZN => n1565);
   U5524 : INV_X1 port map( A => n4479, ZN => n3967);
   U5525 : NAND2_X1 port map( A1 => n4919, A2 => n1793, ZN => n4239);
   U5527 : NAND2_X1 port map( A1 => n1567, A2 => n9023, ZN => n9024);
   U5528 : NAND2_X1 port map( A1 => n8841, A2 => n1567, ZN => n8839);
   U5529 : NAND2_X1 port map( A1 => n1632, A2 => n1566, ZN => n8587);
   U5530 : OR2_X1 port map( A1 => n8836, A2 => n1567, ZN => n1566);
   U5531 : NAND2_X1 port map( A1 => n4721, A2 => n1569, ZN => n5728);
   U5532 : NAND2_X2 port map( A1 => n4704, A2 => n4703, ZN => n6379);
   U5533 : INV_X1 port map( A => n14327, ZN => n14350);
   U5534 : INV_X1 port map( A => n14819, ZN => n1571);
   U5535 : NOR2_X1 port map( A1 => n14353, A2 => n3444, ZN => n1572);
   U5536 : NAND2_X1 port map( A1 => n1574, A2 => n9090, ZN => n8886);
   U5539 : INV_X1 port map( A => n9453, ZN => n1576);
   U5540 : NAND2_X1 port map( A1 => n8562, A2 => n1577, ZN => n9454);
   U5541 : NAND2_X1 port map( A1 => n11953, A2 => n11598, ZN => n11599);
   U5542 : OAI21_X1 port map( B1 => n10953, B2 => n11009, A => n1579, ZN => 
                           n9552);
   U5543 : NAND2_X1 port map( A1 => n11009, A2 => n11149, ZN => n1579);
   U5544 : INV_X1 port map( A => n10953, ZN => n1580);
   U5545 : INV_X1 port map( A => Plaintext(76), ZN => n1581);
   U5547 : MUX2_X1 port map( A => n5024, B => n19788, S => n5022, Z => n5028);
   U5548 : MUX2_X1 port map( A => n8824, B => n8825, S => n9313, Z => n8826);
   U5552 : AND2_X1 port map( A1 => n4217, A2 => n4219, ZN => n1586);
   U5553 : NOR2_X1 port map( A1 => n5826, A2 => n3569, ZN => n1585);
   U5554 : NAND2_X1 port map( A1 => n5823, A2 => n1585, ZN => n3568);
   U5555 : NAND3_X1 port map( A1 => n7866, A2 => n1587, A3 => n9264, ZN => 
                           n8454);
   U5556 : MUX2_X1 port map( A => n9262, B => n7866, S => n9266, Z => n8983);
   U5557 : NAND2_X1 port map( A1 => n10876, A2 => n1588, ZN => n10877);
   U5558 : NOR2_X1 port map( A1 => n1591, A2 => n1589, ZN => n1588);
   U5559 : NAND2_X1 port map( A1 => n11633, A2 => n19755, ZN => n1589);
   U5560 : NAND2_X1 port map( A1 => n14248, A2 => n20377, ZN => n2790);
   U5561 : INV_X1 port map( A => n4574, ZN => n4371);
   U5562 : NAND2_X1 port map( A1 => n12208, A2 => n11808, ZN => n10821);
   U5563 : INV_X1 port map( A => n14656, ZN => n1593);
   U5564 : NAND3_X1 port map( A1 => n5096, A2 => n5098, A3 => n4788, ZN => 
                           n1595);
   U5565 : NAND2_X1 port map( A1 => n5097, A2 => n5096, ZN => n1594);
   U5566 : NAND2_X1 port map( A1 => n20202, A2 => n5088, ZN => n1596);
   U5567 : XNOR2_X2 port map( A => Key(110), B => Plaintext(110), ZN => n5088);
   U5568 : NAND2_X1 port map( A1 => n1598, A2 => n2460, ZN => n1597);
   U5569 : NAND2_X1 port map( A1 => n2461, A2 => n5094, ZN => n1598);
   U5570 : INV_X1 port map( A => n10677, ZN => n1601);
   U5572 : INV_X1 port map( A => n9221, ZN => n1603);
   U5573 : NAND2_X1 port map( A1 => n1603, A2 => n1604, ZN => n8226);
   U5574 : INV_X1 port map( A => n9217, ZN => n1604);
   U5575 : NAND3_X1 port map( A1 => n5172, A2 => n5657, A3 => n6105, ZN => 
                           n2558);
   U5576 : NAND2_X1 port map( A1 => n11093, A2 => n11445, ZN => n1606);
   U5577 : OAI21_X1 port map( B1 => n11093, B2 => n10845, A => n1606, ZN => 
                           n10727);
   U5578 : AOI21_X1 port map( B1 => n1606, B2 => n11444, A => n19920, ZN => 
                           n11450);
   U5579 : NAND2_X1 port map( A1 => n8271, A2 => n1607, ZN => n7720);
   U5580 : NAND2_X1 port map( A1 => n1608, A2 => n8141, ZN => n2156);
   U5583 : NAND3_X1 port map( A1 => n11509, A2 => n10935, A3 => n259, ZN => 
                           n10908);
   U5584 : MUX2_X1 port map( A => n10937, B => n259, S => n19864, Z => n10938);
   U5586 : INV_X1 port map( A => n14935, ZN => n1614);
   U5588 : NAND2_X1 port map( A1 => n15188, A2 => n1611, ZN => n1610);
   U5589 : AND2_X1 port map( A1 => n15503, A2 => n15822, ZN => n1611);
   U5591 : NAND2_X1 port map( A1 => n15504, A2 => n15505, ZN => n1615);
   U5593 : NAND2_X1 port map( A1 => n1620, A2 => n5660, ZN => n1619);
   U5594 : NAND2_X1 port map( A1 => n6111, A2 => n6109, ZN => n1621);
   U5595 : NAND2_X1 port map( A1 => n5658, A2 => n5657, ZN => n1622);
   U5596 : NAND2_X1 port map( A1 => n5659, A2 => n6105, ZN => n1623);
   U5597 : OAI21_X1 port map( B1 => n14303, B2 => n14481, A => n14434, ZN => 
                           n1628);
   U5598 : NAND2_X1 port map( A1 => n14311, A2 => n237, ZN => n1624);
   U5599 : NAND2_X1 port map( A1 => n14310, A2 => n14522, ZN => n1625);
   U5600 : OAI22_X1 port map( A1 => n15553, A2 => n1626, B1 => n14978, B2 => 
                           n15413, ZN => n14907);
   U5601 : NAND2_X1 port map( A1 => n15413, A2 => n15551, ZN => n1626);
   U5602 : NAND2_X1 port map( A1 => n1628, A2 => n1627, ZN => n15409);
   U5603 : NAND2_X1 port map( A1 => n1629, A2 => n14487, ZN => n1627);
   U5604 : NAND2_X1 port map( A1 => n14302, A2 => n14482, ZN => n1629);
   U5605 : INV_X1 port map( A => n15551, ZN => n14905);
   U5606 : NAND2_X1 port map( A1 => n1632, A2 => n19857, ZN => n1630);
   U5607 : INV_X1 port map( A => n8672, ZN => n1632);
   U5608 : NAND2_X1 port map( A1 => n8515, A2 => n1632, ZN => n2024);
   U5609 : MUX2_X1 port map( A => n1632, B => n9024, S => n19857, Z => n9025);
   U5610 : NAND2_X1 port map( A1 => n249, A2 => n12352, ZN => n1633);
   U5611 : NOR2_X2 port map( A1 => n1635, A2 => n1634, ZN => n13070);
   U5612 : NOR2_X1 port map( A1 => n11032, A2 => n1637, ZN => n1636);
   U5613 : INV_X1 port map( A => n19769, ZN => n1637);
   U5614 : INV_X1 port map( A => n1638, ZN => n13414);
   U5615 : NAND2_X1 port map( A1 => n2902, A2 => n2905, ZN => n1638);
   U5616 : NAND2_X1 port map( A1 => n1638, A2 => n15221, ZN => n15770);
   U5617 : NAND2_X1 port map( A1 => n1639, A2 => n15666, ZN => n15668);
   U5618 : AND2_X1 port map( A1 => n234, A2 => n1638, ZN => n15664);
   U5619 : NAND2_X1 port map( A1 => n15772, A2 => n1638, ZN => n15774);
   U5620 : AOI22_X2 port map( A1 => n3254, A2 => n14369, B1 => n3253, B2 => 
                           n3299, ZN => n1640);
   U5621 : NAND2_X1 port map( A1 => n1640, A2 => n15309, ZN => n14177);
   U5622 : OR2_X1 port map( A1 => n15310, A2 => n1640, ZN => n14188);
   U5623 : NAND3_X1 port map( A1 => n3649, A2 => n12685, A3 => n12647, ZN => 
                           n1641);
   U5624 : INV_X1 port map( A => n14731, ZN => n14726);
   U5625 : XNOR2_X2 port map( A => n13402, B => n13401, ZN => n14731);
   U5626 : NAND2_X1 port map( A1 => n255, A2 => n1643, ZN => n12132);
   U5627 : NAND2_X1 port map( A1 => n15498, A2 => n15497, ZN => n1644);
   U5628 : NOR2_X1 port map( A1 => n19512, A2 => n15195, ZN => n15498);
   U5629 : NAND3_X1 port map( A1 => n1647, A2 => n1649, A3 => n19512, ZN => 
                           n1645);
   U5630 : NAND4_X1 port map( A1 => n15508, A2 => n15821, A3 => n15820, A4 => 
                           n1646, ZN => n16374);
   U5631 : NAND3_X1 port map( A1 => n15822, A2 => n13933, A3 => n1758, ZN => 
                           n1646);
   U5632 : NAND2_X1 port map( A1 => n15192, A2 => n15501, ZN => n1647);
   U5633 : NAND2_X1 port map( A1 => n15499, A2 => n15500, ZN => n1649);
   U5634 : NAND2_X1 port map( A1 => n3819, A2 => n15501, ZN => n1650);
   U5635 : NAND3_X2 port map( A1 => n6402, A2 => n3808, A3 => n6401, ZN => 
                           n9453);
   U5636 : NAND2_X1 port map( A1 => n1652, A2 => n1576, ZN => n1651);
   U5638 : NAND2_X1 port map( A1 => n10650, A2 => n20516, ZN => n8400);
   U5639 : MUX2_X1 port map( A => n11161, B => n10649, S => n20516, Z => n10652
                           );
   U5640 : MUX2_X1 port map( A => n10945, B => n11159, S => n11155, Z => n9557)
                           ;
   U5641 : NOR2_X1 port map( A1 => n19872, A2 => n20516, ZN => n9556);
   U5642 : OAI211_X2 port map( C1 => n15133, C2 => n19848, A => n2105, B => 
                           n1655, ZN => n16893);
   U5643 : NAND2_X1 port map( A1 => n1656, A2 => n15132, ZN => n1655);
   U5644 : NAND2_X1 port map( A1 => n9010, A2 => n19490, ZN => n1658);
   U5645 : NAND2_X1 port map( A1 => n9006, A2 => n8895, ZN => n9010);
   U5647 : XNOR2_X1 port map( A => n1659, B => n2423, ZN => Ciphertext(30));
   U5648 : NAND2_X1 port map( A1 => n18518, A2 => n19773, ZN => n18505);
   U5649 : NAND2_X1 port map( A1 => n1662, A2 => n18505, ZN => n1661);
   U5650 : NAND2_X1 port map( A1 => n18504, A2 => n20492, ZN => n1662);
   U5651 : NAND2_X1 port map( A1 => n11091, A2 => n11090, ZN => n1663);
   U5652 : NAND2_X1 port map( A1 => n11086, A2 => n11110, ZN => n1664);
   U5653 : NAND2_X1 port map( A1 => n1665, A2 => n289, ZN => n4871);
   U5654 : NAND2_X1 port map( A1 => n4381, A2 => n4866, ZN => n1665);
   U5655 : INV_X1 port map( A => n4864, ZN => n4865);
   U5657 : XNOR2_X2 port map( A => n1666, B => n1667, ZN => n14148);
   U5658 : XNOR2_X1 port map( A => n13754, B => n13753, ZN => n1666);
   U5659 : XNOR2_X1 port map( A => n13758, B => n13759, ZN => n1667);
   U5660 : NAND2_X1 port map( A1 => n19154, A2 => n19708, ZN => n1668);
   U5663 : NAND2_X1 port map( A1 => n10970, A2 => n11553, ZN => n3488);
   U5664 : OR2_X1 port map( A1 => n18498, A2 => n18497, ZN => n1675);
   U5665 : NAND3_X1 port map( A1 => n16257, A2 => n16256, A3 => n1674, ZN => 
                           n16259);
   U5666 : OAI211_X1 port map( C1 => n1676, C2 => n17640, A => n18500, B => 
                           n1675, ZN => n1674);
   U5667 : INV_X1 port map( A => n18498, ZN => n1676);
   U5668 : NAND2_X1 port map( A1 => n7691, A2 => n7746, ZN => n1677);
   U5669 : NAND2_X1 port map( A1 => n3447, A2 => n7750, ZN => n1678);
   U5670 : AOI21_X1 port map( B1 => n11418, B2 => n10829, A => n1680, ZN => 
                           n3046);
   U5671 : INV_X1 port map( A => n11131, ZN => n1680);
   U5672 : NAND2_X1 port map( A1 => n1681, A2 => n990, ZN => n11423);
   U5673 : NAND2_X1 port map( A1 => n11418, A2 => n11051, ZN => n1681);
   U5674 : INV_X1 port map( A => n15754, ZN => n1683);
   U5676 : NAND2_X1 port map( A1 => n15589, A2 => n14039, ZN => n1682);
   U5677 : NAND2_X1 port map( A1 => n1683, A2 => n15758, ZN => n15589);
   U5679 : NAND2_X1 port map( A1 => n1686, A2 => n14288, ZN => n14024);
   U5680 : INV_X1 port map( A => n14659, ZN => n1686);
   U5681 : NAND2_X1 port map( A1 => n199, A2 => n20266, ZN => n14659);
   U5682 : INV_X1 port map( A => n14547, ZN => n14023);
   U5683 : NAND2_X1 port map( A1 => n2467, A2 => n6046, ZN => n1687);
   U5684 : NAND2_X1 port map( A1 => n12634, A2 => n180, ZN => n1688);
   U5685 : NAND2_X1 port map( A1 => n12633, A2 => n12634, ZN => n1689);
   U5686 : NOR2_X2 port map( A1 => n8796, A2 => n8793, ZN => n9218);
   U5687 : OAI21_X1 port map( B1 => n8176, B2 => n19901, A => n1691, ZN => 
                           n1690);
   U5688 : NAND2_X1 port map( A1 => n1692, A2 => n19901, ZN => n1691);
   U5689 : INV_X1 port map( A => n8178, ZN => n1692);
   U5690 : NAND2_X1 port map( A1 => n282, A2 => n8157, ZN => n8256);
   U5691 : XNOR2_X1 port map( A => n1694, B => n6840, ZN => n1693);
   U5692 : XNOR2_X1 port map( A => n6842, B => n6843, ZN => n1694);
   U5693 : NAND2_X1 port map( A1 => n1695, A2 => n5743, ZN => n5203);
   U5694 : AOI21_X1 port map( B1 => n1695, B2 => n5749, A => n5743, ZN => n5180
                           );
   U5695 : NOR2_X1 port map( A1 => n15645, A2 => n15256, ZN => n15258);
   U5696 : NAND2_X1 port map( A1 => n1699, A2 => n20266, ZN => n1696);
   U5697 : NAND2_X1 port map( A1 => n1698, A2 => n14653, ZN => n1697);
   U5698 : NAND2_X1 port map( A1 => n14653, A2 => n14656, ZN => n3281);
   U5700 : NAND2_X1 port map( A1 => n18425, A2 => n19997, ZN => n2545);
   U5701 : NOR2_X1 port map( A1 => n18427, A2 => n19997, ZN => n18415);
   U5702 : NAND2_X1 port map( A1 => n18427, A2 => n19997, ZN => n18404);
   U5703 : OAI21_X1 port map( B1 => n18412, B2 => n19997, A => n18425, ZN => 
                           n16491);
   U5704 : NAND2_X1 port map( A1 => n18406, A2 => n1701, ZN => n18408);
   U5705 : AND2_X1 port map( A1 => n9532, A2 => n1703, ZN => n1704);
   U5706 : NAND3_X1 port map( A1 => n8592, A2 => n9531, A3 => n9358, ZN => 
                           n1703);
   U5707 : NAND2_X1 port map( A1 => n9533, A2 => n1704, ZN => n9534);
   U5708 : NAND2_X1 port map( A1 => n1706, A2 => n5529, ZN => n1705);
   U5709 : NAND2_X1 port map( A1 => n5562, A2 => n1707, ZN => n1706);
   U5710 : NAND2_X1 port map( A1 => n5563, A2 => n5569, ZN => n1707);
   U5711 : NAND2_X1 port map( A1 => n6036, A2 => n5532, ZN => n6035);
   U5712 : NAND2_X1 port map( A1 => n5562, A2 => n5563, ZN => n6037);
   U5713 : NAND2_X1 port map( A1 => n10958, A2 => n11145, ZN => n1710);
   U5714 : NAND2_X1 port map( A1 => n10959, A2 => n1721, ZN => n1711);
   U5715 : AOI21_X1 port map( B1 => n3486, B2 => n17236, A => n19374, ZN => 
                           n1712);
   U5716 : NAND2_X1 port map( A1 => n1716, A2 => n1715, ZN => n1714);
   U5717 : NAND2_X1 port map( A1 => n18077, A2 => n20111, ZN => n1715);
   U5718 : NAND2_X1 port map( A1 => n2794, A2 => n1717, ZN => n1716);
   U5719 : INV_X1 port map( A => n18394, ZN => n1717);
   U5720 : OAI22_X1 port map( A1 => n17241, A2 => n19823, B1 => n812, B2 => 
                           n20354, ZN => n17242);
   U5721 : NOR2_X1 port map( A1 => n17243, A2 => n1718, ZN => n16463);
   U5722 : NAND2_X1 port map( A1 => n20354, A2 => n19823, ZN => n16461);
   U5723 : NAND2_X1 port map( A1 => n19823, A2 => n17245, ZN => n18541);
   U5724 : AND3_X1 port map( A1 => n17480, A2 => n17479, A3 => n1718, ZN => 
                           n17481);
   U5725 : MUX2_X1 port map( A => n20354, B => n17480, S => n1718, Z => n16809)
                           ;
   U5726 : INV_X1 port map( A => n5879, ZN => n5980);
   U5727 : NAND2_X1 port map( A1 => n5320, A2 => n6068, ZN => n5879);
   U5728 : INV_X1 port map( A => n11145, ZN => n1721);
   U5729 : NAND2_X1 port map( A1 => n14442, A2 => n14168, ZN => n1724);
   U5730 : NAND3_X1 port map( A1 => n1726, A2 => n7978, A3 => n7981, ZN => 
                           n6318);
   U5731 : NAND2_X1 port map( A1 => n1730, A2 => n18078, ZN => n1729);
   U5732 : NAND3_X1 port map( A1 => n1732, A2 => n18376, A3 => n1733, ZN => 
                           n1730);
   U5733 : NAND2_X1 port map( A1 => n19763, A2 => n20361, ZN => n1732);
   U5734 : NAND2_X1 port map( A1 => n11586, A2 => n12128, ZN => n11759);
   U5735 : NAND2_X1 port map( A1 => n11642, A2 => n1734, ZN => n11644);
   U5736 : AND2_X1 port map( A1 => n11586, A2 => n12126, ZN => n1734);
   U5737 : NAND3_X1 port map( A1 => n11642, A2 => n11586, A3 => n882, ZN => 
                           n11643);
   U5738 : NAND3_X1 port map( A1 => n2499, A2 => n8786, A3 => n9145, ZN => 
                           n1736);
   U5739 : NAND2_X1 port map( A1 => n1740, A2 => n3281, ZN => n1739);
   U5740 : NAND2_X1 port map( A1 => n1742, A2 => n14023, ZN => n1741);
   U5741 : NAND2_X1 port map( A1 => n3281, A2 => n3280, ZN => n1742);
   U5742 : NAND2_X1 port map( A1 => n13221, A2 => n1744, ZN => n1743);
   U5743 : NAND2_X1 port map( A1 => n5844, A2 => n1746, ZN => n5850);
   U5744 : NAND3_X1 port map( A1 => n11142, A2 => n20366, A3 => n10960, ZN => 
                           n1747);
   U5746 : NAND2_X1 port map( A1 => n1749, A2 => n11145, ZN => n1748);
   U5747 : XNOR2_X2 port map( A => n9505, B => n9504, ZN => n11145);
   U5749 : INV_X1 port map( A => n8823, ZN => n1751);
   U5750 : NAND3_X1 port map( A1 => n9307, A2 => n9313, A3 => n1754, ZN => 
                           n1753);
   U5752 : NAND2_X1 port map( A1 => n12500, A2 => n12499, ZN => n12347);
   U5753 : AND2_X1 port map( A1 => n1763, A2 => n1762, ZN => n14308);
   U5754 : NAND2_X1 port map( A1 => n14307, A2 => n13868, ZN => n1763);
   U5755 : NAND2_X1 port map( A1 => n1764, A2 => n5115, ZN => n4838);
   U5756 : OAI21_X1 port map( B1 => n169, B2 => n2042, A => n4417, ZN => n1764)
                           ;
   U5757 : NAND2_X1 port map( A1 => n8380, A2 => n8132, ZN => n8389);
   U5758 : NAND2_X1 port map( A1 => n8829, A2 => n9029, ZN => n1765);
   U5760 : NAND2_X1 port map( A1 => n5826, A2 => n3569, ZN => n1832);
   U5762 : NAND2_X1 port map( A1 => n4235, A2 => n4234, ZN => n1769);
   U5763 : NAND2_X1 port map( A1 => n4236, A2 => n4905, ZN => n1768);
   U5764 : OAI21_X1 port map( B1 => n5621, B2 => n6129, A => n1770, ZN => n5262
                           );
   U5766 : NAND2_X1 port map( A1 => n1774, A2 => n1773, ZN => n1772);
   U5767 : INV_X1 port map( A => n19302, ZN => n1773);
   U5768 : MUX2_X1 port map( A => n19292, B => n19284, S => n19299, Z => n1774)
                           ;
   U5769 : NAND2_X1 port map( A1 => n19912, A2 => n1776, ZN => n4181);
   U5770 : NAND2_X1 port map( A1 => n1776, A2 => n5796, ZN => n5793);
   U5771 : OAI22_X1 port map( A1 => n5301, A2 => n5791, B1 => n5428, B2 => 
                           n1776, ZN => n4184);
   U5773 : NAND2_X1 port map( A1 => n1778, A2 => n19663, ZN => n8714);
   U5775 : OAI21_X1 port map( B1 => n11769, B2 => n1779, A => n12288, ZN => 
                           n11465);
   U5776 : INV_X1 port map( A => n182, ZN => n1779);
   U5777 : XNOR2_X1 port map( A => n15739, B => n1780, ZN => n16094);
   U5778 : AND3_X2 port map( A1 => n15278, A2 => n15279, A3 => n15280, ZN => 
                           n15739);
   U5779 : XNOR2_X1 port map( A => n15739, B => n1781, ZN => n16689);
   U5780 : XNOR2_X1 port map( A => n15739, B => n1782, ZN => n15291);
   U5781 : XNOR2_X1 port map( A => n15739, B => n1783, ZN => n16907);
   U5782 : XNOR2_X1 port map( A => n15739, B => n2417, ZN => n17412);
   U5783 : NAND2_X1 port map( A1 => n19521, A2 => n1785, ZN => n1784);
   U5784 : XNOR2_X1 port map( A => n1786, B => n13570, ZN => n13402);
   U5785 : INV_X1 port map( A => n13428, ZN => n1786);
   U5786 : XNOR2_X1 port map( A => n1787, B => n13428, ZN => n11901);
   U5787 : INV_X1 port map( A => n11862, ZN => n1787);
   U5788 : NAND2_X1 port map( A1 => n11480, A2 => n1788, ZN => n2897);
   U5791 : NAND3_X1 port map( A1 => n20206, A2 => n15121, A3 => n14514, ZN => 
                           n1790);
   U5792 : INV_X1 port map( A => n8232, ZN => n1791);
   U5794 : NAND2_X1 port map( A1 => n4966, A2 => n3593, ZN => n1792);
   U5795 : NAND2_X1 port map( A1 => n1793, A2 => n4482, ZN => n4966);
   U5796 : INV_X1 port map( A => n4479, ZN => n1793);
   U5797 : NOR2_X1 port map( A1 => n14450, A2 => n14449, ZN => n1795);
   U5799 : XNOR2_X2 port map( A => n12867, B => n12866, ZN => n14450);
   U5800 : AOI22_X2 port map( A1 => n1794, A2 => n14179, B1 => n14450, B2 => 
                           n13560, ZN => n15237);
   U5801 : AND2_X1 port map( A1 => n19510, A2 => n18682, ZN => n18669);
   U5802 : AND2_X1 port map( A1 => n18688, A2 => n18682, ZN => n1796);
   U5803 : NAND2_X1 port map( A1 => n19510, A2 => n1796, ZN => n1800);
   U5804 : XNOR2_X1 port map( A => n1797, B => n17024, ZN => Ciphertext(68));
   U5805 : NAND3_X1 port map( A1 => n1800, A2 => n1799, A3 => n1798, ZN => 
                           n1797);
   U5806 : NAND2_X1 port map( A1 => n18668, A2 => n19510, ZN => n1798);
   U5807 : OAI21_X1 port map( B1 => n5697, B2 => n19804, A => n1801, ZN => 
                           n5698);
   U5808 : NAND2_X1 port map( A1 => n5699, A2 => n5968, ZN => n1801);
   U5809 : NAND3_X1 port map( A1 => n20272, A2 => n15121, A3 => n1802, ZN => 
                           n15123);
   U5810 : AOI22_X1 port map( A1 => n20206, A2 => n1802, B1 => n15121, B2 => 
                           n14520, ZN => n14185);
   U5811 : MUX2_X1 port map( A => n14516, B => n20206, S => n15120, Z => n14521
                           );
   U5812 : MUX2_X1 port map( A => n14514, B => n13562, S => n15120, Z => n13565
                           );
   U5814 : INV_X1 port map( A => n6184, ZN => n2865);
   U5815 : OR2_X1 port map( A1 => n5846, A2 => n6184, ZN => n1805);
   U5816 : NAND2_X1 port map( A1 => n288, A2 => n6184, ZN => n1806);
   U5817 : NAND2_X1 port map( A1 => n13856, A2 => n954, ZN => n14195);
   U5820 : NAND2_X1 port map( A1 => n1807, A2 => n5717, ZN => n3605);
   U5821 : NAND2_X1 port map( A1 => n14355, A2 => n1808, ZN => n13938);
   U5822 : NAND2_X1 port map( A1 => n14419, A2 => n1808, ZN => n3180);
   U5823 : NAND2_X1 port map( A1 => n8811, A2 => n8813, ZN => n9121);
   U5824 : NAND2_X1 port map( A1 => n11114, A2 => n11458, ZN => n11453);
   U5825 : INV_X1 port map( A => n11458, ZN => n1812);
   U5826 : INV_X1 port map( A => n11110, ZN => n11451);
   U5827 : MUX2_X1 port map( A => n11454, B => n11088, S => n11110, Z => n1814)
                           ;
   U5828 : NAND2_X1 port map( A1 => n15885, A2 => n15335, ZN => n1815);
   U5829 : NAND2_X1 port map( A1 => n1817, A2 => n16016, ZN => n1816);
   U5830 : AOI22_X1 port map( A1 => n13968, A2 => n3473, B1 => n15334, B2 => 
                           n16009, ZN => n1818);
   U5831 : INV_X1 port map( A => n14736, ZN => n1819);
   U5833 : NAND2_X1 port map( A1 => n14270, A2 => n1821, ZN => n1820);
   U5834 : OR2_X1 port map( A1 => n14569, A2 => n14736, ZN => n1821);
   U5835 : NAND2_X1 port map( A1 => n18327, A2 => n19168, ZN => n18320);
   U5836 : NAND2_X1 port map( A1 => n9326, A2 => n9331, ZN => n1822);
   U5838 : OR2_X1 port map( A1 => n954, A2 => n15313, ZN => n11988);
   U5839 : XNOR2_X1 port map( A => n3787, B => n9315, ZN => n1823);
   U5840 : MUX2_X1 port map( A => n7976, B => n7975, S => n7974, Z => n1825);
   U5841 : OAI21_X1 port map( B1 => n12351, B2 => n19768, A => n12350, ZN => 
                           n12357);
   U5842 : NAND2_X1 port map( A1 => n12755, A2 => n245, ZN => n1827);
   U5843 : INV_X1 port map( A => n4034, ZN => n2468);
   U5845 : NAND3_X1 port map( A1 => n3164, A2 => n20363, A3 => n12537, ZN => 
                           n11806);
   U5846 : NAND2_X1 port map( A1 => n11547, A2 => n11548, ZN => n10068);
   U5847 : NAND3_X1 port map( A1 => n19530, A2 => n20424, A3 => n14020, ZN => 
                           n15757);
   U5848 : NAND2_X1 port map( A1 => n5824, A2 => n1832, ZN => n5831);
   U5849 : OR2_X1 port map( A1 => n6129, A2 => n5623, ZN => n5694);
   U5851 : NAND2_X1 port map( A1 => n317, A2 => n8937, ZN => n8944);
   U5852 : NAND2_X1 port map( A1 => n1834, A2 => n1833, ZN => n7583);
   U5853 : NAND2_X1 port map( A1 => n8297, A2 => n5941, ZN => n1833);
   U5855 : NAND2_X1 port map( A1 => n11395, A2 => n11297, ZN => n10860);
   U5856 : NAND2_X1 port map( A1 => n1837, A2 => n1836, ZN => n5254);
   U5857 : NAND2_X1 port map( A1 => n5401, A2 => n5323, ZN => n1836);
   U5858 : NAND2_X1 port map( A1 => n5393, A2 => n1838, ZN => n1837);
   U5859 : NAND3_X1 port map( A1 => n7716, A2 => n7687, A3 => n8131, ZN => 
                           n1839);
   U5860 : OR2_X1 port map( A1 => n4866, A2 => n4651, ZN => n4870);
   U5861 : AND2_X1 port map( A1 => n8291, A2 => n8292, ZN => n3406);
   U5862 : NOR2_X1 port map( A1 => n8381, A2 => n163, ZN => n7714);
   U5864 : OR2_X1 port map( A1 => n12207, A2 => n247, ZN => n12188);
   U5866 : INV_X1 port map( A => n9580, ZN => n9578);
   U5867 : NAND2_X1 port map( A1 => n19519, A2 => n1841, ZN => n9580);
   U5870 : XNOR2_X1 port map( A => n7040, B => n1842, ZN => n4939);
   U5871 : XNOR2_X1 port map( A => n4780, B => n4781, ZN => n1842);
   U5872 : XNOR2_X1 port map( A => n1843, B => n18503, ZN => Ciphertext(29));
   U5875 : NAND2_X1 port map( A1 => n7606, A2 => n8184, ZN => n7892);
   U5876 : NAND2_X1 port map( A1 => n2614, A2 => n2615, ZN => n5982);
   U5877 : NAND2_X1 port map( A1 => n19752, A2 => n15531, ZN => n15082);
   U5878 : INV_X1 port map( A => n3241, ZN => n12358);
   U5879 : NAND2_X1 port map( A1 => n14516, A2 => n14321, ZN => n13562);
   U5880 : NAND2_X1 port map( A1 => n17518, A2 => n17517, ZN => n17581);
   U5881 : XNOR2_X1 port map( A => n1845, B => n18587, ZN => Ciphertext(51));
   U5882 : NAND3_X1 port map( A1 => n3411, A2 => n18586, A3 => n18582, ZN => 
                           n1845);
   U5883 : OAI21_X1 port map( B1 => n5995, B2 => n5999, A => n1846, ZN => n5275
                           );
   U5884 : NAND2_X1 port map( A1 => n5995, A2 => n5998, ZN => n1846);
   U5885 : NAND2_X1 port map( A1 => n1371, A2 => n11722, ZN => n3676);
   U5886 : NAND3_X1 port map( A1 => n11284, A2 => n19779, A3 => n11282, ZN => 
                           n1847);
   U5887 : NAND2_X1 port map( A1 => n10999, A2 => n10947, ZN => n1848);
   U5888 : XOR2_X1 port map( A => n10441, B => n10299, Z => n2900);
   U5889 : XNOR2_X1 port map( A => n13239, B => n3237, ZN => n13240);
   U5891 : NAND2_X1 port map( A1 => n14578, A2 => n14740, ZN => n1849);
   U5893 : NAND2_X2 port map( A1 => n9078, A2 => n9079, ZN => n10382);
   U5894 : NAND2_X1 port map( A1 => n8180, A2 => n8179, ZN => n1851);
   U5896 : NAND3_X1 port map( A1 => n2931, A2 => n2932, A3 => n8359, ZN => 
                           n2933);
   U5897 : XNOR2_X2 port map( A => Key(19), B => Plaintext(19), ZN => n4979);
   U5898 : NAND2_X1 port map( A1 => n1853, A2 => n1852, ZN => n10857);
   U5899 : NAND2_X1 port map( A1 => n11329, A2 => n11330, ZN => n1852);
   U5903 : OAI21_X1 port map( B1 => n14401, B2 => n19908, A => n14400, ZN => 
                           n3047);
   U5904 : NAND3_X1 port map( A1 => n12758, A2 => n3702, A3 => n1856, ZN => 
                           n13002);
   U5905 : AOI22_X1 port map( A1 => n12755, A2 => n12754, B1 => n12756, B2 => 
                           n12759, ZN => n1856);
   U5906 : XOR2_X1 port map( A => n7305, B => n6484, Z => n1863);
   U5907 : NAND3_X2 port map( A1 => n2798, A2 => n2802, A3 => n2801, ZN => 
                           n17098);
   U5908 : NAND3_X1 port map( A1 => n12813, A2 => n19626, A3 => n11803, ZN => 
                           n3169);
   U5909 : NOR2_X1 port map( A1 => n9137, A2 => n263, ZN => n9138);
   U5910 : NOR2_X1 port map( A1 => n15545, A2 => n15406, ZN => n2799);
   U5911 : NAND2_X1 port map( A1 => n4950, A2 => n4912, ZN => n4909);
   U5913 : NAND2_X1 port map( A1 => n1860, A2 => n1859, ZN => n1858);
   U5914 : NAND2_X1 port map( A1 => n201, A2 => n12502, ZN => n1860);
   U5915 : NAND2_X1 port map( A1 => n19775, A2 => n1862, ZN => n18004);
   U5916 : INV_X1 port map( A => n15394, ZN => n2968);
   U5917 : NAND2_X1 port map( A1 => n7420, A2 => n2886, ZN => n7873);
   U5918 : NAND3_X1 port map( A1 => n20157, A2 => n1819, A3 => n14574, ZN => 
                           n13263);
   U5919 : NAND2_X2 port map( A1 => n2403, A2 => n1864, ZN => n7296);
   U5920 : NAND2_X1 port map( A1 => n5417, A2 => n5226, ZN => n1864);
   U5922 : INV_X1 port map( A => n1866, ZN => n1865);
   U5923 : NAND2_X1 port map( A1 => n5842, A2 => n6166, ZN => n1868);
   U5925 : NAND2_X1 port map( A1 => n957, A2 => n5700, ZN => n1870);
   U5926 : OAI21_X1 port map( B1 => n5450, B2 => n5449, A => n5971, ZN => n1871
                           );
   U5927 : NAND2_X1 port map( A1 => n12010, A2 => n12364, ZN => n12011);
   U5930 : NAND3_X2 port map( A1 => n8393, A2 => n8394, A3 => n966, ZN => 
                           n10236);
   U5931 : NAND2_X1 port map( A1 => n12340, A2 => n11974, ZN => n11824);
   U5932 : OAI211_X2 port map( C1 => n14201, C2 => n1262, A => n2790, B => 
                           n1873, ZN => n15071);
   U5933 : NAND2_X1 port map( A1 => n14604, A2 => n20513, ZN => n1873);
   U5934 : INV_X1 port map( A => n4347, ZN => n4540);
   U5935 : INV_X1 port map( A => n10685, ZN => n12101);
   U5936 : XNOR2_X2 port map( A => n3916, B => Key(150), ZN => n4754);
   U5938 : INV_X1 port map( A => n12686, ZN => n12647);
   U5939 : XNOR2_X1 port map( A => n1874, B => n18405, ZN => Ciphertext(12));
   U5940 : NAND3_X1 port map( A1 => n18403, A2 => n18402, A3 => n1875, ZN => 
                           n1874);
   U5941 : XNOR2_X1 port map( A => n10411, B => n10412, ZN => n11129);
   U5943 : AOI21_X1 port map( B1 => n19971, B2 => n12072, A => n12601, ZN => 
                           n2911);
   U5944 : INV_X1 port map( A => n12800, ZN => n14342);
   U5945 : OAI22_X1 port map( A1 => n14306, A2 => n14305, B1 => n19742, B2 => 
                           n1876, ZN => n14309);
   U5946 : INV_X1 port map( A => n14729, ZN => n14728);
   U5947 : INV_X1 port map( A => n5868, ZN => n5386);
   U5948 : INV_X1 port map( A => n5116, ZN => n1916);
   U5950 : OAI21_X1 port map( B1 => n7968, B2 => n7927, A => n7969, ZN => n3386
                           );
   U5952 : NAND2_X1 port map( A1 => n12067, A2 => n1879, ZN => n1878);
   U5954 : NAND2_X1 port map( A1 => n1880, A2 => n8804, ZN => n3501);
   U5955 : NAND2_X1 port map( A1 => n2631, A2 => n9209, ZN => n1880);
   U5956 : INV_X1 port map( A => n1903, ZN => n1902);
   U5957 : NOR2_X2 port map( A1 => n4001, A2 => n1881, ZN => n7264);
   U5958 : AOI21_X1 port map( B1 => n2616, B2 => n4000, A => n3999, ZN => n1881
                           );
   U5959 : NAND2_X1 port map( A1 => n2974, A2 => n15431, ZN => n15084);
   U5960 : NAND2_X1 port map( A1 => n3980, A2 => n2071, ZN => n1882);
   U5962 : NAND2_X1 port map( A1 => n4887, A2 => n4945, ZN => n4116);
   U5964 : OR2_X1 port map( A1 => n11884, A2 => n11120, ZN => n11461);
   U5966 : NAND2_X1 port map( A1 => n11495, A2 => n888, ZN => n10729);
   U5967 : NAND3_X1 port map( A1 => n5473, A2 => n5472, A3 => n6034, ZN => 
                           n1886);
   U5968 : NAND2_X1 port map( A1 => n1888, A2 => n1887, ZN => n11085);
   U5969 : NAND2_X1 port map( A1 => n11081, A2 => n11499, ZN => n1887);
   U5970 : NAND2_X1 port map( A1 => n11505, A2 => n11188, ZN => n1888);
   U5971 : NAND2_X1 port map( A1 => n6217, A2 => n1890, ZN => n6970);
   U5972 : NAND2_X1 port map( A1 => n6203, A2 => n1891, ZN => n6217);
   U5973 : NAND2_X1 port map( A1 => n10890, A2 => n11549, ZN => n1893);
   U5975 : NAND2_X1 port map( A1 => n6033, A2 => n2940, ZN => n1895);
   U5978 : OAI211_X1 port map( C1 => n3389, C2 => n20463, A => n1896, B => 
                           n17219, ZN => n18344);
   U5979 : NAND2_X1 port map( A1 => n19383, A2 => n1897, ZN => n1896);
   U5980 : OR2_X1 port map( A1 => n4518, A2 => n4517, ZN => n4519);
   U5981 : NAND3_X1 port map( A1 => n2174, A2 => n9333, A3 => n9330, ZN => 
                           n9336);
   U5982 : NAND2_X1 port map( A1 => n1939, A2 => n3313, ZN => n1898);
   U5985 : NAND2_X1 port map( A1 => n14846, A2 => n3573, ZN => n1901);
   U5986 : XNOR2_X1 port map( A => n7348, B => n7163, ZN => n6744);
   U5987 : OR2_X1 port map( A1 => n4355, A2 => n4313, ZN => n1908);
   U5988 : NAND2_X1 port map( A1 => n17888, A2 => n19947, ZN => n1905);
   U5989 : NAND2_X1 port map( A1 => n17889, A2 => n1907, ZN => n1906);
   U5991 : NAND2_X1 port map( A1 => n11199, A2 => n3051, ZN => n3048);
   U5992 : NAND2_X1 port map( A1 => n10730, A2 => n11493, ZN => n11199);
   U5994 : NAND3_X1 port map( A1 => n4361, A2 => n4358, A3 => n4547, ZN => 
                           n4359);
   U5995 : NAND2_X1 port map( A1 => n1910, A2 => n1909, ZN => n7636);
   U5996 : NAND2_X1 port map( A1 => n7634, A2 => n8212, ZN => n1909);
   U5998 : NAND2_X1 port map( A1 => n9119, A2 => n8328, ZN => n1912);
   U5999 : AND3_X1 port map( A1 => n12629, A2 => n11722, A3 => n11618, ZN => 
                           n11621);
   U6000 : NAND2_X1 port map( A1 => n4066, A2 => n1914, ZN => n4067);
   U6002 : NAND2_X1 port map( A1 => n11296, A2 => n2724, ZN => n1918);
   U6003 : NAND2_X2 port map( A1 => n3591, A2 => n3043, ZN => n6206);
   U6004 : NAND2_X1 port map( A1 => n1919, A2 => n2115, ZN => n5264);
   U6005 : NAND3_X1 port map( A1 => n5804, A2 => n6194, A3 => n5805, ZN => 
                           n2868);
   U6006 : NAND2_X1 port map( A1 => n8375, A2 => n8376, ZN => n8369);
   U6007 : NAND3_X1 port map( A1 => n9327, A2 => n262, A3 => n20008, ZN => 
                           n9337);
   U6008 : NAND2_X1 port map( A1 => n3265, A2 => n3872, ZN => n1920);
   U6009 : NAND3_X2 port map( A1 => n1922, A2 => n4443, A3 => n4444, ZN => 
                           n6138);
   U6011 : NOR2_X1 port map( A1 => n17899, A2 => n1923, ZN => n17900);
   U6012 : NOR2_X1 port map( A1 => n17897, A2 => n1924, ZN => n1923);
   U6013 : NAND2_X1 port map( A1 => n15148, A2 => n15874, ZN => n1925);
   U6014 : NAND3_X1 port map( A1 => n1926, A2 => n1005, A3 => n2742, ZN => 
                           n11640);
   U6015 : NAND2_X1 port map( A1 => n2743, A2 => n3692, ZN => n1926);
   U6018 : NOR2_X1 port map( A1 => n983, A2 => n2874, ZN => n2873);
   U6019 : OAI21_X1 port map( B1 => n8078, B2 => n3654, A => n3653, ZN => n8082
                           );
   U6020 : OAI21_X1 port map( B1 => n3041, B2 => n15412, A => n14980, ZN => 
                           n1968);
   U6021 : NAND2_X1 port map( A1 => n11147, A2 => n11148, ZN => n10708);
   U6022 : XNOR2_X1 port map( A => n13102, B => n13101, ZN => n3373);
   U6023 : XNOR2_X2 port map( A => n3856, B => Key(95), ZN => n5098);
   U6024 : NOR2_X1 port map( A1 => n8510, A2 => n9021, ZN => n8674);
   U6025 : INV_X1 port map( A => n5612, ZN => n6159);
   U6026 : INV_X1 port map( A => n2523, ZN => n12409);
   U6028 : INV_X1 port map( A => n6300, ZN => n7241);
   U6029 : INV_X1 port map( A => n3995, ZN => n4687);
   U6030 : OAI21_X1 port map( B1 => n10935, B2 => n19864, A => n1928, ZN => 
                           n10744);
   U6031 : NAND2_X1 port map( A1 => n10935, A2 => n11573, ZN => n1928);
   U6036 : NAND2_X1 port map( A1 => n1015, A2 => n8841, ZN => n1929);
   U6037 : OAI211_X2 port map( C1 => n12381, C2 => n11732, A => n1931, B => 
                           n1930, ZN => n13642);
   U6038 : NAND2_X1 port map( A1 => n11731, A2 => n12381, ZN => n1930);
   U6039 : NAND2_X1 port map( A1 => n12371, A2 => n20497, ZN => n1931);
   U6040 : MUX2_X1 port map( A => n9114, B => n9221, S => n9113, Z => n9115);
   U6041 : OAI21_X1 port map( B1 => n4646, B2 => n4647, A => n4645, ZN => n4649
                           );
   U6042 : NAND2_X1 port map( A1 => n4646, A2 => n4319, ZN => n4645);
   U6043 : NAND2_X1 port map( A1 => n12007, A2 => n12008, ZN => n12012);
   U6044 : NAND2_X1 port map( A1 => n1934, A2 => n1933, ZN => n1932);
   U6045 : INV_X1 port map( A => n9046, ZN => n1933);
   U6046 : INV_X1 port map( A => n9045, ZN => n1934);
   U6048 : NAND2_X1 port map( A1 => n1935, A2 => n13877, ZN => n14496);
   U6049 : OAI21_X1 port map( B1 => n14492, B2 => n14491, A => n1936, ZN => 
                           n1935);
   U6050 : NAND3_X1 port map( A1 => n10661, A2 => n11244, A3 => n10662, ZN => 
                           n2859);
   U6051 : NAND2_X1 port map( A1 => n10856, A2 => n20095, ZN => n10662);
   U6052 : XNOR2_X2 port map( A => Key(141), B => Plaintext(141), ZN => n4734);
   U6053 : AND2_X1 port map( A1 => n4633, A2 => n4185, ZN => n3728);
   U6054 : OAI211_X1 port map( C1 => n14081, C2 => n20500, A => n1937, B => 
                           n3497, ZN => n3496);
   U6055 : NAND2_X1 port map( A1 => n1938, A2 => n14801, ZN => n1937);
   U6056 : INV_X1 port map( A => n2628, ZN => n1938);
   U6058 : NAND2_X1 port map( A1 => n3385, A2 => n9046, ZN => n9037);
   U6059 : INV_X1 port map( A => n4708, ZN => n4771);
   U6060 : NOR2_X1 port map( A1 => n19958, A2 => n3315, ZN => n1939);
   U6061 : XNOR2_X1 port map( A => n1940, B => n7213, ZN => n7215);
   U6062 : XNOR2_X1 port map( A => n7210, B => n7360, ZN => n1940);
   U6063 : NAND2_X1 port map( A1 => n19507, A2 => n4969, ZN => n4480);
   U6064 : OR2_X1 port map( A1 => n4908, A2 => n4907, ZN => n1942);
   U6065 : NAND2_X1 port map( A1 => n11111, A2 => n11114, ZN => n1943);
   U6066 : NAND2_X1 port map( A1 => n11112, A2 => n11454, ZN => n1944);
   U6067 : NAND2_X1 port map( A1 => n12387, A2 => n12470, ZN => n1945);
   U6068 : NAND2_X1 port map( A1 => n1948, A2 => n1947, ZN => n6808);
   U6069 : NAND2_X1 port map( A1 => n5215, A2 => n1949, ZN => n1948);
   U6070 : NAND2_X1 port map( A1 => n10710, A2 => n20160, ZN => n10714);
   U6071 : AOI21_X1 port map( B1 => n1950, B2 => n8217, A => n8216, ZN => n8224
                           );
   U6072 : NAND2_X1 port map( A1 => n8219, A2 => n8215, ZN => n1950);
   U6074 : NAND3_X2 port map( A1 => n1954, A2 => n11691, A3 => n1951, ZN => 
                           n13193);
   U6077 : NAND2_X1 port map( A1 => n12123, A2 => n12230, ZN => n1954);
   U6078 : OAI211_X2 port map( C1 => n19809, C2 => n8217, A => n6475, B => 
                           n6474, ZN => n9240);
   U6079 : NOR2_X1 port map( A1 => n15468, A2 => n15469, ZN => n1955);
   U6080 : NAND2_X1 port map( A1 => n4171, A2 => n20143, ZN => n4288);
   U6081 : NAND3_X1 port map( A1 => n151, A2 => n19037, A3 => n1016, ZN => 
                           n19039);
   U6082 : OAI21_X1 port map( B1 => n13275, B2 => n12325, A => n1956, ZN => 
                           n11678);
   U6083 : NAND2_X1 port map( A1 => n13275, A2 => n12513, ZN => n1956);
   U6084 : OAI21_X2 port map( B1 => n6112, B2 => n6113, A => n1957, ZN => n7221
                           );
   U6085 : NAND2_X1 port map( A1 => n6110, A2 => n6109, ZN => n1958);
   U6086 : INV_X1 port map( A => n7711, ZN => n6952);
   U6087 : NAND2_X1 port map( A1 => n6091, A2 => n6088, ZN => n1959);
   U6088 : NAND2_X1 port map( A1 => n2692, A2 => n2693, ZN => n2691);
   U6089 : AND2_X1 port map( A1 => n12417, A2 => n20352, ZN => n12427);
   U6092 : INV_X1 port map( A => n16171, ZN => n3573);
   U6093 : NAND2_X1 port map( A1 => n1963, A2 => n1961, ZN => n9242);
   U6094 : NAND2_X1 port map( A1 => n6610, A2 => n8090, ZN => n1963);
   U6097 : AND2_X1 port map( A1 => n19472, A2 => n17946, ZN => n17774);
   U6098 : OR2_X1 port map( A1 => n7930, A2 => n7933, ZN => n7941);
   U6099 : INV_X1 port map( A => n11211, ZN => n11486);
   U6100 : AND3_X2 port map( A1 => n1965, A2 => n8816, A3 => n1964, ZN => 
                           n10404);
   U6101 : NAND2_X1 port map( A1 => n8819, A2 => n8818, ZN => n1965);
   U6102 : OAI21_X1 port map( B1 => n12535, B2 => n3477, A => n12531, ZN => 
                           n3476);
   U6103 : XNOR2_X1 port map( A => n13136, B => n20170, ZN => n12517);
   U6105 : INV_X1 port map( A => n15127, ZN => n15017);
   U6106 : INV_X1 port map( A => n6031, ZN => n5928);
   U6107 : OAI211_X1 port map( C1 => n14195, C2 => n2731, A => n14194, B => 
                           n14193, ZN => n15615);
   U6108 : NOR2_X1 port map( A1 => n15846, A2 => n15267, ZN => n2529);
   U6110 : XNOR2_X1 port map( A => n3619, B => n6719, ZN => n7286);
   U6111 : XNOR2_X1 port map( A => n2520, B => n2519, ZN => n14012);
   U6112 : OR2_X1 port map( A1 => n15277, A2 => n15601, ZN => n15278);
   U6113 : XNOR2_X1 port map( A => n1966, B => n18428, ZN => Ciphertext(17));
   U6114 : OAI22_X1 port map( A1 => n2546, A2 => n18427, B1 => n18426, B2 => 
                           n18425, ZN => n1966);
   U6115 : AOI21_X1 port map( B1 => n8072, B2 => n2456, A => n585, ZN => n1967)
                           ;
   U6118 : NAND2_X1 port map( A1 => n12591, A2 => n12200, ZN => n11978);
   U6119 : NAND2_X1 port map( A1 => n1968, A2 => n3042, ZN => n16944);
   U6120 : NAND3_X1 port map( A1 => n20313, A2 => n8537, A3 => n9073, ZN => 
                           n8464);
   U6121 : NAND2_X1 port map( A1 => n11429, A2 => n1970, ZN => n10827);
   U6124 : NAND2_X1 port map( A1 => n11151, A2 => n11152, ZN => n1971);
   U6125 : INV_X1 port map( A => n4510, ZN => n4513);
   U6126 : INV_X1 port map( A => n11880, ZN => n3441);
   U6127 : XNOR2_X1 port map( A => n13345, B => n13346, ZN => n1973);
   U6128 : NAND2_X1 port map( A1 => n15860, A2 => n1974, ZN => n15867);
   U6129 : NAND2_X1 port map( A1 => n8263, A2 => n8153, ZN => n8104);
   U6131 : OAI21_X1 port map( B1 => n11976, B2 => n11977, A => n2160, ZN => 
                           n1975);
   U6132 : NAND2_X1 port map( A1 => n6010, A2 => n19979, ZN => n5502);
   U6133 : NAND2_X1 port map( A1 => n5804, A2 => n5805, ZN => n5808);
   U6134 : NAND2_X1 port map( A1 => n3345, A2 => n17879, ZN => n3344);
   U6135 : NAND2_X2 port map( A1 => n2497, A2 => n7913, ZN => n2499);
   U6136 : NAND2_X1 port map( A1 => n4540, A2 => n4541, ZN => n4543);
   U6137 : NAND2_X1 port map( A1 => n3259, A2 => n5101, ZN => n5103);
   U6138 : NAND3_X1 port map( A1 => n7929, A2 => n9149, A3 => n7928, ZN => 
                           n7943);
   U6140 : OAI21_X1 port map( B1 => n5122, B2 => n5917, A => n5916, ZN => n1978
                           );
   U6141 : INV_X1 port map( A => n11377, ZN => n11329);
   U6142 : OAI211_X1 port map( C1 => n8529, C2 => n9038, A => n1979, B => n7657
                           , ZN => n7658);
   U6143 : AOI22_X2 port map( A1 => n11393, A2 => n11392, B1 => n19750, B2 => 
                           n11391, ZN => n12545);
   U6144 : NOR2_X1 port map( A1 => n3764, A2 => n3762, ZN => n3761);
   U6145 : NOR2_X1 port map( A1 => n3030, A2 => n18869, ZN => n18051);
   U6148 : OR2_X1 port map( A1 => n4171, A2 => n4622, ZN => n4627);
   U6149 : NAND2_X1 port map( A1 => n2291, A2 => n3316, ZN => n1983);
   U6150 : OAI21_X1 port map( B1 => n9451, B2 => n8884, A => n8563, ZN => n9455
                           );
   U6151 : INV_X1 port map( A => n7931, ZN => n2030);
   U6152 : INV_X1 port map( A => n10849, ZN => n13114);
   U6153 : INV_X1 port map( A => n4355, ZN => n4547);
   U6154 : AND2_X1 port map( A1 => n5571, A2 => n5581, ZN => n3533);
   U6155 : XNOR2_X2 port map( A => n3881, B => Key(2), ZN => n4171);
   U6156 : NAND2_X1 port map( A1 => n11674, A2 => n11670, ZN => n11843);
   U6157 : NAND2_X1 port map( A1 => n15745, A2 => n15521, ZN => n14982);
   U6158 : NAND3_X1 port map( A1 => n14486, A2 => n14302, A3 => n14480, ZN => 
                           n13554);
   U6159 : NAND2_X1 port map( A1 => n20263, A2 => n14482, ZN => n14486);
   U6160 : NAND2_X1 port map( A1 => n5804, A2 => n1986, ZN => n5380);
   U6163 : AND2_X1 port map( A1 => n11500, A2 => n11193, ZN => n1988);
   U6164 : AND2_X1 port map( A1 => n14673, A2 => n20424, ZN => n13982);
   U6165 : INV_X1 port map( A => n7443, ZN => n8280);
   U6166 : OR2_X2 port map( A1 => n9195, A2 => n9194, ZN => n10107);
   U6168 : NAND2_X1 port map( A1 => n1989, A2 => n3660, ZN => n3659);
   U6170 : INV_X1 port map( A => n2183, ZN => n12564);
   U6171 : NAND2_X1 port map( A1 => n1991, A2 => n1990, ZN => n2183);
   U6172 : NAND2_X1 port map( A1 => n12263, A2 => n12262, ZN => n1990);
   U6173 : NAND2_X1 port map( A1 => n12261, A2 => n12264, ZN => n1991);
   U6174 : NAND2_X1 port map( A1 => n14721, A2 => n1992, ZN => n15566);
   U6175 : OR2_X1 port map( A1 => n14723, A2 => n19843, ZN => n1992);
   U6177 : OR2_X1 port map( A1 => n4541, A2 => n4347, ZN => n4254);
   U6178 : NAND2_X1 port map( A1 => n1995, A2 => n1993, ZN => n7677);
   U6179 : NAND2_X1 port map( A1 => n7676, A2 => n1994, ZN => n1993);
   U6180 : NAND2_X1 port map( A1 => n8362, A2 => n7675, ZN => n1995);
   U6182 : NAND2_X1 port map( A1 => n15700, A2 => n20145, ZN => n1997);
   U6183 : OAI21_X1 port map( B1 => n14344, B2 => n14789, A => n1999, ZN => 
                           n14104);
   U6184 : NAND2_X1 port map( A1 => n2411, A2 => n2412, ZN => n1999);
   U6185 : OAI21_X1 port map( B1 => n2001, B2 => n2000, A => n18996, ZN => 
                           n18998);
   U6186 : NAND2_X1 port map( A1 => n18991, A2 => n18993, ZN => n2000);
   U6187 : NAND2_X1 port map( A1 => n18994, A2 => n18992, ZN => n2001);
   U6188 : NAND2_X1 port map( A1 => n14723, A2 => n14717, ZN => n14719);
   U6189 : XNOR2_X2 port map( A => n6949, B => n7270, ZN => n8341);
   U6190 : NAND2_X1 port map( A1 => n1062, A2 => n3818, ZN => n2002);
   U6191 : NOR2_X1 port map( A1 => n2813, A2 => n14461, ZN => n2812);
   U6192 : NAND3_X1 port map( A1 => n4593, A2 => n4594, A3 => n6194, ZN => 
                           n4595);
   U6194 : OAI21_X1 port map( B1 => n14939, B2 => n14940, A => n20449, ZN => 
                           n2006);
   U6196 : OAI21_X1 port map( B1 => n15160, B2 => n15159, A => n15195, ZN => 
                           n2007);
   U6198 : NAND2_X1 port map( A1 => n20180, A2 => n20441, ZN => n8217);
   U6199 : NAND2_X1 port map( A1 => n11417, A2 => n11129, ZN => n11419);
   U6200 : NAND2_X1 port map( A1 => n16580, A2 => n2008, ZN => n19338);
   U6201 : OR2_X1 port map( A1 => n16657, A2 => n19372, ZN => n2008);
   U6203 : NAND2_X1 port map( A1 => n2009, A2 => n11410, ZN => n3612);
   U6204 : NAND2_X1 port map( A1 => n11408, A2 => n19736, ZN => n2009);
   U6205 : OAI21_X2 port map( B1 => n3879, B2 => n2010, A => n3878, ZN => n5796
                           );
   U6206 : NAND2_X1 port map( A1 => n4980, A2 => n4978, ZN => n2010);
   U6210 : NAND3_X1 port map( A1 => n3626, A2 => n2013, A3 => n2011, ZN => 
                           n13041);
   U6211 : NAND2_X1 port map( A1 => n12120, A2 => n2012, ZN => n2011);
   U6212 : INV_X1 port map( A => n12124, ZN => n2012);
   U6213 : NAND2_X1 port map( A1 => n12123, A2 => n12227, ZN => n2013);
   U6215 : NAND2_X1 port map( A1 => n19663, A2 => n2476, ZN => n2015);
   U6216 : OAI21_X1 port map( B1 => n1859, B2 => n12500, A => n2016, ZN => 
                           n2864);
   U6217 : NAND2_X1 port map( A1 => n9189, A2 => n6656, ZN => n2425);
   U6218 : NAND2_X1 port map( A1 => n3846, A2 => n4676, ZN => n5114);
   U6219 : OAI21_X1 port map( B1 => n8466, B2 => n8545, A => n2330, ZN => n8468
                           );
   U6220 : OAI22_X1 port map( A1 => n2017, A2 => n8602, B1 => n8949, B2 => 
                           n8951, ZN => n7652);
   U6221 : NAND2_X1 port map( A1 => n8949, A2 => n905, ZN => n2017);
   U6222 : XNOR2_X1 port map( A => n13253, B => n13750, ZN => n2189);
   U6223 : NAND3_X1 port map( A1 => n12148, A2 => n3260, A3 => n19952, ZN => 
                           n2104);
   U6226 : INV_X1 port map( A => n18424, ZN => n2019);
   U6227 : XNOR2_X1 port map( A => n2020, B => n10297, ZN => n10302);
   U6228 : XNOR2_X1 port map( A => n10295, B => n10612, ZN => n2020);
   U6229 : MUX2_X1 port map( A => n8194, B => n7456, S => n8051, Z => n2021);
   U6231 : NAND2_X1 port map( A1 => n5115, A2 => n4676, ZN => n3848);
   U6233 : OAI21_X1 port map( B1 => n8215, B2 => n8219, A => n2026, ZN => n3793
                           );
   U6234 : NAND2_X1 port map( A1 => n8220, A2 => n8219, ZN => n2026);
   U6236 : NAND2_X1 port map( A1 => n2028, A2 => n2027, ZN => n4266);
   U6237 : OAI21_X1 port map( B1 => n4754, B2 => n4563, A => n4567, ZN => n2027
                           );
   U6238 : NAND2_X1 port map( A1 => n4265, A2 => n3131, ZN => n2028);
   U6239 : NAND2_X1 port map( A1 => n12004, A2 => n12005, ZN => n2901);
   U6240 : INV_X1 port map( A => n5483, ZN => n4363);
   U6243 : AOI21_X1 port map( B1 => n11358, B2 => n11127, A => n1039, ZN => 
                           n2029);
   U6244 : NAND2_X1 port map( A1 => n4687, A2 => n178, ZN => n4392);
   U6245 : NAND3_X2 port map( A1 => n2034, A2 => n4758, A3 => n3129, ZN => 
                           n5669);
   U6246 : NOR2_X1 port map( A1 => n3112, A2 => n11177, ZN => n3111);
   U6247 : INV_X1 port map( A => n15644, ZN => n2223);
   U6249 : INV_X1 port map( A => n18033, ZN => n18268);
   U6251 : XNOR2_X1 port map( A => n10324, B => n10323, ZN => n11088);
   U6252 : INV_X1 port map( A => n15341, ZN => n15337);
   U6253 : XNOR2_X2 port map( A => Key(33), B => Plaintext(33), ZN => n4912);
   U6254 : NAND2_X1 port map( A1 => n5324, A2 => n5373, ZN => n5325);
   U6255 : NAND2_X1 port map( A1 => n1838, A2 => n5401, ZN => n5373);
   U6256 : OAI21_X1 port map( B1 => n2548, B2 => n7585, A => n2037, ZN => n3611
                           );
   U6257 : NAND2_X1 port map( A1 => n7312, A2 => n2548, ZN => n2037);
   U6258 : NAND2_X1 port map( A1 => n2040, A2 => n2038, ZN => n14754);
   U6259 : NAND3_X1 port map( A1 => n14054, A2 => n13938, A3 => n2039, ZN => 
                           n2038);
   U6260 : NAND2_X1 port map( A1 => n13941, A2 => n13940, ZN => n2040);
   U6261 : OAI21_X1 port map( B1 => n4675, B2 => n2042, A => n2041, ZN => n3842
                           );
   U6262 : NAND2_X1 port map( A1 => n4675, A2 => n4835, ZN => n2041);
   U6263 : AOI21_X1 port map( B1 => n11399, B2 => n11395, A => n11397, ZN => 
                           n2044);
   U6266 : NAND2_X1 port map( A1 => n7645, A2 => n8221, ZN => n7648);
   U6267 : XNOR2_X1 port map( A => n16885, B => n16331, ZN => n16332);
   U6268 : NOR2_X1 port map( A1 => n9371, A2 => n2066, ZN => n2065);
   U6269 : NAND2_X1 port map( A1 => n3500, A2 => n11480, ZN => n11487);
   U6270 : NAND3_X2 port map( A1 => n14158, A2 => n2047, A3 => n3815, ZN => 
                           n14159);
   U6271 : NAND2_X1 port map( A1 => n14248, A2 => n20513, ZN => n2047);
   U6272 : NAND3_X2 port map( A1 => n7596, A2 => n7597, A3 => n7595, ZN => 
                           n8937);
   U6273 : OAI21_X1 port map( B1 => n5996, B2 => n6000, A => n5995, ZN => n2048
                           );
   U6274 : NAND2_X1 port map( A1 => n216, A2 => n3030, ZN => n2049);
   U6275 : NAND2_X1 port map( A1 => n5704, A2 => n5434, ZN => n2051);
   U6276 : NAND2_X1 port map( A1 => n2053, A2 => n1591, ZN => n2052);
   U6277 : NAND2_X1 port map( A1 => n12056, A2 => n12619, ZN => n2054);
   U6278 : NAND2_X1 port map( A1 => n11880, A2 => n11460, ZN => n11879);
   U6279 : XNOR2_X2 port map( A => n10218, B => n10217, ZN => n11880);
   U6280 : NOR2_X1 port map( A1 => n12201, A2 => n12594, ZN => n2056);
   U6281 : NAND2_X1 port map( A1 => n2059, A2 => n2057, ZN => n19006);
   U6282 : NAND2_X1 port map( A1 => n19724, A2 => n2058, ZN => n2057);
   U6283 : NAND2_X1 port map( A1 => n18999, A2 => n19013, ZN => n2059);
   U6284 : NAND2_X1 port map( A1 => n14490, A2 => n20453, ZN => n13877);
   U6285 : NAND2_X1 port map( A1 => n11206, A2 => n11094, ZN => n2060);
   U6286 : NAND2_X1 port map( A1 => n10846, A2 => n11203, ZN => n2061);
   U6288 : NAND2_X1 port map( A1 => n18940, A2 => n18936, ZN => n18933);
   U6290 : NAND3_X1 port map( A1 => n11327, A2 => n11255, A3 => n19886, ZN => 
                           n10309);
   U6292 : OAI211_X2 port map( C1 => n12875, C2 => n20502, A => n2069, B => 
                           n2068, ZN => n17411);
   U6293 : NAND2_X1 port map( A1 => n12874, A2 => n19888, ZN => n2068);
   U6294 : NAND2_X1 port map( A1 => n3979, A2 => n3978, ZN => n2070);
   U6295 : NAND2_X1 port map( A1 => n4420, A2 => n4220, ZN => n3979);
   U6296 : INV_X1 port map( A => n3978, ZN => n2071);
   U6297 : INV_X1 port map( A => n12544, ZN => n12305);
   U6298 : NAND2_X1 port map( A1 => n4866, A2 => n4865, ZN => n2072);
   U6300 : AOI22_X1 port map( A1 => n11405, A2 => n11404, B1 => n11406, B2 => 
                           n19506, ZN => n2810);
   U6301 : NAND2_X1 port map( A1 => n8583, A2 => n9298, ZN => n2073);
   U6302 : NAND2_X1 port map( A1 => n8584, A2 => n8846, ZN => n2074);
   U6303 : XNOR2_X2 port map( A => n16056, B => n16055, ZN => n17876);
   U6304 : OAI21_X1 port map( B1 => n988, B2 => n2075, A => n18597, ZN => 
                           n17626);
   U6305 : NOR2_X1 port map( A1 => n17624, A2 => n19656, ZN => n2075);
   U6306 : INV_X1 port map( A => n3588, ZN => n11403);
   U6307 : NAND3_X1 port map( A1 => n4146, A2 => n4645, A3 => n4325, ZN => 
                           n2076);
   U6308 : NAND2_X1 port map( A1 => n4016, A2 => n4642, ZN => n2077);
   U6310 : OR2_X1 port map( A1 => n3634, A2 => n3551, ZN => n3550);
   U6311 : INV_X1 port map( A => n8074, ZN => n3703);
   U6312 : INV_X1 port map( A => n4638, ZN => n2919);
   U6313 : INV_X1 port map( A => Plaintext(143), ZN => n3153);
   U6314 : INV_X1 port map( A => n18774, ZN => n18749);
   U6315 : XOR2_X1 port map( A => n10552, B => n1969, Z => n3424);
   U6316 : AOI22_X1 port map( A1 => n4276, A2 => n5018, B1 => n5014, B2 => 
                           n4111, ZN => n5276);
   U6317 : XNOR2_X1 port map( A => n9605, B => n10549, ZN => n2570);
   U6318 : XNOR2_X1 port map( A => n4247, B => n4246, ZN => n8060);
   U6319 : XNOR2_X1 port map( A => n13533, B => n2078, ZN => n13140);
   U6320 : XNOR2_X1 port map( A => n13137, B => n13616, ZN => n2078);
   U6322 : NAND2_X1 port map( A1 => n19590, A2 => n9564, ZN => n8703);
   U6323 : OR2_X2 port map( A1 => n14459, A2 => n14458, ZN => n15295);
   U6324 : NAND2_X1 port map( A1 => n2441, A2 => n8384, ZN => n8135);
   U6325 : NAND2_X1 port map( A1 => n7684, A2 => n8380, ZN => n8384);
   U6326 : NAND2_X1 port map( A1 => n2081, A2 => n2080, ZN => n5561);
   U6327 : NAND2_X1 port map( A1 => n5557, A2 => n6048, ZN => n2080);
   U6329 : NAND2_X1 port map( A1 => n5010, A2 => n4204, ZN => n4206);
   U6330 : NOR2_X1 port map( A1 => n14768, A2 => n15107, ZN => n14771);
   U6331 : AOI22_X1 port map( A1 => n17581, A2 => n20433, B1 => n17582, B2 => 
                           n19773, ZN => n17583);
   U6332 : AOI21_X1 port map( B1 => n20618, B2 => n12147, A => n3666, ZN => 
                           n12314);
   U6333 : OAI211_X1 port map( C1 => n14678, C2 => n20120, A => n14279, B => 
                           n14677, ZN => n14683);
   U6334 : NAND3_X1 port map( A1 => n19752, A2 => n15421, A3 => n15420, ZN => 
                           n15083);
   U6335 : NAND2_X1 port map( A1 => n12369, A2 => n12374, ZN => n11856);
   U6336 : NAND2_X1 port map( A1 => n893, A2 => n300, ZN => n2084);
   U6337 : NAND2_X1 port map( A1 => n17737, A2 => n18501, ZN => n17739);
   U6339 : NAND3_X1 port map( A1 => n14210, A2 => n2086, A3 => n2085, ZN => 
                           n15070);
   U6340 : NAND2_X1 port map( A1 => n14207, A2 => n14206, ZN => n2085);
   U6341 : NAND2_X1 port map( A1 => n14209, A2 => n14208, ZN => n2086);
   U6344 : OAI22_X1 port map( A1 => n15500, A2 => n15502, B1 => n15192, B2 => 
                           n15496, ZN => n14042);
   U6345 : AND3_X2 port map( A1 => n2088, A2 => n3173, A3 => n3172, ZN => 
                           n15500);
   U6347 : NAND2_X1 port map( A1 => n7890, A2 => n8190, ZN => n2089);
   U6349 : OR2_X1 port map( A1 => n4094, A2 => n4268, ZN => n4582);
   U6350 : NAND2_X1 port map( A1 => n2093, A2 => n2091, ZN => n4436);
   U6351 : NAND2_X1 port map( A1 => n2092, A2 => n6124, ZN => n2091);
   U6352 : OR2_X1 port map( A1 => n19921, A2 => n14690, ZN => n2094);
   U6355 : XNOR2_X1 port map( A => n13850, B => n13851, ZN => n2095);
   U6357 : NAND3_X1 port map( A1 => n1041, A2 => n9234, A3 => n2097, ZN => 
                           n3059);
   U6358 : NAND2_X1 port map( A1 => n2254, A2 => n2255, ZN => n12644);
   U6359 : XNOR2_X1 port map( A => n13078, B => n19904, ZN => n2200);
   U6360 : XNOR2_X1 port map( A => n13154, B => n13027, ZN => n13078);
   U6361 : NAND2_X1 port map( A1 => n16319, A2 => n2945, ZN => n2127);
   U6362 : NAND2_X1 port map( A1 => n12483, A2 => n12472, ZN => n2552);
   U6363 : XNOR2_X2 port map( A => n15988, B => n15987, ZN => n17676);
   U6364 : AOI21_X1 port map( B1 => n15755, B2 => n2247, A => n2101, ZN => 
                           n2374);
   U6366 : NAND2_X1 port map( A1 => n15760, A2 => n15754, ZN => n2102);
   U6367 : OAI21_X1 port map( B1 => n11363, B2 => n19952, A => n2104, ZN => 
                           n11372);
   U6368 : NAND2_X1 port map( A1 => n15131, A2 => n15285, ZN => n2105);
   U6369 : NAND2_X1 port map( A1 => n8195, A2 => n8055, ZN => n8194);
   U6372 : XNOR2_X1 port map( A => n13052, B => n13051, ZN => n14497);
   U6373 : OR2_X1 port map( A1 => n9081, A2 => n9166, ZN => n2941);
   U6374 : INV_X1 port map( A => n4706, ZN => n3203);
   U6375 : INV_X1 port map( A => Plaintext(124), ZN => n3204);
   U6376 : NOR2_X1 port map( A1 => n11051, A2 => n10829, ZN => n2162);
   U6377 : NOR2_X1 port map( A1 => n15303, A2 => n15302, ZN => n2581);
   U6378 : XNOR2_X1 port map( A => n10351, B => n9908, ZN => n10395);
   U6379 : XNOR2_X1 port map( A => n16555, B => n16236, ZN => n16871);
   U6380 : XNOR2_X1 port map( A => n6410, B => n7288, ZN => n6864);
   U6381 : NAND3_X1 port map( A1 => n5770, A2 => n5766, A3 => n5546, ZN => 
                           n5738);
   U6383 : NAND2_X1 port map( A1 => n2267, A2 => n15338, ZN => n2109);
   U6386 : AOI22_X1 port map( A1 => n20117, A2 => n18850, B1 => n19989, B2 => 
                           n18869, ZN => n18871);
   U6387 : XNOR2_X1 port map( A => n10247, B => n10248, ZN => n10251);
   U6388 : NAND2_X1 port map( A1 => n15039, A2 => n15141, ZN => n2111);
   U6389 : NAND2_X1 port map( A1 => n2113, A2 => n2112, ZN => n14858);
   U6390 : NAND2_X1 port map( A1 => n14857, A2 => n15766, ZN => n2112);
   U6391 : NAND2_X1 port map( A1 => n11155, A2 => n11159, ZN => n2970);
   U6394 : NAND2_X1 port map( A1 => n19710, A2 => n9262, ZN => n2116);
   U6395 : INV_X1 port map( A => n9262, ZN => n2118);
   U6398 : INV_X1 port map( A => n18025, ZN => n2120);
   U6399 : NAND2_X1 port map( A1 => n6143, A2 => n6140, ZN => n4462);
   U6400 : NAND2_X1 port map( A1 => n11718, A2 => n12282, ZN => n2121);
   U6401 : NAND2_X1 port map( A1 => n8071, A2 => n5762, ZN => n8202);
   U6402 : NAND2_X1 port map( A1 => n15664, A2 => n15773, ZN => n15670);
   U6404 : XNOR2_X1 port map( A => n17127, B => n2280, ZN => n15951);
   U6406 : OAI21_X1 port map( B1 => n12392, B2 => n3082, A => n12391, ZN => 
                           n12831);
   U6407 : NAND2_X1 port map( A1 => n4927, A2 => n4932, ZN => n4930);
   U6408 : OAI21_X1 port map( B1 => n13977, B2 => n14284, A => n2125, ZN => 
                           n13978);
   U6409 : NAND3_X1 port map( A1 => n5605, A2 => n5604, A3 => n5714, ZN => 
                           n5607);
   U6410 : OAI21_X1 port map( B1 => n8288, B2 => n7807, A => n2126, ZN => n7400
                           );
   U6411 : NAND2_X1 port map( A1 => n7807, A2 => n8289, ZN => n2126);
   U6412 : OR3_X1 port map( A1 => n8998, A2 => n8997, A3 => n7752, ZN => n7774)
                           ;
   U6413 : XNOR2_X2 port map( A => n3875, B => Key(18), ZN => n4296);
   U6414 : AND2_X1 port map( A1 => n8760, A2 => n265, ZN => n8766);
   U6416 : OAI22_X1 port map( A1 => n17662, A2 => n20185, B1 => n3214, B2 => 
                           n17890, ZN => n3213);
   U6417 : OAI21_X1 port map( B1 => n9299, B2 => n3418, A => n2786, ZN => n3201
                           );
   U6418 : NAND2_X1 port map( A1 => n3652, A2 => n4418, ZN => n3651);
   U6419 : XNOR2_X1 port map( A => n2127, B => n2263, ZN => Ciphertext(152));
   U6420 : OAI21_X1 port map( B1 => n9172, B2 => n8617, A => n8619, ZN => n7806
                           );
   U6422 : NAND3_X1 port map( A1 => n15411, A2 => n15551, A3 => n2129, ZN => 
                           n16050);
   U6423 : NAND2_X1 port map( A1 => n20147, A2 => n15056, ZN => n15411);
   U6424 : NAND2_X1 port map( A1 => n256, A2 => n12179, ZN => n9498);
   U6426 : NOR3_X1 port map( A1 => n12267, A2 => n3734, A3 => n12562, ZN => 
                           n11062);
   U6428 : NAND2_X1 port map( A1 => n2133, A2 => n2132, ZN => n10316);
   U6429 : NAND2_X1 port map( A1 => n12337, A2 => n12336, ZN => n2132);
   U6430 : NAND2_X1 port map( A1 => n11974, A2 => n12334, ZN => n2133);
   U6431 : NOR2_X1 port map( A1 => n2135, A2 => n2134, ZN => n11498);
   U6432 : NAND2_X1 port map( A1 => n2137, A2 => n2136, ZN => n6711);
   U6433 : NAND2_X1 port map( A1 => n5707, A2 => n6002, ZN => n2137);
   U6434 : NAND2_X1 port map( A1 => n3319, A2 => n5880, ZN => n5153);
   U6435 : NAND2_X1 port map( A1 => n19329, A2 => n19324, ZN => n19310);
   U6436 : NAND2_X1 port map( A1 => n12632, A2 => n246, ZN => n2139);
   U6437 : NAND2_X1 port map( A1 => n11618, A2 => n1371, ZN => n2140);
   U6438 : AND3_X2 port map( A1 => n8043, A2 => n2142, A3 => n2141, ZN => n8542
                           );
   U6439 : NAND2_X1 port map( A1 => n8296, A2 => n8300, ZN => n2141);
   U6440 : NAND2_X1 port map( A1 => n8042, A2 => n1835, ZN => n2142);
   U6442 : OR2_X1 port map( A1 => n5781, A2 => n6046, ZN => n2144);
   U6444 : AOI22_X1 port map( A1 => n12072, A2 => n12609, B1 => n12606, B2 => 
                           n12073, ZN => n12076);
   U6445 : XNOR2_X1 port map( A => n929, B => n10369, ZN => n2145);
   U6446 : MUX2_X1 port map( A => n5880, B => n5881, S => n3319, Z => n5882);
   U6447 : OAI21_X2 port map( B1 => n12026, B2 => n12377, A => n12025, ZN => 
                           n13369);
   U6449 : NAND2_X1 port map( A1 => n891, A2 => n9300, ZN => n8584);
   U6451 : NAND2_X1 port map( A1 => n14609, A2 => n14608, ZN => n3226);
   U6452 : NAND2_X1 port map( A1 => n15862, A2 => n15864, ZN => n15860);
   U6453 : NAND2_X1 port map( A1 => n12477, A2 => n12142, ZN => n2148);
   U6454 : AND2_X1 port map( A1 => n14203, A2 => n14012, ZN => n14143);
   U6456 : INV_X1 port map( A => n12542, ZN => n2600);
   U6457 : OR2_X1 port map( A1 => n20357, A2 => n4867, ZN => n4227);
   U6459 : NAND2_X1 port map( A1 => n11569, A2 => n11564, ZN => n2949);
   U6460 : OAI21_X1 port map( B1 => n14159, B2 => n15509, A => n2908, ZN => 
                           n15514);
   U6461 : OAI22_X1 port map( A1 => n8665, A2 => n9204, B1 => n20009, B2 => 
                           n9130, ZN => n9779);
   U6464 : NAND2_X1 port map( A1 => n6041, A2 => n5888, ZN => n2149);
   U6465 : NAND2_X1 port map( A1 => n14649, A2 => n19831, ZN => n2153);
   U6466 : NAND2_X1 port map( A1 => n2154, A2 => n8904, ZN => n8592);
   U6467 : NAND2_X1 port map( A1 => n2756, A2 => n19941, ZN => n2154);
   U6468 : NAND2_X1 port map( A1 => n5865, A2 => n2157, ZN => n6786);
   U6469 : NAND2_X1 port map( A1 => n2158, A2 => n5864, ZN => n2157);
   U6470 : OAI22_X1 port map( A1 => n20464, A2 => n4440, B1 => n5040, B2 => 
                           n4439, ZN => n4441);
   U6471 : NOR2_X1 port map( A1 => n9883, A2 => n11234, ZN => n11367);
   U6473 : NAND2_X1 port map( A1 => n12685, A2 => n12684, ZN => n12687);
   U6474 : AOI21_X1 port map( B1 => n5510, B2 => n5070, A => n5071, ZN => n4665
                           );
   U6475 : NAND2_X1 port map( A1 => n5069, A2 => n4410, ZN => n5510);
   U6476 : NAND2_X1 port map( A1 => n12307, A2 => n12543, ZN => n2159);
   U6477 : OAI21_X1 port map( B1 => n11418, B2 => n11417, A => n2161, ZN => 
                           n10725);
   U6479 : OAI21_X2 port map( B1 => n6203, B2 => n5230, A => n5229, ZN => n7249
                           );
   U6482 : NAND2_X1 port map( A1 => n2236, A2 => n2237, ZN => n18157);
   U6483 : XNOR2_X1 port map( A => n2163, B => n16131, ZN => n16133);
   U6484 : XNOR2_X1 port map( A => n16130, B => n16988, ZN => n2163);
   U6485 : NAND2_X1 port map( A1 => n8032, A2 => n8284, ZN => n2166);
   U6486 : OAI21_X1 port map( B1 => n6139, B2 => n5866, A => n5265, ZN => n5267
                           );
   U6488 : OR2_X1 port map( A1 => n6951, A2 => n8365, ZN => n7676);
   U6489 : OR2_X1 port map( A1 => n11477, A2 => n3482, ZN => n3480);
   U6490 : INV_X1 port map( A => n11311, ZN => n2759);
   U6492 : NAND2_X1 port map( A1 => n2698, A2 => n2167, ZN => n2723);
   U6493 : NAND2_X1 port map( A1 => n2171, A2 => n2168, ZN => n9570);
   U6494 : NAND2_X1 port map( A1 => n9564, A2 => n9563, ZN => n2169);
   U6495 : OR2_X1 port map( A1 => n20105, A2 => n3978, ZN => n4658);
   U6496 : AND2_X1 port map( A1 => n20235, A2 => n11292, ZN => n10979);
   U6497 : INV_X1 port map( A => n3741, ZN => n3103);
   U6498 : XNOR2_X1 port map( A => n17380, B => n2172, ZN => n17381);
   U6499 : XNOR2_X1 port map( A => n17377, B => n17378, ZN => n2172);
   U6501 : XNOR2_X1 port map( A => n10604, B => n2349, ZN => n10606);
   U6502 : AND2_X1 port map( A1 => n8653, A2 => n9265, ZN => n7867);
   U6504 : INV_X1 port map( A => n5815, ZN => n3468);
   U6505 : XNOR2_X1 port map( A => n941, B => n7296, ZN => n7064);
   U6506 : OR2_X1 port map( A1 => n17773, A2 => n18333, ZN => n2177);
   U6507 : OAI21_X1 port map( B1 => n5419, B2 => n5226, A => n5418, ZN => n2404
                           );
   U6508 : XNOR2_X1 port map( A => n16566, B => n17276, ZN => n16091);
   U6511 : NAND2_X1 port map( A1 => n2179, A2 => n2178, ZN => n18798);
   U6512 : NAND2_X1 port map( A1 => n18796, A2 => n18795, ZN => n2178);
   U6514 : INV_X1 port map( A => n18814, ZN => n18811);
   U6515 : NAND2_X1 port map( A1 => n2182, A2 => n2180, ZN => n17058);
   U6516 : NAND2_X1 port map( A1 => n18916, A2 => n2181, ZN => n2180);
   U6517 : NOR2_X1 port map( A1 => n18921, A2 => n18899, ZN => n2181);
   U6518 : NAND2_X1 port map( A1 => n18874, A2 => n19874, ZN => n2182);
   U6522 : INV_X1 port map( A => n17303, ZN => n3205);
   U6523 : OR2_X1 port map( A1 => n11954, A2 => n11951, ZN => n11956);
   U6524 : NOR2_X1 port map( A1 => n3839, A2 => n5782, ZN => n3249);
   U6525 : NOR2_X1 port map( A1 => n3671, A2 => n11145, ZN => n3670);
   U6526 : AND2_X1 port map( A1 => n14465, A2 => n14462, ZN => n14176);
   U6527 : INV_X1 port map( A => n9164, ZN => n8609);
   U6528 : XNOR2_X1 port map( A => n2312, B => n13624, ZN => n13533);
   U6529 : OAI21_X1 port map( B1 => n9158, B2 => n8696, A => n8610, ZN => n8614
                           );
   U6530 : XNOR2_X1 port map( A => n5884, B => n7118, ZN => n6659);
   U6531 : NAND2_X1 port map( A1 => n12565, A2 => n2183, ZN => n12566);
   U6532 : NAND3_X2 port map( A1 => n3536, A2 => n2185, A3 => n2184, ZN => 
                           n13715);
   U6533 : NAND2_X1 port map( A1 => n2737, A2 => n12002, ZN => n2185);
   U6534 : OAI211_X2 port map( C1 => n14696, C2 => n14695, A => n14694, B => 
                           n2186, ZN => n15567);
   U6535 : NAND3_X1 port map( A1 => n2187, A2 => n11639, A3 => n12209, ZN => 
                           n2714);
   U6536 : NAND2_X1 port map( A1 => n12067, A2 => n12206, ZN => n2187);
   U6537 : NAND2_X1 port map( A1 => n9276, A2 => n8991, ZN => n7897);
   U6538 : NAND2_X1 port map( A1 => n11939, A2 => n12110, ZN => n12099);
   U6540 : NAND2_X1 port map( A1 => n8083, A2 => n8232, ZN => n2188);
   U6542 : NAND2_X1 port map( A1 => n6584, A2 => n6585, ZN => n2191);
   U6543 : NOR2_X1 port map( A1 => n4185, A2 => n4633, ZN => n4159);
   U6544 : AOI22_X1 port map( A1 => n15372, A2 => n15567, B1 => n15564, B2 => 
                           n20183, ZN => n15373);
   U6545 : OAI211_X1 port map( C1 => n11329, C2 => n2858, A => n2861, B => 
                           n2857, ZN => n2856);
   U6546 : NAND2_X1 port map( A1 => n3393, A2 => n3457, ZN => n3392);
   U6548 : INV_X1 port map( A => n19113, ZN => n2195);
   U6550 : INV_X1 port map( A => n17533, ZN => n2197);
   U6551 : NAND2_X1 port map( A1 => n4771, A2 => n5035, ZN => n5038);
   U6552 : INV_X1 port map( A => n19386, ZN => n17220);
   U6553 : INV_X1 port map( A => n8167, ZN => n3121);
   U6554 : NAND3_X1 port map( A1 => n19789, A2 => n5926, A3 => n6026, ZN => 
                           n2342);
   U6556 : INV_X1 port map( A => n7750, ZN => n3446);
   U6557 : XNOR2_X1 port map( A => n2199, B => n10588, ZN => n9428);
   U6558 : XNOR2_X1 port map( A => n3184, B => n10430, ZN => n2199);
   U6559 : NAND2_X1 port map( A1 => n3632, A2 => n11599, ZN => n3631);
   U6561 : NAND2_X1 port map( A1 => n1527, A2 => n2201, ZN => n14234);
   U6563 : OAI211_X2 port map( C1 => n5669, C2 => n4880, A => n5677, B => n4879
                           , ZN => n7337);
   U6565 : AND2_X1 port map( A1 => n14556, A2 => n14553, ZN => n14551);
   U6567 : NAND2_X1 port map( A1 => n4588, A2 => n4585, ZN => n5054);
   U6569 : OAI21_X1 port map( B1 => n11421, B2 => n11420, A => n11422, ZN => 
                           n2440);
   U6570 : NAND2_X1 port map( A1 => n2205, A2 => n2204, ZN => n17056);
   U6571 : NAND2_X1 port map( A1 => n19684, A2 => n18961, ZN => n2204);
   U6572 : NAND2_X1 port map( A1 => n17055, A2 => n220, ZN => n2205);
   U6573 : NAND2_X1 port map( A1 => n16674, A2 => n19352, ZN => n2206);
   U6574 : OAI21_X1 port map( B1 => n4368, B2 => n5240, A => n5720, ZN => n2207
                           );
   U6575 : NOR2_X2 port map( A1 => n11068, A2 => n11067, ZN => n13319);
   U6577 : OR2_X2 port map( A1 => n10812, A2 => n10811, ZN => n12211);
   U6579 : NAND2_X1 port map( A1 => n2209, A2 => n11570, ZN => n10752);
   U6580 : NAND2_X1 port map( A1 => n10751, A2 => n2210, ZN => n2209);
   U6581 : INV_X1 port map( A => n11568, ZN => n2210);
   U6582 : XNOR2_X1 port map( A => n6771, B => n6770, ZN => n2211);
   U6583 : NAND2_X1 port map( A1 => n2213, A2 => n2212, ZN => n15359);
   U6584 : NAND2_X1 port map( A1 => n15357, A2 => n15815, ZN => n2212);
   U6585 : NAND2_X1 port map( A1 => n15358, A2 => n3534, ZN => n2213);
   U6589 : NAND2_X1 port map( A1 => n5032, A2 => n4706, ZN => n4709);
   U6591 : NAND2_X1 port map( A1 => n8282, A2 => n8286, ZN => n2217);
   U6593 : XNOR2_X1 port map( A => n13031, B => n12986, ZN => n13733);
   U6594 : INV_X1 port map( A => n18046, ZN => n2586);
   U6595 : INV_X1 port map( A => n5087, ZN => n4801);
   U6596 : OR2_X1 port map( A1 => n4979, A2 => n4296, ZN => n4020);
   U6597 : INV_X1 port map( A => n3305, ZN => n12610);
   U6598 : INV_X1 port map( A => n15295, ZN => n3307);
   U6599 : INV_X1 port map( A => n10926, ZN => n11545);
   U6600 : XNOR2_X1 port map( A => n13707, B => n13002, ZN => n3460);
   U6601 : OAI21_X1 port map( B1 => n5972, B2 => n5971, A => n5970, ZN => n5975
                           );
   U6602 : NAND2_X1 port map( A1 => n5967, A2 => n5697, ZN => n5970);
   U6604 : XNOR2_X1 port map( A => n2224, B => n16518, ZN => n16520);
   U6605 : XNOR2_X1 port map( A => n16602, B => n16517, ZN => n2224);
   U6606 : NAND2_X1 port map( A1 => n8193, A2 => n8197, ZN => n7627);
   U6608 : NAND2_X1 port map( A1 => n18165, A2 => n19292, ZN => n2226);
   U6609 : XNOR2_X1 port map( A => n9946, B => n10071, ZN => n10621);
   U6611 : XNOR2_X1 port map( A => n13513, B => n2228, ZN => n13515);
   U6612 : XNOR2_X1 port map( A => n13514, B => n13512, ZN => n2228);
   U6613 : OAI21_X1 port map( B1 => n10854, B2 => n11230, A => n2229, ZN => 
                           n11233);
   U6614 : NAND2_X1 port map( A1 => n11230, A2 => n11365, ZN => n2229);
   U6615 : XNOR2_X1 port map( A => n2230, B => n13852, ZN => n12249);
   U6616 : XNOR2_X1 port map( A => n13757, B => n12219, ZN => n2230);
   U6617 : INV_X1 port map( A => n873, ZN => n2929);
   U6618 : XNOR2_X2 port map( A => n12783, B => n12782, ZN => n13931);
   U6619 : INV_X1 port map( A => n11176, ZN => n2232);
   U6620 : NAND2_X1 port map( A1 => n10997, A2 => n11289, ZN => n2235);
   U6621 : INV_X1 port map( A => Plaintext(53), ZN => n3543);
   U6624 : OAI21_X1 port map( B1 => n16152, B2 => n20423, A => n16151, ZN => 
                           n2237);
   U6625 : NAND2_X1 port map( A1 => n4545, A2 => n2239, ZN => n4551);
   U6627 : NAND3_X1 port map( A1 => n3710, A2 => n15921, A3 => n15421, ZN => 
                           n14899);
   U6628 : NOR2_X1 port map( A1 => n12212, A2 => n12211, ZN => n2743);
   U6630 : NAND2_X1 port map( A1 => n10854, A2 => n11230, ZN => n9884);
   U6631 : NAND2_X1 port map( A1 => n8618, A2 => n8987, ZN => n2241);
   U6632 : INV_X1 port map( A => n8987, ZN => n2243);
   U6633 : NAND3_X2 port map( A1 => n14628, A2 => n14621, A3 => n14622, ZN => 
                           n15600);
   U6635 : MUX2_X1 port map( A => n8525, B => n8526, S => n9038, Z => n8531);
   U6636 : NAND2_X1 port map( A1 => n15761, A2 => n2247, ZN => n2246);
   U6637 : INV_X1 port map( A => n15760, ZN => n2247);
   U6638 : NAND2_X2 port map( A1 => n3165, A2 => n4794, ZN => n5663);
   U6639 : NAND2_X1 port map( A1 => n12443, A2 => n12440, ZN => n12435);
   U6640 : NAND3_X1 port map( A1 => n20261, A2 => n2697, A3 => n14828, ZN => 
                           n2696);
   U6641 : NOR2_X1 port map( A1 => n7311, A2 => n7312, ZN => n7998);
   U6642 : NAND2_X1 port map( A1 => n210, A2 => n2596, ZN => n2576);
   U6643 : XNOR2_X1 port map( A => n2250, B => n13470, ZN => n13473);
   U6644 : XNOR2_X1 port map( A => n13469, B => n13818, ZN => n2250);
   U6646 : NAND2_X1 port map( A1 => n7905, A2 => n280, ZN => n2252);
   U6647 : AOI21_X1 port map( B1 => n2253, B2 => n4509, A => n4371, ZN => n4374
                           );
   U6648 : NAND2_X1 port map( A1 => n4372, A2 => n4577, ZN => n2253);
   U6649 : INV_X1 port map( A => n15188, ZN => n13933);
   U6650 : XOR2_X1 port map( A => n13778, B => n13059, Z => n2620);
   U6651 : NAND2_X1 port map( A1 => n12637, A2 => n19861, ZN => n2254);
   U6652 : NAND2_X1 port map( A1 => n12638, A2 => n2256, ZN => n2255);
   U6653 : MUX2_X2 port map( A => n10807, B => n10806, S => n11257, Z => n12209
                           );
   U6654 : XNOR2_X2 port map( A => n12764, B => n12763, ZN => n14827);
   U6655 : NAND2_X1 port map( A1 => n2688, A2 => n2703, ZN => n2702);
   U6656 : INV_X1 port map( A => n15052, ZN => n15458);
   U6657 : INV_X1 port map( A => n8993, ZN => n9278);
   U6658 : NAND2_X1 port map( A1 => n13961, A2 => n14924, ZN => n13970);
   U6659 : NAND2_X1 port map( A1 => n6905, A2 => n7909, ZN => n2258);
   U6661 : NAND2_X1 port map( A1 => n19268, A2 => n19267, ZN => n2261);
   U6662 : NAND2_X1 port map( A1 => n19266, A2 => n20444, ZN => n2262);
   U6663 : INV_X1 port map( A => n18354, ZN => n18289);
   U6664 : NOR2_X2 port map( A1 => n6898, A2 => n6897, ZN => n10252);
   U6665 : INV_X1 port map( A => n6107, ZN => n3010);
   U6666 : OAI21_X1 port map( B1 => n11931, B2 => n12480, A => n2265, ZN => 
                           n11708);
   U6667 : NAND2_X1 port map( A1 => n12478, A2 => n12142, ZN => n2265);
   U6668 : NAND4_X2 port map( A1 => n2266, A2 => n3132, A3 => n5062, A4 => 
                           n5061, ZN => n5930);
   U6669 : OAI21_X1 port map( B1 => n13166, B2 => n14664, A => n3367, ZN => 
                           n14671);
   U6671 : NAND2_X1 port map( A1 => n15337, A2 => n15336, ZN => n2267);
   U6672 : NAND3_X1 port map( A1 => n14130, A2 => n14129, A3 => n14128, ZN => 
                           n15607);
   U6674 : INV_X1 port map( A => n2269, ZN => n2268);
   U6675 : OAI22_X1 port map( A1 => n17832, A2 => n17831, B1 => n17833, B2 => 
                           n18959, ZN => n2269);
   U6676 : NAND2_X1 port map( A1 => n11441, A2 => n11440, ZN => n2270);
   U6677 : NAND2_X1 port map( A1 => n11442, A2 => n2272, ZN => n2271);
   U6678 : XNOR2_X2 port map( A => n3930, B => Key(164), ZN => n4347);
   U6679 : NOR2_X1 port map( A1 => n15664, A2 => n2273, ZN => n13460);
   U6680 : INV_X1 port map( A => n15772, ZN => n2273);
   U6681 : NOR2_X2 port map( A1 => n15398, A2 => n15399, ZN => n16761);
   U6682 : AOI21_X1 port map( B1 => n2761, B2 => n2760, A => n2759, ZN => n2758
                           );
   U6683 : NOR2_X1 port map( A1 => n209, A2 => n6068, ZN => n3767);
   U6684 : XNOR2_X1 port map( A => n10507, B => n2506, ZN => n10509);
   U6685 : NAND2_X1 port map( A1 => n4485, A2 => n3996, ZN => n4681);
   U6687 : XNOR2_X2 port map( A => n13728, B => n13729, ZN => n14381);
   U6688 : NOR2_X1 port map( A1 => n20611, A2 => n20361, ZN => n18381);
   U6689 : XNOR2_X1 port map( A => n13191, B => n12825, ZN => n2783);
   U6690 : AOI21_X1 port map( B1 => n2276, B2 => n14502, A => n13040, ZN => 
                           n13056);
   U6691 : NAND2_X1 port map( A1 => n9307, A2 => n9310, ZN => n8824);
   U6692 : NAND2_X1 port map( A1 => n2277, A2 => n20434, ZN => n17615);
   U6693 : INV_X1 port map( A => n19298, ZN => n2277);
   U6694 : AOI21_X2 port map( B1 => n17605, B2 => n17604, A => n17603, ZN => 
                           n19298);
   U6695 : NAND2_X1 port map( A1 => n5749, A2 => n5747, ZN => n2482);
   U6696 : AOI21_X1 port map( B1 => n11369, B2 => n10680, A => n11364, ZN => 
                           n10681);
   U6698 : NOR2_X2 port map( A1 => n7652, A2 => n7651, ZN => n10566);
   U6700 : NAND2_X1 port map( A1 => n5546, A2 => n5736, ZN => n4545);
   U6702 : NAND2_X1 port map( A1 => n15453, A2 => n15683, ZN => n2279);
   U6705 : NAND3_X1 port map( A1 => n4151, A2 => n4312, A3 => n4361, ZN => 
                           n4155);
   U6708 : NAND2_X1 port map( A1 => n13308, A2 => n2282, ZN => n2281);
   U6709 : OAI211_X2 port map( C1 => n7470, C2 => n8031, A => n2283, B => n8030
                           , ZN => n9060);
   U6710 : NAND2_X1 port map( A1 => n8028, A2 => n8029, ZN => n2283);
   U6711 : XNOR2_X1 port map( A => n8509, B => n9445, ZN => n2285);
   U6712 : NAND2_X1 port map( A1 => n16730, A2 => n3755, ZN => n3283);
   U6713 : AOI21_X1 port map( B1 => n6070, B2 => n6072, A => n2286, ZN => n6074
                           );
   U6714 : BUF_X1 port map( A => n3843, Z => n4676);
   U6715 : OAI211_X1 port map( C1 => n5072, C2 => n5071, A => n4816, B => n2287
                           , ZN => n4818);
   U6716 : AND3_X2 port map( A1 => n3650, A2 => n3651, A3 => n4419, ZN => n5868
                           );
   U6717 : XNOR2_X2 port map( A => n16124, B => n16125, ZN => n17840);
   U6718 : INV_X1 port map( A => n15188, ZN => n2288);
   U6719 : INV_X1 port map( A => n2561, ZN => n3385);
   U6720 : XNOR2_X1 port map( A => n3620, B => n7381, ZN => n7388);
   U6721 : MUX2_X1 port map( A => n12532, B => n12534, S => n12162, Z => n11807
                           );
   U6722 : INV_X1 port map( A => n15660, ZN => n15653);
   U6723 : NAND2_X1 port map( A1 => n17774, A2 => n17777, ZN => n2289);
   U6724 : NAND2_X1 port map( A1 => n17449, A2 => n18129, ZN => n2290);
   U6725 : NAND2_X1 port map( A1 => n2292, A2 => n6075, ZN => n2291);
   U6726 : NAND2_X1 port map( A1 => n3318, A2 => n209, ZN => n2292);
   U6727 : NOR2_X2 port map( A1 => n8487, A2 => n8486, ZN => n10402);
   U6728 : NAND2_X1 port map( A1 => n3995, A2 => n4684, ZN => n4226);
   U6729 : NAND2_X1 port map( A1 => n15078, A2 => n15077, ZN => n14371);
   U6731 : NAND2_X1 port map( A1 => n2919, A2 => n20487, ZN => n3634);
   U6733 : INV_X1 port map( A => n15465, ZN => n12768);
   U6734 : OAI211_X2 port map( C1 => n12726, C2 => n12727, A => n13924, B => 
                           n3190, ZN => n15465);
   U6736 : OAI21_X1 port map( B1 => n16461, B2 => n17479, A => n960, ZN => 
                           n2297);
   U6738 : OAI21_X1 port map( B1 => n5717, B2 => n5716, A => n5718, ZN => n3664
                           );
   U6739 : OR2_X1 port map( A1 => n3995, A2 => n3996, ZN => n4851);
   U6742 : XNOR2_X2 port map( A => Key(75), B => Plaintext(75), ZN => n4824);
   U6743 : XNOR2_X1 port map( A => n6982, B => n7050, ZN => n6328);
   U6744 : NAND3_X1 port map( A1 => n619, A2 => n4612, A3 => n3716, ZN => n3714
                           );
   U6747 : OAI21_X2 port map( B1 => n9063, B2 => n9036, A => n9035, ZN => n9991
                           );
   U6748 : NAND3_X2 port map( A1 => n11308, A2 => n11309, A3 => n11307, ZN => 
                           n12809);
   U6749 : OAI21_X1 port map( B1 => n17601, B2 => n17890, A => n2302, ZN => 
                           n17889);
   U6750 : NAND2_X1 port map( A1 => n20019, A2 => n17890, ZN => n2302);
   U6751 : AOI21_X1 port map( B1 => n7853, B2 => n7854, A => n7852, ZN => n2303
                           );
   U6752 : NAND2_X1 port map( A1 => n9029, A2 => n9062, ZN => n8677);
   U6753 : INV_X1 port map( A => n2800, ZN => n15073);
   U6755 : INV_X1 port map( A => n4615, ZN => n3717);
   U6756 : OAI211_X2 port map( C1 => n15797, C2 => n15796, A => n2309, B => 
                           n2308, ZN => n17426);
   U6757 : NAND2_X1 port map( A1 => n15793, A2 => n15796, ZN => n2308);
   U6758 : NAND2_X1 port map( A1 => n16810, A2 => n18546, ZN => n18532);
   U6759 : NAND2_X1 port map( A1 => n13274, A2 => n12324, ZN => n12329);
   U6760 : NAND2_X1 port map( A1 => n12322, A2 => n12323, ZN => n13274);
   U6761 : NAND2_X1 port map( A1 => n13859, A2 => n15443, ZN => n2311);
   U6763 : OAI21_X1 port map( B1 => n14601, B2 => n19918, A => n1262, ZN => 
                           n2314);
   U6764 : NAND2_X1 port map( A1 => n9491, A2 => n12180, ZN => n11845);
   U6767 : OAI21_X1 port map( B1 => n2316, B2 => n14833, A => n14828, ZN => 
                           n12767);
   U6768 : NAND4_X2 port map( A1 => n5162, A2 => n5161, A3 => n5160, A4 => 
                           n5159, ZN => n7365);
   U6769 : INV_X1 port map( A => n2955, ZN => n7610);
   U6770 : OR2_X1 port map( A1 => n14420, A2 => n14355, ZN => n14356);
   U6771 : AND2_X1 port map( A1 => n12315, A2 => n2612, ZN => n2338);
   U6773 : INV_X1 port map( A => n14461, ZN => n15111);
   U6774 : NAND2_X1 port map( A1 => n16780, A2 => n870, ZN => n16779);
   U6775 : XNOR2_X1 port map( A => n2318, B => n16788, ZN => Ciphertext(135));
   U6776 : NAND3_X1 port map( A1 => n3139, A2 => n3142, A3 => n3143, ZN => 
                           n2318);
   U6777 : OAI21_X2 port map( B1 => n11037, B2 => n10523, A => n10522, ZN => 
                           n12514);
   U6778 : NAND3_X1 port map( A1 => n12243, A2 => n12619, A3 => n894, ZN => 
                           n12244);
   U6779 : NAND2_X1 port map( A1 => n14236, A2 => n14239, ZN => n14401);
   U6780 : NAND2_X1 port map( A1 => n3048, A2 => n3052, ZN => n2319);
   U6781 : NAND3_X1 port map( A1 => n4160, A2 => n4517, A3 => n4523, ZN => 
                           n4161);
   U6782 : NAND2_X1 port map( A1 => n12313, A2 => n12153, ZN => n2320);
   U6783 : NAND2_X1 port map( A1 => n3235, A2 => n18104, ZN => n18110);
   U6784 : AND3_X2 port map( A1 => n14152, A2 => n14151, A3 => n14150, ZN => 
                           n3822);
   U6785 : NAND3_X2 port map( A1 => n2322, A2 => n2321, A3 => n5290, ZN => 
                           n7006);
   U6786 : NAND3_X1 port map( A1 => n5289, A2 => n5291, A3 => n5443, ZN => 
                           n2322);
   U6787 : OR2_X2 port map( A1 => n4408, A2 => n4407, ZN => n5873);
   U6788 : INV_X1 port map( A => n7405, ZN => n7402);
   U6790 : NAND2_X1 port map( A1 => n7479, A2 => n7953, ZN => n2324);
   U6791 : INV_X1 port map( A => n7951, ZN => n2325);
   U6792 : INV_X1 port map( A => n7952, ZN => n2326);
   U6793 : MUX2_X1 port map( A => n15282, B => n15128, S => n15127, Z => n15129
                           );
   U6794 : NOR2_X2 port map( A1 => n14528, A2 => n14527, ZN => n15127);
   U6795 : XNOR2_X1 port map( A => n7123, B => n7119, ZN => n3572);
   U6796 : INV_X1 port map( A => n2661, ZN => n2659);
   U6798 : OAI211_X2 port map( C1 => n19789, C2 => n6030, A => n6029, B => 
                           n6028, ZN => n7042);
   U6799 : OAI211_X2 port map( C1 => n12539, C2 => n12538, A => n2328, B => 
                           n2327, ZN => n3159);
   U6800 : NAND2_X1 port map( A1 => n12536, A2 => n12535, ZN => n2327);
   U6802 : NOR2_X1 port map( A1 => n14494, A2 => n3155, ZN => n14495);
   U6804 : NAND3_X1 port map( A1 => n9837, A2 => n20476, A3 => n8542, ZN => 
                           n2330);
   U6808 : INV_X1 port map( A => n12377, ZN => n2333);
   U6809 : XOR2_X1 port map( A => n13581, B => n13582, Z => n3062);
   U6810 : INV_X1 port map( A => n11604, ZN => n11605);
   U6811 : NOR2_X1 port map( A1 => n3669, A2 => n11339, ZN => n11266);
   U6812 : AOI22_X1 port map( A1 => n8068, A2 => n7622, B1 => n8067, B2 => 
                           n8179, ZN => n3526);
   U6813 : AOI22_X2 port map( A1 => n12876, A2 => n14050, B1 => n13932, B2 => 
                           n13931, ZN => n15188);
   U6814 : OR2_X2 port map( A1 => n2334, A2 => n4038, ZN => n5888);
   U6815 : NAND3_X1 port map( A1 => n3729, A2 => n3730, A3 => n18033, ZN => 
                           n3691);
   U6817 : NAND2_X1 port map( A1 => n8617, A2 => n19827, ZN => n8618);
   U6818 : INV_X1 port map( A => n12484, ZN => n12477);
   U6819 : NAND3_X1 port map( A1 => n14275, A2 => n14562, A3 => n14705, ZN => 
                           n2541);
   U6820 : NAND2_X1 port map( A1 => n15635, A2 => n15636, ZN => n15637);
   U6821 : NAND2_X1 port map( A1 => n18593, A2 => n20365, ZN => n17919);
   U6824 : NAND2_X1 port map( A1 => n8873, A2 => n9107, ZN => n8874);
   U6825 : AOI22_X2 port map( A1 => n17162, A2 => n17163, B1 => n17160, B2 => 
                           n17161, ZN => n18589);
   U6826 : INV_X1 port map( A => n13312, ZN => n13161);
   U6828 : OAI211_X1 port map( C1 => n8312, C2 => n8313, A => n2339, B => 
                           n20144, ZN => n8320);
   U6829 : NAND2_X1 port map( A1 => n8312, A2 => n19520, ZN => n2339);
   U6831 : NAND2_X1 port map( A1 => n13141, A2 => n13147, ZN => n12572);
   U6832 : NAND2_X1 port map( A1 => n20157, A2 => n14268, ZN => n14576);
   U6833 : NAND3_X2 port map( A1 => n2717, A2 => n2716, A3 => n14386, ZN => 
                           n15625);
   U6834 : OR2_X1 port map( A1 => n12934, A2 => n14327, ZN => n2535);
   U6835 : OAI211_X2 port map( C1 => n5597, C2 => n6026, A => n2343, B => n2342
                           , ZN => n6819);
   U6836 : NAND2_X1 port map( A1 => n5928, A2 => n5596, ZN => n2343);
   U6837 : NAND2_X1 port map( A1 => n11008, A2 => n12576, ZN => n2346);
   U6838 : OAI21_X2 port map( B1 => n4347, B2 => n4203, A => n4202, ZN => n5670
                           );
   U6839 : NAND3_X1 port map( A1 => n2348, A2 => n18579, A3 => n18578, ZN => 
                           n18580);
   U6840 : OAI21_X1 port map( B1 => n18575, B2 => n18576, A => n19665, ZN => 
                           n2348);
   U6842 : NOR2_X1 port map( A1 => n12082, A2 => n12427, ZN => n12086);
   U6843 : XNOR2_X1 port map( A => n13266, B => n19854, ZN => n13579);
   U6845 : AND2_X1 port map( A1 => n2350, A2 => n12110, ZN => n11622);
   U6846 : INV_X1 port map( A => n12443, ZN => n2350);
   U6847 : MUX2_X1 port map( A => n8671, B => n8586, S => n19857, Z => n2351);
   U6848 : XNOR2_X1 port map( A => n2352, B => n16755, ZN => n16757);
   U6849 : XNOR2_X1 port map( A => n17335, B => n17989, ZN => n2352);
   U6850 : NAND3_X1 port map( A1 => n5735, A2 => n5763, A3 => n5736, ZN => 
                           n5737);
   U6852 : OAI211_X1 port map( C1 => n11193, C2 => n10903, A => n2355, B => 
                           n2354, ZN => n10625);
   U6853 : NAND2_X1 port map( A1 => n10577, A2 => n11193, ZN => n2354);
   U6854 : NAND2_X1 port map( A1 => n10576, A2 => n11186, ZN => n2355);
   U6856 : OR2_X1 port map( A1 => n7908, A2 => n6904, ZN => n7003);
   U6857 : INV_X1 port map( A => n13180, ZN => n15778);
   U6858 : XNOR2_X1 port map( A => n10574, B => n10568, ZN => n2496);
   U6859 : NAND2_X1 port map( A1 => n15336, A2 => n15341, ZN => n15467);
   U6861 : AND3_X2 port map( A1 => n2358, A2 => n14333, A3 => n2357, ZN => 
                           n16300);
   U6862 : NAND2_X1 port map( A1 => n14332, A2 => n20502, ZN => n2357);
   U6864 : OAI21_X1 port map( B1 => n18120, B2 => n19876, A => n2359, ZN => 
                           n18125);
   U6865 : NAND2_X1 port map( A1 => n19876, A2 => n18121, ZN => n2359);
   U6866 : NAND2_X1 port map( A1 => n19069, A2 => n19685, ZN => n19055);
   U6867 : MUX2_X1 port map( A => n10731, B => n10732, S => n11493, Z => n2360)
                           ;
   U6868 : NAND2_X1 port map( A1 => n3117, A2 => n17828, ZN => n3116);
   U6869 : OR2_X1 port map( A1 => n4602, A2 => n4355, ZN => n4605);
   U6870 : NAND2_X1 port map( A1 => n11204, A2 => n11209, ZN => n11097);
   U6871 : NAND2_X1 port map( A1 => n3297, A2 => n3298, ZN => n9381);
   U6872 : XNOR2_X1 port map( A => n2362, B => n2361, ZN => Ciphertext(120));
   U6873 : NAND3_X1 port map( A1 => n20467, A2 => n15167, A3 => n3621, ZN => 
                           n2363);
   U6874 : NAND2_X1 port map( A1 => n15382, A2 => n20103, ZN => n2364);
   U6875 : NAND2_X1 port map( A1 => n17488, A2 => n16800, ZN => n2692);
   U6876 : NAND2_X1 port map( A1 => n2365, A2 => n10862, ZN => n10868);
   U6877 : INV_X1 port map( A => n14518, ZN => n13564);
   U6878 : NAND2_X1 port map( A1 => n20272, A2 => n15121, ZN => n14518);
   U6880 : NAND2_X1 port map( A1 => n2367, A2 => n2366, ZN => n13063);
   U6881 : NAND3_X1 port map( A1 => n4909, A2 => n4910, A3 => n4954, ZN => 
                           n4918);
   U6883 : OAI211_X1 port map( C1 => n4136, C2 => n3231, A => n3230, B => n4377
                           , ZN => n3229);
   U6885 : AOI21_X1 port map( B1 => n8239, B2 => n7862, A => n8111, ZN => n3772
                           );
   U6886 : NAND3_X1 port map( A1 => n7779, A2 => n8007, A3 => n8313, ZN => 
                           n7778);
   U6887 : OR2_X1 port map( A1 => n4361, A2 => n4362, ZN => n2370);
   U6888 : NAND2_X1 port map( A1 => n9176, A2 => n8761, ZN => n8760);
   U6891 : OAI21_X1 port map( B1 => n11960, B2 => n1371, A => n3721, ZN => 
                           n3720);
   U6892 : NOR2_X1 port map( A1 => n16636, A2 => n2372, ZN => n16637);
   U6893 : NAND2_X1 port map( A1 => n16635, A2 => n19348, ZN => n2372);
   U6894 : NAND2_X1 port map( A1 => n14849, A2 => n15655, ZN => n15243);
   U6896 : NOR2_X1 port map( A1 => n15562, A2 => n15510, ZN => n2373);
   U6897 : MUX2_X1 port map( A => n18763, B => n18773, S => n18774, Z => n18767
                           );
   U6899 : AOI22_X2 port map( A1 => n13975, A2 => n14306, B1 => n13871, B2 => 
                           n13870, ZN => n15192);
   U6900 : NOR2_X2 port map( A1 => n2374, A2 => n2814, ZN => n17410);
   U6901 : NOR2_X1 port map( A1 => n3689, A2 => n3690, ZN => n15765);
   U6902 : OAI22_X1 port map( A1 => n12095, A2 => n2805, B1 => n12429, B2 => 
                           n12645, ZN => n2804);
   U6903 : INV_X1 port map( A => n4910, ZN => n3079);
   U6906 : NAND2_X1 port map( A1 => n8203, A2 => n8070, ZN => n2378);
   U6907 : AND2_X1 port map( A1 => n15454, A2 => n15777, ZN => n13095);
   U6908 : AND2_X1 port map( A1 => n231, A2 => n15379, ZN => n15030);
   U6909 : NAND2_X1 port map( A1 => n14418, A2 => n13937, ZN => n14054);
   U6910 : NAND2_X1 port map( A1 => n14377, A2 => n15846, ZN => n2380);
   U6911 : INV_X1 port map( A => n6113, ZN => n6108);
   U6912 : INV_X1 port map( A => n14449, ZN => n14455);
   U6913 : NOR2_X1 port map( A1 => n11646, A2 => n12121, ZN => n12123);
   U6915 : NOR2_X1 port map( A1 => n12919, A2 => n701, ZN => n12926);
   U6916 : INV_X1 port map( A => n7632, ZN => n8094);
   U6919 : INV_X1 port map( A => n5674, ZN => n5673);
   U6920 : OR3_X1 port map( A1 => n8741, A2 => n8743, A3 => n8742, ZN => n7649)
                           ;
   U6921 : NAND3_X1 port map( A1 => n12226, A2 => n12224, A3 => n12220, ZN => 
                           n10934);
   U6922 : NAND2_X1 port map( A1 => n7623, A2 => n8067, ZN => n2387);
   U6923 : NAND4_X2 port map( A1 => n12218, A2 => n12216, A3 => n12215, A4 => 
                           n12217, ZN => n13295);
   U6926 : NAND2_X1 port map( A1 => n4116, A2 => n2389, ZN => n4885);
   U6927 : AOI21_X1 port map( B1 => n12646, B2 => n2805, A => n3647, ZN => 
                           n3646);
   U6928 : NAND2_X1 port map( A1 => n4508, A2 => n4509, ZN => n4515);
   U6929 : NAND2_X1 port map( A1 => n14423, A2 => n14422, ZN => n2390);
   U6930 : NAND2_X1 port map( A1 => n14421, A2 => n2039, ZN => n2391);
   U6931 : OAI21_X1 port map( B1 => n1055, B2 => n1022, A => n2393, ZN => 
                           n17632);
   U6932 : NAND2_X1 port map( A1 => n17631, A2 => n1055, ZN => n2393);
   U6933 : NAND2_X1 port map( A1 => n5767, A2 => n5766, ZN => n5225);
   U6934 : OAI21_X2 port map( B1 => n12564, B2 => n12267, A => n12266, ZN => 
                           n13616);
   U6937 : INV_X1 port map( A => n17878, ZN => n3345);
   U6939 : NAND2_X1 port map( A1 => n8734, A2 => n8736, ZN => n8921);
   U6940 : OAI21_X1 port map( B1 => n7934, B2 => n20195, A => n7936, ZN => 
                           n7520);
   U6941 : XNOR2_X1 port map( A => n17400, B => n3091, ZN => n3090);
   U6942 : XNOR2_X2 port map( A => n6934, B => n2397, ZN => n8166);
   U6943 : XNOR2_X1 port map( A => n6932, B => n6933, ZN => n2397);
   U6946 : NAND2_X1 port map( A1 => n4358, A2 => n4546, ZN => n4311);
   U6947 : AOI21_X1 port map( B1 => n8729, B2 => n2400, A => n8947, ZN => n8594
                           );
   U6950 : INV_X1 port map( A => n11399, ZN => n2725);
   U6951 : NAND2_X1 port map( A1 => n20097, A2 => n18813, ZN => n17991);
   U6952 : NAND2_X1 port map( A1 => n14673, A2 => n3373, ZN => n2402);
   U6953 : INV_X1 port map( A => n2404, ZN => n2403);
   U6954 : NAND2_X1 port map( A1 => n5024, A2 => n4271, ZN => n4581);
   U6955 : AOI21_X2 port map( B1 => n7410, B2 => n7409, A => n2405, ZN => n8749
                           );
   U6956 : OAI211_X2 port map( C1 => n4584, C2 => n5026, A => n4583, B => n4582
                           , ZN => n6189);
   U6957 : OAI21_X1 port map( B1 => n5796, B2 => n2407, A => n2406, ZN => n5431
                           );
   U6958 : NAND2_X1 port map( A1 => n5790, A2 => n5796, ZN => n2406);
   U6959 : OAI21_X1 port map( B1 => n20377, B2 => n19918, A => n2408, ZN => 
                           n3329);
   U6960 : NAND2_X1 port map( A1 => n1262, A2 => n19918, ZN => n2408);
   U6961 : NAND2_X1 port map( A1 => n17592, A2 => n20150, ZN => n17593);
   U6962 : INV_X1 port map( A => n20141, ZN => n2412);
   U6963 : NAND2_X1 port map( A1 => n19361, A2 => n19366, ZN => n2414);
   U6964 : NAND2_X1 port map( A1 => n2415, A2 => n5686, ZN => n5183);
   U6965 : NAND2_X1 port map( A1 => n6084, A2 => n5683, ZN => n2415);
   U6966 : AND3_X1 port map( A1 => n5485, A2 => n5486, A3 => n5487, ZN => n3746
                           );
   U6967 : INV_X1 port map( A => n10897, ZN => n11210);
   U6968 : INV_X1 port map( A => n5888, ZN => n5309);
   U6969 : OR2_X1 port map( A1 => n14823, A2 => n12931, ZN => n3442);
   U6970 : INV_X1 port map( A => n14556, ZN => n14677);
   U6971 : INV_X1 port map( A => n5720, ZN => n3086);
   U6972 : OAI21_X1 port map( B1 => n2419, B2 => n20146, A => n2418, ZN => 
                           n9133);
   U6973 : OAI21_X1 port map( B1 => n11482, B2 => n11211, A => n10059, ZN => 
                           n11073);
   U6974 : OAI21_X1 port map( B1 => n17496, B2 => n17495, A => n2421, ZN => 
                           n3217);
   U6975 : NAND2_X1 port map( A1 => n2422, A2 => n17495, ZN => n2421);
   U6976 : INV_X1 port map( A => n14722, ZN => n13671);
   U6977 : XNOR2_X1 port map( A => n2542, B => n16695, ZN => n16835);
   U6978 : INV_X1 port map( A => n6744, ZN => n6552);
   U6979 : INV_X1 port map( A => n9564, ZN => n9342);
   U6980 : XNOR2_X1 port map( A => n13697, B => n12448, ZN => n12458);
   U6981 : INV_X1 port map( A => n8905, ZN => n3493);
   U6982 : NAND2_X1 port map( A1 => n8720, A2 => n9354, ZN => n8905);
   U6983 : OAI211_X2 port map( C1 => n6656, C2 => n6655, A => n3288, B => n2425
                           , ZN => n10445);
   U6984 : INV_X1 port map( A => n15744, ZN => n15749);
   U6985 : NAND2_X1 port map( A1 => n15593, A2 => n19502, ZN => n15744);
   U6987 : NAND2_X1 port map( A1 => n2429, A2 => n2427, ZN => n2426);
   U6988 : NAND2_X1 port map( A1 => n12207, A2 => n2428, ZN => n2427);
   U6989 : INV_X1 port map( A => n12209, ZN => n2428);
   U6990 : NAND2_X1 port map( A1 => n12189, A2 => n12209, ZN => n2429);
   U6991 : XNOR2_X1 port map( A => n2430, B => n19853, ZN => n8936);
   U6992 : XNOR2_X1 port map( A => n10039, B => n17637, ZN => n2430);
   U6993 : INV_X1 port map( A => n9241, ZN => n8628);
   U6994 : INV_X1 port map( A => n12350, ZN => n2737);
   U6995 : NAND2_X1 port map( A1 => n12467, A2 => n12138, ZN => n2431);
   U6996 : NAND2_X1 port map( A1 => n12139, A2 => n12466, ZN => n2432);
   U6997 : NOR2_X1 port map( A1 => n14327, A2 => n14087, ZN => n14819);
   U6998 : XNOR2_X1 port map( A => n2433, B => n7162, ZN => n7167);
   U6999 : XNOR2_X1 port map( A => n7161, B => n7202, ZN => n2433);
   U7000 : AND2_X2 port map( A1 => n16663, A2 => n16664, ZN => n19453);
   U7001 : OAI21_X1 port map( B1 => n2435, B2 => n2434, A => n5945, ZN => n5461
                           );
   U7003 : INV_X1 port map( A => n15449, ZN => n2438);
   U7004 : NAND2_X1 port map( A1 => n2606, A2 => n10858, ZN => n2602);
   U7005 : NAND2_X1 port map( A1 => n15111, A2 => n15294, ZN => n15108);
   U7006 : NAND2_X1 port map( A1 => n8135, A2 => n8382, ZN => n7498);
   U7008 : AOI21_X1 port map( B1 => n3503, B2 => n9215, A => n9210, ZN => n3502
                           );
   U7009 : NAND2_X1 port map( A1 => n18172, A2 => n19766, ZN => n18812);
   U7010 : NAND2_X1 port map( A1 => n9242, A2 => n2444, ZN => n2443);
   U7012 : OAI22_X1 port map( A1 => n2450, A2 => n2449, B1 => n19435, B2 => 
                           n19448, ZN => n19438);
   U7013 : NOR2_X1 port map( A1 => n3828, A2 => n19434, ZN => n2449);
   U7014 : NOR2_X1 port map( A1 => n3769, A2 => n4499, ZN => n2585);
   U7015 : INV_X1 port map( A => n10833, ZN => n10837);
   U7016 : NAND3_X1 port map( A1 => n2936, A2 => n5346, A3 => n3745, ZN => 
                           n4376);
   U7017 : INV_X1 port map( A => n11527, ZN => n2470);
   U7018 : NAND2_X1 port map( A1 => n3053, A2 => n8054, ZN => n6211);
   U7019 : NAND2_X1 port map( A1 => n16210, A2 => n16790, ZN => n16211);
   U7020 : NAND2_X1 port map( A1 => n7606, A2 => n8185, ZN => n8182);
   U7021 : NAND2_X1 port map( A1 => n3180, A2 => n14358, ZN => n2451);
   U7023 : OAI21_X1 port map( B1 => n15811, B2 => n15815, A => n3374, ZN => 
                           n15819);
   U7024 : NOR2_X1 port map( A1 => n8055, A2 => n8192, ZN => n3054);
   U7025 : AOI22_X1 port map( A1 => n10825, A2 => n11489, B1 => n10824, B2 => 
                           n11069, ZN => n12061);
   U7027 : OR3_X1 port map( A1 => n8993, A2 => n9274, A3 => n20265, ZN => n9279
                           );
   U7029 : NAND2_X1 port map( A1 => n9115, A2 => n9218, ZN => n9116);
   U7032 : OAI21_X1 port map( B1 => n14439, B2 => n14441, A => n238, ZN => 
                           n13557);
   U7033 : NAND2_X1 port map( A1 => n8201, A2 => n8070, ZN => n8072);
   U7034 : NAND2_X1 port map( A1 => n2458, A2 => n11173, ZN => n3359);
   U7035 : OAI21_X1 port map( B1 => n3789, B2 => n11174, A => n3362, ZN => 
                           n2458);
   U7036 : NAND2_X1 port map( A1 => n3358, A2 => n2457, ZN => n12224);
   U7037 : OR2_X1 port map( A1 => n11176, A2 => n2458, ZN => n2457);
   U7040 : OAI21_X1 port map( B1 => n6013, B2 => n6007, A => n6011, ZN => n5208
                           );
   U7041 : INV_X1 port map( A => n5098, ZN => n2460);
   U7042 : INV_X1 port map( A => n5092, ZN => n2461);
   U7043 : AND2_X1 port map( A1 => n5092, A2 => n5093, ZN => n2462);
   U7044 : NAND3_X1 port map( A1 => n2464, A2 => n11080, A3 => n2463, ZN => 
                           n12258);
   U7045 : NAND3_X1 port map( A1 => n11077, A2 => n11474, A3 => n11079, ZN => 
                           n2463);
   U7046 : NAND2_X1 port map( A1 => n3507, A2 => n11076, ZN => n11079);
   U7047 : NAND3_X1 port map( A1 => n2466, A2 => n5311, A3 => n5144, ZN => 
                           n2465);
   U7048 : INV_X1 port map( A => n5781, ZN => n2467);
   U7049 : NAND2_X1 port map( A1 => n11530, A2 => n11528, ZN => n2469);
   U7050 : NAND2_X1 port map( A1 => n15626, A2 => n2472, ZN => n2471);
   U7051 : NAND2_X1 port map( A1 => n15840, A2 => n15625, ZN => n15626);
   U7052 : NAND2_X1 port map( A1 => n2475, A2 => n2473, ZN => n2797);
   U7053 : NAND2_X1 port map( A1 => n2474, A2 => n18130, ZN => n2473);
   U7054 : NAND2_X1 port map( A1 => n18131, A2 => n17946, ZN => n2474);
   U7055 : INV_X1 port map( A => n19974, ZN => n2475);
   U7056 : NAND4_X2 port map( A1 => n7662, A2 => n2479, A3 => n7660, A4 => 
                           n2478, ZN => n10163);
   U7057 : NAND2_X1 port map( A1 => n8747, A2 => n8932, ZN => n8924);
   U7059 : NAND2_X1 port map( A1 => n4491, A2 => n4899, ZN => n2480);
   U7060 : AND2_X1 port map( A1 => n4883, A2 => n2482, ZN => n2481);
   U7061 : NAND2_X1 port map( A1 => n2483, A2 => n2487, ZN => n11892);
   U7062 : NAND2_X1 port map( A1 => n2484, A2 => n2486, ZN => n2483);
   U7063 : INV_X1 port map( A => n11119, ZN => n2486);
   U7064 : NAND2_X1 port map( A1 => n11036, A2 => n11119, ZN => n2487);
   U7066 : INV_X1 port map( A => Plaintext(17), ZN => n2488);
   U7067 : NAND2_X1 port map( A1 => n4986, A2 => n2489, ZN => n4991);
   U7068 : INV_X1 port map( A => n4302, ZN => n2490);
   U7069 : NAND2_X1 port map( A1 => n12513, A2 => n10625, ZN => n13270);
   U7071 : NAND2_X1 port map( A1 => n13275, A2 => n20073, ZN => n2491);
   U7072 : NAND2_X1 port map( A1 => n2493, A2 => n5455, ZN => n2559);
   U7073 : NAND4_X2 port map( A1 => n5173, A2 => n2493, A3 => n5175, A4 => 
                           n5174, ZN => n6634);
   U7074 : NAND2_X1 port map( A1 => n6108, A2 => n5656, ZN => n2493);
   U7075 : XNOR2_X1 port map( A => n10569, B => n10573, ZN => n2495);
   U7076 : NAND2_X1 port map( A1 => n2499, A2 => n8790, ZN => n7928);
   U7077 : NAND2_X1 port map( A1 => n9148, A2 => n2499, ZN => n8785);
   U7078 : NOR2_X1 port map( A1 => n9148, A2 => n2499, ZN => n9150);
   U7079 : NAND2_X1 port map( A1 => n20019, A2 => n17886, ZN => n17665);
   U7080 : AND2_X1 port map( A1 => n20019, A2 => n19947, ZN => n17599);
   U7081 : NAND2_X1 port map( A1 => n3247, A2 => n2500, ZN => n14888);
   U7082 : NAND2_X1 port map( A1 => n2501, A2 => n9145, ZN => n7929);
   U7083 : NAND3_X1 port map( A1 => n9145, A2 => n8786, A3 => n2501, ZN => 
                           n8787);
   U7084 : XNOR2_X1 port map( A => n9960, B => n2505, ZN => n9324);
   U7085 : INV_X1 port map( A => n10026, ZN => n2505);
   U7086 : OR2_X1 port map( A1 => n17094, A2 => n2507, ZN => n2513);
   U7087 : NAND2_X1 port map( A1 => n2517, A2 => n17095, ZN => n2507);
   U7088 : NAND2_X1 port map( A1 => n17092, A2 => n212, ZN => n2517);
   U7089 : OAI21_X1 port map( B1 => n2508, B2 => n17094, A => n2511, ZN => 
                           n2510);
   U7090 : INV_X1 port map( A => n2517, ZN => n2508);
   U7091 : OAI211_X1 port map( C1 => n2513, C2 => n2512, A => n2510, B => n2509
                           , ZN => Ciphertext(190));
   U7092 : INV_X1 port map( A => n17095, ZN => n2511);
   U7093 : INV_X1 port map( A => n2514, ZN => n2512);
   U7094 : NAND2_X1 port map( A1 => n2516, A2 => n2515, ZN => n2514);
   U7095 : XNOR2_X1 port map( A => n12559, B => n2518, ZN => n2519);
   U7096 : XNOR2_X1 port map( A => n12826, B => n12027, ZN => n13213);
   U7097 : XNOR2_X1 port map( A => n12826, B => n2521, ZN => n2520);
   U7099 : NAND2_X1 port map( A1 => n2523, A2 => n12389, ZN => n12391);
   U7100 : OAI211_X1 port map( C1 => n245, C2 => n2523, A => n12389, B => 
                           n11313, ZN => n11314);
   U7101 : NAND2_X1 port map( A1 => n12757, A2 => n2523, ZN => n12758);
   U7102 : NAND2_X1 port map( A1 => n19404, A2 => n17650, ZN => n2527);
   U7104 : INV_X1 port map( A => n15636, ZN => n2530);
   U7105 : XNOR2_X1 port map( A => n2531, B => n17686, ZN => Ciphertext(164));
   U7106 : OAI211_X1 port map( C1 => n20444, C2 => n19261, A => n2534, B => 
                           n2532, ZN => n2531);
   U7107 : OAI211_X1 port map( C1 => n2816, C2 => n19269, A => n2533, B => 
                           n19267, ZN => n2532);
   U7108 : NAND2_X1 port map( A1 => n17685, A2 => n19276, ZN => n2534);
   U7110 : XNOR2_X1 port map( A => n13259, B => n13602, ZN => n12834);
   U7112 : NAND2_X1 port map( A1 => n12393, A2 => n12479, ZN => n2538);
   U7113 : INV_X1 port map( A => n7935, ZN => n2540);
   U7114 : NAND2_X1 port map( A1 => n2540, A2 => n20359, ZN => n7930);
   U7117 : XNOR2_X1 port map( A => n2542, B => n16980, ZN => n16756);
   U7118 : XNOR2_X1 port map( A => n16507, B => n20121, ZN => n16142);
   U7119 : XNOR2_X1 port map( A => n20121, B => n16081, ZN => n16083);
   U7120 : NAND3_X1 port map( A1 => n19802, A2 => n7879, A3 => n3055, ZN => 
                           n2543);
   U7121 : OAI21_X1 port map( B1 => n2546, B2 => n18409, A => n18408, ZN => 
                           n18411);
   U7122 : NAND2_X1 port map( A1 => n8325, A2 => n2548, ZN => n7442);
   U7123 : AOI21_X1 port map( B1 => n7590, B2 => n2548, A => n8322, ZN => n3221
                           );
   U7125 : OAI211_X2 port map( C1 => n2553, C2 => n12394, A => n2549, B => 
                           n2554, ZN => n13528);
   U7126 : NAND3_X1 port map( A1 => n2552, A2 => n2551, A3 => n2550, ZN => 
                           n2549);
   U7127 : NAND2_X1 port map( A1 => n11931, A2 => n12478, ZN => n2551);
   U7128 : NAND2_X1 port map( A1 => n12141, A2 => n12480, ZN => n12394);
   U7129 : NAND2_X1 port map( A1 => n11932, A2 => n11931, ZN => n2554);
   U7130 : OR2_X1 port map( A1 => n5458, A2 => n6097, ZN => n2555);
   U7131 : NAND2_X1 port map( A1 => n1011, A2 => n6097, ZN => n2556);
   U7132 : XNOR2_X1 port map( A => n7070, B => n2557, ZN => n6225);
   U7133 : NAND3_X1 port map( A1 => n2559, A2 => n2560, A3 => n2558, ZN => 
                           n2557);
   U7134 : NAND3_X1 port map( A1 => n6108, A2 => n5656, A3 => n6109, ZN => 
                           n2560);
   U7136 : OAI21_X2 port map( B1 => n13875, B2 => n13874, A => n13873, ZN => 
                           n15496);
   U7137 : XNOR2_X2 port map( A => n10364, B => n10363, ZN => n11110);
   U7139 : XNOR2_X2 port map( A => n10355, B => n10354, ZN => n11452);
   U7142 : NAND2_X1 port map( A1 => n3386, A2 => n7820, ZN => n3384);
   U7143 : MUX2_X1 port map( A => n3387, B => n3386, S => n7820, Z => n2561);
   U7144 : NOR2_X1 port map( A1 => n981, A2 => n2562, ZN => n11831);
   U7145 : NOR2_X1 port map( A1 => n13973, A2 => n2563, ZN => n2564);
   U7146 : NAND2_X1 port map( A1 => n2566, A2 => n20443, ZN => n2565);
   U7147 : NAND2_X1 port map( A1 => n2568, A2 => n2567, ZN => n2566);
   U7148 : NAND2_X1 port map( A1 => n951, A2 => n14525, ZN => n2567);
   U7149 : NAND2_X1 port map( A1 => n19634, A2 => n14648, ZN => n2568);
   U7150 : XNOR2_X1 port map( A => n20216, B => n7035, ZN => n7229);
   U7151 : XNOR2_X1 port map( A => n20216, B => n6735, ZN => n6423);
   U7152 : XNOR2_X1 port map( A => n20216, B => n7360, ZN => n7362);
   U7154 : INV_X1 port map( A => n5611, ZN => n6151);
   U7155 : NAND2_X1 port map( A1 => n2576, A2 => n2595, ZN => n2572);
   U7157 : NAND2_X1 port map( A1 => n2579, A2 => n20533, ZN => n2577);
   U7158 : NAND2_X1 port map( A1 => n2580, A2 => n15905, ZN => n2579);
   U7159 : NAND2_X1 port map( A1 => n15907, A2 => n15909, ZN => n2580);
   U7162 : INV_X1 port map( A => n13838, ZN => n2582);
   U7163 : NAND3_X1 port map( A1 => n2583, A2 => n6153, A3 => n6150, ZN => 
                           n5614);
   U7164 : NAND2_X1 port map( A1 => n5611, A2 => n5349, ZN => n2583);
   U7165 : NAND2_X1 port map( A1 => n4379, A2 => n4857, ZN => n2584);
   U7166 : OR2_X1 port map( A1 => n19933, A2 => n17812, ZN => n17690);
   U7167 : NAND2_X1 port map( A1 => n2587, A2 => n18046, ZN => n17317);
   U7168 : NAND2_X1 port map( A1 => n19933, A2 => n17812, ZN => n2587);
   U7173 : INV_X1 port map( A => n17812, ZN => n2590);
   U7174 : NAND2_X1 port map( A1 => n2592, A2 => n14787, ZN => n2591);
   U7175 : NAND2_X1 port map( A1 => n14343, A2 => n14790, ZN => n2593);
   U7176 : NAND2_X1 port map( A1 => n14103, A2 => n14791, ZN => n2594);
   U7177 : NAND2_X1 port map( A1 => n4377, A2 => n4899, ZN => n2595);
   U7178 : NAND2_X1 port map( A1 => n20205, A2 => n4960, ZN => n2596);
   U7180 : NAND2_X1 port map( A1 => n20057, A2 => n19865, ZN => n2597);
   U7181 : NAND2_X1 port map( A1 => n2598, A2 => n12542, ZN => n12547);
   U7182 : INV_X1 port map( A => n12545, ZN => n2598);
   U7183 : NOR2_X1 port map( A1 => n2601, A2 => n3978, ZN => n3977);
   U7184 : INV_X1 port map( A => n4657, ZN => n2601);
   U7185 : NAND2_X1 port map( A1 => n2603, A2 => n2602, ZN => n12619);
   U7186 : NAND2_X1 port map( A1 => n2610, A2 => n10858, ZN => n2603);
   U7187 : NAND2_X1 port map( A1 => n2604, A2 => n894, ZN => n2608);
   U7189 : NAND2_X1 port map( A1 => n2607, A2 => n10858, ZN => n12057);
   U7190 : NAND3_X1 port map( A1 => n12059, A2 => n12053, A3 => n2608, ZN => 
                           n11634);
   U7191 : AOI21_X1 port map( B1 => n2612, B2 => n11773, A => n3260, ZN => 
                           n11774);
   U7192 : NAND2_X1 port map( A1 => n12313, A2 => n12148, ZN => n2612);
   U7193 : OAI21_X1 port map( B1 => n6069, B2 => n5879, A => n2613, ZN => n5883
                           );
   U7194 : NAND3_X1 port map( A1 => n6069, A2 => n6075, A3 => n6067, ZN => 
                           n2613);
   U7195 : NAND2_X1 port map( A1 => n6069, A2 => n6067, ZN => n2616);
   U7196 : NAND2_X1 port map( A1 => n2616, A2 => n6070, ZN => n2614);
   U7197 : NAND2_X1 port map( A1 => n5979, A2 => n5320, ZN => n2615);
   U7198 : NAND2_X1 port map( A1 => n969, A2 => n2617, ZN => n9643);
   U7199 : XNOR2_X1 port map( A => n10594, B => n10105, ZN => n10106);
   U7200 : XNOR2_X1 port map( A => n2619, B => n12862, ZN => n14452);
   U7201 : XNOR2_X1 port map( A => n13708, B => n2620, ZN => n2619);
   U7202 : XNOR2_X1 port map( A => n2621, B => n6659, ZN => n2622);
   U7203 : INV_X1 port map( A => n6588, ZN => n2621);
   U7205 : XNOR2_X1 port map( A => n13771, B => n13769, ZN => n2624);
   U7206 : NAND2_X1 port map( A1 => n8644, A2 => n8937, ZN => n2955);
   U7207 : OAI211_X1 port map( C1 => n15885, C2 => n2625, A => n16017, B => 
                           n14926, ZN => n14927);
   U7208 : NAND2_X1 port map( A1 => n16012, A2 => n19740, ZN => n2625);
   U7209 : NAND2_X1 port map( A1 => n2627, A2 => n8018, ZN => n7804);
   U7210 : INV_X1 port map( A => n14584, ZN => n2628);
   U7211 : NAND2_X1 port map( A1 => n2629, A2 => n6166, ZN => n5462);
   U7212 : MUX2_X1 port map( A => n1867, B => n170, S => n6172, Z => n4692);
   U7213 : NAND2_X1 port map( A1 => n5843, A2 => n2630, ZN => n7274);
   U7214 : NOR2_X1 port map( A1 => n9135, A2 => n2727, ZN => n2631);
   U7215 : OR2_X1 port map( A1 => n5073, A2 => n291, ZN => n4662);
   U7216 : INV_X1 port map( A => n4816, ZN => n2632);
   U7217 : NAND2_X1 port map( A1 => n20168, A2 => n19814, ZN => n16442);
   U7218 : NAND2_X1 port map( A1 => n2634, A2 => n9218, ZN => n8429);
   U7219 : INV_X1 port map( A => n9118, ZN => n2634);
   U7220 : NAND2_X1 port map( A1 => n9217, A2 => n9221, ZN => n9118);
   U7221 : AOI22_X1 port map( A1 => n267, A2 => n9189, B1 => n8713, B2 => n9241
                           , ZN => n9243);
   U7223 : NAND2_X1 port map( A1 => n2637, A2 => n6587, ZN => n2636);
   U7224 : NAND2_X1 port map( A1 => n987, A2 => n5328, ZN => n2638);
   U7225 : NAND2_X1 port map( A1 => n2641, A2 => n5328, ZN => n2640);
   U7228 : NOR2_X1 port map( A1 => n15297, A2 => n15111, ZN => n2645);
   U7229 : OR2_X1 port map( A1 => n15108, A2 => n15109, ZN => n2646);
   U7230 : INV_X1 port map( A => n12047, ZN => n2647);
   U7231 : NAND2_X1 port map( A1 => n2647, A2 => n12122, ZN => n11647);
   U7232 : INV_X1 port map( A => n12047, ZN => n12229);
   U7234 : NAND2_X1 port map( A1 => n3156, A2 => n14746, ZN => n3155);
   U7235 : OAI21_X1 port map( B1 => n8183, B2 => n8059, A => n2648, ZN => n8065
                           );
   U7236 : NAND2_X1 port map( A1 => n4730, A2 => n2649, ZN => n2648);
   U7237 : NAND2_X1 port map( A1 => n19716, A2 => n8630, ZN => n2652);
   U7238 : OR2_X1 port map( A1 => n13911, A2 => n13907, ZN => n2654);
   U7239 : NOR2_X1 port map( A1 => n15857, A2 => n2655, ZN => n15858);
   U7240 : AOI22_X1 port map( A1 => n15722, A2 => n15864, B1 => n15721, B2 => 
                           n2655, ZN => n13916);
   U7241 : NAND2_X1 port map( A1 => n15859, A2 => n2655, ZN => n15725);
   U7243 : INV_X1 port map( A => n10450, ZN => n11094);
   U7246 : NAND3_X1 port map( A1 => n2662, A2 => n2664, A3 => n2660, ZN => 
                           n16810);
   U7247 : NAND2_X1 port map( A1 => n2661, A2 => n19658, ZN => n2660);
   U7248 : NAND3_X1 port map( A1 => n17552, A2 => n18103, A3 => n2665, ZN => 
                           n2664);
   U7249 : OR2_X1 port map( A1 => n17959, A2 => n17954, ZN => n2665);
   U7250 : INV_X1 port map( A => n16805, ZN => n18105);
   U7251 : NAND2_X1 port map( A1 => n6096, A2 => n6101, ZN => n3589);
   U7253 : NAND2_X1 port map( A1 => n3685, A2 => n2682, ZN => n2666);
   U7254 : NAND2_X1 port map( A1 => n19354, A2 => n20244, ZN => n2668);
   U7255 : AOI21_X2 port map( B1 => n15929, B2 => n2669, A => n15928, ZN => 
                           n18423);
   U7256 : NOR2_X1 port map( A1 => n4797, A2 => n5047, ZN => n2671);
   U7257 : NAND2_X1 port map( A1 => n2675, A2 => n2677, ZN => n2673);
   U7259 : NOR2_X1 port map( A1 => n15870, A2 => n15876, ZN => n15873);
   U7260 : MUX2_X1 port map( A => n14664, B => n14316, S => n14662, Z => n2678)
                           ;
   U7261 : XNOR2_X1 port map( A => n13842, B => n1004, ZN => n2679);
   U7262 : NAND2_X1 port map( A1 => n2680, A2 => n11475, ZN => n3135);
   U7263 : NAND2_X1 port map( A1 => n984, A2 => n2682, ZN => n2681);
   U7267 : NAND2_X1 port map( A1 => n5662, A2 => n6101, ZN => n5948);
   U7268 : INV_X1 port map( A => n8095, ZN => n2687);
   U7269 : OAI21_X1 port map( B1 => n8094, B2 => n8211, A => n2686, ZN => n2688
                           );
   U7270 : NAND2_X1 port map( A1 => n2687, A2 => n8212, ZN => n2686);
   U7271 : XNOR2_X2 port map( A => n6609, B => n6608, ZN => n8212);
   U7272 : XNOR2_X1 port map( A => n10351, B => n2689, ZN => n9724);
   U7273 : NAND2_X1 port map( A1 => n8759, A2 => n8650, ZN => n2690);
   U7277 : NAND2_X1 port map( A1 => n14348, A2 => n19496, ZN => n2695);
   U7278 : NAND2_X1 port map( A1 => n14349, A2 => n19985, ZN => n2698);
   U7279 : NAND2_X1 port map( A1 => n4089, A2 => n2701, ZN => n2699);
   U7281 : NAND2_X1 port map( A1 => n4697, A2 => n5040, ZN => n4799);
   U7282 : AND2_X1 port map( A1 => n4440, A2 => n4439, ZN => n2701);
   U7283 : OAI21_X1 port map( B1 => n11469, B2 => n11568, A => n2705, ZN => 
                           n2704);
   U7284 : AOI21_X1 port map( B1 => n10883, B2 => n11568, A => n11566, ZN => 
                           n2705);
   U7285 : XNOR2_X2 port map( A => n9951, B => n9950, ZN => n11568);
   U7286 : NAND2_X1 port map( A1 => n2707, A2 => n12352, ZN => n3330);
   U7287 : INV_X1 port map( A => n12353, ZN => n2707);
   U7290 : XNOR2_X1 port map( A => n12713, B => n2709, ZN => n12728);
   U7291 : MUX2_X1 port map( A => n7969, B => n7970, S => n7922, Z => n7977);
   U7292 : NAND2_X1 port map( A1 => n2714, A2 => n2711, ZN => n10849);
   U7293 : NAND2_X1 port map( A1 => n15838, A2 => n15625, ZN => n2715);
   U7294 : INV_X1 port map( A => n5279, ZN => n3398);
   U7295 : NAND2_X1 port map( A1 => n5669, A2 => n5425, ZN => n2719);
   U7296 : OAI22_X1 port map( A1 => n14340, A2 => n13931, B1 => n14337, B2 => 
                           n14342, ZN => n3331);
   U7297 : NAND2_X1 port map( A1 => n2722, A2 => n20533, ZN => n2721);
   U7298 : NAND2_X1 port map( A1 => n2725, A2 => n11395, ZN => n11401);
   U7299 : MUX2_X1 port map( A => n10859, B => n10860, S => n11399, Z => n10861
                           );
   U7300 : NAND3_X1 port map( A1 => n9214, A2 => n9209, A3 => n263, ZN => n8394
                           );
   U7301 : NAND3_X1 port map( A1 => n2731, A2 => n14620, A3 => n14192, ZN => 
                           n2730);
   U7302 : INV_X1 port map( A => n14627, ZN => n2731);
   U7303 : XNOR2_X1 port map( A => n13295, B => n2733, ZN => n13135);
   U7304 : OR2_X1 port map( A1 => n12469, A2 => n12470, ZN => n2732);
   U7305 : XNOR2_X1 port map( A => n13063, B => n855, ZN => n13400);
   U7306 : XNOR2_X1 port map( A => n855, B => n13848, ZN => n13851);
   U7307 : XNOR2_X1 port map( A => n13343, B => n2733, ZN => n12864);
   U7308 : INV_X1 port map( A => n10694, ZN => n10995);
   U7310 : NAND2_X1 port map( A1 => n19817, A2 => n19779, ZN => n2734);
   U7312 : OAI21_X1 port map( B1 => n19651, B2 => n7743, A => n2751, ZN => 
                           n7742);
   U7314 : AOI22_X2 port map( A1 => n7744, A2 => n7743, B1 => n7742, B2 => 
                           n7741, ZN => n7752);
   U7315 : NAND2_X1 port map( A1 => n11535, A2 => n11538, ZN => n2736);
   U7316 : OAI21_X1 port map( B1 => n11170, B2 => n11535, A => n2736, ZN => 
                           n8902);
   U7317 : INV_X1 port map( A => Plaintext(79), ZN => n2738);
   U7318 : NAND2_X1 port map( A1 => n3904, A2 => n4554, ZN => n5015);
   U7319 : NAND2_X1 port map( A1 => n3905, A2 => n2740, ZN => n2739);
   U7320 : NAND2_X1 port map( A1 => n5021, A2 => n5018, ZN => n2740);
   U7321 : NAND2_X1 port map( A1 => n3904, A2 => n4555, ZN => n5021);
   U7322 : AOI21_X2 port map( B1 => n15493, B2 => n15587, A => n2741, ZN => 
                           n17109);
   U7323 : MUX2_X1 port map( A => n15492, B => n15761, S => n15760, Z => n2741)
                           ;
   U7324 : NAND2_X1 port map( A1 => n12209, A2 => n12211, ZN => n2742);
   U7325 : XNOR2_X1 port map( A => n9852, B => n10182, ZN => n2745);
   U7326 : NAND2_X1 port map( A1 => n8733, A2 => n8736, ZN => n8920);
   U7327 : NAND2_X1 port map( A1 => n8733, A2 => n8735, ZN => n8332);
   U7328 : NAND2_X1 port map( A1 => n14706, A2 => n20113, ZN => n14564);
   U7329 : AOI21_X1 port map( B1 => n14704, B2 => n20113, A => n14563, ZN => 
                           n14111);
   U7330 : NOR2_X1 port map( A1 => n919, A2 => n20113, ZN => n14709);
   U7331 : OAI21_X1 port map( B1 => n9318, B2 => n2749, A => n9320, ZN => n9319
                           );
   U7332 : NOR2_X1 port map( A1 => n8860, A2 => n2749, ZN => n8864);
   U7333 : NAND2_X1 port map( A1 => n9322, A2 => n2749, ZN => n9838);
   U7334 : NAND2_X1 port map( A1 => n8354, A2 => n7739, ZN => n2751);
   U7335 : NAND2_X1 port map( A1 => n2754, A2 => n2753, ZN => n17309);
   U7336 : OR2_X1 port map( A1 => n18221, A2 => n18016, ZN => n2753);
   U7337 : NAND2_X1 port map( A1 => n17308, A2 => n18221, ZN => n2754);
   U7338 : OAI21_X1 port map( B1 => n224, B2 => n20421, A => n18977, ZN => 
                           n18980);
   U7339 : OAI21_X1 port map( B1 => n18224, B2 => n18223, A => n20421, ZN => 
                           n18721);
   U7340 : NAND2_X1 port map( A1 => n9353, A2 => n8904, ZN => n9357);
   U7341 : INV_X1 port map( A => n8720, ZN => n9353);
   U7342 : OAI21_X1 port map( B1 => n12600, B2 => n12606, A => n2757, ZN => 
                           n11630);
   U7343 : NAND2_X1 port map( A1 => n12609, A2 => n12600, ZN => n2757);
   U7344 : NAND2_X1 port map( A1 => n2762, A2 => n12241, ZN => n12620);
   U7345 : INV_X1 port map( A => n12619, ZN => n2762);
   U7346 : XNOR2_X1 port map( A => n2763, B => n13735, ZN => n13313);
   U7347 : INV_X1 port map( A => n13120, ZN => n2763);
   U7348 : XNOR2_X1 port map( A => n13792, B => n2764, ZN => n13793);
   U7349 : NAND2_X1 port map( A1 => n10818, A2 => n10677, ZN => n11369);
   U7350 : NOR2_X1 port map( A1 => n10676, A2 => n10677, ZN => n9875);
   U7351 : INV_X1 port map( A => n14229, ZN => n2769);
   U7353 : NAND2_X1 port map( A1 => n2769, A2 => n14381, ZN => n2767);
   U7354 : NAND2_X1 port map( A1 => n14697, A2 => n14232, ZN => n2768);
   U7355 : NAND2_X1 port map( A1 => n19503, A2 => n14381, ZN => n14697);
   U7357 : XNOR2_X1 port map( A => n10165, B => n20176, ZN => n2771);
   U7358 : XNOR2_X1 port map( A => n9586, B => n9588, ZN => n2772);
   U7359 : NAND2_X1 port map( A1 => n13919, A2 => n14167, ZN => n2774);
   U7362 : AOI21_X1 port map( B1 => n8568, B2 => n9168, A => n9082, ZN => n2777
                           );
   U7364 : NAND2_X1 port map( A1 => n235, A2 => n14818, ZN => n14823);
   U7365 : XNOR2_X1 port map( A => n12824, B => n12823, ZN => n2784);
   U7368 : NAND2_X1 port map( A1 => n2787, A2 => n9297, ZN => n2786);
   U7369 : NOR2_X1 port map( A1 => n8846, A2 => n9018, ZN => n2787);
   U7370 : NAND2_X1 port map( A1 => n11208, A2 => n2788, ZN => n12142);
   U7371 : NAND2_X1 port map( A1 => n958, A2 => n11445, ZN => n2788);
   U7373 : NAND2_X1 port map( A1 => n15406, A2 => n15547, ZN => n2791);
   U7374 : NAND2_X1 port map( A1 => n15546, A2 => n15071, ZN => n15616);
   U7375 : NAND2_X1 port map( A1 => n15618, A2 => n15405, ZN => n15547);
   U7376 : NAND2_X1 port map( A1 => n8305, A2 => n2792, ZN => n8306);
   U7377 : OAI211_X1 port map( C1 => n8303, C2 => n8301, A => n8044, B => n2792
                           , ZN => n7599);
   U7379 : NAND2_X1 port map( A1 => n5272, A2 => n2792, ZN => n3718);
   U7380 : INV_X1 port map( A => n20361, ZN => n2793);
   U7381 : OAI21_X1 port map( B1 => n5856, B2 => n5855, A => n2796, ZN => n2795
                           );
   U7383 : NAND2_X1 port map( A1 => n2799, A2 => n2800, ZN => n2798);
   U7384 : NAND2_X1 port map( A1 => n15072, A2 => n15620, ZN => n2801);
   U7385 : INV_X1 port map( A => n15546, ZN => n2803);
   U7386 : NAND3_X1 port map( A1 => n19668, A2 => n19682, A3 => n18552, ZN => 
                           n17931);
   U7388 : NAND2_X1 port map( A1 => n2809, A2 => n2807, ZN => n2806);
   U7389 : NAND2_X1 port map( A1 => n13888, A2 => n14593, ZN => n2807);
   U7390 : INV_X1 port map( A => n14590, ZN => n2808);
   U7391 : AND2_X1 port map( A1 => n12544, A2 => n250, ZN => n3462);
   U7392 : AOI21_X2 port map( B1 => n15299, B2 => n15298, A => n2812, ZN => 
                           n16095);
   U7393 : MUX2_X1 port map( A => n15297, B => n15296, S => n15295, Z => n2813)
                           ;
   U7394 : INV_X1 port map( A => n15759, ZN => n2815);
   U7395 : NAND3_X1 port map( A1 => n17661, A2 => n17662, A3 => n17890, ZN => 
                           n2817);
   U7396 : NAND3_X1 port map( A1 => n17665, A2 => n17661, A3 => n17662, ZN => 
                           n2818);
   U7397 : NAND2_X1 port map( A1 => n14027, A2 => n2820, ZN => n15488);
   U7398 : NAND2_X1 port map( A1 => n14574, A2 => n2821, ZN => n2820);
   U7399 : NAND2_X1 port map( A1 => n14268, A2 => n14569, ZN => n2821);
   U7400 : NAND2_X1 port map( A1 => n16262, A2 => n16777, ZN => n2822);
   U7401 : NAND2_X1 port map( A1 => n16264, A2 => n17824, ZN => n2823);
   U7403 : XNOR2_X1 port map( A => n7079, B => n6718, ZN => n2825);
   U7409 : OR2_X1 port map( A1 => n18603, A2 => n18630, ZN => n2830);
   U7411 : XNOR2_X1 port map( A => n13291, B => n2834, ZN => n2833);
   U7412 : NAND2_X1 port map( A1 => n2837, A2 => n2835, ZN => n17551);
   U7413 : XNOR2_X2 port map( A => n17115, B => n17114, ZN => n18233);
   U7415 : NAND2_X1 port map( A1 => n17548, A2 => n19771, ZN => n2837);
   U7416 : NAND2_X1 port map( A1 => n9209, A2 => n2727, ZN => n9212);
   U7417 : NAND3_X1 port map( A1 => n9209, A2 => n9135, A3 => n2727, ZN => 
                           n3454);
   U7418 : INV_X1 port map( A => n14800, ZN => n14081);
   U7419 : AOI21_X1 port map( B1 => n3497, B2 => n14796, A => n14584, ZN => 
                           n2838);
   U7420 : NAND2_X1 port map( A1 => n20380, A2 => n14522, ZN => n14652);
   U7421 : NAND3_X1 port map( A1 => n20380, A2 => n14522, A3 => n19831, ZN => 
                           n2839);
   U7422 : XNOR2_X2 port map( A => n13001, B => n13000, ZN => n14522);
   U7423 : NOR2_X1 port map( A1 => n2840, A2 => n8162, ZN => n8163);
   U7426 : NAND2_X1 port map( A1 => n19872, A2 => n2843, ZN => n2842);
   U7427 : NOR2_X1 port map( A1 => n11160, A2 => n11161, ZN => n2843);
   U7428 : NAND2_X1 port map( A1 => n11161, A2 => n11155, ZN => n2846);
   U7429 : NAND2_X1 port map( A1 => n2848, A2 => n9366, ZN => n2847);
   U7431 : NAND2_X1 port map( A1 => n9364, A2 => n2849, ZN => n2848);
   U7432 : NAND2_X1 port map( A1 => n8960, A2 => n8961, ZN => n2849);
   U7433 : NAND2_X1 port map( A1 => n8961, A2 => n8500, ZN => n9364);
   U7434 : NAND2_X1 port map( A1 => n9361, A2 => n9362, ZN => n8727);
   U7435 : NAND3_X1 port map( A1 => n3421, A2 => n2853, A3 => n2851, ZN => 
                           Ciphertext(28));
   U7436 : NAND2_X1 port map( A1 => n2852, A2 => n2854, ZN => n2851);
   U7437 : NAND2_X1 port map( A1 => n17639, A2 => n19729, ZN => n17647);
   U7438 : NAND3_X1 port map( A1 => n17639, A2 => n19729, A3 => n15134, ZN => 
                           n2853);
   U7439 : NAND2_X1 port map( A1 => n2855, A2 => n893, ZN => n2854);
   U7440 : INV_X1 port map( A => n17914, ZN => n2855);
   U7441 : NAND2_X1 port map( A1 => n18592, A2 => n18585, ZN => n18596);
   U7442 : INV_X1 port map( A => n11376, ZN => n2858);
   U7443 : OR2_X1 port map( A1 => n11330, A2 => n11376, ZN => n2857);
   U7444 : INV_X1 port map( A => n20095, ZN => n2860);
   U7445 : NAND2_X1 port map( A1 => n2860, A2 => n11376, ZN => n10661);
   U7446 : INV_X1 port map( A => n11328, ZN => n11378);
   U7447 : NOR2_X1 port map( A1 => n14811, A2 => n14810, ZN => n14588);
   U7449 : OAI21_X1 port map( B1 => n14589, B2 => n14590, A => n14588, ZN => 
                           n14591);
   U7450 : NAND2_X1 port map( A1 => n2864, A2 => n12498, ZN => n2863);
   U7451 : NAND2_X1 port map( A1 => n5732, A2 => n5802, ZN => n2867);
   U7452 : INV_X1 port map( A => n5045, ZN => n5043);
   U7453 : OAI21_X1 port map( B1 => n2872, B2 => n2871, A => n4796, ZN => n2870
                           );
   U7454 : NOR2_X1 port map( A1 => n4697, A2 => n5040, ZN => n2871);
   U7455 : NOR2_X1 port map( A1 => n3061, A2 => n5045, ZN => n2874);
   U7456 : INV_X1 port map( A => n20247, ZN => n8186);
   U7457 : MUX2_X1 port map( A => n20465, B => n8190, S => n8061, Z => n2875);
   U7458 : XNOR2_X1 port map( A => n3902, B => n7202, ZN => n3963);
   U7459 : NAND2_X1 port map( A1 => n2878, A2 => n2877, ZN => n2876);
   U7460 : NAND2_X1 port map( A1 => n992, A2 => n5429, ZN => n2877);
   U7461 : NAND2_X1 port map( A1 => n2879, A2 => n5793, ZN => n2878);
   U7463 : INV_X1 port map( A => n13243, ZN => n2881);
   U7464 : OAI21_X1 port map( B1 => n19958, B2 => n15583, A => n15811, ZN => 
                           n15584);
   U7465 : INV_X1 port map( A => n8995, ZN => n2883);
   U7466 : NAND2_X1 port map( A1 => n19517, A2 => n8997, ZN => n2884);
   U7467 : NAND2_X1 port map( A1 => n11431, A2 => n11430, ZN => n11042);
   U7469 : MUX2_X1 port map( A => n12269, B => n12374, S => n20497, Z => n11732
                           );
   U7473 : NAND2_X1 port map( A1 => n14697, A2 => n2891, ZN => n2890);
   U7474 : AOI22_X1 port map( A1 => n17903, A2 => n17904, B1 => n19229, B2 => 
                           n2892, ZN => n17905);
   U7475 : AOI22_X1 port map( A1 => n17915, A2 => n19236, B1 => n17916, B2 => 
                           n2892, ZN => n17917);
   U7476 : OAI22_X1 port map( A1 => n19236, A2 => n20124, B1 => n18190, B2 => 
                           n19754, ZN => n2892);
   U7477 : NOR2_X1 port map( A1 => n19166, A2 => n2893, ZN => n17797);
   U7478 : NAND2_X1 port map( A1 => n2895, A2 => n2894, ZN => n2893);
   U7479 : NAND2_X1 port map( A1 => n2918, A2 => n17790, ZN => n2894);
   U7480 : AOI21_X1 port map( B1 => n19165, B2 => n17790, A => n17791, ZN => 
                           n2895);
   U7481 : INV_X1 port map( A => n17791, ZN => n2896);
   U7483 : NAND2_X1 port map( A1 => n10899, A2 => n19897, ZN => n2899);
   U7484 : NAND2_X1 port map( A1 => n11482, A2 => n10746, ZN => n10898);
   U7485 : OAI21_X1 port map( B1 => n12497, B2 => n12499, A => n2901, ZN => 
                           n12503);
   U7486 : INV_X1 port map( A => n2903, ZN => n2902);
   U7489 : NAND2_X1 port map( A1 => n13953, A2 => n14408, ZN => n2905);
   U7490 : NAND2_X1 port map( A1 => n18957, A2 => n2906, ZN => n17068);
   U7493 : NAND2_X1 port map( A1 => n15509, A2 => n3822, ZN => n2908);
   U7494 : NAND3_X1 port map( A1 => n921, A2 => n15559, A3 => n15509, ZN => 
                           n14765);
   U7495 : NOR2_X1 port map( A1 => n15560, A2 => n921, ZN => n15561);
   U7496 : MUX2_X1 port map( A => n15559, B => n921, S => n15558, Z => n15563);
   U7499 : XNOR2_X1 port map( A => n2913, B => n2912, ZN => Ciphertext(142));
   U7500 : INV_X1 port map( A => n2410, ZN => n2912);
   U7501 : NAND3_X1 port map( A1 => n2917, A2 => n2916, A3 => n2914, ZN => 
                           n2913);
   U7502 : OAI211_X1 port map( C1 => n19692, C2 => n19708, A => n2915, B => 
                           n19948, ZN => n2914);
   U7503 : NAND2_X1 port map( A1 => n19692, A2 => n19154, ZN => n2915);
   U7504 : NAND3_X1 port map( A1 => n195, A2 => n19683, A3 => n19165, ZN => 
                           n2916);
   U7505 : NAND2_X1 port map( A1 => n18307, A2 => n2918, ZN => n2917);
   U7506 : AOI21_X1 port map( B1 => n3551, B2 => n2919, A => n4528, ZN => n3624
                           );
   U7507 : NAND2_X1 port map( A1 => n13557, A2 => n13558, ZN => n2920);
   U7508 : NAND2_X1 port map( A1 => n14442, A2 => n14440, ZN => n2921);
   U7509 : AOI21_X2 port map( B1 => n2927, B2 => n2926, A => n2922, ZN => 
                           n15559);
   U7510 : OAI22_X1 port map( A1 => n2925, A2 => n1527, B1 => n2926, B2 => 
                           n2923, ZN => n2922);
   U7511 : INV_X1 port map( A => n14393, ZN => n2924);
   U7512 : NAND2_X1 port map( A1 => n14594, A2 => n19731, ZN => n2925);
   U7513 : NAND2_X1 port map( A1 => n14156, A2 => n14155, ZN => n2927);
   U7514 : NAND2_X1 port map( A1 => n1527, A2 => n14594, ZN => n14156);
   U7515 : INV_X1 port map( A => n9240, ZN => n9186);
   U7516 : NAND2_X1 port map( A1 => n9266, A2 => n9265, ZN => n8981);
   U7518 : NAND2_X1 port map( A1 => n5056, A2 => n4100, ZN => n4590);
   U7519 : NAND2_X1 port map( A1 => n2929, A2 => n5053, ZN => n2928);
   U7520 : NAND2_X1 port map( A1 => n8358, A2 => n8357, ZN => n2932);
   U7521 : NAND2_X1 port map( A1 => n2935, A2 => n8347, ZN => n8273);
   U7522 : NAND2_X1 port map( A1 => n8272, A2 => n8350, ZN => n2935);
   U7523 : XNOR2_X1 port map( A => n9811, B => n9995, ZN => n2938);
   U7524 : MUX2_X1 port map( A => n11418, B => n11051, S => n11417, Z => n11130
                           );
   U7525 : MUX2_X1 port map( A => n11417, B => n11051, S => n205, Z => n10832);
   U7526 : NAND3_X1 port map( A1 => n8707, A2 => n1027, A3 => n2941, ZN => 
                           n9908);
   U7527 : XNOR2_X1 port map( A => n6293, B => n7232, ZN => n7057);
   U7528 : XNOR2_X1 port map( A => n6494, B => n6293, ZN => n6625);
   U7529 : NAND2_X1 port map( A1 => n2944, A2 => n2942, ZN => n2945);
   U7530 : AOI21_X1 port map( B1 => n19197, B2 => n2943, A => n19189, ZN => 
                           n2942);
   U7531 : NAND2_X1 port map( A1 => n19190, A2 => n19202, ZN => n2944);
   U7532 : OAI21_X1 port map( B1 => n8298, B2 => n8040, A => n1835, ZN => n5965
                           );
   U7533 : NOR2_X1 port map( A1 => n7455, A2 => n1835, ZN => n8514);
   U7534 : NAND2_X1 port map( A1 => n12385, A2 => n2946, ZN => n3530);
   U7535 : NOR2_X1 port map( A1 => n12382, A2 => n11915, ZN => n2946);
   U7536 : NAND2_X1 port map( A1 => n898, A2 => n11568, ZN => n11565);
   U7537 : NAND3_X1 port map( A1 => n20349, A2 => n18111, A3 => n18112, ZN => 
                           n2950);
   U7539 : INV_X1 port map( A => n16016, ZN => n15885);
   U7540 : INV_X1 port map( A => n16016, ZN => n3473);
   U7541 : XNOR2_X1 port map( A => n13082, B => n2953, ZN => n13083);
   U7542 : XNOR2_X1 port map( A => n12713, B => n2954, ZN => n2953);
   U7543 : OAI21_X1 port map( B1 => n8004, B2 => n8315, A => n281, ZN => n7593)
                           ;
   U7544 : NAND2_X1 port map( A1 => n19690, A2 => n17927, ZN => n17928);
   U7545 : OAI211_X2 port map( C1 => n5303, C2 => n5302, A => n5301, B => n2956
                           , ZN => n7338);
   U7546 : NAND2_X1 port map( A1 => n2958, A2 => n18568, ZN => n2957);
   U7547 : NOR2_X1 port map( A1 => n18555, A2 => n18565, ZN => n2958);
   U7548 : AND2_X2 port map( A1 => n2959, A2 => n16445, ZN => n18565);
   U7549 : OAI211_X1 port map( C1 => n1060, C2 => n16444, A => n16797, B => 
                           n16443, ZN => n2959);
   U7550 : INV_X1 port map( A => n7728, ZN => n8343);
   U7551 : INV_X1 port map( A => n8166, ZN => n8340);
   U7552 : NAND2_X1 port map( A1 => n2962, A2 => n8166, ZN => n2961);
   U7553 : OAI21_X1 port map( B1 => n7728, B2 => n2964, A => n20274, ZN => 
                           n2962);
   U7555 : INV_X1 port map( A => n8342, ZN => n2964);
   U7556 : NAND2_X1 port map( A1 => n2966, A2 => n2965, ZN => n19405);
   U7557 : NAND2_X1 port map( A1 => n16496, A2 => n2966, ZN => n16501);
   U7558 : NAND2_X1 port map( A1 => n17606, A2 => n19404, ZN => n2966);
   U7560 : XNOR2_X1 port map( A => n17002, B => n16555, ZN => n17141);
   U7563 : AOI22_X1 port map( A1 => n11158, A2 => n11157, B1 => n11156, B2 => 
                           n11155, ZN => n12037);
   U7564 : INV_X1 port map( A => n5069, ZN => n5072);
   U7565 : XNOR2_X2 port map( A => n3836, B => Key(89), ZN => n5069);
   U7566 : INV_X1 port map( A => n5071, ZN => n2971);
   U7567 : NAND2_X1 port map( A1 => n3824, A2 => n2973, ZN => n15414);
   U7568 : OAI21_X1 port map( B1 => n15412, B2 => n2973, A => n15411, ZN => 
                           n15415);
   U7569 : OAI21_X1 port map( B1 => n10855, B2 => n9883, A => n11230, ZN => 
                           n10873);
   U7571 : NAND2_X1 port map( A1 => n14898, A2 => n2974, ZN => n14900);
   U7572 : MUX2_X1 port map( A => n7958, B => n7956, S => n277, Z => n7962);
   U7573 : NAND2_X1 port map( A1 => n8906, A2 => n2976, ZN => n7959);
   U7574 : NAND2_X1 port map( A1 => n7915, A2 => n2975, ZN => n7839);
   U7575 : AND2_X1 port map( A1 => n7956, A2 => n2977, ZN => n2975);
   U7576 : OAI21_X1 port map( B1 => n7835, B2 => n7834, A => n2977, ZN => n7837
                           );
   U7577 : XNOR2_X1 port map( A => n7178, B => n2087, ZN => n6375);
   U7578 : NAND2_X1 port map( A1 => n14236, A2 => n19907, ZN => n2979);
   U7579 : XNOR2_X1 port map( A => n2980, B => n1228, ZN => Ciphertext(64));
   U7581 : AOI22_X1 port map( A1 => n19935, A2 => n18143, B1 => n18144, B2 => 
                           n19934, ZN => n2981);
   U7583 : NOR2_X1 port map( A1 => n2984, A2 => n9296, ZN => n3806);
   U7584 : INV_X1 port map( A => n9295, ZN => n2984);
   U7585 : NAND2_X1 port map( A1 => n2985, A2 => n8845, ZN => n7438);
   U7586 : OAI21_X1 port map( B1 => n20472, B2 => n3418, A => n9018, ZN => 
                           n8522);
   U7587 : NAND2_X1 port map( A1 => n995, A2 => n2987, ZN => n2986);
   U7588 : INV_X1 port map( A => n15379, ZN => n15163);
   U7589 : INV_X1 port map( A => n9158, ZN => n9160);
   U7590 : NAND2_X1 port map( A1 => n9159, A2 => n8696, ZN => n2989);
   U7591 : XNOR2_X1 port map( A => n16744, B => n2993, ZN => n2992);
   U7593 : OAI211_X1 port map( C1 => n3002, C2 => n3000, A => n2998, B => n2995
                           , ZN => Ciphertext(176));
   U7594 : NAND4_X1 port map( A1 => n2997, A2 => n17543, A3 => n2996, A4 => 
                           n17544, ZN => n2995);
   U7595 : INV_X1 port map( A => n3004, ZN => n2997);
   U7596 : NAND3_X1 port map( A1 => n2999, A2 => n3003, A3 => n298, ZN => n2998
                           );
   U7597 : INV_X1 port map( A => n17543, ZN => n2999);
   U7598 : NOR2_X1 port map( A1 => n3004, A2 => n3001, ZN => n3000);
   U7599 : OR2_X1 port map( A1 => n17542, A2 => n17544, ZN => n3001);
   U7600 : XNOR2_X1 port map( A => n3003, B => n17544, ZN => n3002);
   U7601 : NAND2_X1 port map( A1 => n19316, A2 => n19340, ZN => n3003);
   U7602 : OAI21_X1 port map( B1 => n19324, B2 => n19955, A => n17541, ZN => 
                           n3004);
   U7603 : NAND2_X1 port map( A1 => n14809, A2 => n19781, ZN => n3005);
   U7604 : NAND2_X1 port map( A1 => n3007, A2 => n8241, ZN => n8242);
   U7605 : INV_X1 port map( A => n7436, ZN => n3007);
   U7607 : NAND2_X1 port map( A1 => n16684, A2 => n17654, ZN => n17538);
   U7608 : AND2_X1 port map( A1 => n19388, A2 => n20004, ZN => n16684);
   U7609 : AND2_X1 port map( A1 => n3010, A2 => n6113, ZN => n6110);
   U7610 : NAND2_X1 port map( A1 => n4733, A2 => n4732, ZN => n3009);
   U7611 : NAND2_X1 port map( A1 => n3013, A2 => n3011, ZN => n12414);
   U7612 : NAND2_X1 port map( A1 => n12412, A2 => n3012, ZN => n3011);
   U7613 : NAND2_X1 port map( A1 => n12411, A2 => n12754, ZN => n3013);
   U7614 : INV_X1 port map( A => n11174, ZN => n3015);
   U7615 : AOI21_X1 port map( B1 => n11178, B2 => n3789, A => n3014, ZN => 
                           n3016);
   U7616 : OAI21_X1 port map( B1 => n11176, B2 => n11178, A => n3015, ZN => 
                           n3014);
   U7617 : MUX2_X1 port map( A => n3018, B => n11179, S => n9486, Z => n3017);
   U7618 : NOR2_X1 port map( A1 => n3015, A2 => n11177, ZN => n3018);
   U7619 : NAND2_X1 port map( A1 => n3019, A2 => n15504, ZN => n15820);
   U7620 : OAI21_X1 port map( B1 => n3019, B2 => n14069, A => n15822, ZN => 
                           n14072);
   U7621 : XNOR2_X1 port map( A => n3021, B => n6992, ZN => n3020);
   U7622 : XNOR2_X1 port map( A => n3022, B => n6991, ZN => n3021);
   U7623 : INV_X1 port map( A => n7333, ZN => n3022);
   U7625 : AOI22_X2 port map( A1 => n10660, A2 => n11952, B1 => n11828, B2 => 
                           n3024, ZN => n13192);
   U7626 : NAND2_X1 port map( A1 => n13927, A2 => n1364, ZN => n3025);
   U7627 : INV_X1 port map( A => n18868, ZN => n3028);
   U7628 : INV_X1 port map( A => n18868, ZN => n3031);
   U7630 : MUX2_X1 port map( A => n15873, B => n15872, S => n19514, Z => n15878
                           );
   U7631 : XNOR2_X1 port map( A => n3035, B => n1780, ZN => Ciphertext(129));
   U7632 : NAND3_X1 port map( A1 => n20214, A2 => n19109, A3 => n19094, ZN => 
                           n3036);
   U7633 : INV_X1 port map( A => n19089, ZN => n3038);
   U7634 : NAND3_X1 port map( A1 => n18358, A2 => n18341, A3 => n18344, ZN => 
                           n18349);
   U7635 : NAND2_X1 port map( A1 => n17236, A2 => n3461, ZN => n3039);
   U7636 : NAND2_X1 port map( A1 => n10103, A2 => n3040, ZN => n3629);
   U7637 : INV_X1 port map( A => n19949, ZN => n3040);
   U7638 : NAND2_X1 port map( A1 => n14979, A2 => n14978, ZN => n3041);
   U7639 : NAND2_X1 port map( A1 => n6206, A2 => n19492, ZN => n3044);
   U7640 : NAND2_X1 port map( A1 => n4473, A2 => n4472, ZN => n6205);
   U7641 : INV_X1 port map( A => n18442, ZN => n3045);
   U7642 : NAND2_X1 port map( A1 => n20139, A2 => n18467, ZN => n18442);
   U7645 : NAND2_X1 port map( A1 => n8925, A2 => n8748, ZN => n3433);
   U7646 : AOI22_X2 port map( A1 => n7405, A2 => n7948, B1 => n20367, B2 => 
                           n7404, ZN => n8748);
   U7647 : OR2_X2 port map( A1 => n14407, A2 => n3047, ZN => n15628);
   U7648 : NAND2_X1 port map( A1 => n937, A2 => n11278, ZN => n9546);
   U7649 : NAND2_X1 port map( A1 => n10729, A2 => n19913, ZN => n3052);
   U7650 : NOR2_X1 port map( A1 => n8193, A2 => n3054, ZN => n3053);
   U7651 : INV_X1 port map( A => n8193, ZN => n3055);
   U7652 : INV_X1 port map( A => n14714, ZN => n3057);
   U7653 : NAND2_X1 port map( A1 => n3057, A2 => n19843, ZN => n3056);
   U7654 : OAI21_X1 port map( B1 => n3058, B2 => n9238, A => n9233, ZN => n3060
                           );
   U7655 : XNOR2_X1 port map( A => n10319, B => n10029, ZN => n10035);
   U7656 : NAND2_X1 port map( A1 => n20464, A2 => n5046, ZN => n3061);
   U7658 : XNOR2_X1 port map( A => n13762, B => n13616, ZN => n13303);
   U7659 : MUX2_X1 port map( A => n14395, B => n14598, S => n14396, Z => n14398
                           );
   U7661 : NAND3_X1 port map( A1 => n18229, A2 => n18232, A3 => n3066, ZN => 
                           n3064);
   U7662 : NAND3_X1 port map( A1 => n19876, A2 => n18233, A3 => n3066, ZN => 
                           n3065);
   U7663 : NAND3_X1 port map( A1 => n1025, A2 => n3069, A3 => n3070, ZN => 
                           n3068);
   U7664 : NAND2_X1 port map( A1 => n5756, A2 => n287, ZN => n3069);
   U7665 : NAND2_X1 port map( A1 => n5757, A2 => n3071, ZN => n3070);
   U7667 : NAND2_X1 port map( A1 => n8000, A2 => n3074, ZN => n3073);
   U7669 : NAND3_X1 port map( A1 => n14439, A2 => n14442, A3 => n14441, ZN => 
                           n12928);
   U7670 : NAND2_X1 port map( A1 => n139, A2 => n14442, ZN => n3173);
   U7671 : INV_X1 port map( A => n4953, ZN => n3078);
   U7672 : INV_X1 port map( A => n4952, ZN => n4475);
   U7673 : OAI21_X1 port map( B1 => n4399, B2 => n3079, A => n4916, ZN => n4400
                           );
   U7674 : INV_X1 port map( A => n18467, ZN => n18461);
   U7675 : NAND2_X1 port map( A1 => n18465, A2 => n18467, ZN => n3512);
   U7676 : INV_X1 port map( A => n16469, ZN => n3081);
   U7677 : MUX2_X1 port map( A => n14338, B => n14335, S => n12879, Z => n12880
                           );
   U7679 : MUX2_X1 port map( A => n7948, B => n7949, S => n7479, Z => n7955);
   U7680 : NAND3_X1 port map( A1 => n3583, A2 => n7950, A3 => n20367, ZN => 
                           n3581);
   U7681 : INV_X1 port map( A => n16166, ZN => n17505);
   U7682 : NAND3_X1 port map( A1 => n5714, A2 => n3086, A3 => n5715, ZN => 
                           n5724);
   U7683 : NAND2_X1 port map( A1 => n14168, A2 => n14167, ZN => n3088);
   U7685 : NAND2_X1 port map( A1 => n7936, A2 => n7763, ZN => n7519);
   U7687 : XNOR2_X1 port map( A => n3092, B => n20126, ZN => n3091);
   U7688 : INV_X1 port map( A => n16900, ZN => n3092);
   U7689 : XNOR2_X1 port map( A => n16284, B => n16285, ZN => n3093);
   U7691 : OAI22_X1 port map( A1 => n3095, A2 => n4361, B1 => n4608, B2 => 
                           n4601, ZN => n3094);
   U7692 : NAND2_X1 port map( A1 => n3097, A2 => n3096, ZN => n6300);
   U7693 : INV_X1 port map( A => n6089, ZN => n5199);
   U7694 : AOI21_X1 port map( B1 => n6087, B2 => n20149, A => n6089, ZN => 
                           n3098);
   U7696 : INV_X1 port map( A => n12374, ZN => n12376);
   U7697 : OAI21_X1 port map( B1 => n11856, B2 => n12020, A => n3099, ZN => 
                           n11857);
   U7698 : NAND2_X1 port map( A1 => n3100, A2 => n12369, ZN => n3099);
   U7699 : NOR2_X1 port map( A1 => n19504, A2 => n12374, ZN => n3100);
   U7700 : INV_X1 port map( A => n10640, ZN => n11534);
   U7701 : NAND3_X1 port map( A1 => n11535, A2 => n11168, A3 => n11171, ZN => 
                           n3104);
   U7702 : INV_X1 port map( A => n10638, ZN => n11535);
   U7703 : NAND3_X1 port map( A1 => n10640, A2 => n11538, A3 => n11539, ZN => 
                           n3105);
   U7704 : NOR2_X1 port map( A1 => n11535, A2 => n10640, ZN => n11169);
   U7705 : NAND3_X1 port map( A1 => n20146, A2 => n9129, A3 => n9201, ZN => 
                           n3106);
   U7706 : NAND2_X1 port map( A1 => n8276, A2 => n9782, ZN => n3107);
   U7707 : OAI211_X2 port map( C1 => n8244, C2 => n3775, A => n8243, B => n8242
                           , ZN => n9201);
   U7709 : NOR2_X2 port map( A1 => n3113, A2 => n3111, ZN => n12001);
   U7710 : MUX2_X1 port map( A => n9486, B => n11176, S => n11174, Z => n3112);
   U7711 : MUX2_X1 port map( A => n9379, B => n9378, S => n2232, Z => n3113);
   U7712 : XNOR2_X2 port map( A => n9225, B => n9224, ZN => n11176);
   U7713 : INV_X1 port map( A => n17172, ZN => n17826);
   U7714 : NAND2_X1 port map( A1 => n17824, A2 => n17823, ZN => n3114);
   U7715 : INV_X1 port map( A => n17080, ZN => n17822);
   U7716 : NAND2_X1 port map( A1 => n17826, A2 => n17825, ZN => n3117);
   U7718 : AOI22_X1 port map( A1 => n8343, A2 => n2964, B1 => n8166, B2 => 
                           n8344, ZN => n3118);
   U7719 : NAND2_X1 port map( A1 => n3121, A2 => n20274, ZN => n3119);
   U7721 : XNOR2_X1 port map( A => n6946, B => n6945, ZN => n6948);
   U7722 : NAND3_X2 port map( A1 => n3124, A2 => n5281, A3 => n3123, ZN => 
                           n6945);
   U7723 : NAND2_X1 port map( A1 => n3125, A2 => n3128, ZN => n3123);
   U7724 : NAND2_X1 port map( A1 => n3125, A2 => n3126, ZN => n3124);
   U7725 : OR2_X1 port map( A1 => n5280, A2 => n3127, ZN => n3126);
   U7726 : NAND2_X1 port map( A1 => n5282, A2 => n3127, ZN => n3125);
   U7727 : INV_X1 port map( A => n5424, ZN => n3127);
   U7728 : NAND2_X1 port map( A1 => n3130, A2 => n4754, ZN => n3129);
   U7729 : NOR2_X1 port map( A1 => n4565, A2 => n3131, ZN => n3130);
   U7730 : INV_X1 port map( A => n4567, ZN => n3131);
   U7731 : NAND2_X1 port map( A1 => n5518, A2 => n5929, ZN => n3371);
   U7732 : NAND2_X1 port map( A1 => n5053, A2 => n20461, ZN => n3132);
   U7733 : NAND2_X1 port map( A1 => n204, A2 => n11076, ZN => n3133);
   U7734 : NAND2_X1 port map( A1 => n11476, A2 => n3471, ZN => n3134);
   U7735 : NAND3_X1 port map( A1 => n3138, A2 => n15702, A3 => n15696, ZN => 
                           n3137);
   U7736 : NOR2_X1 port map( A1 => n3141, A2 => n3140, ZN => n3139);
   U7737 : NOR2_X1 port map( A1 => n16779, A2 => n19144, ZN => n3140);
   U7739 : NAND2_X1 port map( A1 => n19147, A2 => n19145, ZN => n3143);
   U7742 : NAND2_X1 port map( A1 => n3148, A2 => n14905, ZN => n3146);
   U7743 : NAND3_X1 port map( A1 => n14903, A2 => n15056, A3 => n15413, ZN => 
                           n3147);
   U7744 : INV_X1 port map( A => n14312, ZN => n15549);
   U7745 : NOR2_X1 port map( A1 => n15413, A2 => n15553, ZN => n3148);
   U7746 : INV_X1 port map( A => n14236, ZN => n14114);
   U7747 : NAND2_X1 port map( A1 => n5659, A2 => n6113, ZN => n5660);
   U7748 : NAND2_X1 port map( A1 => n3150, A2 => n17835, ZN => n17844);
   U7749 : NAND2_X1 port map( A1 => n3150, A2 => n3755, ZN => n3285);
   U7750 : NAND2_X1 port map( A1 => n3558, A2 => n11572, ZN => n3151);
   U7751 : NOR2_X1 port map( A1 => n12299, A2 => n12273, ZN => n12033);
   U7752 : OAI21_X1 port map( B1 => n14747, B2 => n1936, A => n3158, ZN => 
                           n13934);
   U7753 : OAI211_X1 port map( C1 => n14427, C2 => n1936, A => n14747, B => 
                           n3158, ZN => n14428);
   U7754 : INV_X1 port map( A => n14747, ZN => n3156);
   U7755 : NAND2_X1 port map( A1 => n14752, A2 => n3157, ZN => n15189);
   U7756 : OR2_X1 port map( A1 => n14753, A2 => n3158, ZN => n3157);
   U7757 : XNOR2_X1 port map( A => n3159, B => n875, ZN => n13474);
   U7758 : XNOR2_X1 port map( A => n3159, B => n18691, ZN => n13360);
   U7759 : XNOR2_X1 port map( A => n3159, B => n538, ZN => n13824);
   U7760 : XNOR2_X1 port map( A => n3159, B => n19467, ZN => n12540);
   U7761 : XNOR2_X1 port map( A => n13368, B => n3159, ZN => n13530);
   U7762 : NAND2_X1 port map( A1 => n11117, A2 => n11435, ZN => n3161);
   U7763 : XNOR2_X1 port map( A => n3162, B => n16019, ZN => n16020);
   U7764 : XNOR2_X1 port map( A => n17406, B => n3162, ZN => n16908);
   U7765 : XNOR2_X1 port map( A => n16770, B => n3162, ZN => n16829);
   U7766 : OAI211_X2 port map( C1 => n15085, C2 => n15086, A => n15084, B => 
                           n15083, ZN => n3162);
   U7767 : NAND2_X1 port map( A1 => n12295, A2 => n3164, ZN => n12163);
   U7768 : MUX2_X1 port map( A => n12534, B => n12531, S => n924, Z => n11772);
   U7769 : INV_X1 port map( A => n3166, ZN => n3165);
   U7770 : NAND2_X1 port map( A1 => n5105, A2 => n5099, ZN => n4792);
   U7771 : NAND2_X1 port map( A1 => n5102, A2 => n5107, ZN => n3598);
   U7772 : NAND2_X1 port map( A1 => n12813, A2 => n11803, ZN => n3171);
   U7773 : OAI211_X1 port map( C1 => n12813, C2 => n19626, A => n3169, B => 
                           n3168, ZN => n12119);
   U7775 : XNOR2_X1 port map( A => n3171, B => n2151, ZN => n13699);
   U7776 : XNOR2_X1 port map( A => n3171, B => n18716, ZN => n11817);
   U7777 : XNOR2_X1 port map( A => n13588, B => n3171, ZN => n12894);
   U7778 : OAI211_X2 port map( C1 => n3177, C2 => n11005, A => n3176, B => 
                           n3175, ZN => n11952);
   U7779 : MUX2_X1 port map( A => n937, B => n19736, S => n9547, Z => n3177);
   U7780 : NAND2_X1 port map( A1 => n14053, A2 => n14422, ZN => n3178);
   U7781 : NAND2_X1 port map( A1 => n2039, A2 => n14359, ZN => n14358);
   U7782 : INV_X1 port map( A => n6345, ZN => n3181);
   U7783 : INV_X1 port map( A => n6345, ZN => n7743);
   U7784 : AOI22_X1 port map( A1 => n3182, A2 => n7741, B1 => n6900, B2 => 
                           n8355, ZN => n6901);
   U7785 : XNOR2_X1 port map( A => n10280, B => n17095, ZN => n3184);
   U7786 : NOR2_X1 port map( A1 => n8697, A2 => n9161, ZN => n3183);
   U7787 : NAND2_X1 port map( A1 => n8698, A2 => n8697, ZN => n3185);
   U7788 : NOR2_X1 port map( A1 => n12103, A2 => n12101, ZN => n3186);
   U7789 : NAND2_X1 port map( A1 => n3449, A2 => n3189, ZN => n3188);
   U7791 : OAI21_X1 port map( B1 => n6148, B2 => n6138, A => n3187, ZN => n5266
                           );
   U7792 : NAND2_X1 port map( A1 => n6138, A2 => n5859, ZN => n3187);
   U7793 : NAND2_X1 port map( A1 => n5616, A2 => n3188, ZN => n5617);
   U7795 : NAND2_X1 port map( A1 => n14176, A2 => n12725, ZN => n3190);
   U7797 : XNOR2_X2 port map( A => Key(101), B => Plaintext(101), ZN => n5080);
   U7798 : NAND2_X1 port map( A1 => n4459, A2 => n5078, ZN => n3450);
   U7800 : NAND3_X1 port map( A1 => n4671, A2 => n4669, A3 => n4670, ZN => 
                           n3192);
   U7801 : NAND2_X1 port map( A1 => n4824, A2 => n4827, ZN => n4670);
   U7802 : XNOR2_X2 port map( A => Key(73), B => Plaintext(73), ZN => n4827);
   U7803 : NAND2_X1 port map( A1 => n3197, A2 => n3195, ZN => n3194);
   U7804 : NAND2_X1 port map( A1 => n3196, A2 => n6184, ZN => n3195);
   U7805 : OAI21_X1 port map( B1 => n6380, B2 => n19476, A => n2865, ZN => 
                           n3197);
   U7806 : NAND2_X1 port map( A1 => n3198, A2 => n20270, ZN => n8020);
   U7807 : NAND2_X1 port map( A1 => n208, A2 => n3198, ZN => n7812);
   U7808 : INV_X1 port map( A => n7801, ZN => n3198);
   U7809 : NAND2_X1 port map( A1 => n8927, A2 => n8928, ZN => n3199);
   U7810 : NAND2_X1 port map( A1 => n8926, A2 => n8925, ZN => n3200);
   U7811 : NAND2_X1 port map( A1 => n5035, A2 => n3203, ZN => n5036);
   U7812 : NAND2_X1 port map( A1 => n4771, A2 => n3203, ZN => n4772);
   U7813 : NAND2_X1 port map( A1 => n4770, A2 => n3203, ZN => n4774);
   U7814 : XNOR2_X1 port map( A => n17266, B => n17265, ZN => n18038);
   U7815 : NAND2_X1 port map( A1 => n3205, A2 => n18038, ZN => n18237);
   U7816 : INV_X1 port map( A => n17303, ZN => n17753);
   U7819 : OAI211_X1 port map( C1 => n630, C2 => n3198, A => n3212, B => n3211,
                           ZN => n3210);
   U7820 : INV_X1 port map( A => n7466, ZN => n3212);
   U7821 : OAI22_X1 port map( A1 => n16260, A2 => n19947, B1 => n17663, B2 => 
                           n3216, ZN => n3215);
   U7824 : NOR2_X1 port map( A1 => n8323, A2 => n3809, ZN => n3220);
   U7827 : OAI211_X1 port map( C1 => n19496, C2 => n14828, A => n3224, B => 
                           n3223, ZN => n3222);
   U7828 : NAND2_X1 port map( A1 => n14828, A2 => n14827, ZN => n3224);
   U7829 : NAND2_X1 port map( A1 => n3225, A2 => n14203, ZN => n14609);
   U7830 : INV_X1 port map( A => n14012, ZN => n3225);
   U7831 : NAND2_X1 port map( A1 => n3226, A2 => n14611, ZN => n14616);
   U7832 : OAI21_X2 port map( B1 => n3228, B2 => n5564, A => n4993, ZN => n7371
                           );
   U7833 : MUX2_X1 port map( A => n5532, B => n6033, S => n5531, Z => n3228);
   U7834 : NAND2_X1 port map( A1 => n4136, A2 => n4960, ZN => n3230);
   U7837 : AND4_X2 port map( A1 => n3241, A2 => n3240, A3 => n3239, A4 => n3238
                           , ZN => n13795);
   U7838 : OR2_X1 port map( A1 => n12175, A2 => n19768, ZN => n3238);
   U7839 : INV_X1 port map( A => n8014, ZN => n7826);
   U7842 : AOI21_X1 port map( B1 => n7829, B2 => n7991, A => n8014, ZN => n3243
                           );
   U7844 : NAND2_X1 port map( A1 => n13008, A2 => n3246, ZN => n3245);
   U7846 : NAND2_X1 port map( A1 => n18762, A2 => n18774, ZN => n18255);
   U7847 : NAND2_X1 port map( A1 => n18250, A2 => n18249, ZN => n3248);
   U7848 : NAND2_X1 port map( A1 => n3249, A2 => n906, ZN => n3867);
   U7849 : NAND2_X1 port map( A1 => n8139, A2 => n8352, ZN => n3251);
   U7850 : INV_X1 port map( A => n13921, ZN => n3252);
   U7853 : INV_X1 port map( A => n11792, ZN => n3256);
   U7854 : NAND2_X1 port map( A1 => n3258, A2 => n3257, ZN => n5846);
   U7855 : NAND2_X1 port map( A1 => n4695, A2 => n3259, ZN => n3257);
   U7856 : NAND2_X1 port map( A1 => n4694, A2 => n5107, ZN => n3258);
   U7857 : NOR2_X1 port map( A1 => n12155, A2 => n3260, ZN => n11908);
   U7858 : NAND2_X1 port map( A1 => n12315, A2 => n3260, ZN => n11712);
   U7860 : OAI21_X1 port map( B1 => n8295, B2 => n7789, A => n7454, ZN => n3261
                           );
   U7861 : NOR2_X1 port map( A1 => n8676, A2 => n8513, ZN => n8516);
   U7862 : XNOR2_X1 port map( A => n10125, B => n10356, ZN => n10130);
   U7863 : NAND3_X1 port map( A1 => n3262, A2 => n5697, A3 => n5522, ZN => 
                           n5523);
   U7864 : NAND2_X1 port map( A1 => n3264, A2 => n3263, ZN => n3262);
   U7865 : NAND2_X1 port map( A1 => n4950, A2 => n4142, ZN => n3263);
   U7866 : NAND2_X1 port map( A1 => n4143, A2 => n3265, ZN => n3264);
   U7867 : NAND2_X1 port map( A1 => n14165, A2 => n14427, ZN => n3266);
   U7868 : NAND2_X1 port map( A1 => n14166, A2 => n14424, ZN => n3268);
   U7869 : INV_X1 port map( A => n12607, ZN => n3269);
   U7870 : XNOR2_X1 port map( A => n12713, B => n18660, ZN => n13392);
   U7871 : NAND3_X1 port map( A1 => n3271, A2 => n280, A3 => n274, ZN => n3270)
                           ;
   U7872 : XNOR2_X2 port map( A => n6282, B => n6281, ZN => n7754);
   U7873 : XNOR2_X1 port map( A => n17377, B => n3273, ZN => n16918);
   U7874 : NAND2_X1 port map( A1 => n14200, A2 => n14590, ZN => n3275);
   U7875 : NAND2_X1 port map( A1 => n11656, A2 => n19768, ZN => n3277);
   U7876 : NAND2_X1 port map( A1 => n14807, A2 => n14813, ZN => n14196);
   U7877 : NAND2_X1 port map( A1 => n12354, A2 => n19768, ZN => n3537);
   U7878 : NAND3_X1 port map( A1 => n3282, A2 => n16734, A3 => n3287, ZN => 
                           n3284);
   U7879 : INV_X1 port map( A => n16730, ZN => n3282);
   U7881 : NAND2_X1 port map( A1 => n3286, A2 => n3284, ZN => n19151);
   U7882 : NAND2_X1 port map( A1 => n16734, A2 => n20423, ZN => n3286);
   U7883 : XNOR2_X1 port map( A => n19760, B => n10445, ZN => n6657);
   U7884 : NAND2_X1 port map( A1 => n3290, A2 => n5035, ZN => n3289);
   U7885 : NAND2_X1 port map( A1 => n3431, A2 => n16128, ZN => n3291);
   U7886 : NAND2_X1 port map( A1 => n15611, A2 => n3291, ZN => n16932);
   U7887 : OAI21_X1 port map( B1 => n9275, B2 => n9278, A => n9272, ZN => n8759
                           );
   U7888 : INV_X1 port map( A => n19144, ZN => n18337);
   U7891 : AND2_X1 port map( A1 => n12429, A2 => n12686, ZN => n12094);
   U7892 : NAND2_X1 port map( A1 => n10718, A2 => n11474, ZN => n3296);
   U7893 : XNOR2_X1 port map( A => n9902, B => n10579, ZN => n8740);
   U7894 : NAND2_X1 port map( A1 => n8731, A2 => n8730, ZN => n3297);
   U7895 : NAND2_X1 port map( A1 => n8732, A2 => n8941, ZN => n3298);
   U7896 : NAND2_X1 port map( A1 => n3301, A2 => n3300, ZN => n12039);
   U7897 : NAND2_X1 port map( A1 => n11169, A2 => n19915, ZN => n3300);
   U7898 : OAI21_X1 port map( B1 => n3303, B2 => n11171, A => n3302, ZN => 
                           n3301);
   U7899 : NAND2_X1 port map( A1 => n3304, A2 => n11171, ZN => n3302);
   U7900 : NOR2_X1 port map( A1 => n11170, A2 => n11168, ZN => n3303);
   U7901 : NAND2_X1 port map( A1 => n11534, A2 => n11170, ZN => n3304);
   U7902 : NAND2_X1 port map( A1 => n3305, A2 => n12237, ZN => n12073);
   U7904 : MUX2_X1 port map( A => n12604, B => n12605, S => n12610, Z => n12613
                           );
   U7905 : XNOR2_X2 port map( A => n12909, B => n12908, ZN => n14442);
   U7906 : NAND2_X1 port map( A1 => n14440, A2 => n14441, ZN => n3306);
   U7907 : NAND3_X1 port map( A1 => n15294, A2 => n15295, A3 => n15109, ZN => 
                           n3308);
   U7908 : OAI211_X2 port map( C1 => n5029, C2 => n5028, A => n3310, B => n3309
                           , ZN => n5927);
   U7909 : NAND3_X1 port map( A1 => n5029, A2 => n5026, A3 => n5025, ZN => 
                           n3310);
   U7910 : NAND2_X1 port map( A1 => n14962, A2 => n3315, ZN => n3314);
   U7911 : INV_X1 port map( A => n15581, ZN => n3315);
   U7912 : NAND2_X1 port map( A1 => n5320, A2 => n3319, ZN => n3318);
   U7913 : INV_X1 port map( A => n5320, ZN => n6070);
   U7914 : NAND2_X1 port map( A1 => n3317, A2 => n5978, ZN => n3316);
   U7915 : NAND2_X1 port map( A1 => n3319, A2 => n6072, ZN => n3317);
   U7916 : AOI21_X1 port map( B1 => n4421, B2 => n20105, A => n3977, ZN => 
                           n3320);
   U7917 : XNOR2_X1 port map( A => n6506, B => n6505, ZN => n3321);
   U7919 : NAND2_X1 port map( A1 => n15617, A2 => n15071, ZN => n14892);
   U7920 : INV_X1 port map( A => n5692, ZN => n4275);
   U7921 : AOI21_X1 port map( B1 => n4254, B2 => n4348, A => n4349, ZN => n3322
                           );
   U7922 : AOI21_X1 port map( B1 => n4256, B2 => n4255, A => n4540, ZN => n3323
                           );
   U7923 : AOI21_X1 port map( B1 => n9884, B2 => n11235, A => n9883, ZN => 
                           n3326);
   U7924 : MUX2_X1 port map( A => n12505, B => n12508, S => n12506, Z => n3565)
                           ;
   U7925 : NAND2_X1 port map( A1 => n9659, A2 => n1330, ZN => n3324);
   U7926 : NOR2_X1 port map( A1 => n12359, A2 => n12509, ZN => n12505);
   U7927 : NOR2_X2 port map( A1 => n3327, A2 => n3326, ZN => n12509);
   U7928 : NAND2_X1 port map( A1 => n9875, A2 => n10818, ZN => n3328);
   U7929 : OAI21_X1 port map( B1 => n14341, B2 => n14339, A => n3333, ZN => 
                           n3332);
   U7930 : NAND2_X1 port map( A1 => n14334, A2 => n19485, ZN => n3333);
   U7932 : NOR2_X1 port map( A1 => n3335, A2 => n7762, ZN => n3334);
   U7933 : NOR2_X1 port map( A1 => n7934, A2 => n7760, ZN => n3335);
   U7935 : MUX2_X1 port map( A => n7765, B => n3337, S => n7932, Z => n3336);
   U7936 : NAND2_X1 port map( A1 => n7934, A2 => n2540, ZN => n3337);
   U7937 : INV_X1 port map( A => n7763, ZN => n7934);
   U7938 : NAND3_X1 port map( A1 => n3339, A2 => n19240, A3 => n3338, ZN => 
                           n19245);
   U7939 : NAND2_X1 port map( A1 => n3340, A2 => n19236, ZN => n3339);
   U7940 : NAND2_X1 port map( A1 => n3341, A2 => n19234, ZN => n3340);
   U7941 : OR2_X1 port map( A1 => n19237, A2 => n19235, ZN => n3341);
   U7942 : NAND2_X1 port map( A1 => n19227, A2 => n19237, ZN => n19234);
   U7943 : OAI22_X2 port map( A1 => n5694, A2 => n5695, B1 => n5693, B2 => 
                           n4275, ZN => n7097);
   U7947 : NAND3_X1 port map( A1 => n16801, A2 => n17489, A3 => n19675, ZN => 
                           n3346);
   U7949 : OAI21_X1 port map( B1 => n1458, B2 => n15052, A => n15350, ZN => 
                           n3348);
   U7951 : OR2_X1 port map( A1 => n4538, A2 => n4539, ZN => n3349);
   U7952 : NAND2_X1 port map( A1 => n3933, A2 => n3932, ZN => n3350);
   U7954 : XNOR2_X1 port map( A => n13440, B => n3352, ZN => n11852);
   U7955 : INV_X1 port map( A => n12993, ZN => n3352);
   U7956 : XNOR2_X1 port map( A => n3353, B => n12993, ZN => n12858);
   U7957 : INV_X1 port map( A => n13078, ZN => n3353);
   U7958 : OAI21_X1 port map( B1 => n3356, B2 => n9255, A => n9252, ZN => n3355
                           );
   U7960 : NAND2_X1 port map( A1 => n11176, A2 => n10912, ZN => n3358);
   U7963 : INV_X1 port map( A => n11177, ZN => n3362);
   U7964 : XNOR2_X1 port map( A => n13569, B => n13134, ZN => n3363);
   U7965 : AND2_X1 port map( A1 => n18489, A2 => n18498, ZN => n17911);
   U7966 : NAND2_X1 port map( A1 => n16166, A2 => n17501, ZN => n16797);
   U7967 : NAND2_X1 port map( A1 => n13166, A2 => n3366, ZN => n13179);
   U7968 : NAND2_X1 port map( A1 => n14665, A2 => n14664, ZN => n3367);
   U7969 : NAND2_X1 port map( A1 => n3369, A2 => n3445, ZN => n3368);
   U7970 : OAI21_X1 port map( B1 => n7748, B2 => n7750, A => n3370, ZN => n3369
                           );
   U7971 : NAND2_X1 port map( A1 => n7749, A2 => n7748, ZN => n3370);
   U7972 : NAND2_X1 port map( A1 => n3948, A2 => n4539, ZN => n4200);
   U7973 : OAI21_X1 port map( B1 => n4350, B2 => n4199, A => n3948, ZN => n3949
                           );
   U7974 : MUX2_X1 port map( A => n4541, B => n3948, S => n4350, Z => n4203);
   U7975 : NAND3_X1 port map( A1 => n4536, A2 => n3948, A3 => n4350, ZN => 
                           n4351);
   U7976 : INV_X1 port map( A => n3373, ZN => n14262);
   U7977 : NOR2_X1 port map( A1 => n13981, A2 => n3373, ZN => n14539);
   U7980 : NOR2_X1 port map( A1 => n7979, A2 => n7921, ZN => n3375);
   U7981 : NAND2_X1 port map( A1 => n7984, A2 => n7981, ZN => n7979);
   U7983 : INV_X1 port map( A => n7921, ZN => n7768);
   U7984 : NAND2_X1 port map( A1 => n7768, A2 => n7978, ZN => n3376);
   U7987 : AND2_X2 port map( A1 => n3380, A2 => n3378, ZN => n10350);
   U7988 : NAND2_X1 port map( A1 => n9050, A2 => n3379, ZN => n3378);
   U7989 : NAND3_X1 port map( A1 => n3395, A2 => n9579, A3 => n3394, ZN => 
                           n3379);
   U7990 : NAND2_X1 port map( A1 => n9052, A2 => n9051, ZN => n3380);
   U7991 : OAI22_X1 port map( A1 => n19519, A2 => n9579, B1 => n8577, B2 => 
                           n19715, ZN => n9052);
   U7992 : NAND2_X1 port map( A1 => n11013, A2 => n3382, ZN => n3381);
   U7993 : OAI22_X1 port map( A1 => n4187, A2 => n4520, B1 => n4343, B2 => 
                           n4524, ZN => n3943);
   U7994 : XNOR2_X2 port map( A => Key(173), B => Plaintext(173), ZN => n4524);
   U7996 : NAND2_X1 port map( A1 => n3387, A2 => n7974, ZN => n3383);
   U7997 : MUX2_X1 port map( A => n278, B => n7922, S => n7967, Z => n3387);
   U7998 : NAND2_X1 port map( A1 => n17222, A2 => n3389, ZN => n3388);
   U7999 : NAND2_X1 port map( A1 => n17219, A2 => n1897, ZN => n3390);
   U8000 : INV_X1 port map( A => n15767, ZN => n15656);
   U8001 : OR2_X2 port map( A1 => n14856, A2 => n11594, ZN => n15767);
   U8003 : NOR2_X1 port map( A1 => n15657, A2 => n15767, ZN => n3393);
   U8005 : AND2_X1 port map( A1 => n13905, A2 => n14782, ZN => n11320);
   U8006 : AND2_X1 port map( A1 => n3397, A2 => n5279, ZN => n5672);
   U8007 : INV_X1 port map( A => n5668, ZN => n3397);
   U8008 : NAND3_X1 port map( A1 => n3398, A2 => n5670, A3 => n5668, ZN => 
                           n5281);
   U8009 : MUX2_X1 port map( A => n3398, B => n5669, S => n5670, Z => n5426);
   U8010 : OAI21_X1 port map( B1 => n5673, B2 => n3398, A => n5670, ZN => n5187
                           );
   U8011 : NAND2_X1 port map( A1 => n4209, A2 => n4208, ZN => n3399);
   U8012 : NAND2_X1 port map( A1 => n12630, A2 => n3401, ZN => n3400);
   U8014 : INV_X1 port map( A => n12630, ZN => n3403);
   U8015 : AOI21_X2 port map( B1 => n8294, B2 => n8293, A => n3406, ZN => n9106
                           );
   U8016 : XNOR2_X1 port map( A => n16707, B => n17143, ZN => n16822);
   U8018 : INV_X1 port map( A => n3408, ZN => n3407);
   U8019 : OAI21_X1 port map( B1 => n6028, B2 => n3410, A => n3409, ZN => n3408
                           );
   U8021 : NAND2_X1 port map( A1 => n3434, A2 => n19790, ZN => n6028);
   U8022 : NAND2_X1 port map( A1 => n16802, A2 => n17492, ZN => n16803);
   U8023 : NAND2_X1 port map( A1 => n16471, A2 => n17492, ZN => n16472);
   U8024 : NAND2_X1 port map( A1 => n7416, A2 => n3525, ZN => n3524);
   U8025 : NAND2_X1 port map( A1 => n3694, A2 => n14562, ZN => n3412);
   U8026 : OAI21_X2 port map( B1 => n14123, B2 => n14122, A => n14121, ZN => 
                           n15608);
   U8027 : NAND2_X1 port map( A1 => n3427, A2 => n997, ZN => n3413);
   U8028 : MUX2_X1 port map( A => n3431, B => n16127, S => n16128, Z => n3415);
   U8029 : XNOR2_X1 port map( A => n10558, B => n10430, ZN => n10242);
   U8031 : NAND2_X1 port map( A1 => n3418, A2 => n9020, ZN => n3416);
   U8032 : NAND3_X1 port map( A1 => n9019, A2 => n9296, A3 => n20159, ZN => 
                           n3417);
   U8033 : XNOR2_X1 port map( A => n13649, B => n3420, ZN => n3419);
   U8034 : INV_X1 port map( A => n13650, ZN => n3420);
   U8035 : NAND3_X1 port map( A1 => n17646, A2 => n3422, A3 => n17647, ZN => 
                           n3421);
   U8036 : NAND2_X1 port map( A1 => n3423, A2 => n17737, ZN => n3422);
   U8037 : NAND2_X1 port map( A1 => n17645, A2 => n17644, ZN => n3423);
   U8038 : XNOR2_X1 port map( A => n10125, B => n3424, ZN => n10412);
   U8039 : NAND2_X1 port map( A1 => n3427, A2 => n3425, ZN => n3426);
   U8040 : OAI21_X1 port map( B1 => n8925, B2 => n8932, A => n3433, ZN => n8754
                           );
   U8044 : NAND3_X1 port map( A1 => n19735, A2 => n18672, A3 => n18666, ZN => 
                           n3436);
   U8045 : NAND3_X1 port map( A1 => n18686, A2 => n19735, A3 => n18671, ZN => 
                           n3437);
   U8047 : NAND2_X1 port map( A1 => n13891, A2 => n3440, ZN => n13892);
   U8048 : NAND3_X1 port map( A1 => n20500, A2 => n14800, A3 => n3440, ZN => 
                           n14802);
   U8049 : OAI22_X1 port map( A1 => n12321, A2 => n3439, B1 => n14797, B2 => 
                           n3440, ZN => n14851);
   U8050 : INV_X1 port map( A => n14801, ZN => n3439);
   U8051 : NAND2_X1 port map( A1 => n11282, A2 => n19779, ZN => n9413);
   U8052 : MUX2_X1 port map( A => n4746, B => n4744, S => n4204, Z => n4751);
   U8053 : NAND2_X1 port map( A1 => n4559, A2 => n4204, ZN => n4250);
   U8054 : MUX2_X1 port map( A => n11881, B => n11048, S => n11880, Z => n11049
                           );
   U8055 : MUX2_X1 port map( A => n11460, B => n11461, S => n11880, Z => n11462
                           );
   U8056 : NAND2_X1 port map( A1 => n14819, A2 => n3444, ZN => n3443);
   U8057 : MUX2_X1 port map( A => n7749, B => n7748, S => n7508, Z => n3447);
   U8058 : XNOR2_X1 port map( A => n3448, B => n16067, ZN => n16068);
   U8059 : XNOR2_X1 port map( A => n16860, B => n3448, ZN => n16765);
   U8060 : XNOR2_X1 port map( A => n16214, B => n3448, ZN => n15855);
   U8061 : OR2_X1 port map( A1 => n15636, A2 => n15846, ZN => n15848);
   U8062 : NAND2_X1 port map( A1 => n3450, A2 => n5077, ZN => n3449);
   U8064 : AOI21_X1 port map( B1 => n20111, B2 => n20361, A => n18384, ZN => 
                           n3456);
   U8066 : INV_X1 port map( A => n15768, ZN => n3457);
   U8067 : OAI21_X1 port map( B1 => n4520, B2 => n4524, A => n4519, ZN => n4521
                           );
   U8070 : NAND2_X1 port map( A1 => n3461, A2 => n19374, ZN => n17598);
   U8071 : OAI22_X1 port map( A1 => n19647, A2 => n19372, B1 => n19380, B2 => 
                           n19666, ZN => n3461);
   U8072 : OAI21_X1 port map( B1 => n3463, B2 => n3462, A => n11757, ZN => 
                           n3464);
   U8073 : INV_X1 port map( A => n12306, ZN => n3463);
   U8074 : INV_X1 port map( A => n9771, ZN => n10298);
   U8075 : NAND2_X1 port map( A1 => n8791, A2 => n9149, ZN => n3465);
   U8076 : NAND2_X1 port map( A1 => n8792, A2 => n8338, ZN => n3466);
   U8077 : NAND2_X1 port map( A1 => n3470, A2 => n5993, ZN => n3469);
   U8078 : NAND2_X1 port map( A1 => n5088, A2 => n5083, ZN => n4090);
   U8079 : NAND3_X1 port map( A1 => n4802, A2 => n5088, A3 => n19777, ZN => 
                           n4700);
   U8080 : NAND3_X1 port map( A1 => n4807, A2 => n5088, A3 => n4804, ZN => 
                           n4805);
   U8081 : INV_X1 port map( A => n8192, ZN => n8051);
   U8083 : NAND2_X1 port map( A1 => n8053, A2 => n8192, ZN => n3472);
   U8084 : XNOR2_X1 port map( A => n6116, B => n6115, ZN => n7457);
   U8085 : AND2_X1 port map( A1 => n15333, A2 => n3473, ZN => n15706);
   U8086 : NAND2_X1 port map( A1 => n2475, A2 => n3475, ZN => n18127);
   U8087 : NAND2_X1 port map( A1 => n17945, A2 => n3475, ZN => n17952);
   U8088 : AND2_X1 port map( A1 => n12532, A2 => n12534, ZN => n3477);
   U8089 : NAND2_X1 port map( A1 => n11477, A2 => n3481, ZN => n3478);
   U8090 : NAND2_X1 port map( A1 => n11478, A2 => n3482, ZN => n3479);
   U8091 : NAND2_X1 port map( A1 => n3483, A2 => n6120, ZN => n5390);
   U8092 : NAND3_X1 port map( A1 => n6128, A2 => n5868, A3 => n3483, ZN => 
                           n4433);
   U8093 : AND2_X1 port map( A1 => n3484, A2 => n20252, ZN => n8146);
   U8094 : NAND2_X1 port map( A1 => n3484, A2 => n7671, ZN => n8371);
   U8095 : NOR2_X1 port map( A1 => n3484, A2 => n20252, ZN => n6750);
   U8097 : NAND2_X1 port map( A1 => n7677, A2 => n3491, ZN => n8722);
   U8099 : NAND2_X1 port map( A1 => n9359, A2 => n3493, ZN => n3492);
   U8100 : MUX2_X1 port map( A => n9358, B => n8904, S => n9359, Z => n3494);
   U8101 : NAND2_X1 port map( A1 => n9352, A2 => n9358, ZN => n3495);
   U8102 : INV_X1 port map( A => n6786, ZN => n6511);
   U8103 : XNOR2_X2 port map( A => Key(68), B => Plaintext(68), ZN => n3978);
   U8104 : INV_X1 port map( A => n13617, ZN => n3498);
   U8105 : OR2_X1 port map( A1 => n11315, A2 => n12409, ZN => n3499);
   U8106 : INV_X1 port map( A => n10746, ZN => n3500);
   U8107 : XNOR2_X1 port map( A => n856, B => n10296, ZN => n10406);
   U8109 : NAND2_X1 port map( A1 => n9211, A2 => n9135, ZN => n3503);
   U8112 : NAND3_X1 port map( A1 => n8923, A2 => n3506, A3 => n3505, ZN => 
                           n3504);
   U8113 : NAND2_X1 port map( A1 => n8733, A2 => n8734, ZN => n3505);
   U8114 : NAND2_X1 port map( A1 => n8916, A2 => n8497, ZN => n3506);
   U8116 : AND2_X1 port map( A1 => n204, A2 => n3711, ZN => n9913);
   U8117 : NAND2_X1 port map( A1 => n11476, A2 => n3507, ZN => n9920);
   U8118 : NAND2_X1 port map( A1 => n204, A2 => n3507, ZN => n10717);
   U8119 : NOR2_X1 port map( A1 => n204, A2 => n3507, ZN => n10894);
   U8120 : OAI21_X1 port map( B1 => n3711, B2 => n11474, A => n3508, ZN => 
                           n11478);
   U8121 : NAND2_X1 port map( A1 => n11474, A2 => n11475, ZN => n3508);
   U8122 : NAND2_X1 port map( A1 => n3509, A2 => n18436, ZN => n16486);
   U8123 : NAND2_X1 port map( A1 => n3512, A2 => n3510, ZN => n3509);
   U8124 : NAND2_X1 port map( A1 => n18453, A2 => n20231, ZN => n3510);
   U8125 : NAND3_X1 port map( A1 => n14574, A2 => n14267, A3 => n14570, ZN => 
                           n14272);
   U8126 : OAI21_X1 port map( B1 => n12430, B2 => n12686, A => n3514, ZN => 
                           n11613);
   U8127 : MUX2_X1 port map( A => n11142, B => n11144, S => n9616, Z => n10958)
                           ;
   U8128 : MUX2_X1 port map( A => n3515, B => n20366, S => n10960, Z => n3671);
   U8129 : INV_X1 port map( A => n12911, ZN => n13865);
   U8130 : OAI21_X1 port map( B1 => n4976, B2 => n4975, A => n4977, ZN => n3517
                           );
   U8131 : NAND3_X1 port map( A1 => n7751, A2 => n3520, A3 => n7752, ZN => 
                           n8658);
   U8132 : INV_X1 port map( A => n7752, ZN => n8999);
   U8134 : NAND2_X1 port map( A1 => n11070, A2 => n3521, ZN => n3638);
   U8135 : INV_X1 port map( A => n14465, ZN => n3522);
   U8136 : NOR2_X1 port map( A1 => n19531, A2 => n3522, ZN => n14364);
   U8137 : NAND2_X1 port map( A1 => n19657, A2 => n3522, ZN => n12726);
   U8138 : OAI22_X1 port map( A1 => n13924, A2 => n3522, B1 => n14363, B2 => 
                           n19538, ZN => n13925);
   U8139 : OAI211_X2 port map( C1 => n3526, C2 => n3525, A => n3524, B => n3523
                           , ZN => n9837);
   U8140 : INV_X1 port map( A => n8069, ZN => n3525);
   U8142 : NAND3_X1 port map( A1 => n5683, A2 => n5682, A3 => n3529, ZN => 
                           n3527);
   U8143 : NAND2_X1 port map( A1 => n5687, A2 => n5686, ZN => n3528);
   U8145 : NAND2_X1 port map( A1 => n11944, A2 => n11945, ZN => n3531);
   U8147 : NAND2_X1 port map( A1 => n3535, A2 => n17538, ZN => n18311);
   U8148 : INV_X1 port map( A => n12001, ZN => n11030);
   U8149 : NAND3_X1 port map( A1 => n14078, A2 => n14217, A3 => n877, ZN => 
                           n3539);
   U8150 : NAND2_X1 port map( A1 => n8235, A2 => n8083, ZN => n3540);
   U8151 : NAND2_X1 port map( A1 => n8234, A2 => n19826, ZN => n3541);
   U8152 : INV_X1 port map( A => n9204, ZN => n3542);
   U8153 : NAND2_X1 port map( A1 => n4233, A2 => n4907, ZN => n4378);
   U8154 : OR2_X1 port map( A1 => n18950, A2 => n18946, ZN => n3548);
   U8155 : INV_X1 port map( A => n18043, ZN => n18047);
   U8156 : NAND2_X1 port map( A1 => n18047, A2 => n3546, ZN => n3545);
   U8157 : NAND2_X1 port map( A1 => n3728, A2 => n20369, ZN => n3549);
   U8158 : XNOR2_X1 port map( A => n8339, B => n9994, ZN => n8396);
   U8159 : NOR2_X1 port map( A1 => n8999, A2 => n8997, ZN => n3557);
   U8162 : NAND2_X1 port map( A1 => n8773, A2 => n3557, ZN => n3556);
   U8163 : NAND3_X1 port map( A1 => n4865, A2 => n4652, A3 => n20356, ZN => 
                           n3561);
   U8165 : AOI21_X1 port map( B1 => n4867, B2 => n4870, A => n4865, ZN => n3564
                           );
   U8166 : OAI21_X1 port map( B1 => n4651, B2 => n3560, A => n3559, ZN => n4655
                           );
   U8167 : NAND2_X1 port map( A1 => n4381, A2 => n20357, ZN => n3559);
   U8168 : INV_X1 port map( A => n4867, ZN => n3560);
   U8169 : OAI21_X1 port map( B1 => n4651, B2 => n3562, A => n3561, ZN => n3563
                           );
   U8171 : NAND2_X1 port map( A1 => n12001, A2 => n12353, ZN => n12350);
   U8173 : NAND2_X1 port map( A1 => n164, A2 => n3978, ZN => n4659);
   U8174 : NAND2_X1 port map( A1 => n9660, A2 => n11383, ZN => n3566);
   U8175 : NAND3_X1 port map( A1 => n5447, A2 => n5825, A3 => n5826, ZN => 
                           n3567);
   U8176 : OAI21_X2 port map( B1 => n4231, B2 => n4230, A => n4229, ZN => n5823
                           );
   U8179 : XNOR2_X1 port map( A => n13864, B => n13184, ZN => n3575);
   U8181 : XNOR2_X1 port map( A => n3578, B => n18012, ZN => Ciphertext(34));
   U8182 : OAI211_X1 port map( C1 => n18010, C2 => n19526, A => n3580, B => 
                           n3579, ZN => n3578);
   U8183 : NAND2_X1 port map( A1 => n994, A2 => n18518, ZN => n3580);
   U8185 : INV_X1 port map( A => n7815, ZN => n3583);
   U8186 : NAND2_X1 port map( A1 => n3587, A2 => n19506, ZN => n3584);
   U8187 : NAND2_X1 port map( A1 => n3588, A2 => n11290, ZN => n11293);
   U8188 : XNOR2_X1 port map( A => n6927, B => n7143, ZN => n3590);
   U8189 : INV_X1 port map( A => n4483, ZN => n3592);
   U8190 : NAND2_X1 port map( A1 => n4968, A2 => n4482, ZN => n3593);
   U8191 : NAND2_X1 port map( A1 => n8265, A2 => n8264, ZN => n3594);
   U8192 : NAND3_X1 port map( A1 => n3596, A2 => n8266, A3 => n3597, ZN => 
                           n3595);
   U8193 : NAND2_X1 port map( A1 => n7864, A2 => n3766, ZN => n3596);
   U8194 : AOI21_X1 port map( B1 => n3598, B2 => n4449, A => n4077, ZN => n4078
                           );
   U8195 : INV_X1 port map( A => n14176, ZN => n3599);
   U8198 : NAND2_X1 port map( A1 => n20496, A2 => n3601, ZN => n11274);
   U8199 : NAND2_X1 port map( A1 => n5813, A2 => n19562, ZN => n3603);
   U8200 : NAND2_X1 port map( A1 => n5716, A2 => n3608, ZN => n5722);
   U8201 : NAND3_X2 port map( A1 => n7478, A2 => n3610, A3 => n3609, ZN => 
                           n8815);
   U8202 : NAND2_X1 port map( A1 => n7476, A2 => n20144, ZN => n3610);
   U8203 : NAND2_X1 port map( A1 => n3612, A2 => n11412, ZN => n3616);
   U8204 : NAND2_X1 port map( A1 => n3614, A2 => n3616, ZN => n12553);
   U8205 : NAND2_X1 port map( A1 => n11977, A2 => n12544, ZN => n11796);
   U8206 : INV_X1 port map( A => n8990, ZN => n9276);
   U8207 : OAI21_X1 port map( B1 => n8649, B2 => n9276, A => n9278, ZN => n3618
                           );
   U8208 : XNOR2_X1 port map( A => n10204, B => n10114, ZN => n9644);
   U8209 : INV_X1 port map( A => n7286, ZN => n6095);
   U8210 : XNOR2_X1 port map( A => n7286, B => n7285, ZN => n7293);
   U8211 : INV_X1 port map( A => n7026, ZN => n3619);
   U8212 : INV_X1 port map( A => n3620, ZN => n7380);
   U8213 : XNOR2_X1 port map( A => n6918, B => n6917, ZN => n3620);
   U8214 : AOI21_X1 port map( B1 => n15031, B2 => n15379, A => n3621, ZN => 
                           n15032);
   U8215 : MUX2_X1 port map( A => n19513, B => n15167, S => n15028, Z => n12936
                           );
   U8216 : NAND2_X1 port map( A1 => n14873, A2 => n3621, ZN => n14878);
   U8217 : OR2_X1 port map( A1 => n4532, A2 => n4528, ZN => n3623);
   U8218 : NAND2_X1 port map( A1 => n12125, A2 => n12230, ZN => n3626);
   U8219 : AND2_X1 port map( A1 => n5435, A2 => n6000, ZN => n3627);
   U8220 : NAND2_X1 port map( A1 => n5996, A2 => n6000, ZN => n5705);
   U8221 : XNOR2_X1 port map( A => n7122, B => n7081, ZN => n6621);
   U8222 : XNOR2_X1 port map( A => n6621, B => n6620, ZN => n6622);
   U8224 : NAND2_X1 port map( A1 => n10921, A2 => n10919, ZN => n10924);
   U8226 : NAND2_X1 port map( A1 => n12222, A2 => n12221, ZN => n10925);
   U8227 : XNOR2_X1 port map( A => n10348, B => n10085, ZN => n3628);
   U8228 : INV_X1 port map( A => n10348, ZN => n10086);
   U8229 : NAND2_X1 port map( A1 => n10104, A2 => n19949, ZN => n3630);
   U8230 : NOR2_X1 port map( A1 => n11658, A2 => n11955, ZN => n3632);
   U8231 : XOR2_X1 port map( A => n13530, B => n13579, Z => n12682);
   U8232 : NAND4_X2 port map( A1 => n12344, A2 => n12343, A3 => n12341, A4 => 
                           n12342, ZN => n13266);
   U8233 : OAI21_X2 port map( B1 => n4535, B2 => n4159, A => n3634, ZN => n5575
                           );
   U8234 : NAND3_X1 port map( A1 => n14357, A2 => n2039, A3 => n14422, ZN => 
                           n3635);
   U8235 : AND2_X2 port map( A1 => n12257, A2 => n3637, ZN => n12250);
   U8236 : NAND2_X1 port map( A1 => n11071, A2 => n11493, ZN => n3639);
   U8237 : INV_X1 port map( A => n5841, ZN => n3640);
   U8238 : NAND2_X1 port map( A1 => n4490, A2 => n210, ZN => n3641);
   U8239 : NAND2_X1 port map( A1 => n14263, A2 => n3642, ZN => n3643);
   U8240 : INV_X1 port map( A => n14262, ZN => n3642);
   U8241 : NAND2_X1 port map( A1 => n14019, A2 => n14262, ZN => n3644);
   U8242 : NAND2_X1 port map( A1 => n3643, A2 => n3644, ZN => n15759);
   U8243 : NAND2_X1 port map( A1 => n15756, A2 => n15754, ZN => n15587);
   U8244 : NAND2_X1 port map( A1 => n3645, A2 => n8917, ZN => n7668);
   U8245 : NAND2_X1 port map( A1 => n4835, A2 => n3846, ZN => n4417);
   U8246 : OAI21_X1 port map( B1 => n20256, B2 => n4676, A => n4417, ZN => 
                           n3652);
   U8247 : NAND2_X1 port map( A1 => n2042, A2 => n19508, ZN => n4418);
   U8248 : NAND2_X1 port map( A1 => n8080, A2 => n20174, ZN => n3653);
   U8249 : NAND2_X1 port map( A1 => n8077, A2 => n3655, ZN => n3654);
   U8250 : NAND2_X1 port map( A1 => n4960, A2 => n292, ZN => n3656);
   U8251 : NAND2_X1 port map( A1 => n3656, A2 => n20205, ZN => n4138);
   U8252 : OAI211_X1 port map( C1 => n3657, C2 => n4899, A => n4898, B => n4892
                           , ZN => n4900);
   U8253 : AND2_X1 port map( A1 => n3658, A2 => n4375, ZN => n3745);
   U8254 : NOR2_X2 port map( A1 => n8422, A2 => n8421, ZN => n9111);
   U8255 : NAND2_X1 port map( A1 => n3659, A2 => n3661, ZN => n8422);
   U8256 : NAND2_X1 port map( A1 => n8285, A2 => n8284, ZN => n3661);
   U8257 : INV_X1 port map( A => n5984, ZN => n3663);
   U8258 : NOR2_X1 port map( A1 => n3665, A2 => n5558, ZN => n5560);
   U8259 : NAND2_X1 port map( A1 => n3665, A2 => n6051, ZN => n5141);
   U8260 : NAND2_X1 port map( A1 => n13164, A2 => n14535, ZN => n13165);
   U8261 : NAND2_X1 port map( A1 => n12311, A2 => n12312, ZN => n3666);
   U8263 : OAI21_X1 port map( B1 => n11340, B2 => n9830, A => n3669, ZN => 
                           n9831);
   U8264 : INV_X1 port map( A => n10673, ZN => n3669);
   U8266 : INV_X1 port map( A => n13618, ZN => n3675);
   U8267 : XNOR2_X1 port map( A => n13085, B => n3675, ZN => n13415);
   U8268 : NAND3_X1 port map( A1 => n10990, A2 => n11869, A3 => n11302, ZN => 
                           n10715);
   U8269 : NAND2_X1 port map( A1 => n3681, A2 => n3678, ZN => n3677);
   U8270 : NAND2_X1 port map( A1 => n3679, A2 => n208, ZN => n3678);
   U8271 : NAND2_X1 port map( A1 => n20490, A2 => n20270, ZN => n3680);
   U8274 : OAI21_X1 port map( B1 => n3689, B2 => n3690, A => n15769, ZN => 
                           n3687);
   U8275 : AND2_X2 port map( A1 => n3687, A2 => n3686, ZN => n16742);
   U8276 : AOI21_X1 port map( B1 => n15766, B2 => n15767, A => n229, ZN => 
                           n3688);
   U8277 : OAI22_X1 port map( A1 => n14273, A2 => n14566, B1 => n14275, B2 => 
                           n14563, ZN => n3694);
   U8278 : AND2_X2 port map( A1 => n3698, A2 => n3695, ZN => n15866);
   U8279 : NAND2_X1 port map( A1 => n3699, A2 => n20518, ZN => n3698);
   U8280 : NAND2_X1 port map( A1 => n13903, A2 => n13902, ZN => n3699);
   U8283 : NAND2_X1 port map( A1 => n14703, A2 => n3705, ZN => n3704);
   U8284 : OAI21_X1 port map( B1 => n6090, B2 => n6089, A => n890, ZN => n6093)
                           ;
   U8285 : NAND2_X1 port map( A1 => n5905, A2 => n4862, ZN => n6089);
   U8286 : NAND2_X1 port map( A1 => n4859, A2 => n3706, ZN => n5905);
   U8287 : NAND2_X1 port map( A1 => n11707, A2 => n12480, ZN => n3707);
   U8288 : XNOR2_X1 port map( A => n12849, B => n13048, ZN => n12998);
   U8289 : NAND2_X1 port map( A1 => n15081, A2 => n15531, ZN => n15916);
   U8290 : NAND2_X1 port map( A1 => n15919, A2 => n15081, ZN => n3709);
   U8292 : NAND2_X1 port map( A1 => n11219, A2 => n204, ZN => n3713);
   U8293 : NAND2_X1 port map( A1 => n4612, A2 => n3716, ZN => n3715);
   U8294 : NAND2_X1 port map( A1 => n20509, A2 => n5742, ZN => n5202);
   U8295 : NAND2_X1 port map( A1 => n5271, A2 => n19865, ZN => n3719);
   U8296 : NAND2_X1 port map( A1 => n11620, A2 => n1371, ZN => n3721);
   U8297 : INV_X1 port map( A => n5743, ZN => n5746);
   U8298 : NAND2_X1 port map( A1 => n15642, A2 => n15256, ZN => n15835);
   U8299 : NAND2_X1 port map( A1 => n15642, A2 => n3722, ZN => n3723);
   U8300 : NAND2_X1 port map( A1 => n3724, A2 => n3723, ZN => n15099);
   U8301 : NAND2_X1 port map( A1 => n15095, A2 => n3725, ZN => n3724);
   U8302 : INV_X1 port map( A => n19931, ZN => n3725);
   U8303 : OR2_X1 port map( A1 => n14664, A2 => n14662, ZN => n14536);
   U8304 : INV_X1 port map( A => n14662, ZN => n3726);
   U8305 : NOR2_X1 port map( A1 => n3726, A2 => n13164, ZN => n14668);
   U8306 : AND3_X1 port map( A1 => n3727, A2 => n14662, A3 => n14664, ZN => 
                           n13178);
   U8307 : NAND2_X1 port map( A1 => n14666, A2 => n14667, ZN => n3727);
   U8308 : NAND2_X1 port map( A1 => n20369, A2 => n4633, ZN => n4637);
   U8309 : INV_X1 port map( A => n18842, ZN => n18813);
   U8310 : NAND2_X1 port map( A1 => n18275, A2 => n221, ZN => n3729);
   U8311 : OR2_X1 port map( A1 => n18275, A2 => n17769, ZN => n3730);
   U8312 : NAND2_X1 port map( A1 => n11888, A2 => n3732, ZN => n3731);
   U8313 : INV_X1 port map( A => n12264, ZN => n3733);
   U8314 : OAI21_X1 port map( B1 => n12261, B2 => n3734, A => n12016, ZN => 
                           n11894);
   U8315 : NOR2_X1 port map( A1 => n11727, A2 => n3734, ZN => n11728);
   U8316 : XNOR2_X1 port map( A => n14914, B => n3735, ZN => n14915);
   U8317 : NAND2_X1 port map( A1 => n3739, A2 => n3737, ZN => n3736);
   U8318 : NAND2_X1 port map( A1 => n3738, A2 => n14900, ZN => n3737);
   U8319 : NOR2_X1 port map( A1 => n3741, A2 => n14901, ZN => n3738);
   U8320 : OAI21_X1 port map( B1 => n3740, B2 => n3741, A => n14901, ZN => 
                           n3739);
   U8321 : INV_X1 port map( A => n14900, ZN => n3740);
   U8322 : OAI21_X1 port map( B1 => n15916, B2 => n15420, A => n14899, ZN => 
                           n3741);
   U8323 : INV_X1 port map( A => n14120, ZN => n14230);
   U8324 : XNOR2_X1 port map( A => n13705, B => n2257, ZN => n3744);
   U8325 : NAND2_X1 port map( A1 => n5484, A2 => n3746, ZN => n7163);
   U8327 : NAND2_X1 port map( A1 => n3748, A2 => n8301, ZN => n7876);
   U8328 : NAND2_X1 port map( A1 => n3747, A2 => n20057, ZN => n5299);
   U8329 : AND2_X1 port map( A1 => n19865, A2 => n8044, ZN => n3747);
   U8330 : NAND3_X1 port map( A1 => n8308, A2 => n8306, A3 => n8307, ZN => 
                           n3750);
   U8332 : NAND2_X1 port map( A1 => n4338, A2 => n3753, ZN => n3752);
   U8333 : NAND2_X1 port map( A1 => n11628, A2 => n11627, ZN => n11969);
   U8334 : INV_X1 port map( A => n17836, ZN => n3755);
   U8335 : INV_X1 port map( A => n16731, ZN => n17838);
   U8336 : OAI21_X1 port map( B1 => n16731, B2 => n3755, A => n17840, ZN => 
                           n16733);
   U8338 : NAND2_X1 port map( A1 => n3951, A2 => n3759, ZN => n5148);
   U8340 : NAND2_X1 port map( A1 => n8264, A2 => n7864, ZN => n3765);
   U8341 : NAND2_X1 port map( A1 => n7569, A2 => n3766, ZN => n7574);
   U8342 : MUX2_X1 port map( A => n6698, B => n6699, S => n8262, Z => n6700);
   U8343 : AOI21_X2 port map( B1 => n5585, B2 => n5586, A => n5584, ZN => n5884
                           );
   U8345 : MUX2_X1 port map( A => n6071, B => n6072, S => n6068, Z => n6073);
   U8346 : OAI21_X1 port map( B1 => n3768, B2 => n9913, A => n9921, ZN => n9930
                           );
   U8347 : MUX2_X1 port map( A => n4902, B => n4497, S => n4856, Z => n3991);
   U8348 : AND2_X1 port map( A1 => n4904, A2 => n4856, ZN => n5901);
   U8349 : AND2_X1 port map( A1 => n4497, A2 => n4498, ZN => n3770);
   U8350 : NAND2_X1 port map( A1 => n4856, A2 => n4907, ZN => n4498);
   U8351 : NAND2_X1 port map( A1 => n3774, A2 => n3772, ZN => n3771);
   U8352 : NAND2_X1 port map( A1 => n20493, A2 => n8099, ZN => n3774);
   U8353 : OR2_X1 port map( A1 => n3776, A2 => n19171, ZN => n16115);
   U8354 : INV_X1 port map( A => n19171, ZN => n18088);
   U8355 : INV_X1 port map( A => n16115, ZN => n16154);
   U8356 : NAND2_X1 port map( A1 => n1003, A2 => n12497, ZN => n3777);
   U8357 : XNOR2_X1 port map( A => n3779, B => n14164, ZN => n16171);
   U8358 : XNOR2_X1 port map( A => n16185, B => n16396, ZN => n3779);
   U8359 : OR2_X1 port map( A1 => n12382, A2 => n12386, ZN => n3782);
   U8360 : NOR2_X1 port map( A1 => n3782, A2 => n11915, ZN => n3781);
   U8363 : NAND2_X1 port map( A1 => n7935, A2 => n7932, ZN => n3784);
   U8364 : NAND2_X1 port map( A1 => n6244, A2 => n20359, ZN => n3785);
   U8365 : NAND2_X1 port map( A1 => n19936, A2 => n19362, ZN => n17860);
   U8367 : MUX2_X1 port map( A => n17863, B => n20212, S => n17672, Z => n17673
                           );
   U8369 : XNOR2_X1 port map( A => n10514, B => n10052, ZN => n3787);
   U8370 : AND2_X1 port map( A1 => n3789, A2 => n11177, ZN => n9378);
   U8371 : INV_X1 port map( A => n10962, ZN => n3789);
   U8374 : INV_X1 port map( A => n7645, ZN => n3795);
   U8375 : INV_X1 port map( A => n4343, ZN => n3925);
   U8378 : OR2_X1 port map( A1 => n12600, A2 => n12601, ZN => n11627);
   U8380 : BUF_X1 port map( A => n19098, Z => n19094);
   U8381 : AND2_X1 port map( A1 => n18834, A2 => n18829, ZN => n18833);
   U8383 : OR2_X1 port map( A1 => n18061, A2 => n19040, ZN => n18081);
   U8384 : XNOR2_X1 port map( A => n16411, B => n16410, ZN => n18097);
   U8386 : OR2_X1 port map( A1 => n15785, A2 => n15783, ZN => n15691);
   U8387 : XNOR2_X1 port map( A => n10180, B => n10030, ZN => n10290);
   U8388 : OR2_X1 port map( A1 => n12209, A2 => n12208, ZN => n12187);
   U8389 : BUF_X1 port map( A => n19441, Z => n19448);
   U8390 : INV_X1 port map( A => n18140, ZN => n17384);
   U8392 : OR2_X1 port map( A1 => n18568, A2 => n18199, ZN => n18561);
   U8393 : OR2_X1 port map( A1 => n18532, A2 => n18529, ZN => n16816);
   U8394 : INV_X1 port map( A => n17705, ZN => n17706);
   U8395 : XNOR2_X1 port map( A => n16082, B => n2392, ZN => n15798);
   U8396 : XNOR2_X1 port map( A => n6829, B => n6828, ZN => n6837);
   U8397 : AND2_X1 port map( A1 => n5967, A2 => n5699, ZN => n5449);
   U8398 : OAI21_X1 port map( B1 => n854, B2 => n17186, A => n17185, ZN => 
                           n19092);
   U8399 : XNOR2_X1 port map( A => n16121, B => n16120, ZN => n17835);
   U8401 : AND2_X1 port map( A1 => n14327, A2 => n14818, ZN => n14086);
   U8403 : XNOR2_X1 port map( A => n13521, B => n13520, ZN => n13522);
   U8406 : OR2_X1 port map( A1 => n15153, A2 => n192, ZN => n15704);
   U8407 : AND2_X1 port map( A1 => n15380, A2 => n15379, ZN => n15382);
   U8408 : INV_X1 port map( A => n6010, ZN => n5590);
   U8409 : NOR2_X2 port map( A1 => n15186, A2 => n15185, ZN => n16608);
   U8410 : AND2_X1 port map( A1 => n14811, A2 => n14810, ZN => n14814);
   U8412 : NAND2_X1 port map( A1 => n12767, A2 => n12766, ZN => n12842);
   U8413 : OR2_X1 port map( A1 => n18495, A2 => n18498, ZN => n17644);
   U8414 : OAI22_X1 port map( A1 => n17617, A2 => n17616, B1 => n17615, B2 => 
                           n1773, ZN => n17621);
   U8415 : OR2_X1 port map( A1 => n19396, A2 => n17656, ZN => n16683);
   U8416 : OR2_X1 port map( A1 => n10663, A2 => n11321, ZN => n10666);
   U8417 : XNOR2_X1 port map( A => n8567, B => n8566, ZN => n10761);
   U8419 : NOR2_X1 port map( A1 => n18358, A2 => n18290, ZN => n18288);
   U8420 : AND2_X1 port map( A1 => n18489, A2 => n18500, ZN => n17735);
   U8421 : AND2_X1 port map( A1 => n18322, A2 => n18321, ZN => n18326);
   U8423 : OR2_X1 port map( A1 => n18700, A2 => n18699, ZN => n18705);
   U8424 : NOR2_X1 port map( A1 => n16493, A2 => n16492, ZN => n16494);
   U8425 : AND3_X1 port map( A1 => n17234, A2 => n17235, A3 => n17233, ZN => 
                           n18382);
   U8426 : AND2_X1 port map( A1 => n16544, A2 => n19955, ZN => n19315);
   U8427 : XNOR2_X1 port map( A => n17044, B => n17043, ZN => n17187);
   U8428 : AND2_X1 port map( A1 => n18362, A2 => n18365, ZN => n17937);
   U8431 : NOR3_X1 port map( A1 => n228, A2 => n19958, A3 => n15581, ZN => 
                           n14834);
   U8433 : OR2_X1 port map( A1 => n17896, A2 => n19707, ZN => n16782);
   U8435 : XNOR2_X1 port map( A => n13235, B => n13236, ZN => n14269);
   U8436 : XNOR2_X1 port map( A => n10244, B => n10243, ZN => n11120);
   U8437 : OR2_X1 port map( A1 => n4827, A2 => n5258, ZN => n4671);
   U8438 : OR2_X1 port map( A1 => n19227, A2 => n19754, ZN => n19219);
   U8439 : OR2_X1 port map( A1 => n11120, A2 => n11880, ZN => n10810);
   U8442 : INV_X1 port map( A => n15295, ZN => n14944);
   U8443 : AND2_X1 port map( A1 => n11871, A2 => n11390, ZN => n11303);
   U8445 : OAI211_X2 port map( C1 => n10193, C2 => n11427, A => n10192, B => 
                           n10191, ZN => n11990);
   U8447 : AOI21_X2 port map( B1 => n9003, B2 => n7776, A => n7775, ZN => n9667
                           );
   U8448 : NOR2_X1 port map( A1 => n12648, A2 => n12686, ZN => n12093);
   U8451 : AOI22_X1 port map( A1 => n16497, A2 => n19403, B1 => n19402, B2 => 
                           n16307, ZN => n19182);
   U8452 : AND2_X1 port map( A1 => n19952, A2 => n12311, ZN => n11905);
   U8453 : AND2_X1 port map( A1 => n4632, A2 => n5743, ZN => n3796);
   U8454 : AND3_X1 port map( A1 => n12362, A2 => n12363, A3 => n12510, ZN => 
                           n3798);
   U8455 : OR2_X1 port map( A1 => n8934, A2 => n8933, ZN => n3799);
   U8456 : AND2_X1 port map( A1 => n9330, A2 => n9328, ZN => n3800);
   U8457 : AND3_X1 port map( A1 => n20215, A2 => n12281, A3 => n12042, ZN => 
                           n3801);
   U8458 : AND2_X1 port map( A1 => n5219, A2 => n5217, ZN => n3802);
   U8459 : XNOR2_X1 port map( A => n3803, B => n7351, ZN => n7470);
   U8460 : XOR2_X1 port map( A => n7350, B => n7349, Z => n3803);
   U8461 : AND2_X1 port map( A1 => n6059, A2 => n906, ZN => n3804);
   U8462 : XOR2_X1 port map( A => n6737, B => n6209, Z => n3805);
   U8463 : OR2_X1 port map( A1 => n7510, A2 => n7675, ZN => n3808);
   U8464 : OR2_X1 port map( A1 => n8325, A2 => n7585, ZN => n3809);
   U8465 : XOR2_X1 port map( A => n9989, B => n9988, Z => n3810);
   U8466 : XOR2_X1 port map( A => n10616, B => n10615, Z => n3812);
   U8467 : OR2_X1 port map( A1 => n12334, A2 => n12332, ZN => n3813);
   U8468 : AND2_X1 port map( A1 => n11495, A2 => n11493, ZN => n3814);
   U8470 : OR2_X1 port map( A1 => n15430, A2 => n15531, ZN => n3817);
   U8471 : OR2_X1 port map( A1 => n20263, A2 => n14482, ZN => n3818);
   U8472 : AND2_X1 port map( A1 => n15496, A2 => n15500, ZN => n3819);
   U8473 : AND3_X1 port map( A1 => n14637, A2 => n20473, A3 => n14512, ZN => 
                           n3820);
   U8474 : AND2_X1 port map( A1 => n19502, A2 => n15516, ZN => n3821);
   U8475 : INV_X1 port map( A => n14316, ZN => n13164);
   U8476 : XOR2_X1 port map( A => n13573, B => n13574, Z => n3823);
   U8477 : AND2_X1 port map( A1 => n15413, A2 => n15553, ZN => n3824);
   U8478 : XNOR2_X1 port map( A => n16074, B => n16073, ZN => n17878);
   U8479 : INV_X1 port map( A => n18519, ZN => n18184);
   U8480 : OR2_X1 port map( A1 => n16101, A2 => n17891, ZN => n3825);
   U8481 : BUF_X1 port map( A => n16155, Z => n18319);
   U8482 : OR2_X1 port map( A1 => n17715, A2 => n17835, ZN => n3826);
   U8483 : OR2_X1 port map( A1 => n19381, A2 => n19439, ZN => n3827);
   U8484 : AND2_X1 port map( A1 => n19441, A2 => n19444, ZN => n3828);
   U8485 : BUF_X1 port map( A => n19182, Z => n19189);
   U8486 : NAND3_X1 port map( A1 => n18666, A2 => n17964, A3 => n19735, ZN => 
                           n3829);
   U8487 : OR2_X1 port map( A1 => n5107, A2 => n5101, ZN => n4450);
   U8489 : OR2_X1 port map( A1 => n5095, A2 => n4405, ZN => n3859);
   U8490 : INV_X1 port map( A => n4319, ZN => n4127);
   U8491 : OR2_X1 port map( A1 => n4518, A2 => n4343, ZN => n4344);
   U8492 : INV_X1 port map( A => Plaintext(23), ZN => n3874);
   U8493 : OR2_X1 port map( A1 => n4011, A2 => n4611, ZN => n4612);
   U8494 : XNOR2_X1 port map( A => Key(159), B => Plaintext(159), ZN => n4575);
   U8496 : OR2_X1 port map( A1 => n4669, A2 => n4214, ZN => n4425);
   U8497 : OR2_X1 port map( A1 => n4627, A2 => n4626, ZN => n4628);
   U8498 : OAI21_X1 port map( B1 => n4125, B2 => n4127, A => n4126, ZN => n4130
                           );
   U8500 : NAND2_X1 port map( A1 => n4838, A2 => n4837, ZN => n5492);
   U8501 : INV_X1 port map( A => n5766, ZN => n5545);
   U8502 : OR2_X1 port map( A1 => n5088, A2 => n19776, ZN => n4438);
   U8504 : OR2_X1 port map( A1 => n4954, A2 => n4953, ZN => n4477);
   U8505 : INV_X1 port map( A => n5559, ZN => n3929);
   U8506 : OR2_X1 port map( A1 => n5997, A2 => n5998, ZN => n5813);
   U8507 : INV_X1 port map( A => n6129, ZN => n5356);
   U8508 : OR2_X1 port map( A1 => n5802, A2 => n5382, ZN => n6190);
   U8509 : INV_X1 port map( A => n6379, ZN => n5730);
   U8510 : AND2_X1 port map( A1 => n6052, A2 => n6048, ZN => n5558);
   U8511 : INV_X1 port map( A => n5393, ZN => n5368);
   U8513 : INV_X1 port map( A => n5502, ZN => n5122);
   U8516 : OR2_X1 port map( A1 => n5317, A2 => n5581, ZN => n5150);
   U8517 : INV_X1 port map( A => n5899, ZN => n5908);
   U8518 : NOR2_X1 port map( A1 => n284, A2 => n5953, ZN => n5950);
   U8519 : OAI211_X1 port map( C1 => n5593, C2 => n5594, A => n5592, B => n5591
                           , ZN => n7115);
   U8520 : OR2_X1 port map( A1 => n5855, A2 => n5612, ZN => n5353);
   U8521 : OR2_X1 port map( A1 => n5363, A2 => n4598, ZN => n5215);
   U8522 : OR2_X1 port map( A1 => n7948, A2 => n7953, ZN => n7168);
   U8523 : XNOR2_X1 port map( A => n6605, B => n6604, ZN => n7632);
   U8525 : OR2_X1 port map( A1 => n20360, A2 => n7936, ZN => n7761);
   U8526 : XNOR2_X1 port map( A => n6671, B => n6670, ZN => n7568);
   U8527 : BUF_X1 port map( A => n7632, Z => n7633);
   U8528 : INV_X1 port map( A => n8029, ZN => n7469);
   U8529 : INV_X1 port map( A => n8011, ZN => n8012);
   U8531 : INV_X1 port map( A => n7407, ZN => n7077);
   U8532 : XNOR2_X1 port map( A => n5238, B => n5239, ZN => n7877);
   U8533 : OR2_X1 port map( A1 => n20180, A2 => n7644, ZN => n6468);
   U8535 : INV_X1 port map( A => n8055, ZN => n8052);
   U8536 : OR2_X1 port map( A1 => n7003, A2 => n7903, ZN => n6284);
   U8537 : XNOR2_X1 port map( A => n6493, B => n6492, ZN => n6702);
   U8538 : INV_X1 port map( A => n6837, ZN => n7724);
   U8539 : INV_X1 port map( A => n8131, ZN => n8138);
   U8540 : XNOR2_X1 port map( A => n6781, B => n6780, ZN => n7684);
   U8541 : OR2_X1 port map( A1 => n7958, A2 => n7956, ZN => n7917);
   U8542 : AND2_X1 port map( A1 => n7749, A2 => n7508, ZN => n6908);
   U8543 : OR2_X1 port map( A1 => n7676, A2 => n7673, ZN => n7513);
   U8544 : AOI22_X1 port map( A1 => n20012, A2 => n7445, B1 => n8280, B2 => 
                           n8286, ZN => n7796);
   U8545 : AOI22_X1 port map( A1 => n8154, A2 => n8153, B1 => n8262, B2 => 
                           n8152, ZN => n8156);
   U8546 : AND2_X1 port map( A1 => n8185, A2 => n8184, ZN => n8187);
   U8547 : INV_X1 port map( A => n9346, ZN => n9567);
   U8548 : INV_X1 port map( A => n8482, ZN => n9368);
   U8549 : NOR2_X1 port map( A1 => n8423, A2 => n19515, ZN => n8327);
   U8550 : INV_X1 port map( A => n9934, ZN => n10037);
   U8551 : INV_X1 port map( A => n11339, ZN => n11340);
   U8552 : XNOR2_X1 port map( A => n9878, B => n9635, ZN => n10462);
   U8553 : INV_X1 port map( A => n11489, ZN => n11494);
   U8554 : INV_X1 port map( A => n9294, ZN => n8680);
   U8555 : XNOR2_X1 port map( A => n9653, B => n9652, ZN => n10684);
   U8556 : AOI21_X1 port map( B1 => n11564, B2 => n11567, A => n11469, ZN => 
                           n11470);
   U8557 : XNOR2_X1 port map( A => n10433, B => n9387, ZN => n9390);
   U8558 : NOR2_X1 port map( A1 => n11253, A2 => n11255, ZN => n11323);
   U8559 : XNOR2_X1 port map( A => n10075, B => n10076, ZN => n10112);
   U8560 : OR2_X1 port map( A1 => n19750, A2 => n11866, ZN => n11304);
   U8561 : OR2_X1 port map( A1 => n11452, A2 => n11110, ZN => n10734);
   U8563 : XNOR2_X1 port map( A => n9990, B => n3810, ZN => n10742);
   U8564 : BUF_X1 port map( A => n10783, Z => n11116);
   U8565 : NOR2_X1 port map( A1 => n19959, A2 => n11133, ZN => n11421);
   U8566 : INV_X1 port map( A => n11445, ZN => n11209);
   U8567 : NOR2_X1 port map( A1 => n11513, A2 => n19864, ZN => n11574);
   U8568 : AND2_X1 port map( A1 => n10704, A2 => n11152, ZN => n10707);
   U8569 : BUF_X1 port map( A => n9666, Z => n11383);
   U8570 : OR2_X1 port map( A1 => n12616, A2 => n12053, ZN => n12055);
   U8571 : NOR2_X1 port map( A1 => n12545, A2 => n12544, ZN => n12555);
   U8572 : INV_X1 port map( A => n12809, ZN => n12487);
   U8573 : OR2_X1 port map( A1 => n12508, A2 => n12359, ZN => n9886);
   U8574 : AND2_X1 port map( A1 => n11686, A2 => n11863, ZN => n11730);
   U8575 : INV_X1 port map( A => n11841, ZN => n12181);
   U8576 : XNOR2_X1 port map( A => n13481, B => n457, ZN => n13432);
   U8577 : OAI21_X1 port map( B1 => n11908, B2 => n11907, A => n11906, ZN => 
                           n13451);
   U8578 : AND2_X1 port map( A1 => n12383, A2 => n12382, ZN => n12388);
   U8579 : OR2_X1 port map( A1 => n12595, A2 => n12201, ZN => n12060);
   U8580 : OR2_X1 port map( A1 => n12333, A2 => n12332, ZN => n12344);
   U8581 : AND2_X1 port map( A1 => n11971, A2 => n11970, ZN => n11972);
   U8582 : INV_X1 port map( A => n13481, ZN => n12984);
   U8584 : OAI21_X1 port map( B1 => n11974, B2 => n11667, A => n11666, ZN => 
                           n11668);
   U8585 : XNOR2_X1 port map( A => n13432, B => n13797, ZN => n13434);
   U8586 : XNOR2_X1 port map( A => n12962, B => n2347, ZN => n12964);
   U8587 : XNOR2_X1 port map( A => n13714, B => n13499, ZN => n11789);
   U8588 : XNOR2_X1 port map( A => n13477, B => n13279, ZN => n13316);
   U8589 : OR2_X1 port map( A1 => n14279, A2 => n14555, ZN => n14280);
   U8591 : OR2_X1 port map( A1 => n14132, A2 => n14729, ZN => n14133);
   U8592 : XNOR2_X1 port map( A => n12970, B => n13207, ZN => n12972);
   U8594 : XNOR2_X1 port map( A => n13015, B => n13014, ZN => n13872);
   U8595 : BUF_X1 port map( A => n13980, Z => n14542);
   U8596 : INV_X1 port map( A => n14543, ZN => n14544);
   U8598 : OR2_X1 port map( A1 => n14304, A2 => n14506, ZN => n13506);
   U8599 : XNOR2_X1 port map( A => n13639, B => n13638, ZN => n14388);
   U8600 : INV_X1 port map( A => n14104, ZN => n14105);
   U8601 : AND2_X1 port map( A1 => n3307, A2 => n15296, ZN => n14768);
   U8602 : OR2_X1 port map( A1 => n15696, A2 => n15695, ZN => n14938);
   U8603 : AND2_X1 port map( A1 => n13907, A2 => n14611, ZN => n14207);
   U8604 : AND2_X1 port map( A1 => n19485, A2 => n12877, ZN => n12878);
   U8605 : INV_X1 port map( A => n14699, ZN => n14122);
   U8606 : AND2_X1 port map( A1 => n14089, A2 => n14088, ZN => n14090);
   U8607 : BUF_X1 port map( A => n12910, Z => n14168);
   U8608 : XNOR2_X1 port map( A => n13472, B => n13473, ZN => n14425);
   U8609 : AND2_X1 port map( A1 => n14508, A2 => n14507, ZN => n14513);
   U8610 : INV_X1 port map( A => n15600, ZN => n15271);
   U8611 : AND2_X1 port map( A1 => n14434, A2 => n14487, ZN => n13881);
   U8612 : NOR2_X1 port map( A1 => n15606, A2 => n16128, ZN => n15201);
   U8613 : INV_X1 port map( A => n13982, ZN => n13133);
   U8614 : BUF_X1 port map( A => n14497, Z => n14501);
   U8615 : OR2_X1 port map( A1 => n15595, A2 => n15748, ZN => n15519);
   U8616 : AND2_X1 port map( A1 => n15636, A2 => n15843, ZN => n15092);
   U8617 : OR2_X1 port map( A1 => n15704, A2 => n13968, ZN => n13969);
   U8618 : OR2_X1 port map( A1 => n15909, A2 => n15907, ZN => n15416);
   U8619 : INV_X1 port map( A => n14964, ZN => n14969);
   U8620 : BUF_X1 port map( A => n15655, Z => n15768);
   U8621 : INV_X1 port map( A => n15532, ZN => n15086);
   U8622 : NAND4_X1 port map( A1 => n15649, A2 => n15648, A3 => n15647, A4 => 
                           n15646, ZN => n15994);
   U8623 : NOR2_X1 port map( A1 => n14876, A2 => n14875, ZN => n14877);
   U8624 : OR2_X1 port map( A1 => n13861, A2 => n13860, ZN => n13862);
   U8625 : OAI21_X1 port map( B1 => n14959, B2 => n15284, A => n14958, ZN => 
                           n15020);
   U8626 : OAI21_X1 port map( B1 => n15290, B2 => n15289, A => n15288, ZN => 
                           n16992);
   U8627 : OR2_X1 port map( A1 => n2005, A2 => n15445, ZN => n15324);
   U8628 : OR2_X1 port map( A1 => n15540, A2 => n15898, ZN => n15541);
   U8629 : XNOR2_X1 port map( A => n16419, B => n16418, ZN => n16422);
   U8630 : INV_X1 port map( A => n18946, ZN => n17687);
   U8631 : XNOR2_X1 port map( A => n16593, B => n16706, ZN => n17357);
   U8632 : BUF_X1 port map( A => n19782, Z => n16420);
   U8633 : XNOR2_X1 port map( A => n15798, B => n17426, ZN => n15810);
   U8634 : AND2_X1 port map( A1 => n17492, A2 => n17491, ZN => n17496);
   U8635 : AND2_X1 port map( A1 => n19943, A2 => n20348, ZN => n17966);
   U8636 : XNOR2_X1 port map( A => n16428, B => n16427, ZN => n17568);
   U8638 : INV_X1 port map( A => n17568, ZN => n18095);
   U8639 : XNOR2_X1 port map( A => n17364, B => n17363, ZN => n17758);
   U8640 : OAI21_X1 port map( B1 => n18115, B2 => n19885, A => n17968, ZN => 
                           n17460);
   U8641 : AND2_X1 port map( A1 => n18033, A2 => n18270, ZN => n17768);
   U8642 : OR2_X1 port map( A1 => n18019, A2 => n18938, ZN => n17705);
   U8643 : XNOR2_X1 port map( A => n16133, B => n16132, ZN => n17063);
   U8644 : INV_X1 port map( A => n17892, ZN => n16784);
   U8645 : OR2_X1 port map( A1 => n17676, A2 => n17078, ZN => n16314);
   U8646 : XNOR2_X1 port map( A => n15790, B => n15789, ZN => n16540);
   U8649 : BUF_X1 port map( A => n17501, Z => n17504);
   U8650 : AOI21_X1 port map( B1 => n17159, B2 => n17158, A => n17157, ZN => 
                           n17623);
   U8651 : AND2_X1 port map( A1 => n20109, A2 => n18097, ZN => n17164);
   U8655 : NOR2_X1 port map( A1 => n20273, A2 => n16673, ZN => n16636);
   U8656 : INV_X1 port map( A => n19432, ZN => n19418);
   U8657 : OR2_X1 port map( A1 => n18240, A2 => n20128, ZN => n18247);
   U8658 : AND2_X1 port map( A1 => n20003, A2 => n18412, ZN => n18406);
   U8659 : BUF_X1 port map( A => n17729, Z => n17640);
   U8660 : OR2_X1 port map( A1 => n17476, A2 => n17475, ZN => n17477);
   U8663 : OR2_X1 port map( A1 => n17719, A2 => n17718, ZN => n17720);
   U8665 : OR2_X1 port map( A1 => n18320, A2 => n16155, ZN => n18321);
   U8666 : BUF_X1 port map( A => n18621, Z => n18613);
   U8667 : OR2_X1 port map( A1 => n19425, A2 => n19409, ZN => n19428);
   U8668 : AND3_X1 port map( A1 => n17789, A2 => n19166, A3 => n17791, ZN => 
                           n17796);
   U8669 : INV_X1 port map( A => Plaintext(71), ZN => n3830);
   U8670 : XNOR2_X1 port map( A => n3830, B => Key(71), ZN => n4220);
   U8671 : NAND2_X1 port map( A1 => n4223, A2 => n164, ZN => n3832);
   U8672 : INV_X1 port map( A => Plaintext(70), ZN => n3831);
   U8673 : XNOR2_X1 port map( A => Key(66), B => Plaintext(66), ZN => n4657);
   U8674 : AOI21_X1 port map( B1 => n3979, B2 => n4657, A => n164, ZN => n3833)
                           ;
   U8675 : INV_X1 port map( A => n3855, ZN => n3839);
   U8677 : INV_X1 port map( A => Plaintext(85), ZN => n3834);
   U8678 : XNOR2_X1 port map( A => n3834, B => Key(85), ZN => n4663);
   U8679 : INV_X1 port map( A => Plaintext(84), ZN => n3835);
   U8680 : XNOR2_X1 port map( A => n3835, B => Key(84), ZN => n4664);
   U8681 : INV_X1 port map( A => n4664, ZN => n4816);
   U8682 : INV_X1 port map( A => Plaintext(89), ZN => n3836);
   U8683 : INV_X1 port map( A => n4410, ZN => n4411);
   U8684 : XNOR2_X1 port map( A => Key(88), B => Plaintext(88), ZN => n5071);
   U8685 : NAND2_X1 port map( A1 => n4411, A2 => n5071, ZN => n4814);
   U8686 : INV_X1 port map( A => Plaintext(80), ZN => n3840);
   U8687 : XNOR2_X1 port map( A => n3840, B => Key(80), ZN => n3843);
   U8688 : INV_X1 port map( A => n3843, ZN => n4835);
   U8689 : INV_X1 port map( A => Plaintext(83), ZN => n3841);
   U8690 : XNOR2_X1 port map( A => n3841, B => Key(83), ZN => n3846);
   U8691 : INV_X1 port map( A => n3846, ZN => n4675);
   U8692 : INV_X1 port map( A => n5117, ZN => n4834);
   U8693 : NAND2_X1 port map( A1 => n3842, A2 => n4834, ZN => n3850);
   U8694 : INV_X1 port map( A => Plaintext(82), ZN => n3844);
   U8695 : XNOR2_X1 port map( A => Key(78), B => Plaintext(78), ZN => n5118);
   U8696 : INV_X1 port map( A => n5118, ZN => n3845);
   U8697 : NAND2_X1 port map( A1 => n3845, A2 => n19508, ZN => n3847);
   U8698 : MUX2_X1 port map( A => n3848, B => n3847, S => n5116, Z => n3849);
   U8699 : INV_X1 port map( A => n3855, ZN => n6058);
   U8700 : INV_X1 port map( A => n4670, ZN => n3854);
   U8701 : INV_X1 port map( A => Plaintext(77), ZN => n3851);
   U8702 : XNOR2_X1 port map( A => Key(74), B => Plaintext(74), ZN => n4669);
   U8703 : INV_X1 port map( A => n4669, ZN => n4828);
   U8704 : INV_X1 port map( A => n4214, ZN => n4673);
   U8705 : INV_X1 port map( A => n5258, ZN => n4668);
   U8706 : NOR2_X1 port map( A1 => n4827, A2 => n4829, ZN => n4213);
   U8707 : INV_X1 port map( A => n4213, ZN => n3852);
   U8708 : OAI211_X1 port map( C1 => n4670, C2 => n4673, A => n4668, B => n3852
                           , ZN => n3853);
   U8709 : NAND3_X1 port map( A1 => n6058, A2 => n906, A3 => n6057, ZN => n3866
                           );
   U8710 : XNOR2_X1 port map( A => Key(99), B => Plaintext(99), ZN => n5081);
   U8711 : XNOR2_X1 port map( A => Key(97), B => Plaintext(97), ZN => n4719);
   U8712 : INV_X1 port map( A => n4719, ZN => n5074);
   U8713 : XNOR2_X1 port map( A => Key(96), B => Plaintext(96), ZN => n5079);
   U8714 : XNOR2_X1 port map( A => Key(100), B => Plaintext(100), ZN => n5077);
   U8715 : INV_X1 port map( A => n5077, ZN => n4081);
   U8718 : INV_X1 port map( A => Plaintext(95), ZN => n3856);
   U8719 : INV_X1 port map( A => Plaintext(90), ZN => n3857);
   U8721 : INV_X1 port map( A => Plaintext(91), ZN => n3858);
   U8722 : OAI211_X1 port map( C1 => n5093, C2 => n4788, A => n3859, B => n2461
                           , ZN => n3862);
   U8723 : INV_X1 port map( A => Plaintext(94), ZN => n3860);
   U8724 : XNOR2_X1 port map( A => n3860, B => Key(94), ZN => n5094);
   U8725 : INV_X1 port map( A => n5094, ZN => n4783);
   U8726 : OAI21_X1 port map( B1 => n5098, B2 => n4783, A => n5092, ZN => n3861
                           );
   U8728 : NAND3_X1 port map( A1 => n6064, A2 => n20670, A3 => n6059, ZN => 
                           n3864);
   U8729 : NAND4_X2 port map( A1 => n3865, A2 => n3867, A3 => n3866, A4 => 
                           n3864, ZN => n7201);
   U8730 : XNOR2_X1 port map( A => n7201, B => n2263, ZN => n3902);
   U8731 : INV_X1 port map( A => Plaintext(32), ZN => n3868);
   U8732 : XNOR2_X1 port map( A => n3868, B => Key(32), ZN => n4953);
   U8733 : INV_X1 port map( A => Plaintext(31), ZN => n3869);
   U8735 : INV_X1 port map( A => n4474, ZN => n4913);
   U8736 : INV_X1 port map( A => Plaintext(34), ZN => n3870);
   U8738 : NAND2_X1 port map( A1 => n3871, A2 => n4952, ZN => n3873);
   U8739 : INV_X1 port map( A => n4911, ZN => n4140);
   U8740 : OAI21_X1 port map( B1 => n4912, B2 => n4913, A => n4140, ZN => n3872
                           );
   U8742 : NAND2_X1 port map( A1 => n4021, A2 => n4928, ZN => n4978);
   U8743 : INV_X1 port map( A => Plaintext(18), ZN => n3875);
   U8744 : NAND2_X1 port map( A1 => n4131, A2 => n4296, ZN => n4980);
   U8745 : XNOR2_X1 port map( A => Key(22), B => Plaintext(22), ZN => n4974);
   U8746 : INV_X1 port map( A => n4297, ZN => n4932);
   U8747 : MUX2_X1 port map( A => n4974, B => n4932, S => n4131, Z => n3879);
   U8748 : INV_X1 port map( A => n4978, ZN => n3877);
   U8749 : AND2_X1 port map( A1 => n4979, A2 => n4928, ZN => n3876);
   U8750 : INV_X1 port map( A => n4622, ZN => n4290);
   U8751 : XNOR2_X1 port map( A => Key(4), B => Plaintext(4), ZN => n4285);
   U8752 : INV_X1 port map( A => n4285, ZN => n3882);
   U8753 : INV_X1 port map( A => Plaintext(0), ZN => n3880);
   U8754 : INV_X1 port map( A => n4169, ZN => n4621);
   U8755 : AOI21_X1 port map( B1 => n4630, B2 => n4621, A => n4623, ZN => n3886
                           );
   U8756 : INV_X1 port map( A => Plaintext(2), ZN => n3881);
   U8757 : NAND2_X1 port map( A1 => n4290, A2 => n4171, ZN => n3884);
   U8758 : XNOR2_X1 port map( A => Key(1), B => Plaintext(1), ZN => n4626);
   U8759 : INV_X1 port map( A => n4626, ZN => n4170);
   U8760 : NAND2_X1 port map( A1 => n4170, A2 => n4623, ZN => n3883);
   U8761 : AOI21_X1 port map( B1 => n3884, B2 => n3883, A => n3882, ZN => n3885
                           );
   U8762 : XNOR2_X1 port map( A => Key(7), B => Plaintext(7), ZN => n4324);
   U8763 : INV_X1 port map( A => n4324, ZN => n4647);
   U8764 : XNOR2_X1 port map( A => Key(6), B => Plaintext(6), ZN => n4318);
   U8765 : INV_X1 port map( A => n4318, ZN => n4646);
   U8766 : NAND2_X1 port map( A1 => n4647, A2 => n4646, ZN => n3888);
   U8767 : XNOR2_X2 port map( A => Key(8), B => Plaintext(8), ZN => n4640);
   U8768 : INV_X1 port map( A => n4640, ZN => n4648);
   U8769 : INV_X1 port map( A => Plaintext(11), ZN => n3887);
   U8770 : XNOR2_X1 port map( A => n3887, B => Key(11), ZN => n4317);
   U8771 : MUX2_X1 port map( A => n3888, B => n4648, S => n4325, Z => n3891);
   U8773 : INV_X1 port map( A => n4125, ZN => n4641);
   U8774 : NAND2_X1 port map( A1 => n4319, A2 => n4324, ZN => n4323);
   U8775 : INV_X1 port map( A => n4323, ZN => n3889);
   U8776 : OAI21_X1 port map( B1 => n4641, B2 => n4325, A => n3889, ZN => n3890
                           );
   U8777 : XNOR2_X1 port map( A => Key(24), B => Plaintext(24), ZN => n4114);
   U8778 : INV_X1 port map( A => n4114, ZN => n4470);
   U8779 : INV_X1 port map( A => n4118, ZN => n4941);
   U8780 : INV_X1 port map( A => n4945, ZN => n4467);
   U8781 : INV_X1 port map( A => n4940, ZN => n4117);
   U8782 : INV_X1 port map( A => Plaintext(28), ZN => n3893);
   U8783 : XNOR2_X1 port map( A => n3893, B => Key(28), ZN => n4946);
   U8784 : NAND3_X1 port map( A1 => n4946, A2 => n4945, A3 => n4947, ZN => 
                           n3894);
   U8785 : OAI211_X1 port map( C1 => n3896, C2 => n4947, A => n3895, B => n3894
                           , ZN => n5795);
   U8786 : XNOR2_X1 port map( A => Key(15), B => Plaintext(15), ZN => n3897);
   U8788 : NAND2_X1 port map( A1 => n4988, A2 => n4982, ZN => n4005);
   U8789 : INV_X1 port map( A => n3897, ZN => n4983);
   U8790 : XNOR2_X1 port map( A => Key(13), B => Plaintext(13), ZN => n4618);
   U8791 : NAND2_X1 port map( A1 => n4983, A2 => n4618, ZN => n3898);
   U8793 : INV_X1 port map( A => n4306, ZN => n4003);
   U8794 : XNOR2_X1 port map( A => Key(16), B => Plaintext(16), ZN => n4305);
   U8795 : NAND2_X1 port map( A1 => n4003, A2 => n4305, ZN => n3900);
   U8796 : NAND2_X1 port map( A1 => n4988, A2 => n4306, ZN => n3899);
   U8797 : INV_X1 port map( A => n5017, ZN => n5014);
   U8799 : INV_X1 port map( A => n5018, ZN => n4736);
   U8800 : XNOR2_X1 port map( A => Key(139), B => Plaintext(139), ZN => n4277);
   U8801 : INV_X1 port map( A => n4277, ZN => n5012);
   U8802 : NAND2_X1 port map( A1 => n5012, A2 => n4734, ZN => n3903);
   U8804 : INV_X1 port map( A => n4734, ZN => n3904);
   U8805 : XNOR2_X1 port map( A => Key(138), B => Plaintext(138), ZN => n4110);
   U8806 : INV_X1 port map( A => n4110, ZN => n4554);
   U8807 : INV_X1 port map( A => Plaintext(161), ZN => n3906);
   U8808 : XNOR2_X2 port map( A => n3906, B => Key(161), ZN => n4370);
   U8809 : INV_X1 port map( A => n4576, ZN => n4570);
   U8811 : XNOR2_X1 port map( A => Key(157), B => Plaintext(157), ZN => n4507);
   U8812 : NAND2_X1 port map( A1 => n4507, A2 => n4575, ZN => n4510);
   U8813 : NAND3_X1 port map( A1 => n4510, A2 => n4576, A3 => n3907, ZN => 
                           n3910);
   U8814 : INV_X1 port map( A => n4370, ZN => n4511);
   U8815 : INV_X1 port map( A => Plaintext(156), ZN => n3908);
   U8816 : INV_X1 port map( A => n4571, ZN => n4573);
   U8817 : NAND3_X1 port map( A1 => n4511, A2 => n4372, A3 => n4573, ZN => 
                           n3909);
   U8818 : INV_X1 port map( A => n6048, ZN => n5139);
   U8819 : NAND2_X1 port map( A1 => n5328, A2 => n5139, ZN => n3920);
   U8820 : INV_X1 port map( A => Plaintext(149), ZN => n3911);
   U8821 : XNOR2_X1 port map( A => n3911, B => Key(149), ZN => n5005);
   U8822 : INV_X1 port map( A => n5005, ZN => n4746);
   U8823 : INV_X1 port map( A => n5010, ZN => n3912);
   U8824 : NAND2_X1 port map( A1 => n4746, A2 => n3912, ZN => n4557);
   U8826 : INV_X1 port map( A => n4206, ZN => n4561);
   U8828 : NAND2_X1 port map( A1 => n4746, A2 => n4745, ZN => n3913);
   U8829 : NAND2_X1 port map( A1 => n4561, A2 => n3913, ZN => n3915);
   U8830 : NAND2_X1 port map( A1 => n4248, A2 => n4744, ZN => n3914);
   U8831 : INV_X1 port map( A => n6049, ZN => n5557);
   U8832 : XNOR2_X2 port map( A => Key(153), B => Plaintext(153), ZN => n4504);
   U8833 : MUX2_X1 port map( A => n4756, B => n4504, S => n4752, Z => n3918);
   U8834 : INV_X1 port map( A => n4504, ZN => n4563);
   U8835 : XNOR2_X1 port map( A => Key(151), B => Plaintext(151), ZN => n4565);
   U8836 : INV_X1 port map( A => n4565, ZN => n4755);
   U8837 : INV_X1 port map( A => Plaintext(150), ZN => n3916);
   U8838 : NAND2_X1 port map( A1 => n4754, A2 => n4504, ZN => n3917);
   U8839 : INV_X1 port map( A => n4567, ZN => n4198);
   U8840 : AOI21_X1 port map( B1 => n3920, B2 => n3919, A => n6052, ZN => n3936
                           );
   U8841 : XNOR2_X1 port map( A => Key(171), B => Plaintext(171), ZN => n4518);
   U8842 : INV_X1 port map( A => n4518, ZN => n3922);
   U8843 : INV_X1 port map( A => Plaintext(169), ZN => n3921);
   U8844 : NAND2_X1 port map( A1 => n3922, A2 => n4517, ZN => n4340);
   U8845 : INV_X1 port map( A => n4340, ZN => n3924);
   U8847 : INV_X1 port map( A => Plaintext(170), ZN => n3923);
   U8848 : OAI21_X1 port map( B1 => n3924, B2 => n4522, A => n4343, ZN => n3928
                           );
   U8849 : INV_X1 port map( A => n4517, ZN => n4520);
   U8850 : INV_X1 port map( A => Plaintext(172), ZN => n3926);
   U8851 : XNOR2_X1 port map( A => n3926, B => Key(172), ZN => n4342);
   U8852 : NAND2_X1 port map( A1 => n3943, A2 => n4342, ZN => n3927);
   U8853 : AND2_X2 port map( A1 => n3928, A2 => n3927, ZN => n5559);
   U8854 : NAND2_X1 port map( A1 => n3929, A2 => n6048, ZN => n4995);
   U8856 : INV_X1 port map( A => n3948, ZN => n4542);
   U8858 : NAND2_X1 port map( A1 => n4539, A2 => n4350, ZN => n3931);
   U8859 : INV_X1 port map( A => Plaintext(164), ZN => n3930);
   U8860 : OAI211_X1 port map( C1 => n4542, C2 => n4539, A => n3931, B => n4347
                           , ZN => n3933);
   U8861 : NAND2_X1 port map( A1 => n5559, A2 => n6050, ZN => n3934);
   U8862 : OAI22_X1 port map( A1 => n6054, A2 => n4995, B1 => n3934, B2 => 
                           n3351, ZN => n3935);
   U8863 : XNOR2_X1 port map( A => Key(175), B => Plaintext(175), ZN => n4532);
   U8864 : XNOR2_X1 port map( A => Key(174), B => Plaintext(174), ZN => n4528);
   U8865 : NAND2_X1 port map( A1 => n19524, A2 => n4529, ZN => n3938);
   U8866 : INV_X1 port map( A => Plaintext(179), ZN => n3937);
   U8867 : XNOR2_X2 port map( A => n3937, B => Key(179), ZN => n4633);
   U8868 : OAI211_X1 port map( C1 => n19524, C2 => n4532, A => n3938, B => 
                           n4633, ZN => n5576);
   U8869 : INV_X1 port map( A => n4633, ZN => n4337);
   U8870 : INV_X1 port map( A => Plaintext(178), ZN => n3939);
   U8872 : NAND2_X2 port map( A1 => n5575, A2 => n5576, ZN => n5408);
   U8873 : NAND2_X1 port map( A1 => n4343, A2 => n4516, ZN => n3942);
   U8875 : AND2_X1 port map( A1 => n4520, A2 => n4523, ZN => n3941);
   U8876 : INV_X1 port map( A => n4342, ZN => n4160);
   U8878 : INV_X1 port map( A => n5581, ZN => n5404);
   U8879 : INV_X1 port map( A => Plaintext(182), ZN => n3944);
   U8880 : INV_X1 port map( A => Plaintext(181), ZN => n3945);
   U8881 : INV_X1 port map( A => n4313, ZN => n4603);
   U8882 : INV_X1 port map( A => Plaintext(183), ZN => n3946);
   U8883 : XNOR2_X1 port map( A => n3946, B => Key(183), ZN => n4152);
   U8884 : INV_X1 port map( A => Plaintext(180), ZN => n3947);
   U8885 : INV_X1 port map( A => n4548, ZN => n4353);
   U8886 : XNOR2_X1 port map( A => Key(185), B => Plaintext(185), ZN => n4602);
   U8887 : XNOR2_X1 port map( A => Key(184), B => Plaintext(184), ZN => n4601);
   U8888 : NAND2_X1 port map( A1 => n4355, A2 => n4601, ZN => n4312);
   U8889 : INV_X1 port map( A => n4602, ZN => n4607);
   U8890 : OAI211_X1 port map( C1 => n4541, C2 => n4349, A => n4542, B => n4539
                           , ZN => n3950);
   U8891 : NAND2_X1 port map( A1 => n3950, A2 => n3949, ZN => n3951);
   U8892 : XNOR2_X1 port map( A => Key(189), B => Plaintext(189), ZN => n4176);
   U8893 : INV_X1 port map( A => n4176, ZN => n4011);
   U8894 : INV_X1 port map( A => Plaintext(186), ZN => n3952);
   U8895 : XNOR2_X1 port map( A => n3952, B => Key(186), ZN => n4611);
   U8896 : NAND2_X1 port map( A1 => n4011, A2 => n4611, ZN => n4010);
   U8897 : INV_X1 port map( A => Plaintext(187), ZN => n3953);
   U8898 : INV_X1 port map( A => n4611, ZN => n4364);
   U8899 : XNOR2_X1 port map( A => Key(190), B => Plaintext(190), ZN => n4013);
   U8900 : NAND2_X1 port map( A1 => n1537, A2 => n748, ZN => n3954);
   U8901 : INV_X1 port map( A => n4365, ZN => n4609);
   U8902 : OR2_X1 port map( A1 => n4010, A2 => n748, ZN => n5574);
   U8903 : NAND2_X1 port map( A1 => n5573, A2 => n5574, ZN => n5405);
   U8904 : AND2_X1 port map( A1 => n4169, A2 => n4623, ZN => n4291);
   U8905 : OAI21_X1 port map( B1 => n4170, B2 => n4621, A => n4171, ZN => n3956
                           );
   U8907 : INV_X1 port map( A => n4171, ZN => n4631);
   U8908 : AOI21_X1 port map( B1 => n4018, B2 => n4627, A => n4285, ZN => n3957
                           );
   U8910 : XNOR2_X1 port map( A => n6693, B => n7304, ZN => n3962);
   U8911 : XNOR2_X1 port map( A => n3963, B => n3962, ZN => n4065);
   U8913 : INV_X1 port map( A => n4968, ZN => n3965);
   U8914 : INV_X1 port map( A => Plaintext(42), ZN => n3964);
   U8915 : XNOR2_X1 port map( A => n3964, B => Key(42), ZN => n4970);
   U8916 : NAND2_X1 port map( A1 => n3965, A2 => n4970, ZN => n4967);
   U8917 : AND2_X1 port map( A1 => n4969, A2 => n4968, ZN => n4483);
   U8919 : NAND2_X1 port map( A1 => n4965, A2 => n4479, ZN => n3966);
   U8920 : NAND2_X1 port map( A1 => n4483, A2 => n3966, ZN => n3968);
   U8922 : OAI211_X1 port map( C1 => n4967, C2 => n3967, A => n3968, B => n4966
                           , ZN => n5978);
   U8923 : INV_X1 port map( A => Plaintext(41), ZN => n3969);
   U8924 : XNOR2_X2 port map( A => n3969, B => Key(41), ZN => n4899);
   U8925 : NAND2_X1 port map( A1 => n4377, A2 => n4899, ZN => n3973);
   U8926 : INV_X1 port map( A => Plaintext(37), ZN => n3970);
   U8928 : XNOR2_X1 port map( A => Key(39), B => Plaintext(39), ZN => n4894);
   U8929 : NAND2_X1 port map( A1 => n4960, A2 => n4894, ZN => n3972);
   U8930 : INV_X1 port map( A => Plaintext(40), ZN => n3971);
   U8931 : AOI21_X1 port map( B1 => n3973, B2 => n3972, A => n4962, ZN => n3976
                           );
   U8932 : AOI21_X1 port map( B1 => n3974, B2 => n4136, A => n3231, ZN => n3975
                           );
   U8933 : NOR2_X1 port map( A1 => n5978, A2 => n6072, ZN => n3993);
   U8934 : NOR2_X1 port map( A1 => n4840, A2 => n4657, ZN => n4421);
   U8935 : INV_X1 port map( A => Plaintext(65), ZN => n3982);
   U8937 : NAND2_X1 port map( A1 => n289, A2 => n4652, ZN => n3986);
   U8938 : INV_X1 port map( A => Plaintext(60), ZN => n3983);
   U8939 : XNOR2_X1 port map( A => n3983, B => Key(60), ZN => n4867);
   U8940 : INV_X1 port map( A => Plaintext(62), ZN => n3984);
   U8941 : NOR2_X1 port map( A1 => n6069, A2 => n5320, ZN => n3992);
   U8942 : INV_X1 port map( A => Plaintext(49), ZN => n3987);
   U8943 : XNOR2_X1 port map( A => n3987, B => Key(49), ZN => n4232);
   U8944 : INV_X1 port map( A => Plaintext(48), ZN => n3988);
   U8945 : XNOR2_X1 port map( A => n3988, B => Key(48), ZN => n4497);
   U8946 : INV_X1 port map( A => n4907, ZN => n4493);
   U8947 : XNOR2_X1 port map( A => Key(52), B => Plaintext(52), ZN => n4855);
   U8948 : NAND2_X1 port map( A1 => n4493, A2 => n4855, ZN => n3989);
   U8951 : INV_X1 port map( A => n3996, ZN => n4853);
   U8952 : INV_X1 port map( A => n176, ZN => n4485);
   U8953 : XNOR2_X1 port map( A => Key(55), B => Plaintext(55), ZN => n4685);
   U8954 : MUX2_X1 port map( A => n4851, B => n4682, S => n4685, Z => n3998);
   U8955 : INV_X1 port map( A => Plaintext(58), ZN => n3994);
   U8957 : XNOR2_X1 port map( A => Key(54), B => Plaintext(54), ZN => n4391);
   U8958 : NAND2_X1 port map( A1 => n178, A2 => n4391, ZN => n4224);
   U8960 : NAND2_X1 port map( A1 => n6068, A2 => n209, ZN => n4000);
   U8961 : OAI21_X1 port map( B1 => n4118, B2 => n4940, A => n4470, ZN => n4002
                           );
   U8962 : INV_X1 port map( A => n4305, ZN => n4989);
   U8963 : MUX2_X1 port map( A => n4005, B => n4004, S => n19822, Z => n4009);
   U8964 : INV_X1 port map( A => n4618, ZN => n4006);
   U8965 : NAND2_X1 port map( A1 => n4988, A2 => n4618, ZN => n4985);
   U8966 : NAND2_X1 port map( A1 => n4007, A2 => n4985, ZN => n4008);
   U8967 : INV_X1 port map( A => n5395, ZN => n5367);
   U8968 : NAND2_X1 port map( A1 => n1537, A2 => n4615, ZN => n4366);
   U8970 : NAND2_X1 port map( A1 => n4012, A2 => n4011, ZN => n4014);
   U8971 : INV_X1 port map( A => n4614, ZN => n4177);
   U8973 : NAND2_X1 port map( A1 => n4640, A2 => n4319, ZN => n4015);
   U8974 : OAI21_X1 port map( B1 => n4641, B2 => n4640, A => n4015, ZN => n4016
                           );
   U8975 : INV_X1 port map( A => n4317, ZN => n4642);
   U8976 : NAND2_X1 port map( A1 => n5368, A2 => n5322, ZN => n4019);
   U8977 : INV_X1 port map( A => n4296, ZN => n4927);
   U8978 : INV_X1 port map( A => n4928, ZN => n4298);
   U8979 : OAI211_X1 port map( C1 => n4927, C2 => n4297, A => n4020, B => n4298
                           , ZN => n4024);
   U8980 : NAND3_X1 port map( A1 => n4975, A2 => n4928, A3 => n4131, ZN => 
                           n4023);
   U8981 : NAND3_X1 port map( A1 => n4932, A2 => n4296, A3 => n4976, ZN => 
                           n4022);
   U8982 : NAND3_X1 port map( A1 => n4282, A2 => n5323, A3 => n5398, ZN => 
                           n4025);
   U8983 : XNOR2_X1 port map( A => n7264, B => n6745, ZN => n4063);
   U8984 : NAND2_X1 port map( A1 => n4796, A2 => n5045, ZN => n4027);
   U8986 : NAND2_X1 port map( A1 => n5042, A2 => n5046, ZN => n4026);
   U8987 : XNOR2_X1 port map( A => Key(115), B => Plaintext(115), ZN => n4440);
   U8988 : INV_X1 port map( A => n4439, ZN => n5048);
   U8989 : INV_X1 port map( A => Plaintext(114), ZN => n4028);
   U8990 : XNOR2_X1 port map( A => Key(119), B => Plaintext(119), ZN => n4088);
   U8991 : INV_X1 port map( A => n4088, ZN => n4698);
   U8992 : INV_X1 port map( A => n6044, ZN => n5144);
   U8994 : NAND2_X1 port map( A1 => n5087, A2 => n5086, ZN => n4032);
   U8996 : INV_X1 port map( A => n5086, ZN => n4802);
   U8997 : INV_X1 port map( A => Plaintext(113), ZN => n4030);
   U8999 : INV_X1 port map( A => n4701, ZN => n4807);
   U9000 : OAI21_X1 port map( B1 => n4032, B2 => n5083, A => n4031, ZN => n4034
                           );
   U9001 : AOI21_X1 port map( B1 => n4032, B2 => n5090, A => n4807, ZN => n4033
                           );
   U9002 : INV_X1 port map( A => Plaintext(132), ZN => n4035);
   U9003 : XNOR2_X1 port map( A => Key(137), B => Plaintext(137), ZN => n4268);
   U9004 : INV_X1 port map( A => n4268, ZN => n5026);
   U9005 : INV_X1 port map( A => Plaintext(134), ZN => n4036);
   U9006 : XNOR2_X1 port map( A => n4036, B => Key(134), ZN => n4094);
   U9007 : INV_X1 port map( A => n4094, ZN => n4761);
   U9008 : NAND2_X1 port map( A1 => n4765, A2 => n4269, ZN => n4037);
   U9009 : AOI21_X1 port map( B1 => n4037, B2 => n4095, A => n4761, ZN => n4038
                           );
   U9010 : INV_X1 port map( A => Plaintext(125), ZN => n4039);
   U9011 : XNOR2_X1 port map( A => n4039, B => Key(125), ZN => n4041);
   U9012 : INV_X1 port map( A => n4041, ZN => n5035);
   U9013 : INV_X1 port map( A => Plaintext(120), ZN => n4040);
   U9014 : XNOR2_X1 port map( A => Key(123), B => Plaintext(123), ZN => n4107);
   U9015 : INV_X1 port map( A => n5031, ZN => n4707);
   U9016 : NAND2_X1 port map( A1 => n4709, A2 => n4707, ZN => n4042);
   U9017 : AND2_X1 port map( A1 => n4107, A2 => n4769, ZN => n5037);
   U9018 : INV_X1 port map( A => n4769, ZN => n4452);
   U9019 : XNOR2_X1 port map( A => Key(105), B => Plaintext(105), ZN => n4048);
   U9020 : INV_X1 port map( A => Plaintext(104), ZN => n4044);
   U9021 : XNOR2_X1 port map( A => n4044, B => Key(104), ZN => n5106);
   U9022 : INV_X1 port map( A => Plaintext(106), ZN => n4045);
   U9024 : INV_X1 port map( A => n5101, ZN => n4077);
   U9025 : MUX2_X1 port map( A => n5105, B => n5102, S => n4077, Z => n4051);
   U9026 : INV_X1 port map( A => Plaintext(107), ZN => n4046);
   U9027 : XNOR2_X2 port map( A => n4046, B => Key(107), ZN => n5107);
   U9028 : XNOR2_X1 port map( A => Key(103), B => Plaintext(103), ZN => n5100);
   U9029 : INV_X1 port map( A => n5100, ZN => n4793);
   U9030 : INV_X1 port map( A => Plaintext(102), ZN => n4047);
   U9031 : XNOR2_X1 port map( A => n4047, B => Key(102), ZN => n5108);
   U9032 : INV_X1 port map( A => n5108, ZN => n5099);
   U9033 : INV_X1 port map( A => n4048, ZN => n4693);
   U9034 : MUX2_X1 port map( A => n4049, B => n5099, S => n4693, Z => n4050);
   U9035 : INV_X1 port map( A => Plaintext(129), ZN => n4053);
   U9036 : XNOR2_X1 port map( A => Key(131), B => Plaintext(131), ZN => n4056);
   U9037 : INV_X1 port map( A => n4056, ZN => n5055);
   U9038 : XNOR2_X1 port map( A => Key(126), B => Plaintext(126), ZN => n4058);
   U9039 : INV_X1 port map( A => Plaintext(130), ZN => n4054);
   U9040 : XNOR2_X1 port map( A => n4054, B => Key(130), ZN => n4445);
   U9041 : INV_X1 port map( A => Plaintext(128), ZN => n4055);
   U9042 : XNOR2_X1 port map( A => n4055, B => Key(128), ZN => n4060);
   U9043 : INV_X1 port map( A => n4060, ZN => n5059);
   U9044 : NAND3_X1 port map( A1 => n4585, A2 => n5059, A3 => n5058, ZN => 
                           n4057);
   U9045 : INV_X1 port map( A => n4058, ZN => n5056);
   U9046 : INV_X1 port map( A => Plaintext(127), ZN => n4059);
   U9047 : INV_X1 port map( A => n5052, ZN => n4739);
   U9048 : NAND2_X1 port map( A1 => n6046, A2 => n5309, ZN => n4061);
   U9049 : NOR2_X1 port map( A1 => n4061, A2 => n6044, ZN => n4062);
   U9050 : XNOR2_X1 port map( A => n4063, B => n7345, ZN => n4064);
   U9051 : XNOR2_X1 port map( A => n4065, B => n4064, ZN => n8061);
   U9052 : INV_X1 port map( A => n4418, ZN => n4066);
   U9053 : INV_X1 port map( A => n5093, ZN => n4715);
   U9054 : INV_X1 port map( A => n4405, ZN => n4713);
   U9055 : NAND3_X1 port map( A1 => n4788, A2 => n4715, A3 => n2460, ZN => 
                           n4069);
   U9057 : OAI21_X1 port map( B1 => n4214, B2 => n4827, A => n4824, ZN => n4072
                           );
   U9058 : INV_X1 port map( A => n4824, ZN => n4426);
   U9059 : NAND2_X1 port map( A1 => n4426, A2 => n4829, ZN => n4071);
   U9060 : AND2_X1 port map( A1 => n4072, A2 => n4071, ZN => n4075);
   U9061 : NAND2_X1 port map( A1 => n4426, A2 => n4214, ZN => n4073);
   U9062 : AOI21_X1 port map( B1 => n4425, B2 => n4073, A => n4668, ZN => n4074
                           );
   U9063 : INV_X1 port map( A => n5434, ZN => n5995);
   U9064 : AOI21_X1 port map( B1 => n5998, B2 => n5997, A => n5995, ZN => n4087
                           );
   U9065 : AOI21_X1 port map( B1 => n4076, B2 => n5108, A => n5102, ZN => n4079
                           );
   U9066 : NAND2_X1 port map( A1 => n4793, A2 => n5108, ZN => n4449);
   U9067 : NAND2_X1 port map( A1 => n5998, A2 => n5434, ZN => n4080);
   U9069 : NAND2_X1 port map( A1 => n4081, A2 => n5075, ZN => n4082);
   U9070 : MUX2_X1 port map( A => n4083, B => n4082, S => n5080, Z => n4086);
   U9071 : NAND2_X1 port map( A1 => n4084, A2 => n4457, ZN => n4085);
   U9072 : INV_X1 port map( A => n6000, ZN => n6002);
   U9073 : NAND2_X1 port map( A1 => n4088, A2 => n5045, ZN => n4089);
   U9074 : NAND2_X1 port map( A1 => n4698, A2 => n5046, ZN => n4798);
   U9075 : INV_X1 port map( A => n5990, ZN => n5708);
   U9076 : MUX2_X1 port map( A => n20202, B => n5086, S => n5087, Z => n4093);
   U9077 : NAND2_X1 port map( A1 => n4090, A2 => n19776, ZN => n4092);
   U9078 : NOR2_X1 port map( A1 => n4801, A2 => n5083, ZN => n4091);
   U9079 : AOI21_X1 port map( B1 => n4093, B2 => n4092, A => n4091, ZN => n5711
                           );
   U9080 : NAND2_X1 port map( A1 => n4765, A2 => n4095, ZN => n4098);
   U9081 : INV_X1 port map( A => n4095, ZN => n4764);
   U9083 : NAND3_X1 port map( A1 => n5025, A2 => n4761, A3 => n5024, ZN => 
                           n4097);
   U9084 : NAND2_X1 port map( A1 => n20461, A2 => n5059, ZN => n4099);
   U9085 : AOI21_X1 port map( B1 => n5054, B2 => n4099, A => n5058, ZN => n4104
                           );
   U9086 : INV_X1 port map( A => n4100, ZN => n5057);
   U9087 : NAND3_X1 port map( A1 => n5057, A2 => n5058, A3 => n873, ZN => n4101
                           );
   U9088 : NAND2_X1 port map( A1 => n4102, A2 => n4101, ZN => n4103);
   U9089 : NAND2_X1 port map( A1 => n4708, A2 => n4107, ZN => n4105);
   U9090 : OAI21_X1 port map( B1 => n4107, B2 => n4769, A => n4105, ZN => n4106
                           );
   U9091 : NAND2_X1 port map( A1 => n4106, A2 => n5032, ZN => n4109);
   U9092 : NAND2_X1 port map( A1 => n303, A2 => n153, ZN => n4108);
   U9093 : INV_X1 port map( A => n5815, ZN => n5709);
   U9094 : OAI21_X1 port map( B1 => n4734, B2 => n4277, A => n4554, ZN => n4111
                           );
   U9095 : INV_X1 port map( A => n5276, ZN => n5986);
   U9096 : NAND2_X1 port map( A1 => n5986, A2 => n5989, ZN => n4112);
   U9097 : XNOR2_X1 port map( A => n6711, B => n7390, ZN => n7016);
   U9098 : AND2_X1 port map( A1 => n4887, A2 => n4946, ZN => n4471);
   U9099 : NAND2_X1 port map( A1 => n4114, A2 => n4118, ZN => n4943);
   U9100 : INV_X1 port map( A => n4943, ZN => n4115);
   U9101 : AOI22_X1 port map( A1 => n4467, A2 => n4471, B1 => n4115, B2 => 
                           n4947, ZN => n4121);
   U9102 : OAI21_X1 port map( B1 => n4467, B2 => n4117, A => n4116, ZN => n4119
                           );
   U9104 : INV_X1 port map( A => n4886, ZN => n4888);
   U9105 : NAND2_X1 port map( A1 => n4119, A2 => n4888, ZN => n4120);
   U9106 : NAND2_X1 port map( A1 => n4003, A2 => n19822, ZN => n4122);
   U9107 : NAND2_X1 port map( A1 => n4620, A2 => n4122, ZN => n4123);
   U9108 : NAND2_X1 port map( A1 => n4125, A2 => n4640, ZN => n4126);
   U9109 : NAND2_X1 port map( A1 => n4647, A2 => n4125, ZN => n4128);
   U9110 : MUX2_X1 port map( A => n4128, B => n4318, S => n4127, Z => n4129);
   U9111 : OAI21_X1 port map( B1 => n4130, B2 => n4642, A => n4129, ZN => n5968
                           );
   U9112 : INV_X1 port map( A => n5968, ZN => n5525);
   U9114 : NAND2_X1 port map( A1 => n4298, A2 => n4975, ZN => n4133);
   U9115 : NAND2_X1 port map( A1 => n4296, A2 => n4297, ZN => n4132);
   U9116 : MUX2_X1 port map( A => n4133, B => n4132, S => n4976, Z => n4134);
   U9117 : OAI21_X2 port map( B1 => n4135, B2 => n4297, A => n4134, ZN => n5697
                           );
   U9118 : INV_X1 port map( A => n5697, ZN => n5294);
   U9120 : NAND2_X1 port map( A1 => n4899, A2 => n4892, ZN => n4137);
   U9121 : INV_X1 port map( A => n4912, ZN => n4914);
   U9124 : NAND2_X1 port map( A1 => n4474, A2 => n4911, ZN => n4141);
   U9126 : NAND2_X1 port map( A1 => n4952, A2 => n4954, ZN => n4142);
   U9127 : INV_X1 port map( A => n4953, ZN => n4950);
   U9128 : OR2_X1 port map( A1 => n4144, A2 => n4954, ZN => n5522);
   U9129 : AOI21_X1 port map( B1 => n4146, B2 => n4646, A => n4640, ZN => n4150
                           );
   U9131 : NAND3_X1 port map( A1 => n4641, A2 => n4325, A3 => n4640, ZN => 
                           n4147);
   U9133 : NAND2_X1 port map( A1 => n4354, A2 => n4547, ZN => n4151);
   U9135 : NAND2_X1 port map( A1 => n19524, A2 => n4532, ZN => n4158);
   U9136 : NAND2_X1 port map( A1 => n4186, A2 => n4637, ZN => n4157);
   U9137 : NAND2_X1 port map( A1 => n4516, A2 => n4342, ZN => n4527);
   U9138 : AOI21_X1 port map( B1 => n4527, B2 => n4522, A => n4523, ZN => n4164
                           );
   U9139 : NAND3_X1 port map( A1 => n4343, A2 => n4516, A3 => n4160, ZN => 
                           n4162);
   U9140 : NAND2_X1 port map( A1 => n4162, A2 => n4161, ZN => n4163);
   U9142 : OAI21_X1 port map( B1 => n5645, B2 => n5443, A => n4165, ZN => n4777
                           );
   U9143 : INV_X1 port map( A => n4623, ZN => n4166);
   U9144 : AOI21_X1 port map( B1 => n4166, B2 => n4169, A => n20143, ZN => 
                           n4175);
   U9145 : NAND2_X1 port map( A1 => n4288, A2 => n4167, ZN => n4174);
   U9146 : INV_X1 port map( A => n4291, ZN => n4168);
   U9147 : OAI21_X1 port map( B1 => n4170, B2 => n4169, A => n4168, ZN => n4172
                           );
   U9148 : NAND3_X1 port map( A1 => n4613, A2 => n4364, A3 => n748, ZN => n4178
                           );
   U9149 : NAND2_X1 port map( A1 => n4179, A2 => n5442, ZN => n4180);
   U9150 : AOI22_X1 port map( A1 => n4777, A2 => n5649, B1 => n4180, B2 => 
                           n5443, ZN => n6352);
   U9151 : INV_X1 port map( A => n6352, ZN => n7298);
   U9152 : XNOR2_X1 port map( A => n7298, B => n7196, ZN => n6858);
   U9153 : XNOR2_X1 port map( A => n7016, B => n6858, ZN => n4247);
   U9154 : NAND2_X1 port map( A1 => n5798, A2 => n5428, ZN => n5301);
   U9155 : INV_X1 port map( A => n5795, ZN => n5791);
   U9156 : AOI21_X1 port map( B1 => n4182, B2 => n4181, A => n5300, ZN => n4183
                           );
   U9157 : INV_X1 port map( A => n4187, ZN => n4339);
   U9158 : NAND2_X1 port map( A1 => n4516, A2 => n4339, ZN => n4191);
   U9159 : NAND2_X1 port map( A1 => n4517, A2 => n4187, ZN => n4188);
   U9160 : OAI211_X1 port map( C1 => n4523, C2 => n4522, A => n4188, B => n4343
                           , ZN => n4190);
   U9161 : NAND2_X1 port map( A1 => n4575, A2 => n4576, ZN => n4257);
   U9162 : NAND2_X1 port map( A1 => n4570, A2 => n4574, ZN => n4192);
   U9163 : AND2_X1 port map( A1 => n4257, A2 => n4192, ZN => n4195);
   U9164 : NAND2_X1 port map( A1 => n20190, A2 => n4575, ZN => n4193);
   U9165 : OAI21_X1 port map( B1 => n4372, B2 => n4507, A => n4193, ZN => n4194
                           );
   U9166 : INV_X1 port map( A => n5424, ZN => n5675);
   U9167 : NAND2_X1 port map( A1 => n4567, A2 => n4756, ZN => n4196);
   U9168 : NAND2_X1 port map( A1 => n4196, A2 => n4504, ZN => n4197);
   U9169 : NAND2_X1 port map( A1 => n4198, A2 => n4752, ZN => n4758);
   U9170 : NAND2_X1 port map( A1 => n4347, A2 => n4199, ZN => n4201);
   U9171 : MUX2_X1 port map( A => n4201, B => n4200, S => n4541, Z => n4202);
   U9172 : NAND3_X1 port map( A1 => n5424, A2 => n5669, A3 => n5670, ZN => 
                           n4211);
   U9173 : INV_X1 port map( A => n4204, ZN => n5003);
   U9174 : NAND2_X1 port map( A1 => n4744, A2 => n4745, ZN => n4207);
   U9175 : NAND2_X1 port map( A1 => n4207, A2 => n4248, ZN => n4208);
   U9176 : NAND2_X1 port map( A1 => n5424, A2 => n5279, ZN => n4210);
   U9177 : XNOR2_X1 port map( A => n6708, B => n6489, ZN => n4245);
   U9178 : NAND2_X1 port map( A1 => n4213, A2 => n4214, ZN => n4219);
   U9179 : AND2_X1 port map( A1 => n4214, A2 => n4669, ZN => n4823);
   U9180 : NAND2_X1 port map( A1 => n4823, A2 => n19688, ZN => n4218);
   U9181 : INV_X1 port map( A => n4829, ZN => n4215);
   U9182 : OAI21_X1 port map( B1 => n4824, B2 => n4827, A => n4215, ZN => n4216
                           );
   U9183 : NAND2_X1 port map( A1 => n4216, A2 => n4828, ZN => n4217);
   U9184 : INV_X1 port map( A => n4220, ZN => n4841);
   U9185 : NAND3_X1 port map( A1 => n4659, A2 => n2601, A3 => n4221, ZN => 
                           n4222);
   U9186 : AND2_X1 port map( A1 => n6016, A2 => n6022, ZN => n5124);
   U9187 : INV_X1 port map( A => n4685, ZN => n4484);
   U9188 : OAI211_X1 port map( C1 => n4484, C2 => n177, A => n4224, B => n4853,
                           ZN => n4225);
   U9189 : INV_X1 port map( A => n5825, ZN => n5824);
   U9190 : NAND2_X1 port map( A1 => n5124, A2 => n5824, ZN => n4243);
   U9191 : NAND2_X1 port map( A1 => n4381, A2 => n4651, ZN => n4228);
   U9192 : INV_X1 port map( A => n4228, ZN => n4231);
   U9193 : OAI21_X1 port map( B1 => n4652, B2 => n4865, A => n20356, ZN => 
                           n4230);
   U9194 : MUX2_X1 port map( A => n4228, B => n4227, S => n896, Z => n4229);
   U9195 : INV_X1 port map( A => n4232, ZN => n4492);
   U9196 : INV_X1 port map( A => n4497, ZN => n4901);
   U9197 : OAI21_X1 port map( B1 => n4492, B2 => n4901, A => n4378, ZN => n4905
                           );
   U9198 : NAND2_X1 port map( A1 => n4493, A2 => n4499, ZN => n4236);
   U9199 : NAND2_X1 port map( A1 => n4492, A2 => n4856, ZN => n4857);
   U9200 : INV_X1 port map( A => n4857, ZN => n4235);
   U9201 : NAND2_X1 port map( A1 => n4855, A2 => n4860, ZN => n4234);
   U9202 : NAND3_X1 port map( A1 => n5823, A2 => n5825, A3 => n3569, ZN => 
                           n4242);
   U9203 : INV_X1 port map( A => n4965, ZN => n4383);
   U9204 : INV_X1 port map( A => n4482, ZN => n4919);
   U9205 : INV_X1 port map( A => n4969, ZN => n4921);
   U9206 : OAI211_X1 port map( C1 => n4965, C2 => n4479, A => n4921, B => 
                           n19507, ZN => n4238);
   U9207 : OAI21_X1 port map( B1 => n4383, B2 => n4968, A => n4969, ZN => n4237
                           );
   U9208 : INV_X1 port map( A => n6017, ZN => n5827);
   U9209 : NAND2_X1 port map( A1 => n5827, A2 => n5825, ZN => n4241);
   U9210 : NAND3_X1 port map( A1 => n3569, A2 => n6017, A3 => n6022, ZN => 
                           n4240);
   U9211 : NAND4_X2 port map( A1 => n4243, A2 => n4242, A3 => n4241, A4 => 
                           n4240, ZN => n7013);
   U9212 : XNOR2_X1 port map( A => n7013, B => n20682, ZN => n4244);
   U9213 : XNOR2_X1 port map( A => n4245, B => n4244, ZN => n4246);
   U9214 : INV_X1 port map( A => n4750, ZN => n5007);
   U9215 : NAND2_X1 port map( A1 => n4248, A2 => n5007, ZN => n4253);
   U9216 : INV_X1 port map( A => n4744, ZN => n5006);
   U9217 : NAND3_X1 port map( A1 => n4559, A2 => n5006, A3 => n4746, ZN => 
                           n4251);
   U9218 : INV_X1 port map( A => n4350, ZN => n4537);
   U9220 : INV_X1 port map( A => n4539, ZN => n4255);
   U9221 : OAI21_X1 port map( B1 => n4370, B2 => n4372, A => n20190, ZN => 
                           n4263);
   U9222 : INV_X1 port map( A => n4257, ZN => n4262);
   U9223 : OAI21_X1 port map( B1 => n4370, B2 => n4574, A => n4576, ZN => n4260
                           );
   U9226 : NAND2_X1 port map( A1 => n4260, A2 => n4259, ZN => n4261);
   U9227 : OAI21_X1 port map( B1 => n4263, B2 => n4262, A => n4261, ZN => n6131
                           );
   U9228 : NAND2_X1 port map( A1 => n4563, A2 => n4752, ZN => n4264);
   U9229 : MUX2_X1 port map( A => n4758, B => n4264, S => n4565, Z => n4267);
   U9230 : INV_X1 port map( A => n4756, ZN => n4566);
   U9231 : INV_X1 port map( A => n4752, ZN => n4564);
   U9232 : NAND2_X1 port map( A1 => n4566, A2 => n4564, ZN => n4265);
   U9233 : NOR2_X1 port map( A1 => n6129, A2 => n5691, ZN => n4274);
   U9234 : NOR2_X1 port map( A1 => n5025, A2 => n5022, ZN => n4270);
   U9235 : NAND2_X1 port map( A1 => n4094, A2 => n4271, ZN => n4763);
   U9236 : NOR2_X1 port map( A1 => n4763, A2 => n5024, ZN => n4272);
   U9237 : AOI22_X2 port map( A1 => n4275, A2 => n6131, B1 => n4274, B2 => 
                           n5621, ZN => n6496);
   U9238 : INV_X1 port map( A => n4276, ZN => n4279);
   U9240 : INV_X1 port map( A => n5691, ZN => n6132);
   U9241 : AOI21_X1 port map( B1 => n5623, B2 => n6132, A => n6133, ZN => n4280
                           );
   U9242 : NAND2_X1 port map( A1 => n4280, A2 => n5694, ZN => n6500);
   U9243 : NAND2_X1 port map( A1 => n6496, A2 => n6500, ZN => n6362);
   U9244 : INV_X1 port map( A => n5322, ZN => n5394);
   U9245 : NAND2_X1 port map( A1 => n5250, A2 => n5322, ZN => n4281);
   U9246 : NAND3_X1 port map( A1 => n5395, A2 => n5368, A3 => n5323, ZN => 
                           n4283);
   U9247 : OAI211_X2 port map( C1 => n5251, C2 => n5373, A => n4284, B => n4283
                           , ZN => n7211);
   U9248 : XNOR2_X1 port map( A => n6362, B => n7211, ZN => n4336);
   U9249 : NAND3_X1 port map( A1 => n20143, A2 => n4171, A3 => n4285, ZN => 
                           n4287);
   U9250 : NAND2_X1 port map( A1 => n4290, A2 => n4626, ZN => n4286);
   U9252 : NAND2_X1 port map( A1 => n4291, A2 => n4290, ZN => n4292);
   U9253 : INV_X1 port map( A => n4979, ZN => n4293);
   U9254 : NAND2_X1 port map( A1 => n4293, A2 => n4296, ZN => n4294);
   U9255 : NAND2_X1 port map( A1 => n4294, A2 => n4978, ZN => n4295);
   U9256 : NAND2_X1 port map( A1 => n4295, A2 => n4975, ZN => n4301);
   U9257 : OAI21_X1 port map( B1 => n4297, B2 => n4979, A => n4296, ZN => n4299
                           );
   U9258 : NAND2_X1 port map( A1 => n4299, A2 => n4298, ZN => n4300);
   U9259 : AND2_X1 port map( A1 => n5628, A2 => n5363, ZN => n5360);
   U9260 : NAND2_X1 port map( A1 => n4983, A2 => n19822, ZN => n4304);
   U9261 : NAND2_X1 port map( A1 => n4003, A2 => n4618, ZN => n4303);
   U9263 : OAI21_X1 port map( B1 => n4983, B2 => n4982, A => n4003, ZN => n4308
                           );
   U9264 : AND2_X1 port map( A1 => n4306, A2 => n4305, ZN => n4987);
   U9265 : INV_X1 port map( A => n4987, ZN => n4307);
   U9266 : INV_X1 port map( A => n4601, ZN => n4358);
   U9267 : AOI21_X1 port map( B1 => n4312, B2 => n4311, A => n4361, ZN => n4316
                           );
   U9268 : NAND2_X1 port map( A1 => n4152, A2 => n4548, ZN => n4362);
   U9270 : OAI21_X1 port map( B1 => n4640, B2 => n4125, A => n4317, ZN => n4322
                           );
   U9271 : NAND2_X1 port map( A1 => n4319, A2 => n4318, ZN => n4320);
   U9272 : NAND2_X1 port map( A1 => n4320, A2 => n4642, ZN => n4321);
   U9273 : NAND2_X1 port map( A1 => n4322, A2 => n4321, ZN => n4327);
   U9274 : OAI211_X1 port map( C1 => n4325, C2 => n4324, A => n4323, B => n4640
                           , ZN => n4326);
   U9275 : AND2_X2 port map( A1 => n4327, A2 => n4326, ZN => n5364);
   U9276 : INV_X1 port map( A => n5364, ZN => n5630);
   U9277 : NOR2_X1 port map( A1 => n5633, A2 => n5630, ZN => n4328);
   U9278 : INV_X1 port map( A => n5363, ZN => n5463);
   U9279 : AOI22_X1 port map( A1 => n5360, A2 => n4598, B1 => n4328, B2 => 
                           n5463, ZN => n4334);
   U9280 : AND2_X1 port map( A1 => n4013, A2 => n3717, ZN => n4331);
   U9281 : NAND2_X1 port map( A1 => n4611, A2 => n4614, ZN => n4367);
   U9282 : MUX2_X1 port map( A => n4367, B => n4365, S => n4615, Z => n4329);
   U9283 : NAND2_X1 port map( A1 => n5631, A2 => n5363, ZN => n4332);
   U9284 : OAI21_X1 port map( B1 => n5364, B2 => n5631, A => n4332, ZN => n4333
                           );
   U9285 : XNOR2_X1 port map( A => n6165, B => n2248, ZN => n4335);
   U9286 : XNOR2_X1 port map( A => n4336, B => n4335, ZN => n4466);
   U9287 : NAND2_X1 port map( A1 => n3551, A2 => n20487, ZN => n4338);
   U9288 : NAND2_X1 port map( A1 => n4518, A2 => n4339, ZN => n4341);
   U9289 : AOI21_X1 port map( B1 => n4341, B2 => n4340, A => n4524, ZN => n4346
                           );
   U9290 : NAND2_X1 port map( A1 => n4343, A2 => n4342, ZN => n4345);
   U9291 : NAND2_X1 port map( A1 => n5605, A2 => n5719, ZN => n5242);
   U9295 : NAND3_X1 port map( A1 => n4603, A2 => n4355, A3 => n4353, ZN => 
                           n4357);
   U9296 : NAND3_X1 port map( A1 => n4355, A2 => n4548, A3 => n4354, ZN => 
                           n4356);
   U9297 : AND2_X1 port map( A1 => n4357, A2 => n4356, ZN => n4360);
   U9298 : OR2_X1 port map( A1 => n4367, A2 => n4013, ZN => n4369);
   U9299 : INV_X1 port map( A => n4507, ZN => n4577);
   U9300 : NAND2_X1 port map( A1 => n4371, A2 => n4370, ZN => n4572);
   U9301 : AOI21_X1 port map( B1 => n4572, B2 => n4573, A => n4372, ZN => n4373
                           );
   U9302 : INV_X1 port map( A => n5715, ZN => n5346);
   U9303 : INV_X1 port map( A => n4962, ZN => n4893);
   U9304 : INV_X1 port map( A => n4855, ZN => n4904);
   U9305 : AOI21_X1 port map( B1 => n4493, B2 => n4904, A => n4860, ZN => n4380
                           );
   U9306 : OAI21_X1 port map( B1 => n4493, B2 => n4902, A => n4378, ZN => n4379
                           );
   U9307 : NOR2_X1 port map( A1 => n5611, A2 => n5349, ZN => n5856);
   U9308 : INV_X1 port map( A => n4864, ZN => n4381);
   U9309 : NAND2_X1 port map( A1 => n4921, A2 => n4482, ZN => n4384);
   U9312 : NAND2_X1 port map( A1 => n4385, A2 => n4968, ZN => n4386);
   U9313 : INV_X1 port map( A => n6150, ZN => n6152);
   U9314 : OAI21_X1 port map( B1 => n6151, B2 => n6155, A => n6152, ZN => n4404
                           );
   U9315 : NAND2_X1 port map( A1 => n6150, A2 => n6155, ZN => n5855);
   U9316 : INV_X1 port map( A => n4684, ZN => n4848);
   U9317 : OAI21_X1 port map( B1 => n4853, B2 => n4848, A => n4687, ZN => n4390
                           );
   U9318 : NAND2_X1 port map( A1 => n4685, A2 => n4391, ZN => n4388);
   U9319 : NAND2_X1 port map( A1 => n4388, A2 => n4387, ZN => n4389);
   U9321 : INV_X1 port map( A => n4391, ZN => n4486);
   U9323 : AND2_X1 port map( A1 => n4475, A2 => n4912, ZN => n4397);
   U9324 : INV_X1 port map( A => n4474, ZN => n4395);
   U9325 : AND2_X1 port map( A1 => n4395, A2 => n4912, ZN => n4958);
   U9326 : INV_X1 port map( A => n4958, ZN => n4396);
   U9327 : OAI21_X1 port map( B1 => n4398, B2 => n4397, A => n4396, ZN => n4401
                           );
   U9328 : NOR2_X1 port map( A1 => n4912, A2 => n4475, ZN => n4399);
   U9329 : INV_X1 port map( A => n4954, ZN => n4916);
   U9330 : INV_X1 port map( A => n6153, ZN => n6149);
   U9331 : NAND3_X1 port map( A1 => n6149, A2 => n20405, A3 => n6156, ZN => 
                           n4402);
   U9332 : AOI21_X1 port map( B1 => n5096, B2 => n5095, A => n5092, ZN => n4408
                           );
   U9333 : NAND2_X1 port map( A1 => n5098, A2 => n5092, ZN => n4786);
   U9334 : NAND2_X1 port map( A1 => n5095, A2 => n4405, ZN => n4406);
   U9335 : AOI21_X1 port map( B1 => n4786, B2 => n4406, A => n4783, ZN => n4407
                           );
   U9336 : OAI21_X1 port map( B1 => n5069, B2 => n5073, A => n2632, ZN => n4416
                           );
   U9337 : INV_X1 port map( A => n4409, ZN => n4415);
   U9338 : OAI21_X1 port map( B1 => n5069, B2 => n5071, A => n4410, ZN => n4413
                           );
   U9339 : NAND2_X1 port map( A1 => n4816, A2 => n291, ZN => n4412);
   U9340 : AND2_X1 port map( A1 => n6123, A2 => n5873, ZN => n5387);
   U9341 : NAND3_X1 port map( A1 => n19508, A2 => n1916, A3 => n169, ZN => 
                           n4419);
   U9342 : INV_X1 port map( A => n4420, ZN => n4844);
   U9343 : AND2_X1 port map( A1 => n4841, A2 => n4844, ZN => n4424);
   U9344 : NAND2_X1 port map( A1 => n4840, A2 => n164, ZN => n4423);
   U9345 : INV_X1 port map( A => n6119, ZN => n5869);
   U9346 : NAND2_X1 port map( A1 => n4824, A2 => n4669, ZN => n4826);
   U9347 : AND2_X1 port map( A1 => n4425, A2 => n4826, ZN => n5257);
   U9348 : NAND2_X1 port map( A1 => n4824, A2 => n4829, ZN => n4667);
   U9349 : NAND3_X1 port map( A1 => n6124, A2 => n5873, A3 => n6119, ZN => 
                           n4434);
   U9350 : INV_X2 port map( A => n5873, ZN => n6128);
   U9351 : NAND2_X1 port map( A1 => n20459, A2 => n20356, ZN => n4654);
   U9353 : NAND2_X1 port map( A1 => n19523, A2 => n896, ZN => n4428);
   U9354 : AOI21_X1 port map( B1 => n4654, B2 => n4428, A => n4652, ZN => n4432
                           );
   U9355 : NAND2_X1 port map( A1 => n20357, A2 => n4652, ZN => n4430);
   U9356 : AOI21_X1 port map( B1 => n4430, B2 => n3560, A => n896, ZN => n4431)
                           ;
   U9357 : OR2_X1 port map( A1 => n4432, A2 => n4431, ZN => n6118);
   U9358 : AND2_X1 port map( A1 => n4433, A2 => n4434, ZN => n4435);
   U9359 : NAND2_X1 port map( A1 => n4436, A2 => n4435, ZN => n6738);
   U9360 : INV_X1 port map( A => n5083, ZN => n4804);
   U9361 : NAND3_X1 port map( A1 => n19776, A2 => n20016, A3 => n5087, ZN => 
                           n4437);
   U9362 : INV_X1 port map( A => n4697, ZN => n5047);
   U9363 : NAND3_X1 port map( A1 => n20464, A2 => n5042, A3 => n5047, ZN => 
                           n4443);
   U9364 : INV_X1 port map( A => n6138, ZN => n5342);
   U9365 : NAND2_X1 port map( A1 => n5056, A2 => n20461, ZN => n4743);
   U9366 : INV_X1 port map( A => n4445, ZN => n4738);
   U9367 : AOI21_X1 port map( B1 => n4743, B2 => n4741, A => n4738, ZN => n4448
                           );
   U9368 : NAND2_X1 port map( A1 => n4100, A2 => n20461, ZN => n4446);
   U9369 : AOI21_X1 port map( B1 => n4446, B2 => n2929, A => n5059, ZN => n4447
                           );
   U9370 : INV_X1 port map( A => n5860, ZN => n6141);
   U9371 : NAND3_X1 port map( A1 => n4450, A2 => n3167, A3 => n5105, ZN => 
                           n4451);
   U9373 : MUX2_X1 port map( A => n303, B => n4452, S => n4771, Z => n4456);
   U9374 : NAND2_X1 port map( A1 => n303, A2 => n4708, ZN => n4454);
   U9375 : MUX2_X1 port map( A => n4454, B => n4453, S => n5035, Z => n4455);
   U9377 : OAI21_X1 port map( B1 => n5080, B2 => n5077, A => n5079, ZN => n4460
                           );
   U9378 : MUX2_X1 port map( A => n4462, B => n4461, S => n6141, Z => n4463);
   U9379 : OAI21_X2 port map( B1 => n4464, B2 => n6143, A => n4463, ZN => n7363
                           );
   U9380 : XNOR2_X1 port map( A => n7363, B => n6738, ZN => n7036);
   U9381 : XNOR2_X1 port map( A => n6881, B => n7036, ZN => n4465);
   U9383 : NOR2_X1 port map( A1 => n4941, A2 => n4940, ZN => n4469);
   U9384 : INV_X1 port map( A => n4946, ZN => n4468);
   U9385 : OAI21_X1 port map( B1 => n4889, B2 => n4469, A => n4468, ZN => n4473
                           );
   U9386 : OAI21_X1 port map( B1 => n4471, B2 => n4470, A => n4941, ZN => n4472
                           );
   U9387 : NAND2_X1 port map( A1 => n4474, A2 => n4954, ZN => n4951);
   U9388 : NAND2_X1 port map( A1 => n4954, A2 => n4475, ZN => n4476);
   U9390 : AOI21_X1 port map( B1 => n4854, B2 => n4851, A => n4848, ZN => n4489
                           );
   U9391 : AOI21_X1 port map( B1 => n4487, B2 => n4486, A => n4687, ZN => n4488
                           );
   U9392 : MUX2_X1 port map( A => n4960, B => n20205, S => n4894, Z => n4491);
   U9393 : MUX2_X1 port map( A => n4962, B => n292, S => n4892, Z => n4490);
   U9394 : OAI21_X1 port map( B1 => n4499, B2 => n4855, A => n4907, ZN => n4496
                           );
   U9395 : NAND2_X1 port map( A1 => n4494, A2 => n4493, ZN => n4495);
   U9396 : AOI21_X1 port map( B1 => n6202, B2 => n6206, A => n6204, ZN => n4502
                           );
   U9397 : MUX2_X1 port map( A => n4504, B => n4752, S => n4756, Z => n4506);
   U9398 : OAI21_X1 port map( B1 => n4566, B2 => n4565, A => n4504, ZN => n4503
                           );
   U9399 : OAI21_X1 port map( B1 => n4754, B2 => n4504, A => n4503, ZN => n4505
                           );
   U9400 : OAI21_X1 port map( B1 => n4507, B2 => n4573, A => n4511, ZN => n4508
                           );
   U9401 : NAND2_X1 port map( A1 => n4574, A2 => n4511, ZN => n4512);
   U9402 : NAND2_X1 port map( A1 => n4513, A2 => n4512, ZN => n4514);
   U9404 : NAND3_X1 port map( A1 => n4524, A2 => n4523, A3 => n4522, ZN => 
                           n4525);
   U9405 : MUX2_X1 port map( A => n5545, B => n5734, S => n5765, Z => n4552);
   U9406 : INV_X1 port map( A => n4528, ZN => n4529);
   U9408 : OAI21_X1 port map( B1 => n4529, B2 => n4532, A => n20369, ZN => 
                           n4533);
   U9409 : NAND2_X1 port map( A1 => n4636, A2 => n4533, ZN => n4534);
   U9410 : OAI21_X1 port map( B1 => n4636, B2 => n3753, A => n4534, ZN => n5539
                           );
   U9411 : NAND2_X1 port map( A1 => n4535, A2 => n4185, ZN => n5540);
   U9412 : NAND2_X1 port map( A1 => n5539, A2 => n5540, ZN => n5763);
   U9413 : OAI22_X1 port map( A1 => n4538, A2 => n4537, B1 => n4536, B2 => 
                           n4540, ZN => n5537);
   U9414 : INV_X1 port map( A => n5765, ZN => n5546);
   U9415 : NAND2_X1 port map( A1 => n4313, A2 => n4548, ZN => n4608);
   U9416 : NAND2_X1 port map( A1 => n4546, A2 => n4313, ZN => n4549);
   U9417 : AOI21_X1 port map( B1 => n4549, B2 => n4548, A => n4547, ZN => n4550
                           );
   U9418 : INV_X1 port map( A => n5768, ZN => n5735);
   U9419 : MUX2_X2 port map( A => n4552, B => n4551, S => n5735, Z => n7288);
   U9420 : NAND2_X1 port map( A1 => n4734, A2 => n20229, ZN => n4553);
   U9421 : INV_X1 port map( A => n4555, ZN => n5016);
   U9422 : OAI211_X1 port map( C1 => n5018, C2 => n20229, A => n4553, B => 
                           n5016, ZN => n4556);
   U9423 : NAND2_X1 port map( A1 => n4557, A2 => n4744, ZN => n4562);
   U9424 : MUX2_X1 port map( A => n4559, B => n4558, S => n4746, Z => n4560);
   U9425 : OAI21_X2 port map( B1 => n4562, B2 => n4561, A => n4560, ZN => n5805
                           );
   U9426 : NAND2_X1 port map( A1 => n5378, A2 => n5805, ZN => n6191);
   U9427 : OAI21_X1 port map( B1 => n4754, B2 => n4565, A => n4564, ZN => n4569
                           );
   U9428 : NAND2_X1 port map( A1 => n4566, A2 => n4752, ZN => n4568);
   U9429 : NAND2_X1 port map( A1 => n5803, A2 => n5802, ZN => n6195);
   U9430 : MUX2_X1 port map( A => n4572, B => n20190, S => n4570, Z => n4580);
   U9431 : OAI22_X1 port map( A1 => n4576, A2 => n4575, B1 => n4574, B2 => 
                           n4573, ZN => n4578);
   U9432 : NAND2_X1 port map( A1 => n4578, A2 => n4577, ZN => n4579);
   U9433 : NAND3_X1 port map( A1 => n6191, A2 => n6195, A3 => n5382, ZN => 
                           n4596);
   U9434 : AND2_X1 port map( A1 => n5805, A2 => n6189, ZN => n5379);
   U9435 : INV_X1 port map( A => n5379, ZN => n4594);
   U9436 : INV_X1 port map( A => n5805, ZN => n6193);
   U9437 : NAND3_X1 port map( A1 => n5060, A2 => n5055, A3 => n4585, ZN => 
                           n4587);
   U9438 : NAND2_X1 port map( A1 => n5057, A2 => n4738, ZN => n4586);
   U9439 : AOI22_X1 port map( A1 => n4587, A2 => n4586, B1 => n4739, B2 => 
                           n4738, ZN => n4592);
   U9440 : NAND3_X1 port map( A1 => n4588, A2 => n5055, A3 => n4738, ZN => 
                           n4589);
   U9441 : NAND2_X1 port map( A1 => n4590, A2 => n4589, ZN => n4591);
   U9442 : NOR2_X2 port map( A1 => n4592, A2 => n4591, ZN => n6192);
   U9443 : INV_X1 port map( A => n6192, ZN => n5804);
   U9445 : XNOR2_X1 port map( A => n6477, B => n19180, ZN => n4597);
   U9446 : XNOR2_X1 port map( A => n6864, B => n4597, ZN => n4729);
   U9447 : MUX2_X1 port map( A => n5631, B => n5633, S => n5364, Z => n4599);
   U9448 : MUX2_X1 port map( A => n4599, B => n5465, S => n5463, Z => n4600);
   U9449 : NAND2_X1 port map( A1 => n4602, A2 => n4601, ZN => n4604);
   U9450 : INV_X1 port map( A => n4982, ZN => n4617);
   U9451 : OAI21_X1 port map( B1 => n4988, B2 => n4618, A => n4617, ZN => n4619
                           );
   U9452 : AOI22_X1 port map( A1 => n4620, A2 => n4989, B1 => n4003, B2 => 
                           n4619, ZN => n4882);
   U9453 : NAND2_X1 port map( A1 => n4631, A2 => n4626, ZN => n4625);
   U9454 : MUX2_X1 port map( A => n4625, B => n4624, S => n4623, Z => n4629);
   U9455 : OAI211_X1 port map( C1 => n4631, C2 => n4630, A => n4629, B => n4628
                           , ZN => n5744);
   U9456 : INV_X1 port map( A => n5744, ZN => n4632);
   U9457 : NAND2_X1 port map( A1 => n3551, A2 => n19524, ZN => n4635);
   U9458 : NAND2_X1 port map( A1 => n4633, A2 => n4185, ZN => n4634);
   U9459 : NAND2_X1 port map( A1 => n4185, A2 => n19524, ZN => n4639);
   U9460 : NAND2_X1 port map( A1 => n4127, A2 => n4646, ZN => n4644);
   U9461 : NAND2_X1 port map( A1 => n4641, A2 => n4640, ZN => n4643);
   U9462 : NOR2_X1 port map( A1 => n5201, A2 => n5747, ZN => n5496);
   U9463 : INV_X1 port map( A => n6719, ZN => n4650);
   U9464 : XNOR2_X1 port map( A => n4650, B => n20203, ZN => n4727);
   U9465 : AND2_X1 port map( A1 => n4651, A2 => n896, ZN => n4653);
   U9466 : NAND2_X1 port map( A1 => n4659, A2 => n4658, ZN => n4660);
   U9467 : AOI21_X1 port map( B1 => n4662, B2 => n2632, A => n4410, ZN => n4666
                           );
   U9468 : NAND2_X1 port map( A1 => n4664, A2 => n4663, ZN => n5070);
   U9469 : INV_X1 port map( A => n6171, ZN => n4691);
   U9470 : MUX2_X1 port map( A => n4675, B => n4835, S => n19508, Z => n4680);
   U9471 : NAND2_X1 port map( A1 => n5115, A2 => n4675, ZN => n4678);
   U9472 : NAND2_X1 port map( A1 => n2042, A2 => n169, ZN => n4677);
   U9473 : MUX2_X1 port map( A => n4678, B => n4677, S => n4676, Z => n4679);
   U9474 : NAND2_X1 port map( A1 => n1867, A2 => n6166, ZN => n4689);
   U9475 : OAI21_X1 port map( B1 => n4682, B2 => n4684, A => n4681, ZN => n4683
                           );
   U9476 : NAND2_X1 port map( A1 => n4683, A2 => n4391, ZN => n5219);
   U9477 : NAND2_X1 port map( A1 => n4684, A2 => n177, ZN => n5217);
   U9478 : AND2_X1 port map( A1 => n178, A2 => n4685, ZN => n4850);
   U9479 : OAI21_X1 port map( B1 => n3996, B2 => n4687, A => n4850, ZN => n5218
                           );
   U9480 : OAI21_X2 port map( B1 => n4692, B2 => n4691, A => n4690, ZN => n7216
                           );
   U9481 : MUX2_X1 port map( A => n5101, B => n4693, S => n5102, Z => n4695);
   U9482 : NAND2_X1 port map( A1 => n4693, A2 => n5100, ZN => n4790);
   U9483 : AND2_X1 port map( A1 => n4790, A2 => n4792, ZN => n4694);
   U9484 : NOR2_X1 port map( A1 => n6183, A2 => n5847, ZN => n6182);
   U9485 : AND2_X1 port map( A1 => n4699, A2 => n4700, ZN => n4704);
   U9486 : NAND2_X1 port map( A1 => n4804, A2 => n19777, ZN => n5091);
   U9487 : NAND2_X1 port map( A1 => n4801, A2 => n5086, ZN => n4702);
   U9488 : MUX2_X1 port map( A => n5091, B => n4702, S => n5088, Z => n4703);
   U9489 : NOR2_X1 port map( A1 => n5846, A2 => n5730, ZN => n4705);
   U9490 : NOR2_X1 port map( A1 => n6182, A2 => n4705, ZN => n6382);
   U9491 : INV_X1 port map( A => n6382, ZN => n4725);
   U9492 : AOI22_X1 port map( A1 => n303, A2 => n4707, B1 => n4706, B2 => n4708
                           , ZN => n4711);
   U9493 : MUX2_X1 port map( A => n4709, B => n4708, S => n4707, Z => n4710);
   U9494 : OAI211_X1 port map( C1 => n5093, C2 => n4713, A => n4712, B => n4783
                           , ZN => n4718);
   U9495 : NAND2_X1 port map( A1 => n4714, A2 => n5094, ZN => n4717);
   U9496 : NOR2_X1 port map( A1 => n4788, A2 => n4715, ZN => n4716);
   U9498 : AND2_X1 port map( A1 => n5080, A2 => n5077, ZN => n4722);
   U9499 : NAND2_X1 port map( A1 => n5081, A2 => n4719, ZN => n5076);
   U9500 : NAND2_X1 port map( A1 => n4720, A2 => n5078, ZN => n4721);
   U9501 : INV_X1 port map( A => n5383, ZN => n4723);
   U9502 : OAI211_X1 port map( C1 => n19476, C2 => n6379, A => n4723, B => 
                           n6184, ZN => n4724);
   U9503 : OAI21_X1 port map( B1 => n4725, B2 => n6184, A => n4724, ZN => n4726
                           );
   U9504 : XNOR2_X1 port map( A => n7216, B => n4726, ZN => n6562);
   U9505 : XNOR2_X1 port map( A => n4727, B => n6562, ZN => n4728);
   U9507 : MUX2_X1 port map( A => n7461, B => n4730, S => n8190, Z => n5137);
   U9508 : OAI21_X1 port map( B1 => n5012, B2 => n5014, A => n4731, ZN => n4733
                           );
   U9509 : NAND2_X1 port map( A1 => n5058, A2 => n4738, ZN => n4740);
   U9510 : NAND3_X1 port map( A1 => n4740, A2 => n4739, A3 => n5057, ZN => 
                           n4742);
   U9511 : INV_X1 port map( A => n6104, ZN => n5659);
   U9512 : INV_X1 port map( A => n4745, ZN => n5004);
   U9513 : NAND2_X1 port map( A1 => n4750, A2 => n5010, ZN => n4747);
   U9514 : MUX2_X1 port map( A => n4748, B => n4747, S => n5006, Z => n4749);
   U9515 : AOI21_X1 port map( B1 => n4753, B2 => n4754, A => n4752, ZN => n4760
                           );
   U9516 : NAND2_X1 port map( A1 => n4755, A2 => n4754, ZN => n4757);
   U9517 : AOI21_X1 port map( B1 => n4758, B2 => n4757, A => n4756, ZN => n4759
                           );
   U9518 : NOR2_X1 port map( A1 => n5172, A2 => n6109, ZN => n4776);
   U9519 : NAND2_X1 port map( A1 => n4761, A2 => n19788, ZN => n4762);
   U9520 : NAND2_X1 port map( A1 => n4763, A2 => n4762, ZN => n4768);
   U9521 : NAND2_X1 port map( A1 => n4765, A2 => n5022, ZN => n4766);
   U9522 : NAND2_X1 port map( A1 => n5027, A2 => n4766, ZN => n4767);
   U9523 : MUX2_X2 port map( A => n4768, B => n4767, S => n5026, Z => n6105);
   U9524 : OAI22_X1 port map( A1 => n153, A2 => n5035, B1 => n303, B2 => n4769,
                           ZN => n4770);
   U9525 : NAND3_X1 port map( A1 => n5038, A2 => n303, A3 => n4772, ZN => n4773
                           );
   U9526 : INV_X1 port map( A => n6107, ZN => n5656);
   U9527 : NAND3_X1 port map( A1 => n5657, A2 => n6104, A3 => n5656, ZN => 
                           n4775);
   U9528 : XNOR2_X1 port map( A => n7384, B => n2122, ZN => n4781);
   U9529 : NOR2_X1 port map( A1 => n5649, A2 => n5643, ZN => n4779);
   U9531 : NAND2_X1 port map( A1 => n4777, A2 => n5648, ZN => n4778);
   U9532 : INV_X1 port map( A => n7336, ZN => n4780);
   U9533 : INV_X1 port map( A => n4782, ZN => n4785);
   U9534 : NAND2_X1 port map( A1 => n2460, A2 => n4783, ZN => n4784);
   U9535 : NAND2_X1 port map( A1 => n4785, A2 => n4784, ZN => n4787);
   U9536 : OAI211_X1 port map( C1 => n4789, C2 => n4788, A => n4787, B => n4786
                           , ZN => n5952);
   U9537 : NAND2_X1 port map( A1 => n5101, A2 => n5107, ZN => n4791);
   U9538 : MUX2_X1 port map( A => n4791, B => n4790, S => n5102, Z => n4794);
   U9539 : INV_X1 port map( A => n4795, ZN => n4797);
   U9540 : NAND2_X1 port map( A1 => n4799, A2 => n4798, ZN => n4800);
   U9541 : NAND2_X1 port map( A1 => n4801, A2 => n20016, ZN => n4808);
   U9542 : NAND2_X1 port map( A1 => n4802, A2 => n20202, ZN => n4803);
   U9543 : NAND3_X1 port map( A1 => n4808, A2 => n5090, A3 => n4803, ZN => 
                           n4806);
   U9544 : OAI211_X1 port map( C1 => n4808, C2 => n4807, A => n4806, B => n4805
                           , ZN => n5949);
   U9545 : NOR2_X1 port map( A1 => n6101, A2 => n5949, ZN => n4822);
   U9546 : NAND2_X1 port map( A1 => n20431, A2 => n5075, ZN => n4811);
   U9547 : OAI21_X1 port map( B1 => n5075, B2 => n5077, A => n4811, ZN => n4812
                           );
   U9548 : INV_X1 port map( A => n6097, ZN => n5662);
   U9549 : INV_X1 port map( A => n4814, ZN => n4815);
   U9550 : NAND2_X1 port map( A1 => n4815, A2 => n5069, ZN => n4820);
   U9551 : OAI21_X1 port map( B1 => n2971, B2 => n291, A => n5073, ZN => n4817)
                           ;
   U9552 : NAND2_X1 port map( A1 => n4818, A2 => n4817, ZN => n4819);
   U9553 : NAND2_X1 port map( A1 => n5950, A2 => n5664, ZN => n4821);
   U9554 : INV_X1 port map( A => n4823, ZN => n4833);
   U9555 : NAND2_X1 port map( A1 => n4828, A2 => n4827, ZN => n4830);
   U9556 : MUX2_X1 port map( A => n4831, B => n4830, S => n4829, Z => n4832);
   U9557 : OAI21_X1 port map( B1 => n19688, B2 => n4833, A => n4832, ZN => 
                           n5200);
   U9558 : AOI21_X1 port map( B1 => n20256, B2 => n4834, A => n169, ZN => n4836
                           );
   U9559 : OR2_X1 port map( A1 => n4836, A2 => n4835, ZN => n4837);
   U9560 : INV_X1 port map( A => n6092, ZN => n5912);
   U9561 : INV_X1 port map( A => n4839, ZN => n4843);
   U9562 : NOR2_X1 port map( A1 => n4841, A2 => n4840, ZN => n4842);
   U9563 : NOR2_X1 port map( A1 => n4846, A2 => n4845, ZN => n5902);
   U9564 : INV_X1 port map( A => n5902, ZN => n4847);
   U9566 : INV_X1 port map( A => n6090, ZN => n5493);
   U9567 : NAND2_X1 port map( A1 => n4850, A2 => n4849, ZN => n4852);
   U9568 : OAI211_X1 port map( C1 => n4854, C2 => n4853, A => n4852, B => n4851
                           , ZN => n6087);
   U9569 : INV_X1 port map( A => n6087, ZN => n5176);
   U9570 : NAND2_X1 port map( A1 => n5493, A2 => n5176, ZN => n4876);
   U9572 : INV_X1 port map( A => n4856, ZN => n4903);
   U9573 : NAND2_X1 port map( A1 => n4903, A2 => n4901, ZN => n4858);
   U9574 : NAND2_X1 port map( A1 => n4858, A2 => n4857, ZN => n4859);
   U9575 : INV_X1 port map( A => n5901, ZN => n4862);
   U9576 : NAND3_X1 port map( A1 => n20357, A2 => n4867, A3 => n896, ZN => 
                           n4869);
   U9577 : NAND3_X1 port map( A1 => n4871, A2 => n4870, A3 => n4869, ZN => 
                           n4872);
   U9578 : NAND2_X1 port map( A1 => n890, A2 => n5899, ZN => n4874);
   U9579 : XNOR2_X1 port map( A => n7184, B => n6918, ZN => n7040);
   U9580 : INV_X1 port map( A => n5670, ZN => n5185);
   U9581 : NAND2_X1 port map( A1 => n5185, A2 => n5425, ZN => n4880);
   U9582 : NAND2_X1 port map( A1 => n5675, A2 => n5668, ZN => n5677);
   U9583 : INV_X1 port map( A => n5669, ZN => n5676);
   U9584 : OAI21_X1 port map( B1 => n3397, B2 => n5670, A => n5676, ZN => n4878
                           );
   U9585 : OAI21_X1 port map( B1 => n5279, B2 => n5668, A => n5669, ZN => n4877
                           );
   U9586 : NAND2_X1 port map( A1 => n4878, A2 => n4877, ZN => n4879);
   U9587 : NOR2_X1 port map( A1 => n20509, A2 => n5745, ZN => n5497);
   U9588 : NAND2_X1 port map( A1 => n5201, A2 => n5741, ZN => n4881);
   U9589 : NAND2_X1 port map( A1 => n5497, A2 => n4881, ZN => n4884);
   U9590 : INV_X1 port map( A => n4882, ZN => n5749);
   U9591 : NAND3_X1 port map( A1 => n5741, A2 => n5743, A3 => n5745, ZN => 
                           n4883);
   U9592 : XNOR2_X1 port map( A => n7188, B => n7337, ZN => n4938);
   U9593 : INV_X1 port map( A => n4885, ZN => n4891);
   U9594 : OAI21_X1 port map( B1 => n4946, B2 => n4887, A => n4886, ZN => n4890
                           );
   U9596 : OAI21_X1 port map( B1 => n4892, B2 => n4893, A => n4899, ZN => n4897
                           );
   U9598 : AOI21_X1 port map( B1 => n4903, B2 => n4902, A => n4901, ZN => n4908
                           );
   U9599 : NAND2_X1 port map( A1 => n4905, A2 => n4904, ZN => n4906);
   U9600 : NAND2_X1 port map( A1 => n4912, A2 => n4911, ZN => n4955);
   U9602 : NAND3_X1 port map( A1 => n4955, A2 => n4916, A3 => n4915, ZN => 
                           n4917);
   U9603 : NAND2_X1 port map( A1 => n5684, A2 => n5476, ZN => n5680);
   U9604 : NAND2_X1 port map( A1 => n4968, A2 => n19507, ZN => n4920);
   U9605 : OAI211_X1 port map( C1 => n4921, C2 => n19507, A => n4920, B => 
                           n4919, ZN => n4923);
   U9606 : OAI21_X1 port map( B1 => n3967, B2 => n4965, A => n4482, ZN => n4922
                           );
   U9607 : NAND2_X1 port map( A1 => n4923, A2 => n4922, ZN => n4924);
   U9608 : OAI21_X1 port map( B1 => n4926, B2 => n19507, A => n4924, ZN => 
                           n6083);
   U9609 : INV_X1 port map( A => n6083, ZN => n5411);
   U9610 : AOI22_X1 port map( A1 => n5686, A2 => n5680, B1 => n5411, B2 => 
                           n3529, ZN => n4936);
   U9611 : NAND2_X1 port map( A1 => n4928, A2 => n4974, ZN => n4929);
   U9612 : AOI22_X1 port map( A1 => n4931, A2 => n4930, B1 => n4929, B2 => 
                           n4976, ZN => n4934);
   U9613 : NOR2_X1 port map( A1 => n4932, A2 => n4974, ZN => n4933);
   U9614 : OR2_X1 port map( A1 => n5683, A2 => n5410, ZN => n5412);
   U9615 : NOR2_X1 port map( A1 => n5412, A2 => n5684, ZN => n4935);
   U9616 : OR2_X1 port map( A1 => n4936, A2 => n4935, ZN => n7383);
   U9617 : INV_X1 port map( A => n7383, ZN => n4937);
   U9618 : XNOR2_X1 port map( A => n4938, B => n4937, ZN => n6877);
   U9619 : XNOR2_X1 port map( A => n4939, B => n6877, ZN => n8185);
   U9620 : INV_X1 port map( A => n8062, ZN => n7606);
   U9623 : NAND2_X1 port map( A1 => n4945, A2 => n4118, ZN => n4944);
   U9624 : OAI21_X1 port map( B1 => n4946, B2 => n4945, A => n4944, ZN => n4948
                           );
   U9625 : NAND2_X1 port map( A1 => n4951, A2 => n4950, ZN => n4959);
   U9626 : NAND2_X1 port map( A1 => n292, A2 => n20205, ZN => n4964);
   U9627 : NAND2_X1 port map( A1 => n4962, A2 => n4892, ZN => n4963);
   U9628 : AOI21_X1 port map( B1 => n4967, B2 => n4966, A => n4965, ZN => n4973
                           );
   U9629 : AOI21_X1 port map( B1 => n4971, B2 => n4970, A => n4482, ZN => n4972
                           );
   U9630 : INV_X1 port map( A => n6036, ZN => n5564);
   U9631 : INV_X1 port map( A => n5531, ZN => n4981);
   U9632 : INV_X1 port map( A => n4974, ZN => n4975);
   U9633 : NAND3_X1 port map( A1 => n6033, A2 => n4981, A3 => n20241, ZN => 
                           n4992);
   U9634 : NAND2_X1 port map( A1 => n4983, A2 => n4982, ZN => n4984);
   U9635 : NAND2_X1 port map( A1 => n4985, A2 => n4984, ZN => n4986);
   U9636 : NAND2_X1 port map( A1 => n4989, A2 => n4988, ZN => n4990);
   U9637 : AND2_X1 port map( A1 => n4992, A2 => n5471, ZN => n4993);
   U9638 : NAND2_X1 port map( A1 => n5328, A2 => n6048, ZN => n4999);
   U9639 : NOR2_X1 port map( A1 => n5559, A2 => n6050, ZN => n4994);
   U9640 : NAND2_X1 port map( A1 => n3351, A2 => n4994, ZN => n4998);
   U9642 : NAND3_X1 port map( A1 => n5139, A2 => n5138, A3 => n6049, ZN => 
                           n4996);
   U9644 : XNOR2_X1 port map( A => n7318, B => n7371, ZN => n6889);
   U9645 : AOI21_X1 port map( B1 => n5405, B2 => n3959, A => n5148, ZN => n5002
                           );
   U9646 : NOR2_X1 port map( A1 => n5408, A2 => n5580, ZN => n5318);
   U9647 : OAI21_X1 port map( B1 => n5318, B2 => n5000, A => n946, ZN => n5001)
                           ;
   U9648 : AOI22_X1 port map( A1 => n5007, A2 => n5004, B1 => n5003, B2 => 
                           n5006, ZN => n5011);
   U9649 : NAND2_X1 port map( A1 => n4248, A2 => n5004, ZN => n5008);
   U9651 : NAND3_X1 port map( A1 => n5015, A2 => n5014, A3 => n5013, ZN => 
                           n5020);
   U9652 : NAND3_X1 port map( A1 => n5018, A2 => n20229, A3 => n5016, ZN => 
                           n5019);
   U9653 : NAND2_X1 port map( A1 => n5030, A2 => n5927, ZN => n5066);
   U9654 : INV_X1 port map( A => n6027, ZN => n5192);
   U9655 : NAND2_X1 port map( A1 => n5032, A2 => n153, ZN => n5033);
   U9656 : NAND2_X1 port map( A1 => n5034, A2 => n5033, ZN => n5039);
   U9657 : INV_X1 port map( A => n6025, ZN => n5520);
   U9658 : NAND3_X1 port map( A1 => n6026, A2 => n5192, A3 => n5520, ZN => 
                           n5065);
   U9659 : NAND2_X1 port map( A1 => n5040, A2 => n5045, ZN => n5041);
   U9660 : OAI211_X1 port map( C1 => n5044, C2 => n5043, A => n5042, B => n5041
                           , ZN => n5051);
   U9661 : AND2_X1 port map( A1 => n5046, A2 => n5045, ZN => n5049);
   U9662 : OAI211_X1 port map( C1 => n5049, C2 => n20464, A => n5048, B => 
                           n5047, ZN => n5050);
   U9663 : NAND2_X1 port map( A1 => n5927, A2 => n5926, ZN => n5064);
   U9664 : NAND3_X1 port map( A1 => n5057, A2 => n5056, A3 => n5055, ZN => 
                           n5062);
   U9665 : NAND3_X1 port map( A1 => n5060, A2 => n5059, A3 => n5058, ZN => 
                           n5061);
   U9666 : NAND3_X1 port map( A1 => n5192, A2 => n19789, A3 => n5930, ZN => 
                           n5063);
   U9667 : INV_X1 port map( A => n7373, ZN => n5067);
   U9668 : XNOR2_X1 port map( A => n7088, B => n5067, ZN => n5068);
   U9669 : XNOR2_X1 port map( A => n5068, B => n6889, ZN => n5134);
   U9670 : OR2_X1 port map( A1 => n5070, A2 => n5069, ZN => n5504);
   U9671 : AND3_X1 port map( A1 => n5080, A2 => n3451, A3 => n5079, ZN => n5508
                           );
   U9673 : OAI21_X1 port map( B1 => n5083, B2 => n5086, A => n20016, ZN => 
                           n5085);
   U9674 : OR3_X1 port map( A1 => n5088, A2 => n5087, A3 => n5086, ZN => n5089)
                           ;
   U9675 : INV_X1 port map( A => n19979, ZN => n5921);
   U9676 : OAI22_X1 port map( A1 => n6007, A2 => n5914, B1 => n5921, B2 => n861
                           , ZN => n5111);
   U9678 : MUX2_X1 port map( A => n5107, B => n5106, S => n4048, Z => n5109);
   U9679 : NAND2_X1 port map( A1 => n5109, A2 => n5108, ZN => n5110);
   U9680 : NAND2_X1 port map( A1 => n5111, A2 => n5590, ZN => n5123);
   U9681 : NAND2_X1 port map( A1 => n20256, A2 => n19508, ZN => n5113);
   U9682 : AOI21_X1 port map( B1 => n5114, B2 => n5113, A => n5115, ZN => n5121
                           );
   U9683 : NAND2_X1 port map( A1 => n5116, A2 => n5115, ZN => n5119);
   U9684 : AOI21_X1 port map( B1 => n5119, B2 => n169, A => n19508, ZN => n5120
                           );
   U9685 : INV_X1 port map( A => n5823, ZN => n5828);
   U9686 : NAND3_X1 port map( A1 => n5828, A2 => n5447, A3 => n3569, ZN => 
                           n5127);
   U9687 : NAND2_X1 port map( A1 => n5124, A2 => n5823, ZN => n5126);
   U9688 : NAND3_X1 port map( A1 => n5447, A2 => n5825, A3 => n6016, ZN => 
                           n5125);
   U9689 : XNOR2_X1 port map( A => n7046, B => n7179, ZN => n6579);
   U9690 : NAND2_X1 port map( A1 => n5647, A2 => n5641, ZN => n5128);
   U9691 : AOI21_X1 port map( B1 => n5128, B2 => n5648, A => n5649, ZN => n5131
                           );
   U9692 : NAND2_X1 port map( A1 => n5442, A2 => n5444, ZN => n5291);
   U9693 : NAND3_X1 port map( A1 => n5649, A2 => n5444, A3 => n5643, ZN => 
                           n5129);
   U9694 : NAND2_X1 port map( A1 => n5291, A2 => n5129, ZN => n5130);
   U9695 : XNOR2_X1 port map( A => n7144, B => n1840, ZN => n5132);
   U9696 : XNOR2_X1 port map( A => n6579, B => n5132, ZN => n5133);
   U9697 : AOI21_X1 port map( B1 => n20465, B2 => n8184, A => n8060, ZN => 
                           n5135);
   U9698 : AND2_X1 port map( A1 => n8182, A2 => n5135, ZN => n5136);
   U9699 : INV_X1 port map( A => n5559, ZN => n6051);
   U9702 : AND2_X1 port map( A1 => n5559, A2 => n6049, ZN => n5329);
   U9703 : NOR3_X1 port map( A1 => n5329, A2 => n3351, A3 => n5330, ZN => n5142
                           );
   U9704 : NAND2_X1 port map( A1 => n6044, A2 => n5888, ZN => n5781);
   U9705 : INV_X1 port map( A => n6041, ZN => n5776);
   U9706 : NAND3_X1 port map( A1 => n135, A2 => n5776, A3 => n5309, ZN => n5145
                           );
   U9707 : XNOR2_X1 port map( A => n6674, B => n6494, ZN => n7228);
   U9708 : NAND3_X1 port map( A1 => n5571, A2 => n5580, A3 => n5582, ZN => 
                           n5151);
   U9709 : NAND2_X1 port map( A1 => n5408, A2 => n3959, ZN => n5317);
   U9710 : NAND3_X2 port map( A1 => n5152, A2 => n5151, A3 => n5150, ZN => 
                           n7212);
   U9711 : OAI21_X1 port map( B1 => n6068, B2 => n5978, A => n6069, ZN => n5155
                           );
   U9712 : INV_X1 port map( A => n5978, ZN => n6075);
   U9713 : NOR2_X1 port map( A1 => n6067, A2 => n6072, ZN => n5880);
   U9714 : XNOR2_X1 port map( A => n7212, B => n7232, ZN => n6801);
   U9715 : XNOR2_X1 port map( A => n6801, B => n7228, ZN => n5166);
   U9716 : INV_X1 port map( A => n5796, ZN => n5792);
   U9717 : XNOR2_X1 port map( A => n7364, B => n7211, ZN => n5164);
   U9718 : INV_X1 port map( A => n6057, ZN => n6056);
   U9719 : NAND3_X1 port map( A1 => n6064, A2 => n6056, A3 => n5891, ZN => 
                           n5162);
   U9720 : NAND3_X1 port map( A1 => n6064, A2 => n6057, A3 => n6055, ZN => 
                           n5161);
   U9721 : INV_X1 port map( A => n5782, ZN => n5895);
   U9722 : NAND3_X1 port map( A1 => n6058, A2 => n20670, A3 => n5895, ZN => 
                           n5160);
   U9723 : NAND3_X1 port map( A1 => n906, A2 => n5891, A3 => n6059, ZN => n5159
                           );
   U9724 : XNOR2_X1 port map( A => n7365, B => n2096, ZN => n5163);
   U9725 : XNOR2_X1 port map( A => n5164, B => n5163, ZN => n5165);
   U9726 : NAND2_X1 port map( A1 => n5663, A2 => n5953, ZN => n5167);
   U9727 : NAND2_X1 port map( A1 => n5661, A2 => n5167, ZN => n5171);
   U9728 : OAI21_X1 port map( B1 => n6097, B2 => n5949, A => n6101, ZN => n5170
                           );
   U9729 : INV_X1 port map( A => n5949, ZN => n5168);
   U9730 : NOR2_X1 port map( A1 => n5663, A2 => n5168, ZN => n5169);
   U9731 : AOI21_X2 port map( B1 => n5171, B2 => n5170, A => n5169, ZN => n6679
                           );
   U9732 : INV_X1 port map( A => n6105, ZN => n5955);
   U9733 : NAND3_X1 port map( A1 => n5955, A2 => n5957, A3 => n6109, ZN => 
                           n5175);
   U9734 : NAND3_X1 port map( A1 => n5172, A2 => n6108, A3 => n6109, ZN => 
                           n5174);
   U9735 : NAND3_X1 port map( A1 => n6113, A2 => n5957, A3 => n6104, ZN => 
                           n5173);
   U9736 : XNOR2_X1 port map( A => n6679, B => n6634, ZN => n7279);
   U9737 : INV_X1 port map( A => n7279, ZN => n6926);
   U9738 : OAI21_X1 port map( B1 => n5199, B2 => n890, A => n20149, ZN => n5177
                           );
   U9739 : INV_X1 port map( A => n5200, ZN => n5494);
   U9740 : NAND3_X1 port map( A1 => n5742, A2 => n5201, A3 => n5749, ZN => 
                           n5178);
   U9741 : XNOR2_X1 port map( A => n6926, B => n7377, ZN => n5191);
   U9742 : INV_X1 port map( A => n5682, ZN => n6084);
   U9743 : INV_X1 port map( A => n5476, ZN => n6082);
   U9744 : OAI21_X1 port map( B1 => n6082, B2 => n6083, A => n5684, ZN => n5182
                           );
   U9745 : AND2_X1 port map( A1 => n5682, A2 => n6083, ZN => n5181);
   U9746 : INV_X1 port map( A => n5425, ZN => n5184);
   U9747 : NAND2_X1 port map( A1 => n5668, A2 => n5184, ZN => n5188);
   U9748 : NAND3_X1 port map( A1 => n5669, A2 => n5185, A3 => n5184, ZN => 
                           n5186);
   U9749 : XNOR2_X1 port map( A => n7144, B => n19205, ZN => n5189);
   U9750 : XNOR2_X1 port map( A => n6838, B => n5189, ZN => n5190);
   U9751 : INV_X1 port map( A => n5926, ZN => n5931);
   U9752 : OR2_X1 port map( A1 => n5931, A2 => n6025, ZN => n6030);
   U9753 : AOI21_X1 port map( B1 => n6028, B2 => n6030, A => n5192, ZN => n5195
                           );
   U9755 : AOI21_X1 port map( B1 => n5193, B2 => n5926, A => n5929, ZN => n5194
                           );
   U9756 : NAND2_X1 port map( A1 => n5736, A2 => n5768, ZN => n5224);
   U9758 : INV_X1 port map( A => n5763, ZN => n5769);
   U9759 : AOI21_X1 port map( B1 => n5224, B2 => n5225, A => n5769, ZN => n5198
                           );
   U9760 : NAND2_X1 port map( A1 => n5765, A2 => n5767, ZN => n5196);
   U9761 : AOI21_X1 port map( B1 => n5766, B2 => n5196, A => n5736, ZN => n5197
                           );
   U9762 : NAND2_X1 port map( A1 => n5203, A2 => n5202, ZN => n5204);
   U9763 : NAND2_X1 port map( A1 => n5204, A2 => n5745, ZN => n5206);
   U9764 : NAND2_X1 port map( A1 => n5742, A2 => n5746, ZN => n5205);
   U9766 : XNOR2_X1 port map( A => n7238, B => n6824, ZN => n5214);
   U9767 : INV_X1 port map( A => n6007, ZN => n5207);
   U9768 : INV_X1 port map( A => n5917, ZN => n6013);
   U9769 : AOI21_X1 port map( B1 => n5916, B2 => n5207, A => n6013, ZN => n5210
                           );
   U9770 : NAND2_X1 port map( A1 => n5208, A2 => n6010, ZN => n5209);
   U9771 : XNOR2_X1 port map( A => n7392, B => n6854, ZN => n5212);
   U9772 : INV_X1 port map( A => n20672, ZN => n18660);
   U9773 : XNOR2_X1 port map( A => n7196, B => n18660, ZN => n5211);
   U9774 : XNOR2_X1 port map( A => n5212, B => n5211, ZN => n5213);
   U9775 : NOR2_X1 port map( A1 => n8304, A2 => n8301, ZN => n5272);
   U9777 : AOI21_X1 port map( B1 => n5631, B2 => n5633, A => n5363, ZN => n5216
                           );
   U9778 : INV_X1 port map( A => n6808, ZN => n5222);
   U9779 : INV_X1 port map( A => n6167, ZN => n6176);
   U9780 : AND2_X1 port map( A1 => n5218, A2 => n5217, ZN => n5220);
   U9782 : NAND2_X1 port map( A1 => n6176, A2 => n5945, ZN => n5943);
   U9783 : NAND2_X1 port map( A1 => n6172, A2 => n6168, ZN => n6175);
   U9784 : INV_X1 port map( A => n6171, ZN => n5842);
   U9785 : OAI211_X1 port map( C1 => n6166, C2 => n6172, A => n170, B => n5842,
                           ZN => n5221);
   U9786 : XNOR2_X1 port map( A => n5222, B => n6873, ZN => n7381);
   U9787 : INV_X1 port map( A => n7381, ZN => n6464);
   U9788 : OAI211_X1 port map( C1 => n5763, C2 => n5768, A => n5546, B => n5734
                           , ZN => n5223);
   U9790 : INV_X1 port map( A => n5839, ZN => n6203);
   U9792 : NOR2_X1 port map( A1 => n6204, A2 => n19968, ZN => n5230);
   U9793 : NAND3_X1 port map( A1 => n6218, A2 => n6205, A3 => n19492, ZN => 
                           n5227);
   U9794 : OAI21_X1 port map( B1 => n5226, B2 => n6218, A => n5227, ZN => n5228
                           );
   U9795 : INV_X1 port map( A => n5228, ZN => n5229);
   U9796 : XNOR2_X1 port map( A => n7187, B => n7249, ZN => n6810);
   U9797 : XNOR2_X1 port map( A => n6810, B => n6464, ZN => n5239);
   U9798 : NAND2_X1 port map( A1 => n5382, A2 => n6189, ZN => n5234);
   U9799 : INV_X1 port map( A => n6190, ZN => n5232);
   U9800 : NOR2_X1 port map( A1 => n5805, A2 => n6189, ZN => n5231);
   U9801 : OAI22_X1 port map( A1 => n5232, A2 => n5231, B1 => n6194, B2 => 
                           n5803, ZN => n5233);
   U9802 : INV_X1 port map( A => n6919, ZN => n6513);
   U9803 : NOR2_X1 port map( A1 => n6184, A2 => n5845, ZN => n5235);
   U9804 : INV_X1 port map( A => n5728, ZN => n6380);
   U9805 : XNOR2_X1 port map( A => n6513, B => n7248, ZN => n5237);
   U9806 : XNOR2_X1 port map( A => n7188, B => n2221, ZN => n5236);
   U9807 : XNOR2_X1 port map( A => n5237, B => n5236, ZN => n5238);
   U9808 : NOR2_X1 port map( A1 => n8046, A2 => n8044, ZN => n5271);
   U9809 : INV_X1 port map( A => n5240, ZN => n5241);
   U9810 : OAI211_X1 port map( C1 => n5346, C2 => n5605, A => n5243, B => n5720
                           , ZN => n5244);
   U9811 : NAND2_X1 port map( A1 => n6150, A2 => n5612, ZN => n5246);
   U9813 : XNOR2_X1 port map( A => n7254, B => n5249, ZN => n6590);
   U9814 : INV_X1 port map( A => n6590, ZN => n6818);
   U9815 : NAND2_X1 port map( A1 => n5401, A2 => n5251, ZN => n5252);
   U9816 : INV_X1 port map( A => n6123, ZN => n5338);
   U9817 : NAND2_X1 port map( A1 => n6128, A2 => n5338, ZN => n5870);
   U9818 : OAI21_X1 port map( B1 => n6128, B2 => n6119, A => n5386, ZN => n5260
                           );
   U9819 : NAND2_X1 port map( A1 => n5255, A2 => n19688, ZN => n5256);
   U9820 : OAI211_X1 port map( C1 => n19688, C2 => n5257, A => n6128, B => 
                           n5256, ZN => n5259);
   U9821 : OAI211_X1 port map( C1 => n6117, C2 => n6128, A => n5260, B => n5259
                           , ZN => n5261);
   U9822 : XNOR2_X1 port map( A => n6818, B => n7353, ZN => n5270);
   U9823 : XNOR2_X1 port map( A => n20203, B => n2296, ZN => n5268);
   U9824 : MUX2_X1 port map( A => n6129, B => n6131, S => n6133, Z => n5263);
   U9826 : NAND2_X1 port map( A1 => n6139, A2 => n6138, ZN => n5265);
   U9827 : MUX2_X1 port map( A => n5267, B => n5266, S => n5860, Z => n6285);
   U9828 : XNOR2_X1 port map( A => n6285, B => n6520, ZN => n7256);
   U9829 : XNOR2_X1 port map( A => n7256, B => n5268, ZN => n5269);
   U9830 : AND2_X1 port map( A1 => n5704, A2 => n5997, ZN => n5433);
   U9831 : NAND2_X1 port map( A1 => n5433, A2 => n5434, ZN => n5274);
   U9832 : NAND3_X1 port map( A1 => n19562, A2 => n5996, A3 => n6002, ZN => 
                           n5273);
   U9833 : XNOR2_X1 port map( A => n6850, B => n19222, ZN => n5278);
   U9834 : NAND2_X1 port map( A1 => n5711, A2 => n5985, ZN => n5993);
   U9835 : INV_X1 port map( A => n5711, ZN => n5817);
   U9836 : NAND2_X1 port map( A1 => n5818, A2 => n5989, ZN => n5277);
   U9837 : XNOR2_X1 port map( A => n5278, B => n6947, ZN => n5284);
   U9838 : NAND2_X1 port map( A1 => n3397, A2 => n5425, ZN => n5282);
   U9839 : NOR2_X1 port map( A1 => n5670, A2 => n5279, ZN => n5280);
   U9840 : XNOR2_X1 port map( A => n7202, B => n6945, ZN => n5283);
   U9841 : XNOR2_X1 port map( A => n5284, B => n5283, ZN => n5297);
   U9842 : NOR2_X1 port map( A1 => n3569, A2 => n6017, ZN => n5286);
   U9843 : NOR2_X1 port map( A1 => n5823, A2 => n5827, ZN => n5285);
   U9844 : OAI21_X1 port map( B1 => n5286, B2 => n5285, A => n5825, ZN => n5288
                           );
   U9845 : NAND3_X1 port map( A1 => n5824, A2 => n5826, A3 => n6022, ZN => 
                           n5287);
   U9846 : INV_X1 port map( A => n5442, ZN => n5646);
   U9847 : NAND2_X1 port map( A1 => n5646, A2 => n5641, ZN => n5289);
   U9848 : INV_X1 port map( A => n5443, ZN => n5642);
   U9849 : NAND3_X1 port map( A1 => n5645, A2 => n5649, A3 => n5642, ZN => 
                           n5290);
   U9850 : XNOR2_X1 port map( A => n7006, B => n7266, ZN => n5296);
   U9851 : MUX2_X1 port map( A => n5699, B => n5971, S => n5968, Z => n5295);
   U9852 : INV_X1 port map( A => n5524, ZN => n5967);
   U9853 : NOR2_X1 port map( A1 => n5697, A2 => n5967, ZN => n5450);
   U9854 : NAND2_X1 port map( A1 => n5450, A2 => n5973, ZN => n5293);
   U9855 : NAND2_X1 port map( A1 => n957, A2 => n5971, ZN => n5292);
   U9856 : OAI211_X1 port map( C1 => n5295, C2 => n5294, A => n5293, B => n5292
                           , ZN => n6348);
   U9857 : INV_X1 port map( A => n6348, ZN => n7344);
   U9858 : XNOR2_X1 port map( A => n7344, B => n5296, ZN => n6835);
   U9859 : NAND3_X1 port map( A1 => n20001, A2 => n8301, A3 => n8303, ZN => 
                           n5298);
   U9860 : NAND2_X1 port map( A1 => n5792, A2 => n5300, ZN => n5303);
   U9861 : NOR2_X1 port map( A1 => n5798, A2 => n19912, ZN => n5302);
   U9862 : INV_X1 port map( A => n5300, ZN => n5790);
   U9863 : OAI211_X1 port map( C1 => n5304, C2 => n6059, A => n5895, B => n6057
                           , ZN => n5307);
   U9864 : INV_X1 port map( A => n6061, ZN => n5306);
   U9865 : XNOR2_X1 port map( A => n6687, B => n7338, ZN => n5315);
   U9866 : OAI21_X1 port map( B1 => n6044, B2 => n5309, A => n5308, ZN => n6047
                           );
   U9867 : NOR2_X1 port map( A1 => n6046, A2 => n5888, ZN => n5310);
   U9868 : NOR2_X1 port map( A1 => n5311, A2 => n5310, ZN => n5313);
   U9869 : INV_X1 port map( A => n5311, ZN => n5312);
   U9870 : INV_X1 port map( A => n6728, ZN => n5314);
   U9871 : XNOR2_X1 port map( A => n5315, B => n5314, ZN => n6630);
   U9872 : OAI21_X1 port map( B1 => n5582, B2 => n5581, A => n5317, ZN => n5406
                           );
   U9873 : INV_X1 port map( A => n5318, ZN => n5319);
   U9874 : INV_X1 port map( A => n6782, ZN => n5321);
   U9875 : XNOR2_X1 port map( A => n5321, B => n7134, ZN => n5690);
   U9876 : NOR2_X1 port map( A1 => n1838, A2 => n5398, ZN => n5327);
   U9877 : NAND2_X1 port map( A1 => n5397, A2 => n5323, ZN => n5324);
   U9878 : XNOR2_X1 port map( A => n7041, B => n18691, ZN => n5335);
   U9879 : NAND2_X1 port map( A1 => n5329, A2 => n5328, ZN => n5334);
   U9880 : NAND2_X1 port map( A1 => n6052, A2 => n6051, ZN => n5333);
   U9881 : NAND2_X1 port map( A1 => n5330, A2 => n6050, ZN => n5332);
   U9882 : NAND2_X1 port map( A1 => n5330, A2 => n6051, ZN => n5331);
   U9883 : NAND4_X1 port map( A1 => n5334, A2 => n5333, A3 => n5332, A4 => 
                           n5331, ZN => n6573);
   U9884 : INV_X1 port map( A => n6573, ZN => n6038);
   U9885 : XNOR2_X1 port map( A => n5335, B => n6038, ZN => n5336);
   U9886 : XNOR2_X1 port map( A => n5690, B => n5336, ZN => n5337);
   U9888 : NAND3_X1 port map( A1 => n5868, A2 => n5338, A3 => n6119, ZN => 
                           n5339);
   U9889 : NAND2_X1 port map( A1 => n5386, A2 => n6118, ZN => n6127);
   U9890 : AND2_X1 port map( A1 => n6127, A2 => n5339, ZN => n5340);
   U9891 : OAI21_X2 port map( B1 => n6128, B2 => n5341, A => n5340, ZN => n7087
                           );
   U9892 : INV_X1 port map( A => n6140, ZN => n5866);
   U9893 : NAND2_X1 port map( A1 => n5866, A2 => n5860, ZN => n5345);
   U9894 : OAI21_X1 port map( B1 => n20334, B2 => n6140, A => n5342, ZN => 
                           n5344);
   U9895 : INV_X1 port map( A => n6724, ZN => n6633);
   U9896 : XNOR2_X1 port map( A => n6633, B => n7087, ZN => n6237);
   U9897 : INV_X1 port map( A => n6237, ZN => n5354);
   U9898 : MUX2_X1 port map( A => n5604, B => n5605, S => n5716, Z => n5348);
   U9899 : NAND2_X1 port map( A1 => n5605, A2 => n5346, ZN => n5347);
   U9900 : OR2_X1 port map( A1 => n5610, A2 => n1277, ZN => n5352);
   U9901 : NAND2_X1 port map( A1 => n6153, A2 => n5349, ZN => n5351);
   U9902 : NAND3_X1 port map( A1 => n5611, A2 => n6156, A3 => n6159, ZN => 
                           n5350);
   U9903 : XNOR2_X1 port map( A => n5354, B => n6506, ZN => n5377);
   U9904 : NAND2_X1 port map( A1 => n5356, A2 => n5623, ZN => n5355);
   U9905 : AOI21_X1 port map( B1 => n5355, B2 => n5692, A => n6131, ZN => n5359
                           );
   U9906 : NAND2_X1 port map( A1 => n5691, A2 => n6131, ZN => n5357);
   U9907 : AOI21_X1 port map( B1 => n5621, B2 => n5357, A => n5356, ZN => n5358
                           );
   U9908 : INV_X1 port map( A => n7142, ZN => n6469);
   U9909 : INV_X1 port map( A => n5360, ZN => n5362);
   U9910 : NAND2_X1 port map( A1 => n5631, A2 => n5364, ZN => n5361);
   U9911 : AOI21_X1 port map( B1 => n5362, B2 => n5361, A => n4598, ZN => n5366
                           );
   U9912 : NAND2_X1 port map( A1 => n4598, A2 => n5363, ZN => n5629);
   U9913 : INV_X1 port map( A => n5633, ZN => n5466);
   U9914 : AOI21_X1 port map( B1 => n5629, B2 => n5466, A => n5364, ZN => n5365
                           );
   U9915 : NOR2_X1 port map( A1 => n5366, A2 => n5365, ZN => n7048);
   U9916 : INV_X1 port map( A => n7048, ZN => n6680);
   U9917 : XNOR2_X1 port map( A => n6469, B => n6680, ZN => n5375);
   U9918 : NAND2_X1 port map( A1 => n5392, A2 => n5367, ZN => n5372);
   U9919 : OAI21_X1 port map( B1 => n5394, B2 => n5398, A => n5395, ZN => n5370
                           );
   U9920 : NAND2_X1 port map( A1 => n5370, A2 => n5369, ZN => n5371);
   U9921 : XNOR2_X1 port map( A => n7316, B => n2123, ZN => n5374);
   U9922 : XNOR2_X1 port map( A => n5375, B => n5374, ZN => n5376);
   U9923 : OAI21_X1 port map( B1 => n5379, B2 => n6192, A => n5802, ZN => n5381
                           );
   U9924 : OAI211_X1 port map( C1 => n5733, C2 => n5382, A => n5381, B => n5380
                           , ZN => n6714);
   U9925 : NAND2_X1 port map( A1 => n5728, A2 => n5845, ZN => n5385);
   U9926 : NAND3_X1 port map( A1 => n6183, A2 => n5845, A3 => n6184, ZN => 
                           n5384);
   U9927 : XNOR2_X1 port map( A => n7065, B => n6714, ZN => n6640);
   U9928 : INV_X1 port map( A => n6640, ZN => n5403);
   U9929 : NAND3_X1 port map( A1 => n6120, A2 => n5386, A3 => n6119, ZN => 
                           n5391);
   U9930 : AND2_X1 port map( A1 => n6118, A2 => n6119, ZN => n5867);
   U9931 : NAND2_X1 port map( A1 => n5867, A2 => n6123, ZN => n5389);
   U9932 : NAND2_X1 port map( A1 => n5387, A2 => n6124, ZN => n5388);
   U9933 : INV_X1 port map( A => n5392, ZN => n5402);
   U9934 : OAI21_X1 port map( B1 => n5395, B2 => n5394, A => n5393, ZN => n5396
                           );
   U9935 : NAND2_X1 port map( A1 => n5396, A2 => n5401, ZN => n5400);
   U9936 : OAI211_X2 port map( C1 => n5402, C2 => n5401, A => n5400, B => n5399
                           , ZN => n6777);
   U9937 : XNOR2_X1 port map( A => n7128, B => n6777, ZN => n6488);
   U9938 : XNOR2_X1 port map( A => n5403, B => n6488, ZN => n5423);
   U9939 : NAND2_X1 port map( A1 => n5406, A2 => n5405, ZN => n5407);
   U9940 : OR2_X1 port map( A1 => n5410, A2 => n5682, ZN => n6081);
   U9941 : INV_X1 port map( A => n5683, ZN => n5479);
   U9942 : AOI21_X1 port map( B1 => n6081, B2 => n5479, A => n5476, ZN => n5414
                           );
   U9943 : AOI21_X1 port map( B1 => n5412, B2 => n5680, A => n5411, ZN => n5413
                           );
   U9944 : INV_X1 port map( A => n7014, ZN => n5415);
   U9945 : XNOR2_X1 port map( A => n19855, B => n5415, ZN => n5421);
   U9946 : NAND2_X1 port map( A1 => n6204, A2 => n19968, ZN => n5419);
   U9947 : INV_X1 port map( A => n19492, ZN => n5416);
   U9948 : OAI21_X1 port map( B1 => n19522, B2 => n5416, A => n6205, ZN => 
                           n5417);
   U9949 : NAND3_X1 port map( A1 => n6205, A2 => n19492, A3 => n3640, ZN => 
                           n5418);
   U9950 : XNOR2_X1 port map( A => n7296, B => n2376, ZN => n5420);
   U9951 : XNOR2_X1 port map( A => n5421, B => n5420, ZN => n5422);
   U9952 : MUX2_X1 port map( A => n5670, B => n5425, S => n5424, Z => n5427);
   U9953 : MUX2_X1 port map( A => n19912, B => n5796, S => n5428, Z => n5430);
   U9954 : MUX2_X2 port map( A => n5431, B => n5430, S => n5429, Z => n7253);
   U9955 : XNOR2_X1 port map( A => n7116, B => n7253, ZN => n5441);
   U9956 : INV_X1 port map( A => n5998, ZN => n5432);
   U9957 : NAND2_X1 port map( A1 => n5437, A2 => n5436, ZN => n7081);
   U9958 : MUX2_X1 port map( A => n5711, B => n5990, S => n5985, Z => n5440);
   U9959 : NOR2_X1 port map( A1 => n5815, A2 => n5989, ZN => n5988);
   U9960 : NOR2_X1 port map( A1 => n5988, A2 => n5438, ZN => n5439);
   U9961 : MUX2_X2 port map( A => n5440, B => n5439, S => n5818, Z => n7122);
   U9962 : XNOR2_X1 port map( A => n5441, B => n6621, ZN => n5454);
   U9963 : MUX2_X1 port map( A => n5442, B => n5641, S => n5444, Z => n5446);
   U9964 : MUX2_X1 port map( A => n5444, B => n5649, S => n5443, Z => n5445);
   U9965 : MUX2_X1 port map( A => n5825, B => n6017, S => n6016, Z => n5448);
   U9966 : XNOR2_X1 port map( A => n7257, B => n7121, ZN => n5599);
   U9968 : NAND3_X1 port map( A1 => n5973, A2 => n19804, A3 => n20673, ZN => 
                           n5451);
   U9969 : XNOR2_X1 port map( A => n7289, B => n2455, ZN => n5452);
   U9970 : XNOR2_X1 port map( A => n5599, B => n5452, ZN => n5453);
   U9971 : AOI21_X1 port map( B1 => n6107, B2 => n6104, A => n6105, ZN => n5455
                           );
   U9972 : NAND2_X1 port map( A1 => n5663, A2 => n6101, ZN => n5456);
   U9973 : OAI21_X1 port map( B1 => n5662, B2 => n5663, A => n5456, ZN => n5457
                           );
   U9974 : NAND2_X1 port map( A1 => n5457, A2 => n283, ZN => n5459);
   U9975 : INV_X1 port map( A => n6225, ZN => n6646);
   U9976 : INV_X1 port map( A => n5945, ZN => n6173);
   U9977 : NAND3_X1 port map( A1 => n1867, A2 => n170, A3 => n6173, ZN => n5460
                           );
   U9978 : NAND2_X1 port map( A1 => n5463, A2 => n4598, ZN => n5470);
   U9979 : NAND3_X1 port map( A1 => n5467, A2 => n5466, A3 => n31, ZN => n5468)
                           ;
   U9980 : XNOR2_X1 port map( A => n7160, B => n7263, ZN => n6484);
   U9981 : XNOR2_X1 port map( A => n6646, B => n6484, ZN => n5491);
   U9982 : INV_X1 port map( A => n5532, ZN => n5529);
   U9983 : OAI21_X1 port map( B1 => n5562, B2 => n2940, A => n5529, ZN => n5474
                           );
   U9984 : NOR2_X1 port map( A1 => n5532, A2 => n6036, ZN => n5565);
   U9985 : INV_X1 port map( A => n5565, ZN => n5473);
   U9986 : INV_X1 port map( A => n5566, ZN => n6034);
   U9987 : NAND2_X1 port map( A1 => n5476, A2 => n6083, ZN => n5478);
   U9988 : MUX2_X1 port map( A => n5478, B => n5477, S => n5684, Z => n5482);
   U9989 : NAND2_X1 port map( A1 => n5682, A2 => n5479, ZN => n6080);
   U9990 : OAI21_X1 port map( B1 => n5681, B2 => n5479, A => n6080, ZN => n5480
                           );
   U9991 : NAND2_X1 port map( A1 => n5480, A2 => n6082, ZN => n5481);
   U9992 : XNOR2_X1 port map( A => n7267, B => n7306, ZN => n5489);
   U9993 : NOR2_X1 port map( A1 => n5719, A2 => n5715, ZN => n5603);
   U9994 : NAND2_X1 port map( A1 => n5603, A2 => n5717, ZN => n5487);
   U9995 : NAND3_X1 port map( A1 => n5605, A2 => n5715, A3 => n5720, ZN => 
                           n5486);
   U9996 : AND2_X1 port map( A1 => n5719, A2 => n5483, ZN => n5602);
   U9997 : NAND3_X1 port map( A1 => n5718, A2 => n5604, A3 => n5715, ZN => 
                           n5484);
   U9998 : XNOR2_X1 port map( A => n7163, B => n2395, ZN => n5488);
   U9999 : XNOR2_X1 port map( A => n5489, B => n5488, ZN => n5490);
   U10000 : INV_X1 port map( A => n8034, ZN => n7603);
   U10001 : INV_X1 port map( A => n5492, ZN => n5900);
   U10003 : INV_X1 port map( A => n5497, ZN => n5498);
   U10004 : NAND3_X1 port map( A1 => n4632, A2 => n5741, A3 => n5746, ZN => 
                           n5499);
   U10007 : INV_X1 port map( A => n862, ZN => n5919);
   U10008 : NAND2_X1 port map( A1 => n5502, A2 => n5919, ZN => n5515);
   U10009 : INV_X1 port map( A => n5503, ZN => n5513);
   U10010 : INV_X1 port map( A => n5504, ZN => n5507);
   U10011 : INV_X1 port map( A => n5505, ZN => n5506);
   U10012 : NOR2_X1 port map( A1 => n5507, A2 => n5506, ZN => n5512);
   U10013 : INV_X1 port map( A => n5508, ZN => n5509);
   U10014 : AND2_X1 port map( A1 => n5510, A2 => n5509, ZN => n5511);
   U10015 : NAND4_X1 port map( A1 => n5513, A2 => n862, A3 => n5512, A4 => 
                           n5511, ZN => n5514);
   U10016 : NAND3_X1 port map( A1 => n6014, A2 => n5515, A3 => n5514, ZN => 
                           n5517);
   U10017 : NAND2_X1 port map( A1 => n5517, A2 => n5516, ZN => n6420);
   U10018 : NAND2_X1 port map( A1 => n5927, A2 => n6025, ZN => n5518);
   U10019 : NOR2_X1 port map( A1 => n5926, A2 => n6031, ZN => n5519);
   U10020 : XNOR2_X1 port map( A => n6420, B => n6736, ZN => n6626);
   U10021 : XNOR2_X1 port map( A => n6495, B => n6626, ZN => n5553);
   U10022 : NAND3_X1 port map( A1 => n5528, A2 => n5967, A3 => n5523, ZN => 
                           n5527);
   U10023 : NAND3_X1 port map( A1 => n5700, A2 => n5525, A3 => n19804, ZN => 
                           n5526);
   U10024 : OAI211_X1 port map( C1 => n5700, C2 => n5528, A => n5527, B => 
                           n5526, ZN => n7035);
   U10025 : NAND2_X1 port map( A1 => n6036, A2 => n20241, ZN => n5530);
   U10026 : NAND2_X1 port map( A1 => n5531, A2 => n6036, ZN => n5533);
   U10027 : OAI22_X1 port map( A1 => n5534, A2 => n5569, B1 => n5533, B2 => 
                           n5532, ZN => n5535);
   U10028 : NOR2_X1 port map( A1 => n5536, A2 => n5535, ZN => n6293);
   U10029 : INV_X1 port map( A => n6293, ZN => n7326);
   U10030 : XNOR2_X1 port map( A => n7326, B => n7035, ZN => n5551);
   U10031 : NAND2_X1 port map( A1 => n5736, A2 => n5734, ZN => n5544);
   U10032 : INV_X1 port map( A => n5537, ZN => n5542);
   U10033 : INV_X1 port map( A => n5538, ZN => n5541);
   U10034 : NAND4_X1 port map( A1 => n5542, A2 => n5541, A3 => n5540, A4 => 
                           n5539, ZN => n5543);
   U10035 : NAND3_X1 port map( A1 => n5544, A2 => n5768, A3 => n5543, ZN => 
                           n5549);
   U10036 : NAND3_X1 port map( A1 => n5736, A2 => n5734, A3 => n5765, ZN => 
                           n5548);
   U10037 : NAND3_X1 port map( A1 => n5546, A2 => n5735, A3 => n5545, ZN => 
                           n5547);
   U10039 : XNOR2_X1 port map( A => n7155, B => n2222, ZN => n5550);
   U10040 : XNOR2_X1 port map( A => n5551, B => n5550, ZN => n5552);
   U10041 : XNOR2_X1 port map( A => n5553, B => n5552, ZN => n8033);
   U10042 : OAI21_X1 port map( B1 => n7600, B2 => n8033, A => n7445, ZN => 
                           n5554);
   U10043 : INV_X1 port map( A => n8286, ZN => n7444);
   U10044 : NAND2_X1 port map( A1 => n5554, A2 => n7444, ZN => n5555);
   U10045 : OAI21_X1 port map( B1 => n7796, B2 => n8034, A => n5555, ZN => 
                           n5556);
   U10047 : NAND2_X1 port map( A1 => n5562, A2 => n6036, ZN => n5570);
   U10048 : OAI21_X1 port map( B1 => n5564, B2 => n20241, A => n5569, ZN => 
                           n5567);
   U10049 : MUX2_X1 port map( A => n5567, B => n5566, S => n5565, Z => n5568);
   U10050 : XNOR2_X1 port map( A => n7080, B => n7287, ZN => n6759);
   U10051 : NAND2_X1 port map( A1 => n5572, A2 => n5571, ZN => n5586);
   U10052 : INV_X1 port map( A => n5573, ZN => n5578);
   U10053 : NAND3_X1 port map( A1 => n5576, A2 => n5575, A3 => n5574, ZN => 
                           n5577);
   U10054 : OAI21_X1 port map( B1 => n5578, B2 => n5577, A => n5580, ZN => 
                           n5579);
   U10055 : OAI21_X1 port map( B1 => n5581, B2 => n5580, A => n5579, ZN => 
                           n5585);
   U10056 : XNOR2_X1 port map( A => n5884, B => n19158, ZN => n5587);
   U10057 : XNOR2_X1 port map( A => n6759, B => n5587, ZN => n5601);
   U10059 : NAND2_X1 port map( A1 => n20368, A2 => n5588, ZN => n5594);
   U10060 : NOR2_X1 port map( A1 => n5920, A2 => n19980, ZN => n5593);
   U10061 : NAND3_X1 port map( A1 => n5916, A2 => n6007, A3 => n19980, ZN => 
                           n5592);
   U10062 : INV_X1 port map( A => n7115, ZN => n5598);
   U10063 : INV_X1 port map( A => n5927, ZN => n5595);
   U10064 : XNOR2_X1 port map( A => n5598, B => n6819, ZN => n7285);
   U10065 : XNOR2_X1 port map( A => n7285, B => n5599, ZN => n5600);
   U10066 : XNOR2_X1 port map( A => n5600, B => n5601, ZN => n7420);
   U10067 : NAND2_X1 port map( A1 => n5602, A2 => n5720, ZN => n5609);
   U10068 : INV_X1 port map( A => n5603, ZN => n5608);
   U10069 : NAND3_X1 port map( A1 => n20034, A2 => n5715, A3 => n5483, ZN => 
                           n5606);
   U10072 : XNOR2_X1 port map( A => n6558, B => n7297, ZN => n6526);
   U10073 : INV_X1 port map( A => n6526, ZN => n6774);
   U10075 : NAND2_X1 port map( A1 => n5615, A2 => n6140, ZN => n5619);
   U10076 : NAND2_X1 port map( A1 => n6138, A2 => n5859, ZN => n5616);
   U10077 : NAND2_X1 port map( A1 => n5617, A2 => n6143, ZN => n5618);
   U10078 : INV_X1 port map( A => n6133, ZN => n6130);
   U10079 : AOI22_X1 port map( A1 => n5623, A2 => n5622, B1 => n6130, B2 => 
                           n5691, ZN => n5693);
   U10080 : INV_X1 port map( A => n6131, ZN => n5626);
   U10081 : OAI21_X1 port map( B1 => n5624, B2 => n5621, A => n6133, ZN => 
                           n5625);
   U10082 : OAI21_X1 port map( B1 => n5693, B2 => n5626, A => n5625, ZN => 
                           n6855);
   U10083 : XNOR2_X1 port map( A => n6855, B => n6713, ZN => n7295);
   U10084 : XNOR2_X1 port map( A => n6774, B => n7295, ZN => n5639);
   U10085 : NAND3_X1 port map( A1 => n5631, A2 => n4598, A3 => n5633, ZN => 
                           n5627);
   U10086 : OAI21_X1 port map( B1 => n5629, B2 => n5628, A => n5627, ZN => 
                           n5636);
   U10087 : AOI21_X1 port map( B1 => n5634, B2 => n5633, A => n5632, ZN => 
                           n5635);
   U10088 : INV_X1 port map( A => n6301, ZN => n6936);
   U10089 : XNOR2_X1 port map( A => n6936, B => n404, ZN => n5637);
   U10090 : XNOR2_X1 port map( A => n6488, B => n5637, ZN => n5638);
   U10091 : INV_X1 port map( A => n5640, ZN => n5654);
   U10092 : INV_X1 port map( A => n5641, ZN => n5644);
   U10093 : OAI21_X1 port map( B1 => n5644, B2 => n5643, A => n5642, ZN => 
                           n5653);
   U10094 : NAND3_X1 port map( A1 => n5647, A2 => n5646, A3 => n5645, ZN => 
                           n5652);
   U10096 : NAND2_X1 port map( A1 => n5650, A2 => n5649, ZN => n5651);
   U10098 : XNOR2_X1 port map( A => n6912, B => n18203, ZN => n5655);
   U10099 : XNOR2_X1 port map( A => n6495, B => n5655, ZN => n5689);
   U10100 : OAI21_X1 port map( B1 => n284, B2 => n6101, A => n5662, ZN => n5666
                           );
   U10101 : NAND2_X1 port map( A1 => n6097, A2 => n5949, ZN => n6096);
   U10103 : XNOR2_X1 port map( A => n6966, B => n6735, ZN => n7323);
   U10104 : NOR2_X1 port map( A1 => n5424, A2 => n5669, ZN => n5671);
   U10106 : OAI22_X1 port map( A1 => n5677, A2 => n5676, B1 => n3127, B2 => 
                           n5674, ZN => n5678);
   U10108 : OAI21_X1 port map( B1 => n5681, B2 => n6082, A => n5680, ZN => 
                           n5687);
   U10109 : NAND3_X1 port map( A1 => n5684, A2 => n6082, A3 => n6083, ZN => 
                           n5685);
   U10110 : XNOR2_X1 port map( A => n19765, B => n19698, ZN => n6752);
   U10111 : XNOR2_X1 port map( A => n7323, B => n6752, ZN => n5688);
   U10112 : XNOR2_X1 port map( A => n5689, B => n5688, ZN => n5762);
   U10113 : NOR2_X1 port map( A1 => n5691, A2 => n6131, ZN => n5695);
   U10114 : NAND2_X1 port map( A1 => n5698, A2 => n5970, ZN => n5702);
   U10115 : INV_X1 port map( A => n5699, ZN => n5972);
   U10116 : OAI211_X1 port map( C1 => n5973, C2 => n5967, A => n5972, B => 
                           n5700, ZN => n5701);
   U10117 : INV_X1 port map( A => n7332, ZN => n5703);
   U10118 : XNOR2_X1 port map( A => n5703, B => n7097, ZN => n6534);
   U10119 : INV_X1 port map( A => n5813, ZN => n5706);
   U10120 : AOI22_X1 port map( A1 => n5707, A2 => n6003, B1 => n5706, B2 => 
                           n5705, ZN => n7133);
   U10121 : INV_X1 port map( A => n7133, ZN => n6512);
   U10122 : NAND2_X1 port map( A1 => n5708, A2 => n5989, ZN => n5713);
   U10123 : OAI21_X1 port map( B1 => n5985, B2 => n5990, A => n3468, ZN => 
                           n5710);
   U10124 : NAND3_X1 port map( A1 => n5276, A2 => n5711, A3 => n5990, ZN => 
                           n5712);
   U10125 : INV_X1 port map( A => n6872, ZN => n6811);
   U10126 : NAND3_X1 port map( A1 => n5718, A2 => n5717, A3 => n5720, ZN => 
                           n5723);
   U10127 : NAND2_X1 port map( A1 => n5719, A2 => n5720, ZN => n5721);
   U10128 : XNOR2_X1 port map( A => n6917, B => n17637, ZN => n5725);
   U10129 : XNOR2_X1 port map( A => n7334, B => n5725, ZN => n5726);
   U10130 : NOR2_X1 port map( A1 => n8205, A2 => n8204, ZN => n5760);
   U10131 : MUX2_X1 port map( A => n6379, B => n5728, S => n19475, Z => n5729);
   U10132 : NOR2_X1 port map( A1 => n5729, A2 => n6183, ZN => n5731);
   U10133 : NAND2_X1 port map( A1 => n6192, A2 => n6189, ZN => n5732);
   U10134 : INV_X1 port map( A => n5736, ZN => n5770);
   U10136 : AND2_X1 port map( A1 => n5765, A2 => n5768, ZN => n5764);
   U10137 : NAND2_X1 port map( A1 => n5764, A2 => n5766, ZN => n5739);
   U10139 : XNOR2_X1 port map( A => n6767, B => n17089, ZN => n5754);
   U10140 : NAND2_X1 port map( A1 => n5742, A2 => n5741, ZN => n5753);
   U10141 : NAND2_X1 port map( A1 => n5750, A2 => n5749, ZN => n5751);
   U10142 : MUX2_X1 port map( A => n5226, B => n6204, S => n6206, Z => n5757);
   U10143 : NOR2_X1 port map( A1 => n6202, A2 => n19492, ZN => n5756);
   U10144 : NAND2_X1 port map( A1 => n6218, A2 => n19968, ZN => n5758);
   U10145 : INV_X1 port map( A => n5762, ZN => n7871);
   U10146 : NAND2_X1 port map( A1 => n5764, A2 => n5763, ZN => n5774);
   U10147 : NAND2_X1 port map( A1 => n5766, A2 => n5765, ZN => n5773);
   U10148 : NAND3_X1 port map( A1 => n5769, A2 => n5546, A3 => n5767, ZN => 
                           n5772);
   U10149 : NAND3_X1 port map( A1 => n5770, A2 => n5769, A3 => n5768, ZN => 
                           n5771);
   U10150 : XNOR2_X1 port map( A => n6927, B => n19140, ZN => n5775);
   U10151 : XNOR2_X1 port map( A => n6506, B => n5775, ZN => n5812);
   U10152 : NAND2_X1 port map( A1 => n6041, A2 => n6042, ZN => n5778);
   U10153 : NAND3_X1 port map( A1 => n6046, A2 => n6041, A3 => n5888, ZN => 
                           n5780);
   U10154 : NAND2_X1 port map( A1 => n6059, A2 => n5782, ZN => n5783);
   U10155 : OAI21_X1 port map( B1 => n6064, B2 => n6059, A => n5783, ZN => 
                           n5784);
   U10156 : NAND2_X1 port map( A1 => n5784, A2 => n5891, ZN => n5789);
   U10157 : NOR2_X1 port map( A1 => n6057, A2 => n6055, ZN => n5787);
   U10158 : INV_X1 port map( A => n6059, ZN => n5786);
   U10159 : AOI22_X1 port map( A1 => n5787, A2 => n5786, B1 => n5785, B2 => 
                           n6055, ZN => n5788);
   U10160 : NAND2_X1 port map( A1 => n5789, A2 => n5788, ZN => n6723);
   U10161 : XNOR2_X1 port map( A => n6839, B => n6723, ZN => n7313);
   U10162 : AND2_X1 port map( A1 => n5794, A2 => n5793, ZN => n5801);
   U10163 : MUX2_X1 port map( A => n5797, B => n5796, S => n19912, Z => n5799);
   U10164 : NAND2_X1 port map( A1 => n5799, A2 => n5798, ZN => n5800);
   U10165 : NAND2_X1 port map( A1 => n5801, A2 => n5800, ZN => n7317);
   U10166 : INV_X1 port map( A => n5803, ZN => n5806);
   U10167 : NOR2_X1 port map( A1 => n5806, A2 => n5805, ZN => n5810);
   U10168 : OAI21_X1 port map( B1 => n5803, B2 => n5802, A => n6194, ZN => 
                           n5809);
   U10169 : NAND3_X1 port map( A1 => n6193, A2 => n5806, A3 => n6189, ZN => 
                           n5807);
   U10170 : OAI211_X2 port map( C1 => n5809, C2 => n5810, A => n5808, B => 
                           n5807, ZN => n7091);
   U10171 : XNOR2_X1 port map( A => n7317, B => n7091, ZN => n6790);
   U10172 : XNOR2_X1 port map( A => n6790, B => n7313, ZN => n5811);
   U10173 : XNOR2_X1 port map( A => n5812, B => n5811, ZN => n7615);
   U10174 : INV_X1 port map( A => n5997, ZN => n5999);
   U10175 : NAND2_X1 port map( A1 => n5816, A2 => n5986, ZN => n5821);
   U10176 : NAND3_X1 port map( A1 => n5818, A2 => n285, A3 => n5817, ZN => 
                           n5819);
   U10177 : OAI211_X1 port map( C1 => n5988, C2 => n5821, A => n5820, B => 
                           n5819, ZN => n6754);
   U10178 : XNOR2_X1 port map( A => n7231, B => n6754, ZN => n6268);
   U10179 : INV_X1 port map( A => n6268, ZN => n6603);
   U10180 : XNOR2_X1 port map( A => n19765, B => n7364, ZN => n5822);
   U10181 : XNOR2_X1 port map( A => n6603, B => n5822, ZN => n5834);
   U10182 : NOR2_X1 port map( A1 => n3569, A2 => n5823, ZN => n6018);
   U10183 : AND2_X1 port map( A1 => n5825, A2 => n6016, ZN => n6020);
   U10184 : NAND2_X1 port map( A1 => n6020, A2 => n6022, ZN => n5830);
   U10185 : XNOR2_X1 port map( A => n6912, B => n7154, ZN => n6676);
   U10186 : XNOR2_X1 port map( A => n7035, B => n2284, ZN => n5832);
   U10187 : XNOR2_X1 port map( A => n6676, B => n5832, ZN => n5833);
   U10188 : XNOR2_X1 port map( A => n5833, B => n5834, ZN => n7453);
   U10189 : OAI21_X1 port map( B1 => n5226, B2 => n19968, A => n6204, ZN => 
                           n5837);
   U10190 : OAI21_X1 port map( B1 => n5839, B2 => n5838, A => n5837, ZN => 
                           n5840);
   U10191 : OAI21_X1 port map( B1 => n5846, B2 => n5845, A => n6184, ZN => 
                           n5849);
   U10192 : XNOR2_X1 port map( A => n6680, B => n7091, ZN => n5852);
   U10193 : XNOR2_X1 port map( A => n6985, B => n19243, ZN => n5851);
   U10194 : XNOR2_X1 port map( A => n5852, B => n5851, ZN => n5853);
   U10195 : NAND2_X1 port map( A1 => n7453, A2 => n8040, ZN => n7788);
   U10197 : INV_X1 port map( A => n5856, ZN => n5857);
   U10198 : XNOR2_X1 port map( A => n19780, B => n6917, ZN => n6686);
   U10199 : XNOR2_X1 port map( A => n7097, B => n6808, ZN => n5858);
   U10200 : XNOR2_X1 port map( A => n6686, B => n5858, ZN => n5878);
   U10201 : NAND2_X1 port map( A1 => n6143, A2 => n5860, ZN => n5863);
   U10202 : NAND2_X1 port map( A1 => n5861, A2 => n6141, ZN => n5862);
   U10203 : OAI21_X1 port map( B1 => n5864, B2 => n5863, A => n5862, ZN => 
                           n5865);
   U10204 : INV_X1 port map( A => n5867, ZN => n5874);
   U10205 : NAND3_X1 port map( A1 => n5870, A2 => n5869, A3 => n5868, ZN => 
                           n5872);
   U10206 : NAND2_X1 port map( A1 => n6124, A2 => n5873, ZN => n5871);
   U10207 : XNOR2_X1 port map( A => n6249, B => n6786, ZN => n6598);
   U10208 : INV_X1 port map( A => n2306, ZN => n5875);
   U10209 : XNOR2_X1 port map( A => n7041, B => n5875, ZN => n5876);
   U10210 : XNOR2_X1 port map( A => n6598, B => n5876, ZN => n5877);
   U10211 : XNOR2_X1 port map( A => n5878, B => n5877, ZN => n8041);
   U10212 : INV_X1 port map( A => n8041, ZN => n8298);
   U10213 : NOR2_X1 port map( A1 => n6068, A2 => n6067, ZN => n5881);
   U10214 : NOR2_X2 port map( A1 => n5883, A2 => n5882, ZN => n7118);
   U10215 : NAND3_X1 port map( A1 => n6044, A2 => n1007, A3 => n5885, ZN => 
                           n5886);
   U10216 : OAI21_X1 port map( B1 => n6041, B2 => n6044, A => n5886, ZN => 
                           n5887);
   U10217 : INV_X1 port map( A => n5887, ZN => n5890);
   U10219 : XNOR2_X1 port map( A => n6761, B => n7258, ZN => n6588);
   U10220 : XNOR2_X1 port map( A => n7080, B => n7253, ZN => n5897);
   U10221 : XNOR2_X1 port map( A => n6977, B => n2347, ZN => n5896);
   U10222 : XNOR2_X1 port map( A => n5897, B => n5896, ZN => n5898);
   U10223 : INV_X1 port map( A => n6942, ZN => n5913);
   U10224 : NAND2_X1 port map( A1 => n5900, A2 => n5899, ZN => n6091);
   U10225 : NOR2_X1 port map( A1 => n5902, A2 => n5901, ZN => n5906);
   U10226 : NAND4_X1 port map( A1 => n5906, A2 => n5905, A3 => n5904, A4 => 
                           n5903, ZN => n5907);
   U10227 : OAI21_X1 port map( B1 => n5199, B2 => n6087, A => n5907, ZN => 
                           n5909);
   U10228 : NAND2_X1 port map( A1 => n5909, A2 => n5908, ZN => n5911);
   U10229 : NAND3_X1 port map( A1 => n20149, A2 => n5199, A3 => n890, ZN => 
                           n5910);
   U10230 : OAI211_X1 port map( C1 => n5912, C2 => n6091, A => n5911, B => 
                           n5910, ZN => n7164);
   U10231 : XNOR2_X1 port map( A => n5913, B => n7164, ZN => n6692);
   U10233 : OAI21_X1 port map( B1 => n5914, B2 => n861, A => n5915, ZN => n5918
                           );
   U10234 : NAND2_X1 port map( A1 => n5918, A2 => n5917, ZN => n5925);
   U10235 : NAND3_X1 port map( A1 => n5919, A2 => n6007, A3 => n6013, ZN => 
                           n5923);
   U10236 : NAND3_X1 port map( A1 => n5921, A2 => n6010, A3 => n862, ZN => 
                           n5922);
   U10237 : AND2_X1 port map( A1 => n5923, A2 => n5922, ZN => n5924);
   U10238 : NAND2_X1 port map( A1 => n5925, A2 => n5924, ZN => n6946);
   U10239 : OAI21_X1 port map( B1 => n5595, B2 => n19790, A => n5926, ZN => 
                           n5935);
   U10240 : NOR2_X1 port map( A1 => n5927, A2 => n5930, ZN => n5934);
   U10241 : XNOR2_X1 port map( A => n6946, B => n6768, ZN => n6611);
   U10242 : INV_X1 port map( A => n6611, ZN => n5936);
   U10243 : XNOR2_X1 port map( A => n6692, B => n5936, ZN => n5940);
   U10244 : XNOR2_X1 port map( A => n6348, B => n7267, ZN => n5938);
   U10245 : XNOR2_X1 port map( A => n20225, B => n17686, ZN => n5937);
   U10246 : XNOR2_X1 port map( A => n5938, B => n5937, ZN => n5939);
   U10247 : INV_X1 port map( A => n7787, ZN => n5963);
   U10248 : INV_X1 port map( A => n6166, ZN => n5942);
   U10249 : AOI21_X1 port map( B1 => n5943, B2 => n6175, A => n5942, ZN => 
                           n5947);
   U10250 : NAND2_X1 port map( A1 => n6176, A2 => n6171, ZN => n5944);
   U10251 : AOI21_X1 port map( B1 => n5945, B2 => n5944, A => n6168, ZN => 
                           n5946);
   U10252 : XNOR2_X1 port map( A => n7127, B => n6936, ZN => n6665);
   U10253 : INV_X1 port map( A => n5948, ZN => n5951);
   U10254 : XNOR2_X1 port map( A => n7240, B => n941, ZN => n6606);
   U10255 : XNOR2_X1 port map( A => n6665, B => n6606, ZN => n5962);
   U10256 : INV_X1 port map( A => n7392, ZN => n5958);
   U10257 : XNOR2_X1 port map( A => n7014, B => n5958, ZN => n5960);
   U10258 : XNOR2_X1 port map( A => n6558, B => n2401, ZN => n5959);
   U10259 : XNOR2_X1 port map( A => n5960, B => n5959, ZN => n5961);
   U10262 : AND2_X1 port map( A1 => n5967, A2 => n5971, ZN => n5969);
   U10263 : INV_X1 port map( A => n5973, ZN => n5974);
   U10264 : NAND2_X1 port map( A1 => n5975, A2 => n5974, ZN => n5976);
   U10265 : XNOR2_X1 port map( A => n7372, B => n7142, ZN => n6721);
   U10266 : INV_X1 port map( A => n6721, ZN => n5983);
   U10267 : NAND2_X1 port map( A1 => n209, A2 => n5978, ZN => n5979);
   U10268 : AOI22_X1 port map( A1 => n5980, A2 => n6069, B1 => n6072, B2 => 
                           n6067, ZN => n5981);
   U10269 : XNOR2_X1 port map( A => n7047, B => n7088, ZN => n7315);
   U10270 : XNOR2_X1 port map( A => n7315, B => n5983, ZN => n6006);
   U10271 : XNOR2_X1 port map( A => n7272, B => n2410, ZN => n6004);
   U10272 : AND2_X1 port map( A1 => n5985, A2 => n5989, ZN => n5987);
   U10273 : OAI21_X1 port map( B1 => n5988, B2 => n5987, A => n5986, ZN => 
                           n5994);
   U10274 : INV_X1 port map( A => n5989, ZN => n5991);
   U10275 : NAND3_X1 port map( A1 => n5991, A2 => n285, A3 => n5990, ZN => 
                           n5992);
   U10276 : NAND3_X1 port map( A1 => n6000, A2 => n5999, A3 => n5998, ZN => 
                           n6001);
   U10277 : INV_X1 port map( A => n6328, ZN => n7177);
   U10278 : XNOR2_X1 port map( A => n7177, B => n6004, ZN => n6005);
   U10279 : OAI211_X1 port map( C1 => n6010, C2 => n19980, A => n20368, B => 
                           n6007, ZN => n6012);
   U10280 : INV_X1 port map( A => n2349, ZN => n6015);
   U10281 : XNOR2_X1 port map( A => n6990, B => n6015, ZN => n6024);
   U10282 : AOI21_X1 port map( B1 => n3569, B2 => n6017, A => n6016, ZN => 
                           n6021);
   U10283 : INV_X1 port map( A => n6021, ZN => n6023);
   U10285 : OAI211_X1 port map( C1 => n6027, C2 => n19789, A => n5595, B => 
                           n6025, ZN => n6029);
   U10286 : XNOR2_X1 port map( A => n6782, B => n7042, ZN => n6032);
   U10287 : XNOR2_X1 port map( A => n7382, B => n7336, ZN => n6039);
   U10288 : XNOR2_X1 port map( A => n6039, B => n6038, ZN => n6732);
   U10289 : NAND2_X1 port map( A1 => n6043, A2 => n6042, ZN => n6045);
   U10290 : AOI22_X2 port map( A1 => n6047, A2 => n6046, B1 => n6045, B2 => 
                           n6044, ZN => n6997);
   U10292 : XNOR2_X1 port map( A => n6997, B => n7018, ZN => n7193);
   U10293 : INV_X1 port map( A => n7193, ZN => n6066);
   U10294 : AOI21_X1 port map( B1 => n6056, B2 => n5782, A => n6058, ZN => 
                           n6063);
   U10295 : NOR2_X1 port map( A1 => n6058, A2 => n6057, ZN => n6060);
   U10296 : XNOR2_X1 port map( A => n7017, B => n6708, ZN => n7294);
   U10297 : INV_X1 port map( A => n7294, ZN => n6065);
   U10298 : XNOR2_X1 port map( A => n6065, B => n6066, ZN => n6079);
   U10299 : XNOR2_X1 port map( A => n6707, B => n7391, ZN => n6077);
   U10300 : XNOR2_X1 port map( A => n6777, B => n1148, ZN => n6076);
   U10301 : XNOR2_X1 port map( A => n6077, B => n6076, ZN => n6078);
   U10302 : NAND2_X1 port map( A1 => n6081, A2 => n6080, ZN => n6086);
   U10303 : MUX2_X1 port map( A => n6084, B => n6083, S => n6082, Z => n6085);
   U10305 : NAND2_X1 port map( A1 => n890, A2 => n6087, ZN => n6088);
   U10306 : NAND3_X1 port map( A1 => n6093, A2 => n6092, A3 => n6091, ZN => 
                           n6094);
   U10307 : XNOR2_X1 port map( A => n6095, B => n6718, ZN => n6116);
   U10308 : OAI21_X1 port map( B1 => n6098, B2 => n6097, A => n6096, ZN => 
                           n6103);
   U10309 : NAND2_X1 port map( A1 => n6100, A2 => n6099, ZN => n6102);
   U10310 : MUX2_X1 port map( A => n6105, B => n6104, S => n6109, Z => n6106);
   U10311 : INV_X1 port map( A => n6106, ZN => n6112);
   U10312 : XNOR2_X1 port map( A => n7218, B => n7221, ZN => n6337);
   U10313 : XNOR2_X1 port map( A => n7257, B => n2368, ZN => n6114);
   U10314 : XNOR2_X1 port map( A => n6337, B => n6114, ZN => n6115);
   U10315 : NAND2_X1 port map( A1 => n8196, A2 => n20198, ZN => n7628);
   U10316 : NOR2_X1 port map( A1 => n6119, A2 => n6118, ZN => n6121);
   U10317 : OAI21_X1 port map( B1 => n6122, B2 => n6121, A => n6120, ZN => 
                           n6126);
   U10318 : NAND3_X1 port map( A1 => n6124, A2 => n6128, A3 => n6123, ZN => 
                           n6125);
   U10319 : OAI211_X1 port map( C1 => n6128, C2 => n6127, A => n6126, B => 
                           n6125, ZN => n7009);
   U10320 : XNOR2_X1 port map( A => n7009, B => n6745, ZN => n7308);
   U10321 : MUX2_X1 port map( A => n6130, B => n6132, S => n6129, Z => n6137);
   U10322 : NAND2_X1 port map( A1 => n6132, A2 => n6131, ZN => n6135);
   U10323 : MUX2_X1 port map( A => n6135, B => n6134, S => n6133, Z => n6136);
   U10324 : OAI21_X2 port map( B1 => n6137, B2 => n5621, A => n6136, ZN => 
                           n7007);
   U10325 : MUX2_X1 port map( A => n6139, B => n6141, S => n6138, Z => n6147);
   U10326 : NAND2_X1 port map( A1 => n6141, A2 => n6140, ZN => n6145);
   U10327 : NAND2_X1 port map( A1 => n6148, A2 => n20334, ZN => n6144);
   U10328 : MUX2_X1 port map( A => n6145, B => n6144, S => n6143, Z => n6146);
   U10329 : XNOR2_X1 port map( A => n7007, B => n7206, ZN => n6349);
   U10330 : XNOR2_X1 port map( A => n6349, B => n7308, ZN => n6164);
   U10331 : NAND3_X1 port map( A1 => n6151, A2 => n6150, A3 => n6149, ZN => 
                           n6158);
   U10332 : OAI211_X1 port map( C1 => n6156, C2 => n6155, A => n6154, B => 
                           n6153, ZN => n6157);
   U10334 : INV_X1 port map( A => n2445, ZN => n6161);
   U10335 : XNOR2_X1 port map( A => n7263, B => n6161, ZN => n6162);
   U10336 : XNOR2_X1 port map( A => n6744, B => n6162, ZN => n6163);
   U10337 : XNOR2_X1 port map( A => n6164, B => n6163, ZN => n8192);
   U10338 : INV_X1 port map( A => n6165, ZN => n6180);
   U10339 : NAND2_X1 port map( A1 => n6167, A2 => n6171, ZN => n6169);
   U10340 : MUX2_X1 port map( A => n6170, B => n6169, S => n6168, Z => n6179);
   U10341 : NOR2_X1 port map( A1 => n6172, A2 => n6171, ZN => n6174);
   U10342 : NAND2_X1 port map( A1 => n6174, A2 => n6173, ZN => n6178);
   U10343 : XNOR2_X1 port map( A => n6180, B => n7032, ZN => n7324);
   U10344 : INV_X1 port map( A => n7324, ZN => n6546);
   U10345 : NOR2_X1 port map( A1 => n6379, A2 => n288, ZN => n6181);
   U10346 : OAI21_X1 port map( B1 => n6380, B2 => n6184, A => n6183, ZN => 
                           n6185);
   U10347 : NOR2_X1 port map( A1 => n6186, A2 => n6185, ZN => n6187);
   U10349 : MUX2_X1 port map( A => n6191, B => n6190, S => n6189, Z => n6198);
   U10350 : NAND2_X1 port map( A1 => n6193, A2 => n6192, ZN => n6196);
   U10352 : XNOR2_X1 port map( A => n19778, B => n7031, ZN => n6199);
   U10353 : XNOR2_X1 port map( A => n6546, B => n6199, ZN => n6210);
   U10354 : XNOR2_X1 port map( A => n7230, B => n484, ZN => n6209);
   U10355 : NAND2_X1 port map( A1 => n6218, A2 => n19492, ZN => n6201);
   U10356 : NAND2_X1 port map( A1 => n6220, A2 => n6204, ZN => n6208);
   U10357 : NOR2_X1 port map( A1 => n6206, A2 => n6205, ZN => n6219);
   U10358 : NAND2_X1 port map( A1 => n6219, A2 => n6218, ZN => n6207);
   U10359 : XNOR2_X1 port map( A => n6970, B => n7155, ZN => n6737);
   U10361 : NAND3_X1 port map( A1 => n9238, A2 => n9233, A3 => n8708, ZN => 
                           n6213);
   U10362 : XNOR2_X1 port map( A => n9819, B => n17791, ZN => n6658);
   U10363 : XNOR2_X1 port map( A => n7151, B => n19840, ZN => n6911);
   U10364 : XNOR2_X1 port map( A => n6165, B => n17791, ZN => n6216);
   U10365 : XNOR2_X1 port map( A => n6911, B => n6216, ZN => n6224);
   U10366 : XNOR2_X1 port map( A => n6736, B => n7360, ZN => n6222);
   U10367 : XNOR2_X1 port map( A => n6420, B => n19764, ZN => n7058);
   U10368 : XNOR2_X1 port map( A => n7058, B => n6222, ZN => n6223);
   U10369 : XNOR2_X1 port map( A => n20224, B => n6745, ZN => n7073);
   U10370 : XNOR2_X1 port map( A => n6225, B => n7073, ZN => n6228);
   U10371 : INV_X1 port map( A => n7160, ZN => n6226);
   U10372 : XNOR2_X1 port map( A => n6228, B => n6227, ZN => n7931);
   U10373 : XNOR2_X1 port map( A => n7080, B => n7354, ZN => n6565);
   U10374 : XNOR2_X1 port map( A => n6565, B => n19847, ZN => n6233);
   U10375 : XNOR2_X1 port map( A => n6719, B => n7121, ZN => n6231);
   U10376 : XNOR2_X1 port map( A => n7258, B => n18006, ZN => n6230);
   U10377 : XNOR2_X1 port map( A => n6231, B => n6230, ZN => n6232);
   U10378 : INV_X1 port map( A => n7372, ZN => n6234);
   U10379 : XNOR2_X1 port map( A => n7088, B => n6234, ZN => n6236);
   U10380 : XNOR2_X1 port map( A => n7091, B => n17932, ZN => n6235);
   U10381 : XNOR2_X1 port map( A => n6236, B => n6235, ZN => n6239);
   U10382 : XNOR2_X1 port map( A => n7146, B => n7274, ZN => n6925);
   U10383 : XNOR2_X1 port map( A => n6237, B => n6925, ZN => n6238);
   U10384 : INV_X1 port map( A => n7936, ZN => n7933);
   U10385 : XNOR2_X1 port map( A => n7240, B => n7128, ZN => n6935);
   U10386 : XNOR2_X1 port map( A => n6935, B => n6640, ZN => n6243);
   U10387 : XNOR2_X1 port map( A => n6558, B => n6708, ZN => n7066);
   U10388 : INV_X1 port map( A => n7066, ZN => n6241);
   U10389 : XNOR2_X1 port map( A => n7391, B => n18304, ZN => n6240);
   U10390 : XNOR2_X1 port map( A => n6241, B => n6240, ZN => n6242);
   U10391 : XNOR2_X1 port map( A => n6687, B => n649, ZN => n6246);
   U10392 : INV_X1 port map( A => n7097, ZN => n6783);
   U10393 : XNOR2_X1 port map( A => n6246, B => n6783, ZN => n6248);
   U10394 : XNOR2_X1 port map( A => n6728, B => n7382, ZN => n6247);
   U10395 : XNOR2_X1 port map( A => n6248, B => n6247, ZN => n6252);
   U10396 : XNOR2_X1 port map( A => n943, B => n7336, ZN => n6250);
   U10397 : XNOR2_X1 port map( A => n6250, B => n7134, ZN => n6251);
   U10398 : XNOR2_X1 port map( A => n6252, B => n6251, ZN => n7763);
   U10399 : NOR2_X1 port map( A1 => n7930, A2 => n1063, ZN => n6438);
   U10400 : INV_X1 port map( A => n7297, ZN => n6253);
   U10401 : XNOR2_X1 port map( A => n941, B => n6253, ZN => n6255);
   U10403 : XNOR2_X1 port map( A => n6777, B => n16788, ZN => n6254);
   U10404 : XNOR2_X1 port map( A => n6255, B => n6254, ZN => n6258);
   U10405 : XNOR2_X1 port map( A => n7240, B => n6641, ZN => n6256);
   U10406 : XNOR2_X1 port map( A => n7127, B => n6854, ZN => n6398);
   U10407 : XNOR2_X1 port map( A => n6256, B => n6398, ZN => n6257);
   U10408 : XNOR2_X2 port map( A => n6257, B => n6258, ZN => n7903);
   U10409 : XNOR2_X1 port map( A => n6611, B => n7305, ZN => n6262);
   U10410 : XNOR2_X1 port map( A => n7263, B => Key(63), ZN => n6259);
   U10411 : XNOR2_X1 port map( A => n6259, B => n6945, ZN => n6260);
   U10412 : XNOR2_X1 port map( A => n7164, B => n6850, ZN => n6393);
   U10413 : XNOR2_X1 port map( A => n6260, B => n6393, ZN => n6261);
   U10414 : XNOR2_X1 port map( A => n6261, B => n6262, ZN => n7530);
   U10415 : XNOR2_X1 port map( A => n7332, B => n2216, ZN => n6263);
   U10416 : XNOR2_X1 port map( A => n6263, B => n6598, ZN => n6266);
   U10417 : XNOR2_X1 port map( A => n6782, B => n6919, ZN => n7247);
   U10418 : XNOR2_X1 port map( A => n6873, B => n7137, ZN => n6368);
   U10419 : INV_X1 port map( A => n6368, ZN => n6264);
   U10420 : XNOR2_X1 port map( A => n6264, B => n7247, ZN => n6265);
   U10421 : XNOR2_X1 port map( A => n6265, B => n6266, ZN => n6904);
   U10422 : INV_X1 port map( A => n6904, ZN => n7902);
   U10423 : INV_X1 port map( A => n6494, ZN => n6545);
   U10424 : XNOR2_X1 port map( A => n6545, B => n7230, ZN => n6267);
   U10425 : XNOR2_X1 port map( A => n6268, B => n6267, ZN => n6271);
   U10426 : XNOR2_X1 port map( A => n19699, B => n18338, ZN => n6269);
   U10427 : XNOR2_X1 port map( A => n7154, B => n7365, ZN => n6364);
   U10428 : XNOR2_X1 port map( A => n6269, B => n6364, ZN => n6270);
   U10429 : XNOR2_X1 port map( A => n6271, B => n6270, ZN => n7002);
   U10430 : BUF_X2 port map( A => n7002, Z => n7909);
   U10431 : NOR2_X1 port map( A1 => n7902, A2 => n7909, ZN => n6272);
   U10432 : XNOR2_X1 port map( A => n7272, B => n7317, ZN => n6274);
   U10433 : XNOR2_X1 port map( A => n6634, B => n18011, ZN => n6273);
   U10434 : XNOR2_X1 port map( A => n6274, B => n6273, ZN => n6276);
   U10435 : XNOR2_X1 port map( A => n6593, B => n6374, ZN => n6275);
   U10436 : XNOR2_X1 port map( A => n6276, B => n6275, ZN => n7908);
   U10437 : INV_X1 port map( A => n7118, ZN => n6384);
   U10438 : XNOR2_X1 port map( A => n6384, B => n6520, ZN => n6277);
   U10439 : XNOR2_X1 port map( A => n6277, B => n6588, ZN => n6282);
   U10440 : INV_X1 port map( A => n7257, ZN => n6278);
   U10441 : XNOR2_X1 port map( A => n6278, B => n1053, ZN => n6280);
   U10442 : XNOR2_X1 port map( A => n19730, B => n17587, ZN => n6279);
   U10443 : XNOR2_X1 port map( A => n6280, B => n6279, ZN => n6281);
   U10444 : NAND2_X1 port map( A1 => n7754, A2 => n7903, ZN => n6283);
   U10445 : XNOR2_X1 port map( A => n5884, B => n6477, ZN => n7356);
   U10446 : XNOR2_X1 port map( A => n7254, B => n7289, ZN => n7078);
   U10447 : XNOR2_X1 port map( A => n7356, B => n7078, ZN => n6289);
   U10448 : INV_X1 port map( A => n6285, ZN => n6661);
   U10449 : XNOR2_X1 port map( A => n6661, B => n7216, ZN => n6287);
   U10450 : XNOR2_X1 port map( A => n19730, B => n2423, ZN => n6286);
   U10451 : XNOR2_X1 port map( A => n6287, B => n6286, ZN => n6288);
   U10452 : XNOR2_X1 port map( A => n6289, B => n6288, ZN => n7919);
   U10454 : XNOR2_X1 port map( A => n6942, B => n6693, ZN => n7346);
   U10455 : XNOR2_X1 port map( A => n6850, B => n6947, ZN => n6446);
   U10456 : XNOR2_X1 port map( A => n7346, B => n6446, ZN => n6292);
   U10457 : XNOR2_X1 port map( A => n7201, B => n7266, ZN => n6346);
   U10458 : XNOR2_X1 port map( A => n7306, B => n2375, ZN => n6290);
   U10459 : XNOR2_X1 port map( A => n6346, B => n6290, ZN => n6291);
   U10460 : XNOR2_X1 port map( A => n6362, B => n6912, ZN => n7361);
   U10461 : INV_X1 port map( A => n7057, ZN => n6294);
   U10462 : XNOR2_X1 port map( A => n6294, B => n7361, ZN => n6298);
   U10463 : XNOR2_X1 port map( A => n6674, B => n6738, ZN => n6296);
   U10464 : XNOR2_X1 port map( A => n7365, B => n16035, ZN => n6295);
   U10465 : XNOR2_X1 port map( A => n6296, B => n6295, ZN => n6297);
   U10466 : INV_X1 port map( A => n7978, ZN => n6299);
   U10467 : XNOR2_X1 port map( A => n6711, B => n6300, ZN => n6355);
   U10468 : XNOR2_X1 port map( A => n6301, B => n6489, ZN => n7395);
   U10469 : XNOR2_X1 port map( A => n7395, B => n6355, ZN => n6305);
   U10470 : XNOR2_X1 port map( A => n6776, B => n6854, ZN => n6303);
   U10471 : XNOR2_X1 port map( A => n7296, B => n1911, ZN => n6302);
   U10472 : XNOR2_X1 port map( A => n6303, B => n6302, ZN => n6304);
   U10474 : INV_X1 port map( A => n6679, ZN => n6307);
   U10475 : XNOR2_X1 port map( A => n6927, B => n645, ZN => n6308);
   U10476 : XNOR2_X1 port map( A => n6309, B => n6308, ZN => n6311);
   U10477 : XNOR2_X1 port map( A => n7316, B => n7373, ZN => n6505);
   U10478 : XNOR2_X1 port map( A => n7273, B => n7179, ZN => n6327);
   U10479 : XNOR2_X1 port map( A => n6505, B => n6327, ZN => n6310);
   U10480 : NAND2_X1 port map( A1 => n7982, A2 => n7984, ZN => n7110);
   U10481 : XNOR2_X1 port map( A => n7249, B => n7184, ZN => n6334);
   U10482 : INV_X1 port map( A => n7338, ZN => n6313);
   U10483 : XNOR2_X1 port map( A => n7384, B => n6313, ZN => n6514);
   U10484 : XNOR2_X1 port map( A => n6514, B => n6334, ZN => n6317);
   U10485 : XNOR2_X1 port map( A => n6873, B => n6917, ZN => n6315);
   U10486 : XNOR2_X1 port map( A => n7248, B => n2341, ZN => n6314);
   U10487 : XNOR2_X1 port map( A => n6314, B => n6315, ZN => n6316);
   U10489 : NAND2_X1 port map( A1 => n7110, A2 => n6318, ZN => n6319);
   U10491 : NAND2_X1 port map( A1 => n8470, A2 => n20010, ZN => n6442);
   U10492 : XNOR2_X1 port map( A => n7325, B => n1904, ZN => n6321);
   U10493 : XNOR2_X1 port map( A => n6321, B => n6735, ZN => n6323);
   U10494 : XNOR2_X1 port map( A => n7232, B => n7364, ZN => n6322);
   U10495 : XNOR2_X1 port map( A => n6323, B => n6322, ZN => n6326);
   U10496 : XNOR2_X1 port map( A => n6738, B => n7031, ZN => n6325);
   U10497 : INV_X1 port map( A => n19778, ZN => n6324);
   U10498 : XNOR2_X1 port map( A => n6325, B => n6324, ZN => n7214);
   U10499 : XNOR2_X1 port map( A => n7214, B => n6326, ZN => n6344);
   U10500 : INV_X1 port map( A => n6344, ZN => n8355);
   U10501 : XNOR2_X1 port map( A => n6328, B => n6327, ZN => n6332);
   U10502 : XNOR2_X1 port map( A => n6723, B => n7318, ZN => n6330);
   U10503 : XNOR2_X1 port map( A => n6985, B => n2392, ZN => n6329);
   U10504 : XNOR2_X1 port map( A => n6330, B => n6329, ZN => n6331);
   U10505 : NAND2_X1 port map( A1 => n8355, A2 => n7739, ZN => n7501);
   U10506 : INV_X1 port map( A => n7501, ZN => n6343);
   U10507 : XNOR2_X1 port map( A => n899, B => n2257, ZN => n6333);
   U10508 : XNOR2_X1 port map( A => n7042, B => n6990, ZN => n7185);
   U10509 : XNOR2_X1 port map( A => n7185, B => n6333, ZN => n6336);
   U10510 : XNOR2_X1 port map( A => n6808, B => n7337, ZN => n6992);
   U10511 : XNOR2_X1 port map( A => n6334, B => n6992, ZN => n6335);
   U10512 : NOR2_X1 port map( A1 => n8354, A2 => n7739, ZN => n6342);
   U10513 : XNOR2_X1 port map( A => n6478, B => n7216, ZN => n6717);
   U10514 : XNOR2_X1 port map( A => n6717, B => n6337, ZN => n6341);
   U10515 : XNOR2_X1 port map( A => n7254, B => n7288, ZN => n6339);
   U10516 : XNOR2_X1 port map( A => n6977, B => n2100, ZN => n6338);
   U10517 : XNOR2_X1 port map( A => n6339, B => n6338, ZN => n6340);
   U10518 : XNOR2_X1 port map( A => n6341, B => n6340, ZN => n6345);
   U10519 : OAI21_X1 port map( B1 => n6343, B2 => n6342, A => n7743, ZN => 
                           n6361);
   U10520 : NAND2_X1 port map( A1 => n8359, A2 => n7739, ZN => n6359);
   U10521 : XNOR2_X1 port map( A => n6743, B => n2420, ZN => n6347);
   U10522 : XNOR2_X1 port map( A => n6346, B => n6347, ZN => n6351);
   U10524 : XNOR2_X1 port map( A => n6961, B => n6349, ZN => n6350);
   U10525 : XNOR2_X1 port map( A => n6350, B => n6351, ZN => n7741);
   U10526 : NAND2_X1 port map( A1 => n7504, A2 => n7741, ZN => n6358);
   U10527 : XNOR2_X1 port map( A => n7392, B => n6352, ZN => n6995);
   U10528 : INV_X1 port map( A => n6995, ZN => n6354);
   U10529 : XNOR2_X1 port map( A => n6713, B => n1996, ZN => n6353);
   U10530 : XNOR2_X1 port map( A => n6354, B => n6353, ZN => n6357);
   U10531 : XNOR2_X1 port map( A => n7193, B => n6355, ZN => n6356);
   U10532 : MUX2_X1 port map( A => n6359, B => n6358, S => n8358, Z => n6360);
   U10533 : NOR2_X1 port map( A1 => n8128, A2 => n8884, ZN => n9089);
   U10534 : XNOR2_X1 port map( A => n6967, B => n7363, ZN => n6363);
   U10535 : XNOR2_X1 port map( A => n6362, B => n7035, ZN => n6672);
   U10536 : XNOR2_X1 port map( A => n6672, B => n6363, ZN => n6367);
   U10537 : XNOR2_X1 port map( A => n7212, B => n1857, ZN => n6365);
   U10538 : XNOR2_X1 port map( A => n6365, B => n6364, ZN => n6366);
   U10539 : XNOR2_X1 port map( A => n6367, B => n6366, ZN => n6951);
   U10540 : INV_X1 port map( A => n6951, ZN => n8361);
   U10541 : XNOR2_X1 port map( A => n7041, B => n7384, ZN => n6689);
   U10542 : XNOR2_X1 port map( A => n6368, B => n6689, ZN => n6372);
   U10543 : XNOR2_X1 port map( A => n6918, B => n19944, ZN => n6370);
   U10544 : XNOR2_X1 port map( A => n6990, B => n19216, ZN => n6369);
   U10545 : XNOR2_X1 port map( A => n6370, B => n6369, ZN => n6371);
   U10546 : INV_X1 port map( A => n7709, ZN => n8360);
   U10547 : XNOR2_X1 port map( A => n6982, B => n6680, ZN => n6373);
   U10548 : XNOR2_X1 port map( A => n6374, B => n6373, ZN => n6378);
   U10549 : XNOR2_X1 port map( A => n7046, B => n7373, ZN => n6376);
   U10550 : XNOR2_X1 port map( A => n6376, B => n6375, ZN => n6377);
   U10551 : XNOR2_X1 port map( A => n6378, B => n6377, ZN => n7673);
   U10552 : OAI21_X1 port map( B1 => n8361, B2 => n8360, A => n7673, ZN => 
                           n6390);
   U10553 : MUX2_X1 port map( A => n19476, B => n6380, S => n6379, Z => n6383);
   U10554 : XNOR2_X1 port map( A => n6384, B => n7355, ZN => n6385);
   U10556 : XNOR2_X1 port map( A => n6385, B => n6660, ZN => n6389);
   U10557 : XNOR2_X1 port map( A => n6867, B => n7218, ZN => n6387);
   U10558 : XNOR2_X1 port map( A => n6386, B => n6387, ZN => n6388);
   U10559 : XNOR2_X2 port map( A => n6389, B => n6388, ZN => n7675);
   U10560 : NAND2_X1 port map( A1 => n6390, A2 => n7675, ZN => n6402);
   U10561 : AND2_X1 port map( A1 => n7709, A2 => n7673, ZN => n8364);
   U10562 : XNOR2_X1 port map( A => n7006, B => n18284, ZN => n6391);
   U10563 : XNOR2_X1 port map( A => n6391, B => n7206, ZN => n6392);
   U10564 : XNOR2_X1 port map( A => n6693, B => n7267, ZN => n6612);
   U10565 : XNOR2_X1 port map( A => n6392, B => n6612, ZN => n6395);
   U10566 : XNOR2_X1 port map( A => n7345, B => n6393, ZN => n6394);
   U10567 : NAND2_X1 port map( A1 => n8364, A2 => n7674, ZN => n6401);
   U10568 : XNOR2_X1 port map( A => n6997, B => n632, ZN => n6397);
   U10569 : XNOR2_X1 port map( A => n7195, B => n7390, ZN => n6396);
   U10570 : XNOR2_X1 port map( A => n6397, B => n6396, ZN => n6400);
   U10571 : XNOR2_X1 port map( A => n6489, B => n7014, ZN => n6666);
   U10572 : XNOR2_X1 port map( A => n6666, B => n6398, ZN => n6399);
   U10573 : NOR2_X1 port map( A1 => n9453, A2 => n6438, ZN => n6403);
   U10574 : NAND2_X1 port map( A1 => n9089, A2 => n6403, ZN => n6441);
   U10575 : XNOR2_X1 port map( A => n6404, B => n7196, ZN => n7126);
   U10576 : INV_X1 port map( A => n7126, ZN => n6557);
   U10577 : XNOR2_X1 port map( A => n6557, B => n7295, ZN => n6407);
   U10578 : XNOR2_X1 port map( A => n7017, B => n7065, ZN => n6773);
   U10579 : XNOR2_X1 port map( A => n7013, B => n2424, ZN => n6405);
   U10580 : XNOR2_X1 port map( A => n6773, B => n6405, ZN => n6406);
   U10581 : XNOR2_X2 port map( A => n6407, B => n6406, ZN => n7749);
   U10582 : INV_X1 port map( A => n7116, ZN => n6409);
   U10583 : XNOR2_X1 port map( A => n7115, B => n17170, ZN => n6408);
   U10584 : XNOR2_X1 port map( A => n6408, B => n6409, ZN => n6412);
   U10585 : XNOR2_X1 port map( A => n6410, B => n7081, ZN => n6411);
   U10586 : XNOR2_X1 port map( A => n6412, B => n6411, ZN => n6415);
   U10587 : XNOR2_X1 port map( A => n7026, B => n6819, ZN => n6413);
   U10588 : XNOR2_X1 port map( A => n6413, B => n20203, ZN => n6414);
   U10589 : XNOR2_X1 port map( A => n7070, B => n7202, ZN => n6416);
   U10590 : XNOR2_X1 port map( A => n7303, B => n6416, ZN => n6419);
   U10591 : XNOR2_X1 port map( A => n7163, B => n7264, ZN => n6443);
   U10592 : XNOR2_X1 port map( A => n179, B => n2344, ZN => n6417);
   U10593 : XNOR2_X1 port map( A => n6443, B => n6417, ZN => n6418);
   U10594 : XNOR2_X1 port map( A => n6419, B => n6418, ZN => n7914);
   U10595 : INV_X1 port map( A => n7914, ZN => n7746);
   U10596 : INV_X1 port map( A => n6420, ZN => n6675);
   U10597 : XNOR2_X1 port map( A => n6675, B => n7032, ZN => n6422);
   U10598 : XNOR2_X1 port map( A => n7155, B => n18090, ZN => n6421);
   U10599 : XNOR2_X1 port map( A => n6422, B => n6421, ZN => n6425);
   U10600 : XNOR2_X1 port map( A => n6883, B => n6423, ZN => n6424);
   U10601 : XNOR2_X1 port map( A => n7383, B => n7333, ZN => n6426);
   U10602 : XNOR2_X1 port map( A => n7334, B => n6426, ZN => n6431);
   U10603 : XNOR2_X1 port map( A => n6427, B => n6573, ZN => n7135);
   U10604 : INV_X1 port map( A => n7135, ZN => n6429);
   U10605 : XNOR2_X1 port map( A => n6687, B => n875, ZN => n6428);
   U10606 : XNOR2_X1 port map( A => n6429, B => n6428, ZN => n6430);
   U10607 : XNOR2_X1 port map( A => n6431, B => n6430, ZN => n7508);
   U10608 : INV_X1 port map( A => n7087, ZN => n6432);
   U10609 : XNOR2_X1 port map( A => n7047, B => n6432, ZN => n6433);
   U10610 : XNOR2_X1 port map( A => n7313, B => n6433, ZN => n6437);
   U10611 : XNOR2_X1 port map( A => n7371, B => n6469, ZN => n6435);
   U10612 : XNOR2_X1 port map( A => n7144, B => n17999, ZN => n6434);
   U10613 : XNOR2_X1 port map( A => n6435, B => n6434, ZN => n6436);
   U10614 : INV_X1 port map( A => n6438, ZN => n8126);
   U10615 : INV_X1 port map( A => n6443, ZN => n6445);
   U10616 : XNOR2_X1 port map( A => n7007, B => n17851, ZN => n6444);
   U10617 : XNOR2_X1 port map( A => n6445, B => n6444, ZN => n6448);
   U10618 : XNOR2_X1 port map( A => n6446, B => n6961, ZN => n6447);
   U10619 : XNOR2_X1 port map( A => n7116, B => n7221, ZN => n6449);
   U10620 : XNOR2_X1 port map( A => n6864, B => n6449, ZN => n6452);
   U10621 : XNOR2_X1 port map( A => n6661, B => n610, ZN => n6450);
   U10622 : XNOR2_X1 port map( A => n7353, B => n6450, ZN => n6451);
   U10623 : XNOR2_X1 port map( A => n6452, B => n6451, ZN => n6467);
   U10624 : XNOR2_X1 port map( A => n6707, B => n2023, ZN => n6453);
   U10625 : XNOR2_X1 port map( A => n6776, B => n7018, ZN => n6669);
   U10626 : XNOR2_X1 port map( A => n6453, B => n6669, ZN => n6455);
   U10627 : XNOR2_X1 port map( A => n7013, B => n6854, ZN => n7397);
   U10628 : XNOR2_X1 port map( A => n7397, B => n6995, ZN => n6454);
   U10629 : XNOR2_X1 port map( A => n7364, B => n7031, ZN => n6456);
   U10630 : XNOR2_X1 port map( A => n6881, B => n6456, ZN => n6460);
   U10631 : XNOR2_X1 port map( A => n6674, B => n7155, ZN => n6458);
   U10632 : XNOR2_X1 port map( A => n7365, B => n18478, ZN => n6457);
   U10633 : XNOR2_X1 port map( A => n6458, B => n6457, ZN => n6459);
   U10634 : XNOR2_X1 port map( A => n7383, B => n6573, ZN => n6463);
   U10635 : INV_X1 port map( A => n20593, ZN => n6461);
   U10636 : XNOR2_X1 port map( A => n7337, B => n6461, ZN => n6462);
   U10637 : XNOR2_X1 port map( A => n6463, B => n6462, ZN => n6466);
   U10638 : XNOR2_X1 port map( A => n7248, B => n7042, ZN => n6685);
   U10639 : XNOR2_X1 port map( A => n6464, B => n6685, ZN => n6465);
   U10640 : XNOR2_X1 port map( A => n6466, B => n6465, ZN => n7644);
   U10641 : NAND2_X1 port map( A1 => n8219, A2 => n7644, ZN => n7646);
   U10642 : INV_X1 port map( A => n6467, ZN => n8079);
   U10643 : NAND3_X1 port map( A1 => n7646, A2 => n8079, A3 => n6468, ZN => 
                           n6475);
   U10644 : INV_X1 port map( A => n8076, ZN => n7645);
   U10645 : XNOR2_X1 port map( A => n7377, B => n6889, ZN => n6473);
   U10646 : XNOR2_X1 port map( A => n6679, B => n6469, ZN => n6471);
   U10647 : XNOR2_X1 port map( A => n7050, B => n19052, ZN => n6470);
   U10648 : XNOR2_X1 port map( A => n6471, B => n6470, ZN => n6472);
   U10649 : NAND3_X1 port map( A1 => n8220, A2 => n7645, A3 => n8219, ZN => 
                           n6474);
   U10650 : XNOR2_X1 port map( A => n7289, B => n6520, ZN => n6619);
   U10651 : XNOR2_X1 port map( A => n6761, B => n20227, ZN => n6476);
   U10652 : XNOR2_X1 port map( A => n6619, B => n6476, ZN => n6482);
   U10653 : XNOR2_X1 port map( A => n6477, B => n7257, ZN => n6480);
   U10654 : XNOR2_X1 port map( A => n6478, B => n2151, ZN => n6479);
   U10655 : XNOR2_X1 port map( A => n6480, B => n6479, ZN => n6481);
   U10656 : XNOR2_X1 port map( A => n6743, B => n6693, ZN => n6483);
   U10657 : XNOR2_X1 port map( A => n6768, B => n7306, ZN => n7074);
   U10658 : XNOR2_X1 port map( A => n7074, B => n6483, ZN => n6487);
   U10659 : XNOR2_X1 port map( A => n6945, B => n2446, ZN => n6485);
   U10660 : XNOR2_X1 port map( A => n6485, B => n6484, ZN => n6486);
   U10661 : XNOR2_X1 port map( A => n6487, B => n6486, ZN => n8113);
   U10662 : XNOR2_X1 port map( A => n7064, B => n6488, ZN => n6493);
   U10663 : XNOR2_X1 port map( A => n6489, B => n6641, ZN => n6491);
   U10664 : INV_X1 port map( A => n2305, ZN => n18389);
   U10665 : XNOR2_X1 port map( A => n6713, B => n18389, ZN => n6490);
   U10666 : XNOR2_X1 port map( A => n6491, B => n6490, ZN => n6492);
   U10667 : NAND3_X1 port map( A1 => n8253, A2 => n7844, A3 => n8114, ZN => 
                           n6519);
   U10668 : AND2_X1 port map( A1 => n6702, A2 => n8113, ZN => n8254);
   U10669 : XNOR2_X1 port map( A => n6495, B => n6625, ZN => n6504);
   U10670 : XNOR2_X1 port map( A => n6735, B => n19850, ZN => n6502);
   U10671 : NAND3_X1 port map( A1 => n6496, A2 => n641, A3 => n6500, ZN => 
                           n6499);
   U10672 : INV_X1 port map( A => n6496, ZN => n6497);
   U10673 : INV_X1 port map( A => n641, ZN => n18379);
   U10674 : NAND2_X1 port map( A1 => n6497, A2 => n18379, ZN => n6498);
   U10675 : OAI211_X1 port map( C1 => n641, C2 => n6500, A => n6499, B => n6498
                           , ZN => n6501);
   U10676 : XNOR2_X1 port map( A => n6502, B => n6501, ZN => n6503);
   U10677 : XNOR2_X1 port map( A => n6504, B => n6503, ZN => n6510);
   U10678 : NAND2_X1 port map( A1 => n8254, A2 => n7560, ZN => n6518);
   U10679 : XNOR2_X1 port map( A => n6723, B => n6793, ZN => n6508);
   U10680 : XNOR2_X1 port map( A => n6634, B => n18863, ZN => n6507);
   U10681 : XNOR2_X1 port map( A => n6508, B => n6507, ZN => n6509);
   U10682 : NAND2_X1 port map( A1 => n7560, A2 => n8245, ZN => n6517);
   U10683 : XNOR2_X1 port map( A => n6512, B => n6511, ZN => n6730);
   U10684 : XNOR2_X1 port map( A => n6513, B => n16651, ZN => n6515);
   U10685 : NAND3_X1 port map( A1 => n8248, A2 => n8251, A3 => n7844, ZN => 
                           n6516);
   U10686 : NAND4_X1 port map( A1 => n6519, A2 => n6518, A3 => n6517, A4 => 
                           n6516, ZN => n8713);
   U10687 : XNOR2_X1 port map( A => n7286, B => n6759, ZN => n6524);
   U10688 : XNOR2_X1 port map( A => n6520, B => n7218, ZN => n6522);
   U10689 : XNOR2_X1 port map( A => n7122, B => n18984, ZN => n6521);
   U10690 : XNOR2_X1 port map( A => n6522, B => n6521, ZN => n6523);
   U10691 : INV_X1 port map( A => n6997, ZN => n6525);
   U10692 : XNOR2_X1 port map( A => n6525, B => n6714, ZN => n6856);
   U10693 : XNOR2_X1 port map( A => n6526, B => n6856, ZN => n6529);
   U10694 : XNOR2_X1 port map( A => n6641, B => n2035, ZN => n6527);
   U10695 : XNOR2_X1 port map( A => n7294, B => n6527, ZN => n6528);
   U10696 : XNOR2_X1 port map( A => n6529, B => n6528, ZN => n8087);
   U10697 : XNOR2_X1 port map( A => n6982, B => n6633, ZN => n6887);
   U10698 : XNOR2_X1 port map( A => n20455, B => n7315, ZN => n6533);
   U10699 : INV_X1 port map( A => n17060, ZN => n6530);
   U10700 : XNOR2_X1 port map( A => n6634, B => n6530, ZN => n6531);
   U10701 : XNOR2_X1 port map( A => n6790, B => n6531, ZN => n6532);
   U10702 : XNOR2_X1 port map( A => n6533, B => n6532, ZN => n8085);
   U10703 : XNOR2_X1 port map( A => n6728, B => n6990, ZN => n6876);
   U10704 : XNOR2_X1 port map( A => n6534, B => n6876, ZN => n6538);
   U10705 : XNOR2_X1 port map( A => n7333, B => n6919, ZN => n6536);
   U10706 : XNOR2_X1 port map( A => n7336, B => n18396, ZN => n6535);
   U10707 : XNOR2_X1 port map( A => n6536, B => n6535, ZN => n6537);
   U10708 : XNOR2_X1 port map( A => n6538, B => n6537, ZN => n8086);
   U10709 : AOI22_X1 port map( A1 => n19826, A2 => n20254, B1 => n8085, B2 => 
                           n8086, ZN => n7556);
   U10710 : INV_X1 port map( A => n8087, ZN => n6539);
   U10711 : XNOR2_X1 port map( A => n6742, B => n7206, ZN => n6849);
   U10712 : XNOR2_X1 port map( A => n6767, B => n18997, ZN => n6540);
   U10713 : XNOR2_X1 port map( A => n6540, B => n6945, ZN => n6541);
   U10714 : XNOR2_X1 port map( A => n6541, B => n6849, ZN => n6544);
   U10715 : INV_X1 port map( A => n7308, ZN => n6542);
   U10716 : XNOR2_X1 port map( A => n7305, B => n6542, ZN => n6543);
   U10717 : XNOR2_X1 port map( A => n6545, B => n2382, ZN => n6547);
   U10718 : XNOR2_X1 port map( A => n6546, B => n6547, ZN => n6549);
   U10719 : XNOR2_X1 port map( A => n19778, B => n6736, ZN => n6879);
   U10720 : XNOR2_X1 port map( A => n6879, B => n6752, ZN => n6548);
   U10722 : INV_X1 port map( A => n8086, ZN => n8230);
   U10723 : OAI211_X1 port map( C1 => n20254, C2 => n8232, A => n20108, B => 
                           n8230, ZN => n6550);
   U10724 : XNOR2_X1 port map( A => n7201, B => n18084, ZN => n6551);
   U10725 : XNOR2_X1 port map( A => n7202, B => n6551, ZN => n6553);
   U10726 : XNOR2_X1 port map( A => n6552, B => n6553, ZN => n6556);
   U10727 : XNOR2_X1 port map( A => n7345, B => n6554, ZN => n6555);
   U10728 : XNOR2_X2 port map( A => n6556, B => n6555, ZN => n8241);
   U10729 : XNOR2_X1 port map( A => n6855, B => n7391, ZN => n6996);
   U10730 : XNOR2_X1 port map( A => n6557, B => n6996, ZN => n6561);
   U10731 : XNOR2_X1 port map( A => n6558, B => n347, ZN => n6559);
   U10732 : XNOR2_X1 port map( A => n7016, B => n6559, ZN => n6560);
   U10733 : XNOR2_X1 port map( A => n7116, B => n20203, ZN => n6563);
   U10734 : XNOR2_X1 port map( A => n6562, B => n6563, ZN => n6567);
   U10735 : XNOR2_X1 port map( A => n6819, B => n18208, ZN => n6564);
   U10736 : XNOR2_X1 port map( A => n6565, B => n6564, ZN => n6566);
   U10737 : XNOR2_X1 port map( A => n6567, B => n6566, ZN => n7862);
   U10738 : XNOR2_X1 port map( A => n6883, B => n7036, ZN => n6571);
   U10739 : XNOR2_X1 port map( A => n19764, B => n18433, ZN => n6569);
   U10740 : XNOR2_X1 port map( A => n6569, B => n6737, ZN => n6570);
   U10741 : XNOR2_X1 port map( A => n6570, B => n6571, ZN => n6578);
   U10742 : NOR2_X1 port map( A1 => n8239, A2 => n8100, ZN => n6572);
   U10743 : NAND2_X1 port map( A1 => n6572, A2 => n7862, ZN => n6586);
   U10744 : XNOR2_X1 port map( A => n7097, B => n6573, ZN => n6574);
   U10745 : XNOR2_X1 port map( A => n7040, B => n6574, ZN => n6577);
   U10746 : XNOR2_X1 port map( A => n7382, B => n6872, ZN => n6993);
   U10747 : XNOR2_X1 port map( A => n7188, B => n2280, ZN => n6575);
   U10748 : XNOR2_X1 port map( A => n6993, B => n6575, ZN => n6576);
   U10749 : XNOR2_X1 port map( A => n6577, B => n6576, ZN => n8098);
   U10750 : INV_X1 port map( A => n6578, ZN => n8099);
   U10751 : OAI21_X1 port map( B1 => n20493, B2 => n8238, A => n8099, ZN => 
                           n6585);
   U10752 : XNOR2_X1 port map( A => n6721, B => n6579, ZN => n6583);
   U10753 : XNOR2_X1 port map( A => n6839, B => n7091, ZN => n6581);
   U10754 : XNOR2_X1 port map( A => n7144, B => n19018, ZN => n6580);
   U10755 : XNOR2_X1 port map( A => n6581, B => n6580, ZN => n6582);
   U10756 : OAI21_X1 port map( B1 => n8112, B2 => n8111, A => n8239, ZN => 
                           n6584);
   U10757 : OAI21_X1 port map( B1 => n8628, B2 => n8713, A => n6587, ZN => 
                           n6655);
   U10758 : XNOR2_X1 port map( A => n6588, B => n6660, ZN => n6592);
   U10759 : XNOR2_X1 port map( A => n7288, B => n17535, ZN => n6589);
   U10760 : XNOR2_X1 port map( A => n6590, B => n6589, ZN => n6591);
   U10761 : XNOR2_X2 port map( A => n6592, B => n6591, ZN => n8095);
   U10762 : XNOR2_X1 port map( A => n6593, B => n6838, ZN => n6597);
   U10763 : XNOR2_X1 port map( A => n6680, B => n7318, ZN => n6595);
   U10764 : XNOR2_X1 port map( A => n7373, B => n1386, ZN => n6594);
   U10765 : XNOR2_X1 port map( A => n6595, B => n6594, ZN => n6596);
   U10766 : XNOR2_X1 port map( A => n6597, B => n6596, ZN => n8090);
   U10768 : XNOR2_X1 port map( A => n6810, B => n6598, ZN => n6601);
   U10769 : INV_X1 port map( A => n2369, ZN => n18503);
   U10770 : XNOR2_X1 port map( A => n7337, B => n18503, ZN => n6599);
   U10771 : XNOR2_X1 port map( A => n6689, B => n6599, ZN => n6600);
   U10772 : NAND2_X1 port map( A1 => n20511, A2 => n8211, ZN => n6618);
   U10773 : XNOR2_X1 port map( A => n883, B => n2307, ZN => n6602);
   U10774 : XOR2_X1 port map( A => n6801, B => n6602, Z => n6605);
   U10775 : XNOR2_X1 port map( A => n6672, B => n6603, ZN => n6604);
   U10776 : XNOR2_X1 port map( A => n6824, B => n6606, ZN => n6609);
   U10777 : XNOR2_X1 port map( A => n7298, B => n2954, ZN => n6607);
   U10778 : XNOR2_X1 port map( A => n6666, B => n6607, ZN => n6608);
   U10779 : NAND2_X1 port map( A1 => n8094, A2 => n8212, ZN => n7898);
   U10780 : OAI21_X1 port map( B1 => n8095, B2 => n8094, A => n7898, ZN => 
                           n6610);
   U10781 : XNOR2_X1 port map( A => n6611, B => n6612, ZN => n6616);
   U10782 : XNOR2_X1 port map( A => n7304, B => n7266, ZN => n6614);
   U10783 : XNOR2_X1 port map( A => n7006, B => n19102, ZN => n6613);
   U10784 : XNOR2_X1 port map( A => n6614, B => n6613, ZN => n6615);
   U10785 : XNOR2_X1 port map( A => n6616, B => n6615, ZN => n7631);
   U10786 : NAND3_X1 port map( A1 => n8095, A2 => n7631, A3 => n8209, ZN => 
                           n6617);
   U10787 : XNOR2_X1 port map( A => n6659, B => n6619, ZN => n6623);
   U10789 : INV_X1 port map( A => n8175, ZN => n8067);
   U10790 : XNOR2_X1 port map( A => n7212, B => n2233, ZN => n6624);
   U10791 : XNOR2_X1 port map( A => n6676, B => n6624, ZN => n6629);
   U10792 : INV_X1 port map( A => n6625, ZN => n6627);
   U10793 : XNOR2_X1 port map( A => n6627, B => n6626, ZN => n6628);
   U10794 : XNOR2_X1 port map( A => n7187, B => n538, ZN => n6631);
   U10795 : XNOR2_X1 port map( A => n20250, B => n6631, ZN => n6632);
   U10796 : NAND3_X1 port map( A1 => n8067, A2 => n8178, A3 => n8068, ZN => 
                           n6639);
   U10797 : XNOR2_X1 port map( A => n6633, B => n7178, ZN => n6636);
   U10798 : INV_X1 port map( A => n2385, ZN => n19123);
   U10799 : XNOR2_X1 port map( A => n6634, B => n19123, ZN => n6635);
   U10800 : XNOR2_X1 port map( A => n6636, B => n6635, ZN => n6637);
   U10801 : OR2_X1 port map( A1 => n19901, A2 => n8066, ZN => n7417);
   U10802 : NAND2_X1 port map( A1 => n6639, A2 => n7417, ZN => n6654);
   U10803 : XNOR2_X1 port map( A => n6665, B => n6640, ZN => n6645);
   U10804 : XNOR2_X1 port map( A => n6641, B => n7195, ZN => n6643);
   U10805 : XNOR2_X1 port map( A => n7296, B => n2337, ZN => n6642);
   U10806 : XNOR2_X1 port map( A => n6643, B => n6642, ZN => n6644);
   U10807 : XNOR2_X2 port map( A => n6645, B => n6644, ZN => n8179);
   U10808 : NAND2_X1 port map( A1 => n8068, A2 => n923, ZN => n6652);
   U10809 : INV_X1 port map( A => n6692, ZN => n6647);
   U10810 : XNOR2_X1 port map( A => n6647, B => n6646, ZN => n6651);
   U10811 : XNOR2_X1 port map( A => n7306, B => n6945, ZN => n6649);
   U10812 : XNOR2_X1 port map( A => n7006, B => n2079, ZN => n6648);
   U10813 : XNOR2_X1 port map( A => n6649, B => n6648, ZN => n6650);
   U10814 : XNOR2_X1 port map( A => n6651, B => n6650, ZN => n7621);
   U10815 : AOI21_X1 port map( B1 => n7887, B2 => n6652, A => n8069, ZN => 
                           n6653);
   U10817 : XNOR2_X1 port map( A => n6659, B => n6660, ZN => n6664);
   U10818 : XNOR2_X1 port map( A => n6661, B => n7081, ZN => n6760);
   U10819 : XNOR2_X1 port map( A => n7221, B => n18848, ZN => n6662);
   U10820 : XNOR2_X1 port map( A => n6760, B => n6662, ZN => n6663);
   U10821 : XNOR2_X2 port map( A => n6664, B => n6663, ZN => n8262);
   U10822 : INV_X1 port map( A => n6665, ZN => n6667);
   U10823 : XNOR2_X1 port map( A => n7065, B => n621, ZN => n6668);
   U10824 : XNOR2_X1 port map( A => n6669, B => n6668, ZN => n6670);
   U10825 : XNOR2_X1 port map( A => n7031, B => n15479, ZN => n6673);
   U10826 : XNOR2_X1 port map( A => n6672, B => n6673, ZN => n6678);
   U10827 : XNOR2_X1 port map( A => n6675, B => n6674, ZN => n6751);
   U10828 : XNOR2_X1 port map( A => n6751, B => n6676, ZN => n6677);
   U10829 : XNOR2_X1 port map( A => n6678, B => n6677, ZN => n7571);
   U10830 : INV_X1 port map( A => n7571, ZN => n8264);
   U10831 : XNOR2_X1 port map( A => n6679, B => n7087, ZN => n6794);
   U10832 : XNOR2_X1 port map( A => n7050, B => n18830, ZN => n6682);
   U10833 : XNOR2_X1 port map( A => n6680, B => n7373, ZN => n6681);
   U10834 : XNOR2_X1 port map( A => n6682, B => n6681, ZN => n6683);
   U10836 : XNOR2_X1 port map( A => n6686, B => n6685, ZN => n6691);
   U10837 : XNOR2_X1 port map( A => n6687, B => n19467, ZN => n6688);
   U10838 : XNOR2_X1 port map( A => n6689, B => n6688, ZN => n6690);
   U10839 : XNOR2_X1 port map( A => n6690, B => n6691, ZN => n8150);
   U10840 : NAND2_X1 port map( A1 => n8261, A2 => n8150, ZN => n6699);
   U10841 : XNOR2_X1 port map( A => n6692, B => n6770, ZN => n6697);
   U10842 : XNOR2_X1 port map( A => n6693, B => n7007, ZN => n6695);
   U10843 : XNOR2_X1 port map( A => n7267, B => n18308, ZN => n6694);
   U10844 : XNOR2_X1 port map( A => n6695, B => n6694, ZN => n6696);
   U10845 : XNOR2_X1 port map( A => n6697, B => n6696, ZN => n8153);
   U10846 : INV_X1 port map( A => n6702, ZN => n8246);
   U10847 : NOR2_X1 port map( A1 => n8253, A2 => n8246, ZN => n8252);
   U10849 : NAND3_X1 port map( A1 => n8253, A2 => n7560, A3 => n8251, ZN => 
                           n6705);
   U10850 : AND2_X1 port map( A1 => n9313, A2 => n9305, ZN => n6896);
   U10851 : INV_X1 port map( A => n941, ZN => n6706);
   U10852 : XNOR2_X1 port map( A => n19855, B => n6706, ZN => n6710);
   U10853 : XNOR2_X1 port map( A => n6708, B => n2323, ZN => n6709);
   U10854 : XNOR2_X1 port map( A => n6710, B => n6709, ZN => n6716);
   U10855 : INV_X1 port map( A => n6711, ZN => n6712);
   U10856 : XNOR2_X1 port map( A => n6712, B => n7391, ZN => n7194);
   U10857 : XNOR2_X1 port map( A => n6713, B => n6714, ZN => n7125);
   U10858 : XNOR2_X1 port map( A => n7194, B => n7125, ZN => n6715);
   U10859 : XNOR2_X1 port map( A => n6716, B => n6715, ZN => n6734);
   U10860 : XNOR2_X1 port map( A => n7122, B => n18716, ZN => n6720);
   U10861 : XNOR2_X1 port map( A => n6722, B => n6721, ZN => n6727);
   U10862 : XNOR2_X1 port map( A => n6724, B => n6723, ZN => n7148);
   U10863 : XNOR2_X1 port map( A => n7179, B => n2317, ZN => n6725);
   U10864 : XNOR2_X1 port map( A => n7148, B => n6725, ZN => n6726);
   U10865 : XNOR2_X1 port map( A => n6727, B => n6726, ZN => n7671);
   U10866 : INV_X1 port map( A => n7671, ZN => n8375);
   U10867 : XNOR2_X1 port map( A => n6729, B => n7184, ZN => n6731);
   U10868 : INV_X1 port map( A => n6734, ZN => n8377);
   U10870 : XNOR2_X1 port map( A => n6736, B => n6735, ZN => n7152);
   U10871 : XNOR2_X1 port map( A => n7152, B => n6737, ZN => n6741);
   U10872 : XNOR2_X1 port map( A => n6738, B => n19321, ZN => n6739);
   U10873 : XNOR2_X1 port map( A => n6754, B => n6165, ZN => n7060);
   U10874 : XNOR2_X1 port map( A => n6739, B => n7060, ZN => n6740);
   U10876 : XNOR2_X1 port map( A => n6743, B => n6742, ZN => n7162);
   U10877 : XNOR2_X1 port map( A => n6744, B => n7162, ZN => n6749);
   U10878 : XNOR2_X1 port map( A => n6768, B => n6745, ZN => n6747);
   U10879 : XNOR2_X1 port map( A => n7201, B => n2381, ZN => n6746);
   U10880 : XNOR2_X1 port map( A => n6747, B => n6746, ZN => n6748);
   U10881 : XNOR2_X1 port map( A => n6749, B => n6748, ZN => n7542);
   U10882 : NAND2_X1 port map( A1 => n7542, A2 => n6734, ZN => n8142);
   U10883 : INV_X1 port map( A => n6751, ZN => n6753);
   U10884 : XNOR2_X1 port map( A => n6753, B => n6752, ZN => n6758);
   U10885 : XNOR2_X1 port map( A => n7230, B => n7032, ZN => n6756);
   U10886 : XNOR2_X1 port map( A => n19850, B => n16366, ZN => n6755);
   U10887 : XNOR2_X1 port map( A => n6756, B => n6755, ZN => n6757);
   U10889 : XNOR2_X1 port map( A => n6759, B => n6760, ZN => n6765);
   U10890 : XNOR2_X1 port map( A => n6761, B => n7257, ZN => n6763);
   U10891 : XNOR2_X1 port map( A => n7026, B => n17466, ZN => n6762);
   U10892 : XNOR2_X1 port map( A => n6763, B => n6762, ZN => n6764);
   U10893 : XNOR2_X1 port map( A => n6765, B => n6764, ZN => n8380);
   U10894 : XNOR2_X1 port map( A => n179, B => n7263, ZN => n6766);
   U10895 : XNOR2_X1 port map( A => n7305, B => n6766, ZN => n6772);
   U10896 : XNOR2_X1 port map( A => n20225, B => n18075, ZN => n6769);
   U10897 : XNOR2_X1 port map( A => n6769, B => n6768, ZN => n6771);
   U10898 : MUX2_X1 port map( A => n8387, B => n163, S => n19925, Z => n6800);
   U10899 : INV_X1 port map( A => n6773, ZN => n6775);
   U10900 : XNOR2_X1 port map( A => n6775, B => n6774, ZN => n6781);
   U10901 : XNOR2_X1 port map( A => n941, B => n6776, ZN => n6779);
   U10902 : XNOR2_X1 port map( A => n6777, B => n573, ZN => n6778);
   U10903 : XNOR2_X1 port map( A => n6779, B => n6778, ZN => n6780);
   U10904 : INV_X1 port map( A => n7684, ZN => n8385);
   U10905 : XNOR2_X1 port map( A => n6782, B => n7332, ZN => n6785);
   U10906 : XNOR2_X1 port map( A => n6783, B => n7333, ZN => n6784);
   U10907 : XNOR2_X1 port map( A => n6784, B => n6785, ZN => n6789);
   U10908 : XNOR2_X1 port map( A => n7248, B => n16242, ZN => n6787);
   U10909 : XNOR2_X1 port map( A => n7098, B => n6787, ZN => n6788);
   U10910 : NAND3_X1 port map( A1 => n19925, A2 => n8387, A3 => n7497, ZN => 
                           n6799);
   U10911 : XNOR2_X1 port map( A => n7272, B => n17989, ZN => n6792);
   U10913 : XNOR2_X1 port map( A => n19852, B => n6792, ZN => n6798);
   U10914 : XNOR2_X1 port map( A => n7047, B => n6793, ZN => n6796);
   U10915 : INV_X1 port map( A => n6794, ZN => n6795);
   U10916 : XNOR2_X1 port map( A => n6795, B => n6796, ZN => n6797);
   U10918 : XNOR2_X1 port map( A => n6966, B => n7031, ZN => n6803);
   U10919 : INV_X1 port map( A => n6801, ZN => n6802);
   U10920 : XNOR2_X1 port map( A => n6802, B => n6803, ZN => n6807);
   U10921 : XNOR2_X1 port map( A => n7364, B => n19457, ZN => n6805);
   U10922 : XNOR2_X1 port map( A => n7363, B => n19840, ZN => n6804);
   U10923 : XNOR2_X1 port map( A => n6805, B => n6804, ZN => n6806);
   U10924 : XNOR2_X1 port map( A => n6808, B => n7042, ZN => n6809);
   U10925 : XNOR2_X1 port map( A => n6810, B => n6809, ZN => n6815);
   U10926 : XNOR2_X1 port map( A => n6918, B => n6811, ZN => n6813);
   U10927 : XNOR2_X1 port map( A => n943, B => n620, ZN => n6812);
   U10928 : XNOR2_X1 port map( A => n6813, B => n6812, ZN => n6814);
   U10929 : XNOR2_X1 port map( A => n6815, B => n6814, ZN => n6830);
   U10930 : INV_X1 port map( A => n7221, ZN => n6816);
   U10931 : XNOR2_X1 port map( A => n7355, B => n6816, ZN => n6817);
   U10932 : XNOR2_X1 port map( A => n6818, B => n6817, ZN => n6823);
   U10933 : XNOR2_X1 port map( A => n6977, B => n6819, ZN => n6821);
   U10934 : XNOR2_X1 port map( A => n7258, B => n2055, ZN => n6820);
   U10935 : XNOR2_X1 port map( A => n6821, B => n6820, ZN => n6822);
   U10936 : XNOR2_X1 port map( A => n7240, B => n6855, ZN => n6825);
   U10937 : XNOR2_X1 port map( A => n6824, B => n6825, ZN => n6829);
   U10938 : XNOR2_X1 port map( A => n7392, B => n7390, ZN => n6827);
   U10939 : XNOR2_X1 port map( A => n7018, B => n457, ZN => n6826);
   U10940 : XOR2_X1 port map( A => n6827, B => n6826, Z => n6828);
   U10941 : NAND2_X1 port map( A1 => n7852, A2 => n282, ZN => n6831);
   U10942 : XNOR2_X1 port map( A => n6832, B => n7345, ZN => n6834);
   U10943 : XNOR2_X1 port map( A => n6946, B => n7007, ZN => n6833);
   U10944 : XNOR2_X1 port map( A => n6834, B => n6833, ZN => n6836);
   U10945 : XNOR2_X1 port map( A => n6836, B => n6835, ZN => n8162);
   U10946 : INV_X1 port map( A => n8162, ZN => n7856);
   U10947 : INV_X1 port map( A => n8159, ZN => n7851);
   U10948 : NAND3_X1 port map( A1 => n7856, A2 => n7724, A3 => n7851, ZN => 
                           n6846);
   U10949 : INV_X1 port map( A => n6838, ZN => n6841);
   U10950 : XNOR2_X1 port map( A => n7274, B => n6839, ZN => n6840);
   U10951 : XNOR2_X1 port map( A => n7050, B => n18801, ZN => n6843);
   U10952 : XNOR2_X1 port map( A => n6985, B => n7046, ZN => n6842);
   U10953 : INV_X1 port map( A => n8157, ZN => n6844);
   U10954 : OAI21_X1 port map( B1 => n1751, B2 => n20011, A => n8824, ZN => 
                           n6895);
   U10955 : INV_X1 port map( A => n16424, ZN => n18792);
   U10956 : XNOR2_X1 port map( A => n6849, B => n6848, ZN => n6853);
   U10957 : XNOR2_X1 port map( A => n6850, B => n7264, ZN => n7350);
   U10958 : XNOR2_X1 port map( A => n7202, B => n7304, ZN => n6851);
   U10959 : XNOR2_X1 port map( A => n7350, B => n6851, ZN => n6852);
   U10960 : XNOR2_X1 port map( A => n6853, B => n6852, ZN => n8350);
   U10961 : XNOR2_X1 port map( A => n6855, B => n6854, ZN => n6857);
   U10962 : INV_X1 port map( A => n6858, ZN => n6860);
   U10963 : XNOR2_X1 port map( A => n7013, B => n2275, ZN => n6859);
   U10964 : XNOR2_X1 port map( A => n6860, B => n6859, ZN => n6861);
   U10967 : NAND2_X1 port map( A1 => n8350, A2 => n8140, ZN => n7722);
   U10968 : INV_X1 port map( A => n7122, ZN => n6863);
   U10969 : XNOR2_X1 port map( A => n20203, B => n6863, ZN => n6866);
   U10971 : XNOR2_X1 port map( A => n19741, B => n6866, ZN => n6870);
   U10972 : XNOR2_X1 port map( A => n6819, B => n7218, ZN => n6976);
   U10973 : XNOR2_X1 port map( A => n19730, B => n17787, ZN => n6868);
   U10974 : XNOR2_X1 port map( A => n6976, B => n6868, ZN => n6869);
   U10976 : XNOR2_X1 port map( A => n6874, B => n6873, ZN => n6875);
   U10977 : XNOR2_X1 port map( A => n6875, B => n6876, ZN => n6878);
   U10978 : XNOR2_X1 port map( A => n6878, B => n6877, ZN => n8348);
   U10980 : NAND2_X1 port map( A1 => n19914, A2 => n8272, ZN => n6886);
   U10981 : INV_X1 port map( A => n6879, ZN => n6880);
   U10982 : XNOR2_X1 port map( A => n6880, B => n6881, ZN => n6885);
   U10983 : XNOR2_X1 port map( A => n7365, B => n2298, ZN => n6882);
   U10984 : XNOR2_X1 port map( A => n6883, B => n6882, ZN => n6884);
   U10985 : OAI211_X1 port map( C1 => n8352, C2 => n8272, A => n6886, B => 
                           n8349, ZN => n6894);
   U10986 : INV_X1 port map( A => n6887, ZN => n6888);
   U10987 : XNOR2_X1 port map( A => n6888, B => n6889, ZN => n6893);
   U10988 : XNOR2_X1 port map( A => n7144, B => n18278, ZN => n6890);
   U10989 : XNOR2_X1 port map( A => n6891, B => n6890, ZN => n6892);
   U10990 : INV_X1 port map( A => n20200, ZN => n8141);
   U10991 : MUX2_X1 port map( A => n6896, B => n6895, S => n9228, Z => n6898);
   U10992 : INV_X1 port map( A => n9307, ZN => n9309);
   U10993 : AND3_X1 port map( A1 => n20011, A2 => n9309, A3 => n9053, ZN => 
                           n6897);
   U10996 : NOR2_X1 port map( A1 => n7500, A2 => n7739, ZN => n6900);
   U10997 : OAI211_X1 port map( C1 => n7931, C2 => n20360, A => n1063, B => 
                           n20195, ZN => n6903);
   U10998 : INV_X1 port map( A => n9162, ZN => n8696);
   U10999 : NAND2_X1 port map( A1 => n7904, A2 => n7908, ZN => n6905);
   U11001 : INV_X1 port map( A => n20166, ZN => n7755);
   U11002 : NOR2_X1 port map( A1 => n7914, A2 => n7750, ZN => n6907);
   U11003 : NOR2_X1 port map( A1 => n7748, A2 => n7507, ZN => n6906);
   U11004 : MUX2_X1 port map( A => n6907, B => n6906, S => n7749, Z => n6910);
   U11005 : XNOR2_X1 port map( A => n7228, B => n6911, ZN => n6916);
   U11006 : XNOR2_X1 port map( A => n7326, B => n7363, ZN => n6914);
   U11007 : XNOR2_X1 port map( A => n6912, B => n2356, ZN => n6913);
   U11008 : XNOR2_X1 port map( A => n6914, B => n6913, ZN => n6915);
   U11009 : XNOR2_X1 port map( A => n7338, B => Key(60), ZN => n6920);
   U11010 : XNOR2_X1 port map( A => n6920, B => n20250, ZN => n6921);
   U11011 : XNOR2_X1 port map( A => n7380, B => n6921, ZN => n6924);
   U11012 : XNOR2_X1 port map( A => n7248, B => n943, ZN => n6922);
   U11013 : XNOR2_X1 port map( A => n6922, B => n7134, ZN => n6923);
   U11014 : XNOR2_X1 port map( A => n6924, B => n6923, ZN => n7728);
   U11015 : XNOR2_X1 port map( A => n6926, B => n6925, ZN => n6930);
   U11016 : XNOR2_X1 port map( A => n6927, B => n7046, ZN => n7376);
   U11017 : XNOR2_X1 port map( A => n7316, B => n18146, ZN => n6928);
   U11018 : XNOR2_X1 port map( A => n7376, B => n6928, ZN => n6929);
   U11020 : XNOR2_X1 port map( A => n5884, B => n7355, ZN => n6931);
   U11021 : XNOR2_X1 port map( A => n6931, B => n7256, ZN => n6934);
   U11022 : XNOR2_X1 port map( A => n7258, B => n7121, ZN => n6933);
   U11023 : XNOR2_X1 port map( A => n6935, B => n7238, ZN => n6940);
   U11024 : XNOR2_X1 port map( A => n7390, B => n7296, ZN => n6938);
   U11025 : INV_X1 port map( A => n20064, ZN => n17683);
   U11026 : XNOR2_X1 port map( A => n6936, B => n17683, ZN => n6937);
   U11027 : XNOR2_X1 port map( A => n6938, B => n6937, ZN => n6939);
   U11028 : XNOR2_X1 port map( A => n6940, B => n6939, ZN => n7493);
   U11029 : OAI22_X1 port map( A1 => n8166, A2 => n7679, B1 => n8165, B2 => 
                           n7728, ZN => n7729);
   U11030 : INV_X1 port map( A => n17024, ZN => n18670);
   U11031 : XNOR2_X1 port map( A => n7160, B => n18670, ZN => n6941);
   U11032 : XNOR2_X1 port map( A => n7345, B => n6941, ZN => n6944);
   U11033 : XNOR2_X1 port map( A => n6942, B => n7306, ZN => n6943);
   U11034 : XNOR2_X1 port map( A => n6944, B => n6943, ZN => n6949);
   U11035 : XNOR2_X1 port map( A => n6948, B => n6947, ZN => n7270);
   U11036 : NAND2_X1 port map( A1 => n7729, A2 => n8341, ZN => n6950);
   U11037 : NAND2_X1 port map( A1 => n6951, A2 => n7673, ZN => n7711);
   U11038 : NAND2_X1 port map( A1 => n6952, A2 => n8365, ZN => n6957);
   U11039 : INV_X1 port map( A => n7673, ZN => n6953);
   U11040 : NAND2_X1 port map( A1 => n7709, A2 => n6953, ZN => n6954);
   U11041 : NAND3_X1 port map( A1 => n7711, A2 => n7675, A3 => n6954, ZN => 
                           n6956);
   U11042 : INV_X1 port map( A => n7675, ZN => n8366);
   U11043 : INV_X1 port map( A => n8365, ZN => n8363);
   U11044 : NAND3_X1 port map( A1 => n1994, A2 => n8363, A3 => n7674, ZN => 
                           n6955);
   U11045 : INV_X1 port map( A => n9163, ZN => n9161);
   U11046 : NAND3_X1 port map( A1 => n8611, A2 => n8609, A3 => n9161, ZN => 
                           n6959);
   U11047 : NAND3_X1 port map( A1 => n9164, A2 => n9158, A3 => n1230, ZN => 
                           n6958);
   U11048 : XNOR2_X1 port map( A => n6961, B => n6960, ZN => n6965);
   U11049 : XNOR2_X1 port map( A => n7009, B => n18439, ZN => n6963);
   U11050 : XNOR2_X1 port map( A => n6963, B => n6962, ZN => n6964);
   U11052 : XNOR2_X1 port map( A => n6966, B => n6967, ZN => n6969);
   U11053 : XNOR2_X1 port map( A => n7151, B => n7032, ZN => n6968);
   U11054 : XNOR2_X1 port map( A => n6969, B => n6968, ZN => n6974);
   U11055 : XNOR2_X1 port map( A => n6970, B => n7364, ZN => n6972);
   U11056 : XNOR2_X1 port map( A => n883, B => n18065, ZN => n6971);
   U11057 : XNOR2_X1 port map( A => n6972, B => n6971, ZN => n6973);
   U11058 : XNOR2_X2 port map( A => n6974, B => n6973, ZN => n7967);
   U11059 : XNOR2_X1 port map( A => n7354, B => n7288, ZN => n6975);
   U11060 : XNOR2_X1 port map( A => n20209, B => n6975, ZN => n6981);
   U11061 : XNOR2_X1 port map( A => n6977, B => n20227, ZN => n6979);
   U11062 : XNOR2_X1 port map( A => n7026, B => n16487, ZN => n6978);
   U11063 : XNOR2_X1 port map( A => n6979, B => n6978, ZN => n6980);
   U11064 : XNOR2_X1 port map( A => n6981, B => n6980, ZN => n7487);
   U11065 : XNOR2_X1 port map( A => n6982, B => n7047, ZN => n6984);
   U11066 : XNOR2_X1 port map( A => n903, B => n6839, ZN => n6983);
   U11067 : XNOR2_X1 port map( A => n6984, B => n6983, ZN => n6989);
   U11068 : XNOR2_X1 port map( A => n7146, B => n7318, ZN => n6987);
   U11069 : XNOR2_X1 port map( A => n6985, B => n18420, ZN => n6986);
   U11070 : XNOR2_X1 port map( A => n6987, B => n6986, ZN => n6988);
   U11071 : XNOR2_X1 port map( A => n6989, B => n6988, ZN => n7971);
   U11072 : XNOR2_X1 port map( A => n6990, B => n19027, ZN => n6991);
   U11073 : XNOR2_X1 port map( A => n6993, B => n7134, ZN => n6994);
   U11074 : XNOR2_X1 port map( A => n6995, B => n6996, ZN => n7001);
   U11075 : XNOR2_X1 port map( A => n7017, B => n2417, ZN => n6999);
   U11076 : XNOR2_X1 port map( A => n6997, B => n7128, ZN => n6998);
   U11077 : XNOR2_X1 port map( A => n6999, B => n6998, ZN => n7000);
   U11078 : INV_X1 port map( A => n8527, ZN => n8849);
   U11079 : INV_X1 port map( A => n7002, ZN => n7753);
   U11080 : INV_X1 port map( A => n9046, ZN => n8852);
   U11081 : XNOR2_X1 port map( A => n7201, B => n17733, ZN => n7005);
   U11082 : XNOR2_X1 port map( A => n7005, B => n7264, ZN => n7008);
   U11083 : XNOR2_X1 port map( A => n7006, B => n7007, ZN => n7204);
   U11084 : XNOR2_X1 port map( A => n7008, B => n7204, ZN => n7012);
   U11085 : XNOR2_X1 port map( A => n179, B => n7267, ZN => n7010);
   U11086 : XNOR2_X1 port map( A => n7010, B => n7345, ZN => n7011);
   U11087 : INV_X1 port map( A => n20165, ZN => n7915);
   U11088 : INV_X1 port map( A => n7013, ZN => n7015);
   U11089 : XNOR2_X1 port map( A => n7015, B => n7014, ZN => n7237);
   U11090 : XNOR2_X1 port map( A => n7016, B => n7237, ZN => n7022);
   U11091 : XNOR2_X1 port map( A => n7017, B => n1869, ZN => n7020);
   U11092 : XNOR2_X1 port map( A => n7195, B => n7018, ZN => n7019);
   U11093 : XNOR2_X1 port map( A => n7020, B => n7019, ZN => n7021);
   U11094 : XNOR2_X2 port map( A => n7022, B => n7021, ZN => n8910);
   U11095 : INV_X1 port map( A => n8910, ZN => n8906);
   U11096 : XNOR2_X1 port map( A => n7355, B => n7216, ZN => n7024);
   U11097 : XNOR2_X1 port map( A => n7253, B => n7221, ZN => n7023);
   U11098 : XNOR2_X1 port map( A => n7024, B => n7023, ZN => n7030);
   U11099 : XNOR2_X1 port map( A => n7026, B => n7025, ZN => n7028);
   U11100 : XNOR2_X1 port map( A => n7028, B => n7027, ZN => n7029);
   U11102 : INV_X1 port map( A => n7836, ZN => n7961);
   U11103 : XNOR2_X1 port map( A => n7212, B => n7031, ZN => n7034);
   U11104 : XNOR2_X1 port map( A => n7032, B => n2384, ZN => n7033);
   U11105 : XNOR2_X1 port map( A => n7034, B => n7033, ZN => n7038);
   U11106 : XNOR2_X1 port map( A => n7036, B => n7229, ZN => n7037);
   U11108 : XNOR2_X1 port map( A => n19944, B => n7333, ZN => n7039);
   U11109 : XNOR2_X1 port map( A => n7040, B => n7039, ZN => n7045);
   U11110 : XNOR2_X1 port map( A => n7041, B => n7383, ZN => n7246);
   U11111 : XNOR2_X1 port map( A => n7042, B => n642, ZN => n7043);
   U11112 : XNOR2_X1 port map( A => n7246, B => n7043, ZN => n7044);
   U11113 : XNOR2_X1 port map( A => n7045, B => n7044, ZN => n7956);
   U11114 : XNOR2_X1 port map( A => n7046, B => n7047, ZN => n7049);
   U11115 : XNOR2_X1 port map( A => n7048, B => n7371, ZN => n7277);
   U11116 : XNOR2_X1 port map( A => n7277, B => n7049, ZN => n7054);
   U11117 : XNOR2_X1 port map( A => n7050, B => n7178, ZN => n7052);
   U11118 : XNOR2_X1 port map( A => n7179, B => n2448, ZN => n7051);
   U11119 : XNOR2_X1 port map( A => n7052, B => n7051, ZN => n7053);
   U11120 : INV_X1 port map( A => n7958, ZN => n7835);
   U11121 : NAND3_X1 port map( A1 => n277, A2 => n7835, A3 => n8910, ZN => 
                           n7055);
   U11122 : XNOR2_X1 port map( A => n7057, B => n7058, ZN => n7062);
   U11123 : XNOR2_X1 port map( A => n7154, B => n18887, ZN => n7059);
   U11124 : XNOR2_X1 port map( A => n7060, B => n7059, ZN => n7061);
   U11125 : XNOR2_X1 port map( A => n7062, B => n7061, ZN => n7096);
   U11126 : INV_X1 port map( A => n7096, ZN => n7830);
   U11127 : XNOR2_X1 port map( A => n7127, B => n7241, ZN => n7063);
   U11128 : XNOR2_X1 port map( A => n7064, B => n7063, ZN => n7069);
   U11129 : XNOR2_X1 port map( A => n7065, B => n2203, ZN => n7067);
   U11130 : XNOR2_X1 port map( A => n7066, B => n7067, ZN => n7068);
   U11131 : XNOR2_X1 port map( A => n7070, B => n17365, ZN => n7072);
   U11132 : XNOR2_X1 port map( A => n7164, B => n7266, ZN => n7071);
   U11133 : XNOR2_X1 port map( A => n7072, B => n7071, ZN => n7076);
   U11134 : XNOR2_X1 port map( A => n7074, B => n7073, ZN => n7075);
   U11135 : XNOR2_X1 port map( A => n7078, B => n7079, ZN => n7085);
   U11136 : XNOR2_X1 port map( A => n7118, B => n7080, ZN => n7083);
   U11137 : XNOR2_X1 port map( A => n7081, B => n2413, ZN => n7082);
   U11138 : XNOR2_X1 port map( A => n7083, B => n7082, ZN => n7084);
   U11139 : NAND2_X1 port map( A1 => n8014, A2 => n7086, ZN => n7106);
   U11140 : XNOR2_X1 port map( A => n7087, B => n7088, ZN => n7090);
   U11141 : XNOR2_X1 port map( A => n7090, B => n7089, ZN => n7095);
   U11142 : XNOR2_X1 port map( A => n7273, B => n7316, ZN => n7093);
   U11143 : XNOR2_X1 port map( A => n7091, B => n18366, ZN => n7092);
   U11144 : XNOR2_X1 port map( A => n7093, B => n7092, ZN => n7094);
   U11145 : XNOR2_X1 port map( A => n7095, B => n7094, ZN => n8011);
   U11146 : NAND2_X1 port map( A1 => n7830, A2 => n8012, ZN => n7105);
   U11147 : XNOR2_X1 port map( A => n7097, B => n19780, ZN => n7099);
   U11148 : XNOR2_X1 port map( A => n7098, B => n7099, ZN => n7103);
   U11149 : XNOR2_X1 port map( A => n7249, B => n7336, ZN => n7101);
   U11150 : XNOR2_X1 port map( A => n7338, B => n2164, ZN => n7100);
   U11151 : XNOR2_X1 port map( A => n7101, B => n7100, ZN => n7102);
   U11152 : XNOR2_X1 port map( A => n7103, B => n7102, ZN => n7990);
   U11153 : INV_X1 port map( A => n7990, ZN => n7829);
   U11154 : NAND3_X1 port map( A1 => n7096, A2 => n7829, A3 => n8015, ZN => 
                           n7104);
   U11155 : INV_X1 port map( A => n8851, ZN => n7656);
   U11156 : NAND2_X1 port map( A1 => n7919, A2 => n7768, ZN => n7113);
   U11157 : INV_X1 port map( A => n7984, ZN => n7534);
   U11158 : NAND2_X1 port map( A1 => n7534, A2 => n7981, ZN => n7108);
   U11159 : NAND3_X1 port map( A1 => n7110, A2 => n19812, A3 => n7108, ZN => 
                           n7112);
   U11160 : NAND3_X1 port map( A1 => n505, A2 => n7921, A3 => n7984, ZN => 
                           n7111);
   U11161 : OAI211_X1 port map( C1 => n7978, C2 => n7113, A => n7112, B => 
                           n7111, ZN => n8848);
   U11162 : INV_X1 port map( A => n8848, ZN => n7659);
   U11163 : NOR2_X1 port map( A1 => n9046, A2 => n7659, ZN => n7114);
   U11164 : NAND2_X1 port map( A1 => n7114, A2 => n8849, ZN => n7173);
   U11165 : XNOR2_X1 port map( A => n6478, B => n2394, ZN => n7117);
   U11167 : XNOR2_X1 port map( A => n7118, B => n1053, ZN => n7119);
   U11168 : XNOR2_X1 port map( A => n7122, B => n20227, ZN => n7123);
   U11169 : XNOR2_X1 port map( A => n7126, B => n7125, ZN => n7132);
   U11170 : XNOR2_X1 port map( A => n7127, B => n19953, ZN => n7130);
   U11171 : XNOR2_X1 port map( A => n7128, B => n1782, ZN => n7129);
   U11172 : XNOR2_X1 port map( A => n7130, B => n7129, ZN => n7131);
   U11173 : XNOR2_X1 port map( A => n899, B => n7134, ZN => n7136);
   U11174 : XNOR2_X1 port map( A => n7136, B => n7135, ZN => n7141);
   U11175 : XNOR2_X1 port map( A => n6728, B => n2442, ZN => n7139);
   U11176 : XNOR2_X1 port map( A => n7137, B => n7332, ZN => n7138);
   U11177 : XNOR2_X1 port map( A => n7139, B => n7138, ZN => n7140);
   U11178 : XNOR2_X1 port map( A => n7141, B => n7140, ZN => n7952);
   U11179 : XNOR2_X1 port map( A => n7143, B => n7142, ZN => n7145);
   U11180 : XNOR2_X1 port map( A => n7317, B => n7144, ZN => n7176);
   U11181 : XNOR2_X1 port map( A => n7176, B => n7145, ZN => n7150);
   U11182 : XNOR2_X1 port map( A => n7146, B => n18078, ZN => n7147);
   U11183 : XNOR2_X1 port map( A => n7148, B => n7147, ZN => n7149);
   U11184 : XNOR2_X1 port map( A => n7149, B => n7150, ZN => n7951);
   U11185 : XNOR2_X1 port map( A => n7151, B => n7211, ZN => n7153);
   U11186 : XNOR2_X1 port map( A => n7152, B => n7153, ZN => n7159);
   U11187 : XNOR2_X1 port map( A => n19699, B => n7154, ZN => n7157);
   U11188 : XNOR2_X1 port map( A => n7155, B => n18988, ZN => n7156);
   U11189 : XNOR2_X1 port map( A => n7157, B => n7156, ZN => n7158);
   U11190 : XNOR2_X1 port map( A => n7159, B => n7158, ZN => n7481);
   U11191 : INV_X1 port map( A => n7481, ZN => n7950);
   U11193 : INV_X1 port map( A => n7814, ZN => n7169);
   U11194 : XNOR2_X1 port map( A => n7160, B => n311, ZN => n7161);
   U11195 : XNOR2_X1 port map( A => n7164, B => n7163, ZN => n7165);
   U11196 : XNOR2_X1 port map( A => n7305, B => n7165, ZN => n7166);
   U11197 : XNOR2_X2 port map( A => n7167, B => n7166, ZN => n7948);
   U11198 : NAND2_X1 port map( A1 => n7169, A2 => n7168, ZN => n7171);
   U11199 : INV_X1 port map( A => n7818, ZN => n7170);
   U11201 : INV_X1 port map( A => n9039, ZN => n8529);
   U11202 : NAND3_X1 port map( A1 => n8529, A2 => n8527, A3 => n7656, ZN => 
                           n7172);
   U11203 : NAND2_X1 port map( A1 => n7173, A2 => n7172, ZN => n7174);
   U11204 : XNOR2_X1 port map( A => n7177, B => n7176, ZN => n7183);
   U11205 : XNOR2_X1 port map( A => n903, B => n7178, ZN => n7181);
   U11206 : XNOR2_X1 port map( A => n7179, B => n19336, ZN => n7180);
   U11207 : XNOR2_X1 port map( A => n7181, B => n7180, ZN => n7182);
   U11208 : XNOR2_X1 port map( A => n7183, B => n7182, ZN => n7475);
   U11209 : XNOR2_X1 port map( A => n7332, B => n7184, ZN => n7186);
   U11210 : XNOR2_X1 port map( A => n7186, B => n7185, ZN => n7192);
   U11211 : XNOR2_X1 port map( A => n19944, B => n7382, ZN => n7190);
   U11212 : XNOR2_X1 port map( A => n7188, B => n18779, ZN => n7189);
   U11213 : XNOR2_X1 port map( A => n7190, B => n7189, ZN => n7191);
   U11215 : INV_X1 port map( A => n8315, ZN => n8003);
   U11216 : INV_X1 port map( A => n7594, ZN => n7227);
   U11217 : XNOR2_X1 port map( A => n7193, B => n7194, ZN => n7200);
   U11218 : XNOR2_X1 port map( A => n7195, B => n19953, ZN => n7198);
   U11219 : XNOR2_X1 port map( A => n7196, B => n2329, ZN => n7197);
   U11220 : XNOR2_X1 port map( A => n7198, B => n7197, ZN => n7199);
   U11222 : XNOR2_X1 port map( A => n7201, B => n16030, ZN => n7203);
   U11223 : XNOR2_X1 port map( A => n7203, B => n7202, ZN => n7205);
   U11224 : XNOR2_X1 port map( A => n7205, B => n7204, ZN => n7209);
   U11225 : XNOR2_X1 port map( A => n7348, B => n7206, ZN => n7207);
   U11226 : XNOR2_X1 port map( A => n7305, B => n7207, ZN => n7208);
   U11227 : XNOR2_X1 port map( A => n7209, B => n7208, ZN => n7591);
   U11228 : XNOR2_X1 port map( A => n7212, B => n7211, ZN => n7213);
   U11229 : OAI211_X1 port map( C1 => n7592, C2 => n8313, A => n8004, B => 
                           n8315, ZN => n7226);
   U11230 : XNOR2_X1 port map( A => n7217, B => n7216, ZN => n7220);
   U11231 : XNOR2_X1 port map( A => n7218, B => n7354, ZN => n7219);
   U11232 : XNOR2_X1 port map( A => n7220, B => n7219, ZN => n7224);
   U11233 : XNOR2_X1 port map( A => n1052, B => n7221, ZN => n7222);
   U11234 : XNOR2_X1 port map( A => n20203, B => n7222, ZN => n7223);
   U11235 : XNOR2_X1 port map( A => n7224, B => n7223, ZN => n8316);
   U11237 : NAND2_X1 port map( A1 => n19520, A2 => n8313, ZN => n7225);
   U11238 : XNOR2_X1 port map( A => n7228, B => n7229, ZN => n7236);
   U11239 : XNOR2_X1 port map( A => n7230, B => n18854, ZN => n7234);
   U11240 : XNOR2_X1 port map( A => n19841, B => n7232, ZN => n7233);
   U11241 : XNOR2_X1 port map( A => n7234, B => n7233, ZN => n7235);
   U11242 : INV_X1 port map( A => n7237, ZN => n7239);
   U11243 : XNOR2_X1 port map( A => n7239, B => n7238, ZN => n7245);
   U11244 : XNOR2_X1 port map( A => n7240, B => n7241, ZN => n7243);
   U11245 : XNOR2_X1 port map( A => n6777, B => n18055, ZN => n7242);
   U11246 : XNOR2_X1 port map( A => n7243, B => n7242, ZN => n7244);
   U11247 : XNOR2_X1 port map( A => n7249, B => n7248, ZN => n7251);
   U11248 : XNOR2_X1 port map( A => n6249, B => n2108, ZN => n7250);
   U11249 : XNOR2_X1 port map( A => n7251, B => n7250, ZN => n7252);
   U11250 : XNOR2_X1 port map( A => n7254, B => n7253, ZN => n7255);
   U11251 : XNOR2_X1 port map( A => n7256, B => n7255, ZN => n7262);
   U11252 : XNOR2_X1 port map( A => n7025, B => n7257, ZN => n7260);
   U11253 : XNOR2_X1 port map( A => n7258, B => n2032, ZN => n7259);
   U11254 : XNOR2_X1 port map( A => n7260, B => n7259, ZN => n7261);
   U11255 : XNOR2_X1 port map( A => n7261, B => n7262, ZN => n7466);
   U11256 : INV_X1 port map( A => n7963, ZN => n7283);
   U11257 : INV_X1 port map( A => n2192, ZN => n17940);
   U11258 : XNOR2_X1 port map( A => n7263, B => n17940, ZN => n7265);
   U11259 : XNOR2_X1 port map( A => n7265, B => n7264, ZN => n7269);
   U11260 : XNOR2_X1 port map( A => n7266, B => n7267, ZN => n7268);
   U11261 : XNOR2_X1 port map( A => n7269, B => n7268, ZN => n7271);
   U11262 : XNOR2_X1 port map( A => n7271, B => n7270, ZN => n7965);
   U11263 : INV_X1 port map( A => n7965, ZN => n8018);
   U11264 : XNOR2_X1 port map( A => n7272, B => n17095, ZN => n7276);
   U11265 : XNOR2_X1 port map( A => n7273, B => n7274, ZN => n7275);
   U11266 : XNOR2_X1 port map( A => n7276, B => n7275, ZN => n7281);
   U11267 : INV_X1 port map( A => n7277, ZN => n7278);
   U11268 : XNOR2_X1 port map( A => n7279, B => n7278, ZN => n7280);
   U11271 : NOR2_X1 port map( A1 => n20347, A2 => n20490, ZN => n7282);
   U11272 : AOI22_X1 port map( A1 => n7283, A2 => n8018, B1 => n208, B2 => 
                           n7282, ZN => n7284);
   U11273 : XNOR2_X1 port map( A => n1052, B => n7288, ZN => n7291);
   U11274 : XNOR2_X1 port map( A => n7289, B => n2310, ZN => n7290);
   U11275 : XNOR2_X1 port map( A => n7291, B => n7290, ZN => n7292);
   U11276 : XNOR2_X1 port map( A => n7295, B => n7294, ZN => n7302);
   U11277 : XNOR2_X1 port map( A => n7296, B => n19953, ZN => n7300);
   U11278 : XNOR2_X1 port map( A => n7298, B => n18768, ZN => n7299);
   U11279 : XNOR2_X1 port map( A => n7300, B => n7299, ZN => n7301);
   U11280 : XNOR2_X1 port map( A => n7302, B => n7301, ZN => n7312);
   U11281 : NAND2_X1 port map( A1 => n1425, A2 => n7312, ZN => n7343);
   U11282 : XNOR2_X1 port map( A => n7306, B => n17544, ZN => n7307);
   U11283 : XNOR2_X1 port map( A => n7308, B => n7307, ZN => n7309);
   U11284 : XNOR2_X1 port map( A => n7310, B => n7309, ZN => n7311);
   U11285 : INV_X1 port map( A => n7312, ZN => n8001);
   U11286 : INV_X1 port map( A => n7313, ZN => n7314);
   U11287 : XNOR2_X1 port map( A => n7314, B => n7315, ZN => n7322);
   U11288 : XNOR2_X1 port map( A => n7317, B => n7316, ZN => n7320);
   U11289 : XNOR2_X1 port map( A => n7318, B => n345, ZN => n7319);
   U11290 : XNOR2_X1 port map( A => n7320, B => n7319, ZN => n7321);
   U11291 : XNOR2_X1 port map( A => n7323, B => n7324, ZN => n7331);
   U11292 : XNOR2_X1 port map( A => n883, B => n18726, ZN => n7329);
   U11293 : XNOR2_X1 port map( A => n7326, B => n19698, ZN => n7328);
   U11294 : XNOR2_X1 port map( A => n7328, B => n7329, ZN => n7330);
   U11295 : XNOR2_X1 port map( A => n7331, B => n7330, ZN => n7585);
   U11296 : XNOR2_X1 port map( A => n7332, B => n7333, ZN => n7335);
   U11297 : XNOR2_X1 port map( A => n7335, B => n7334, ZN => n7342);
   U11298 : XNOR2_X1 port map( A => n7337, B => n7336, ZN => n7340);
   U11299 : XNOR2_X1 port map( A => n7338, B => n17804, ZN => n7339);
   U11300 : XNOR2_X1 port map( A => n7340, B => n7339, ZN => n7341);
   U11301 : MUX2_X1 port map( A => n8925, B => n8932, S => n8928, Z => n7413);
   U11302 : XNOR2_X1 port map( A => n7345, B => n7344, ZN => n7347);
   U11303 : XNOR2_X1 port map( A => n7346, B => n7347, ZN => n7351);
   U11304 : XNOR2_X1 port map( A => n7348, B => n18070, ZN => n7349);
   U11305 : XNOR2_X1 port map( A => n7025, B => n2383, ZN => n7352);
   U11306 : XNOR2_X1 port map( A => n7352, B => n7353, ZN => n7359);
   U11307 : XNOR2_X1 port map( A => n7355, B => n7354, ZN => n7357);
   U11308 : XNOR2_X1 port map( A => n7357, B => n7356, ZN => n7358);
   U11309 : XNOR2_X1 port map( A => n7359, B => n7358, ZN => n8025);
   U11310 : XNOR2_X1 port map( A => n7361, B => n7362, ZN => n7369);
   U11311 : XNOR2_X1 port map( A => n7364, B => n7363, ZN => n7367);
   U11312 : XNOR2_X1 port map( A => n7365, B => n17993, ZN => n7366);
   U11313 : XNOR2_X1 port map( A => n7367, B => n7366, ZN => n7368);
   U11314 : XNOR2_X1 port map( A => n7368, B => n7369, ZN => n7389);
   U11315 : INV_X1 port map( A => n7389, ZN => n8290);
   U11316 : OAI21_X1 port map( B1 => n8293, B2 => n20189, A => n7370, ZN => 
                           n7401);
   U11317 : XNOR2_X1 port map( A => n7371, B => n903, ZN => n7375);
   U11318 : XNOR2_X1 port map( A => n7373, B => n19436, ZN => n7374);
   U11319 : XNOR2_X1 port map( A => n7375, B => n7374, ZN => n7379);
   U11320 : XNOR2_X1 port map( A => n7377, B => n7376, ZN => n7378);
   U11321 : XNOR2_X1 port map( A => n7378, B => n7379, ZN => n8288);
   U11322 : XNOR2_X1 port map( A => n7382, B => n7383, ZN => n7386);
   U11323 : XNOR2_X1 port map( A => n7384, B => n18809, ZN => n7385);
   U11324 : XNOR2_X1 port map( A => n7386, B => n7385, ZN => n7387);
   U11325 : XNOR2_X1 port map( A => n7390, B => n7391, ZN => n7394);
   U11326 : XNOR2_X1 port map( A => n7392, B => n18819, ZN => n7393);
   U11327 : XNOR2_X1 port map( A => n7394, B => n7393, ZN => n7399);
   U11328 : INV_X1 port map( A => n7395, ZN => n7396);
   U11329 : XNOR2_X1 port map( A => n7397, B => n7396, ZN => n7398);
   U11330 : NAND2_X1 port map( A1 => n8928, A2 => n8932, ZN => n7662);
   U11331 : OAI21_X1 port map( B1 => n7950, B2 => n2326, A => n7951, ZN => 
                           n7404);
   U11332 : NAND2_X1 port map( A1 => n8596, A2 => n8931, ZN => n7406);
   U11333 : OAI21_X1 port map( B1 => n7662, B2 => n8931, A => n7406, ZN => 
                           n7411);
   U11334 : OAI211_X1 port map( C1 => n7826, C2 => n7830, A => n7407, B => 
                           n8012, ZN => n7410);
   U11335 : OAI21_X1 port map( B1 => n7826, B2 => n7829, A => n8011, ZN => 
                           n7409);
   U11336 : NAND2_X1 port map( A1 => n8749, A2 => n8748, ZN => n8640);
   U11337 : NAND2_X1 port map( A1 => n7411, A2 => n8640, ZN => n7412);
   U11338 : OAI21_X1 port map( B1 => n7413, B2 => n8596, A => n7412, ZN => 
                           n10299);
   U11339 : NOR2_X1 port map( A1 => n8178, A2 => n19901, ZN => n7415);
   U11340 : OAI21_X1 port map( B1 => n7416, B2 => n7415, A => n923, ZN => n7419
                           );
   U11341 : NOR2_X1 port map( A1 => n8069, A2 => n8179, ZN => n7418);
   U11342 : INV_X1 port map( A => n7420, ZN => n8201);
   U11344 : AOI21_X1 port map( B1 => n7615, B2 => n7422, A => n8201, ZN => 
                           n7423);
   U11345 : NAND2_X1 port map( A1 => n9300, A2 => n9018, ZN => n7424);
   U11346 : INV_X1 port map( A => n7644, ZN => n8215);
   U11348 : NAND2_X1 port map( A1 => n20108, A2 => n8086, ZN => n7425);
   U11349 : NOR2_X1 port map( A1 => n20107, A2 => n6539, ZN => n7426);
   U11350 : INV_X1 port map( A => n20108, ZN => n8084);
   U11351 : NAND2_X1 port map( A1 => n8084, A2 => n8085, ZN => n8236);
   U11352 : INV_X1 port map( A => n8236, ZN => n7428);
   U11353 : NAND2_X1 port map( A1 => n7631, A2 => n8212, ZN => n7431);
   U11354 : NAND2_X1 port map( A1 => n8094, A2 => n8211, ZN => n7430);
   U11355 : MUX2_X1 port map( A => n7431, B => n7430, S => n8095, Z => n7435);
   U11357 : INV_X1 port map( A => n8211, ZN => n8093);
   U11358 : INV_X1 port map( A => n8098, ZN => n7638);
   U11359 : INV_X1 port map( A => n8111, ZN => n8237);
   U11360 : MUX2_X1 port map( A => n3775, B => n7436, S => n20493, Z => n7437);
   U11362 : INV_X1 port map( A => n9304, ZN => n8845);
   U11364 : MUX2_X1 port map( A => n8323, B => n7441, S => n1425, Z => n8512);
   U11365 : OAI21_X1 port map( B1 => n7590, B2 => n7442, A => n7584, ZN => 
                           n8513);
   U11366 : BUF_X2 port map( A => n7443, Z => n8282);
   U11367 : NAND3_X1 port map( A1 => n8286, A2 => n7603, A3 => n8282, ZN => 
                           n7449);
   U11368 : NAND3_X1 port map( A1 => n7444, A2 => n3660, A3 => n7445, ZN => 
                           n7448);
   U11369 : NAND3_X1 port map( A1 => n7444, A2 => n8281, A3 => n7600, ZN => 
                           n7447);
   U11370 : INV_X1 port map( A => n8033, ZN => n8284);
   U11371 : NAND3_X1 port map( A1 => n8284, A2 => n8280, A3 => n7445, ZN => 
                           n7446);
   U11372 : AND4_X1 port map( A1 => n7448, A2 => n7449, A3 => n7447, A4 => 
                           n7446, ZN => n9021);
   U11373 : INV_X1 port map( A => n7877, ZN => n8305);
   U11376 : INV_X1 port map( A => n20257, ZN => n7789);
   U11378 : INV_X1 port map( A => n8040, ZN => n7581);
   U11379 : NAND3_X1 port map( A1 => n8297, A2 => n20243, A3 => n7581, ZN => 
                           n7454);
   U11380 : MUX2_X1 port map( A => n20243, B => n8297, S => n8298, Z => n7455);
   U11381 : INV_X1 port map( A => n8676, ZN => n8841);
   U11382 : NAND2_X1 port map( A1 => n8054, A2 => n8193, ZN => n7456);
   U11383 : NOR2_X1 port map( A1 => n8052, A2 => n8192, ZN => n7458);
   U11384 : AOI22_X1 port map( A1 => n7458, A2 => n19802, B1 => n19474, B2 => 
                           n8197, ZN => n7459);
   U11385 : INV_X1 port map( A => n8060, ZN => n7460);
   U11386 : NAND2_X1 port map( A1 => n7460, A2 => n8190, ZN => n8183);
   U11387 : INV_X1 port map( A => n8185, ZN => n8059);
   U11388 : NAND3_X1 port map( A1 => n7462, A2 => n20465, A3 => n8059, ZN => 
                           n7464);
   U11389 : NAND3_X1 port map( A1 => n8185, A2 => n7893, A3 => n8184, ZN => 
                           n7463);
   U11390 : XNOR2_X1 port map( A => n9602, B => n10482, ZN => n9984);
   U11391 : INV_X1 port map( A => n8025, ZN => n8292);
   U11392 : INV_X1 port map( A => n8026, ZN => n8024);
   U11393 : INV_X1 port map( A => n8288, ZN => n7468);
   U11394 : NAND2_X1 port map( A1 => n8292, A2 => n8026, ZN => n8031);
   U11395 : NAND2_X1 port map( A1 => n8290, A2 => n8289, ZN => n8029);
   U11396 : NAND2_X1 port map( A1 => n7470, A2 => n8024, ZN => n7471);
   U11397 : NAND2_X1 port map( A1 => n7096, A2 => n7990, ZN => n7994);
   U11398 : NAND3_X1 port map( A1 => n7096, A2 => n8011, A3 => n20154, ZN => 
                           n7472);
   U11399 : NAND2_X1 port map( A1 => n8316, A2 => n7591, ZN => n8007);
   U11400 : INV_X1 port map( A => n8007, ZN => n7474);
   U11401 : NOR2_X1 port map( A1 => n8004, A2 => n7591, ZN => n7473);
   U11402 : OAI21_X1 port map( B1 => n7474, B2 => n7473, A => n8313, ZN => 
                           n7478);
   U11404 : INV_X1 port map( A => n8004, ZN => n7476);
   U11405 : OAI21_X1 port map( B1 => n8811, B2 => n8810, A => n8815, ZN => 
                           n7486);
   U11407 : NAND3_X1 port map( A1 => n7479, A2 => n20013, A3 => n7948, ZN => 
                           n7484);
   U11408 : NOR2_X1 port map( A1 => n7952, A2 => n7951, ZN => n7480);
   U11409 : INV_X1 port map( A => n7951, ZN => n7815);
   U11410 : NAND3_X1 port map( A1 => n7949, A2 => n7951, A3 => n7953, ZN => 
                           n7482);
   U11411 : AND2_X1 port map( A1 => n8812, A2 => n8815, ZN => n7485);
   U11412 : INV_X1 port map( A => n8811, ZN => n9119);
   U11413 : AOI22_X1 port map( A1 => n8818, A2 => n7486, B1 => n7485, B2 => 
                           n9119, ZN => n7492);
   U11414 : NAND2_X1 port map( A1 => n7487, A2 => n7974, ZN => n7970);
   U11415 : INV_X1 port map( A => n7972, ZN => n7927);
   U11416 : OAI22_X1 port map( A1 => n7970, A2 => n7927, B1 => n278, B2 => 
                           n7968, ZN => n7490);
   U11417 : INV_X1 port map( A => n7487, ZN => n7973);
   U11418 : NAND2_X1 port map( A1 => n7973, A2 => n7967, ZN => n7489);
   U11419 : NAND2_X1 port map( A1 => n7972, A2 => n278, ZN => n7488);
   U11420 : NOR2_X1 port map( A1 => n8550, A2 => n9122, ZN => n9120);
   U11421 : NAND2_X1 port map( A1 => n9120, A2 => n8812, ZN => n7491);
   U11422 : INV_X1 port map( A => n7493, ZN => n8344);
   U11423 : MUX2_X1 port map( A => n8166, B => n8344, S => n8342, Z => n7495);
   U11424 : NOR2_X1 port map( A1 => n8340, A2 => n8343, ZN => n7494);
   U11426 : AND3_X1 port map( A1 => n8340, A2 => n8341, A3 => n7679, ZN => 
                           n9048);
   U11427 : INV_X1 port map( A => n9289, ZN => n9577);
   U11428 : INV_X1 port map( A => n8387, ZN => n7496);
   U11429 : AOI21_X1 port map( B1 => n7497, B2 => n7496, A => n20177, ZN => 
                           n7499);
   U11430 : INV_X1 port map( A => n7686, ZN => n8382);
   U11431 : NAND2_X1 port map( A1 => n8359, A2 => n8354, ZN => n7740);
   U11432 : NAND3_X1 port map( A1 => n7501, A2 => n7740, A3 => n7500, ZN => 
                           n7503);
   U11433 : NAND3_X1 port map( A1 => n8355, A2 => n8358, A3 => n7504, ZN => 
                           n7502);
   U11435 : AOI22_X1 port map( A1 => n2031, A2 => n20360, B1 => n20195, B2 => 
                           n7763, ZN => n7505);
   U11436 : NAND2_X1 port map( A1 => n2540, A2 => n7936, ZN => n7506);
   U11437 : OAI211_X1 port map( C1 => n7746, C2 => n7749, A => n7911, B => 
                           n7910, ZN => n7509);
   U11438 : NAND2_X1 port map( A1 => n7510, A2 => n7675, ZN => n7511);
   U11439 : NAND3_X1 port map( A1 => n8366, A2 => n7709, A3 => n8365, ZN => 
                           n7514);
   U11440 : NAND2_X1 port map( A1 => n9049, A2 => n9576, ZN => n7515);
   U11441 : AOI21_X1 port map( B1 => n9287, B2 => n7515, A => n19896, ZN => 
                           n7516);
   U11442 : AOI21_X2 port map( B1 => n9577, B2 => n20196, A => n7516, ZN => 
                           n9983);
   U11443 : XNOR2_X1 port map( A => n10028, B => n9983, ZN => n7517);
   U11444 : XNOR2_X1 port map( A => n9984, B => n7517, ZN => n7580);
   U11445 : INV_X1 port map( A => n7956, ZN => n7834);
   U11446 : MUX2_X1 port map( A => n277, B => n7834, S => n7958, Z => n8907);
   U11449 : AOI21_X1 port map( B1 => n7760, B2 => n7519, A => n2030, ZN => 
                           n8908);
   U11450 : AND2_X1 port map( A1 => n7520, A2 => n2031, ZN => n8909);
   U11451 : NAND2_X1 port map( A1 => n8923, A2 => n8917, ZN => n7533);
   U11452 : INV_X1 port map( A => n7974, ZN => n7820);
   U11454 : NAND2_X1 port map( A1 => n7523, A2 => n7970, ZN => n8733);
   U11455 : INV_X1 port map( A => n7948, ZN => n7819);
   U11456 : OAI21_X1 port map( B1 => n7819, B2 => n20013, A => n7815, ZN => 
                           n7524);
   U11457 : NAND2_X1 port map( A1 => n7524, A2 => n7949, ZN => n7526);
   U11458 : NAND3_X1 port map( A1 => n7819, A2 => n7950, A3 => n7952, ZN => 
                           n7525);
   U11459 : OAI211_X1 port map( C1 => n7818, C2 => n7948, A => n7526, B => 
                           n7525, ZN => n8735);
   U11460 : NAND2_X1 port map( A1 => n7909, A2 => n7903, ZN => n7527);
   U11461 : OAI21_X1 port map( B1 => n7909, B2 => n7754, A => n7527, ZN => 
                           n7529);
   U11462 : NOR2_X1 port map( A1 => n7754, A2 => n7902, ZN => n7528);
   U11463 : AND3_X1 port map( A1 => n7754, A2 => n19521, A3 => n7530, ZN => 
                           n7531);
   U11464 : INV_X1 port map( A => n7981, ZN => n7766);
   U11465 : NAND3_X1 port map( A1 => n7920, A2 => n7536, A3 => n7921, ZN => 
                           n7535);
   U11466 : AOI21_X1 port map( B1 => n9158, B2 => n8696, A => n9159, ZN => 
                           n7540);
   U11467 : INV_X1 port map( A => n9164, ZN => n7537);
   U11468 : NOR2_X1 port map( A1 => n7537, A2 => n9163, ZN => n9157);
   U11469 : NAND2_X1 port map( A1 => n9157, A2 => n8611, ZN => n7539);
   U11470 : NAND3_X1 port map( A1 => n1230, A2 => n8696, A3 => n9161, ZN => 
                           n7538);
   U11472 : XNOR2_X1 port map( A => n10620, B => n9947, ZN => n9416);
   U11474 : NOR2_X1 port map( A1 => n7541, A2 => n8372, ZN => n7546);
   U11475 : INV_X1 port map( A => n8376, ZN => n7703);
   U11476 : NAND3_X1 port map( A1 => n8372, A2 => n20252, A3 => n8377, ZN => 
                           n7543);
   U11477 : NAND3_X1 port map( A1 => n7544, A2 => n7543, A3 => n8369, ZN => 
                           n7545);
   U11478 : INV_X1 port map( A => n8352, ZN => n7717);
   U11479 : OAI22_X1 port map( A1 => n7717, A2 => n8140, B1 => n19914, B2 => 
                           n8347, ZN => n8351);
   U11480 : INV_X1 port map( A => n8270, ZN => n7549);
   U11481 : NOR2_X1 port map( A1 => n8349, A2 => n8348, ZN => n7548);
   U11482 : INV_X1 port map( A => n8350, ZN => n8268);
   U11483 : NAND2_X1 port map( A1 => n8268, A2 => n8140, ZN => n7547);
   U11484 : NAND2_X1 port map( A1 => n7724, A2 => n282, ZN => n7551);
   U11485 : NAND2_X1 port map( A1 => n7552, A2 => n7855, ZN => n7555);
   U11486 : NAND3_X1 port map( A1 => n7856, A2 => n7851, A3 => n7852, ZN => 
                           n7553);
   U11488 : NAND2_X1 port map( A1 => n7559, A2 => n9364, ZN => n7567);
   U11489 : AND2_X1 port map( A1 => n7560, A2 => n8114, ZN => n7843);
   U11490 : NOR2_X1 port map( A1 => n7560, A2 => n6704, ZN => n7561);
   U11491 : OAI21_X1 port map( B1 => n7843, B2 => n7561, A => n8245, ZN => 
                           n7566);
   U11493 : NOR2_X1 port map( A1 => n7844, A2 => n8114, ZN => n7563);
   U11494 : AOI22_X1 port map( A1 => n7564, A2 => n20251, B1 => n7563, B2 => 
                           n6704, ZN => n7565);
   U11495 : NAND2_X1 port map( A1 => n7567, A2 => n9362, ZN => n7577);
   U11496 : NOR2_X1 port map( A1 => n8961, A2 => n8960, ZN => n7575);
   U11497 : MUX2_X1 port map( A => n8264, B => n8263, S => n895, Z => n7569);
   U11498 : INV_X1 port map( A => n8104, ZN => n7570);
   U11499 : NAND2_X1 port map( A1 => n7570, A2 => n8262, ZN => n7573);
   U11500 : AND3_X2 port map( A1 => n7574, A2 => n7573, A3 => n7572, ZN => 
                           n8958);
   U11501 : INV_X1 port map( A => n8958, ZN => n7653);
   U11502 : AOI22_X1 port map( A1 => n7575, A2 => n7653, B1 => n8959, B2 => 
                           n8726, ZN => n7576);
   U11503 : XNOR2_X1 port map( A => n9802, B => n2344, ZN => n7578);
   U11504 : XNOR2_X1 port map( A => n9416, B => n7578, ZN => n7579);
   U11505 : XNOR2_X1 port map( A => n7580, B => n7579, ZN => n9492);
   U11506 : INV_X1 port map( A => n9492, ZN => n11160);
   U11507 : MUX2_X2 port map( A => n7583, B => n7582, S => n8299, Z => n8947);
   U11509 : INV_X1 port map( A => n7585, ZN => n8322);
   U11510 : NAND2_X1 port map( A1 => n8322, A2 => n8001, ZN => n7586);
   U11511 : OAI211_X1 port map( C1 => n1425, C2 => n8322, A => n7586, B => 
                           n8325, ZN => n7587);
   U11513 : INV_X1 port map( A => n8644, ZN => n7608);
   U11514 : INV_X1 port map( A => n7591, ZN => n7592);
   U11515 : NAND2_X1 port map( A1 => n7593, A2 => n8316, ZN => n7596);
   U11516 : NAND2_X1 port map( A1 => n7594, A2 => n7592, ZN => n7595);
   U11517 : NAND2_X1 port map( A1 => n7608, A2 => n8937, ZN => n7613);
   U11518 : NAND3_X1 port map( A1 => n8304, A2 => n8046, A3 => n8305, ZN => 
                           n7598);
   U11519 : NOR2_X1 port map( A1 => n8286, A2 => n19686, ZN => n7795);
   U11521 : NAND3_X1 port map( A1 => n8033, A2 => n8282, A3 => n8281, ZN => 
                           n7604);
   U11523 : NAND3_X1 port map( A1 => n8185, A2 => n20247, A3 => n20465, ZN => 
                           n7607);
   U11525 : NAND2_X1 port map( A1 => n7610, A2 => n8730, ZN => n7611);
   U11526 : XNOR2_X1 port map( A => n10054, B => n1782, ZN => n7655);
   U11527 : INV_X1 port map( A => n7615, ZN => n8203);
   U11528 : NAND3_X1 port map( A1 => n8201, A2 => n7421, A3 => n8204, ZN => 
                           n7617);
   U11529 : INV_X1 port map( A => n8743, ZN => n8949);
   U11530 : INV_X1 port map( A => n7887, ZN => n7620);
   U11531 : NOR2_X1 port map( A1 => n8179, A2 => n923, ZN => n7619);
   U11532 : AOI22_X1 port map( A1 => n7620, A2 => n8068, B1 => n7622, B2 => 
                           n7619, ZN => n7625);
   U11533 : INV_X1 port map( A => n7621, ZN => n8176);
   U11534 : NAND2_X1 port map( A1 => n8176, A2 => n8179, ZN => n7623);
   U11535 : INV_X1 port map( A => n8178, ZN => n7622);
   U11536 : INV_X1 port map( A => n8197, ZN => n7879);
   U11537 : AOI21_X1 port map( B1 => n7628, B2 => n7627, A => n8051, ZN => 
                           n7629);
   U11539 : NAND2_X1 port map( A1 => n8090, A2 => n7633, ZN => n7634);
   U11540 : NOR2_X1 port map( A1 => n8241, A2 => n8112, ZN => n7637);
   U11541 : NAND2_X1 port map( A1 => n7637, A2 => n3775, ZN => n7643);
   U11542 : INV_X1 port map( A => n8241, ZN => n7639);
   U11543 : NAND3_X1 port map( A1 => n8239, A2 => n7639, A3 => n7638, ZN => 
                           n7642);
   U11544 : NAND3_X1 port map( A1 => n8099, A2 => n8100, A3 => n8241, ZN => 
                           n7641);
   U11545 : NAND2_X1 port map( A1 => n8099, A2 => n8237, ZN => n7640);
   U11546 : AND2_X1 port map( A1 => n8603, A2 => n8741, ZN => n8485);
   U11547 : INV_X1 port map( A => n8485, ZN => n7650);
   U11548 : INV_X1 port map( A => n8741, ZN => n8953);
   U11549 : OAI22_X1 port map( A1 => n20441, A2 => n7645, B1 => n8220, B2 => 
                           n7644, ZN => n7847);
   U11550 : INV_X1 port map( A => n7646, ZN => n7647);
   U11551 : INV_X1 port map( A => n8742, ZN => n8950);
   U11552 : NAND2_X1 port map( A1 => n7650, A2 => n7649, ZN => n7651);
   U11553 : INV_X1 port map( A => n9362, ZN => n7654);
   U11554 : XNOR2_X1 port map( A => n10566, B => n10456, ZN => n10017);
   U11555 : XNOR2_X1 port map( A => n7655, B => n10017, ZN => n7664);
   U11556 : OAI21_X1 port map( B1 => n8527, B2 => n8848, A => n9046, ZN => 
                           n7657);
   U11557 : NAND2_X1 port map( A1 => n8749, A2 => n8747, ZN => n7661);
   U11558 : INV_X1 port map( A => n8932, ZN => n8638);
   U11559 : NAND3_X1 port map( A1 => n8638, A2 => n8749, A3 => n8925, ZN => 
                           n7660);
   U11560 : XNOR2_X1 port map( A => n9430, B => n10163, ZN => n7663);
   U11561 : INV_X1 port map( A => n8499, ZN => n7666);
   U11562 : INV_X1 port map( A => n8733, ZN => n8497);
   U11563 : NOR2_X1 port map( A1 => n8499, A2 => n8734, ZN => n8738);
   U11564 : MUX2_X1 port map( A => n7665, B => n8738, S => n8736, Z => n7670);
   U11565 : NAND2_X1 port map( A1 => n19518, A2 => n8736, ZN => n7667);
   U11566 : INV_X1 port map( A => n8736, ZN => n8916);
   U11567 : AOI22_X1 port map( A1 => n7668, A2 => n7667, B1 => n7666, B2 => 
                           n8916, ZN => n7669);
   U11569 : OAI21_X1 port map( B1 => n8146, B2 => n7671, A => n8370, ZN => 
                           n7672);
   U11570 : MUX2_X1 port map( A => n7673, B => n7709, S => n6951, Z => n7678);
   U11571 : INV_X1 port map( A => n7674, ZN => n7708);
   U11572 : INV_X1 port map( A => n8342, ZN => n8167);
   U11573 : MUX2_X1 port map( A => n2964, B => n7679, S => n8343, Z => n7682);
   U11574 : NAND3_X1 port map( A1 => n8167, A2 => n8165, A3 => n7679, ZN => 
                           n7681);
   U11575 : NOR2_X1 port map( A1 => n8340, A2 => n7679, ZN => n7733);
   U11576 : NAND2_X1 port map( A1 => n7733, A2 => n8341, ZN => n7680);
   U11579 : INV_X1 port map( A => n8386, ZN => n7683);
   U11580 : INV_X1 port map( A => n8380, ZN => n8133);
   U11581 : OAI21_X1 port map( B1 => n8132, B2 => n7683, A => n8133, ZN => 
                           n7688);
   U11583 : INV_X1 port map( A => n7714, ZN => n7687);
   U11584 : MUX2_X1 port map( A => n9358, B => n19941, S => n9528, Z => n7702);
   U11585 : OAI21_X1 port map( B1 => n7746, B2 => n3445, A => n7748, ZN => 
                           n7693);
   U11586 : NOR2_X1 port map( A1 => n7748, A2 => n7910, ZN => n7690);
   U11587 : OAI21_X1 port map( B1 => n7691, B2 => n7690, A => n7914, ZN => 
                           n7692);
   U11589 : NAND2_X1 port map( A1 => n9354, A2 => n8904, ZN => n8492);
   U11592 : NAND3_X1 port map( A1 => n7696, A2 => n7695, A3 => n8355, ZN => 
                           n7697);
   U11593 : AOI21_X2 port map( B1 => n9359, B2 => n7702, A => n7701, ZN => 
                           n10203);
   U11594 : XNOR2_X1 port map( A => n10200, B => n10203, ZN => n10596);
   U11596 : NAND2_X1 port map( A1 => n7703, A2 => n7671, ZN => n7704);
   U11597 : MUX2_X1 port map( A => n7705, B => n7704, S => n8373, Z => n7706);
   U11599 : MUX2_X1 port map( A => n8366, B => n8361, S => n7674, Z => n7712);
   U11600 : NAND3_X1 port map( A1 => n8361, A2 => n7709, A3 => n7708, ZN => 
                           n7710);
   U11601 : INV_X1 port map( A => n8879, ZN => n9255);
   U11602 : AOI21_X1 port map( B1 => n8132, B2 => n8381, A => n8387, ZN => 
                           n7713);
   U11603 : OAI22_X1 port map( A1 => n7714, A2 => n7713, B1 => n163, B2 => 
                           n8131, ZN => n7715);
   U11604 : OAI21_X1 port map( B1 => n20177, B2 => n7716, A => n7715, ZN => 
                           n9250);
   U11605 : NAND2_X1 port map( A1 => n20200, A2 => n8271, ZN => n7719);
   U11606 : NAND2_X1 port map( A1 => n8348, A2 => n8347, ZN => n7718);
   U11607 : NAND3_X1 port map( A1 => n7723, A2 => n7719, A3 => n7718, ZN => 
                           n7721);
   U11608 : OAI211_X1 port map( C1 => n7723, C2 => n7722, A => n7721, B => 
                           n7720, ZN => n8972);
   U11609 : AND2_X1 port map( A1 => n9252, A2 => n8972, ZN => n7727);
   U11610 : NAND2_X1 port map( A1 => n8167, A2 => n7728, ZN => n7732);
   U11611 : NOR2_X1 port map( A1 => n8341, A2 => n8344, ZN => n7731);
   U11612 : INV_X1 port map( A => n7729, ZN => n7730);
   U11613 : OAI21_X1 port map( B1 => n7732, B2 => n7731, A => n7730, ZN => 
                           n7735);
   U11614 : NAND2_X1 port map( A1 => n7733, A2 => n7732, ZN => n7734);
   U11615 : INV_X1 port map( A => n9249, ZN => n8971);
   U11619 : NOR2_X1 port map( A1 => n7736, A2 => n19516, ZN => n7737);
   U11620 : NAND2_X1 port map( A1 => n7740, A2 => n7739, ZN => n7744);
   U11621 : NAND2_X1 port map( A1 => n7746, A2 => n7745, ZN => n7747);
   U11622 : NOR2_X1 port map( A1 => n7747, A2 => n7912, ZN => n8124);
   U11623 : INV_X1 port map( A => n8125, ZN => n7751);
   U11624 : OAI21_X1 port map( B1 => n7002, B2 => n7908, A => n7903, ZN => 
                           n7757);
   U11625 : NAND3_X1 port map( A1 => n7754, A2 => n7753, A3 => n19521, ZN => 
                           n7756);
   U11626 : NAND2_X1 port map( A1 => n7752, A2 => n8657, ZN => n7759);
   U11627 : NAND2_X1 port map( A1 => n8658, A2 => n7759, ZN => n9003);
   U11628 : NOR2_X1 port map( A1 => n7761, A2 => n2540, ZN => n7762);
   U11629 : NAND2_X1 port map( A1 => n7931, A2 => n20359, ZN => n7765);
   U11630 : NAND2_X1 port map( A1 => n8998, A2 => n8657, ZN => n7776);
   U11631 : NAND2_X1 port map( A1 => n8999, A2 => n8998, ZN => n8443);
   U11632 : NAND2_X1 port map( A1 => n7919, A2 => n7921, ZN => n7980);
   U11634 : INV_X1 port map( A => n8998, ZN => n8773);
   U11635 : NOR2_X1 port map( A1 => n7958, A2 => n7834, ZN => n7770);
   U11636 : NAND3_X1 port map( A1 => n7836, A2 => n20165, A3 => n8906, ZN => 
                           n7771);
   U11637 : OAI21_X1 port map( B1 => n8443, B2 => n19517, A => n7774, ZN => 
                           n7775);
   U11638 : XNOR2_X1 port map( A => n9792, B => n9667, ZN => n10603);
   U11639 : NAND2_X1 port map( A1 => n19520, A2 => n8315, ZN => n7779);
   U11640 : INV_X1 port map( A => n8313, ZN => n8314);
   U11641 : NAND3_X1 port map( A1 => n8312, A2 => n8314, A3 => n19942, ZN => 
                           n7777);
   U11642 : NAND2_X1 port map( A1 => n7807, A2 => n8288, ZN => n7780);
   U11643 : INV_X1 port map( A => n7780, ZN => n7784);
   U11644 : OAI21_X1 port map( B1 => n934, B2 => n8289, A => n8292, ZN => n7783
                           );
   U11645 : NAND2_X1 port map( A1 => n8293, A2 => n20189, ZN => n7781);
   U11646 : MUX2_X1 port map( A => n7781, B => n7780, S => n8026, Z => n7782);
   U11648 : AND2_X1 port map( A1 => n7585, A2 => n8001, ZN => n8324);
   U11649 : NAND2_X1 port map( A1 => n7787, A2 => n8299, ZN => n8043);
   U11650 : NAND3_X1 port map( A1 => n8043, A2 => n8295, A3 => n7788, ZN => 
                           n7792);
   U11651 : NAND2_X1 port map( A1 => n8297, A2 => n20257, ZN => n7791);
   U11652 : AND3_X1 port map( A1 => n8297, A2 => n7789, A3 => n20485, ZN => 
                           n7790);
   U11653 : NAND2_X1 port map( A1 => n8034, A2 => n8282, ZN => n8287);
   U11654 : NAND2_X1 port map( A1 => n7793, A2 => n8287, ZN => n7794);
   U11655 : OAI21_X1 port map( B1 => n7796, B2 => n7795, A => n7794, ZN => 
                           n8761);
   U11656 : OAI21_X1 port map( B1 => n19827, B2 => n9176, A => n8760, ZN => 
                           n7805);
   U11657 : NAND2_X1 port map( A1 => n3212, A2 => n20490, ZN => n7800);
   U11658 : NAND2_X1 port map( A1 => n20347, A2 => n7801, ZN => n7799);
   U11659 : AOI21_X1 port map( B1 => n8016, B2 => n7801, A => n20270, ZN => 
                           n7802);
   U11660 : OR2_X1 port map( A1 => n7802, A2 => n3212, ZN => n7803);
   U11661 : NAND2_X1 port map( A1 => n8293, A2 => n8026, ZN => n7808);
   U11662 : NAND2_X1 port map( A1 => n8293, A2 => n8290, ZN => n7810);
   U11664 : NAND3_X1 port map( A1 => n7950, A2 => n20013, A3 => n7815, ZN => 
                           n7817);
   U11665 : MUX2_X1 port map( A => n9006, B => n8890, S => n8895, Z => n7842);
   U11666 : NAND2_X1 port map( A1 => n7972, A2 => n7820, ZN => n7825);
   U11667 : NAND2_X1 port map( A1 => n7974, A2 => n7967, ZN => n7821);
   U11668 : OAI211_X1 port map( C1 => n7967, C2 => n7968, A => n7821, B => n278
                           , ZN => n7823);
   U11669 : OAI21_X1 port map( B1 => n7922, B2 => n7968, A => n7971, ZN => 
                           n7822);
   U11670 : NAND2_X1 port map( A1 => n7823, A2 => n7822, ZN => n7824);
   U11671 : OAI21_X1 port map( B1 => n7973, B2 => n7825, A => n7824, ZN => 
                           n9008);
   U11672 : NAND3_X1 port map( A1 => n7828, A2 => n7827, A3 => n20154, ZN => 
                           n7832);
   U11673 : MUX2_X1 port map( A => n9008, B => n8895, S => n9007, Z => n7841);
   U11674 : NOR2_X1 port map( A1 => n7836, A2 => n7833, ZN => n7957);
   U11675 : INV_X1 port map( A => n7957, ZN => n7840);
   U11676 : NAND2_X1 port map( A1 => n7837, A2 => n90, ZN => n7838);
   U11677 : INV_X1 port map( A => n9009, ZN => n8623);
   U11678 : XNOR2_X1 port map( A => n9420, B => n10262, ZN => n8407);
   U11679 : XNOR2_X1 port map( A => n10603, B => n8407, ZN => n7947);
   U11680 : INV_X1 port map( A => n7843, ZN => n7846);
   U11681 : NAND2_X1 port map( A1 => n8248, A2 => n8245, ZN => n7845);
   U11682 : INV_X1 port map( A => n9271, ZN => n8984);
   U11683 : INV_X1 port map( A => n8221, ZN => n8216);
   U11684 : NAND2_X1 port map( A1 => n7847, A2 => n8216, ZN => n7850);
   U11685 : INV_X1 port map( A => n8219, ZN => n8218);
   U11686 : AOI21_X1 port map( B1 => n8215, B2 => n8218, A => n8220, ZN => 
                           n7848);
   U11688 : NOR2_X1 port map( A1 => n8984, A2 => n9265, ZN => n7870);
   U11689 : NAND2_X1 port map( A1 => n8162, A2 => n7851, ZN => n7854);
   U11690 : NAND2_X1 port map( A1 => n7856, A2 => n7855, ZN => n7853);
   U11691 : OAI21_X1 port map( B1 => n7857, B2 => n7856, A => n8160, ZN => 
                           n7858);
   U11692 : MUX2_X1 port map( A => n20108, B => n6539, S => n8086, Z => n7861);
   U11695 : INV_X1 port map( A => n7866, ZN => n9267);
   U11696 : NAND2_X1 port map( A1 => n8981, A2 => n9267, ZN => n7869);
   U11697 : NAND2_X1 port map( A1 => n8238, A2 => n8111, ZN => n7863);
   U11698 : NOR2_X1 port map( A1 => n8979, A2 => n9265, ZN => n8652);
   U11699 : OAI22_X1 port map( A1 => n8262, A2 => n7864, B1 => n8150, B2 => 
                           n8261, ZN => n8154);
   U11700 : NOR2_X1 port map( A1 => n8264, A2 => n895, ZN => n7865);
   U11701 : INV_X1 port map( A => n8153, ZN => n8107);
   U11702 : NAND2_X1 port map( A1 => n8107, A2 => n7864, ZN => n8266);
   U11703 : AOI22_X1 port map( A1 => n8154, A2 => n8106, B1 => n7865, B2 => 
                           n8266, ZN => n8653);
   U11704 : INV_X1 port map( A => n8653, ZN => n9262);
   U11705 : AOI22_X1 port map( A1 => n19880, A2 => n8652, B1 => n7867, B2 => 
                           n7866, ZN => n7868);
   U11706 : INV_X1 port map( A => n8200, ZN => n8071);
   U11707 : MUX2_X1 port map( A => n7873, B => n7872, S => n8070, Z => n7875);
   U11709 : NOR2_X1 port map( A1 => n8195, A2 => n20198, ZN => n7880);
   U11710 : AOI22_X1 port map( A1 => n7880, A2 => n7879, B1 => n7878, B2 => 
                           n8053, ZN => n7884);
   U11711 : AOI21_X1 port map( B1 => n8052, B2 => n8193, A => n8053, ZN => 
                           n7882);
   U11712 : NAND2_X1 port map( A1 => n7882, A2 => n7881, ZN => n7883);
   U11713 : NAND2_X1 port map( A1 => n1850, A2 => n923, ZN => n7886);
   U11714 : OAI21_X1 port map( B1 => n8179, B2 => n8176, A => n7622, ZN => 
                           n7885);
   U11715 : MUX2_X1 port map( A => n7886, B => n7885, S => n8181, Z => n7888);
   U11716 : NAND2_X1 port map( A1 => n9275, A2 => n20265, ZN => n7889);
   U11717 : NAND3_X1 port map( A1 => n7897, A2 => n9274, A3 => n7889, ZN => 
                           n7901);
   U11718 : NAND2_X1 port map( A1 => n8186, A2 => n7893, ZN => n7890);
   U11719 : INV_X1 port map( A => n7892, ZN => n7894);
   U11720 : NAND2_X1 port map( A1 => n7894, A2 => n7460, ZN => n7895);
   U11721 : INV_X1 port map( A => n9274, ZN => n9277);
   U11722 : NAND3_X1 port map( A1 => n19732, A2 => n9277, A3 => n20265, ZN => 
                           n7899);
   U11723 : XNOR2_X1 port map( A => n10528, B => n10264, ZN => n9974);
   U11725 : INV_X1 port map( A => n7904, ZN => n7905);
   U11726 : INV_X1 port map( A => n9149, ZN => n9144);
   U11727 : NAND2_X1 port map( A1 => n7961, A2 => n8906, ZN => n7916);
   U11729 : NAND2_X1 port map( A1 => n9144, A2 => n8337, ZN => n7944);
   U11730 : OAI21_X1 port map( B1 => n7972, B2 => n7973, A => n7974, ZN => 
                           n7925);
   U11731 : NAND2_X1 port map( A1 => n7967, A2 => n278, ZN => n7924);
   U11732 : NAND3_X1 port map( A1 => n7925, A2 => n7924, A3 => n7923, ZN => 
                           n7926);
   U11733 : OAI21_X1 port map( B1 => n7927, B2 => n7967, A => n7926, ZN => 
                           n8790);
   U11734 : NAND3_X1 port map( A1 => n7932, A2 => n1452, A3 => n7931, ZN => 
                           n7940);
   U11735 : NAND3_X1 port map( A1 => n2031, A2 => n1063, A3 => n7933, ZN => 
                           n7939);
   U11736 : NAND3_X1 port map( A1 => n2031, A2 => n7936, A3 => n20195, ZN => 
                           n7938);
   U11738 : AOI21_X2 port map( B1 => n7944, B2 => n7943, A => n7942, ZN => 
                           n9937);
   U11739 : XNOR2_X1 port map( A => n9937, B => n2341, ZN => n7945);
   U11740 : XNOR2_X1 port map( A => n9974, B => n7945, ZN => n7946);
   U11741 : INV_X1 port map( A => n11161, ZN => n10650);
   U11742 : MUX2_X1 port map( A => n9555, B => n10945, S => n10650, Z => n8402)
                           ;
   U11743 : MUX2_X1 port map( A => n7952, B => n7951, S => n7950, Z => n7954);
   U11744 : NAND2_X1 port map( A1 => n7957, A2 => n8910, ZN => n7960);
   U11745 : OAI211_X1 port map( C1 => n7962, C2 => n7961, A => n7960, B => 
                           n7959, ZN => n9171);
   U11746 : INV_X1 port map( A => n9171, ZN => n9080);
   U11747 : OAI21_X1 port map( B1 => n7965, B2 => n8017, A => n20270, ZN => 
                           n7964);
   U11748 : AOI22_X1 port map( A1 => n7966, A2 => n7965, B1 => n8016, B2 => 
                           n7964, ZN => n8568);
   U11749 : NAND2_X1 port map( A1 => n7968, A2 => n7967, ZN => n7969);
   U11750 : NAND2_X1 port map( A1 => n7973, A2 => n7972, ZN => n7975);
   U11751 : NOR2_X1 port map( A1 => n269, A2 => n8569, ZN => n7988);
   U11752 : AOI21_X1 port map( B1 => n7980, B2 => n7979, A => n7978, ZN => 
                           n7987);
   U11753 : NAND2_X1 port map( A1 => n7982, A2 => n7981, ZN => n7985);
   U11754 : AOI21_X1 port map( B1 => n7985, B2 => n7984, A => n7919, ZN => 
                           n7986);
   U11756 : OAI22_X1 port map( A1 => n8014, A2 => n20154, B1 => n8011, B2 => 
                           n7990, ZN => n8010);
   U11757 : OAI21_X1 port map( B1 => n7995, B2 => n7994, A => n7993, ZN => 
                           n9168);
   U11758 : NOR2_X2 port map( A1 => n7997, A2 => n7996, ZN => n10150);
   U11759 : NOR2_X1 port map( A1 => n7998, A2 => n8322, ZN => n8000);
   U11761 : NOR2_X1 port map( A1 => n1425, A2 => n8001, ZN => n8002);
   U11762 : NAND2_X1 port map( A1 => n19520, A2 => n8004, ZN => n8006);
   U11763 : AND2_X1 port map( A1 => n8006, A2 => n8007, ZN => n8008);
   U11765 : MUX2_X1 port map( A => n3212, B => n8017, S => n8016, Z => n8023);
   U11766 : MUX2_X1 port map( A => n8020, B => n8019, S => n3212, Z => n8021);
   U11767 : OAI21_X1 port map( B1 => n8023, B2 => n20270, A => n8021, ZN => 
                           n9062);
   U11768 : INV_X1 port map( A => n8677, ZN => n8037);
   U11769 : NAND3_X1 port map( A1 => n8290, A2 => n8024, A3 => n7468, ZN => 
                           n8030);
   U11770 : OAI21_X1 port map( B1 => n8026, B2 => n8289, A => n20189, ZN => 
                           n8027);
   U11771 : INV_X1 port map( A => n8027, ZN => n8028);
   U11772 : NAND2_X1 port map( A1 => n8034, A2 => n8280, ZN => n8035);
   U11773 : OAI21_X1 port map( B1 => n8034, B2 => n8282, A => n8281, ZN => 
                           n8032);
   U11774 : NOR3_X1 port map( A1 => n9029, A2 => n9060, A3 => n8833, ZN => 
                           n8036);
   U11775 : AOI21_X1 port map( B1 => n8037, B2 => n8831, A => n8036, ZN => 
                           n8039);
   U11776 : NAND3_X1 port map( A1 => n9031, A2 => n8829, A3 => n9060, ZN => 
                           n8038);
   U11777 : XNOR2_X1 port map( A => n10270, B => n10150, ZN => n8524);
   U11778 : OAI21_X1 port map( B1 => n8297, B2 => n8298, A => n8040, ZN => 
                           n8042);
   U11779 : AND2_X1 port map( A1 => n8040, A2 => n20485, ZN => n8296);
   U11780 : INV_X1 port map( A => n8303, ZN => n8309);
   U11781 : NAND3_X1 port map( A1 => n20001, A2 => n8045, A3 => n8044, ZN => 
                           n8049);
   U11782 : OAI211_X1 port map( C1 => n20057, C2 => n20001, A => n8047, B => 
                           n8304, ZN => n8048);
   U11783 : NAND2_X1 port map( A1 => n9836, A2 => n9066, ZN => n9069);
   U11784 : NAND2_X1 port map( A1 => n8054, A2 => n8197, ZN => n8056);
   U11785 : NAND2_X1 port map( A1 => n8056, A2 => n20198, ZN => n8057);
   U11786 : NOR2_X1 port map( A1 => n20247, A2 => n8060, ZN => n8064);
   U11787 : NOR2_X1 port map( A1 => n8185, A2 => n20465, ZN => n8063);
   U11789 : INV_X1 port map( A => n8066, ZN => n8177);
   U11791 : NOR2_X1 port map( A1 => n7421, A2 => n8070, ZN => n8073);
   U11793 : NOR2_X1 port map( A1 => n3795, A2 => n8219, ZN => n8078);
   U11794 : NOR2_X1 port map( A1 => n8079, A2 => n8215, ZN => n8080);
   U11795 : NOR3_X1 port map( A1 => n19809, A2 => n20441, A3 => n3795, ZN => 
                           n8081);
   U11796 : MUX2_X1 port map( A => n8086, B => n8085, S => n20107, Z => n8088);
   U11797 : AND2_X1 port map( A1 => n8093, A2 => n8090, ZN => n8210);
   U11798 : AOI21_X1 port map( B1 => n8094, B2 => n8093, A => n20511, ZN => 
                           n8096);
   U11799 : OR2_X1 port map( A1 => n8096, A2 => n8095, ZN => n8097);
   U11800 : NAND2_X1 port map( A1 => n9333, A2 => n9328, ZN => n8869);
   U11801 : MUX2_X1 port map( A => n8100, B => n8099, S => n8098, Z => n8102);
   U11802 : NAND2_X1 port map( A1 => n8241, A2 => n8100, ZN => n8244);
   U11803 : INV_X1 port map( A => n8244, ZN => n8101);
   U11804 : MUX2_X1 port map( A => n8102, B => n8101, S => n3775, Z => n8463);
   U11805 : INV_X1 port map( A => n8463, ZN => n8119);
   U11807 : AND2_X1 port map( A1 => n8104, A2 => n8261, ZN => n8110);
   U11808 : NAND2_X1 port map( A1 => n8151, A2 => n895, ZN => n8105);
   U11809 : NAND2_X1 port map( A1 => n8106, A2 => n8105, ZN => n8108);
   U11810 : NAND2_X1 port map( A1 => n8108, A2 => n8107, ZN => n8109);
   U11811 : INV_X1 port map( A => n9330, ZN => n9074);
   U11812 : AND3_X1 port map( A1 => n8112, A2 => n8239, A3 => n8111, ZN => 
                           n8462);
   U11813 : INV_X1 port map( A => n8462, ZN => n8118);
   U11814 : NAND4_X1 port map( A1 => n8119, A2 => n20008, A3 => n9074, A4 => 
                           n8118, ZN => n8123);
   U11815 : NAND2_X1 port map( A1 => n8245, A2 => n8246, ZN => n8117);
   U11816 : OAI21_X1 port map( B1 => n8114, B2 => n8113, A => n8248, ZN => 
                           n8116);
   U11817 : MUX2_X1 port map( A => n8117, B => n8116, S => n20251, Z => n8120);
   U11818 : NAND4_X1 port map( A1 => n8119, A2 => n900, A3 => n8120, A4 => 
                           n8118, ZN => n8121);
   U11819 : XNOR2_X1 port map( A => n10552, B => n10271, ZN => n9998);
   U11820 : XNOR2_X1 port map( A => n9998, B => n8524, ZN => n8173);
   U11821 : OR2_X1 port map( A1 => n7752, A2 => n8657, ZN => n8660);
   U11822 : XNOR2_X1 port map( A => n9635, B => n17587, ZN => n8171);
   U11823 : INV_X1 port map( A => n8470, ZN => n9091);
   U11824 : NAND2_X1 port map( A1 => n8884, A2 => n9453, ZN => n8889);
   U11825 : NAND2_X1 port map( A1 => n8387, A2 => n8132, ZN => n8137);
   U11826 : NAND2_X1 port map( A1 => n8133, A2 => n8381, ZN => n8134);
   U11827 : MUX2_X1 port map( A => n20200, B => n8272, S => n8348, Z => n8139);
   U11828 : OAI21_X1 port map( B1 => n8370, B2 => n8377, A => n8142, ZN => 
                           n8144);
   U11829 : NAND2_X1 port map( A1 => n20294, A2 => n20252, ZN => n8143);
   U11830 : NAND2_X1 port map( A1 => n8144, A2 => n8143, ZN => n8148);
   U11831 : INV_X1 port map( A => n8261, ZN => n8149);
   U11832 : OAI21_X1 port map( B1 => n7571, B2 => n8150, A => n8149, ZN => 
                           n8152);
   U11833 : INV_X1 port map( A => n8156, ZN => n9341);
   U11834 : NAND2_X1 port map( A1 => n9341, A2 => n9346, ZN => n8701);
   U11835 : NOR2_X1 port map( A1 => n8157, A2 => n6830, ZN => n8158);
   U11836 : NOR2_X1 port map( A1 => n8159, A2 => n8158, ZN => n8161);
   U11837 : NOR2_X1 port map( A1 => n9341, A2 => n9563, ZN => n9191);
   U11838 : NAND2_X1 port map( A1 => n9191, A2 => n9564, ZN => n8168);
   U11839 : XNOR2_X1 port map( A => n9999, B => n918, ZN => n10584);
   U11840 : XNOR2_X1 port map( A => n10584, B => n8171, ZN => n8172);
   U11841 : INV_X1 port map( A => n10945, ZN => n8174);
   U11842 : NAND2_X1 port map( A1 => n8174, A2 => n11158, ZN => n8399);
   U11843 : NOR2_X1 port map( A1 => n8178, A2 => n8177, ZN => n8180);
   U11844 : AND2_X1 port map( A1 => n8182, A2 => n8184, ZN => n8191);
   U11845 : INV_X1 port map( A => n8183, ZN => n8188);
   U11846 : OAI21_X1 port map( B1 => n8188, B2 => n8187, A => n8186, ZN => 
                           n8189);
   U11847 : NAND2_X1 port map( A1 => n9218, A2 => n908, ZN => n8228);
   U11848 : OAI21_X1 port map( B1 => n8196, B2 => n8195, A => n8194, ZN => 
                           n8198);
   U11849 : NAND2_X1 port map( A1 => n8198, A2 => n8197, ZN => n8199);
   U11850 : INV_X1 port map( A => n9221, ZN => n8795);
   U11851 : NAND3_X1 port map( A1 => n8205, A2 => n819, A3 => n8203, ZN => 
                           n8206);
   U11852 : NAND2_X1 port map( A1 => n8210, A2 => n8209, ZN => n8214);
   U11853 : OAI211_X1 port map( C1 => n7631, C2 => n8212, A => n7633, B => 
                           n8211, ZN => n8213);
   U11854 : NOR2_X1 port map( A1 => n9114, A2 => n9113, ZN => n8225);
   U11855 : NAND2_X1 port map( A1 => n8218, A2 => n20180, ZN => n8222);
   U11856 : OAI22_X1 port map( A1 => n8222, A2 => n19809, B1 => n8219, B2 => 
                           n20174, ZN => n8223);
   U11857 : AND2_X1 port map( A1 => n8797, A2 => n9113, ZN => n8428);
   U11858 : AOI22_X1 port map( A1 => n8226, A2 => n8225, B1 => n8428, B2 => 
                           n8795, ZN => n8227);
   U11859 : NAND2_X1 port map( A1 => n8228, A2 => n8227, ZN => n9769);
   U11860 : MUX2_X1 port map( A => n20107, B => n8230, S => n20495, Z => n8235)
                           ;
   U11861 : AND2_X1 port map( A1 => n6539, A2 => n8232, ZN => n8234);
   U11862 : OAI21_X1 port map( B1 => n8239, B2 => n8098, A => n8237, ZN => 
                           n8240);
   U11863 : NAND2_X1 port map( A1 => n8240, A2 => n3775, ZN => n8243);
   U11864 : NOR3_X1 port map( A1 => n8435, A2 => n8434, A3 => n9201, ZN => 
                           n8279);
   U11865 : NAND2_X1 port map( A1 => n8247, A2 => n8246, ZN => n8249);
   U11866 : OR2_X1 port map( A1 => n8256, A2 => n7724, ZN => n8257);
   U11868 : NOR2_X1 port map( A1 => n8349, A2 => n19914, ZN => n8269);
   U11869 : OAI21_X1 port map( B1 => n8270, B2 => n8269, A => n8268, ZN => 
                           n8275);
   U11870 : NAND2_X1 port map( A1 => n8273, A2 => n20200, ZN => n8274);
   U11871 : NAND2_X1 port map( A1 => n9129, A2 => n8276, ZN => n8432);
   U11872 : OR2_X1 port map( A1 => n8432, A2 => n9201, ZN => n8277);
   U11874 : XNOR2_X1 port map( A => n9769, B => n10431, ZN => n9996);
   U11875 : NOR2_X1 port map( A1 => n20012, A2 => n8282, ZN => n8285);
   U11876 : NOR2_X1 port map( A1 => n8287, A2 => n8286, ZN => n8421);
   U11877 : OAI21_X1 port map( B1 => n8290, B2 => n8289, A => n934, ZN => n8291
                           );
   U11878 : OAI211_X1 port map( C1 => n8300, C2 => n8299, A => n8298, B => 
                           n8297, ZN => n9099);
   U11879 : OAI21_X1 port map( B1 => n8303, B2 => n20001, A => n8301, ZN => 
                           n8308);
   U11880 : NAND2_X1 port map( A1 => n20057, A2 => n8304, ZN => n8307);
   U11882 : NAND2_X1 port map( A1 => n7592, A2 => n8314, ZN => n8318);
   U11883 : NAND2_X1 port map( A1 => n19942, A2 => n8315, ZN => n8317);
   U11884 : MUX2_X1 port map( A => n8318, B => n8317, S => n8316, Z => n8319);
   U11885 : NAND2_X1 port map( A1 => n8872, A2 => n9106, ZN => n8559);
   U11886 : NAND3_X1 port map( A1 => n8559, A2 => n9107, A3 => n20000, ZN => 
                           n8326);
   U11888 : INV_X1 port map( A => n9120, ZN => n8331);
   U11889 : INV_X1 port map( A => n9122, ZN => n8814);
   U11890 : NAND2_X1 port map( A1 => n8815, A2 => n9122, ZN => n8328);
   U11891 : XNOR2_X1 port map( A => n9861, B => n19990, ZN => n8469);
   U11892 : XNOR2_X1 port map( A => n8469, B => n9996, ZN => n8398);
   U11893 : AND2_X1 port map( A1 => n8332, A2 => n8734, ZN => n8335);
   U11894 : INV_X1 port map( A => n9648, ZN => n8339);
   U11895 : INV_X1 port map( A => n9143, ZN => n8338);
   U11896 : MUX2_X1 port map( A => n8341, B => n3121, S => n8340, Z => n8346);
   U11897 : MUX2_X1 port map( A => n20274, B => n8343, S => n8342, Z => n8345);
   U11898 : AOI21_X1 port map( B1 => n8349, B2 => n8348, A => n8347, ZN => 
                           n8353);
   U11899 : NAND2_X1 port map( A1 => n8355, A2 => n8354, ZN => n8356);
   U11900 : NAND2_X1 port map( A1 => n8364, A2 => n8363, ZN => n8368);
   U11901 : NAND2_X1 port map( A1 => n1994, A2 => n8365, ZN => n8367);
   U11902 : NAND3_X1 port map( A1 => n20294, A2 => n8373, A3 => n8372, ZN => 
                           n8379);
   U11903 : NAND3_X1 port map( A1 => n8377, A2 => n20252, A3 => n8375, ZN => 
                           n8378);
   U11904 : INV_X1 port map( A => n8389, ZN => n8392);
   U11907 : NAND2_X1 port map( A1 => n8386, A2 => n8385, ZN => n8388);
   U11908 : MUX2_X1 port map( A => n8389, B => n8388, S => n8387, Z => n8390);
   U11909 : NAND3_X1 port map( A1 => n9212, A2 => n9211, A3 => n8420, ZN => 
                           n8393);
   U11910 : XNOR2_X1 port map( A => n10236, B => n2448, ZN => n8395);
   U11911 : XNOR2_X1 port map( A => n8396, B => n8395, ZN => n8397);
   U11913 : AOI21_X1 port map( B1 => n8400, B2 => n8399, A => n11159, ZN => 
                           n8401);
   U11914 : MUX2_X1 port map( A => n8569, B => n9171, S => n9167, Z => n8404);
   U11915 : MUX2_X1 port map( A => n9163, B => n9160, S => n8611, Z => n8406);
   U11916 : MUX2_X1 port map( A => n9159, B => n9162, S => n9158, Z => n8405);
   U11917 : XNOR2_X1 port map( A => n9794, B => n10472, ZN => n8408);
   U11918 : XNOR2_X1 port map( A => n8408, B => n8407, ZN => n8418);
   U11919 : MUX2_X1 port map( A => n8713, B => n9241, S => n9240, Z => n8410);
   U11920 : MUX2_X1 port map( A => n9240, B => n9242, S => n6587, Z => n8409);
   U11921 : MUX2_X1 port map( A => n8410, B => n8409, S => n266, Z => n10526);
   U11925 : XNOR2_X1 port map( A => n10425, B => n10526, ZN => n9459);
   U11926 : NAND2_X1 port map( A1 => n9564, A2 => n9338, ZN => n8413);
   U11927 : MUX2_X1 port map( A => n8699, B => n8413, S => n9567, Z => n8414);
   U11928 : OAI21_X2 port map( B1 => n8415, B2 => n9338, A => n8414, ZN => 
                           n10265);
   U11929 : XNOR2_X1 port map( A => n10265, B => n2257, ZN => n8416);
   U11930 : XNOR2_X1 port map( A => n9459, B => n8416, ZN => n8417);
   U11931 : XNOR2_X1 port map( A => n8418, B => n8417, ZN => n10756);
   U11932 : NOR2_X1 port map( A1 => n9111, A2 => n9106, ZN => n8424);
   U11933 : OAI21_X1 port map( B1 => n8555, B2 => n9105, A => n9111, ZN => 
                           n8425);
   U11934 : XNOR2_X1 port map( A => n10620, B => n18075, ZN => n8426);
   U11935 : XNOR2_X1 port map( A => n8427, B => n8426, ZN => n8441);
   U11936 : NOR2_X1 port map( A1 => n9219, A2 => n9112, ZN => n8431);
   U11937 : NAND2_X1 port map( A1 => n8428, A2 => n9217, ZN => n8430);
   U11938 : AND2_X1 port map( A1 => n8433, A2 => n8432, ZN => n8437);
   U11939 : AOI21_X1 port map( B1 => n9130, B2 => n8276, A => n8805, ZN => 
                           n8436);
   U11940 : OAI22_X1 port map( A1 => n8437, A2 => n9780, B1 => n9204, B2 => 
                           n8436, ZN => n9535);
   U11941 : XNOR2_X1 port map( A => n10072, B => n9535, ZN => n10543);
   U11942 : NAND2_X1 port map( A1 => n9151, A2 => n9143, ZN => n8438);
   U11943 : NAND2_X1 port map( A1 => n9151, A2 => n8790, ZN => n8789);
   U11944 : XNOR2_X1 port map( A => n10028, B => n8769, ZN => n10480);
   U11945 : XNOR2_X1 port map( A => n10480, B => n10543, ZN => n8440);
   U11946 : OAI21_X1 port map( B1 => n8995, B2 => n8443, A => n8442, ZN => 
                           n9923);
   U11947 : NOR2_X1 port map( A1 => n9209, A2 => n8445, ZN => n8446);
   U11948 : XNOR2_X1 port map( A => n10303, B => n9923, ZN => n9738);
   U11949 : OAI21_X1 port map( B1 => n9275, B2 => n9274, A => n8650, ZN => 
                           n8449);
   U11950 : XNOR2_X1 port map( A => n8450, B => n10114, ZN => n8451);
   U11951 : XNOR2_X1 port map( A => n9738, B => n8451, ZN => n8461);
   U11952 : OAI21_X1 port map( B1 => n8979, B2 => n2118, A => n9267, ZN => 
                           n8453);
   U11953 : NOR2_X1 port map( A1 => n8979, A2 => n19710, ZN => n8452);
   U11954 : INV_X1 port map( A => n8550, ZN => n9128);
   U11956 : NAND3_X1 port map( A1 => n9119, A2 => n8552, A3 => n8810, ZN => 
                           n8455);
   U11957 : OAI211_X2 port map( C1 => n9128, C2 => n8457, A => n8456, B => 
                           n8455, ZN => n10572);
   U11958 : XNOR2_X1 port map( A => n10570, B => n10572, ZN => n8459);
   U11959 : XNOR2_X1 port map( A => n10054, B => n2067, ZN => n8458);
   U11960 : XNOR2_X1 port map( A => n8459, B => n8458, ZN => n8460);
   U11961 : XNOR2_X1 port map( A => n8461, B => n8460, ZN => n11526);
   U11962 : INV_X1 port map( A => n9331, ZN => n9073);
   U11963 : NOR2_X1 port map( A1 => n9836, A2 => n9066, ZN => n8545);
   U11964 : INV_X1 port map( A => n9834, ZN => n9317);
   U11965 : XNOR2_X1 port map( A => n9647, B => n10557, ZN => n9470);
   U11966 : XNOR2_X1 port map( A => n9470, B => n8469, ZN => n8481);
   U11967 : NAND2_X1 port map( A1 => n9451, A2 => n9453, ZN => n8474);
   U11968 : NAND3_X1 port map( A1 => n1576, A2 => n9090, A3 => n9091, ZN => 
                           n8473);
   U11969 : NAND3_X1 port map( A1 => n8474, A2 => n8473, A3 => n8472, ZN => 
                           n9812);
   U11971 : OAI21_X1 port map( B1 => n670, B2 => n8972, A => n8971, ZN => n8476
                           );
   U11972 : NAND3_X1 port map( A1 => n9249, A2 => n9256, A3 => n8879, ZN => 
                           n8475);
   U11973 : XNOR2_X1 port map( A => n10281, B => n9812, ZN => n9722);
   U11974 : INV_X1 port map( A => n9007, ZN => n9004);
   U11975 : NAND2_X1 port map( A1 => n9004, A2 => n19490, ZN => n8477);
   U11976 : INV_X1 port map( A => n8895, ZN => n8891);
   U11977 : OAI211_X1 port map( C1 => n19490, C2 => n9008, A => n8891, B => 
                           n9005, ZN => n8478);
   U11978 : XNOR2_X1 port map( A => n10497, B => n17999, ZN => n8479);
   U11979 : XNOR2_X1 port map( A => n9722, B => n8479, ZN => n8480);
   U11981 : NOR2_X1 port map( A1 => n10756, A2 => n11527, ZN => n10635);
   U11983 : MUX2_X1 port map( A => n8485, B => n8483, S => n9368, Z => n8487);
   U11984 : NOR2_X1 port map( A1 => n8603, A2 => n8742, ZN => n8484);
   U11985 : MUX2_X1 port map( A => n8945, B => n8941, S => n8729, Z => n8489);
   U11986 : NOR2_X1 port map( A1 => n8944, A2 => n8939, ZN => n8490);
   U11988 : XNOR2_X1 port map( A => n10442, B => n10402, ZN => n9445);
   U11989 : INV_X1 port map( A => n8492, ZN => n8496);
   U11990 : OAI21_X1 port map( B1 => n8904, B2 => n8720, A => n9358, ZN => 
                           n8495);
   U11991 : NAND2_X1 port map( A1 => n8722, A2 => n9528, ZN => n8493);
   U11992 : MUX2_X1 port map( A => n8493, B => n8492, S => n9359, Z => n8494);
   U11994 : XNOR2_X1 port map( A => n10506, B => n9817, ZN => n8507);
   U11995 : NAND2_X1 port map( A1 => n9361, A2 => n207, ZN => n8505);
   U11996 : NAND2_X1 port map( A1 => n9363, A2 => n9362, ZN => n8501);
   U11997 : MUX2_X1 port map( A => n8502, B => n8501, S => n8961, Z => n8504);
   U11998 : NAND3_X1 port map( A1 => n8958, A2 => n8726, A3 => n207, ZN => 
                           n8503);
   U11999 : XNOR2_X1 port map( A => n19785, B => n2356, ZN => n8506);
   U12000 : XNOR2_X1 port map( A => n8507, B => n8506, ZN => n8508);
   U12001 : INV_X1 port map( A => n11527, ZN => n10919);
   U12002 : INV_X1 port map( A => n11521, ZN => n11530);
   U12003 : NOR2_X1 port map( A1 => n8676, A2 => n9023, ZN => n9022);
   U12006 : INV_X1 port map( A => n8512, ZN => n8517);
   U12007 : NAND3_X1 port map( A1 => n8517, A2 => n8516, A3 => n8515, ZN => 
                           n8518);
   U12008 : NOR2_X1 port map( A1 => n8846, A2 => n9300, ZN => n8523);
   U12009 : NOR2_X1 port map( A1 => n9018, A2 => n9295, ZN => n8842);
   U12010 : AOI22_X1 port map( A1 => n9304, A2 => n8842, B1 => n8520, B2 => 
                           n8846, ZN => n8521);
   U12011 : XNOR2_X1 port map( A => n10551, B => n10461, ZN => n9476);
   U12012 : XNOR2_X1 port map( A => n9476, B => n8524, ZN => n8536);
   U12013 : NOR2_X1 port map( A1 => n8527, A2 => n9039, ZN => n8526);
   U12014 : NOR2_X1 port map( A1 => n9046, A2 => n8851, ZN => n8525);
   U12015 : NAND3_X1 port map( A1 => n8527, A2 => n9046, A3 => n8848, ZN => 
                           n8528);
   U12016 : OAI21_X1 port map( B1 => n9037, B2 => n8529, A => n8528, ZN => 
                           n8530);
   U12017 : NOR2_X2 port map( A1 => n8531, A2 => n8530, ZN => n10491);
   U12018 : NOR2_X1 port map( A1 => n9291, A2 => n9576, ZN => n8532);
   U12019 : XNOR2_X1 port map( A => n9824, B => n10491, ZN => n8534);
   U12020 : NAND2_X1 port map( A1 => n8823, A2 => n9307, ZN => n9054);
   U12021 : XNOR2_X1 port map( A => n10274, B => n2218, ZN => n8533);
   U12022 : XNOR2_X1 port map( A => n8534, B => n8533, ZN => n8535);
   U12024 : NOR2_X1 port map( A1 => n9331, A2 => n9326, ZN => n8538);
   U12025 : AOI22_X1 port map( A1 => n8539, A2 => n9333, B1 => n8538, B2 => 
                           n9329, ZN => n8540);
   U12027 : NOR2_X1 port map( A1 => n8543, A2 => n8542, ZN => n8547);
   U12028 : XNOR2_X1 port map( A => n872, B => n10604, ZN => n9503);
   U12030 : INV_X1 port map( A => n9420, ZN => n10173);
   U12031 : XNOR2_X1 port map( A => n10173, B => n2442, ZN => n8548);
   U12033 : NOR2_X1 port map( A1 => n8550, A2 => n8813, ZN => n8551);
   U12034 : AOI21_X1 port map( B1 => n8552, B2 => n8818, A => n8551, ZN => 
                           n8554);
   U12035 : INV_X1 port map( A => n9107, ZN => n8871);
   U12036 : OAI21_X1 port map( B1 => n8871, B2 => n9111, A => n9106, ZN => 
                           n8558);
   U12037 : INV_X1 port map( A => n8555, ZN => n8557);
   U12038 : INV_X1 port map( A => n8780, ZN => n8556);
   U12039 : INV_X1 port map( A => n8559, ZN => n8560);
   U12040 : NAND2_X1 port map( A1 => n9111, A2 => n8560, ZN => n8561);
   U12041 : XNOR2_X1 port map( A => n10171, B => n10421, ZN => n9208);
   U12042 : INV_X1 port map( A => n9087, ZN => n8562);
   U12043 : OAI211_X1 port map( C1 => n9451, C2 => n8884, A => n8563, B => 
                           n1576, ZN => n8564);
   U12044 : OAI21_X1 port map( B1 => n1576, B2 => n9454, A => n8564, ZN => 
                           n9500);
   U12045 : XNOR2_X1 port map( A => n9500, B => n19767, ZN => n9750);
   U12046 : XNOR2_X1 port map( A => n9208, B => n9750, ZN => n8566);
   U12048 : NOR3_X1 port map( A1 => n9167, A2 => n9080, A3 => n9166, ZN => 
                           n8570);
   U12049 : INV_X1 port map( A => n8833, ZN => n9059);
   U12050 : INV_X1 port map( A => n9029, ZN => n8571);
   U12051 : MUX2_X1 port map( A => n8829, B => n8571, S => n9060, Z => n8575);
   U12053 : MUX2_X1 port map( A => n8573, B => n8572, S => n8829, Z => n8574);
   U12054 : XNOR2_X1 port map( A => n10254, B => n10186, ZN => n9325);
   U12055 : NAND2_X1 port map( A1 => n9579, A2 => n19896, ZN => n8581);
   U12056 : NAND3_X1 port map( A1 => n8577, A2 => n19519, A3 => n19715, ZN => 
                           n8580);
   U12057 : AND2_X1 port map( A1 => n9291, A2 => n9576, ZN => n9290);
   U12058 : NOR2_X1 port map( A1 => n19896, A2 => n9576, ZN => n8578);
   U12059 : OAI21_X1 port map( B1 => n9290, B2 => n8578, A => n9287, ZN => 
                           n8579);
   U12060 : OAI211_X1 port map( C1 => n9289, C2 => n8581, A => n8580, B => 
                           n8579, ZN => n9844);
   U12061 : XNOR2_X1 port map( A => n9844, B => n10252, ZN => n9773);
   U12062 : XNOR2_X1 port map( A => n9325, B => n9773, ZN => n8591);
   U12063 : MUX2_X1 port map( A => n891, B => n8846, S => n2984, Z => n8585);
   U12064 : NAND2_X1 port map( A1 => n9304, A2 => n9296, ZN => n8583);
   U12065 : INV_X1 port map( A => n8671, ZN => n8588);
   U12066 : INV_X1 port map( A => n9023, ZN => n8836);
   U12067 : INV_X1 port map( A => n9021, ZN => n8837);
   U12068 : NAND2_X1 port map( A1 => n8672, A2 => n8837, ZN => n8586);
   U12069 : XNOR2_X1 port map( A => n10612, B => n10367, ZN => n9512);
   U12070 : XNOR2_X1 port map( A => n9842, B => n2384, ZN => n8589);
   U12071 : XNOR2_X1 port map( A => n9512, B => n8589, ZN => n8590);
   U12072 : XNOR2_X1 port map( A => n9754, B => n8593, ZN => n10182);
   U12073 : NAND2_X1 port map( A1 => n8947, A2 => n8937, ZN => n8728);
   U12074 : OAI21_X1 port map( B1 => n8939, B2 => n8945, A => n8728, ZN => 
                           n8648);
   U12075 : AOI21_X2 port map( B1 => n8644, B2 => n8648, A => n8594, ZN => 
                           n10320);
   U12076 : XNOR2_X1 port map( A => n10320, B => n2375, ZN => n8595);
   U12077 : XNOR2_X1 port map( A => n10182, B => n8595, ZN => n8608);
   U12078 : INV_X1 port map( A => n8928, ZN => n8752);
   U12079 : INV_X1 port map( A => n8925, ZN => n8639);
   U12081 : OAI22_X1 port map( A1 => n8752, A2 => n8639, B1 => n8933, B2 => 
                           n8931, ZN => n8643);
   U12082 : INV_X1 port map( A => n8749, ZN => n8929);
   U12083 : NAND2_X1 port map( A1 => n8932, A2 => n8925, ZN => n8597);
   U12085 : NAND2_X1 port map( A1 => n9037, A2 => n9045, ZN => n8601);
   U12086 : NAND2_X1 port map( A1 => n9039, A2 => n9038, ZN => n8599);
   U12087 : AOI21_X1 port map( B1 => n8599, B2 => n8851, A => n8849, ZN => 
                           n8600);
   U12088 : AOI21_X1 port map( B1 => n8601, B2 => n8848, A => n8600, ZN => 
                           n9402);
   U12089 : XNOR2_X1 port map( A => n9402, B => n10179, ZN => n9232);
   U12090 : INV_X1 port map( A => n9232, ZN => n8606);
   U12091 : NAND2_X1 port map( A1 => n9372, A2 => n9367, ZN => n8605);
   U12092 : OAI21_X1 port map( B1 => n8953, B2 => n8742, A => n8603, ZN => 
                           n8604);
   U12093 : AOI22_X1 port map( A1 => n8605, A2 => n8743, B1 => n8956, B2 => 
                           n8604, ZN => n9537);
   U12094 : INV_X1 port map( A => n9537, ZN => n10286);
   U12096 : INV_X1 port map( A => n9756, ZN => n10619);
   U12097 : XNOR2_X1 port map( A => n10619, B => n8606, ZN => n8607);
   U12098 : OAI21_X1 port map( B1 => n11544, B2 => n11545, A => n11550, ZN => 
                           n8692);
   U12100 : NAND3_X1 port map( A1 => n9160, A2 => n8609, A3 => n9159, ZN => 
                           n8612);
   U12101 : INV_X1 port map( A => n9879, ZN => n8615);
   U12102 : XNOR2_X1 port map( A => n8615, B => n10150, ZN => n8627);
   U12103 : NOR2_X1 port map( A1 => n9172, A2 => n8761, ZN => n8616);
   U12105 : NAND2_X1 port map( A1 => n9172, A2 => n9177, ZN => n8619);
   U12106 : INV_X1 port map( A => n9176, ZN => n8617);
   U12107 : NAND3_X1 port map( A1 => n9005, A2 => n8895, A3 => n9007, ZN => 
                           n8625);
   U12108 : NAND3_X1 port map( A1 => n8623, A2 => n8891, A3 => n8622, ZN => 
                           n8624);
   U12110 : INV_X1 port map( A => n8713, ZN => n9239);
   U12111 : NAND3_X1 port map( A1 => n266, A2 => n9239, A3 => n9186, ZN => 
                           n8629);
   U12112 : OAI21_X1 port map( B1 => n9233, B2 => n1041, A => n19716, ZN => 
                           n8634);
   U12113 : XNOR2_X1 port map( A => n10359, B => n10582, ZN => n9508);
   U12114 : XNOR2_X1 port map( A => n917, B => n16487, ZN => n8635);
   U12117 : NAND2_X1 port map( A1 => n8933, A2 => n8747, ZN => n8642);
   U12118 : AND3_X1 port map( A1 => n8640, A2 => n8639, A3 => n8638, ZN => 
                           n8641);
   U12120 : NAND2_X1 port map( A1 => n111, A2 => n8937, ZN => n8647);
   U12121 : OAI211_X1 port map( C1 => n8644, C2 => n8937, A => n8941, B => 
                           n8945, ZN => n8645);
   U12122 : INV_X1 port map( A => n8645, ZN => n8646);
   U12123 : AOI21_X2 port map( B1 => n8648, B2 => n8647, A => n8646, ZN => 
                           n10157);
   U12124 : XNOR2_X1 port map( A => n10157, B => n10240, ZN => n9360);
   U12125 : INV_X1 port map( A => n8649, ZN => n9273);
   U12126 : OAI211_X1 port map( C1 => n9273, C2 => n20265, A => n9277, B => 
                           n9275, ZN => n8651);
   U12127 : NAND2_X1 port map( A1 => n8771, A2 => n19710, ZN => n8654);
   U12129 : XNOR2_X1 port map( A => n10351, B => n10589, ZN => n9523);
   U12130 : INV_X1 port map( A => n9523, ZN => n8656);
   U12131 : XNOR2_X1 port map( A => n8656, B => n9360, ZN => n8664);
   U12132 : NOR2_X1 port map( A1 => n8998, A2 => n19517, ZN => n8659);
   U12133 : XNOR2_X1 port map( A => n9861, B => n9862, ZN => n8662);
   U12134 : XNOR2_X1 port map( A => n10236, B => n18366, ZN => n8661);
   U12135 : XNOR2_X1 port map( A => n8662, B => n8661, ZN => n8663);
   U12136 : XNOR2_X1 port map( A => n8664, B => n8663, ZN => n10760);
   U12137 : INV_X1 port map( A => n10760, ZN => n11549);
   U12138 : INV_X1 port map( A => n10928, ZN => n8689);
   U12140 : NOR2_X1 port map( A1 => n20146, A2 => n8805, ZN => n9781);
   U12143 : NAND3_X1 port map( A1 => n9217, A2 => n1428, A3 => n9114, ZN => 
                           n8668);
   U12144 : XNOR2_X1 port map( A => n10595, B => n20161, ZN => n9518);
   U12145 : OAI21_X1 port map( B1 => n19857, B2 => n8672, A => n8671, ZN => 
                           n8673);
   U12147 : NAND2_X1 port map( A1 => n8831, A2 => n9029, ZN => n9032);
   U12148 : OAI21_X1 port map( B1 => n9031, B2 => n9060, A => n9032, ZN => 
                           n8679);
   U12149 : INV_X1 port map( A => n9062, ZN => n8830);
   U12150 : NAND2_X1 port map( A1 => n8677, A2 => n9059, ZN => n8678);
   U12152 : XNOR2_X1 port map( A => n10567, B => n19806, ZN => n9294);
   U12153 : XNOR2_X1 port map( A => n8680, B => n9518, ZN => n8687);
   U12154 : XNOR2_X1 port map( A => n10163, B => n10203, ZN => n8685);
   U12155 : NOR2_X1 port map( A1 => n8338, A2 => n8786, ZN => n8682);
   U12156 : XNOR2_X1 port map( A => n9777, B => n18819, ZN => n8684);
   U12157 : XNOR2_X1 port map( A => n8685, B => n8684, ZN => n8686);
   U12158 : XNOR2_X1 port map( A => n8687, B => n8686, ZN => n11548);
   U12160 : NAND2_X1 port map( A1 => n647, A2 => n11546, ZN => n8688);
   U12161 : NAND2_X1 port map( A1 => n8689, A2 => n8688, ZN => n8691);
   U12162 : NOR2_X1 port map( A1 => n10926, A2 => n11546, ZN => n8690);
   U12164 : NAND2_X1 port map( A1 => n8987, A2 => n8761, ZN => n8695);
   U12165 : OAI21_X1 port map( B1 => n19827, B2 => n8695, A => n8694, ZN => 
                           n10043);
   U12166 : INV_X1 port map( A => n10497, ZN => n9589);
   U12167 : XNOR2_X1 port map( A => n10043, B => n9589, ZN => n9524);
   U12168 : OAI21_X1 port map( B1 => n9159, B2 => n9162, A => n8609, ZN => 
                           n8697);
   U12169 : INV_X1 port map( A => n8699, ZN => n8704);
   U12170 : OAI21_X1 port map( B1 => n19590, B2 => n9340, A => n8700, ZN => 
                           n9072);
   U12171 : NAND2_X1 port map( A1 => n9072, A2 => n8701, ZN => n8702);
   U12172 : OAI21_X1 port map( B1 => n8704, B2 => n8703, A => n8702, ZN => 
                           n9685);
   U12173 : XNOR2_X1 port map( A => n10280, B => n9685, ZN => n9651);
   U12174 : XNOR2_X1 port map( A => n9524, B => n9651, ZN => n8719);
   U12175 : NAND2_X1 port map( A1 => n269, A2 => n9168, ZN => n9081);
   U12176 : INV_X1 port map( A => n9168, ZN => n8706);
   U12177 : OAI211_X1 port map( C1 => n9171, C2 => n9166, A => n264, B => n8706
                           , ZN => n8707);
   U12178 : NAND3_X1 port map( A1 => n2097, A2 => n8411, A3 => n1041, ZN => 
                           n8710);
   U12179 : OAI211_X1 port map( C1 => n8712, C2 => n8711, A => n8710, B => 
                           n9236, ZN => n10088);
   U12180 : XNOR2_X1 port map( A => n9908, B => n10088, ZN => n8717);
   U12181 : XNOR2_X1 port map( A => n8717, B => n8716, ZN => n8718);
   U12182 : OAI22_X1 port map( A1 => n8721, A2 => n8720, B1 => n8905, B2 => 
                           n9358, ZN => n8725);
   U12183 : NOR2_X1 port map( A1 => n19941, A2 => n8904, ZN => n8723);
   U12184 : XNOR2_X1 port map( A => n10273, B => n10126, ZN => n9632);
   U12185 : NOR2_X1 port map( A1 => n8729, A2 => n8937, ZN => n8732);
   U12186 : NOR3_X1 port map( A1 => n8917, A2 => n8736, A3 => n8735, ZN => 
                           n8737);
   U12187 : AOI21_X1 port map( B1 => n8738, B2 => n3645, A => n8737, ZN => 
                           n8739);
   U12188 : XNOR2_X1 port map( A => n9632, B => n8740, ZN => n8757);
   U12189 : NOR2_X1 port map( A1 => n8741, A2 => n8950, ZN => n9371);
   U12190 : NAND2_X1 port map( A1 => n8482, A2 => n8743, ZN => n8744);
   U12192 : XNOR2_X1 port map( A => n10213, B => n2151, ZN => n8755);
   U12193 : NOR2_X1 port map( A1 => n8932, A2 => n8747, ZN => n8751);
   U12194 : NOR2_X1 port map( A1 => n8749, A2 => n8748, ZN => n8750);
   U12196 : XNOR2_X1 port map( A => n9952, B => n10491, ZN => n9507);
   U12197 : XNOR2_X1 port map( A => n8755, B => n9507, ZN => n8756);
   U12199 : INV_X1 port map( A => n9172, ZN => n8765);
   U12200 : INV_X1 port map( A => n8761, ZN => n9178);
   U12201 : NOR2_X1 port map( A1 => n19827, A2 => n9178, ZN => n8762);
   U12202 : OAI21_X1 port map( B1 => n8763, B2 => n8762, A => n9177, ZN => 
                           n8764);
   U12203 : OAI21_X1 port map( B1 => n8766, B2 => n8765, A => n8764, ZN => 
                           n10071);
   U12204 : XNOR2_X1 port map( A => n9894, B => n10071, ZN => n8770);
   U12205 : AOI22_X1 port map( A1 => n8768, A2 => n9008, B1 => n8767, B2 => 
                           n9004, ZN => n9710);
   U12206 : XNOR2_X1 port map( A => n9600, B => n9710, ZN => n9538);
   U12207 : XNOR2_X1 port map( A => n8770, B => n9538, ZN => n8778);
   U12208 : OAI21_X1 port map( B1 => n8773, B2 => n8772, A => n8997, ZN => 
                           n8774);
   U12209 : NAND2_X1 port map( A1 => n8774, A2 => n3518, ZN => n8775);
   U12211 : XNOR2_X1 port map( A => n8777, B => n8778, ZN => n10640);
   U12212 : NOR2_X1 port map( A1 => n9107, A2 => n9105, ZN => n8784);
   U12213 : OAI21_X1 port map( B1 => n8779, B2 => n20000, A => n9111, ZN => 
                           n8783);
   U12214 : INV_X1 port map( A => n8872, ZN => n8781);
   U12215 : NAND3_X1 port map( A1 => n1960, A2 => n8781, A3 => n9106, ZN => 
                           n8782);
   U12217 : INV_X1 port map( A => n8790, ZN => n9148);
   U12218 : INV_X1 port map( A => n8789, ZN => n8792);
   U12219 : NOR2_X1 port map( A1 => n9145, A2 => n8790, ZN => n8791);
   U12220 : XNOR2_X1 port map( A => n20211, B => n9771, ZN => n8802);
   U12221 : INV_X1 port map( A => n8793, ZN => n8794);
   U12222 : AND3_X1 port map( A1 => n1603, A2 => n8794, A3 => n9217, ZN => 
                           n8800);
   U12223 : INV_X1 port map( A => n8796, ZN => n8799);
   U12224 : AND2_X1 port map( A1 => n9114, A2 => n8797, ZN => n8798);
   U12225 : XNOR2_X1 port map( A => n10247, B => n2382, ZN => n8801);
   U12226 : XNOR2_X1 port map( A => n8802, B => n8801, ZN => n8822);
   U12227 : NAND2_X1 port map( A1 => n8803, A2 => n9135, ZN => n8804);
   U12228 : NAND2_X1 port map( A1 => n9204, A2 => n8665, ZN => n8809);
   U12229 : NOR2_X1 port map( A1 => n9129, A2 => n8276, ZN => n8806);
   U12230 : OAI21_X1 port map( B1 => n9202, B2 => n8806, A => n3542, ZN => 
                           n8808);
   U12231 : NAND2_X1 port map( A1 => n9782, A2 => n9129, ZN => n8807);
   U12232 : OAI211_X1 port map( C1 => n9780, C2 => n8809, A => n8808, B => 
                           n8807, ZN => n9691);
   U12233 : XNOR2_X1 port map( A => n9691, B => n10296, ZN => n8820);
   U12234 : MUX2_X1 port map( A => n8811, B => n8810, S => n8815, Z => n8819);
   U12235 : NAND2_X1 port map( A1 => n9122, A2 => n8812, ZN => n8817);
   U12236 : NAND3_X1 port map( A1 => n8815, A2 => n8814, A3 => n8813, ZN => 
                           n8816);
   U12237 : XNOR2_X1 port map( A => n10506, B => n10404, ZN => n9514);
   U12238 : XNOR2_X1 port map( A => n9514, B => n8820, ZN => n8821);
   U12239 : MUX2_X1 port map( A => n8823, B => n9228, S => n9313, Z => n8827);
   U12240 : NAND2_X1 port map( A1 => n9305, A2 => n9228, ZN => n8825);
   U12241 : OAI21_X1 port map( B1 => n9307, B2 => n8827, A => n8826, ZN => 
                           n9668);
   U12242 : XNOR2_X1 port map( A => n10261, B => n9668, ZN => n9625);
   U12243 : INV_X1 port map( A => n9031, ZN => n9061);
   U12244 : NAND3_X1 port map( A1 => n9061, A2 => n9060, A3 => n9029, ZN => 
                           n8835);
   U12245 : INV_X1 port map( A => n9060, ZN => n9028);
   U12246 : NAND2_X1 port map( A1 => n8831, A2 => n8830, ZN => n8832);
   U12247 : NAND3_X1 port map( A1 => n8833, A2 => n9029, A3 => n9028, ZN => 
                           n8834);
   U12248 : XNOR2_X1 port map( A => n9934, B => n10472, ZN => n9499);
   U12249 : XNOR2_X1 port map( A => n9625, B => n9499, ZN => n8859);
   U12250 : MUX2_X1 port map( A => n8839, B => n8838, S => n19857, Z => n8840);
   U12251 : NAND2_X1 port map( A1 => n2984, A2 => n9018, ZN => n8844);
   U12252 : INV_X1 port map( A => n8842, ZN => n8843);
   U12253 : OAI22_X1 port map( A1 => n8845, A2 => n8844, B1 => n8843, B2 => 
                           n20472, ZN => n8847);
   U12255 : XNOR2_X1 port map( A => n9623, B => n10422, ZN => n9407);
   U12256 : NOR2_X1 port map( A1 => n9046, A2 => n8848, ZN => n9040);
   U12257 : NOR2_X1 port map( A1 => n9046, A2 => n9038, ZN => n8850);
   U12258 : MUX2_X1 port map( A => n9040, B => n8850, S => n8849, Z => n8856);
   U12259 : NOR2_X1 port map( A1 => n8852, A2 => n8851, ZN => n8854);
   U12260 : NOR2_X1 port map( A1 => n1933, A2 => n9039, ZN => n8853);
   U12262 : XNOR2_X1 port map( A => n20483, B => n19467, ZN => n8857);
   U12263 : XNOR2_X1 port map( A => n9407, B => n8857, ZN => n8858);
   U12264 : XNOR2_X1 port map( A => n8858, B => n8859, ZN => n10638);
   U12265 : INV_X1 port map( A => n9066, ZN => n9321);
   U12266 : NOR2_X1 port map( A1 => n9837, A2 => n9065, ZN => n8862);
   U12267 : OR2_X1 port map( A1 => n9317, A2 => n9066, ZN => n8861);
   U12268 : AOI22_X1 port map( A1 => n8862, A2 => n9069, B1 => n8861, B2 => 
                           n9065, ZN => n8863);
   U12269 : INV_X1 port map( A => n8866, ZN => n9327);
   U12270 : OAI21_X1 port map( B1 => n8866, B2 => n9326, A => n9074, ZN => 
                           n8865);
   U12271 : NAND2_X1 port map( A1 => n8865, A2 => n9329, ZN => n8868);
   U12273 : OAI211_X2 port map( C1 => n8869, C2 => n9327, A => n8868, B => 
                           n8867, ZN => n10204);
   U12274 : XNOR2_X1 port map( A => n10594, B => n10204, ZN => n8878);
   U12276 : NAND2_X1 port map( A1 => n8872, A2 => n19515, ZN => n8876);
   U12277 : OAI21_X1 port map( B1 => n8872, B2 => n9106, A => n9105, ZN => 
                           n8870);
   U12278 : NAND2_X1 port map( A1 => n8871, A2 => n8870, ZN => n8875);
   U12279 : NOR2_X1 port map( A1 => n8781, A2 => n20000, ZN => n8873);
   U12280 : OAI211_X2 port map( C1 => n1960, C2 => n8876, A => n8875, B => 
                           n8874, ZN => n10388);
   U12281 : INV_X1 port map( A => n10572, ZN => n8877);
   U12282 : XNOR2_X1 port map( A => n8877, B => n10388, ZN => n9520);
   U12283 : XNOR2_X1 port map( A => n8878, B => n9520, ZN => n8900);
   U12284 : INV_X1 port map( A => n8972, ZN => n9251);
   U12285 : NAND2_X1 port map( A1 => n19516, A2 => n9249, ZN => n8883);
   U12286 : NAND2_X1 port map( A1 => n8974, A2 => n8879, ZN => n8882);
   U12287 : OAI21_X1 port map( B1 => n9252, B2 => n8972, A => n670, ZN => n8881
                           );
   U12288 : INV_X1 port map( A => n8884, ZN => n9452);
   U12289 : AND3_X1 port map( A1 => n8887, A2 => n8886, A3 => n8885, ZN => 
                           n8888);
   U12290 : XNOR2_X1 port map( A => n9429, B => n9922, ZN => n8898);
   U12291 : INV_X1 port map( A => n9008, ZN => n8896);
   U12292 : OAI21_X1 port map( B1 => n9004, B2 => n9008, A => n19490, ZN => 
                           n8893);
   U12293 : NAND2_X1 port map( A1 => n8891, A2 => n8890, ZN => n8892);
   U12294 : OAI21_X1 port map( B1 => n8896, B2 => n8895, A => n8894, ZN => 
                           n9926);
   U12295 : XNOR2_X1 port map( A => n9926, B => n2323, ZN => n8897);
   U12296 : XNOR2_X1 port map( A => n8898, B => n8897, ZN => n8899);
   U12297 : NAND2_X1 port map( A1 => n11538, A2 => n11532, ZN => n8901);
   U12298 : MUX2_X1 port map( A => n8902, B => n8901, S => n11534, Z => n8903);
   U12299 : NAND2_X1 port map( A1 => n8907, A2 => n8906, ZN => n8915);
   U12300 : INV_X1 port map( A => n8908, ZN => n8914);
   U12301 : INV_X1 port map( A => n8909, ZN => n8913);
   U12302 : NAND2_X1 port map( A1 => n8911, A2 => n8910, ZN => n8912);
   U12303 : NAND4_X1 port map( A1 => n8915, A2 => n8914, A3 => n8913, A4 => 
                           n8912, ZN => n8919);
   U12304 : NAND4_X1 port map( A1 => n8921, A2 => n8920, A3 => n8919, A4 => 
                           n8918, ZN => n8922);
   U12305 : NOR2_X1 port map( A1 => n8932, A2 => n8931, ZN => n8927);
   U12306 : INV_X1 port map( A => n8924, ZN => n8926);
   U12309 : NAND2_X1 port map( A1 => n8932, A2 => n8931, ZN => n8934);
   U12310 : XNOR2_X1 port map( A => n9624, B => n20484, ZN => n9456);
   U12311 : XNOR2_X1 port map( A => n8936, B => n9456, ZN => n8969);
   U12313 : NAND2_X1 port map( A1 => n8953, A2 => n904, ZN => n8955);
   U12314 : NAND3_X1 port map( A1 => n8953, A2 => n8952, A3 => n8482, ZN => 
                           n8954);
   U12315 : OAI21_X1 port map( B1 => n8956, B2 => n8955, A => n8954, ZN => 
                           n8957);
   U12316 : XNOR2_X1 port map( A => n10527, B => n9670, ZN => n9421);
   U12317 : NOR2_X1 port map( A1 => n9362, A2 => n8961, ZN => n8962);
   U12318 : NAND2_X1 port map( A1 => n8962, A2 => n9363, ZN => n8963);
   U12319 : NAND2_X1 port map( A1 => n8964, A2 => n8963, ZN => n8967);
   U12320 : NOR2_X1 port map( A1 => n8965, A2 => n8726, ZN => n8966);
   U12321 : NOR2_X2 port map( A1 => n8967, A2 => n8966, ZN => n9869);
   U12322 : XNOR2_X1 port map( A => n9421, B => n9869, ZN => n8968);
   U12323 : XNOR2_X1 port map( A => n8969, B => n8968, ZN => n9017);
   U12324 : NOR2_X1 port map( A1 => n9256, A2 => n9255, ZN => n8973);
   U12325 : AND2_X1 port map( A1 => n8973, A2 => n8974, ZN => n8975);
   U12326 : AND2_X1 port map( A1 => n8979, A2 => n19710, ZN => n8980);
   U12327 : NAND2_X1 port map( A1 => n8984, A2 => n8980, ZN => n8982);
   U12328 : OAI211_X1 port map( C1 => n8984, C2 => n8983, A => n8982, B => 
                           n3797, ZN => n9398);
   U12329 : INV_X1 port map( A => n9398, ZN => n10094);
   U12330 : XNOR2_X1 port map( A => n9692, B => n10094, ZN => n8994);
   U12331 : NAND2_X1 port map( A1 => n9177, A2 => n8987, ZN => n8989);
   U12332 : OAI21_X1 port map( B1 => n265, B2 => n9178, A => n9172, ZN => n8986
                           );
   U12333 : NAND2_X1 port map( A1 => n265, A2 => n9176, ZN => n9175);
   U12334 : MUX2_X1 port map( A => n8987, B => n8986, S => n9175, Z => n8988);
   U12335 : OAI21_X1 port map( B1 => n9172, B2 => n8989, A => n8988, ZN => 
                           n10613);
   U12336 : XNOR2_X1 port map( A => n10441, B => n10613, ZN => n10257);
   U12337 : XNOR2_X1 port map( A => n10257, B => n8994, ZN => n9016);
   U12338 : MUX2_X1 port map( A => n19517, B => n8998, S => n8997, Z => n9001);
   U12339 : NAND3_X1 port map( A1 => n8999, A2 => n8998, A3 => n8997, ZN => 
                           n9000);
   U12340 : OAI21_X1 port map( B1 => n9001, B2 => n8657, A => n9000, ZN => 
                           n9002);
   U12341 : XNOR2_X1 port map( A => n10026, B => n2248, ZN => n9014);
   U12342 : INV_X1 port map( A => n9010, ZN => n9013);
   U12343 : OAI21_X1 port map( B1 => n9006, B2 => n9005, A => n9004, ZN => 
                           n9012);
   U12344 : XNOR2_X1 port map( A => n10008, B => n9771, ZN => n9446);
   U12345 : XNOR2_X1 port map( A => n9446, B => n9014, ZN => n9015);
   U12346 : XNOR2_X1 port map( A => n9016, B => n9015, ZN => n11553);
   U12348 : NOR2_X1 port map( A1 => n9304, A2 => n9018, ZN => n9020);
   U12349 : AND2_X1 port map( A1 => n19857, A2 => n9021, ZN => n9027);
   U12350 : INV_X1 port map( A => n9022, ZN => n9026);
   U12351 : NOR2_X1 port map( A1 => n9062, A2 => n9029, ZN => n9030);
   U12352 : NOR2_X1 port map( A1 => n9034, A2 => n9030, ZN => n9036);
   U12353 : INV_X1 port map( A => n9032, ZN => n9033);
   U12354 : NAND2_X1 port map( A1 => n9034, A2 => n9033, ZN => n9035);
   U12355 : XNOR2_X1 port map( A => n9908, B => n9991, ZN => n9469);
   U12356 : XNOR2_X1 port map( A => n10242, B => n9469, ZN => n9058);
   U12357 : INV_X1 port map( A => n9037, ZN => n9043);
   U12358 : NOR2_X1 port map( A1 => n9039, A2 => n9038, ZN => n9042);
   U12359 : INV_X1 port map( A => n9040, ZN => n9041);
   U12360 : OAI21_X1 port map( B1 => n9043, B2 => n9042, A => n9041, ZN => 
                           n9044);
   U12361 : NOR2_X1 port map( A1 => n9049, A2 => n9576, ZN => n9050);
   U12362 : XNOR2_X1 port map( A => n10046, B => n10350, ZN => n9056);
   U12363 : NAND2_X1 port map( A1 => n1751, A2 => n20011, ZN => n9226);
   U12365 : XNOR2_X1 port map( A => n10087, B => n2385, ZN => n9055);
   U12366 : XNOR2_X1 port map( A => n9056, B => n9055, ZN => n9057);
   U12367 : XNOR2_X1 port map( A => n9058, B => n9057, ZN => n10913);
   U12368 : AOI21_X1 port map( B1 => n9061, B2 => n9060, A => n9059, ZN => 
                           n9064);
   U12369 : OAI21_X1 port map( B1 => n9317, B2 => n9065, A => n9837, ZN => 
                           n9068);
   U12370 : AND3_X1 port map( A1 => n20476, A2 => n9837, A3 => n9066, ZN => 
                           n9067);
   U12371 : XNOR2_X1 port map( A => n865, B => n10220, ZN => n9415);
   U12372 : INV_X1 port map( A => n9070, ZN => n9339);
   U12373 : OAI21_X1 port map( B1 => n19590, B2 => n9564, A => n9563, ZN => 
                           n9071);
   U12374 : AOI22_X1 port map( A1 => n9075, A2 => n9329, B1 => n9074, B2 => 
                           n9333, ZN => n9079);
   U12377 : XNOR2_X1 port map( A => n9414, B => n10382, ZN => n9674);
   U12378 : XNOR2_X1 port map( A => n9415, B => n9674, ZN => n9097);
   U12379 : AOI21_X1 port map( B1 => n1027, B2 => n9081, A => n9080, ZN => 
                           n9084);
   U12381 : XNOR2_X1 port map( A => n20134, B => n9986, ZN => n9464);
   U12382 : NOR2_X1 port map( A1 => n9087, A2 => n20010, ZN => n9094);
   U12383 : NAND2_X1 port map( A1 => n9089, A2 => n9088, ZN => n9093);
   U12384 : NAND3_X1 port map( A1 => n9452, A2 => n9091, A3 => n9090, ZN => 
                           n9092);
   U12386 : XNOR2_X1 port map( A => n10027, B => n19222, ZN => n9095);
   U12387 : XNOR2_X1 port map( A => n9464, B => n9095, ZN => n9096);
   U12390 : AOI21_X1 port map( B1 => n19564, B2 => n10913, A => n19957, ZN => 
                           n9098);
   U12391 : NAND3_X1 port map( A1 => n9107, A2 => n9106, A3 => n9105, ZN => 
                           n9108);
   U12392 : OAI211_X1 port map( C1 => n9111, C2 => n9110, A => n9109, B => 
                           n9108, ZN => n10578);
   U12393 : NAND3_X1 port map( A1 => n1056, A2 => n8795, A3 => n9112, ZN => 
                           n9117);
   U12394 : XNOR2_X1 port map( A => n10578, B => n10154, ZN => n10210);
   U12395 : NAND2_X1 port map( A1 => n9120, A2 => n9119, ZN => n9126);
   U12396 : AOI22_X1 port map( A1 => n9124, A2 => n9128, B1 => n9123, B2 => 
                           n9122, ZN => n9125);
   U12397 : XNOR2_X1 port map( A => n10079, B => n9902, ZN => n9477);
   U12398 : XNOR2_X1 port map( A => n20491, B => n9477, ZN => n9156);
   U12399 : NAND2_X1 port map( A1 => n9780, A2 => n3542, ZN => n9132);
   U12402 : INV_X1 port map( A => n9134, ZN => n9142);
   U12403 : NOR2_X1 port map( A1 => n9211, A2 => n9214, ZN => n9136);
   U12404 : NAND2_X1 port map( A1 => n9213, A2 => n9136, ZN => n9141);
   U12405 : AND2_X1 port map( A1 => n9137, A2 => n9214, ZN => n9139);
   U12406 : AOI22_X1 port map( A1 => n9213, A2 => n9139, B1 => n9138, B2 => 
                           n9211, ZN => n9140);
   U12407 : XNOR2_X1 port map( A => n19945, B => n10358, ZN => n9154);
   U12408 : NOR2_X1 port map( A1 => n9144, A2 => n9143, ZN => n9152);
   U12410 : XNOR2_X1 port map( A => n10061, B => n20394, ZN => n9153);
   U12411 : XNOR2_X1 port map( A => n9154, B => n9153, ZN => n9155);
   U12412 : NAND2_X1 port map( A1 => n10913, A2 => n11556, ZN => n10645);
   U12413 : OR2_X1 port map( A1 => n10645, A2 => n9017, ZN => n9200);
   U12414 : INV_X1 port map( A => n11556, ZN => n11162);
   U12415 : AND2_X1 port map( A1 => n9164, A2 => n9163, ZN => n9165);
   U12416 : OAI21_X1 port map( B1 => n9167, B2 => n9171, A => n9166, ZN => 
                           n9170);
   U12417 : NAND2_X1 port map( A1 => n264, A2 => n9168, ZN => n9169);
   U12418 : NAND2_X1 port map( A1 => n264, A2 => n9171, ZN => n10328);
   U12420 : XNOR2_X1 port map( A => n9587, B => n10052, ZN => n9179);
   U12421 : OAI21_X1 port map( B1 => n9172, B2 => n9177, A => n2243, ZN => 
                           n9174);
   U12422 : INV_X1 port map( A => n9177, ZN => n9173);
   U12423 : XNOR2_X1 port map( A => n9926, B => n9643, ZN => n9480);
   U12424 : XNOR2_X1 port map( A => n9480, B => n9179, ZN => n9198);
   U12425 : NAND2_X1 port map( A1 => n9234, A2 => n19716, ZN => n9180);
   U12426 : AOI21_X1 port map( B1 => n9183, B2 => n9182, A => n9234, ZN => 
                           n9184);
   U12427 : NAND2_X1 port map( A1 => n9186, A2 => n9241, ZN => n9187);
   U12428 : AOI21_X1 port map( B1 => n9188, B2 => n9187, A => n9242, ZN => 
                           n9703);
   U12429 : OR2_X1 port map( A1 => n9703, A2 => n9700, ZN => n10166);
   U12430 : XNOR2_X1 port map( A => n10166, B => n10571, ZN => n10201);
   U12431 : OAI21_X1 port map( B1 => n9339, B2 => n9563, A => n9342, ZN => 
                           n9192);
   U12432 : NOR2_X1 port map( A1 => n9192, A2 => n9191, ZN => n9195);
   U12433 : AOI21_X1 port map( B1 => n8701, B2 => n9193, A => n9339, ZN => 
                           n9194);
   U12434 : XNOR2_X1 port map( A => n10107, B => n2023, ZN => n9196);
   U12435 : XNOR2_X1 port map( A => n10201, B => n9196, ZN => n9197);
   U12436 : XNOR2_X1 port map( A => n9197, B => n9198, ZN => n11559);
   U12437 : INV_X1 port map( A => n11559, ZN => n10914);
   U12438 : NAND3_X1 port map( A1 => n19957, A2 => n11162, A3 => n10914, ZN => 
                           n9199);
   U12439 : NAND2_X1 port map( A1 => n12354, A2 => n12349, ZN => n11032);
   U12440 : XNOR2_X1 port map( A => n10229, B => n18779, ZN => n9206);
   U12441 : XNOR2_X1 port map( A => n19746, B => n9206, ZN => n9207);
   U12442 : XNOR2_X1 port map( A => n9208, B => n9207, ZN => n9225);
   U12443 : XNOR2_X1 port map( A => n9977, B => n9937, ZN => n10098);
   U12444 : NAND2_X1 port map( A1 => n9218, A2 => n1056, ZN => n9216);
   U12445 : OAI21_X1 port map( B1 => n9218, B2 => n9217, A => n9216, ZN => 
                           n9223);
   U12446 : NOR2_X1 port map( A1 => n9220, A2 => n9219, ZN => n9222);
   U12447 : XNOR2_X1 port map( A => n10098, B => n10473, ZN => n9224);
   U12448 : INV_X1 port map( A => n9305, ZN => n9308);
   U12449 : AOI21_X1 port map( B1 => n9227, B2 => n9226, A => n9308, ZN => 
                           n9231);
   U12450 : INV_X1 port map( A => n9228, ZN => n9306);
   U12451 : AOI21_X1 port map( B1 => n9229, B2 => n20011, A => n9306, ZN => 
                           n9230);
   U12452 : XNOR2_X1 port map( A => n10417, B => n9232, ZN => n9248);
   U12453 : INV_X1 port map( A => n9234, ZN => n9235);
   U12454 : XNOR2_X1 port map( A => n10484, B => n10027, ZN => n9246);
   U12456 : XNOR2_X1 port map( A => n9854, B => n17365, ZN => n9245);
   U12457 : XNOR2_X1 port map( A => n9246, B => n9245, ZN => n9247);
   U12458 : XNOR2_X1 port map( A => n9248, B => n9247, ZN => n9351);
   U12459 : NAND2_X1 port map( A1 => n9252, A2 => n9251, ZN => n9253);
   U12460 : NAND3_X1 port map( A1 => n9260, A2 => n670, A3 => n9253, ZN => 
                           n9258);
   U12461 : NAND3_X1 port map( A1 => n19516, A2 => n9256, A3 => n9255, ZN => 
                           n9257);
   U12462 : XNOR2_X1 port map( A => n10462, B => n9261, ZN => n9286);
   U12463 : INV_X1 port map( A => n9264, ZN => n9269);
   U12464 : NOR2_X1 port map( A1 => n9266, A2 => n9265, ZN => n9268);
   U12466 : XNOR2_X1 port map( A => n19718, B => n10360, ZN => n9284);
   U12467 : XNOR2_X1 port map( A => n10061, B => n2383, ZN => n9283);
   U12468 : XNOR2_X1 port map( A => n9284, B => n9283, ZN => n9285);
   U12469 : XNOR2_X2 port map( A => n9286, B => n9285, ZN => n11174);
   U12470 : NOR2_X1 port map( A1 => n19715, A2 => n9576, ZN => n9288);
   U12471 : AOI22_X1 port map( A1 => n9578, A2 => n9291, B1 => n9577, B2 => 
                           n9290, ZN => n9292);
   U12472 : NAND2_X1 port map( A1 => n9582, A2 => n9292, ZN => n9293);
   U12473 : XNOR2_X1 port map( A => n9293, B => n9430, ZN => n10453);
   U12474 : XNOR2_X1 port map( A => n9294, B => n10453, ZN => n9316);
   U12475 : INV_X1 port map( A => n9299, ZN => n9301);
   U12476 : NAND2_X1 port map( A1 => n9301, A2 => n9300, ZN => n9302);
   U12477 : MUX2_X1 port map( A => n9306, B => n9307, S => n9305, Z => n9314);
   U12478 : NAND3_X1 port map( A1 => n9308, A2 => n9307, A3 => n1751, ZN => 
                           n9312);
   U12479 : NAND2_X1 port map( A1 => n20011, A2 => n9309, ZN => n9311);
   U12480 : XNOR2_X1 port map( A => n10205, B => n2401, ZN => n9315);
   U12481 : NAND2_X1 port map( A1 => n20505, A2 => n9837, ZN => n9320);
   U12482 : NOR2_X1 port map( A1 => n9837, A2 => n9317, ZN => n9318);
   U12483 : NOR2_X1 port map( A1 => n9321, A2 => n9836, ZN => n9322);
   U12484 : XNOR2_X1 port map( A => n9324, B => n9325, ZN => n9350);
   U12485 : NAND2_X1 port map( A1 => n9329, A2 => n3800, ZN => n9335);
   U12486 : NOR2_X1 port map( A1 => n9331, A2 => n9330, ZN => n9332);
   U12487 : NAND2_X1 port map( A1 => n9333, A2 => n9332, ZN => n9334);
   U12488 : XNOR2_X1 port map( A => n10248, B => n18854, ZN => n9348);
   U12489 : NAND2_X1 port map( A1 => n9339, A2 => n9338, ZN => n9566);
   U12490 : NAND3_X1 port map( A1 => n19590, A2 => n9346, A3 => n9340, ZN => 
                           n9343);
   U12491 : NAND3_X1 port map( A1 => n9342, A2 => n9341, A3 => n9563, ZN => 
                           n9568);
   U12492 : AND2_X1 port map( A1 => n9343, A2 => n9568, ZN => n9345);
   U12493 : NAND3_X1 port map( A1 => n9564, A2 => n9346, A3 => n9563, ZN => 
                           n9344);
   U12494 : OAI211_X1 port map( C1 => n9346, C2 => n9566, A => n9345, B => 
                           n9344, ZN => n9347);
   U12495 : XNOR2_X1 port map( A => n9957, B => n9347, ZN => n10447);
   U12496 : XNOR2_X1 port map( A => n9348, B => n10447, ZN => n9349);
   U12497 : XNOR2_X1 port map( A => n9350, B => n9349, ZN => n11175);
   U12498 : NOR2_X1 port map( A1 => n11175, A2 => n11178, ZN => n9379);
   U12499 : NOR2_X1 port map( A1 => n19941, A2 => n2756, ZN => n9355);
   U12500 : XNOR2_X1 port map( A => n10436, B => n9648, ZN => n10085);
   U12501 : XNOR2_X1 port map( A => n10085, B => n9360, ZN => n9377);
   U12502 : NOR2_X1 port map( A1 => n9362, A2 => n9361, ZN => n9365);
   U12503 : XNOR2_X1 port map( A => n10349, B => n10046, ZN => n9375);
   U12504 : INV_X1 port map( A => n9367, ZN => n9369);
   U12505 : NAND2_X1 port map( A1 => n9373, A2 => n9372, ZN => n10498);
   U12506 : XNOR2_X1 port map( A => n10498, B => n345, ZN => n9374);
   U12507 : XNOR2_X1 port map( A => n9375, B => n9374, ZN => n9376);
   U12508 : NOR3_X1 port map( A1 => n12002, A2 => n12001, A3 => n19769, ZN => 
                           n9380);
   U12509 : XNOR2_X1 port map( A => n9383, B => n10002, ZN => n9679);
   U12510 : XNOR2_X1 port map( A => n10077, B => n10273, ZN => n10409);
   U12511 : XNOR2_X1 port map( A => n10409, B => n9679, ZN => n9386);
   U12512 : XNOR2_X1 port map( A => n9824, B => n10061, ZN => n9728);
   U12513 : XNOR2_X1 port map( A => n10213, B => n2347, ZN => n9384);
   U12514 : XNOR2_X1 port map( A => n9728, B => n9384, ZN => n9385);
   U12515 : XNOR2_X1 port map( A => n9386, B => n9385, ZN => n11283);
   U12516 : INV_X1 port map( A => n11283, ZN => n11282);
   U12517 : XNOR2_X1 port map( A => n10240, B => n10088, ZN => n10433);
   U12518 : XNOR2_X1 port map( A => n9812, B => n10046, ZN => n9387);
   U12519 : XNOR2_X1 port map( A => n10397, B => n9388, ZN => n9389);
   U12520 : INV_X1 port map( A => n10199, ZN => n9392);
   U12521 : XNOR2_X1 port map( A => n10107, B => n9429, ZN => n10392);
   U12522 : XNOR2_X1 port map( A => n10392, B => n10454, ZN => n9396);
   U12523 : XNOR2_X1 port map( A => n9923, B => n10204, ZN => n9394);
   U12524 : XNOR2_X1 port map( A => n10052, B => n404, ZN => n9393);
   U12525 : XNOR2_X1 port map( A => n9394, B => n9393, ZN => n9395);
   U12526 : XNOR2_X1 port map( A => n9396, B => n9395, ZN => n10693);
   U12527 : INV_X1 port map( A => n10693, ZN => n11281);
   U12529 : INV_X1 port map( A => n20210, ZN => n9397);
   U12530 : XNOR2_X1 port map( A => n9397, B => n10254, ZN => n10444);
   U12531 : XNOR2_X1 port map( A => n10026, B => n9817, ZN => n9717);
   U12532 : XNOR2_X1 port map( A => n10444, B => n9717, ZN => n9401);
   U12533 : XNOR2_X1 port map( A => n10247, B => n2222, ZN => n9399);
   U12534 : XNOR2_X1 port map( A => n10406, B => n9399, ZN => n9400);
   U12535 : XNOR2_X1 port map( A => n9401, B => n9400, ZN => n9559);
   U12536 : XNOR2_X1 port map( A => n10027, B => n9799, ZN => n9713);
   U12537 : INV_X1 port map( A => n9402, ZN => n10219);
   U12538 : XNOR2_X1 port map( A => n10219, B => n19818, ZN => n10416);
   U12539 : XNOR2_X1 port map( A => n20268, B => n9713, ZN => n9406);
   U12540 : XNOR2_X1 port map( A => n9894, B => n10382, ZN => n9403);
   U12541 : XNOR2_X1 port map( A => n9404, B => n9403, ZN => n9405);
   U12542 : NAND2_X1 port map( A1 => n9559, A2 => n10995, ZN => n9411);
   U12543 : XNOR2_X1 port map( A => n9869, B => n10261, ZN => n10036);
   U12544 : XNOR2_X1 port map( A => n10036, B => n9407, ZN => n9410);
   U12545 : XNOR2_X1 port map( A => n10421, B => n2221, ZN => n9408);
   U12546 : INV_X1 port map( A => n9794, ZN => n9458);
   U12547 : XNOR2_X1 port map( A => n20608, B => n19746, ZN => n9733);
   U12548 : XNOR2_X1 port map( A => n9408, B => n9733, ZN => n9409);
   U12549 : XNOR2_X1 port map( A => n9415, B => n10321, ZN => n9419);
   U12550 : XNOR2_X1 port map( A => n9416, B => n9417, ZN => n9418);
   U12551 : XNOR2_X2 port map( A => n9419, B => n9418, ZN => n11278);
   U12552 : INV_X1 port map( A => n11278, ZN => n10688);
   U12553 : XNOR2_X1 port map( A => n9420, B => n10261, ZN => n9422);
   U12554 : INV_X1 port map( A => n9421, ZN => n10233);
   U12555 : XNOR2_X1 port map( A => n9422, B => n10233, ZN => n9425);
   U12556 : XNOR2_X1 port map( A => n10229, B => n9669, ZN => n10342);
   U12557 : XNOR2_X1 port map( A => n9937, B => n2164, ZN => n9423);
   U12558 : XNOR2_X1 port map( A => n10342, B => n9423, ZN => n9424);
   U12559 : INV_X1 port map( A => n9861, ZN => n9426);
   U12560 : XNOR2_X1 port map( A => n9426, B => n10558, ZN => n10588);
   U12561 : XNOR2_X1 port map( A => n9648, B => n10349, ZN => n9427);
   U12562 : XNOR2_X1 port map( A => n9427, B => n10350, ZN => n9944);
   U12563 : XNOR2_X1 port map( A => n9697, B => n9856, ZN => n10334);
   U12564 : XNOR2_X1 port map( A => n10334, B => n10201, ZN => n9431);
   U12565 : XNOR2_X1 port map( A => n9432, B => n9431, ZN => n11413);
   U12566 : INV_X1 port map( A => n11413, ZN => n9547);
   U12567 : INV_X1 port map( A => n10248, ZN => n9846);
   U12568 : XNOR2_X1 port map( A => n9846, B => n9692, ZN => n10371);
   U12569 : XNOR2_X1 port map( A => n10296, B => n19760, ZN => n9661);
   U12570 : XNOR2_X1 port map( A => n9842, B => n18065, ZN => n9433);
   U12571 : XNOR2_X1 port map( A => n9661, B => n9433, ZN => n9434);
   U12572 : XNOR2_X1 port map( A => n10257, B => n9434, ZN => n9435);
   U12573 : XNOR2_X1 port map( A => n9435, B => n10371, ZN => n11411);
   U12574 : NAND2_X1 port map( A1 => n11276, A2 => n11411, ZN => n9444);
   U12575 : XNOR2_X1 port map( A => n10210, B => n10150, ZN => n9438);
   U12576 : INV_X1 port map( A => n10273, ZN => n9436);
   U12577 : XNOR2_X1 port map( A => n9436, B => n2394, ZN => n9437);
   U12578 : XNOR2_X1 port map( A => n9438, B => n9437, ZN => n9441);
   U12579 : XNOR2_X1 port map( A => n928, B => n9635, ZN => n9440);
   U12580 : INV_X1 port map( A => n10360, ZN => n9439);
   U12581 : XNOR2_X1 port map( A => n9441, B => n926, ZN => n9545);
   U12582 : INV_X1 port map( A => n9545, ZN => n11408);
   U12583 : OAI21_X1 port map( B1 => n11408, B2 => n11277, A => n11413, ZN => 
                           n9442);
   U12584 : NAND2_X1 port map( A1 => n9442, A2 => n19851, ZN => n9443);
   U12585 : NOR2_X1 port map( A1 => n11841, A2 => n11674, ZN => n9543);
   U12586 : XNOR2_X1 port map( A => n9691, B => n9817, ZN => n10508);
   U12587 : XNOR2_X1 port map( A => n9445, B => n10508, ZN => n9450);
   U12588 : INV_X1 port map( A => n9446, ZN => n9448);
   U12589 : XNOR2_X1 port map( A => n9844, B => n2307, ZN => n9447);
   U12590 : XNOR2_X1 port map( A => n9448, B => n9447, ZN => n9449);
   U12591 : XNOR2_X1 port map( A => n9450, B => n9449, ZN => n11011);
   U12592 : XNOR2_X1 port map( A => n9868, B => n2280, ZN => n9457);
   U12593 : XNOR2_X1 port map( A => n9457, B => n9456, ZN => n9461);
   U12594 : XNOR2_X1 port map( A => n9458, B => n9668, ZN => n10475);
   U12595 : XNOR2_X1 port map( A => n10475, B => n9459, ZN => n9460);
   U12597 : XNOR2_X1 port map( A => n10072, B => n2079, ZN => n9463);
   U12598 : XNOR2_X1 port map( A => n10481, B => n9463, ZN => n9467);
   U12599 : XNOR2_X1 port map( A => n9464, B => n9465, ZN => n9466);
   U12600 : XNOR2_X1 port map( A => n9467, B => n9466, ZN => n9548);
   U12601 : NOR2_X1 port map( A1 => n10953, A2 => n10952, ZN => n11013);
   U12602 : INV_X1 port map( A => n9812, ZN => n9468);
   U12603 : XNOR2_X1 port map( A => n9468, B => n9685, ZN => n10501);
   U12604 : XNOR2_X1 port map( A => n10501, B => n9469, ZN => n9474);
   U12605 : INV_X1 port map( A => n9470, ZN => n9472);
   U12606 : XNOR2_X1 port map( A => n9862, B => n17060, ZN => n9471);
   U12607 : XNOR2_X1 port map( A => n9472, B => n9471, ZN => n9473);
   U12610 : XNOR2_X1 port map( A => n9879, B => n610, ZN => n9475);
   U12611 : XNOR2_X1 port map( A => n9476, B => n9475, ZN => n9478);
   U12612 : INV_X1 port map( A => n9551, ZN => n11147);
   U12613 : XNOR2_X1 port map( A => n9923, B => n10114, ZN => n9479);
   U12614 : XNOR2_X1 port map( A => n9479, B => n9480, ZN => n9484);
   U12615 : XNOR2_X1 port map( A => n9922, B => n10570, ZN => n9482);
   U12616 : INV_X1 port map( A => n621, ZN => n18355);
   U12617 : XNOR2_X1 port map( A => n9777, B => n18355, ZN => n9481);
   U12618 : XNOR2_X1 port map( A => n9482, B => n9481, ZN => n9483);
   U12619 : XNOR2_X1 port map( A => n9484, B => n9483, ZN => n11149);
   U12620 : INV_X1 port map( A => n11149, ZN => n10951);
   U12621 : NAND3_X1 port map( A1 => n11016, A2 => n10952, A3 => n10951, ZN => 
                           n9485);
   U12622 : NOR2_X1 port map( A1 => n11175, A2 => n9351, ZN => n10657);
   U12623 : INV_X1 port map( A => n10657, ZN => n10912);
   U12624 : NAND2_X1 port map( A1 => n11174, A2 => n10962, ZN => n9487);
   U12627 : NAND2_X1 port map( A1 => n11175, A2 => n11178, ZN => n9488);
   U12628 : OAI22_X1 port map( A1 => n9488, A2 => n11176, B1 => n11177, B2 => 
                           n11174, ZN => n9489);
   U12629 : NOR2_X1 port map( A1 => n11161, A2 => n10649, ZN => n11157);
   U12630 : INV_X1 port map( A => n11157, ZN => n9495);
   U12631 : INV_X1 port map( A => n11156, ZN => n9494);
   U12632 : NAND2_X1 port map( A1 => n10649, A2 => n11159, ZN => n9493);
   U12633 : NAND3_X1 port map( A1 => n9495, A2 => n9494, A3 => n9493, ZN => 
                           n9497);
   U12634 : OAI211_X1 port map( C1 => n11158, C2 => n11160, A => n11155, B => 
                           n11159, ZN => n9496);
   U12635 : INV_X1 port map( A => n9499, ZN => n9501);
   U12636 : XNOR2_X1 port map( A => n9500, B => n10265, ZN => n10524);
   U12637 : XNOR2_X1 port map( A => n10524, B => n9501, ZN => n9505);
   U12638 : XNOR2_X1 port map( A => n9667, B => n16242, ZN => n9502);
   U12639 : XNOR2_X1 port map( A => n9503, B => n9502, ZN => n9504);
   U12640 : INV_X1 port map( A => n10274, ZN => n9506);
   U12641 : XNOR2_X1 port map( A => n9879, B => n9506, ZN => n10548);
   U12642 : XNOR2_X1 port map( A => n10548, B => n9507, ZN => n9511);
   U12643 : XNOR2_X1 port map( A => n9999, B => n18716, ZN => n9509);
   U12644 : XNOR2_X1 port map( A => n9509, B => n9508, ZN => n9510);
   U12645 : NOR2_X1 port map( A1 => n1721, A2 => n20366, ZN => n9517);
   U12646 : XNOR2_X1 port map( A => n9844, B => n19786, ZN => n10535);
   U12647 : XNOR2_X1 port map( A => n10535, B => n9512, ZN => n9516);
   U12648 : XNOR2_X1 port map( A => n10249, B => n2298, ZN => n9513);
   U12649 : XNOR2_X1 port map( A => n9514, B => n9513, ZN => n9515);
   U12650 : XNOR2_X1 port map( A => n9516, B => n9515, ZN => n10642);
   U12651 : XNOR2_X1 port map( A => n20176, B => n1996, ZN => n9519);
   U12652 : XNOR2_X1 port map( A => n9518, B => n9519, ZN => n9522);
   U12653 : XNOR2_X1 port map( A => n10303, B => n9777, ZN => n10568);
   U12654 : XNOR2_X1 port map( A => n10568, B => n9520, ZN => n9521);
   U12655 : XNOR2_X1 port map( A => n9524, B => n9523, ZN => n9525);
   U12656 : XNOR2_X1 port map( A => n9526, B => n9525, ZN => n9616);
   U12657 : NAND3_X1 port map( A1 => n9527, A2 => n18177, A3 => n9530, ZN => 
                           n9533);
   U12658 : INV_X1 port map( A => n18177, ZN => n9531);
   U12659 : NAND3_X1 port map( A1 => n9529, A2 => n9531, A3 => n9528, ZN => 
                           n9532);
   U12660 : XNOR2_X1 port map( A => n9534, B => n9983, ZN => n9536);
   U12661 : INV_X1 port map( A => n9535, ZN => n10180);
   U12662 : XNOR2_X1 port map( A => n10180, B => n10320, ZN => n9711);
   U12663 : XNOR2_X1 port map( A => n9711, B => n9536, ZN => n9541);
   U12664 : INV_X1 port map( A => n9538, ZN => n9539);
   U12665 : XNOR2_X1 port map( A => n10483, B => n9539, ZN => n9540);
   U12666 : INV_X1 port map( A => n13042, ZN => n9544);
   U12667 : XNOR2_X1 port map( A => n9544, B => n13070, ZN => n11801);
   U12669 : INV_X1 port map( A => n11000, ZN => n11005);
   U12670 : INV_X1 port map( A => n11952, ZN => n11827);
   U12671 : INV_X1 port map( A => n11011, ZN => n11153);
   U12672 : NOR2_X1 port map( A1 => n10953, A2 => n11153, ZN => n9550);
   U12673 : NOR2_X1 port map( A1 => n20470, A2 => n11147, ZN => n9549);
   U12674 : INV_X1 port map( A => n9548, ZN => n11009);
   U12675 : MUX2_X1 port map( A => n9550, B => n9549, S => n11009, Z => n9554);
   U12676 : NOR2_X1 port map( A1 => n9552, A2 => n11010, ZN => n9553);
   U12677 : NOR2_X1 port map( A1 => n11157, A2 => n9555, ZN => n9558);
   U12678 : NAND2_X1 port map( A1 => n10947, A2 => n10694, ZN => n11289);
   U12679 : INV_X1 port map( A => n9559, ZN => n10950);
   U12680 : NAND3_X1 port map( A1 => n10995, A2 => n11283, A3 => n11281, ZN => 
                           n9562);
   U12681 : INV_X1 port map( A => n10946, ZN => n11284);
   U12682 : NAND2_X1 port map( A1 => n11284, A2 => n11283, ZN => n10998);
   U12683 : NAND3_X1 port map( A1 => n19817, A2 => n10998, A3 => n9560, ZN => 
                           n9561);
   U12684 : XNOR2_X1 port map( A => n10506, B => n10186, ZN => n10533);
   U12685 : INV_X1 port map( A => n9568, ZN => n9569);
   U12686 : XNOR2_X1 port map( A => n10249, B => n1857, ZN => n9571);
   U12687 : XNOR2_X1 port map( A => n9571, B => n9843, ZN => n9572);
   U12688 : XNOR2_X1 port map( A => n10533, B => n9572, ZN => n9575);
   U12689 : XNOR2_X1 port map( A => n9960, B => n10445, ZN => n9573);
   U12693 : NAND2_X1 port map( A1 => n9577, A2 => n9576, ZN => n9581);
   U12694 : AOI21_X1 port map( B1 => n9581, B2 => n9580, A => n9579, ZN => 
                           n9584);
   U12695 : XNOR2_X1 port map( A => n10572, B => n1911, ZN => n9585);
   U12696 : XNOR2_X1 port map( A => n9585, B => n10016, ZN => n9586);
   U12697 : XNOR2_X1 port map( A => n10567, B => n10456, ZN => n10165);
   U12698 : XNOR2_X1 port map( A => n10514, B => n9587, ZN => n9588);
   U12699 : XNOR2_X1 port map( A => n10157, B => n10350, ZN => n9591);
   U12700 : XNOR2_X1 port map( A => n10498, B => n9589, ZN => n9590);
   U12701 : XNOR2_X1 port map( A => n9591, B => n9590, ZN => n9595);
   U12702 : XNOR2_X1 port map( A => n9994, B => n10431, ZN => n9593);
   U12703 : XNOR2_X1 port map( A => n10436, B => n17932, ZN => n9592);
   U12704 : XNOR2_X1 port map( A => n9593, B => n9592, ZN => n9594);
   U12705 : XNOR2_X1 port map( A => n9595, B => n9594, ZN => n11294);
   U12706 : INV_X1 port map( A => n11406, ZN => n9612);
   U12707 : INV_X1 port map( A => n10264, ZN => n9597);
   U12708 : XNOR2_X1 port map( A => n9597, B => n9667, ZN => n9598);
   U12709 : XNOR2_X1 port map( A => n9598, B => n10473, ZN => n9599);
   U12710 : XNOR2_X1 port map( A => n10179, B => n9600, ZN => n9800);
   U12711 : INV_X1 port map( A => n9987, ZN => n9601);
   U12712 : XNOR2_X1 port map( A => n9601, B => n10484, ZN => n9853);
   U12713 : XNOR2_X1 port map( A => n9853, B => n9800, ZN => n9604);
   U12714 : NOR2_X1 port map( A1 => n11292, A2 => n19506, ZN => n9610);
   U12715 : XNOR2_X1 port map( A => n9999, B => n10271, ZN => n9605);
   U12716 : XNOR2_X1 port map( A => n10358, B => n2100, ZN => n9607);
   U12717 : XNOR2_X1 port map( A => n878, B => n19717, ZN => n9606);
   U12718 : XNOR2_X1 port map( A => n9607, B => n9606, ZN => n9608);
   U12719 : INV_X1 port map( A => n11294, ZN => n11402);
   U12720 : OAI21_X1 port map( B1 => n11403, B2 => n11402, A => n10980, ZN => 
                           n9609);
   U12722 : MUX2_X1 port map( A => n9613, B => n981, S => n11951, Z => n9622);
   U12723 : INV_X1 port map( A => n10958, ZN => n9615);
   U12724 : NAND2_X1 port map( A1 => n9615, A2 => n9614, ZN => n9619);
   U12725 : NAND2_X1 port map( A1 => n11145, A2 => n11142, ZN => n9618);
   U12726 : INV_X1 port map( A => n10642, ZN => n11140);
   U12727 : AND3_X1 port map( A1 => n1749, A2 => n11140, A3 => n10701, ZN => 
                           n9617);
   U12728 : INV_X1 port map( A => n11830, ZN => n11953);
   U12729 : OAI21_X1 port map( B1 => n11659, B2 => n11953, A => n11828, ZN => 
                           n9620);
   U12730 : NOR2_X1 port map( A1 => n9620, A2 => n981, ZN => n9621);
   U12731 : INV_X1 port map( A => n10343, ZN => n9626);
   U12732 : XNOR2_X1 port map( A => n9626, B => n9625, ZN => n9631);
   U12733 : INV_X1 port map( A => n9937, ZN => n9627);
   U12734 : XNOR2_X1 port map( A => n10265, B => n9627, ZN => n9629);
   U12735 : XNOR2_X1 port map( A => n10425, B => n17804, ZN => n9628);
   U12736 : XNOR2_X1 port map( A => n9629, B => n9628, ZN => n9630);
   U12738 : INV_X1 port map( A => n9632, ZN => n9634);
   U12739 : XNOR2_X1 port map( A => n10461, B => n10079, ZN => n9633);
   U12740 : XNOR2_X1 port map( A => n9634, B => n9633, ZN => n9639);
   U12741 : XNOR2_X1 port map( A => n10213, B => n9635, ZN => n9637);
   U12742 : XNOR2_X1 port map( A => n10274, B => n19410, ZN => n9636);
   U12743 : XNOR2_X1 port map( A => n9637, B => n9636, ZN => n9638);
   U12744 : XNOR2_X1 port map( A => n9639, B => n9638, ZN => n10685);
   U12745 : NOR2_X1 port map( A1 => n20496, A2 => n12101, ZN => n9660);
   U12746 : XNOR2_X1 port map( A => n10303, B => n20672, ZN => n9640);
   U12747 : XNOR2_X1 port map( A => n10304, B => n9640, ZN => n9642);
   U12748 : XNOR2_X1 port map( A => n9967, B => n9922, ZN => n9641);
   U12749 : XNOR2_X1 port map( A => n9642, B => n9641, ZN => n9645);
   U12750 : XNOR2_X1 port map( A => n9644, B => n10105, ZN => n10337);
   U12751 : XNOR2_X1 port map( A => n10337, B => n9645, ZN => n10683);
   U12753 : XNOR2_X1 port map( A => n20156, B => n9648, ZN => n10438);
   U12754 : INV_X1 port map( A => n10438, ZN => n9649);
   U12755 : XNOR2_X1 port map( A => n10086, B => n9649, ZN => n9653);
   U12756 : XNOR2_X1 port map( A => n10281, B => n2123, ZN => n9650);
   U12757 : XNOR2_X1 port map( A => n9651, B => n9650, ZN => n9652);
   U12758 : INV_X1 port map( A => n10684, ZN => n10864);
   U12759 : INV_X1 port map( A => n10290, ZN => n9655);
   U12760 : XNOR2_X1 port map( A => n9947, B => n2192, ZN => n9654);
   U12761 : XNOR2_X1 port map( A => n9655, B => n9654, ZN => n9658);
   U12762 : XNOR2_X1 port map( A => n9894, B => n9986, ZN => n10318);
   U12763 : XNOR2_X1 port map( A => n9656, B => n10318, ZN => n9657);
   U12764 : XNOR2_X1 port map( A => n9658, B => n9657, ZN => n9666);
   U12765 : XNOR2_X1 port map( A => n10442, B => n9691, ZN => n9662);
   U12766 : XNOR2_X1 port map( A => n9662, B => n9661, ZN => n9665);
   U12768 : XNOR2_X1 port map( A => n19786, B => n17993, ZN => n9663);
   U12769 : XNOR2_X1 port map( A => n929, B => n9663, ZN => n9664);
   U12770 : XNOR2_X1 port map( A => n9664, B => n9665, ZN => n11380);
   U12771 : INV_X1 port map( A => n11380, ZN => n11275);
   U12772 : NAND2_X1 port map( A1 => n11275, A2 => n11383, ZN => n12100);
   U12773 : INV_X1 port map( A => n10422, ZN => n10605);
   U12774 : XNOR2_X1 port map( A => n9869, B => n10605, ZN => n10099);
   U12775 : XNOR2_X1 port map( A => n9667, B => n10421, ZN => n9975);
   U12776 : XNOR2_X1 port map( A => n10099, B => n9975, ZN => n9673);
   U12777 : XNOR2_X1 port map( A => n19853, B => n9668, ZN => n10138);
   U12778 : INV_X1 port map( A => n9670, ZN => n10174);
   U12779 : XNOR2_X1 port map( A => n10174, B => n642, ZN => n9671);
   U12780 : XNOR2_X1 port map( A => n10138, B => n9671, ZN => n9672);
   U12781 : XNOR2_X1 port map( A => n9673, B => n9672, ZN => n11328);
   U12782 : XNOR2_X1 port map( A => n10416, B => n9674, ZN => n9678);
   U12783 : XNOR2_X1 port map( A => n10220, B => n9983, ZN => n9676);
   U12784 : XNOR2_X1 port map( A => n9462, B => n2208, ZN => n9675);
   U12785 : XNOR2_X1 port map( A => n9676, B => n9675, ZN => n9677);
   U12786 : XNOR2_X1 port map( A => n9678, B => n9677, ZN => n11244);
   U12787 : XNOR2_X1 port map( A => n10077, B => n10126, ZN => n9680);
   U12788 : INV_X1 port map( A => n9679, ZN => n10465);
   U12789 : XNOR2_X1 port map( A => n10465, B => n9680, ZN => n9684);
   U12790 : XNOR2_X1 port map( A => n9999, B => n1057, ZN => n9682);
   U12791 : XNOR2_X1 port map( A => n928, B => n2423, ZN => n9681);
   U12792 : XNOR2_X1 port map( A => n9682, B => n9681, ZN => n9683);
   U12793 : XNOR2_X2 port map( A => n9684, B => n9683, ZN => n11376);
   U12794 : XNOR2_X1 port map( A => n10350, B => n9685, ZN => n10122);
   U12795 : INV_X1 port map( A => n10122, ZN => n9687);
   U12796 : XNOR2_X1 port map( A => n9994, B => n18420, ZN => n9686);
   U12797 : XNOR2_X1 port map( A => n9687, B => n9686, ZN => n9690);
   U12798 : XNOR2_X1 port map( A => n10430, B => n10087, ZN => n9688);
   U12799 : XNOR2_X1 port map( A => n10433, B => n9688, ZN => n9689);
   U12800 : MUX2_X1 port map( A => n11375, B => n10661, S => n11329, Z => 
                           n12363);
   U12801 : XNOR2_X1 port map( A => n9692, B => n9691, ZN => n10134);
   U12802 : XNOR2_X1 port map( A => n10444, B => n10134, ZN => n9696);
   U12803 : XNOR2_X1 port map( A => n10441, B => n10094, ZN => n9694);
   U12804 : XNOR2_X1 port map( A => n10249, B => n18338, ZN => n9693);
   U12805 : XNOR2_X1 port map( A => n9694, B => n9693, ZN => n9695);
   U12806 : XNOR2_X1 port map( A => n9696, B => n9695, ZN => n11373);
   U12807 : INV_X1 port map( A => n11373, ZN => n10856);
   U12808 : INV_X1 port map( A => n11376, ZN => n11332);
   U12809 : XNOR2_X1 port map( A => n9697, B => n9922, ZN => n10118);
   U12810 : INV_X1 port map( A => n10118, ZN => n9698);
   U12811 : XNOR2_X1 port map( A => n9698, B => n20176, ZN => n9708);
   U12812 : INV_X1 port map( A => n9700, ZN => n9699);
   U12813 : NAND2_X1 port map( A1 => n9699, A2 => n2203, ZN => n9704);
   U12814 : INV_X1 port map( A => n2203, ZN => n18909);
   U12815 : NAND2_X1 port map( A1 => n9703, A2 => n18909, ZN => n9702);
   U12816 : NAND2_X1 port map( A1 => n9700, A2 => n18909, ZN => n9701);
   U12817 : OAI211_X1 port map( C1 => n9704, C2 => n9703, A => n9702, B => 
                           n9701, ZN => n9705);
   U12818 : XNOR2_X1 port map( A => n9705, B => n10107, ZN => n9706);
   U12819 : XNOR2_X1 port map( A => n10454, B => n9706, ZN => n9707);
   U12820 : NAND2_X1 port map( A1 => n2858, A2 => n11330, ZN => n9709);
   U12821 : MUX2_X1 port map( A => n10662, B => n9709, S => n11244, Z => n12362
                           );
   U12822 : INV_X1 port map( A => n9710, ZN => n10031);
   U12823 : XNOR2_X1 port map( A => n10072, B => n10031, ZN => n10379);
   U12824 : XNOR2_X1 port map( A => n10379, B => n9711, ZN => n9715);
   U12825 : XNOR2_X1 port map( A => n9802, B => n2263, ZN => n9712);
   U12826 : XNOR2_X1 port map( A => n9713, B => n9712, ZN => n9714);
   U12827 : XNOR2_X2 port map( A => n9715, B => n9714, ZN => n11399);
   U12828 : INV_X1 port map( A => n10404, ZN => n9716);
   U12829 : XNOR2_X1 port map( A => n9716, B => n10402, ZN => n10131);
   U12830 : XNOR2_X1 port map( A => n10131, B => n9717, ZN => n9721);
   U12831 : XNOR2_X1 port map( A => n10252, B => n10367, ZN => n9719);
   U12832 : XNOR2_X1 port map( A => n19785, B => n484, ZN => n9718);
   U12833 : XNOR2_X1 port map( A => n9719, B => n9718, ZN => n9720);
   U12834 : XNOR2_X1 port map( A => n9721, B => n9720, ZN => n11297);
   U12835 : XNOR2_X1 port map( A => n10043, B => n10557, ZN => n10396);
   U12836 : XNOR2_X1 port map( A => n10396, B => n9722, ZN => n9726);
   U12837 : XNOR2_X1 port map( A => n10236, B => n1386, ZN => n9723);
   U12838 : XNOR2_X1 port map( A => n9724, B => n9723, ZN => n9725);
   U12839 : XNOR2_X1 port map( A => n9726, B => n9725, ZN => n10667);
   U12840 : INV_X1 port map( A => n10667, ZN => n11394);
   U12841 : INV_X1 port map( A => n9952, ZN => n9727);
   U12842 : XNOR2_X1 port map( A => n9727, B => n10551, ZN => n10125);
   U12843 : XNOR2_X1 port map( A => n10125, B => n9728, ZN => n9732);
   U12844 : XNOR2_X1 port map( A => n10359, B => n917, ZN => n9730);
   U12845 : XNOR2_X1 port map( A => n10274, B => n19158, ZN => n9729);
   U12846 : XNOR2_X1 port map( A => n9730, B => n9729, ZN => n9731);
   U12847 : NAND2_X1 port map( A1 => n11394, A2 => n11397, ZN => n9746);
   U12848 : XNOR2_X1 port map( A => n19767, B => n10339, ZN => n9734);
   U12849 : XNOR2_X1 port map( A => n9734, B => n9733, ZN => n9737);
   U12850 : XNOR2_X1 port map( A => n10037, B => n10526, ZN => n10376);
   U12851 : XNOR2_X1 port map( A => n10265, B => n538, ZN => n9735);
   U12852 : XNOR2_X1 port map( A => n10376, B => n9735, ZN => n9736);
   U12853 : XNOR2_X1 port map( A => n20161, B => n10052, ZN => n9739);
   U12854 : XNOR2_X1 port map( A => n9738, B => n9739, ZN => n9743);
   U12855 : XNOR2_X1 port map( A => n10388, B => n10203, ZN => n9741);
   U12856 : XNOR2_X1 port map( A => n10570, B => n347, ZN => n9740);
   U12857 : XNOR2_X1 port map( A => n9741, B => n9740, ZN => n9742);
   U12858 : XNOR2_X1 port map( A => n9743, B => n9742, ZN => n10986);
   U12859 : NAND2_X1 port map( A1 => n10667, A2 => n10986, ZN => n9744);
   U12860 : OAI21_X1 port map( B1 => n11395, B2 => n11399, A => n9744, ZN => 
                           n10985);
   U12861 : NAND2_X1 port map( A1 => n10985, A2 => n11401, ZN => n9745);
   U12863 : INV_X1 port map( A => n12009, ZN => n12510);
   U12864 : XNOR2_X1 port map( A => n9748, B => n620, ZN => n9749);
   U12865 : XNOR2_X1 port map( A => n20483, B => n9749, ZN => n9751);
   U12866 : XNOR2_X1 port map( A => n9750, B => n9751, ZN => n9753);
   U12867 : XNOR2_X1 port map( A => n10528, B => n10262, ZN => n9752);
   U12868 : XNOR2_X1 port map( A => n10137, B => n9752, ZN => n10477);
   U12869 : XNOR2_X1 port map( A => n9753, B => n10477, ZN => n11871);
   U12870 : XNOR2_X1 port map( A => n9754, B => n10482, ZN => n10540);
   U12871 : XNOR2_X1 port map( A => n9987, B => n18997, ZN => n9755);
   U12872 : XNOR2_X1 port map( A => n10540, B => n9755, ZN => n9758);
   U12873 : XNOR2_X1 port map( A => n20134, B => n10028, ZN => n10287);
   U12874 : XNOR2_X1 port map( A => n9756, B => n10287, ZN => n9757);
   U12876 : INV_X1 port map( A => n11303, ZN => n10862);
   U12879 : XNOR2_X1 port map( A => n9760, B => n10270, ZN => n10489);
   U12881 : XNOR2_X1 port map( A => n9761, B => n9902, ZN => n9763);
   U12882 : XNOR2_X1 port map( A => n9879, B => n878, ZN => n9762);
   U12883 : XNOR2_X1 port map( A => n9763, B => n9762, ZN => n9764);
   U12884 : XNOR2_X1 port map( A => n10489, B => n9764, ZN => n11389);
   U12886 : XNOR2_X1 port map( A => n10236, B => n18278, ZN => n9766);
   U12887 : INV_X1 port map( A => n9908, ZN => n9765);
   U12888 : XNOR2_X1 port map( A => n9766, B => n9765, ZN => n9768);
   U12889 : XNOR2_X1 port map( A => n9862, B => n10436, ZN => n9767);
   U12890 : XNOR2_X1 port map( A => n9768, B => n9767, ZN => n9770);
   U12891 : XNOR2_X1 port map( A => n10589, B => n10048, ZN => n10279);
   U12892 : INV_X1 port map( A => n9769, ZN => n10561);
   U12893 : XNOR2_X1 port map( A => n10279, B => n10561, ZN => n10503);
   U12895 : INV_X1 port map( A => n11866, ZN => n10990);
   U12896 : XNOR2_X1 port map( A => n9772, B => n9843, ZN => n9774);
   U12897 : INV_X1 port map( A => n9819, ZN => n10401);
   U12898 : XNOR2_X1 port map( A => n10401, B => n10612, ZN => n9775);
   U12899 : XNOR2_X1 port map( A => n9775, B => n19871, ZN => n10510);
   U12900 : NAND2_X1 port map( A1 => n11302, A2 => n19750, ZN => n10711);
   U12901 : INV_X1 port map( A => n9777, ZN => n9778);
   U12902 : INV_X1 port map( A => n9779, ZN => n9785);
   U12904 : AOI21_X1 port map( B1 => n19553, B2 => n9782, A => n9781, ZN => 
                           n9783);
   U12905 : OAI21_X1 port map( B1 => n9785, B2 => n19553, A => n9783, ZN => 
                           n9786);
   U12906 : XNOR2_X1 port map( A => n9786, B => n10054, ZN => n10517);
   U12907 : XNOR2_X1 port map( A => n10517, B => n9860, ZN => n9790);
   U12908 : INV_X1 port map( A => n10566, ZN => n10387);
   U12909 : INV_X1 port map( A => n10203, ZN => n9787);
   U12910 : XNOR2_X1 port map( A => n9926, B => n573, ZN => n9788);
   U12911 : XNOR2_X1 port map( A => n9789, B => n9790, ZN => n10709);
   U12912 : AOI21_X1 port map( B1 => n10711, B2 => n20517, A => n20601, ZN => 
                           n9791);
   U12913 : MUX2_X1 port map( A => n12008, B => n12510, S => n12508, Z => n9887
                           );
   U12914 : XNOR2_X1 port map( A => n10171, B => n10472, ZN => n10525);
   U12915 : XNOR2_X1 port map( A => n10525, B => n9974, ZN => n9798);
   U12918 : XNOR2_X1 port map( A => n10229, B => n18396, ZN => n9795);
   U12919 : XNOR2_X1 port map( A => n9796, B => n9795, ZN => n9797);
   U12920 : XNOR2_X1 port map( A => n10482, B => n9799, ZN => n9801);
   U12921 : INV_X1 port map( A => n9800, ZN => n10541);
   U12922 : XNOR2_X1 port map( A => n10541, B => n9801, ZN => n9805);
   U12923 : XNOR2_X1 port map( A => n9854, B => n9802, ZN => n10223);
   U12924 : XNOR2_X1 port map( A => n10289, B => n19102, ZN => n9803);
   U12925 : XNOR2_X1 port map( A => n9803, B => n10223, ZN => n9804);
   U12926 : XNOR2_X1 port map( A => n9805, B => n9804, ZN => n10194);
   U12927 : INV_X1 port map( A => n10194, ZN => n11337);
   U12928 : XNOR2_X1 port map( A => n10203, B => n9923, ZN => n9806);
   U12929 : XNOR2_X1 port map( A => n10165, B => n9806, ZN => n9810);
   U12930 : XNOR2_X1 port map( A => n10387, B => n10205, ZN => n9808);
   U12931 : XNOR2_X1 port map( A => n10572, B => n457, ZN => n9807);
   U12932 : XNOR2_X1 port map( A => n9808, B => n9807, ZN => n9809);
   U12933 : XNOR2_X1 port map( A => n9809, B => n9810, ZN => n10673);
   U12934 : XNOR2_X1 port map( A => n10497, B => n10157, ZN => n10559);
   U12935 : INV_X1 port map( A => n9996, ZN => n9811);
   U12936 : XNOR2_X1 port map( A => n9811, B => n10559, ZN => n9816);
   U12937 : XNOR2_X1 port map( A => n9812, B => n10349, ZN => n9814);
   U12938 : XNOR2_X1 port map( A => n10236, B => n18863, ZN => n9813);
   U12939 : XNOR2_X1 port map( A => n9814, B => n9813, ZN => n9815);
   U12940 : INV_X1 port map( A => n9830, ZN => n11264);
   U12941 : XNOR2_X1 port map( A => n10252, B => n9817, ZN => n9818);
   U12942 : XNOR2_X1 port map( A => n10533, B => n9818, ZN => n9823);
   U12943 : XNOR2_X1 port map( A => n10248, B => n18478, ZN => n9821);
   U12944 : INV_X1 port map( A => n10445, ZN => n9820);
   U12945 : XNOR2_X1 port map( A => n9819, B => n9820, ZN => n10011);
   U12946 : XNOR2_X1 port map( A => n9821, B => n10011, ZN => n9822);
   U12947 : INV_X1 port map( A => n11267, ZN => n11343);
   U12948 : XNOR2_X1 port map( A => n9998, B => n10549, ZN => n9829);
   U12949 : XNOR2_X1 port map( A => n9824, B => n10360, ZN => n9827);
   U12950 : XNOR2_X1 port map( A => n918, B => n18208, ZN => n9826);
   U12951 : XNOR2_X1 port map( A => n9827, B => n9826, ZN => n9828);
   U12952 : MUX2_X1 port map( A => n20505, B => n20476, S => n19606, Z => n9840
                           );
   U12953 : NAND3_X1 port map( A1 => n9837, A2 => n9836, A3 => n20505, ZN => 
                           n9839);
   U12954 : XNOR2_X1 port map( A => n9842, B => n9841, ZN => n10611);
   U12955 : XNOR2_X1 port map( A => n10613, B => n9843, ZN => n10010);
   U12956 : XNOR2_X1 port map( A => n10010, B => n10611, ZN => n9850);
   U12957 : INV_X1 port map( A => n9844, ZN => n9845);
   U12958 : XNOR2_X1 port map( A => n9845, B => n10094, ZN => n9848);
   U12959 : XNOR2_X1 port map( A => n9846, B => n19321, ZN => n9847);
   U12960 : XNOR2_X1 port map( A => n9848, B => n9847, ZN => n9849);
   U12961 : INV_X1 port map( A => n11365, ZN => n10676);
   U12962 : INV_X1 port map( A => n10382, ZN => n9851);
   U12963 : XNOR2_X1 port map( A => n9851, B => n10542, ZN => n9852);
   U12964 : XNOR2_X1 port map( A => n9854, B => n16424, ZN => n9855);
   U12965 : XNOR2_X1 port map( A => n10598, B => n10205, ZN => n9858);
   U12966 : XNOR2_X1 port map( A => n10107, B => n2424, ZN => n9857);
   U12967 : XNOR2_X1 port map( A => n9857, B => n9858, ZN => n9859);
   U12968 : XNOR2_X1 port map( A => n10571, B => n10163, ZN => n10600);
   U12969 : INV_X1 port map( A => n9883, ZN => n10852);
   U12970 : XNOR2_X1 port map( A => n10558, B => n10436, ZN => n9992);
   U12971 : XNOR2_X1 port map( A => n10498, B => n9861, ZN => n10158);
   U12973 : XNOR2_X1 port map( A => n9862, B => n2087, ZN => n9864);
   U12974 : XNOR2_X1 port map( A => n10087, B => n10349, ZN => n9863);
   U12976 : INV_X1 port map( A => n11234, ZN => n10851);
   U12977 : NOR2_X1 port map( A1 => n10852, A2 => n10851, ZN => n9874);
   U12978 : XNOR2_X1 port map( A => n10229, B => Key(60), ZN => n9867);
   U12979 : XNOR2_X1 port map( A => n9867, B => n9868, ZN => n9871);
   U12980 : XNOR2_X1 port map( A => n9977, B => n9869, ZN => n9870);
   U12981 : XNOR2_X1 port map( A => n9871, B => n9870, ZN => n9873);
   U12982 : XNOR2_X1 port map( A => n20115, B => n10173, ZN => n9872);
   U12983 : XNOR2_X1 port map( A => n9872, B => n10473, ZN => n10609);
   U12984 : XNOR2_X1 port map( A => n9873, B => n10609, ZN => n10675);
   U12985 : BUF_X2 port map( A => n10675, Z => n11230);
   U12986 : INV_X1 port map( A => n10490, ZN => n9876);
   U12987 : XNOR2_X1 port map( A => n9876, B => n10150, ZN => n10580);
   U12988 : XNOR2_X1 port map( A => n19945, B => n10360, ZN => n9877);
   U12990 : INV_X1 port map( A => n10578, ZN => n10550);
   U12991 : XNOR2_X1 port map( A => n878, B => n10550, ZN => n10004);
   U12992 : XNOR2_X1 port map( A => n9879, B => n17466, ZN => n9880);
   U12994 : INV_X1 port map( A => n11231, ZN => n10854);
   U12995 : INV_X1 port map( A => n12509, ZN => n11834);
   U12996 : NAND2_X1 port map( A1 => n11834, A2 => n12359, ZN => n9885);
   U12997 : XNOR2_X1 port map( A => n13746, B => n12696, ZN => n13444);
   U12998 : XNOR2_X1 port map( A => n11801, B => n13444, ZN => n10634);
   U12999 : XNOR2_X1 port map( A => n10171, B => n10262, ZN => n9889);
   U13000 : XNOR2_X1 port map( A => n10231, B => n2216, ZN => n9888);
   U13001 : XNOR2_X1 port map( A => n9889, B => n9888, ZN => n9893);
   U13002 : XNOR2_X1 port map( A => n872, B => n20484, ZN => n10373);
   U13003 : INV_X1 port map( A => n10373, ZN => n9891);
   U13004 : XNOR2_X1 port map( A => n9891, B => n10475, ZN => n9892);
   U13006 : INV_X1 port map( A => n9894, ZN => n10222);
   U13007 : XNOR2_X1 port map( A => n10222, B => n2420, ZN => n9895);
   U13008 : XNOR2_X1 port map( A => n20228, B => n9895, ZN => n9900);
   U13009 : XNOR2_X1 port map( A => n20134, B => n10320, ZN => n10381);
   U13010 : XNOR2_X1 port map( A => n19839, B => n10028, ZN => n9898);
   U13011 : XNOR2_X1 port map( A => n10381, B => n9898, ZN => n9899);
   U13012 : XNOR2_X1 port map( A => n9900, B => n9899, ZN => n9919);
   U13013 : INV_X1 port map( A => n10359, ZN => n9901);
   U13014 : XNOR2_X1 port map( A => n9901, B => n9902, ZN => n10410);
   U13015 : XNOR2_X1 port map( A => n19829, B => n10410, ZN => n9907);
   U13016 : XNOR2_X1 port map( A => n10151, B => n10270, ZN => n9905);
   U13017 : XNOR2_X1 port map( A => n10213, B => n18006, ZN => n9904);
   U13018 : XNOR2_X1 port map( A => n9905, B => n9904, ZN => n9906);
   U13019 : XNOR2_X1 port map( A => n10395, B => n10501, ZN => n9912);
   U13020 : XNOR2_X1 port map( A => n19990, B => n645, ZN => n9909);
   U13021 : XNOR2_X1 port map( A => n9910, B => n9909, ZN => n9911);
   U13022 : XNOR2_X1 port map( A => n9912, B => n9911, ZN => n11216);
   U13023 : XNOR2_X1 port map( A => n10186, B => n19871, ZN => n9914);
   U13024 : XNOR2_X1 port map( A => n9914, B => n10508, ZN => n9918);
   U13025 : XNOR2_X1 port map( A => n10298, B => n10367, ZN => n10403);
   U13026 : INV_X1 port map( A => n10403, ZN => n9916);
   U13027 : XNOR2_X1 port map( A => n10247, B => n18090, ZN => n9915);
   U13028 : XNOR2_X1 port map( A => n9916, B => n9915, ZN => n9917);
   U13029 : XNOR2_X1 port map( A => n9918, B => n9917, ZN => n11475);
   U13030 : NAND2_X1 port map( A1 => n9920, A2 => n11475, ZN => n9921);
   U13031 : XNOR2_X1 port map( A => n10567, B => n10204, ZN => n9925);
   U13032 : XNOR2_X1 port map( A => n9923, B => n9922, ZN => n10515);
   U13033 : INV_X1 port map( A => n10515, ZN => n9924);
   U13034 : XNOR2_X1 port map( A => n9925, B => n9924, ZN => n9929);
   U13035 : XNOR2_X1 port map( A => n9926, B => n10332, ZN => n10391);
   U13036 : XNOR2_X1 port map( A => n10054, B => n2417, ZN => n9927);
   U13037 : XNOR2_X1 port map( A => n10391, B => n9927, ZN => n9928);
   U13038 : NAND2_X1 port map( A1 => n9930, A2 => n11079, ZN => n12498);
   U13039 : INV_X1 port map( A => n10755, ZN => n11522);
   U13040 : OAI21_X1 port map( B1 => n11528, B2 => n11530, A => n19999, ZN => 
                           n9931);
   U13041 : XNOR2_X1 port map( A => n10422, B => n9935, ZN => n9936);
   U13042 : XNOR2_X1 port map( A => n9936, B => n10342, ZN => n9940);
   U13043 : XNOR2_X1 port map( A => n9937, B => n9978, ZN => n9938);
   U13044 : XNOR2_X1 port map( A => n10473, B => n9938, ZN => n9939);
   U13045 : XNOR2_X1 port map( A => n10043, B => n19018, ZN => n9942);
   U13046 : INV_X1 port map( A => n9991, ZN => n9941);
   U13047 : XNOR2_X1 port map( A => n9942, B => n9941, ZN => n9943);
   U13048 : XNOR2_X1 port map( A => n10088, B => n10498, ZN => n10587);
   U13049 : XNOR2_X1 port map( A => n9943, B => n10587, ZN => n9945);
   U13050 : XNOR2_X1 port map( A => n9945, B => n9944, ZN => n10883);
   U13051 : INV_X1 port map( A => n10484, ZN => n9946);
   U13052 : XNOR2_X1 port map( A => n10031, B => n9986, ZN => n9949);
   U13053 : XNOR2_X1 port map( A => n9947, B => n17089, ZN => n9948);
   U13054 : XNOR2_X1 port map( A => n9949, B => n9948, ZN => n9950);
   U13055 : XNOR2_X1 port map( A => n9952, B => n10579, ZN => n9955);
   U13056 : XNOR2_X1 port map( A => n19717, B => n17535, ZN => n9953);
   U13057 : XNOR2_X1 port map( A => n9953, B => n10079, ZN => n9954);
   U13058 : XNOR2_X1 port map( A => n9954, B => n9955, ZN => n9956);
   U13059 : XNOR2_X1 port map( A => n9957, B => n20211, ZN => n9959);
   U13060 : XNOR2_X1 port map( A => n10008, B => n2233, ZN => n9958);
   U13061 : XNOR2_X1 port map( A => n9958, B => n9959, ZN => n9962);
   U13062 : XNOR2_X1 port map( A => n9960, B => n10404, ZN => n9961);
   U13063 : XNOR2_X1 port map( A => n9962, B => n9961, ZN => n9964);
   U13064 : INV_X1 port map( A => n10371, ZN => n9963);
   U13065 : NAND2_X1 port map( A1 => n11182, A2 => n10882, ZN => n9972);
   U13066 : XNOR2_X1 port map( A => n10514, B => n10105, ZN => n9966);
   U13067 : XNOR2_X1 port map( A => n10594, B => n10388, ZN => n9965);
   U13068 : XNOR2_X1 port map( A => n9965, B => n9966, ZN => n9970);
   U13069 : XNOR2_X1 port map( A => n9967, B => n2305, ZN => n9968);
   U13070 : XNOR2_X1 port map( A => n10334, B => n9968, ZN => n9969);
   U13071 : NAND2_X1 port map( A1 => n11566, A2 => n11466, ZN => n9971);
   U13072 : MUX2_X1 port map( A => n9972, B => n9971, S => n11568, Z => n9973);
   U13073 : INV_X1 port map( A => n9974, ZN => n9976);
   U13074 : XNOR2_X1 port map( A => n9976, B => n9975, ZN => n9982);
   U13075 : XNOR2_X1 port map( A => n9977, B => n20115, ZN => n9980);
   U13076 : XNOR2_X1 port map( A => n9978, B => n2306, ZN => n9979);
   U13077 : XNOR2_X1 port map( A => n9979, B => n9980, ZN => n9981);
   U13078 : XNOR2_X1 port map( A => n10542, B => n9983, ZN => n10618);
   U13079 : INV_X1 port map( A => n9984, ZN => n9985);
   U13080 : XNOR2_X1 port map( A => n10618, B => n9985, ZN => n9990);
   U13081 : XNOR2_X1 port map( A => n10219, B => n9986, ZN => n9989);
   U13082 : XNOR2_X1 port map( A => n9987, B => n16030, ZN => n9988);
   U13083 : NAND2_X1 port map( A1 => n11515, A2 => n10742, ZN => n11575);
   U13084 : XNOR2_X1 port map( A => n10240, B => n9991, ZN => n9993);
   U13085 : XNOR2_X1 port map( A => n9992, B => n9993, ZN => n9997);
   U13086 : XNOR2_X1 port map( A => n9994, B => n19205, ZN => n9995);
   U13087 : INV_X1 port map( A => n9998, ZN => n10001);
   U13088 : XNOR2_X1 port map( A => n9999, B => n10079, ZN => n10000);
   U13089 : XNOR2_X1 port map( A => n10001, B => n10000, ZN => n10006);
   U13090 : INV_X1 port map( A => n10002, ZN => n10214);
   U13091 : XNOR2_X1 port map( A => n10214, B => n2455, ZN => n10003);
   U13092 : XNOR2_X1 port map( A => n10004, B => n10003, ZN => n10005);
   U13094 : XNOR2_X1 port map( A => n10254, B => n10008, ZN => n10009);
   U13095 : XNOR2_X1 port map( A => n10010, B => n10009, ZN => n10015);
   U13096 : INV_X1 port map( A => n10011, ZN => n10013);
   U13097 : XNOR2_X1 port map( A => n10249, B => n18726, ZN => n10012);
   U13098 : XNOR2_X1 port map( A => n10013, B => n10012, ZN => n10014);
   U13101 : XNOR2_X1 port map( A => n10016, B => n20176, ZN => n10018);
   U13102 : XNOR2_X1 port map( A => n10018, B => n10017, ZN => n10022);
   U13103 : XNOR2_X1 port map( A => n10105, B => n19806, ZN => n10020);
   U13104 : XNOR2_X1 port map( A => n10571, B => n1148, ZN => n10019);
   U13105 : XNOR2_X1 port map( A => n10020, B => n10019, ZN => n10021);
   U13106 : XNOR2_X1 port map( A => n10022, B => n10021, ZN => n11510);
   U13107 : NOR2_X1 port map( A1 => n11510, A2 => n11514, ZN => n10740);
   U13108 : INV_X1 port map( A => n12498, ZN => n12497);
   U13109 : XNOR2_X1 port map( A => n10404, B => n19457, ZN => n10024);
   U13110 : XNOR2_X1 port map( A => n10406, B => n10024, ZN => n10025);
   U13111 : XNOR2_X1 port map( A => n10026, B => n10442, ZN => n10370);
   U13112 : XNOR2_X1 port map( A => n10028, B => n10382, ZN => n10029);
   U13113 : XNOR2_X1 port map( A => n10220, B => n10030, ZN => n10033);
   U13114 : XNOR2_X1 port map( A => n10031, B => n18308, ZN => n10032);
   U13115 : XNOR2_X1 port map( A => n10033, B => n10032, ZN => n10034);
   U13116 : XNOR2_X1 port map( A => n10035, B => n10034, ZN => n10060);
   U13117 : INV_X1 port map( A => n10060, ZN => n11482);
   U13118 : INV_X1 port map( A => n10036, ZN => n10374);
   U13119 : XNOR2_X1 port map( A => n10037, B => n10262, ZN => n10038);
   U13120 : XNOR2_X1 port map( A => n10374, B => n10038, ZN => n10042);
   U13121 : XNOR2_X1 port map( A => n10174, B => n456, ZN => n10040);
   U13122 : XNOR2_X1 port map( A => n10340, B => n10040, ZN => n10041);
   U13123 : INV_X1 port map( A => n10043, ZN => n10044);
   U13124 : XNOR2_X1 port map( A => n10044, B => n10430, ZN => n10047);
   U13125 : XNOR2_X1 port map( A => n10347, B => n10047, ZN => n10051);
   U13126 : XNOR2_X1 port map( A => n19990, B => n17989, ZN => n10049);
   U13127 : XNOR2_X1 port map( A => n10397, B => n10049, ZN => n10050);
   U13128 : XNOR2_X1 port map( A => n10051, B => n10050, ZN => n10745);
   U13129 : XNOR2_X1 port map( A => n10052, B => n10388, ZN => n10115);
   U13130 : INV_X1 port map( A => n10392, ZN => n10053);
   U13131 : XNOR2_X1 port map( A => n10115, B => n10053, ZN => n10058);
   U13132 : XNOR2_X1 port map( A => n10114, B => n10166, ZN => n10458);
   U13133 : INV_X1 port map( A => n10458, ZN => n10056);
   U13134 : XNOR2_X1 port map( A => n10054, B => n632, ZN => n10055);
   U13135 : XNOR2_X1 port map( A => n10056, B => n10055, ZN => n10057);
   U13136 : XNOR2_X1 port map( A => n10058, B => n10057, ZN => n10896);
   U13137 : NAND2_X1 port map( A1 => n19897, A2 => n11480, ZN => n10748);
   U13138 : NAND2_X1 port map( A1 => n11073, A2 => n10748, ZN => n10066);
   U13139 : INV_X1 port map( A => n10745, ZN => n11481);
   U13140 : XNOR2_X1 port map( A => n10409, B => n10356, ZN => n10065);
   U13141 : XNOR2_X1 port map( A => n1057, B => n10270, ZN => n10063);
   U13142 : XNOR2_X1 port map( A => n9952, B => n17787, ZN => n10062);
   U13143 : XNOR2_X1 port map( A => n10063, B => n10062, ZN => n10064);
   U13144 : NAND2_X1 port map( A1 => n11481, A2 => n10897, ZN => n11479);
   U13145 : NAND2_X1 port map( A1 => n10066, A2 => n11479, ZN => n10067);
   U13146 : INV_X1 port map( A => n10761, ZN => n10889);
   U13147 : INV_X1 port map( A => n11546, ZN => n11547);
   U13148 : NAND2_X1 port map( A1 => n11546, A2 => n11550, ZN => n10069);
   U13149 : NAND3_X1 port map( A1 => n1859, A2 => n12005, A3 => n12502, ZN => 
                           n10070);
   U13150 : XNOR2_X1 port map( A => n19818, B => n18284, ZN => n10074);
   U13151 : XNOR2_X1 port map( A => n10072, B => n10382, ZN => n10073);
   U13152 : XNOR2_X1 port map( A => n10074, B => n10073, ZN => n10076);
   U13153 : XNOR2_X1 port map( A => n10318, B => n10417, ZN => n10075);
   U13154 : INV_X1 port map( A => n10112, ZN => n11125);
   U13155 : INV_X1 port map( A => n19945, ZN => n10078);
   U13156 : XNOR2_X1 port map( A => n10078, B => n10579, ZN => n10081);
   U13157 : INV_X1 port map( A => n10213, ZN => n10080);
   U13158 : XNOR2_X1 port map( A => n10080, B => n10079, ZN => n10357);
   U13159 : XNOR2_X1 port map( A => n10357, B => n10081, ZN => n10084);
   U13160 : XNOR2_X1 port map( A => n10551, B => n17170, ZN => n10082);
   U13161 : XNOR2_X1 port map( A => n10462, B => n10082, ZN => n10083);
   U13162 : XNOR2_X1 port map( A => n10557, B => n10087, ZN => n10090);
   U13163 : XNOR2_X1 port map( A => n10088, B => n18011, ZN => n10089);
   U13164 : XNOR2_X1 port map( A => n10090, B => n10089, ZN => n10091);
   U13165 : MUX2_X1 port map( A => n11125, B => n10814, S => n1317, Z => n10104
                           );
   U13166 : XNOR2_X1 port map( A => n20210, B => n1904, ZN => n10093);
   U13167 : INV_X1 port map( A => n929, ZN => n10092);
   U13168 : XNOR2_X1 port map( A => n10093, B => n10092, ZN => n10097);
   U13169 : XNOR2_X1 port map( A => n10094, B => n10402, ZN => n10095);
   U13170 : XNOR2_X1 port map( A => n10447, B => n10095, ZN => n10096);
   U13171 : INV_X1 port map( A => n11358, ZN => n10103);
   U13173 : XNOR2_X1 port map( A => n20456, B => n10099, ZN => n10102);
   U13174 : XNOR2_X1 port map( A => n10526, B => n649, ZN => n10100);
   U13175 : XNOR2_X1 port map( A => n10343, B => n10100, ZN => n10101);
   U13176 : XNOR2_X1 port map( A => n10453, B => n10106, ZN => n10111);
   U13177 : XNOR2_X1 port map( A => n10204, B => n10570, ZN => n10109);
   U13178 : XNOR2_X1 port map( A => n10107, B => n1869, ZN => n10108);
   U13179 : XNOR2_X1 port map( A => n10109, B => n10108, ZN => n10110);
   U13180 : XNOR2_X1 port map( A => n10111, B => n10110, ZN => n11356);
   U13181 : INV_X1 port map( A => n11356, ZN => n11127);
   U13182 : NAND2_X1 port map( A1 => n11127, A2 => n10813, ZN => n10113);
   U13183 : XNOR2_X1 port map( A => n10595, B => n10114, ZN => n10116);
   U13184 : XNOR2_X1 port map( A => n10116, B => n10115, ZN => n10120);
   U13185 : XNOR2_X1 port map( A => n10570, B => n18768, ZN => n10117);
   U13186 : XNOR2_X1 port map( A => n10118, B => n10117, ZN => n10119);
   U13187 : XNOR2_X1 port map( A => n10120, B => n10119, ZN => n11238);
   U13188 : INV_X1 port map( A => n11238, ZN => n11355);
   U13189 : XNOR2_X1 port map( A => n10589, B => n19436, ZN => n10121);
   U13190 : XNOR2_X1 port map( A => n10396, B => n10121, ZN => n10124);
   U13191 : XNOR2_X1 port map( A => n10347, B => n10122, ZN => n10123);
   U13192 : XNOR2_X1 port map( A => n10123, B => n10124, ZN => n10779);
   U13193 : INV_X1 port map( A => n10779, ZN => n11239);
   U13194 : XNOR2_X1 port map( A => n10126, B => n10358, ZN => n10128);
   U13195 : XNOR2_X1 port map( A => n10582, B => n2413, ZN => n10127);
   U13196 : XNOR2_X1 port map( A => n10128, B => n10127, ZN => n10129);
   U13197 : XNOR2_X1 port map( A => n10130, B => n10129, ZN => n11240);
   U13198 : INV_X1 port map( A => n10131, ZN => n10133);
   U13199 : XNOR2_X1 port map( A => n10612, B => n18988, ZN => n10132);
   U13200 : XNOR2_X1 port map( A => n10133, B => n10132, ZN => n10136);
   U13201 : XNOR2_X1 port map( A => n10134, B => n10370, ZN => n10135);
   U13202 : INV_X1 port map( A => n11349, ZN => n11055);
   U13203 : INV_X1 port map( A => n10604, ZN => n10137);
   U13204 : XNOR2_X1 port map( A => n10137, B => n2108, ZN => n10139);
   U13205 : XNOR2_X1 port map( A => n10139, B => n10138, ZN => n10141);
   U13206 : XNOR2_X1 port map( A => n10376, B => n10340, ZN => n10140);
   U13207 : XNOR2_X1 port map( A => n10140, B => n10141, ZN => n11347);
   U13208 : INV_X1 port map( A => n11347, ZN => n11350);
   U13209 : NAND2_X1 port map( A1 => n11347, A2 => n10798, ZN => n10142);
   U13210 : NAND2_X1 port map( A1 => n11060, A2 => n10142, ZN => n10148);
   U13211 : XNOR2_X1 port map( A => n10379, B => n10319, ZN => n10147);
   U13212 : XNOR2_X1 port map( A => n10286, B => n9462, ZN => n10145);
   U13213 : XNOR2_X1 port map( A => n10143, B => n18439, ZN => n10144);
   U13214 : XNOR2_X1 port map( A => n10145, B => n10144, ZN => n10146);
   U13215 : INV_X1 port map( A => n11057, ZN => n11348);
   U13216 : MUX2_X2 port map( A => n10149, B => n10148, S => n11348, Z => 
                           n12334);
   U13217 : XNOR2_X1 port map( A => n10151, B => n10150, ZN => n10153);
   U13218 : XNOR2_X1 port map( A => n19718, B => n2082, ZN => n10152);
   U13219 : XNOR2_X1 port map( A => n10153, B => n10152, ZN => n10156);
   U13220 : XNOR2_X1 port map( A => n1057, B => n10271, ZN => n10464);
   U13221 : XNOR2_X1 port map( A => n10548, B => n10464, ZN => n10155);
   U13222 : XNOR2_X1 port map( A => n260, B => n10430, ZN => n10159);
   U13223 : XNOR2_X1 port map( A => n10158, B => n10159, ZN => n10162);
   U13224 : XNOR2_X1 port map( A => n10431, B => n19052, ZN => n10160);
   U13225 : XNOR2_X1 port map( A => n10563, B => n10160, ZN => n10161);
   U13226 : INV_X1 port map( A => n11428, ZN => n11425);
   U13227 : XNOR2_X1 port map( A => n10514, B => n10163, ZN => n10164);
   U13228 : XNOR2_X1 port map( A => n10165, B => n10164, ZN => n10170);
   U13229 : INV_X1 port map( A => n10568, ZN => n10168);
   U13230 : XNOR2_X1 port map( A => n10166, B => n2035, ZN => n10167);
   U13231 : XNOR2_X1 port map( A => n10168, B => n10167, ZN => n10169);
   U13232 : AOI21_X1 port map( B1 => n11105, B2 => n11425, A => n11106, ZN => 
                           n10193);
   U13233 : XNOR2_X1 port map( A => n10473, B => n10171, ZN => n10172);
   U13234 : XNOR2_X1 port map( A => n10524, B => n10172, ZN => n10177);
   U13235 : XNOR2_X1 port map( A => n10173, B => n2369, ZN => n10175);
   U13236 : XNOR2_X1 port map( A => n10264, B => n10174, ZN => n10427);
   U13237 : XNOR2_X1 port map( A => n10427, B => n10175, ZN => n10176);
   U13238 : XNOR2_X1 port map( A => n10177, B => n10176, ZN => n11104);
   U13239 : INV_X1 port map( A => n11104, ZN => n11427);
   U13240 : XNOR2_X1 port map( A => n10289, B => n10220, ZN => n10415);
   U13241 : XNOR2_X1 port map( A => n10484, B => n2445, ZN => n10178);
   U13242 : XNOR2_X1 port map( A => n10415, B => n10178, ZN => n10184);
   U13243 : XNOR2_X1 port map( A => n19839, B => n10180, ZN => n10181);
   U13244 : XNOR2_X1 port map( A => n10182, B => n10181, ZN => n10183);
   U13245 : XNOR2_X1 port map( A => n10185, B => n10186, ZN => n10187);
   U13246 : XNOR2_X1 port map( A => n10187, B => n10611, ZN => n10190);
   U13247 : XNOR2_X1 port map( A => n10445, B => n18203, ZN => n10188);
   U13248 : XNOR2_X1 port map( A => n10535, B => n10188, ZN => n10189);
   U13249 : INV_X1 port map( A => n11106, ZN => n11424);
   U13250 : NAND3_X1 port map( A1 => n11425, A2 => n11430, A3 => n11424, ZN => 
                           n10191);
   U13251 : NAND2_X1 port map( A1 => n12334, A2 => n11990, ZN => n12333);
   U13252 : OAI21_X1 port map( B1 => n12338, B2 => n12334, A => n12333, ZN => 
                           n10317);
   U13254 : AOI21_X1 port map( B1 => n11337, B2 => n11263, A => n3669, ZN => 
                           n10198);
   U13255 : NOR2_X1 port map( A1 => n11267, A2 => n11265, ZN => n10797);
   U13256 : NOR2_X1 port map( A1 => n11339, A2 => n9830, ZN => n10196);
   U13257 : INV_X1 port map( A => n11263, ZN => n10195);
   U13258 : OAI21_X1 port map( B1 => n10797, B2 => n10196, A => n10195, ZN => 
                           n10197);
   U13259 : INV_X1 port map( A => n11992, ZN => n12337);
   U13260 : XNOR2_X1 port map( A => n19806, B => n10200, ZN => n10202);
   U13261 : XNOR2_X1 port map( A => n10201, B => n10202, ZN => n10209);
   U13262 : XNOR2_X1 port map( A => n10203, B => n10204, ZN => n10207);
   U13263 : XNOR2_X1 port map( A => n10205, B => n20064, ZN => n10206);
   U13264 : XNOR2_X1 port map( A => n10207, B => n10206, ZN => n10208);
   U13265 : XNOR2_X1 port map( A => n10209, B => n10208, ZN => n11460);
   U13266 : INV_X1 port map( A => n11460, ZN => n11048);
   U13270 : XNOR2_X1 port map( A => n10213, B => n10360, ZN => n10216);
   U13271 : XNOR2_X1 port map( A => n10214, B => n2055, ZN => n10215);
   U13272 : XNOR2_X1 port map( A => n10216, B => n10215, ZN => n10217);
   U13274 : XNOR2_X1 port map( A => n10219, B => n10220, ZN => n10221);
   U13275 : XNOR2_X1 port map( A => n10618, B => n10221, ZN => n10227);
   U13276 : XNOR2_X1 port map( A => n10222, B => n2446, ZN => n10225);
   U13277 : INV_X1 port map( A => n10223, ZN => n10224);
   U13278 : XNOR2_X1 port map( A => n10225, B => n10224, ZN => n10226);
   U13279 : XNOR2_X1 port map( A => n10226, B => n10227, ZN => n10259);
   U13280 : XNOR2_X1 port map( A => n10229, B => n10421, ZN => n10230);
   U13281 : XNOR2_X1 port map( A => n10603, B => n10230, ZN => n10235);
   U13282 : XNOR2_X1 port map( A => n10231, B => n106, ZN => n10232);
   U13283 : XNOR2_X1 port map( A => n10233, B => n10232, ZN => n10234);
   U13284 : XNOR2_X1 port map( A => n10235, B => n10234, ZN => n10808);
   U13285 : XNOR2_X1 port map( A => n10237, B => n10236, ZN => n10591);
   U13286 : INV_X1 port map( A => n10591, ZN => n10239);
   U13287 : XNOR2_X1 port map( A => n10239, B => n10238, ZN => n10244);
   U13288 : XNOR2_X1 port map( A => n10240, B => n10349, ZN => n10241);
   U13289 : XNOR2_X1 port map( A => n10242, B => n10241, ZN => n10243);
   U13290 : INV_X1 port map( A => n11120, ZN => n11881);
   U13291 : NAND2_X1 port map( A1 => n11881, A2 => n11460, ZN => n10245);
   U13292 : NAND3_X1 port map( A1 => n10246, A2 => n10788, A3 => n10245, ZN => 
                           n10260);
   U13293 : XNOR2_X1 port map( A => n10249, B => n15479, ZN => n10250);
   U13294 : XNOR2_X1 port map( A => n10251, B => n10250, ZN => n10256);
   U13295 : INV_X1 port map( A => n10252, ZN => n10253);
   U13296 : XNOR2_X1 port map( A => n10254, B => n10253, ZN => n10255);
   U13297 : XNOR2_X1 port map( A => n10256, B => n10255, ZN => n10258);
   U13298 : XNOR2_X1 port map( A => n10258, B => n10257, ZN => n11884);
   U13299 : NAND2_X1 port map( A1 => n10786, A2 => n10259, ZN => n11050);
   U13300 : INV_X1 port map( A => n11884, ZN => n11459);
   U13301 : INV_X1 port map( A => n12339, ZN => n11974);
   U13302 : INV_X1 port map( A => n12338, ZN => n10314);
   U13303 : XNOR2_X1 port map( A => n10261, B => n10262, ZN => n10263);
   U13304 : XNOR2_X1 port map( A => n10373, B => n10263, ZN => n10269);
   U13305 : XNOR2_X1 port map( A => n10604, B => n10264, ZN => n10267);
   U13306 : XNOR2_X1 port map( A => n10265, B => n2122, ZN => n10266);
   U13307 : XNOR2_X1 port map( A => n10267, B => n10266, ZN => n10268);
   U13308 : INV_X1 port map( A => n190, ZN => n11254);
   U13309 : XNOR2_X1 port map( A => n10271, B => n10270, ZN => n10272);
   U13310 : XNOR2_X1 port map( A => n10410, B => n10272, ZN => n10278);
   U13311 : XNOR2_X1 port map( A => n10273, B => n10582, ZN => n10276);
   U13312 : XNOR2_X1 port map( A => n10274, B => n2296, ZN => n10275);
   U13313 : XNOR2_X1 port map( A => n10276, B => n10275, ZN => n10277);
   U13314 : XNOR2_X1 port map( A => n10395, B => n10279, ZN => n10285);
   U13315 : XNOR2_X1 port map( A => n10280, B => n10431, ZN => n10283);
   U13316 : XNOR2_X1 port map( A => n10281, B => n2410, ZN => n10282);
   U13317 : XNOR2_X1 port map( A => n10283, B => n10282, ZN => n10284);
   U13318 : XNOR2_X1 port map( A => n10285, B => n10284, ZN => n11321);
   U13319 : XNOR2_X1 port map( A => n10286, B => n10320, ZN => n10288);
   U13320 : XNOR2_X1 port map( A => n10287, B => n10288, ZN => n10293);
   U13321 : XNOR2_X1 port map( A => n10289, B => n2395, ZN => n10291);
   U13322 : XNOR2_X1 port map( A => n10290, B => n10291, ZN => n10292);
   U13324 : INV_X1 port map( A => n11257, ZN => n11327);
   U13325 : INV_X1 port map( A => n2284, ZN => n18664);
   U13326 : XNOR2_X1 port map( A => n19785, B => n18664, ZN => n10295);
   U13327 : XNOR2_X1 port map( A => n10296, B => n10367, ZN => n10297);
   U13328 : XNOR2_X1 port map( A => n10298, B => n10445, ZN => n10300);
   U13329 : XNOR2_X1 port map( A => n10300, B => n19871, ZN => n10301);
   U13330 : XNOR2_X1 port map( A => n10302, B => n10301, ZN => n11256);
   U13331 : INV_X1 port map( A => n11256, ZN => n11322);
   U13332 : XNOR2_X1 port map( A => n10517, B => n10391, ZN => n10308);
   U13333 : XNOR2_X1 port map( A => n10303, B => n2337, ZN => n10306);
   U13334 : XNOR2_X1 port map( A => n10304, B => n10456, ZN => n10305);
   U13335 : XNOR2_X1 port map( A => n10306, B => n10305, ZN => n10307);
   U13336 : OAI21_X1 port map( B1 => n10310, B2 => n11322, A => n10309, ZN => 
                           n10311);
   U13337 : NOR2_X1 port map( A1 => n11992, A2 => n12335, ZN => n10313);
   U13338 : XNOR2_X1 port map( A => n13588, B => n13352, ZN => n13289);
   U13339 : INV_X1 port map( A => n13289, ZN => n10632);
   U13340 : XNOR2_X1 port map( A => n10318, B => n10319, ZN => n10324);
   U13341 : XNOR2_X1 port map( A => n10320, B => n2381, ZN => n10322);
   U13342 : XNOR2_X1 port map( A => n10321, B => n10322, ZN => n10323);
   U13344 : INV_X1 port map( A => n10328, ZN => n10326);
   U13345 : INV_X1 port map( A => n18304, ZN => n10325);
   U13346 : OAI21_X1 port map( B1 => n10327, B2 => n10326, A => n10325, ZN => 
                           n10331);
   U13347 : NAND3_X1 port map( A1 => n10329, A2 => n18304, A3 => n10328, ZN => 
                           n10330);
   U13348 : NAND2_X1 port map( A1 => n10331, A2 => n10330, ZN => n10333);
   U13349 : XNOR2_X1 port map( A => n10333, B => n20161, ZN => n10336);
   U13350 : INV_X1 port map( A => n10334, ZN => n10335);
   U13351 : XNOR2_X1 port map( A => n10336, B => n10335, ZN => n10338);
   U13352 : XNOR2_X1 port map( A => n10339, B => n19216, ZN => n10341);
   U13353 : XNOR2_X1 port map( A => n10341, B => n10340, ZN => n10345);
   U13354 : XNOR2_X1 port map( A => n10343, B => n10342, ZN => n10344);
   U13355 : XNOR2_X1 port map( A => n10345, B => n10344, ZN => n11087);
   U13356 : NAND2_X1 port map( A1 => n11455, A2 => n11454, ZN => n10346);
   U13357 : OAI21_X1 port map( B1 => n11455, B2 => n1812, A => n10346, ZN => 
                           n10366);
   U13358 : XNOR2_X1 port map( A => n10348, B => n10347, ZN => n10355);
   U13359 : XNOR2_X1 port map( A => n10349, B => n2392, ZN => n10353);
   U13360 : XNOR2_X1 port map( A => n10351, B => n10350, ZN => n10352);
   U13361 : XNOR2_X1 port map( A => n10353, B => n10352, ZN => n10354);
   U13362 : NOR2_X1 port map( A1 => n11452, A2 => n11455, ZN => n10365);
   U13363 : XNOR2_X1 port map( A => n10357, B => n10356, ZN => n10364);
   U13364 : XNOR2_X1 port map( A => n928, B => n18170, ZN => n10362);
   U13365 : XNOR2_X1 port map( A => n10359, B => n10360, ZN => n10361);
   U13366 : XNOR2_X1 port map( A => n10362, B => n10361, ZN => n10363);
   U13367 : XNOR2_X1 port map( A => n10367, B => n16366, ZN => n10369);
   U13368 : BUF_X2 port map( A => n11088, Z => n11455);
   U13369 : NAND2_X1 port map( A1 => n11455, A2 => n11114, ZN => n10372);
   U13370 : XNOR2_X1 port map( A => n10374, B => n10373, ZN => n10378);
   U13371 : XNOR2_X1 port map( A => n10528, B => n19027, ZN => n10375);
   U13372 : XNOR2_X1 port map( A => n10376, B => n10375, ZN => n10377);
   U13373 : INV_X1 port map( A => n10379, ZN => n10380);
   U13374 : XNOR2_X1 port map( A => n10380, B => n10381, ZN => n10386);
   U13375 : XNOR2_X1 port map( A => n10482, B => n10382, ZN => n10384);
   U13376 : XNOR2_X1 port map( A => n10384, B => n10383, ZN => n10385);
   U13377 : XNOR2_X1 port map( A => n10387, B => n10388, ZN => n10390);
   U13378 : XNOR2_X1 port map( A => n10570, B => n18055, ZN => n10389);
   U13379 : XNOR2_X1 port map( A => n10390, B => n10389, ZN => n10394);
   U13380 : XNOR2_X1 port map( A => n10392, B => n10391, ZN => n10393);
   U13381 : XNOR2_X1 port map( A => n10394, B => n10393, ZN => n11132);
   U13382 : XNOR2_X1 port map( A => n10395, B => n10396, ZN => n10400);
   U13383 : XNOR2_X1 port map( A => n10561, B => n18078, ZN => n10398);
   U13384 : XNOR2_X1 port map( A => n10397, B => n10398, ZN => n10399);
   U13385 : XNOR2_X1 port map( A => n10400, B => n10399, ZN => n10724);
   U13386 : AOI22_X1 port map( A1 => n11133, A2 => n11131, B1 => n19837, B2 => 
                           n10724, ZN => n11054);
   U13387 : INV_X1 port map( A => n11131, ZN => n11420);
   U13388 : NOR2_X1 port map( A1 => n11133, A2 => n11420, ZN => n10414);
   U13389 : XNOR2_X1 port map( A => n10401, B => n10402, ZN => n10534);
   U13390 : XNOR2_X1 port map( A => n10534, B => n10403, ZN => n10408);
   U13391 : XNOR2_X1 port map( A => n10404, B => n16035, ZN => n10405);
   U13392 : XNOR2_X1 port map( A => n10406, B => n10405, ZN => n10407);
   U13394 : XNOR2_X1 port map( A => n10409, B => n10410, ZN => n10411);
   U13395 : OAI21_X1 port map( B1 => n11054, B2 => n10414, A => n10413, ZN => 
                           n11997);
   U13396 : INV_X1 port map( A => n11997, ZN => n12515);
   U13397 : XNOR2_X1 port map( A => n10416, B => n10415, ZN => n10420);
   U13398 : XNOR2_X1 port map( A => n10417, B => n10418, ZN => n10419);
   U13399 : XNOR2_X1 port map( A => n10420, B => n10419, ZN => n10450);
   U13400 : XNOR2_X1 port map( A => n10422, B => n10421, ZN => n10424);
   U13401 : XNOR2_X1 port map( A => n10424, B => n20456, ZN => n10429);
   U13402 : XNOR2_X1 port map( A => n10425, B => n16651, ZN => n10426);
   U13403 : XNOR2_X1 port map( A => n10427, B => n10426, ZN => n10428);
   U13404 : INV_X1 port map( A => n10430, ZN => n10432);
   U13405 : XNOR2_X1 port map( A => n10432, B => n10431, ZN => n10434);
   U13406 : XNOR2_X1 port map( A => n10434, B => n10433, ZN => n10440);
   U13407 : INV_X1 port map( A => n18830, ZN => n10435);
   U13408 : XNOR2_X1 port map( A => n10436, B => n10435, ZN => n10437);
   U13409 : XOR2_X1 port map( A => n10438, B => n10437, Z => n10439);
   U13411 : XNOR2_X1 port map( A => n10441, B => n10442, ZN => n10443);
   U13412 : XNOR2_X1 port map( A => n10444, B => n10443, ZN => n10449);
   U13413 : XNOR2_X1 port map( A => n10445, B => n18433, ZN => n10446);
   U13414 : XNOR2_X1 port map( A => n10447, B => n10446, ZN => n10448);
   U13415 : XNOR2_X1 port map( A => n10449, B => n10448, ZN => n11446);
   U13416 : NOR2_X1 port map( A1 => n11446, A2 => n11202, ZN => n10452);
   U13417 : INV_X1 port map( A => n19920, ZN => n10451);
   U13418 : INV_X1 port map( A => n10453, ZN => n10455);
   U13419 : XNOR2_X1 port map( A => n10455, B => n10454, ZN => n10460);
   U13420 : XNOR2_X1 port map( A => n10456, B => n2275, ZN => n10457);
   U13421 : XNOR2_X1 port map( A => n10458, B => n10457, ZN => n10459);
   U13422 : NAND2_X1 port map( A1 => n11202, A2 => n10845, ZN => n10468);
   U13423 : XNOR2_X1 port map( A => n10461, B => n18984, ZN => n10463);
   U13424 : XNOR2_X1 port map( A => n10463, B => n10462, ZN => n10467);
   U13425 : XNOR2_X1 port map( A => n10464, B => n10465, ZN => n10466);
   U13426 : XNOR2_X1 port map( A => n10467, B => n10466, ZN => n10726);
   U13427 : INV_X1 port map( A => n11995, ZN => n12325);
   U13428 : XNOR2_X1 port map( A => n10472, B => n18691, ZN => n10474);
   U13429 : XNOR2_X1 port map( A => n10474, B => n10473, ZN => n10476);
   U13430 : XNOR2_X1 port map( A => n10476, B => n10475, ZN => n10479);
   U13431 : INV_X1 port map( A => n10477, ZN => n10478);
   U13432 : XNOR2_X1 port map( A => n10480, B => n10481, ZN => n10488);
   U13433 : XNOR2_X1 port map( A => n10482, B => n10483, ZN => n10486);
   U13434 : XNOR2_X1 port map( A => n10484, B => n18070, ZN => n10485);
   U13435 : XNOR2_X1 port map( A => n10486, B => n10485, ZN => n10487);
   U13436 : XNOR2_X1 port map( A => n10488, B => n10487, ZN => n10513);
   U13437 : INV_X1 port map( A => n10489, ZN => n10496);
   U13438 : XNOR2_X1 port map( A => n10490, B => n2310, ZN => n10492);
   U13439 : XNOR2_X1 port map( A => n10492, B => n10491, ZN => n10493);
   U13440 : XNOR2_X1 port map( A => n10494, B => n10493, ZN => n10495);
   U13441 : XNOR2_X1 port map( A => n10497, B => n19243, ZN => n10500);
   U13442 : INV_X1 port map( A => n10498, ZN => n10499);
   U13443 : XNOR2_X1 port map( A => n10500, B => n10499, ZN => n10502);
   U13444 : XNOR2_X1 port map( A => n10502, B => n10501, ZN => n10504);
   U13445 : XNOR2_X1 port map( A => n10504, B => n10503, ZN => n11115);
   U13446 : NOR2_X1 port map( A1 => n11116, A2 => n11115, ZN => n10505);
   U13447 : XNOR2_X1 port map( A => n10506, B => n2454, ZN => n10507);
   U13448 : XNOR2_X1 port map( A => n10509, B => n10508, ZN => n10512);
   U13449 : INV_X1 port map( A => n10510, ZN => n10511);
   U13450 : AND2_X1 port map( A1 => n11037, A2 => n11440, ZN => n11117);
   U13451 : XNOR2_X1 port map( A => n10566, B => n10514, ZN => n10516);
   U13452 : XNOR2_X1 port map( A => n10515, B => n10516, ZN => n10521);
   U13453 : INV_X1 port map( A => n10517, ZN => n10519);
   U13454 : XNOR2_X1 port map( A => n10572, B => n20682, ZN => n10518);
   U13455 : XNOR2_X1 port map( A => n10519, B => n10518, ZN => n10520);
   U13457 : OAI21_X1 port map( B1 => n11117, B2 => n11035, A => n11116, ZN => 
                           n10522);
   U13459 : XNOR2_X1 port map( A => n10524, B => n10525, ZN => n10532);
   U13460 : XNOR2_X1 port map( A => n10527, B => n10526, ZN => n10530);
   U13461 : XNOR2_X1 port map( A => n10528, B => n18809, ZN => n10529);
   U13462 : XNOR2_X1 port map( A => n10530, B => n10529, ZN => n10531);
   U13463 : XNOR2_X2 port map( A => n10532, B => n10531, ZN => n11193);
   U13464 : XNOR2_X1 port map( A => n10534, B => n10533, ZN => n10539);
   U13465 : XNOR2_X1 port map( A => n10613, B => n18887, ZN => n10537);
   U13466 : INV_X1 port map( A => n10535, ZN => n10536);
   U13467 : XNOR2_X1 port map( A => n10536, B => n10537, ZN => n10538);
   U13468 : XNOR2_X1 port map( A => n10540, B => n10541, ZN => n10547);
   U13469 : XNOR2_X1 port map( A => n865, B => n311, ZN => n10545);
   U13470 : INV_X1 port map( A => n10543, ZN => n10544);
   U13471 : XNOR2_X1 port map( A => n10544, B => n10545, ZN => n10546);
   U13472 : NAND2_X1 port map( A1 => n11186, A2 => n19983, ZN => n10903);
   U13473 : XNOR2_X1 port map( A => n10548, B => n10549, ZN => n10556);
   U13474 : XNOR2_X1 port map( A => n10550, B => n2032, ZN => n10554);
   U13475 : XNOR2_X1 port map( A => n10552, B => n10551, ZN => n10553);
   U13476 : XNOR2_X1 port map( A => n10554, B => n10553, ZN => n10555);
   U13477 : XNOR2_X1 port map( A => n10557, B => n10558, ZN => n10560);
   U13478 : XNOR2_X1 port map( A => n10560, B => n10559, ZN => n10565);
   U13479 : XNOR2_X1 port map( A => n10561, B => n19336, ZN => n10562);
   U13480 : XNOR2_X1 port map( A => n10562, B => n10563, ZN => n10564);
   U13481 : XNOR2_X1 port map( A => n10564, B => n10565, ZN => n10575);
   U13482 : XNOR2_X1 port map( A => n10566, B => n10567, ZN => n10569);
   U13483 : XNOR2_X1 port map( A => n10571, B => n10570, ZN => n10574);
   U13484 : XNOR2_X1 port map( A => n10572, B => n2376, ZN => n10573);
   U13485 : OAI21_X1 port map( B1 => n11500, B2 => n11499, A => n11192, ZN => 
                           n10577);
   U13486 : INV_X1 port map( A => n10575, ZN => n11188);
   U13487 : NAND2_X1 port map( A1 => n11188, A2 => n11192, ZN => n11502);
   U13488 : INV_X1 port map( A => n11502, ZN => n10576);
   U13489 : NAND2_X1 port map( A1 => n11995, A2 => n11820, ZN => n10627);
   U13490 : XNOR2_X1 port map( A => n10578, B => n10579, ZN => n10581);
   U13491 : XNOR2_X1 port map( A => n10581, B => n10580, ZN => n10586);
   U13492 : XNOR2_X1 port map( A => n10582, B => n19180, ZN => n10583);
   U13493 : XNOR2_X1 port map( A => n10584, B => n10583, ZN => n10585);
   U13494 : INV_X1 port map( A => n11491, ZN => n11495);
   U13495 : XNOR2_X1 port map( A => n10588, B => n10587, ZN => n10593);
   U13496 : XNOR2_X1 port map( A => n10589, B => n19140, ZN => n10590);
   U13497 : XNOR2_X1 port map( A => n10591, B => n10590, ZN => n10592);
   U13498 : XNOR2_X1 port map( A => n10594, B => n10595, ZN => n10597);
   U13499 : XNOR2_X1 port map( A => n10596, B => n10597, ZN => n10602);
   U13500 : INV_X1 port map( A => Key(124), ZN => n18517);
   U13501 : XNOR2_X1 port map( A => n10598, B => n18517, ZN => n10599);
   U13502 : XNOR2_X1 port map( A => n10600, B => n10599, ZN => n10601);
   U13504 : INV_X1 port map( A => n10603, ZN => n10608);
   U13505 : XNOR2_X1 port map( A => n10606, B => n10605, ZN => n10607);
   U13506 : XNOR2_X1 port map( A => n10608, B => n10607, ZN => n10610);
   U13507 : XNOR2_X1 port map( A => n961, B => n10611, ZN => n10617);
   U13508 : XNOR2_X1 port map( A => n10613, B => n10612, ZN => n10616);
   U13509 : XNOR2_X1 port map( A => n20210, B => n2096, ZN => n10615);
   U13510 : XNOR2_X1 port map( A => n10619, B => n10618, ZN => n10622);
   U13511 : NOR2_X1 port map( A1 => n11494, A2 => n11493, ZN => n10623);
   U13513 : INV_X1 port map( A => n10625, ZN => n12326);
   U13514 : NAND2_X1 port map( A1 => n12513, A2 => n12326, ZN => n10626);
   U13515 : OAI22_X1 port map( A1 => n20073, A2 => n10627, B1 => n10626, B2 => 
                           n13275, ZN => n10629);
   U13516 : AOI21_X1 port map( B1 => n13275, B2 => n10630, A => n10629, ZN => 
                           n12962);
   U13517 : INV_X1 port map( A => n12962, ZN => n13590);
   U13518 : INV_X1 port map( A => n2100, ZN => n15021);
   U13519 : XNOR2_X1 port map( A => n13590, B => n15021, ZN => n10631);
   U13520 : XNOR2_X1 port map( A => n10632, B => n10631, ZN => n10633);
   U13521 : XNOR2_X1 port map( A => n10633, B => n10634, ZN => n14775);
   U13522 : INV_X1 port map( A => n14775, ZN => n14057);
   U13523 : AOI21_X1 port map( B1 => n11528, B2 => n11521, A => n10635, ZN => 
                           n10636);
   U13524 : INV_X1 port map( A => n11528, ZN => n10921);
   U13525 : MUX2_X1 port map( A => n10636, B => n10924, S => n10755, Z => 
                           n10637);
   U13526 : NOR2_X1 port map( A1 => n10638, A2 => n10640, ZN => n10932);
   U13527 : NOR2_X1 port map( A1 => n11168, A2 => n11539, ZN => n10639);
   U13528 : OAI211_X1 port map( C1 => n11534, C2 => n11170, A => n11538, B => 
                           n11168, ZN => n10641);
   U13529 : OAI21_X1 port map( B1 => n10737, B2 => n11169, A => n10641, ZN => 
                           n12422);
   U13530 : NAND2_X1 port map( A1 => n12415, A2 => n12422, ZN => n11312);
   U13531 : AOI22_X1 port map( A1 => n1721, A2 => n20366, B1 => n10642, B2 => 
                           n10960, ZN => n10644);
   U13532 : NAND2_X1 port map( A1 => n11142, A2 => n10642, ZN => n10957);
   U13533 : MUX2_X1 port map( A => n10960, B => n10957, S => n11145, Z => 
                           n10643);
   U13534 : OAI21_X2 port map( B1 => n10644, B2 => n10701, A => n10643, ZN => 
                           n12416);
   U13537 : NAND2_X1 port map( A1 => n12416, A2 => n20352, ZN => n11311);
   U13538 : NAND2_X1 port map( A1 => n11161, A2 => n10649, ZN => n10654);
   U13539 : NAND2_X1 port map( A1 => n10650, A2 => n11159, ZN => n10651);
   U13540 : MUX2_X1 port map( A => n10652, B => n10651, S => n10945, Z => 
                           n10653);
   U13542 : INV_X1 port map( A => n11602, ZN => n12419);
   U13543 : AOI21_X1 port map( B1 => n11312, B2 => n11311, A => n12419, ZN => 
                           n10659);
   U13546 : AOI21_X1 port map( B1 => n12083, B2 => n12415, A => n20352, ZN => 
                           n10658);
   U13548 : NAND2_X1 port map( A1 => n11659, A2 => n11830, ZN => n11954);
   U13549 : NAND2_X1 port map( A1 => n11957, A2 => n11954, ZN => n10660);
   U13550 : XNOR2_X1 port map( A => n13088, B => n13192, ZN => n11975);
   U13551 : AOI22_X1 port map( A1 => n11254, A2 => n11253, B1 => n11256, B2 => 
                           n11255, ZN => n10663);
   U13552 : NAND2_X1 port map( A1 => n11256, A2 => n11257, ZN => n10664);
   U13553 : MUX2_X1 port map( A => n11255, B => n10664, S => n191, Z => n10665)
                           ;
   U13554 : INV_X1 port map( A => n11395, ZN => n11296);
   U13555 : NAND2_X1 port map( A1 => n2724, A2 => n10667, ZN => n10668);
   U13556 : INV_X1 port map( A => n10986, ZN => n11398);
   U13557 : INV_X1 port map( A => n11397, ZN => n11295);
   U13558 : MUX2_X1 port map( A => n10668, B => n11398, S => n11295, Z => 
                           n10669);
   U13559 : NAND2_X1 port map( A1 => n12099, A2 => n12435, ZN => n10687);
   U13560 : MUX2_X1 port map( A => n11267, B => n11265, S => n11339, Z => 
                           n10674);
   U13561 : NAND2_X1 port map( A1 => n11263, A2 => n11265, ZN => n10671);
   U13562 : NAND2_X1 port map( A1 => n10673, A2 => n9830, ZN => n10670);
   U13563 : MUX2_X1 port map( A => n10671, B => n10670, S => n11343, Z => 
                           n10672);
   U13564 : INV_X1 port map( A => n10675, ZN => n10818);
   U13565 : NOR2_X1 port map( A1 => n10852, A2 => n11231, ZN => n10678);
   U13566 : MUX2_X1 port map( A => n10679, B => n10678, S => n11366, Z => 
                           n10682);
   U13567 : NAND2_X1 port map( A1 => n10818, A2 => n11234, ZN => n10680);
   U13568 : NOR2_X1 port map( A1 => n12437, A2 => n12440, ZN => n11065);
   U13569 : AOI21_X2 port map( B1 => n10687, B2 => n10686, A => n11065, ZN => 
                           n13618);
   U13570 : MUX2_X1 port map( A => n11408, B => n10688, S => n19736, Z => 
                           n10692);
   U13571 : NAND2_X1 port map( A1 => n11000, A2 => n11278, ZN => n11410);
   U13572 : INV_X1 port map( A => n11410, ZN => n10690);
   U13573 : NOR2_X1 port map( A1 => n11278, A2 => n11413, ZN => n10689);
   U13574 : AOI22_X1 port map( A1 => n10690, A2 => n11411, B1 => n10689, B2 => 
                           n11408, ZN => n10691);
   U13575 : INV_X1 port map( A => n12631, ZN => n12629);
   U13576 : MUX2_X1 port map( A => n10947, B => n10693, S => n19779, Z => 
                           n10695);
   U13577 : NOR2_X1 port map( A1 => n9559, A2 => n10694, ZN => n10999);
   U13578 : NOR2_X1 port map( A1 => n10980, A2 => n11294, ZN => n10697);
   U13579 : NOR2_X1 port map( A1 => n20235, A2 => n11290, ZN => n10696);
   U13581 : NAND2_X1 port map( A1 => n11292, A2 => n11403, ZN => n10698);
   U13582 : AOI21_X1 port map( B1 => n10698, B2 => n11293, A => n11291, ZN => 
                           n10699);
   U13583 : NOR2_X2 port map( A1 => n10700, A2 => n10699, ZN => n12634);
   U13584 : OAI22_X1 port map( A1 => n11145, A2 => n1749, B1 => n20366, B2 => 
                           n10701, ZN => n10703);
   U13586 : NAND3_X1 port map( A1 => n11148, A2 => n11147, A3 => n11009, ZN => 
                           n10704);
   U13587 : NAND2_X1 port map( A1 => n11009, A2 => n10953, ZN => n11152);
   U13589 : INV_X1 port map( A => n10709, ZN => n11869);
   U13590 : OAI21_X1 port map( B1 => n20601, B2 => n11866, A => n11869, ZN => 
                           n10710);
   U13591 : INV_X1 port map( A => n10711, ZN => n10712);
   U13592 : INV_X1 port map( A => n11871, ZN => n11388);
   U13593 : NAND2_X1 port map( A1 => n10712, A2 => n11388, ZN => n10713);
   U13594 : INV_X1 port map( A => n12634, ZN => n10716);
   U13595 : XNOR2_X1 port map( A => n13415, B => n11975, ZN => n10795);
   U13596 : NAND2_X1 port map( A1 => n10717, A2 => n11076, ZN => n10718);
   U13597 : INV_X1 port map( A => n11191, ZN => n11501);
   U13598 : NOR2_X1 port map( A1 => n11500, A2 => n11501, ZN => n10719);
   U13600 : NOR2_X1 port map( A1 => n11193, A2 => n19983, ZN => n10721);
   U13601 : NOR2_X1 port map( A1 => n11192, A2 => n11188, ZN => n10720);
   U13602 : AOI22_X1 port map( A1 => n10721, A2 => n11186, B1 => n10720, B2 => 
                           n11193, ZN => n10722);
   U13603 : INV_X1 port map( A => n12648, ZN => n12645);
   U13604 : INV_X1 port map( A => n11132, ZN => n11417);
   U13605 : INV_X1 port map( A => n11446, ZN => n10847);
   U13606 : MUX2_X1 port map( A => n10847, B => n11093, S => n19920, Z => 
                           n10728);
   U13607 : MUX2_X2 port map( A => n10728, B => n10727, S => n11094, Z => 
                           n12684);
   U13608 : INV_X1 port map( A => n10730, ZN => n11069);
   U13609 : NAND2_X1 port map( A1 => n11069, A2 => n11489, ZN => n10732);
   U13610 : NAND2_X1 port map( A1 => n19505, A2 => n19719, ZN => n10731);
   U13611 : INV_X1 port map( A => n11456, ZN => n11091);
   U13612 : OAI21_X1 port map( B1 => n10734, B2 => n11091, A => n10733, ZN => 
                           n10736);
   U13613 : AOI21_X1 port map( B1 => n10734, B2 => n11114, A => n11455, ZN => 
                           n10735);
   U13614 : NOR2_X1 port map( A1 => n10736, A2 => n10735, ZN => n12430);
   U13615 : AND2_X2 port map( A1 => n10739, A2 => n10738, ZN => n12759);
   U13616 : INV_X1 port map( A => n12759, ZN => n12410);
   U13617 : INV_X1 port map( A => n11514, ZN => n10906);
   U13618 : INV_X1 port map( A => n11515, ZN => n10935);
   U13619 : INV_X1 port map( A => n10740, ZN => n10741);
   U13620 : OAI21_X1 port map( B1 => n10906, B2 => n11513, A => n10741, ZN => 
                           n10743);
   U13622 : INV_X1 port map( A => n10896, ZN => n11483);
   U13623 : AOI21_X1 port map( B1 => n11487, B2 => n11483, A => n20233, ZN => 
                           n10750);
   U13624 : NAND2_X1 port map( A1 => n10745, A2 => n20233, ZN => n10747);
   U13625 : AOI21_X1 port map( B1 => n10748, B2 => n10747, A => n3500, ZN => 
                           n10749);
   U13626 : NOR2_X1 port map( A1 => n898, A2 => n11568, ZN => n10754);
   U13627 : NAND2_X1 port map( A1 => n10883, A2 => n11566, ZN => n10753);
   U13628 : INV_X1 port map( A => n10883, ZN => n11567);
   U13629 : NAND2_X1 port map( A1 => n11567, A2 => n11466, ZN => n10751);
   U13631 : AOI22_X1 port map( A1 => n12410, A2 => n12754, B1 => n254, B2 => 
                           n12407, ZN => n11315);
   U13633 : NAND2_X1 port map( A1 => n10755, A2 => n11527, ZN => n10757);
   U13634 : INV_X1 port map( A => n12754, ZN => n10766);
   U13635 : NAND3_X1 port map( A1 => n10889, A2 => n10760, A3 => n11546, ZN => 
                           n10763);
   U13636 : INV_X1 port map( A => n12407, ZN => n11313);
   U13637 : OAI21_X1 port map( B1 => n12389, B2 => n11313, A => n254, ZN => 
                           n10765);
   U13638 : NAND2_X1 port map( A1 => n10766, A2 => n10765, ZN => n10767);
   U13639 : INV_X1 port map( A => n11430, ZN => n10768);
   U13640 : NOR2_X1 port map( A1 => n19830, A2 => n10768, ZN => n10770);
   U13641 : MUX2_X1 port map( A => n10770, B => n10769, S => n11041, Z => 
                           n10773);
   U13642 : INV_X1 port map( A => n11105, ZN => n11429);
   U13644 : NAND2_X1 port map( A1 => n11105, A2 => n19830, ZN => n11109);
   U13646 : NOR2_X2 port map( A1 => n10773, A2 => n10772, ZN => n12639);
   U13647 : OAI21_X1 port map( B1 => n10802, B2 => n10774, A => n11257, ZN => 
                           n10778);
   U13648 : INV_X1 port map( A => n11255, ZN => n10775);
   U13649 : MUX2_X1 port map( A => n10776, B => n10775, S => n11253, Z => 
                           n10777);
   U13650 : NAND2_X1 port map( A1 => n10778, A2 => n10777, ZN => n12453);
   U13651 : NAND2_X1 port map( A1 => n11238, A2 => n10779, ZN => n11236);
   U13652 : OAI211_X1 port map( C1 => n11349, C2 => n11057, A => n11239, B => 
                           n10798, ZN => n10780);
   U13653 : NAND2_X1 port map( A1 => n11347, A2 => n11057, ZN => n11237);
   U13654 : OAI211_X1 port map( C1 => n11057, C2 => n11236, A => n10780, B => 
                           n11237, ZN => n12449);
   U13655 : NAND2_X1 port map( A1 => n12453, A2 => n12449, ZN => n11946);
   U13656 : INV_X1 port map( A => n11115, ZN => n11439);
   U13657 : NAND2_X1 port map( A1 => n11439, A2 => n11035, ZN => n10782);
   U13658 : NAND2_X1 port map( A1 => n11034, A2 => n11440, ZN => n10781);
   U13659 : NAND2_X1 port map( A1 => n10782, A2 => n10781, ZN => n10833);
   U13660 : OAI21_X1 port map( B1 => n11438, B2 => n11115, A => n11035, ZN => 
                           n10784);
   U13661 : NAND2_X1 port map( A1 => n12637, A2 => n12642, ZN => n10792);
   U13662 : MUX2_X1 port map( A => n11886, B => n11880, S => n11120, Z => 
                           n10789);
   U13663 : NAND2_X1 port map( A1 => n12636, A2 => n12449, ZN => n12089);
   U13664 : INV_X1 port map( A => n12089, ZN => n10790);
   U13665 : INV_X1 port map( A => n12453, ZN => n12450);
   U13666 : INV_X1 port map( A => n12642, ZN => n12452);
   U13667 : OAI21_X1 port map( B1 => n10790, B2 => n12450, A => n12452, ZN => 
                           n10791);
   U13669 : XNOR2_X1 port map( A => n13617, B => n13336, ZN => n13305);
   U13670 : XNOR2_X1 port map( A => n13305, B => n10793, ZN => n10794);
   U13671 : NOR2_X1 port map( A1 => n11337, A2 => n11263, ZN => n10796);
   U13672 : AND2_X1 port map( A1 => n11355, A2 => n10798, ZN => n10799);
   U13673 : AND2_X1 port map( A1 => n11239, A2 => n11347, ZN => n10800);
   U13674 : INV_X1 port map( A => n10800, ZN => n10801);
   U13675 : NAND2_X1 port map( A1 => n12212, A2 => n12208, ZN => n11639);
   U13676 : NAND2_X1 port map( A1 => n10805, A2 => n10804, ZN => n10807);
   U13677 : AND2_X1 port map( A1 => n11321, A2 => n11253, ZN => n11324);
   U13678 : AOI21_X1 port map( B1 => n11124, B2 => n10809, A => n11459, ZN => 
                           n10812);
   U13679 : AOI21_X1 port map( B1 => n10810, B2 => n11048, A => n11883, ZN => 
                           n10811);
   U13680 : NOR2_X1 port map( A1 => n20099, A2 => n11125, ZN => n10816);
   U13681 : NOR2_X1 port map( A1 => n11127, A2 => n10813, ZN => n10815);
   U13682 : OAI22_X1 port map( A1 => n10818, A2 => n1601, B1 => n11231, B2 => 
                           n11234, ZN => n10820);
   U13683 : INV_X1 port map( A => n11235, ZN => n10819);
   U13684 : NOR2_X1 port map( A1 => n9883, A2 => n10854, ZN => n11638);
   U13685 : INV_X1 port map( A => n11638, ZN => n11808);
   U13686 : NOR2_X1 port map( A1 => n11811, A2 => n10821, ZN => n10822);
   U13687 : NAND2_X1 port map( A1 => n913, A2 => n3051, ZN => n11200);
   U13688 : NAND2_X1 port map( A1 => n11199, A2 => n11200, ZN => n10825);
   U13689 : OAI21_X1 port map( B1 => n19719, B2 => n19913, A => n913, ZN => 
                           n10824);
   U13690 : INV_X1 port map( A => n12061, ZN => n11637);
   U13691 : NAND3_X1 port map( A1 => n11042, A2 => n11106, A3 => n11105, ZN => 
                           n10828);
   U13693 : NOR2_X1 port map( A1 => n1378, A2 => n11430, ZN => n10826);
   U13695 : INV_X1 port map( A => n12202, ZN => n12591);
   U13696 : NOR2_X1 port map( A1 => n11637, A2 => n12591, ZN => n10844);
   U13699 : INV_X1 port map( A => n12594, ZN => n12590);
   U13700 : OAI211_X1 port map( C1 => n11037, C2 => n11440, A => n11115, B => 
                           n11438, ZN => n10835);
   U13701 : NAND2_X1 port map( A1 => n11451, A2 => n11455, ZN => n10843);
   U13702 : INV_X1 port map( A => n11088, ZN => n10839);
   U13703 : NAND2_X1 port map( A1 => n10839, A2 => n11452, ZN => n10838);
   U13704 : OAI21_X1 port map( B1 => n11451, B2 => n11452, A => n10838, ZN => 
                           n10841);
   U13705 : NAND2_X1 port map( A1 => n10839, A2 => n11113, ZN => n11112);
   U13706 : NAND2_X1 port map( A1 => n11112, A2 => n11114, ZN => n10840);
   U13707 : OAI21_X1 port map( B1 => n10841, B2 => n11114, A => n10840, ZN => 
                           n10842);
   U13708 : AOI21_X1 port map( B1 => n10845, B2 => n11445, A => n11443, ZN => 
                           n10846);
   U13709 : INV_X1 port map( A => n10845, ZN => n11444);
   U13710 : XNOR2_X1 port map( A => n13577, B => n10849, ZN => n13357);
   U13711 : INV_X1 port map( A => n13357, ZN => n10881);
   U13712 : INV_X1 port map( A => n11670, ZN => n12185);
   U13713 : NOR2_X1 port map( A1 => n11841, A2 => n20427, ZN => n11844);
   U13714 : NAND2_X1 port map( A1 => n11844, A2 => n11670, ZN => n10850);
   U13715 : INV_X1 port map( A => n11369, ZN => n10853);
   U13716 : NOR2_X1 port map( A1 => n10854, A2 => n11234, ZN => n10855);
   U13718 : NAND2_X1 port map( A1 => n10986, A2 => n11397, ZN => n10859);
   U13719 : AOI21_X1 port map( B1 => n19756, B2 => n12057, A => n874, ZN => 
                           n10879);
   U13720 : INV_X1 port map( A => n19750, ZN => n11867);
   U13721 : NAND2_X1 port map( A1 => n20601, A2 => n11866, ZN => n11305);
   U13722 : INV_X1 port map( A => n11305, ZN => n10863);
   U13724 : NAND2_X1 port map( A1 => n10868, A2 => n10867, ZN => n12615);
   U13725 : NAND2_X1 port map( A1 => n11380, A2 => n12103, ZN => n10866);
   U13726 : NAND2_X1 port map( A1 => n10864, A2 => n12101, ZN => n10865);
   U13727 : MUX2_X1 port map( A => n10866, B => n10865, S => n11381, Z => 
                           n11632);
   U13728 : NAND4_X1 port map( A1 => n11632, A2 => n10868, A3 => n11633, A4 => 
                           n10867, ZN => n10869);
   U13729 : OAI22_X1 port map( A1 => n19756, A2 => n12053, B1 => n10869, B2 => 
                           n12240, ZN => n10878);
   U13730 : OAI22_X1 port map( A1 => n10978, A2 => n19506, B1 => n11402, B2 => 
                           n3588, ZN => n10871);
   U13731 : OAI22_X1 port map( A1 => n11293, A2 => n20235, B1 => n11403, B2 => 
                           n11291, ZN => n10870);
   U13732 : INV_X1 port map( A => n11632, ZN => n10875);
   U13733 : INV_X1 port map( A => n10873, ZN => n10874);
   U13734 : NOR2_X1 port map( A1 => n10875, A2 => n10874, ZN => n10876);
   U13735 : XNOR2_X1 port map( A => n13827, B => n19854, ZN => n10880);
   U13736 : XNOR2_X1 port map( A => n10881, B => n10880, ZN => n10977);
   U13737 : INV_X1 port map( A => n10882, ZN => n11469);
   U13738 : MUX2_X1 port map( A => n11568, B => n10884, S => n10883, Z => 
                           n10888);
   U13739 : NAND2_X1 port map( A1 => n11565, A2 => n11569, ZN => n10887);
   U13740 : INV_X1 port map( A => n927, ZN => n11467);
   U13741 : INV_X1 port map( A => n11466, ZN => n11564);
   U13742 : NOR2_X1 port map( A1 => n11467, A2 => n10885, ZN => n10886);
   U13744 : OAI22_X1 port map( A1 => n647, A2 => n10926, B1 => n10889, B2 => 
                           n11547, ZN => n10890);
   U13745 : NAND2_X1 port map( A1 => n11544, A2 => n647, ZN => n10892);
   U13746 : INV_X1 port map( A => n11217, ZN => n10895);
   U13747 : MUX2_X1 port map( A => n19897, B => n10896, S => n10060, Z => 
                           n10900);
   U13748 : INV_X1 port map( A => n10898, ZN => n10899);
   U13749 : AOI22_X1 port map( A1 => n11193, A2 => n19983, B1 => n11188, B2 => 
                           n11500, ZN => n10901);
   U13750 : NOR2_X1 port map( A1 => n10901, A2 => n11186, ZN => n10905);
   U13751 : AOI21_X1 port map( B1 => n10903, B2 => n19998, A => n11500, ZN => 
                           n10904);
   U13752 : NOR2_X1 port map( A1 => n10905, A2 => n10904, ZN => n12601);
   U13753 : NAND2_X1 port map( A1 => n12609, A2 => n12601, ZN => n10911);
   U13755 : NAND3_X1 port map( A1 => n20106, A2 => n20639, A3 => n11572, ZN => 
                           n10910);
   U13756 : NAND3_X1 port map( A1 => n11510, A2 => n19864, A3 => n10936, ZN => 
                           n10909);
   U13757 : NAND3_X1 port map( A1 => n10935, A2 => n11510, A3 => n10906, ZN => 
                           n10907);
   U13759 : INV_X1 port map( A => n10913, ZN => n11557);
   U13760 : MUX2_X1 port map( A => n11556, B => n11557, S => n10914, Z => 
                           n10918);
   U13761 : INV_X1 port map( A => n11553, ZN => n11163);
   U13762 : NAND2_X1 port map( A1 => n11556, A2 => n11559, ZN => n10915);
   U13763 : MUX2_X1 port map( A => n10916, B => n10915, S => n20479, Z => 
                           n10917);
   U13764 : OAI21_X1 port map( B1 => n10918, B2 => n19564, A => n10917, ZN => 
                           n12232);
   U13765 : NAND2_X1 port map( A1 => n12230, A2 => n12232, ZN => n12048);
   U13766 : MUX2_X1 port map( A => n11523, B => n19999, S => n2470, Z => n10922
                           );
   U13767 : NOR2_X1 port map( A1 => n10922, A2 => n10921, ZN => n12223);
   U13768 : INV_X1 port map( A => n12121, ZN => n10944);
   U13769 : NAND2_X1 port map( A1 => n258, A2 => n10926, ZN => n10927);
   U13770 : NAND3_X1 port map( A1 => n11548, A2 => n258, A3 => n11549, ZN => 
                           n10929);
   U13771 : AND3_X2 port map( A1 => n10931, A2 => n10930, A3 => n10929, ZN => 
                           n12122);
   U13772 : INV_X1 port map( A => n12122, ZN => n12226);
   U13773 : NAND2_X1 port map( A1 => n10932, A2 => n11533, ZN => n10933);
   U13774 : NOR2_X1 port map( A1 => n20639, A2 => n10935, ZN => n10940);
   U13775 : OAI21_X1 port map( B1 => n11573, B2 => n19864, A => n10936, ZN => 
                           n10939);
   U13776 : NAND2_X1 port map( A1 => n11573, A2 => n11513, ZN => n10937);
   U13778 : INV_X1 port map( A => n12228, ZN => n10941);
   U13780 : XNOR2_X1 port map( A => n13058, B => n13580, ZN => n12791);
   U13781 : NAND2_X1 port map( A1 => n10946, A2 => n10693, ZN => n10996);
   U13782 : OAI21_X1 port map( B1 => n11284, B2 => n11283, A => n10693, ZN => 
                           n10948);
   U13783 : NAND2_X1 port map( A1 => n10948, A2 => n10947, ZN => n10949);
   U13784 : NAND2_X1 port map( A1 => n12130, A2 => n12126, ZN => n11760);
   U13785 : MUX2_X1 port map( A => n11010, B => n20470, S => n10951, Z => 
                           n10955);
   U13786 : NAND2_X1 port map( A1 => n3382, A2 => n10952, ZN => n10954);
   U13787 : MUX2_X1 port map( A => n10955, B => n10954, S => n10953, Z => 
                           n10956);
   U13788 : INV_X1 port map( A => n12127, ZN => n11701);
   U13789 : INV_X1 port map( A => n10957, ZN => n10959);
   U13791 : NAND2_X1 port map( A1 => n11176, A2 => n11178, ZN => n10965);
   U13792 : OAI211_X1 port map( C1 => n19878, C2 => n11178, A => n11174, B => 
                           n3789, ZN => n10964);
   U13793 : OAI211_X1 port map( C1 => n10966, C2 => n11178, A => n10965, B => 
                           n10964, ZN => n12128);
   U13794 : NOR2_X1 port map( A1 => n11586, A2 => n12128, ZN => n10967);
   U13795 : AND2_X1 port map( A1 => n12126, A2 => n12128, ZN => n10972);
   U13796 : AOI21_X1 port map( B1 => n11163, B2 => n20479, A => n11559, ZN => 
                           n10971);
   U13797 : OAI22_X1 port map( A1 => n19957, A2 => n19564, B1 => n10913, B2 => 
                           n11556, ZN => n10970);
   U13798 : OAI211_X2 port map( C1 => n11701, C2 => n11760, A => n10974, B => 
                           n10973, ZN => n13020);
   U13799 : XNOR2_X1 port map( A => n13020, B => n2164, ZN => n10975);
   U13800 : XNOR2_X1 port map( A => n12791, B => n10975, ZN => n10976);
   U13801 : XNOR2_X1 port map( A => n10977, B => n10976, ZN => n13901);
   U13802 : NOR2_X1 port map( A1 => n11292, A2 => n11294, ZN => n10982);
   U13803 : NOR2_X1 port map( A1 => n10980, A2 => n11290, ZN => n10981);
   U13804 : MUX2_X1 port map( A => n10982, B => n10981, S => n11403, Z => 
                           n10983);
   U13805 : NAND2_X1 port map( A1 => n10985, A2 => n11297, ZN => n10989);
   U13806 : OAI21_X1 port map( B1 => n11394, B2 => n11397, A => n10986, ZN => 
                           n10987);
   U13807 : NAND2_X1 port map( A1 => n10987, A2 => n11395, ZN => n10988);
   U13808 : NAND2_X1 port map( A1 => n11686, A2 => n11683, ZN => n11018);
   U13809 : NOR2_X1 port map( A1 => n11388, A2 => n10990, ZN => n10992);
   U13811 : MUX2_X1 port map( A => n10992, B => n10991, S => n11869, Z => 
                           n10994);
   U13812 : NOR2_X1 port map( A1 => n11871, A2 => n11390, ZN => n11385);
   U13813 : NAND2_X1 port map( A1 => n11385, A2 => n11302, ZN => n11874);
   U13814 : INV_X1 port map( A => n11874, ZN => n10993);
   U13815 : NAND2_X1 port map( A1 => n20462, A2 => n11922, ZN => n11007);
   U13816 : NOR2_X1 port map( A1 => n19851, A2 => n11278, ZN => n11002);
   U13817 : NOR2_X1 port map( A1 => n11277, A2 => n10688, ZN => n11001);
   U13818 : OAI21_X1 port map( B1 => n11002, B2 => n11001, A => n937, ZN => 
                           n11004);
   U13819 : NAND3_X1 port map( A1 => n11408, A2 => n11278, A3 => n11413, ZN => 
                           n11003);
   U13820 : NAND2_X1 port map( A1 => n11007, A2 => n12579, ZN => n11008);
   U13821 : AOI21_X1 port map( B1 => n11009, B2 => n3382, A => n11149, ZN => 
                           n11015);
   U13822 : NOR2_X1 port map( A1 => n11148, A2 => n11010, ZN => n11012);
   U13823 : OAI21_X1 port map( B1 => n11013, B2 => n11012, A => n11011, ZN => 
                           n11014);
   U13824 : OAI21_X1 port map( B1 => n11016, B2 => n11015, A => n11014, ZN => 
                           n11863);
   U13825 : INV_X1 port map( A => n12502, ZN => n11020);
   U13826 : NAND3_X1 port map( A1 => n11020, A2 => n12004, A3 => n201, ZN => 
                           n11022);
   U13827 : INV_X1 port map( A => n12499, ZN => n11019);
   U13828 : OAI211_X1 port map( C1 => n12497, C2 => n12500, A => n11022, B => 
                           n11021, ZN => n11024);
   U13829 : NOR2_X1 port map( A1 => n12345, A2 => n12500, ZN => n11023);
   U13830 : NAND2_X1 port map( A1 => n12419, A2 => n20351, ZN => n11025);
   U13831 : OAI21_X1 port map( B1 => n12419, B2 => n12084, A => n11025, ZN => 
                           n11028);
   U13832 : INV_X1 port map( A => n12416, ZN => n12418);
   U13833 : INV_X1 port map( A => n12422, ZN => n11603);
   U13834 : NOR2_X1 port map( A1 => n11603, A2 => n12084, ZN => n11026);
   U13835 : AOI22_X1 port map( A1 => n11026, A2 => n12419, B1 => n12415, B2 => 
                           n12084, ZN => n11027);
   U13836 : OAI21_X2 port map( B1 => n11028, B2 => n12418, A => n11027, ZN => 
                           n13657);
   U13837 : XNOR2_X1 port map( A => n11029, B => n13657, ZN => n13076);
   U13838 : INV_X1 port map( A => n13076, ZN => n11103);
   U13839 : INV_X1 port map( A => n12354, ZN => n11031);
   U13840 : NAND3_X1 port map( A1 => n12001, A2 => n12352, A3 => n11031, ZN => 
                           n11033);
   U13841 : XNOR2_X1 port map( A => n13715, B => n2344, ZN => n11064);
   U13842 : NOR2_X1 port map( A1 => n11034, A2 => n11439, ZN => n11036);
   U13843 : INV_X1 port map( A => n11035, ZN => n11119);
   U13844 : INV_X1 port map( A => n11037, ZN => n11436);
   U13845 : NOR3_X1 port map( A1 => n11435, A2 => n11440, A3 => n11436, ZN => 
                           n11891);
   U13846 : INV_X1 port map( A => n11038, ZN => n11040);
   U13847 : NAND2_X1 port map( A1 => n1039, A2 => n1317, ZN => n11039);
   U13848 : INV_X1 port map( A => n12261, ZN => n12563);
   U13849 : NAND2_X1 port map( A1 => n11428, A2 => n11105, ZN => n11043);
   U13850 : MUX2_X1 port map( A => n11043, B => n11042, S => n11041, Z => 
                           n11047);
   U13851 : NOR2_X1 port map( A1 => n11428, A2 => n1378, ZN => n11045);
   U13852 : NOR2_X1 port map( A1 => n19830, A2 => n11105, ZN => n11044);
   U13853 : AOI22_X1 port map( A1 => n11045, A2 => n11427, B1 => n11044, B2 => 
                           n11106, ZN => n11046);
   U13854 : NAND2_X1 port map( A1 => n11047, A2 => n11046, ZN => n11061);
   U13855 : OAI21_X1 port map( B1 => n11129, B2 => n11051, A => n19837, ZN => 
                           n11052);
   U13856 : OAI21_X2 port map( B1 => n11054, B2 => n19959, A => n11053, ZN => 
                           n12262);
   U13857 : OAI21_X1 port map( B1 => n12563, B2 => n12016, A => n12565, ZN => 
                           n11063);
   U13858 : NOR2_X1 port map( A1 => n11346, A2 => n11239, ZN => n11056);
   U13859 : AOI22_X1 port map( A1 => n11056, A2 => n11055, B1 => n11346, B2 => 
                           n11238, ZN => n11059);
   U13860 : NAND3_X1 port map( A1 => n11349, A2 => n11057, A3 => n11346, ZN => 
                           n11058);
   U13861 : OAI211_X1 port map( C1 => n11060, C2 => n11348, A => n11059, B => 
                           n11058, ZN => n12264);
   U13862 : INV_X1 port map( A => n11061, ZN => n12562);
   U13864 : XNOR2_X1 port map( A => n11064, B => n13321, ZN => n11101);
   U13865 : NAND2_X1 port map( A1 => n11943, A2 => n12441, ZN => n11066);
   U13866 : NOR2_X1 port map( A1 => n11066, A2 => n11065, ZN => n11068);
   U13867 : MUX2_X1 port map( A => n19505, B => n19913, S => n11495, Z => 
                           n11071);
   U13869 : INV_X1 port map( A => n11198, ZN => n11072);
   U13870 : AND2_X1 port map( A1 => n11072, A2 => n20539, ZN => n12252);
   U13871 : AOI21_X1 port map( B1 => n10745, B2 => n11210, A => n11483, ZN => 
                           n11075);
   U13872 : NAND2_X1 port map( A1 => n11073, A2 => n3500, ZN => n11074);
   U13874 : NAND2_X1 port map( A1 => n12250, A2 => n20153, ZN => n12570);
   U13875 : INV_X1 port map( A => n12570, ZN => n13144);
   U13876 : INV_X1 port map( A => n11076, ZN => n11218);
   U13877 : NAND2_X1 port map( A1 => n11218, A2 => n204, ZN => n11077);
   U13878 : NAND2_X1 port map( A1 => n11475, A2 => n11219, ZN => n11078);
   U13879 : INV_X1 port map( A => n12253, ZN => n13145);
   U13880 : NOR2_X1 port map( A1 => n11501, A2 => n11193, ZN => n11505);
   U13881 : NOR2_X1 port map( A1 => n11193, A2 => n11500, ZN => n11081);
   U13882 : INV_X1 port map( A => n11193, ZN => n11187);
   U13883 : INV_X1 port map( A => n11186, ZN => n11503);
   U13884 : MUX2_X1 port map( A => n11083, B => n11082, S => n11501, Z => 
                           n11084);
   U13886 : NAND2_X1 port map( A1 => n11112, A2 => n11458, ZN => n11086);
   U13887 : INV_X1 port map( A => n11452, ZN => n11089);
   U13888 : OAI22_X1 port map( A1 => n11089, A2 => n11110, B1 => n11455, B2 => 
                           n11454, ZN => n11090);
   U13889 : NOR2_X1 port map( A1 => n13147, A2 => n12255, ZN => n11092);
   U13890 : OAI21_X1 port map( B1 => n13146, B2 => n13145, A => n11092, ZN => 
                           n11099);
   U13891 : NAND3_X1 port map( A1 => n11209, A2 => n11201, A3 => n11094, ZN => 
                           n11096);
   U13892 : NAND3_X1 port map( A1 => n11445, A2 => n11202, A3 => n11444, ZN => 
                           n11095);
   U13893 : NAND4_X1 port map( A1 => n11097, A2 => n11448, A3 => n11096, A4 => 
                           n11095, ZN => n12254);
   U13894 : INV_X1 port map( A => n12254, ZN => n13141);
   U13895 : OAI21_X1 port map( B1 => n13141, B2 => n12258, A => n13147, ZN => 
                           n11098);
   U13896 : XNOR2_X1 port map( A => n13319, B => n13280, ZN => n11100);
   U13897 : XNOR2_X1 port map( A => n11101, B => n11100, ZN => n11102);
   U13898 : INV_X1 port map( A => n14780, ZN => n14077);
   U13899 : NOR2_X1 port map( A1 => n14077, A2 => n20518, ZN => n11319);
   U13901 : NOR2_X1 port map( A1 => n11106, A2 => n11105, ZN => n11107);
   U13902 : NAND2_X1 port map( A1 => n11452, A2 => n11110, ZN => n11111);
   U13903 : NAND2_X1 port map( A1 => n12138, A2 => n12137, ZN => n11139);
   U13904 : AND2_X1 port map( A1 => n11120, A2 => n11880, ZN => n11121);
   U13905 : OAI21_X1 port map( B1 => n11121, B2 => n11883, A => n85, ZN => 
                           n11123);
   U13906 : NAND2_X1 port map( A1 => n11121, A2 => n909, ZN => n11122);
   U13907 : NAND3_X1 port map( A1 => n12470, A2 => n11915, A3 => n12137, ZN => 
                           n11138);
   U13908 : NAND2_X1 port map( A1 => n20099, A2 => n11125, ZN => n11126);
   U13909 : NAND3_X1 port map( A1 => n205, A2 => n19837, A3 => n11131, ZN => 
                           n11135);
   U13910 : NOR2_X1 port map( A1 => n12463, A2 => n12386, ZN => n11136);
   U13911 : NAND2_X1 port map( A1 => n12470, A2 => n11136, ZN => n11137);
   U13912 : INV_X1 port map( A => n12281, ZN => n11167);
   U13913 : OAI21_X1 port map( B1 => n11148, B2 => n11147, A => n11149, ZN => 
                           n11154);
   U13914 : NAND2_X1 port map( A1 => n20470, A2 => n11149, ZN => n11151);
   U13916 : NAND2_X1 port map( A1 => n11557, A2 => n11559, ZN => n11554);
   U13917 : OR2_X1 port map( A1 => n11554, A2 => n20479, ZN => n11165);
   U13918 : NAND2_X1 port map( A1 => n19564, A2 => n10968, ZN => n11555);
   U13919 : OAI211_X1 port map( C1 => n11163, C2 => n20479, A => n10913, B => 
                           n11162, ZN => n11164);
   U13920 : AND3_X1 port map( A1 => n11555, A2 => n11165, A3 => n11164, ZN => 
                           n12279);
   U13921 : NAND2_X1 port map( A1 => n11717, A2 => n12279, ZN => n12044);
   U13922 : INV_X1 port map( A => n12044, ZN => n11166);
   U13923 : OAI21_X1 port map( B1 => n11167, B2 => n12040, A => n11166, ZN => 
                           n11181);
   U13924 : NAND2_X1 port map( A1 => n11171, A2 => n11532, ZN => n12035);
   U13925 : INV_X1 port map( A => n12035, ZN => n11172);
   U13926 : INV_X1 port map( A => n12279, ZN => n12042);
   U13927 : AOI21_X1 port map( B1 => n12282, B2 => n12042, A => n12040, ZN => 
                           n11180);
   U13928 : NOR2_X1 port map( A1 => n11176, A2 => n11175, ZN => n11179);
   U13929 : AND2_X1 port map( A1 => n12040, A2 => n12041, ZN => n11775);
   U13930 : XNOR2_X1 port map( A => n13330, B => n13833, ZN => n11229);
   U13931 : INV_X1 port map( A => n11182, ZN => n11183);
   U13932 : OAI22_X1 port map( A1 => n11183, A2 => n11564, B1 => n11566, B2 => 
                           n11469, ZN => n11184);
   U13933 : NAND2_X1 port map( A1 => n11184, A2 => n11567, ZN => n11185);
   U13935 : NOR2_X1 port map( A1 => n11500, A2 => n11188, ZN => n11189);
   U13937 : MUX2_X1 port map( A => n11193, B => n11192, S => n11191, Z => 
                           n11194);
   U13938 : AOI21_X1 port map( B1 => n11446, B2 => n19920, A => n11202, ZN => 
                           n11207);
   U13939 : INV_X1 port map( A => n11203, ZN => n11206);
   U13940 : INV_X1 port map( A => n11204, ZN => n11205);
   U13941 : OAI21_X1 port map( B1 => n11207, B2 => n11206, A => n11205, ZN => 
                           n11208);
   U13942 : NAND2_X1 port map( A1 => n11708, A2 => n12394, ZN => n12785);
   U13943 : INV_X1 port map( A => n12785, ZN => n11225);
   U13944 : NAND2_X1 port map( A1 => n3500, A2 => n11482, ZN => n11213);
   U13945 : NAND2_X1 port map( A1 => n11481, A2 => n11483, ZN => n11212);
   U13946 : MUX2_X1 port map( A => n11213, B => n11212, S => n19897, Z => 
                           n11214);
   U13947 : NAND2_X1 port map( A1 => n11217, A2 => n11475, ZN => n11221);
   U13948 : OAI211_X1 port map( C1 => n11474, C2 => n11222, A => n11221, B => 
                           n11220, ZN => n11930);
   U13949 : BUF_X2 port map( A => n11930, Z => n12473);
   U13950 : NOR2_X1 port map( A1 => n12478, A2 => n12473, ZN => n11223);
   U13951 : INV_X1 port map( A => n12784, ZN => n11224);
   U13952 : OAI21_X1 port map( B1 => n11225, B2 => n11224, A => n18355, ZN => 
                           n11227);
   U13953 : NAND3_X1 port map( A1 => n12785, A2 => n621, A3 => n12784, ZN => 
                           n11226);
   U13954 : NAND2_X1 port map( A1 => n11227, A2 => n11226, ZN => n11228);
   U13955 : XNOR2_X1 port map( A => n11229, B => n11228, ZN => n11318);
   U13956 : NOR2_X1 port map( A1 => n9883, A2 => n11231, ZN => n11232);
   U13957 : NOR2_X1 port map( A1 => n11235, A2 => n11234, ZN => n11243);
   U13958 : NAND2_X1 port map( A1 => n11237, A2 => n11236, ZN => n11242);
   U13959 : OAI21_X1 port map( B1 => n11239, B2 => n10798, A => n11238, ZN => 
                           n11241);
   U13960 : NOR2_X1 port map( A1 => n12381, A2 => n20191, ZN => n11270);
   U13961 : NOR2_X1 port map( A1 => n20191, A2 => n11243, ZN => n11251);
   U13962 : AOI21_X1 port map( B1 => n11373, B2 => n11244, A => n11376, ZN => 
                           n11246);
   U13963 : NOR2_X1 port map( A1 => n2861, A2 => n11330, ZN => n11245);
   U13964 : MUX2_X1 port map( A => n11246, B => n11245, S => n11377, Z => 
                           n11248);
   U13965 : INV_X1 port map( A => n11375, ZN => n11247);
   U13966 : MUX2_X1 port map( A => n11381, B => n11271, S => n11380, Z => 
                           n11250);
   U13967 : AOI22_X1 port map( A1 => n11252, A2 => n11251, B1 => n12269, B2 => 
                           n20497, ZN => n12271);
   U13969 : NAND2_X1 port map( A1 => n11253, A2 => n11255, ZN => n11258);
   U13970 : INV_X1 port map( A => n11258, ZN => n11262);
   U13971 : OAI21_X1 port map( B1 => n11321, B2 => n11255, A => n11254, ZN => 
                           n11261);
   U13972 : NAND2_X1 port map( A1 => n191, A2 => n11256, ZN => n11259);
   U13973 : MUX2_X1 port map( A => n11259, B => n11258, S => n11257, Z => 
                           n11260);
   U13974 : NOR2_X1 port map( A1 => n11267, A2 => n11263, ZN => n11336);
   U13975 : OAI21_X1 port map( B1 => n11343, B2 => n11264, A => n11337, ZN => 
                           n11268);
   U13976 : AND2_X1 port map( A1 => n11339, A2 => n9830, ZN => n11335);
   U13977 : OAI21_X1 port map( B1 => n12369, B2 => n12373, A => n12377, ZN => 
                           n11269);
   U13978 : OAI21_X1 port map( B1 => n11270, B2 => n12271, A => n11269, ZN => 
                           n13120);
   U13979 : NAND2_X1 port map( A1 => n11276, A2 => n11410, ZN => n11280);
   U13980 : OAI211_X1 port map( C1 => n11411, C2 => n11278, A => n11408, B => 
                           n11277, ZN => n11279);
   U13982 : OAI21_X1 port map( B1 => n11284, B2 => n9559, A => n11283, ZN => 
                           n11285);
   U13983 : OAI21_X1 port map( B1 => n11287, B2 => n11286, A => n11285, ZN => 
                           n11288);
   U13984 : MUX2_X1 port map( A => n11296, B => n11399, S => n11295, Z => 
                           n11301);
   U13985 : NAND2_X1 port map( A1 => n11297, A2 => n11399, ZN => n11299);
   U13986 : NAND2_X1 port map( A1 => n11394, A2 => n11398, ZN => n11298);
   U13987 : MUX2_X1 port map( A => n11299, B => n11298, S => n11395, Z => 
                           n11300);
   U13988 : INV_X1 port map( A => n12488, ZN => n12812);
   U13989 : NAND2_X1 port map( A1 => n11303, A2 => n11302, ZN => n11309);
   U13990 : NAND3_X1 port map( A1 => n11305, A2 => n11388, A3 => n11304, ZN => 
                           n11308);
   U13991 : NAND3_X1 port map( A1 => n20517, A2 => n11867, A3 => n20601, ZN => 
                           n11307);
   U13992 : OAI211_X1 port map( C1 => n12399, C2 => n12807, A => n12812, B => 
                           n12487, ZN => n11310);
   U13993 : OAI211_X1 port map( C1 => n12807, C2 => n11693, A => n11911, B => 
                           n11310, ZN => n13431);
   U13994 : XNOR2_X1 port map( A => n13120, B => n13431, ZN => n13329);
   U13995 : INV_X1 port map( A => n13329, ZN => n11316);
   U13996 : NOR2_X1 port map( A1 => n12754, A2 => n12759, ZN => n12757);
   U13997 : OAI21_X1 port map( B1 => n11315, B2 => n12757, A => n11314, ZN => 
                           n13079);
   U13998 : XNOR2_X1 port map( A => n13031, B => n13079, ZN => n11965);
   U13999 : XNOR2_X1 port map( A => n11316, B => n11965, ZN => n11317);
   U14002 : AOI22_X1 port map( A1 => n191, A2 => n11324, B1 => n11323, B2 => 
                           n11327, ZN => n11326);
   U14003 : INV_X1 port map( A => n11709, ZN => n12311);
   U14004 : OAI21_X1 port map( B1 => n11331, B2 => n2611, A => n2861, ZN => 
                           n11334);
   U14005 : MUX2_X1 port map( A => n11330, B => n11329, S => n11332, Z => 
                           n11333);
   U14006 : NAND2_X1 port map( A1 => n12311, A2 => n20486, ZN => n11363);
   U14007 : NAND2_X1 port map( A1 => n11341, A2 => n11340, ZN => n11342);
   U14008 : AOI21_X1 port map( B1 => n11343, B2 => n11265, A => n11342, ZN => 
                           n11344);
   U14009 : MUX2_X1 port map( A => n11347, B => n11348, S => n11346, Z => 
                           n11354);
   U14011 : NAND2_X1 port map( A1 => n11355, A2 => n11239, ZN => n11351);
   U14012 : MUX2_X1 port map( A => n11352, B => n11351, S => n11350, Z => 
                           n11353);
   U14013 : NAND2_X1 port map( A1 => n11358, A2 => n19949, ZN => n11361);
   U14014 : NAND2_X1 port map( A1 => n11367, A2 => n11366, ZN => n11368);
   U14015 : MUX2_X1 port map( A => n12312, B => n12148, S => n19952, Z => 
                           n11370);
   U14016 : NOR2_X1 port map( A1 => n11370, A2 => n12311, ZN => n11371);
   U14017 : INV_X1 port map( A => n13099, ZN => n11416);
   U14018 : NAND2_X1 port map( A1 => n202, A2 => n11377, ZN => n11374);
   U14019 : NAND2_X1 port map( A1 => n11377, A2 => n11376, ZN => n11379);
   U14020 : AOI21_X1 port map( B1 => n11379, B2 => n202, A => n11378, ZN => 
                           n12548);
   U14022 : NOR2_X1 port map( A1 => n12542, A2 => n12543, ZN => n12310);
   U14023 : INV_X1 port map( A => n11385, ZN => n11386);
   U14025 : NAND2_X1 port map( A1 => n11388, A2 => n11870, ZN => n11392);
   U14026 : MUX2_X1 port map( A => n20517, B => n11866, S => n11389, Z => 
                           n11391);
   U14027 : MUX2_X1 port map( A => n11399, B => n11397, S => n11394, Z => 
                           n11396);
   U14028 : NAND3_X1 port map( A1 => n11399, A2 => n11398, A3 => n11397, ZN => 
                           n11400);
   U14029 : NOR2_X1 port map( A1 => n10978, A2 => n11405, ZN => n11407);
   U14030 : AOI22_X1 port map( A1 => n12310, A2 => n2160, B1 => n11795, B2 => 
                           n12305, ZN => n11415);
   U14031 : INV_X1 port map( A => n11411, ZN => n11412);
   U14032 : AND2_X1 port map( A1 => n11413, A2 => n937, ZN => n12549);
   U14033 : NAND2_X1 port map( A1 => n11415, A2 => n11414, ZN => n13756);
   U14034 : XNOR2_X1 port map( A => n11416, B => n13756, ZN => n13347);
   U14035 : NAND2_X1 port map( A1 => n11419, A2 => n1680, ZN => n11422);
   U14036 : INV_X1 port map( A => n12524, ZN => n12165);
   U14037 : AOI21_X1 port map( B1 => n11425, B2 => n11424, A => n19830, ZN => 
                           n11434);
   U14038 : NOR2_X1 port map( A1 => n11427, A2 => n1378, ZN => n11433);
   U14039 : OAI211_X1 port map( C1 => n19830, C2 => n11430, A => n11429, B => 
                           n11428, ZN => n11432);
   U14041 : INV_X1 port map( A => n12167, ZN => n12520);
   U14042 : MUX2_X1 port map( A => n11438, B => n11436, S => n11435, Z => 
                           n11442);
   U14043 : NAND2_X1 port map( A1 => n11445, A2 => n11444, ZN => n11447);
   U14044 : NAND3_X1 port map( A1 => n11456, A2 => n11455, A3 => n11454, ZN => 
                           n11457);
   U14045 : MUX2_X1 port map( A => n11883, B => n11880, S => n11884, Z => 
                           n11463);
   U14046 : INV_X1 port map( A => n12168, ZN => n11464);
   U14047 : NAND2_X1 port map( A1 => n898, A2 => n11469, ZN => n11468);
   U14048 : NAND2_X1 port map( A1 => n11467, A2 => n11466, ZN => n11471);
   U14049 : MUX2_X1 port map( A => n11468, B => n11471, S => n11568, Z => 
                           n11473);
   U14050 : NAND2_X1 port map( A1 => n11471, A2 => n11470, ZN => n11472);
   U14051 : OAI211_X1 port map( C1 => n11481, C2 => n11480, A => n11486, B => 
                           n11479, ZN => n11485);
   U14052 : NAND3_X1 port map( A1 => n11483, A2 => n20233, A3 => n11482, ZN => 
                           n11484);
   U14053 : OAI211_X2 port map( C1 => n11486, C2 => n11487, A => n11485, B => 
                           n11484, ZN => n12534);
   U14054 : NAND2_X1 port map( A1 => n19719, A2 => n3051, ZN => n11490);
   U14055 : NAND2_X1 port map( A1 => n20539, A2 => n11493, ZN => n11497);
   U14056 : NOR2_X1 port map( A1 => n11495, A2 => n11494, ZN => n11496);
   U14057 : NAND2_X1 port map( A1 => n11500, A2 => n11499, ZN => n11504);
   U14058 : MUX2_X1 port map( A => n11504, B => n11502, S => n11501, Z => 
                           n11508);
   U14059 : NOR2_X1 port map( A1 => n11504, A2 => n11503, ZN => n11506);
   U14060 : NOR2_X1 port map( A1 => n11506, A2 => n11505, ZN => n11507);
   U14061 : NAND2_X1 port map( A1 => n11508, A2 => n11507, ZN => n12532);
   U14062 : MUX2_X1 port map( A => n12535, B => n243, S => n12534, Z => n11519)
                           ;
   U14063 : NAND2_X1 port map( A1 => n11512, A2 => n20639, ZN => n11518);
   U14065 : XNOR2_X1 port map( A => n13569, B => n13347, ZN => n11593);
   U14066 : NOR2_X1 port map( A1 => n11528, A2 => n11521, ZN => n11525);
   U14067 : NOR2_X1 port map( A1 => n11522, A2 => n11527, ZN => n11524);
   U14068 : NAND3_X1 port map( A1 => n11528, A2 => n11527, A3 => n11526, ZN => 
                           n11529);
   U14069 : OAI21_X1 port map( B1 => n11531, B2 => n11530, A => n11529, ZN => 
                           n11742);
   U14070 : NOR2_X2 port map( A1 => n11741, A2 => n11742, ZN => n12299);
   U14072 : NAND2_X1 port map( A1 => n731, A2 => n11538, ZN => n11541);
   U14074 : MUX2_X1 port map( A => n11549, B => n11548, S => n11547, Z => 
                           n11551);
   U14076 : AOI21_X1 port map( B1 => n11555, B2 => n11554, A => n11553, ZN => 
                           n11562);
   U14077 : NAND2_X1 port map( A1 => n11557, A2 => n11556, ZN => n11560);
   U14078 : AOI21_X1 port map( B1 => n11560, B2 => n11559, A => n19564, ZN => 
                           n11561);
   U14079 : INV_X1 port map( A => n11563, ZN => n12304);
   U14080 : NOR2_X1 port map( A1 => n12299, A2 => n11782, ZN => n11739);
   U14081 : AOI21_X1 port map( B1 => n11565, B2 => n11564, A => n927, ZN => 
                           n11744);
   U14082 : NAND2_X1 port map( A1 => n11567, A2 => n927, ZN => n11571);
   U14083 : NAND2_X1 port map( A1 => n11569, A2 => n11568, ZN => n11570);
   U14084 : AOI21_X1 port map( B1 => n11571, B2 => n11570, A => n898, ZN => 
                           n11740);
   U14085 : AND2_X1 port map( A1 => n12304, A2 => n12274, ZN => n11578);
   U14086 : INV_X1 port map( A => n12033, ZN => n11577);
   U14087 : INV_X1 port map( A => n13063, ZN => n11585);
   U14088 : NAND2_X1 port map( A1 => n12281, A2 => n12041, ZN => n11581);
   U14089 : AND2_X1 port map( A1 => n11580, A2 => n11581, ZN => n11584);
   U14090 : OAI21_X1 port map( B1 => n11582, B2 => n11776, A => n12278, ZN => 
                           n11583);
   U14091 : XNOR2_X1 port map( A => n11585, B => n12863, ZN => n11862);
   U14092 : INV_X1 port map( A => n12128, ZN => n11642);
   U14093 : OAI21_X1 port map( B1 => n882, B2 => n12126, A => n12130, ZN => 
                           n11588);
   U14094 : INV_X1 port map( A => n11586, ZN => n11763);
   U14095 : NAND2_X1 port map( A1 => n11588, A2 => n11587, ZN => n11589);
   U14096 : XNOR2_X1 port map( A => n13425, B => n1840, ZN => n11591);
   U14097 : XNOR2_X1 port map( A => n11862, B => n11591, ZN => n11592);
   U14098 : NAND2_X1 port map( A1 => n14216, A2 => n14781, ZN => n14852);
   U14099 : INV_X1 port map( A => n14852, ZN => n11594);
   U14100 : AND2_X1 port map( A1 => n12408, A2 => n12389, ZN => n12756);
   U14101 : NOR2_X1 port map( A1 => n12409, A2 => n12759, ZN => n11595);
   U14102 : NOR2_X1 port map( A1 => n12389, A2 => n12407, ZN => n12755);
   U14103 : XNOR2_X1 port map( A => n19792, B => n19027, ZN => n11609);
   U14104 : INV_X1 port map( A => n11951, ZN => n11955);
   U14105 : INV_X1 port map( A => n11659, ZN => n11600);
   U14106 : NAND3_X1 port map( A1 => n11955, A2 => n1578, A3 => n11600, ZN => 
                           n11601);
   U14107 : NOR2_X1 port map( A1 => n11602, A2 => n20351, ZN => n12082);
   U14110 : NAND2_X1 port map( A1 => n11605, A2 => n12084, ZN => n11606);
   U14111 : XNOR2_X1 port map( A => n13368, B => n13277, ZN => n13582);
   U14112 : XNOR2_X1 port map( A => n13582, B => n11609, ZN => n11626);
   U14114 : NAND2_X1 port map( A1 => n12684, A2 => n12648, ZN => n11610);
   U14115 : MUX2_X1 port map( A => n11611, B => n11610, S => n12686, Z => 
                           n11612);
   U14116 : INV_X1 port map( A => n13707, ZN => n13019);
   U14117 : INV_X1 port map( A => n12449, ZN => n12635);
   U14118 : NAND2_X1 port map( A1 => n11948, A2 => n12642, ZN => n11617);
   U14119 : INV_X1 port map( A => n12455, ZN => n12640);
   U14120 : NOR2_X1 port map( A1 => n12640, A2 => n12635, ZN => n11616);
   U14121 : NAND3_X1 port map( A1 => n20458, A2 => n2256, A3 => n12450, ZN => 
                           n11615);
   U14122 : NAND2_X1 port map( A1 => n12637, A2 => n12452, ZN => n11614);
   U14124 : XNOR2_X1 port map( A => n13019, B => n13774, ZN => n13233);
   U14125 : NOR2_X1 port map( A1 => n12634, A2 => n11618, ZN => n11620);
   U14126 : NAND2_X1 port map( A1 => n11618, A2 => n12630, ZN => n11619);
   U14127 : MUX2_X1 port map( A => n11942, B => n12437, S => n12440, Z => 
                           n11624);
   U14128 : NOR2_X1 port map( A1 => n12440, A2 => n11942, ZN => n11623);
   U14129 : XNOR2_X1 port map( A => n13706, B => n13776, ZN => n13475);
   U14130 : XNOR2_X1 port map( A => n13233, B => n13475, ZN => n11625);
   U14131 : AOI21_X1 port map( B1 => n12603, B2 => n12237, A => n12072, ZN => 
                           n11631);
   U14132 : INV_X1 port map( A => n11628, ZN => n11629);
   U14133 : NAND2_X1 port map( A1 => n12242, A2 => n12240, ZN => n12054);
   U14134 : INV_X1 port map( A => n12054, ZN => n11635);
   U14135 : INV_X1 port map( A => n12616, ZN => n12059);
   U14136 : XNOR2_X1 port map( A => n12986, B => n13734, ZN => n11641);
   U14137 : INV_X1 port map( A => n12201, ZN => n12593);
   U14138 : INV_X1 port map( A => n12200, ZN => n12592);
   U14139 : OAI211_X1 port map( C1 => n11637, C2 => n12593, A => n193, B => 
                           n12592, ZN => n11636);
   U14140 : OAI211_X1 port map( C1 => n11978, C2 => n11637, A => n11636, B => 
                           n11979, ZN => n13029);
   U14141 : NOR2_X1 port map( A1 => n12211, A2 => n19726, ZN => n12214);
   U14142 : XNOR2_X1 port map( A => n13029, B => n11640, ZN => n13237);
   U14143 : XNOR2_X1 port map( A => n11641, B => n13237, ZN => n11655);
   U14144 : NAND2_X1 port map( A1 => n12129, A2 => n12128, ZN => n11702);
   U14145 : OR2_X1 port map( A1 => n11702, A2 => n12126, ZN => n11645);
   U14146 : NAND4_X1 port map( A1 => n11703, A2 => n11645, A3 => n11644, A4 => 
                           n11643, ZN => n12671);
   U14147 : INV_X1 port map( A => n12671, ZN => n13391);
   U14148 : NAND2_X1 port map( A1 => n12121, A2 => n12230, ZN => n12049);
   U14150 : INV_X1 port map( A => n12232, ZN => n11646);
   U14151 : OAI21_X1 port map( B1 => n12049, B2 => n19694, A => n11648, ZN => 
                           n13484);
   U14152 : XNOR2_X1 port map( A => n13391, B => n13484, ZN => n13612);
   U14153 : NOR2_X1 port map( A1 => n12180, A2 => n256, ZN => n11652);
   U14154 : NAND2_X1 port map( A1 => n11841, A2 => n20427, ZN => n11651);
   U14155 : XNOR2_X1 port map( A => n13612, B => n11653, ZN => n11654);
   U14156 : XNOR2_X1 port map( A => n11654, B => n11655, ZN => n14806);
   U14158 : NOR2_X1 port map( A1 => n11828, A2 => n11829, ZN => n11657);
   U14159 : MUX2_X1 port map( A => n11659, B => n11830, S => n11829, Z => 
                           n11660);
   U14160 : INV_X1 port map( A => n13134, ZN => n12087);
   U14161 : XNOR2_X1 port map( A => n12087, B => n13572, ZN => n13464);
   U14162 : MUX2_X1 port map( A => n12008, B => n12509, S => n12506, Z => 
                           n11663);
   U14163 : INV_X1 port map( A => n12359, ZN => n11661);
   U14165 : NAND2_X1 port map( A1 => n11992, A2 => n965, ZN => n11664);
   U14166 : XNOR2_X1 port map( A => n12940, B => n13651, ZN => n13243);
   U14167 : NAND2_X1 port map( A1 => n11841, A2 => n11670, ZN => n11671);
   U14168 : MUX2_X1 port map( A => n12179, B => n11673, S => n12180, Z => 
                           n11675);
   U14169 : MUX2_X1 port map( A => n12514, B => n11997, S => n11995, Z => 
                           n11677);
   U14170 : XNOR2_X1 port map( A => n13397, B => n13687, ZN => n11681);
   U14171 : MUX2_X1 port map( A => n201, B => n12499, S => n12004, Z => n11679)
                           ;
   U14172 : XNOR2_X1 port map( A => n12979, B => n19243, ZN => n11680);
   U14173 : XNOR2_X1 port map( A => n11681, B => n11680, ZN => n11682);
   U14174 : INV_X1 port map( A => n14806, ZN => n14811);
   U14175 : NAND2_X1 port map( A1 => n11863, A2 => n11922, ZN => n12578);
   U14176 : INV_X1 port map( A => n12578, ZN => n11685);
   U14177 : NOR2_X1 port map( A1 => n11926, A2 => n12577, ZN => n11684);
   U14179 : NAND2_X1 port map( A1 => n11686, A2 => n11922, ZN => n11865);
   U14180 : INV_X1 port map( A => n11863, ZN => n11923);
   U14181 : NAND2_X1 port map( A1 => n11865, A2 => n11863, ZN => n11687);
   U14182 : NAND2_X1 port map( A1 => n11687, A2 => n11926, ZN => n11688);
   U14183 : OAI21_X1 port map( B1 => n12229, B2 => n12122, A => n12228, ZN => 
                           n11690);
   U14184 : NAND2_X1 port map( A1 => n11690, A2 => n12121, ZN => n11691);
   U14185 : XNOR2_X1 port map( A => n13622, B => n13193, ZN => n11698);
   U14186 : NAND2_X1 port map( A1 => n11911, A2 => n11693, ZN => n11696);
   U14187 : NAND2_X1 port map( A1 => n12488, A2 => n12809, ZN => n11694);
   U14188 : NAND2_X1 port map( A1 => n11694, A2 => n12811, ZN => n11695);
   U14189 : XNOR2_X1 port map( A => n13339, B => n18433, ZN => n11697);
   U14190 : XNOR2_X1 port map( A => n11698, B => n11697, ZN => n11716);
   U14191 : INV_X1 port map( A => n12386, ZN => n12384);
   U14192 : NAND2_X1 port map( A1 => n12384, A2 => n12137, ZN => n12383);
   U14193 : INV_X1 port map( A => n12138, ZN => n12468);
   U14194 : NOR2_X1 port map( A1 => n12138, A2 => n857, ZN => n11699);
   U14195 : OR3_X1 port map( A1 => n12138, A2 => n12470, A3 => n11915, ZN => 
                           n11700);
   U14198 : XNOR2_X1 port map( A => n13222, B => n13623, ZN => n11714);
   U14199 : NAND2_X1 port map( A1 => n12478, A2 => n11930, ZN => n11706);
   U14200 : NAND2_X1 port map( A1 => n11706, A2 => n12142, ZN => n11707);
   U14201 : INV_X1 port map( A => n12312, ZN => n12154);
   U14202 : INV_X1 port map( A => n12152, ZN => n11710);
   U14203 : AOI21_X1 port map( B1 => n12153, B2 => n20186, A => n11710, ZN => 
                           n11713);
   U14204 : INV_X1 port map( A => n12148, ZN => n12155);
   U14205 : OAI21_X1 port map( B1 => n12148, B2 => n19952, A => n11711, ZN => 
                           n12315);
   U14206 : XNOR2_X1 port map( A => n13138, B => n13048, ZN => n13227);
   U14207 : INV_X1 port map( A => n13227, ZN => n13727);
   U14208 : XNOR2_X1 port map( A => n13727, B => n11714, ZN => n11715);
   U14210 : NAND2_X1 port map( A1 => n12041, A2 => n12279, ZN => n11721);
   U14211 : OR2_X1 port map( A1 => n11717, A2 => n12280, ZN => n11777);
   U14212 : OAI21_X1 port map( B1 => n12283, B2 => n11776, A => n11777, ZN => 
                           n11718);
   U14213 : NOR2_X1 port map( A1 => n12281, A2 => n12040, ZN => n11719);
   U14214 : NAND2_X1 port map( A1 => n11719, A2 => n876, ZN => n11720);
   U14215 : XNOR2_X1 port map( A => n13491, B => n18170, ZN => n11724);
   U14216 : NAND2_X1 port map( A1 => n12634, A2 => n11618, ZN => n11962);
   U14217 : NAND2_X1 port map( A1 => n12630, A2 => n11722, ZN => n11961);
   U14218 : NAND3_X1 port map( A1 => n11961, A2 => n12632, A3 => n1371, ZN => 
                           n11723);
   U14219 : XNOR2_X1 port map( A => n11724, B => n13517, ZN => n11729);
   U14220 : NOR2_X1 port map( A1 => n12267, A2 => n12262, ZN => n11725);
   U14221 : INV_X1 port map( A => n11726, ZN => n11727);
   U14222 : XNOR2_X1 port map( A => n11729, B => n13248, ZN => n11756);
   U14223 : NAND2_X1 port map( A1 => n12373, A2 => n20191, ZN => n11855);
   U14224 : INV_X1 port map( A => n11855, ZN => n11731);
   U14225 : INV_X1 port map( A => n11856, ZN => n12371);
   U14226 : XNOR2_X1 port map( A => n13745, B => n13642, ZN => n11754);
   U14227 : INV_X1 port map( A => n13149, ZN => n11734);
   U14228 : NAND2_X1 port map( A1 => n244, A2 => n12254, ZN => n11733);
   U14229 : NOR2_X1 port map( A1 => n13146, A2 => n20153, ZN => n11735);
   U14230 : NOR2_X1 port map( A1 => n12029, A2 => n12304, ZN => n11738);
   U14231 : INV_X1 port map( A => n12275, ZN => n12272);
   U14232 : AOI22_X1 port map( A1 => n11739, A2 => n12274, B1 => n11738, B2 => 
                           n12272, ZN => n11752);
   U14233 : INV_X1 port map( A => n12299, ZN => n12028);
   U14234 : INV_X1 port map( A => n11740, ZN => n11749);
   U14235 : INV_X1 port map( A => n11741, ZN => n11746);
   U14236 : INV_X1 port map( A => n11742, ZN => n11743);
   U14237 : AND2_X1 port map( A1 => n11744, A2 => n11743, ZN => n11745);
   U14238 : NAND2_X1 port map( A1 => n11746, A2 => n11745, ZN => n11747);
   U14239 : OAI211_X1 port map( C1 => n12028, C2 => n11749, A => n11748, B => 
                           n11747, ZN => n11750);
   U14240 : NAND2_X1 port map( A1 => n11750, A2 => n920, ZN => n11751);
   U14241 : NAND2_X1 port map( A1 => n11752, A2 => n11751, ZN => n12846);
   U14242 : XNOR2_X1 port map( A => n13695, B => n12846, ZN => n11753);
   U14243 : XNOR2_X1 port map( A => n11754, B => n11753, ZN => n11755);
   U14244 : NOR2_X1 port map( A1 => n14807, A2 => n14593, ZN => n14809);
   U14245 : INV_X1 port map( A => n14593, ZN => n14590);
   U14247 : INV_X1 port map( A => n12543, ZN => n11757);
   U14248 : NAND2_X1 port map( A1 => n11795, A2 => n12543, ZN => n11758);
   U14249 : AOI21_X1 port map( B1 => n11760, B2 => n11759, A => n882, ZN => 
                           n11767);
   U14250 : INV_X1 port map( A => n11761, ZN => n11762);
   U14251 : NAND2_X1 port map( A1 => n11763, A2 => n11762, ZN => n11765);
   U14252 : NOR2_X1 port map( A1 => n882, A2 => n12129, ZN => n11764);
   U14253 : NOR2_X1 port map( A1 => n11765, A2 => n11764, ZN => n11766);
   U14254 : NOR2_X1 port map( A1 => n11767, A2 => n11766, ZN => n12077);
   U14255 : XNOR2_X1 port map( A => n13717, B => n12077, ZN => n13153);
   U14256 : INV_X1 port map( A => n13153, ZN => n13499);
   U14257 : OAI21_X1 port map( B1 => n11768, B2 => n12522, A => n12525, ZN => 
                           n11771);
   U14258 : NOR2_X1 port map( A1 => n12528, A2 => n12288, ZN => n12292);
   U14259 : NAND2_X1 port map( A1 => n12165, A2 => n182, ZN => n11770);
   U14260 : XNOR2_X1 port map( A => n19697, B => n13255, ZN => n13714);
   U14261 : NAND2_X1 port map( A1 => n12311, A2 => n20186, ZN => n11773);
   U14263 : NOR2_X1 port map( A1 => n11777, A2 => n12281, ZN => n11778);
   U14264 : NOR2_X1 port map( A1 => n3801, A2 => n11778, ZN => n11779);
   U14265 : XNOR2_X1 port map( A => n13601, B => n13539, ZN => n11787);
   U14266 : OAI211_X1 port map( C1 => n12029, C2 => n11782, A => n12028, B => 
                           n11781, ZN => n11785);
   U14267 : INV_X1 port map( A => n12029, ZN => n12300);
   U14268 : OAI21_X1 port map( B1 => n12300, B2 => n12298, A => n12299, ZN => 
                           n11784);
   U14269 : NOR2_X1 port map( A1 => n12300, A2 => n11782, ZN => n11783);
   U14270 : XNOR2_X1 port map( A => n13602, B => n18284, ZN => n11786);
   U14271 : XNOR2_X1 port map( A => n11787, B => n11786, ZN => n11788);
   U14272 : NOR2_X1 port map( A1 => n907, A2 => n12167, ZN => n11794);
   U14273 : INV_X1 port map( A => n11795, ZN => n11800);
   U14274 : OAI211_X1 port map( C1 => n11977, C2 => n250, A => n11796, B => 
                           n2160, ZN => n11799);
   U14275 : XNOR2_X1 port map( A => n13126, B => n13810, ZN => n13641);
   U14276 : XNOR2_X1 port map( A => n13641, B => n11801, ZN => n11819);
   U14277 : INV_X1 port map( A => n12807, ZN => n12490);
   U14278 : OAI21_X1 port map( B1 => n12812, B2 => n12811, A => n953, ZN => 
                           n11802);
   U14279 : NAND2_X1 port map( A1 => n12811, A2 => n12809, ZN => n12397);
   U14280 : MUX2_X1 port map( A => n12490, B => n11802, S => n12397, Z => 
                           n11803);
   U14282 : INV_X1 port map( A => n13519, ZN => n11816);
   U14283 : NAND3_X1 port map( A1 => n11810, A2 => n11809, A3 => n11808, ZN => 
                           n11812);
   U14284 : INV_X1 port map( A => n12209, ZN => n12213);
   U14285 : OAI21_X1 port map( B1 => n11812, B2 => n11811, A => n2428, ZN => 
                           n11815);
   U14286 : NAND3_X1 port map( A1 => n12209, A2 => n12206, A3 => n19726, ZN => 
                           n11813);
   U14287 : OAI211_X2 port map( C1 => n11815, C2 => n12065, A => n11814, B => 
                           n11813, ZN => n13351);
   U14288 : XNOR2_X1 port map( A => n13351, B => n11816, ZN => n13447);
   U14289 : INV_X1 port map( A => n13447, ZN => n13375);
   U14290 : XNOR2_X1 port map( A => n13375, B => n11817, ZN => n11818);
   U14291 : INV_X1 port map( A => n12513, ZN => n11996);
   U14292 : NAND2_X1 port map( A1 => n13275, A2 => n11820, ZN => n11822);
   U14293 : NAND2_X1 port map( A1 => n12514, A2 => n11995, ZN => n11821);
   U14294 : OAI21_X1 port map( B1 => n11996, B2 => n11995, A => n11823, ZN => 
                           n13404);
   U14295 : AOI21_X1 port map( B1 => n12339, B2 => n11990, A => n11992, ZN => 
                           n11826);
   U14296 : NAND3_X1 port map( A1 => n12338, A2 => n11974, A3 => n12335, ZN => 
                           n11825);
   U14297 : OAI211_X1 port map( C1 => n12338, C2 => n11826, A => n11825, B => 
                           n11824, ZN => n13108);
   U14298 : XNOR2_X1 port map( A => n13404, B => n13108, ZN => n13440);
   U14299 : NOR2_X1 port map( A1 => n11827, A2 => n11829, ZN => n11833);
   U14300 : OAI21_X1 port map( B1 => n11952, B2 => n11828, A => n11951, ZN => 
                           n11832);
   U14301 : NAND2_X1 port map( A1 => n12509, A2 => n12009, ZN => n11836);
   U14302 : NAND2_X1 port map( A1 => n12008, A2 => n11836, ZN => n11838);
   U14303 : NAND2_X1 port map( A1 => n12507, A2 => n12508, ZN => n11837);
   U14304 : NAND2_X1 port map( A1 => n11838, A2 => n11837, ZN => n11839);
   U14305 : NAND2_X1 port map( A1 => n11840, A2 => n11839, ZN => n13405);
   U14306 : XNOR2_X1 port map( A => n13843, B => n13405, ZN => n12993);
   U14307 : NAND2_X1 port map( A1 => n252, A2 => n256, ZN => n11842);
   U14308 : AOI21_X1 port map( B1 => n11843, B2 => n11842, A => n12181, ZN => 
                           n11848);
   U14309 : INV_X1 port map( A => n11844, ZN => n11846);
   U14310 : OAI21_X1 port map( B1 => n11846, B2 => n252, A => n11845, ZN => 
                           n11847);
   U14311 : XNOR2_X1 port map( A => n13409, B => n13711, ZN => n11850);
   U14312 : XNOR2_X1 port map( A => n13715, B => n18075, ZN => n11849);
   U14313 : XNOR2_X1 port map( A => n11850, B => n11849, ZN => n11851);
   U14314 : AND2_X1 port map( A1 => n12374, A2 => n20191, ZN => n11853);
   U14315 : NAND2_X1 port map( A1 => n12381, A2 => n11853, ZN => n11854);
   U14316 : OAI21_X1 port map( B1 => n12381, B2 => n11855, A => n11854, ZN => 
                           n11858);
   U14317 : NOR2_X1 port map( A1 => n13147, A2 => n13141, ZN => n12251);
   U14318 : INV_X1 port map( A => n12251, ZN => n11860);
   U14319 : AOI21_X1 port map( B1 => n13147, B2 => n12255, A => n13145, ZN => 
                           n11859);
   U14320 : NAND2_X1 port map( A1 => n11860, A2 => n11859, ZN => n11861);
   U14321 : NOR2_X1 port map( A1 => n12258, A2 => n20153, ZN => n12573);
   U14322 : XNOR2_X1 port map( A => n13064, B => n12471, ZN => n13428);
   U14323 : NAND2_X1 port map( A1 => n20462, A2 => n11863, ZN => n11864);
   U14324 : NAND2_X1 port map( A1 => n11865, A2 => n11864, ZN => n11878);
   U14325 : NAND3_X1 port map( A1 => n20517, A2 => n11866, A3 => n20160, ZN => 
                           n11873);
   U14326 : NAND2_X1 port map( A1 => n11870, A2 => n11867, ZN => n11868);
   U14327 : OAI211_X1 port map( C1 => n20160, C2 => n11870, A => n11869, B => 
                           n11868, ZN => n11872);
   U14328 : NAND3_X1 port map( A1 => n11874, A2 => n11873, A3 => n11872, ZN => 
                           n11875);
   U14329 : NAND2_X1 port map( A1 => n11926, A2 => n11875, ZN => n11876);
   U14330 : OAI21_X1 port map( B1 => n20462, B2 => n11926, A => n11876, ZN => 
                           n11877);
   U14331 : XNOR2_X1 port map( A => n13848, B => n345, ZN => n11899);
   U14332 : INV_X1 port map( A => n11879, ZN => n11890);
   U14333 : OAI21_X1 port map( B1 => n11881, B2 => n11880, A => n85, ZN => 
                           n11889);
   U14334 : NOR2_X1 port map( A1 => n11883, A2 => n85, ZN => n11885);
   U14335 : AOI22_X1 port map( A1 => n11887, A2 => n11886, B1 => n11885, B2 => 
                           n909, ZN => n11888);
   U14336 : NOR3_X1 port map( A1 => n11892, A2 => n11891, A3 => n12262, ZN => 
                           n12568);
   U14337 : MUX2_X1 port map( A => n3401, B => n12630, S => n12631, Z => n11897
                           );
   U14338 : XNOR2_X1 port map( A => n13422, B => n13686, ZN => n11898);
   U14339 : XNOR2_X1 port map( A => n11899, B => n11898, ZN => n11900);
   U14340 : OAI21_X1 port map( B1 => n12148, B2 => n20186, A => n12313, ZN => 
                           n11907);
   U14341 : NAND2_X1 port map( A1 => n11709, A2 => n12312, ZN => n11903);
   U14343 : AOI21_X1 port map( B1 => n11905, B2 => n11710, A => n11904, ZN => 
                           n11906);
   U14344 : NOR2_X1 port map( A1 => n12807, A2 => n12811, ZN => n11909);
   U14345 : MUX2_X1 port map( A => n11910, B => n11909, S => n12487, Z => 
                           n11914);
   U14347 : NOR2_X2 port map( A1 => n11914, A2 => n11913, ZN => n13230);
   U14348 : XNOR2_X1 port map( A => n12859, B => n13230, ZN => n13005);
   U14349 : INV_X1 port map( A => n13005, ZN => n11929);
   U14350 : INV_X1 port map( A => n12470, ZN => n12139);
   U14351 : NOR2_X1 port map( A1 => n12139, A2 => n12463, ZN => n11921);
   U14352 : OAI21_X1 port map( B1 => n11915, B2 => n12137, A => n12138, ZN => 
                           n11920);
   U14353 : NAND4_X1 port map( A1 => n12459, A2 => n12460, A3 => n12382, A4 => 
                           n11916, ZN => n11917);
   U14354 : INV_X1 port map( A => n11918, ZN => n11919);
   U14355 : INV_X1 port map( A => n11922, ZN => n12574);
   U14356 : MUX2_X1 port map( A => n12577, B => n20462, S => n12574, Z => 
                           n11927);
   U14357 : NAND3_X1 port map( A1 => n20462, A2 => n12577, A3 => n11923, ZN => 
                           n11925);
   U14358 : XNOR2_X1 port map( A => n20155, B => n13453, ZN => n11928);
   U14359 : XNOR2_X1 port map( A => n11929, B => n11928, ZN => n11936);
   U14360 : INV_X1 port map( A => n11930, ZN => n12472);
   U14361 : NOR2_X1 port map( A1 => n12142, A2 => n12473, ZN => n11932);
   U14362 : XNOR2_X1 port map( A => n13058, B => n13528, ZN => n11934);
   U14363 : XNOR2_X1 port map( A => n13020, B => n2341, ZN => n11933);
   U14364 : XNOR2_X1 port map( A => n11934, B => n11933, ZN => n11935);
   U14366 : AOI22_X1 port map( A1 => n14627, A2 => n14146, B1 => n14192, B2 => 
                           n19875, ZN => n11989);
   U14367 : NOR2_X1 port map( A1 => n12110, A2 => n11942, ZN => n11937);
   U14368 : NAND2_X1 port map( A1 => n11939, A2 => n12441, ZN => n11940);
   U14369 : INV_X1 port map( A => n12093, ZN => n11945);
   U14370 : XNOR2_X1 port map( A => n13390, B => n12713, ZN => n11950);
   U14371 : NAND2_X1 port map( A1 => n20457, A2 => n12639, ZN => n12088);
   U14372 : INV_X1 port map( A => n12088, ZN => n11949);
   U14373 : OAI21_X1 port map( B1 => n11949, B2 => n11948, A => n11947, ZN => 
                           n13121);
   U14374 : INV_X1 port map( A => n13121, ZN => n13672);
   U14375 : XNOR2_X1 port map( A => n11950, B => n13672, ZN => n13436);
   U14376 : INV_X1 port map( A => n13436, ZN => n11968);
   U14377 : NOR2_X1 port map( A1 => n11952, A2 => n11951, ZN => n11959);
   U14378 : NAND2_X1 port map( A1 => n1578, A2 => n11953, ZN => n11958);
   U14380 : XNOR2_X1 port map( A => n13736, B => n2023, ZN => n11964);
   U14381 : OAI211_X1 port map( C1 => n11962, C2 => n12630, A => n11961, B => 
                           n11960, ZN => n11963);
   U14382 : XNOR2_X1 port map( A => n11964, B => n20222, ZN => n11966);
   U14383 : XNOR2_X1 port map( A => n11966, B => n11965, ZN => n11967);
   U14384 : XNOR2_X2 port map( A => n11968, B => n11967, ZN => n14623);
   U14385 : OR2_X1 port map( A1 => n12338, A2 => n3813, ZN => n11973);
   U14386 : XNOR2_X1 port map( A => n13534, B => n19887, ZN => n13416);
   U14387 : XNOR2_X1 port map( A => n13416, B => n11975, ZN => n11987);
   U14388 : NOR2_X1 port map( A1 => n250, A2 => n12305, ZN => n11976);
   U14389 : OAI21_X1 port map( B1 => n11977, B2 => n12305, A => n12547, ZN => 
                           n12307);
   U14390 : AOI21_X1 port map( B1 => n12589, B2 => n12200, A => n12202, ZN => 
                           n11981);
   U14392 : XNOR2_X1 port map( A => n13103, B => n13725, ZN => n11985);
   U14393 : AND2_X1 port map( A1 => n12616, A2 => n12615, ZN => n12246);
   U14394 : OAI21_X1 port map( B1 => n12246, B2 => n19784, A => n12240, ZN => 
                           n11982);
   U14395 : XNOR2_X1 port map( A => n20260, B => n2307, ZN => n11984);
   U14396 : XNOR2_X1 port map( A => n11985, B => n11984, ZN => n11986);
   U14397 : XNOR2_X1 port map( A => n11987, B => n11986, ZN => n14000);
   U14398 : OR2_X1 port map( A1 => n12339, A2 => n11990, ZN => n11991);
   U14399 : NAND3_X1 port map( A1 => n11991, A2 => n12338, A3 => n12332, ZN => 
                           n11994);
   U14400 : OAI21_X1 port map( B1 => n13275, B2 => n12326, A => n12322, ZN => 
                           n12000);
   U14401 : NAND2_X1 port map( A1 => n11996, A2 => n12326, ZN => n11999);
   U14404 : NAND2_X1 port map( A1 => n12352, A2 => n12349, ZN => n12175);
   U14405 : OR2_X1 port map( A1 => n12352, A2 => n12354, ZN => n12003);
   U14406 : XNOR2_X1 port map( A => n13736, B => n13795, ZN => n12913);
   U14407 : OR2_X1 port map( A1 => n12499, A2 => n12004, ZN => n12346);
   U14408 : AOI21_X1 port map( B1 => n12509, B2 => n12359, A => n12009, ZN => 
                           n12007);
   U14409 : AND2_X1 port map( A1 => n12359, A2 => n12009, ZN => n12364);
   U14410 : INV_X1 port map( A => n12508, ZN => n12010);
   U14411 : XNOR2_X1 port map( A => n13673, B => n2417, ZN => n12013);
   U14412 : XNOR2_X1 port map( A => n12014, B => n12013, ZN => n12015);
   U14413 : INV_X1 port map( A => n14203, ZN => n14206);
   U14414 : NAND2_X1 port map( A1 => n13145, A2 => n12254, ZN => n12017);
   U14416 : OAI21_X1 port map( B1 => n12020, B2 => n12369, A => n12381, ZN => 
                           n12026);
   U14417 : NAND2_X1 port map( A1 => n12373, A2 => n12369, ZN => n12023);
   U14418 : NAND3_X1 port map( A1 => n12376, A2 => n19504, A3 => n20191, ZN => 
                           n12022);
   U14419 : OAI21_X1 port map( B1 => n12381, B2 => n12023, A => n12022, ZN => 
                           n12024);
   U14420 : INV_X1 port map( A => n12024, ZN => n12025);
   U14421 : INV_X1 port map( A => n13369, ZN => n12027);
   U14422 : NOR2_X1 port map( A1 => n12028, A2 => n12274, ZN => n12031);
   U14423 : NOR2_X1 port map( A1 => n12272, A2 => n12029, ZN => n12030);
   U14424 : AND2_X1 port map( A1 => n12304, A2 => n12273, ZN => n12032);
   U14425 : NAND3_X1 port map( A1 => n12037, A2 => n12036, A3 => n12035, ZN => 
                           n12038);
   U14426 : OAI21_X1 port map( B1 => n12039, B2 => n12038, A => n12280, ZN => 
                           n12046);
   U14427 : OAI21_X1 port map( B1 => n12281, B2 => n876, A => n12040, ZN => 
                           n12045);
   U14428 : AOI21_X1 port map( B1 => n12280, B2 => n12042, A => n12041, ZN => 
                           n12043);
   U14429 : AOI22_X2 port map( A1 => n12046, A2 => n12045, B1 => n12044, B2 => 
                           n12043, ZN => n13783);
   U14430 : XNOR2_X1 port map( A => n13018, B => n13783, ZN => n12559);
   U14431 : NAND2_X1 port map( A1 => n12047, A2 => n12228, ZN => n12120);
   U14432 : NAND3_X1 port map( A1 => n12049, A2 => n12120, A3 => n12048, ZN => 
                           n12052);
   U14433 : NAND2_X1 port map( A1 => n12229, A2 => n1952, ZN => n12051);
   U14434 : NOR3_X1 port map( A1 => n1952, A2 => n12047, A3 => n12122, ZN => 
                           n12050);
   U14435 : INV_X1 port map( A => n12615, ZN => n12053);
   U14436 : NAND2_X1 port map( A1 => n12055, A2 => n12054, ZN => n12056);
   U14437 : NAND3_X1 port map( A1 => n12057, A2 => n2053, A3 => n19756, ZN => 
                           n12058);
   U14438 : XNOR2_X1 port map( A => n13658, B => n13260, ZN => n12920);
   U14439 : OAI21_X1 port map( B1 => n12592, B2 => n12593, A => n193, ZN => 
                           n12063);
   U14441 : NOR2_X1 port map( A1 => n12595, A2 => n20430, ZN => n12062);
   U14442 : INV_X1 port map( A => n13027, ZN => n12071);
   U14443 : INV_X1 port map( A => n12065, ZN => n12069);
   U14444 : NOR2_X1 port map( A1 => n2712, A2 => n19726, ZN => n12066);
   U14445 : AND2_X1 port map( A1 => n948, A2 => n12211, ZN => n12189);
   U14447 : INV_X1 port map( A => n13710, ZN => n12070);
   U14448 : XNOR2_X1 port map( A => n13206, B => n12920, ZN => n12081);
   U14449 : NOR2_X1 port map( A1 => n19971, A2 => n12237, ZN => n12075);
   U14450 : INV_X1 port map( A => n12601, ZN => n12608);
   U14451 : INV_X1 port map( A => n12077, ZN => n13772);
   U14452 : XNOR2_X1 port map( A => n13772, B => n17686, ZN => n12078);
   U14453 : XNOR2_X1 port map( A => n12079, B => n12078, ZN => n12080);
   U14454 : XNOR2_X1 port map( A => n12081, B => n12080, ZN => n13908);
   U14455 : INV_X1 port map( A => n13908, ZN => n12196);
   U14456 : MUX2_X1 port map( A => n14206, B => n14612, S => n12196, Z => 
                           n12199);
   U14457 : XNOR2_X1 port map( A => n12087, B => n12906, ZN => n13754);
   U14458 : NAND2_X1 port map( A1 => n12642, A2 => n20458, ZN => n12457);
   U14459 : NAND2_X1 port map( A1 => n12457, A2 => n12088, ZN => n12092);
   U14460 : NAND2_X1 port map( A1 => n12642, A2 => n19861, ZN => n12091);
   U14461 : AOI21_X1 port map( B1 => n2256, B2 => n12453, A => n20458, ZN => 
                           n12090);
   U14463 : AOI22_X1 port map( A1 => n12095, A2 => n12094, B1 => n12093, B2 => 
                           n12684, ZN => n12098);
   U14464 : NOR2_X1 port map( A1 => n12684, A2 => n12686, ZN => n12096);
   U14465 : NAND2_X1 port map( A1 => n12096, A2 => n12095, ZN => n12097);
   U14466 : XNOR2_X1 port map( A => n13065, B => n13462, ZN => n13218);
   U14467 : XNOR2_X1 port map( A => n13754, B => n13218, ZN => n12117);
   U14468 : XNOR2_X1 port map( A => n940, B => n13427, ZN => n12115);
   U14469 : INV_X1 port map( A => n12099, ZN => n12438);
   U14470 : INV_X1 port map( A => n12100, ZN => n12102);
   U14471 : NOR2_X1 port map( A1 => n12102, A2 => n12101, ZN => n12106);
   U14472 : MUX2_X1 port map( A => n12106, B => n12105, S => n12104, Z => 
                           n12108);
   U14473 : NOR2_X1 port map( A1 => n12108, A2 => n12107, ZN => n12109);
   U14474 : NAND3_X1 port map( A1 => n1099, A2 => n12440, A3 => n12110, ZN => 
                           n12111);
   U14475 : XNOR2_X1 port map( A => n13398, B => n17989, ZN => n12114);
   U14476 : XNOR2_X1 port map( A => n12115, B => n12114, ZN => n12116);
   U14477 : XNOR2_X1 port map( A => n12117, B => n12116, ZN => n14011);
   U14478 : INV_X1 port map( A => n13745, ZN => n12118);
   U14479 : XNOR2_X1 port map( A => n12119, B => n12118, ZN => n12135);
   U14480 : INV_X1 port map( A => n12120, ZN => n12125);
   U14481 : OAI21_X1 port map( B1 => n12122, B2 => n12228, A => n12121, ZN => 
                           n12124);
   U14483 : NOR2_X1 port map( A1 => n12129, A2 => n12128, ZN => n12131);
   U14484 : XNOR2_X1 port map( A => n12697, B => n13250, ZN => n12614);
   U14485 : XNOR2_X1 port map( A => n12135, B => n12614, ZN => n12161);
   U14486 : AOI21_X1 port map( B1 => n12382, B2 => n12463, A => n12138, ZN => 
                           n12136);
   U14487 : OAI21_X1 port map( B1 => n12470, B2 => n12382, A => n12136, ZN => 
                           n12140);
   U14488 : AND2_X1 port map( A1 => n857, A2 => n12137, ZN => n12466);
   U14489 : NOR2_X1 port map( A1 => n12137, A2 => n12386, ZN => n12467);
   U14490 : NAND2_X1 port map( A1 => n2550, A2 => n12479, ZN => n12145);
   U14491 : INV_X1 port map( A => n12142, ZN => n12474);
   U14492 : NAND2_X1 port map( A1 => n12478, A2 => n12474, ZN => n12143);
   U14493 : NAND3_X1 port map( A1 => n12480, A2 => n12393, A3 => n12143, ZN => 
                           n12144);
   U14496 : NOR2_X1 port map( A1 => n12148, A2 => n12147, ZN => n12151);
   U14498 : MUX2_X1 port map( A => n12154, B => n12153, S => n20486, Z => 
                           n12156);
   U14499 : NOR2_X1 port map( A1 => n12156, A2 => n12155, ZN => n12157);
   U14501 : XNOR2_X1 port map( A => n12159, B => n13643, ZN => n13187);
   U14502 : INV_X1 port map( A => n13187, ZN => n12160);
   U14504 : NAND2_X1 port map( A1 => n19488, A2 => n14011, ZN => n14614);
   U14505 : NAND2_X1 port map( A1 => n3811, A2 => n12537, ZN => n12164);
   U14506 : AND2_X1 port map( A1 => n12162, A2 => n12532, ZN => n12295);
   U14507 : OAI21_X1 port map( B1 => n12165, B2 => n12520, A => n907, ZN => 
                           n12166);
   U14508 : NOR2_X1 port map( A1 => n3256, A2 => n12166, ZN => n12171);
   U14509 : NAND2_X1 port map( A1 => n12168, A2 => n12167, ZN => n12289);
   U14510 : INV_X1 port map( A => n12289, ZN => n12169);
   U14511 : NAND2_X1 port map( A1 => n12169, A2 => n182, ZN => n12170);
   U14513 : XNOR2_X1 port map( A => n13721, B => n12173, ZN => n13191);
   U14514 : INV_X1 port map( A => n13191, ZN => n12186);
   U14515 : AND2_X1 port map( A1 => n11030, A2 => n19769, ZN => n12177);
   U14516 : INV_X1 port map( A => n12175, ZN => n12176);
   U14517 : AOI22_X1 port map( A1 => n12355, A2 => n12177, B1 => n12176, B2 => 
                           n11030, ZN => n12178);
   U14518 : AOI21_X1 port map( B1 => n12180, B2 => n256, A => n12179, ZN => 
                           n12184);
   U14519 : INV_X1 port map( A => n12745, ZN => n12889);
   U14520 : XNOR2_X1 port map( A => n13047, B => n12889, ZN => n12504);
   U14521 : XNOR2_X1 port map( A => n12186, B => n12504, ZN => n12195);
   U14522 : AOI21_X1 port map( B1 => n12188, B2 => n12187, A => n12212, ZN => 
                           n12190);
   U14523 : XNOR2_X1 port map( A => n13383, B => n13725, ZN => n12193);
   U14524 : XNOR2_X1 port map( A => n13339, B => n2384, ZN => n12192);
   U14525 : XNOR2_X1 port map( A => n12193, B => n12192, ZN => n12194);
   U14526 : XNOR2_X2 port map( A => n12195, B => n12194, ZN => n14611);
   U14527 : INV_X1 port map( A => n14611, ZN => n14208);
   U14528 : NAND3_X1 port map( A1 => n14614, A2 => n14208, A3 => n19488, ZN => 
                           n12198);
   U14529 : NAND3_X1 port map( A1 => n14612, A2 => n12196, A3 => n14611, ZN => 
                           n12197);
   U14531 : NOR2_X1 port map( A1 => n15474, A2 => n15769, ZN => n15245);
   U14532 : MUX2_X1 port map( A => n12200, B => n20430, S => n12595, Z => 
                           n12205);
   U14533 : NAND3_X1 port map( A1 => n12209, A2 => n2712, A3 => n12208, ZN => 
                           n12217);
   U14534 : NAND3_X1 port map( A1 => n12212, A2 => n12211, A3 => n12210, ZN => 
                           n12216);
   U14535 : NAND2_X1 port map( A1 => n12214, A2 => n12213, ZN => n12215);
   U14536 : XNOR2_X1 port map( A => n13295, B => n2087, ZN => n12219);
   U14537 : NAND2_X1 port map( A1 => n12225, A2 => n12224, ZN => n12231);
   U14538 : NAND2_X1 port map( A1 => n12231, A2 => n12047, ZN => n12236);
   U14539 : NAND3_X1 port map( A1 => n12230, A2 => n12229, A3 => n12228, ZN => 
                           n12234);
   U14540 : XNOR2_X1 port map( A => n13425, B => n19869, ZN => n13852);
   U14541 : MUX2_X1 port map( A => n12600, B => n12601, S => n12609, Z => 
                           n12238);
   U14542 : OAI21_X1 port map( B1 => n12616, B2 => n19784, A => n12242, ZN => 
                           n12618);
   U14543 : NAND2_X1 port map( A1 => n12241, A2 => n12243, ZN => n12245);
   U14544 : OAI211_X1 port map( C1 => n12618, C2 => n12246, A => n12245, B => 
                           n12244, ZN => n13688);
   U14545 : XNOR2_X1 port map( A => n13688, B => n13755, ZN => n12247);
   U14546 : XNOR2_X1 port map( A => n13397, B => n12247, ZN => n12248);
   U14547 : OAI21_X1 port map( B1 => n12251, B2 => n244, A => n12250, ZN => 
                           n12260);
   U14548 : AOI22_X1 port map( A1 => n12255, A2 => n12254, B1 => n12253, B2 => 
                           n12252, ZN => n12256);
   U14549 : OAI21_X1 port map( B1 => n13145, B2 => n12257, A => n12256, ZN => 
                           n12569);
   U14551 : OAI21_X1 port map( B1 => n12563, B2 => n12562, A => n12264, ZN => 
                           n12265);
   U14552 : NAND2_X1 port map( A1 => n12265, A2 => n248, ZN => n12266);
   U14553 : INV_X1 port map( A => n12373, ZN => n12370);
   U14554 : AOI21_X1 port map( B1 => n12374, B2 => n12269, A => n19504, ZN => 
                           n12270);
   U14555 : OAI22_X1 port map( A1 => n12271, A2 => n12370, B1 => n12381, B2 => 
                           n12270, ZN => n13724);
   U14556 : NAND2_X1 port map( A1 => n12272, A2 => n12304, ZN => n12302);
   U14557 : NAND2_X1 port map( A1 => n12274, A2 => n12273, ZN => n12303);
   U14558 : NAND2_X1 port map( A1 => n12302, A2 => n12303, ZN => n12276);
   U14559 : XNOR2_X1 port map( A => n19883, B => n13724, ZN => n12277);
   U14560 : XNOR2_X1 port map( A => n13303, B => n12277, ZN => n12287);
   U14561 : XNOR2_X1 port map( A => n13335, B => n12284, ZN => n13817);
   U14564 : INV_X1 port map( A => n12522, ZN => n12291);
   U14565 : OAI21_X1 port map( B1 => n12531, B2 => n20363, A => n12293, ZN => 
                           n12297);
   U14566 : NAND2_X1 port map( A1 => n924, A2 => n20363, ZN => n12296);
   U14567 : XNOR2_X1 port map( A => n19946, B => n13791, ZN => n12957);
   U14568 : OAI211_X1 port map( C1 => n12300, C2 => n12304, A => n12299, B => 
                           n12298, ZN => n12301);
   U14569 : OAI211_X1 port map( C1 => n12304, C2 => n12303, A => n12302, B => 
                           n12301, ZN => n13328);
   U14570 : NAND2_X1 port map( A1 => n250, A2 => n12305, ZN => n12309);
   U14571 : NAND2_X1 port map( A1 => n12307, A2 => n12306, ZN => n12308);
   U14572 : OAI21_X1 port map( B1 => n12310, B2 => n12309, A => n12308, ZN => 
                           n13735);
   U14573 : XNOR2_X1 port map( A => n13735, B => n13328, ZN => n13551);
   U14574 : XNOR2_X1 port map( A => n13551, B => n12957, ZN => n12319);
   U14575 : XNOR2_X1 port map( A => n13309, B => n13833, ZN => n12317);
   U14576 : XNOR2_X1 port map( A => n13391, B => n2203, ZN => n12316);
   U14577 : XNOR2_X1 port map( A => n12317, B => n12316, ZN => n12318);
   U14578 : INV_X1 port map( A => n13275, ZN => n12324);
   U14579 : NAND2_X1 port map( A1 => n13270, A2 => n13275, ZN => n12328);
   U14582 : XNOR2_X1 port map( A => n19796, B => n18396, ZN => n12331);
   U14583 : XNOR2_X1 port map( A => n13368, B => n13827, ZN => n12330);
   U14584 : XNOR2_X1 port map( A => n12330, B => n12331, ZN => n12368);
   U14585 : INV_X1 port map( A => n12334, ZN => n12336);
   U14586 : NAND2_X1 port map( A1 => n12340, A2 => n12339, ZN => n12341);
   U14588 : NOR2_X1 port map( A1 => n12354, A2 => n12349, ZN => n12351);
   U14590 : INV_X1 port map( A => n12506, ZN => n12361);
   U14591 : NAND2_X1 port map( A1 => n12508, A2 => n12359, ZN => n12360);
   U14592 : OAI22_X1 port map( A1 => n916, A2 => n12361, B1 => n12507, B2 => 
                           n12360, ZN => n12366);
   U14593 : NOR3_X1 port map( A1 => n12506, A2 => n12364, A3 => n3798, ZN => 
                           n12365);
   U14594 : XNOR2_X1 port map( A => n13826, B => n13781, ZN => n13527);
   U14595 : NAND2_X1 port map( A1 => n12370, A2 => n12369, ZN => n12380);
   U14596 : NAND2_X1 port map( A1 => n12371, A2 => n12373, ZN => n12379);
   U14597 : AND2_X1 port map( A1 => n12386, A2 => n12463, ZN => n12387);
   U14598 : INV_X1 port map( A => n12992, ZN => n13768);
   U14600 : AOI21_X1 port map( B1 => n12754, B2 => n12409, A => n12759, ZN => 
                           n12392);
   U14601 : NAND2_X1 port map( A1 => n12389, A2 => n12407, ZN => n12390);
   U14602 : XNOR2_X1 port map( A => n13544, B => n13657, ZN => n13846);
   U14603 : XNOR2_X1 port map( A => n13282, B => n13846, ZN => n12406);
   U14604 : NAND2_X1 port map( A1 => n12472, A2 => n12478, ZN => n12396);
   U14605 : NAND3_X1 port map( A1 => n12479, A2 => n12473, A3 => n19833, ZN => 
                           n12395);
   U14606 : XNOR2_X1 port map( A => n13601, B => n13259, ZN => n12404);
   U14607 : OAI21_X1 port map( B1 => n953, B2 => n12399, A => n12807, ZN => 
                           n12402);
   U14608 : NAND2_X1 port map( A1 => n12487, A2 => n12488, ZN => n12398);
   U14609 : AND2_X1 port map( A1 => n12398, A2 => n12397, ZN => n12401);
   U14610 : NOR2_X1 port map( A1 => n253, A2 => n12809, ZN => n12400);
   U14611 : AOI21_X1 port map( B1 => n12402, B2 => n12401, A => n12400, ZN => 
                           n13541);
   U14612 : INV_X1 port map( A => n13541, ZN => n13716);
   U14613 : XNOR2_X1 port map( A => n13716, B => n2263, ZN => n12403);
   U14614 : XNOR2_X1 port map( A => n12404, B => n12403, ZN => n12405);
   U14615 : XNOR2_X1 port map( A => n12406, B => n12405, ZN => n13891);
   U14616 : NOR2_X1 port map( A1 => n12412, A2 => n12759, ZN => n12413);
   U14617 : NOR2_X2 port map( A1 => n12414, A2 => n12413, ZN => n13251);
   U14618 : OAI21_X1 port map( B1 => n12417, B2 => n12416, A => n12415, ZN => 
                           n12426);
   U14619 : NAND2_X1 port map( A1 => n12418, A2 => n20351, ZN => n12420);
   U14620 : OR2_X1 port map( A1 => n12420, A2 => n12419, ZN => n12425);
   U14621 : NOR2_X1 port map( A1 => n12422, A2 => n20352, ZN => n12423);
   U14622 : NAND2_X1 port map( A1 => n257, A2 => n12423, ZN => n12424);
   U14623 : OAI211_X1 port map( C1 => n12427, C2 => n12426, A => n12425, B => 
                           n12424, ZN => n13168);
   U14624 : XNOR2_X1 port map( A => n12696, B => n13168, ZN => n13807);
   U14625 : NOR3_X1 port map( A1 => n12684, A2 => n12645, A3 => n12686, ZN => 
                           n12432);
   U14626 : AND3_X1 port map( A1 => n12684, A2 => n12430, A3 => n12429, ZN => 
                           n12431);
   U14627 : AOI21_X1 port map( B1 => n12434, B2 => n12685, A => n12433, ZN => 
                           n12448);
   U14628 : INV_X1 port map( A => n12435, ZN => n12436);
   U14629 : NAND2_X1 port map( A1 => n12440, A2 => n12439, ZN => n12445);
   U14630 : MUX2_X1 port map( A => n12445, B => n12444, S => n12443, Z => 
                           n12446);
   U14631 : NAND2_X1 port map( A1 => n12450, A2 => n12449, ZN => n12451);
   U14632 : NAND2_X1 port map( A1 => n19861, A2 => n12453, ZN => n12641);
   U14633 : MUX2_X1 port map( A => n20457, B => n12454, S => n12641, Z => 
                           n12456);
   U14634 : XNOR2_X1 port map( A => n12458, B => n19689, ZN => n13291);
   U14635 : NOR2_X1 port map( A1 => n14850, A2 => n14851, ZN => n15655);
   U14636 : INV_X1 port map( A => n15655, ZN => n15658);
   U14637 : INV_X1 port map( A => n12459, ZN => n12462);
   U14638 : NAND2_X1 port map( A1 => n12460, A2 => n991, ZN => n12461);
   U14639 : NOR2_X1 port map( A1 => n12462, A2 => n12461, ZN => n12464);
   U14640 : AOI22_X1 port map( A1 => n12465, A2 => n12464, B1 => n12463, B2 => 
                           n12137, ZN => n12469);
   U14641 : INV_X1 port map( A => n12471, ZN => n13343);
   U14642 : XNOR2_X1 port map( A => n12863, B => n13427, ZN => n13035);
   U14643 : XNOR2_X1 port map( A => n12864, B => n13035, ZN => n12496);
   U14644 : NOR2_X1 port map( A1 => n12480, A2 => n12472, ZN => n12476);
   U14645 : NOR2_X1 port map( A1 => n12474, A2 => n12473, ZN => n12475);
   U14647 : INV_X1 port map( A => n12478, ZN => n12483);
   U14648 : NAND2_X1 port map( A1 => n12480, A2 => n12479, ZN => n12482);
   U14649 : OAI22_X1 port map( A1 => n12484, A2 => n12483, B1 => n12482, B2 => 
                           n19833, ZN => n12485);
   U14650 : NOR2_X2 port map( A1 => n12486, A2 => n12485, ZN => n13512);
   U14651 : XNOR2_X1 port map( A => n13512, B => n12906, ZN => n12494);
   U14652 : NOR2_X1 port map( A1 => n953, A2 => n12487, ZN => n12491);
   U14653 : MUX2_X1 port map( A => n12811, B => n12488, S => n12809, Z => 
                           n12489);
   U14654 : XNOR2_X1 port map( A => n13396, B => n17999, ZN => n12493);
   U14655 : XNOR2_X1 port map( A => n12494, B => n12493, ZN => n12495);
   U14656 : INV_X1 port map( A => n14789, ZN => n14343);
   U14657 : OAI21_X1 port map( B1 => n12500, B2 => n12499, A => n12498, ZN => 
                           n12501);
   U14658 : XNOR2_X1 port map( A => n19887, B => n13468, ZN => n13340);
   U14659 : XNOR2_X1 port map( A => n13340, B => n12504, ZN => n12519);
   U14660 : OR2_X1 port map( A1 => n12509, A2 => n12508, ZN => n12511);
   U14661 : XNOR2_X1 port map( A => n13192, B => n18854, ZN => n12516);
   U14662 : XNOR2_X1 port map( A => n12517, B => n12516, ZN => n12518);
   U14663 : XNOR2_X1 port map( A => n12519, B => n12518, ZN => n14792);
   U14664 : NOR2_X1 port map( A1 => n12523, A2 => n12520, ZN => n12521);
   U14665 : NOR2_X1 port map( A1 => n12522, A2 => n12521, ZN => n12529);
   U14666 : NOR3_X1 port map( A1 => n12524, A2 => n907, A3 => n12523, ZN => 
                           n12527);
   U14667 : AOI211_X4 port map( C1 => n12529, C2 => n3256, A => n12527, B => 
                           n12526, ZN => n13173);
   U14668 : XNOR2_X1 port map( A => n13173, B => n13020, ZN => n12541);
   U14669 : INV_X1 port map( A => n12530, ZN => n12539);
   U14670 : OAI21_X1 port map( B1 => n12531, B2 => n12532, A => n12533, ZN => 
                           n12538);
   U14671 : NOR2_X1 port map( A1 => n12534, A2 => n12533, ZN => n12536);
   U14672 : XNOR2_X1 port map( A => n12541, B => n12540, ZN => n12561);
   U14673 : NAND2_X1 port map( A1 => n12543, A2 => n12542, ZN => n12546);
   U14674 : AOI21_X1 port map( B1 => n12547, B2 => n12546, A => n12555, ZN => 
                           n12558);
   U14675 : INV_X1 port map( A => n12548, ZN => n12550);
   U14676 : NAND2_X1 port map( A1 => n12550, A2 => n3615, ZN => n12551);
   U14677 : NOR3_X1 port map( A1 => n12553, A2 => n12552, A3 => n12551, ZN => 
                           n12556);
   U14678 : MUX2_X1 port map( A => n12556, B => n12555, S => n12554, Z => 
                           n12557);
   U14679 : INV_X1 port map( A => n13451, ZN => n13359);
   U14680 : XNOR2_X1 port map( A => n13017, B => n13359, ZN => n13366);
   U14681 : XNOR2_X1 port map( A => n12559, B => n13366, ZN => n12560);
   U14682 : INV_X1 port map( A => n14790, ZN => n13897);
   U14683 : NAND2_X1 port map( A1 => n12563, A2 => n12562, ZN => n12567);
   U14684 : OAI21_X1 port map( B1 => n12568, B2 => n12567, A => n12566, ZN => 
                           n13834);
   U14685 : XNOR2_X1 port map( A => n13834, B => n13390, ZN => n12870);
   U14687 : AND2_X1 port map( A1 => n20462, A2 => n12574, ZN => n12582);
   U14688 : NAND2_X1 port map( A1 => n12576, A2 => n12577, ZN => n12581);
   U14689 : NAND2_X1 port map( A1 => n12578, A2 => n12577, ZN => n12580);
   U14690 : AOI22_X1 port map( A1 => n12582, A2 => n12581, B1 => n12580, B2 => 
                           n12579, ZN => n12715);
   U14691 : INV_X1 port map( A => n12715, ZN => n13607);
   U14692 : XNOR2_X1 port map( A => n13479, B => n13607, ZN => n12583);
   U14693 : XNOR2_X1 port map( A => n12870, B => n12583, ZN => n12588);
   U14694 : XNOR2_X1 port map( A => n13795, B => n18819, ZN => n12586);
   U14695 : INV_X1 port map( A => n13031, ZN => n12584);
   U14696 : XNOR2_X1 port map( A => n12584, B => n13677, ZN => n12585);
   U14697 : XNOR2_X1 port map( A => n12586, B => n12585, ZN => n12587);
   U14699 : AOI22_X1 port map( A1 => n14343, A2 => n20141, B1 => n13897, B2 => 
                           n14787, ZN => n12657);
   U14700 : INV_X1 port map( A => n12596, ZN => n12599);
   U14701 : OAI21_X1 port map( B1 => n12592, B2 => n12591, A => n12590, ZN => 
                           n12598);
   U14702 : OAI21_X1 port map( B1 => n12599, B2 => n12598, A => n12597, ZN => 
                           n13376);
   U14703 : NAND2_X1 port map( A1 => n12601, A2 => n12600, ZN => n12605);
   U14704 : NAND2_X1 port map( A1 => n12607, A2 => n12606, ZN => n12612);
   U14705 : NAND3_X1 port map( A1 => n12610, A2 => n12609, A3 => n12608, ZN => 
                           n12611);
   U14706 : XNOR2_X1 port map( A => n13042, B => n13351, ZN => n12624);
   U14707 : MUX2_X1 port map( A => n12616, B => n12615, S => n19784, Z => 
                           n12622);
   U14708 : OR2_X1 port map( A1 => n12618, A2 => n19784, ZN => n12621);
   U14709 : XNOR2_X1 port map( A => n20253, B => n2368, ZN => n12623);
   U14710 : XNOR2_X1 port map( A => n12624, B => n12623, ZN => n12625);
   U14711 : NAND2_X1 port map( A1 => n12627, A2 => n14791, ZN => n14344);
   U14712 : INV_X1 port map( A => n14344, ZN => n12655);
   U14713 : NOR2_X1 port map( A1 => n3403, A2 => n20184, ZN => n12633);
   U14714 : XNOR2_X1 port map( A => n13405, B => n13659, ZN => n13437);
   U14715 : INV_X1 port map( A => n13437, ZN => n12652);
   U14718 : NAND2_X1 port map( A1 => n12645, A2 => n3649, ZN => n12651);
   U14719 : NOR2_X1 port map( A1 => n12648, A2 => n12647, ZN => n12649);
   U14720 : NAND2_X1 port map( A1 => n12684, A2 => n12649, ZN => n12650);
   U14721 : XNOR2_X1 port map( A => n20489, B => n13543, ZN => n13844);
   U14722 : XNOR2_X1 port map( A => n13844, B => n12652, ZN => n12653);
   U14723 : XNOR2_X1 port map( A => n12653, B => n12654, ZN => n14103);
   U14727 : INV_X1 port map( A => n14849, ZN => n15660);
   U14729 : NAND2_X1 port map( A1 => n15659, A2 => n15655, ZN => n12660);
   U14730 : NAND2_X1 port map( A1 => n12660, A2 => n15660, ZN => n12661);
   U14731 : XNOR2_X1 port map( A => n13397, B => n13512, ZN => n13097);
   U14732 : XNOR2_X1 port map( A => n13757, B => n13427, ZN => n12665);
   U14733 : XNOR2_X1 port map( A => n12665, B => n13097, ZN => n12668);
   U14734 : XNOR2_X1 port map( A => n13756, B => n13295, ZN => n13573);
   U14735 : XNOR2_X1 port map( A => n13063, B => n2448, ZN => n12666);
   U14736 : XNOR2_X1 port map( A => n13573, B => n12666, ZN => n12667);
   U14737 : XNOR2_X1 port map( A => n12668, B => n12667, ZN => n13940);
   U14738 : XNOR2_X1 port map( A => n13079, B => n13791, ZN => n12670);
   U14739 : XNOR2_X1 port map( A => n13677, B => n2401, ZN => n12669);
   U14740 : XNOR2_X1 port map( A => n12670, B => n12669, ZN => n12672);
   U14741 : XNOR2_X1 port map( A => n13479, B => n12671, ZN => n13550);
   U14742 : XNOR2_X1 port map( A => n13309, B => n13431, ZN => n13080);
   U14743 : XNOR2_X1 port map( A => n13468, B => n13622, ZN => n13536);
   U14744 : XNOR2_X1 port map( A => n13536, B => n19899, ZN => n12678);
   U14747 : XNOR2_X1 port map( A => n13088, B => n13618, ZN => n12675);
   U14748 : XNOR2_X1 port map( A => n12676, B => n12675, ZN => n12677);
   U14749 : MUX2_X1 port map( A => n2039, B => n19939, S => n14052, Z => n12695
                           );
   U14750 : INV_X1 port map( A => n19797, ZN => n12679);
   U14751 : XNOR2_X1 port map( A => n13058, B => n16242, ZN => n12680);
   U14752 : XNOR2_X1 port map( A => n13070, B => n13517, ZN => n13374);
   U14753 : INV_X1 port map( A => n13746, ZN => n12683);
   U14754 : XNOR2_X1 port map( A => n12683, B => n13518, ZN => n13353);
   U14755 : XNOR2_X1 port map( A => n13353, B => n13374, ZN => n12691);
   U14756 : XNOR2_X1 port map( A => n12697, B => n13584, ZN => n12689);
   U14757 : XNOR2_X1 port map( A => n13747, B => n610, ZN => n12688);
   U14758 : XNOR2_X1 port map( A => n12689, B => n12688, ZN => n12690);
   U14759 : XNOR2_X1 port map( A => n12691, B => n12690, ZN => n13939);
   U14760 : XNOR2_X1 port map( A => n13543, B => n13767, ZN => n13322);
   U14761 : XNOR2_X1 port map( A => n13282, B => n13322, ZN => n12694);
   U14762 : XNOR2_X1 port map( A => n13409, B => n13601, ZN => n13110);
   U14763 : XNOR2_X1 port map( A => n13659, B => n18084, ZN => n12692);
   U14764 : XNOR2_X1 port map( A => n13110, B => n12692, ZN => n12693);
   U14765 : XNOR2_X1 port map( A => n12694, B => n12693, ZN => n14355);
   U14766 : INV_X1 port map( A => n14355, ZN => n14418);
   U14767 : XNOR2_X1 port map( A => n12697, B => n12696, ZN => n13640);
   U14768 : XNOR2_X1 port map( A => n13352, B => n13585, ZN => n13812);
   U14769 : XNOR2_X1 port map( A => n13812, B => n13640, ZN => n12701);
   U14770 : XNOR2_X1 port map( A => n13590, B => n12846, ZN => n12699);
   U14771 : XNOR2_X1 port map( A => n19892, B => n16487, ZN => n12698);
   U14772 : XNOR2_X1 port map( A => n12699, B => n12698, ZN => n12700);
   U14773 : XNOR2_X1 port map( A => n12701, B => n12700, ZN => n14469);
   U14774 : INV_X1 port map( A => n14469, ZN => n14369);
   U14775 : XNOR2_X1 port map( A => n13085, B => n13047, ZN => n13633);
   U14776 : XNOR2_X1 port map( A => n13619, B => n13336, ZN => n13816);
   U14777 : XNOR2_X1 port map( A => n13816, B => n13633, ZN => n12706);
   U14778 : INV_X1 port map( A => n13534, ZN => n12702);
   U14779 : XNOR2_X1 port map( A => n12702, B => n13624, ZN => n12704);
   U14780 : XNOR2_X1 port map( A => n13193, B => n2356, ZN => n12703);
   U14781 : XNOR2_X1 port map( A => n12704, B => n12703, ZN => n12705);
   U14782 : NOR2_X1 port map( A1 => n14369, A2 => n14468, ZN => n12727);
   U14783 : XNOR2_X1 port map( A => n13017, B => n2306, ZN => n12707);
   U14784 : XNOR2_X1 port map( A => n12707, B => n19792, ZN => n12708);
   U14785 : XNOR2_X1 port map( A => n12708, B => n13357, ZN => n12712);
   U14786 : XNOR2_X1 port map( A => n13528, B => n12709, ZN => n13057);
   U14791 : XNOR2_X1 port map( A => n12986, B => n632, ZN => n12714);
   U14792 : XNOR2_X1 port map( A => n13120, B => n12715, ZN => n13838);
   U14793 : XNOR2_X1 port map( A => n13404, B => n13321, ZN => n13542);
   U14794 : XNOR2_X1 port map( A => n13842, B => n13542, ZN => n12719);
   U14795 : XNOR2_X1 port map( A => n13657, B => n13659, ZN => n12717);
   U14796 : XNOR2_X1 port map( A => n19697, B => n311, ZN => n12716);
   U14797 : XNOR2_X1 port map( A => n12717, B => n12716, ZN => n12718);
   U14798 : XNOR2_X1 port map( A => n12719, B => n12718, ZN => n14462);
   U14799 : INV_X1 port map( A => n14468, ZN => n12725);
   U14800 : XNOR2_X1 port map( A => n13344, B => n13064, ZN => n13510);
   U14801 : XNOR2_X1 port map( A => n13396, B => n13099, ZN => n13853);
   U14802 : INV_X1 port map( A => n13853, ZN => n12720);
   U14803 : XNOR2_X1 port map( A => n12720, B => n13510, ZN => n12724);
   U14804 : XNOR2_X1 port map( A => n13427, B => n12979, ZN => n12722);
   U14805 : XNOR2_X1 port map( A => n13425, B => n19018, ZN => n12721);
   U14806 : XNOR2_X1 port map( A => n12722, B => n12721, ZN => n12723);
   U14807 : XNOR2_X1 port map( A => n12724, B => n12723, ZN => n13921);
   U14808 : XNOR2_X1 port map( A => n13484, B => n13795, ZN => n12729);
   U14809 : XNOR2_X1 port map( A => n12729, B => n12728, ZN => n12733);
   U14810 : XNOR2_X1 port map( A => n12986, B => n20222, ZN => n12731);
   U14811 : XNOR2_X1 port map( A => n13673, B => n13121, ZN => n12915);
   U14812 : INV_X1 port map( A => n12915, ZN => n12730);
   U14813 : XNOR2_X1 port map( A => n12730, B => n12731, ZN => n12732);
   U14814 : XNOR2_X1 port map( A => n12732, B => n12733, ZN => n14826);
   U14815 : INV_X1 port map( A => n13440, ZN => n12734);
   U14816 : XNOR2_X1 port map( A => n12734, B => n12920, ZN => n12739);
   U14817 : INV_X1 port map( A => n19697, ZN => n12735);
   U14818 : INV_X1 port map( A => n13843, ZN => n13258);
   U14819 : XNOR2_X1 port map( A => n13258, B => n12735, ZN => n12737);
   U14820 : XNOR2_X1 port map( A => n13602, B => Key(63), ZN => n12736);
   U14821 : XNOR2_X1 port map( A => n12737, B => n12736, ZN => n12738);
   U14822 : XNOR2_X1 port map( A => n13572, B => n12979, ZN => n12741);
   U14825 : XNOR2_X1 port map( A => n20237, B => n12741, ZN => n12744);
   U14827 : XNOR2_X1 port map( A => n13064, B => n19140, ZN => n12742);
   U14828 : XNOR2_X1 port map( A => n13649, B => n12742, ZN => n12743);
   U14829 : INV_X1 port map( A => n12996, ZN => n12746);
   U14830 : XNOR2_X1 port map( A => n13631, B => n12746, ZN => n12750);
   U14831 : XNOR2_X1 port map( A => n20482, B => n13623, ZN => n12748);
   U14832 : XNOR2_X1 port map( A => n13193, B => n19457, ZN => n12747);
   U14833 : XNOR2_X1 port map( A => n12748, B => n12747, ZN => n12749);
   U14834 : NOR2_X1 port map( A1 => n14347, A2 => n2684, ZN => n14833);
   U14835 : XNOR2_X1 port map( A => n13491, B => n13643, ZN => n12961);
   U14836 : XNOR2_X1 port map( A => n13641, B => n12961, ZN => n12753);
   U14837 : XNOR2_X1 port map( A => n12846, B => n13250, ZN => n13012);
   U14838 : XNOR2_X1 port map( A => n19892, B => n18006, ZN => n12751);
   U14839 : XNOR2_X1 port map( A => n13012, B => n12751, ZN => n12752);
   U14840 : XNOR2_X1 port map( A => n13453, B => n13369, ZN => n13668);
   U14841 : XNOR2_X1 port map( A => n13002, B => n13277, ZN => n12760);
   U14842 : XNOR2_X1 port map( A => n933, B => n12760, ZN => n12764);
   U14843 : XNOR2_X1 port map( A => n13230, B => n13528, ZN => n12762);
   U14844 : XNOR2_X1 port map( A => n13783, B => n18809, ZN => n12761);
   U14845 : XNOR2_X1 port map( A => n12762, B => n12761, ZN => n12763);
   U14846 : OAI21_X1 port map( B1 => n14827, B2 => n14826, A => n19985, ZN => 
                           n12765);
   U14847 : NAND2_X1 port map( A1 => n19496, A2 => n12765, ZN => n12766);
   U14848 : MUX2_X1 port map( A => n15341, B => n12768, S => n12842, Z => 
                           n12875);
   U14849 : XNOR2_X1 port map( A => n13248, B => n12769, ZN => n13744);
   U14850 : XNOR2_X1 port map( A => n13168, B => n2423, ZN => n12771);
   U14851 : XNOR2_X1 port map( A => n13490, B => n12771, ZN => n12773);
   U14852 : XNOR2_X1 port map( A => n13070, B => n20123, ZN => n12772);
   U14853 : XNOR2_X1 port map( A => n12773, B => n12772, ZN => n12774);
   U14854 : XNOR2_X1 port map( A => n12774, B => n13744, ZN => n12876);
   U14855 : INV_X1 port map( A => n12876, ZN => n14094);
   U14856 : XNOR2_X1 port map( A => n13617, B => n13088, ZN => n12775);
   U14857 : XNOR2_X1 port map( A => n13761, B => n12775, ZN => n12779);
   U14858 : XNOR2_X1 port map( A => n13335, B => n13048, ZN => n12777);
   U14859 : XNOR2_X1 port map( A => n13339, B => n19321, ZN => n12776);
   U14860 : XOR2_X1 port map( A => n12777, B => n12776, Z => n12778);
   U14862 : XNOR2_X1 port map( A => n13293, B => n13687, ZN => n12905);
   U14863 : INV_X1 port map( A => n12905, ZN => n12780);
   U14864 : XNOR2_X1 port map( A => n13134, B => n19869, ZN => n13348);
   U14865 : XNOR2_X1 port map( A => n12780, B => n13348, ZN => n12783);
   U14866 : XNOR2_X1 port map( A => n12940, B => n13688, ZN => n13753);
   U14867 : XNOR2_X1 port map( A => n13063, B => n1386, ZN => n12781);
   U14868 : XNOR2_X1 port map( A => n13753, B => n12781, ZN => n12782);
   U14869 : NAND2_X1 port map( A1 => n19485, A2 => n13931, ZN => n14093);
   U14870 : XNOR2_X1 port map( A => n13312, B => n13079, ZN => n12787);
   U14871 : XNOR2_X1 port map( A => n12787, B => n12786, ZN => n12790);
   U14872 : INV_X1 port map( A => n13551, ZN => n12788);
   U14873 : XNOR2_X1 port map( A => n12788, B => n13237, ZN => n12789);
   U14874 : XNOR2_X1 port map( A => n13233, B => n13527, ZN => n12794);
   U14875 : XNOR2_X1 port map( A => n13776, B => n17804, ZN => n12792);
   U14876 : XNOR2_X1 port map( A => n12791, B => n12792, ZN => n12793);
   U14877 : XNOR2_X1 port map( A => n12794, B => n12793, ZN => n13930);
   U14879 : INV_X1 port map( A => n13930, ZN => n14336);
   U14880 : XNOR2_X1 port map( A => n13255, B => n13280, ZN => n12921);
   U14881 : XNOR2_X1 port map( A => n13772, B => n13544, ZN => n13325);
   U14882 : XNOR2_X1 port map( A => n13325, B => n12921, ZN => n12799);
   U14883 : INV_X1 port map( A => n13409, ZN => n12795);
   U14884 : XNOR2_X1 port map( A => n12795, B => n13539, ZN => n12797);
   U14885 : XNOR2_X1 port map( A => n13716, B => n17733, ZN => n12796);
   U14886 : XNOR2_X1 port map( A => n12797, B => n12796, ZN => n12798);
   U14887 : XNOR2_X1 port map( A => n12798, B => n12799, ZN => n12879);
   U14888 : INV_X1 port map( A => n12879, ZN => n14092);
   U14889 : NAND2_X1 port map( A1 => n14334, A2 => n14342, ZN => n12801);
   U14891 : XNOR2_X1 port map( A => n13511, B => n18011, ZN => n12803);
   U14892 : XNOR2_X1 port map( A => n12803, B => n13572, ZN => n12804);
   U14893 : XNOR2_X1 port map( A => n13755, B => n940, ZN => n12938);
   U14894 : XNOR2_X1 port map( A => n12938, B => n12804, ZN => n12806);
   U14895 : XNOR2_X1 port map( A => n13651, B => n13218, ZN => n12805);
   U14896 : NAND2_X1 port map( A1 => n12807, A2 => n12809, ZN => n12808);
   U14897 : OAI211_X1 port map( C1 => n3586, C2 => n12809, A => n12811, B => 
                           n12808, ZN => n12810);
   U14898 : INV_X1 port map( A => n12810, ZN => n12815);
   U14899 : AOI21_X1 port map( B1 => n953, B2 => n12812, A => n12811, ZN => 
                           n12814);
   U14900 : XNOR2_X1 port map( A => n13251, B => n13287, ZN => n12965);
   U14901 : INV_X1 port map( A => n12965, ZN => n12817);
   U14902 : INV_X1 port map( A => n13446, ZN => n12816);
   U14903 : XNOR2_X1 port map( A => n12816, B => n13642, ZN => n13489);
   U14904 : INV_X1 port map( A => n13489, ZN => n13694);
   U14905 : XNOR2_X1 port map( A => n12817, B => n13694, ZN => n12822);
   U14906 : INV_X1 port map( A => n13168, ZN => n12818);
   U14907 : XNOR2_X1 port map( A => n13491, B => n12818, ZN => n12820);
   U14908 : XNOR2_X1 port map( A => n13644, B => n2082, ZN => n12819);
   U14909 : XNOR2_X1 port map( A => n12820, B => n12819, ZN => n12821);
   U14910 : XNOR2_X1 port map( A => n12822, B => n12821, ZN => n14087);
   U14911 : INV_X1 port map( A => n14087, ZN => n14821);
   U14912 : XNOR2_X1 port map( A => n19883, B => n13725, ZN => n12823);
   U14913 : XNOR2_X1 port map( A => n13335, B => n2454, ZN => n12825);
   U14914 : INV_X1 port map( A => n13138, ZN => n13635);
   U14915 : XNOR2_X1 port map( A => n13635, B => n13623, ZN => n12824);
   U14916 : NOR2_X1 port map( A1 => n14821, A2 => n14818, ZN => n14328);
   U14917 : XNOR2_X1 port map( A => n13778, B => n13702, ZN => n12950);
   U14918 : XNOR2_X1 port map( A => n12826, B => n12950, ZN => n12830);
   U14919 : XNOR2_X1 port map( A => n20440, B => n13706, ZN => n12828);
   U14920 : XNOR2_X1 port map( A => n13277, B => n106, ZN => n12827);
   U14921 : XNOR2_X1 port map( A => n12828, B => n12827, ZN => n12829);
   U14922 : XNOR2_X1 port map( A => n12831, B => n19102, ZN => n12832);
   U14923 : XNOR2_X1 port map( A => n12832, B => n13717, ZN => n12833);
   U14924 : XNOR2_X1 port map( A => n13206, B => n12833, ZN => n12835);
   U14925 : XNOR2_X1 port map( A => n12834, B => n13711, ZN => n12971);
   U14926 : XNOR2_X1 port map( A => n12835, B => n12971, ZN => n14325);
   U14927 : NOR2_X1 port map( A1 => n14823, A2 => n14352, ZN => n14330);
   U14928 : AOI21_X1 port map( B1 => n19693, B2 => n14328, A => n14330, ZN => 
                           n12841);
   U14929 : INV_X1 port map( A => n14325, ZN => n12932);
   U14931 : XNOR2_X1 port map( A => n12914, B => n13734, ZN => n13238);
   U14932 : XNOR2_X1 port map( A => n13199, B => n13238, ZN => n12838);
   U14933 : XNOR2_X1 port map( A => n13736, B => n13484, ZN => n13311);
   U14934 : XNOR2_X1 port map( A => n13328, B => n18768, ZN => n12836);
   U14935 : XNOR2_X1 port map( A => n13311, B => n12836, ZN => n12837);
   U14936 : XNOR2_X1 port map( A => n12838, B => n12837, ZN => n12931);
   U14937 : INV_X1 port map( A => n12931, ZN => n14326);
   U14938 : NOR2_X1 port map( A1 => n14352, A2 => n912, ZN => n14817);
   U14939 : INV_X1 port map( A => n14817, ZN => n12839);
   U14940 : OAI211_X1 port map( C1 => n12932, C2 => n14326, A => n14350, B => 
                           n12839, ZN => n12840);
   U14941 : INV_X1 port map( A => n12842, ZN => n15468);
   U14942 : INV_X1 port map( A => n13351, ZN => n12843);
   U14943 : XNOR2_X1 port map( A => n13251, B => n12843, ZN => n12845);
   U14944 : XNOR2_X1 port map( A => n13810, B => n18984, ZN => n12844);
   U14945 : XNOR2_X1 port map( A => n12845, B => n12844, ZN => n12848);
   U14946 : XNOR2_X1 port map( A => n13644, B => n13376, ZN => n13073);
   U14947 : XNOR2_X1 port map( A => n13042, B => n12846, ZN => n13693);
   U14948 : XNOR2_X1 port map( A => n13073, B => n13693, ZN => n12847);
   U14949 : INV_X1 port map( A => n14453, ZN => n14179);
   U14950 : XNOR2_X1 port map( A => n20260, B => n13136, ZN => n13815);
   U14951 : XNOR2_X1 port map( A => n13193, B => n13192, ZN => n13722);
   U14952 : XNOR2_X1 port map( A => n13815, B => n13722, ZN => n12853);
   U14953 : INV_X1 port map( A => n12997, ZN => n12849);
   U14954 : XNOR2_X1 port map( A => n12945, B => n12849, ZN => n12851);
   U14955 : XNOR2_X1 port map( A => n12851, B => n12850, ZN => n12852);
   U14956 : INV_X1 port map( A => n13715, ZN => n12854);
   U14957 : XNOR2_X1 port map( A => n19697, B => n12854, ZN => n12856);
   U14958 : XNOR2_X1 port map( A => n13259, B => n2446, ZN => n12855);
   U14959 : XNOR2_X1 port map( A => n12856, B => n12855, ZN => n12857);
   U14961 : AOI21_X1 port map( B1 => n14179, B2 => n1364, A => n14451, ZN => 
                           n12873);
   U14962 : XNOR2_X1 port map( A => n13173, B => n13230, ZN => n13823);
   U14963 : XNOR2_X1 port map( A => n12859, B => n19216, ZN => n12860);
   U14964 : XNOR2_X1 port map( A => n13823, B => n12860, ZN => n12862);
   U14965 : XNOR2_X1 port map( A => n12863, B => n12979, ZN => n13684);
   U14966 : XNOR2_X1 port map( A => n12864, B => n13684, ZN => n12867);
   U14967 : XNOR2_X1 port map( A => n13065, B => n13848, ZN => n13650);
   U14968 : XNOR2_X1 port map( A => n13755, B => n18078, ZN => n12865);
   U14969 : XNOR2_X1 port map( A => n13650, B => n12865, ZN => n12866);
   U14970 : INV_X1 port map( A => n14450, ZN => n14454);
   U14971 : XNOR2_X1 port map( A => n12914, B => n20682, ZN => n12868);
   U14972 : XNOR2_X1 port map( A => n13733, B => n12868, ZN => n12872);
   U14973 : INV_X1 port map( A => n13081, ZN => n12869);
   U14974 : XNOR2_X1 port map( A => n12869, B => n20223, ZN => n13676);
   U14975 : XNOR2_X1 port map( A => n13676, B => n12870, ZN => n12871);
   U14976 : INV_X1 port map( A => n15339, ZN => n14896);
   U14977 : NAND2_X1 port map( A1 => n14092, A2 => n14336, ZN => n12877);
   U14978 : NAND2_X1 port map( A1 => n12880, A2 => n13931, ZN => n12881);
   U14979 : INV_X1 port map( A => n14052, ZN => n14357);
   U14980 : MUX2_X1 port map( A => n14357, B => n14419, S => n19939, Z => 
                           n12884);
   U14981 : NAND3_X1 port map( A1 => n14357, A2 => n14355, A3 => n14419, ZN => 
                           n12883);
   U14982 : NAND3_X1 port map( A1 => n2039, A2 => n14359, A3 => n14422, ZN => 
                           n12882);
   U14985 : MUX2_X1 port map( A => n14369, B => n19531, S => n3252, Z => n12887
                           );
   U14986 : MUX2_X1 port map( A => n14465, B => n19819, S => n19657, Z => 
                           n12886);
   U14987 : INV_X1 port map( A => n12888, ZN => n15165);
   U14988 : XNOR2_X1 port map( A => n12889, B => n12945, ZN => n13764);
   U14989 : XNOR2_X1 port map( A => n13764, B => n13631, ZN => n12893);
   U14990 : XNOR2_X1 port map( A => n13617, B => n13725, ZN => n12891);
   U14991 : XNOR2_X1 port map( A => n13048, B => n1904, ZN => n12890);
   U14992 : XNOR2_X1 port map( A => n12891, B => n12890, ZN => n12892);
   U14993 : XNOR2_X1 port map( A => n12893, B => n12892, ZN => n12910);
   U14994 : INV_X1 port map( A => n12910, ZN => n14441);
   U14995 : XNOR2_X1 port map( A => n20123, B => n13643, ZN => n12895);
   U14996 : XNOR2_X1 port map( A => n12895, B => n12894, ZN => n12899);
   U14997 : XNOR2_X1 port map( A => n13250, B => n2413, ZN => n12897);
   U14998 : INV_X1 port map( A => n13251, ZN => n12896);
   U14999 : XNOR2_X1 port map( A => n12898, B => n12899, ZN => n12911);
   U15000 : XNOR2_X1 port map( A => n13019, B => n13580, ZN => n12901);
   U15001 : XNOR2_X1 port map( A => n13783, B => n2122, ZN => n12900);
   U15002 : XNOR2_X1 port map( A => n12901, B => n12900, ZN => n12904);
   U15003 : INV_X1 port map( A => n12950, ZN => n12902);
   U15004 : XNOR2_X1 port map( A => n13668, B => n12902, ZN => n12903);
   U15005 : XNOR2_X1 port map( A => n12905, B => n12938, ZN => n12909);
   U15006 : XNOR2_X1 port map( A => n12906, B => n18863, ZN => n12907);
   U15007 : XNOR2_X1 port map( A => n13649, B => n12907, ZN => n12908);
   U15008 : XNOR2_X1 port map( A => n13312, B => n19734, ZN => n12912);
   U15009 : XNOR2_X1 port map( A => n12912, B => n12913, ZN => n12918);
   U15010 : XNOR2_X1 port map( A => n12914, B => n2424, ZN => n12916);
   U15011 : XNOR2_X1 port map( A => n12915, B => n12916, ZN => n12917);
   U15012 : XNOR2_X1 port map( A => n12918, B => n12917, ZN => n14167);
   U15013 : INV_X1 port map( A => n14167, ZN => n12919);
   U15014 : XNOR2_X1 port map( A => n12921, B => n12920, ZN => n12925);
   U15016 : XNOR2_X1 port map( A => n13259, B => n2192, ZN => n12922);
   U15017 : XNOR2_X1 port map( A => n12923, B => n12922, ZN => n12924);
   U15018 : XNOR2_X1 port map( A => n12925, B => n12924, ZN => n13918);
   U15019 : AOI22_X1 port map( A1 => n14439, A2 => n12926, B1 => n3516, B2 => 
                           n20262, ZN => n12927);
   U15020 : NAND2_X1 port map( A1 => n15165, A2 => n15379, ZN => n15375);
   U15021 : MUX2_X1 port map( A => n13559, B => n1363, S => n14455, Z => n12930
                           );
   U15023 : NAND2_X1 port map( A1 => n231, A2 => n19513, ZN => n15031);
   U15024 : NAND2_X1 port map( A1 => n15375, A2 => n15031, ZN => n12935);
   U15025 : AOI21_X1 port map( B1 => n235, B2 => n12931, A => n14352, ZN => 
                           n12934);
   U15026 : AND2_X1 port map( A1 => n12932, A2 => n12931, ZN => n14085);
   U15027 : OAI21_X1 port map( B1 => n14086, B2 => n14085, A => n19821, ZN => 
                           n12933);
   U15029 : XNOR2_X1 port map( A => n12937, B => n13572, ZN => n12939);
   U15030 : XNOR2_X1 port map( A => n12938, B => n12939, ZN => n12943);
   U15031 : XNOR2_X1 port map( A => n13398, B => n12940, ZN => n13215);
   U15032 : XNOR2_X1 port map( A => n13757, B => n18146, ZN => n12941);
   U15033 : XNOR2_X1 port map( A => n13215, B => n12941, ZN => n12942);
   U15034 : XNOR2_X1 port map( A => n13222, B => n13762, ZN => n12944);
   U15035 : XNOR2_X1 port map( A => n13725, B => n13623, ZN => n13302);
   U15036 : XNOR2_X1 port map( A => n13302, B => n12944, ZN => n12949);
   U15037 : XNOR2_X1 port map( A => n13624, B => n19923, ZN => n12947);
   U15038 : XNOR2_X1 port map( A => n19883, B => n18065, ZN => n12946);
   U15039 : XNOR2_X1 port map( A => n12947, B => n12946, ZN => n12948);
   U15040 : XNOR2_X1 port map( A => n12949, B => n12948, ZN => n12973);
   U15041 : INV_X1 port map( A => n12973, ZN => n14509);
   U15042 : NOR2_X1 port map( A1 => n20473, A2 => n14509, ZN => n14636);
   U15043 : XNOR2_X1 port map( A => n13577, B => n13774, ZN => n13525);
   U15044 : XNOR2_X1 port map( A => n12950, B => n13525, ZN => n12954);
   U15045 : XNOR2_X1 port map( A => n13369, B => n13277, ZN => n12952);
   U15046 : XNOR2_X1 port map( A => n19796, B => n2280, ZN => n12951);
   U15047 : XNOR2_X1 port map( A => n12952, B => n12951, ZN => n12953);
   U15049 : XNOR2_X1 port map( A => n13792, B => n12955, ZN => n12956);
   U15050 : XNOR2_X1 port map( A => n12956, B => n12957, ZN => n12960);
   U15051 : XNOR2_X1 port map( A => n13673, B => Key(94), ZN => n12958);
   U15052 : XNOR2_X1 port map( A => n13311, B => n12958, ZN => n12959);
   U15053 : XNOR2_X1 port map( A => n12960, B => n12959, ZN => n14642);
   U15054 : NOR2_X1 port map( A1 => n14642, A2 => n14641, ZN => n14031);
   U15055 : AOI22_X1 port map( A1 => n14636, A2 => n19703, B1 => n14031, B2 => 
                           n14509, ZN => n12976);
   U15056 : XNOR2_X1 port map( A => n12961, B => n13248, ZN => n12968);
   U15057 : XNOR2_X1 port map( A => n12964, B => n13747, ZN => n12966);
   U15058 : XNOR2_X1 port map( A => n12965, B => n12966, ZN => n12967);
   U15060 : XNOR2_X1 port map( A => n12992, B => n19222, ZN => n12969);
   U15061 : XNOR2_X1 port map( A => n12969, B => n13321, ZN => n12970);
   U15062 : XNOR2_X1 port map( A => n13658, B => n13539, ZN => n13207);
   U15064 : XNOR2_X1 port map( A => n12977, B => n13687, ZN => n12978);
   U15065 : XNOR2_X1 port map( A => n20442, B => n12978, ZN => n12983);
   U15066 : XNOR2_X1 port map( A => n12471, B => n2123, ZN => n12981);
   U15067 : XNOR2_X1 port map( A => n12979, B => n13462, ZN => n12980);
   U15068 : XNOR2_X1 port map( A => n12981, B => n12980, ZN => n12982);
   U15070 : XNOR2_X1 port map( A => n13791, B => n20223, ZN => n12985);
   U15071 : XNOR2_X1 port map( A => n13029, B => n12984, ZN => n13732);
   U15072 : XNOR2_X1 port map( A => n12985, B => n13732, ZN => n12990);
   U15073 : XNOR2_X1 port map( A => n13795, B => n12986, ZN => n12988);
   U15074 : XNOR2_X1 port map( A => n13390, B => n347, ZN => n12987);
   U15075 : XNOR2_X1 port map( A => n12987, B => n12988, ZN => n12989);
   U15076 : XNOR2_X1 port map( A => n12990, B => n12989, ZN => n14525);
   U15077 : NOR2_X1 port map( A1 => n20443, A2 => n19831, ZN => n13008);
   U15078 : XNOR2_X1 port map( A => n13260, B => n17024, ZN => n12991);
   U15079 : XNOR2_X1 port map( A => n13714, B => n12991, ZN => n12995);
   U15080 : XNOR2_X1 port map( A => n13710, B => n12992, ZN => n13497);
   U15081 : XNOR2_X1 port map( A => n12993, B => n13497, ZN => n12994);
   U15082 : XNOR2_X1 port map( A => n13721, B => n13762, ZN => n13470);
   U15083 : XNOR2_X1 port map( A => n13470, B => n12996, ZN => n13001);
   U15084 : XNOR2_X1 port map( A => n12999, B => n12998, ZN => n13000);
   U15086 : XNOR2_X1 port map( A => n13783, B => n642, ZN => n13004);
   U15087 : XNOR2_X1 port map( A => n13005, B => n13004, ZN => n13006);
   U15089 : XNOR2_X1 port map( A => n13695, B => n13810, ZN => n13011);
   U15090 : XNOR2_X1 port map( A => n13747, B => n17466, ZN => n13010);
   U15091 : XNOR2_X1 port map( A => n13011, B => n13010, ZN => n13015);
   U15092 : XNOR2_X1 port map( A => n13446, B => n13351, ZN => n13013);
   U15093 : XOR2_X1 port map( A => n13013, B => n13012, Z => n13014);
   U15094 : NAND3_X1 port map( A1 => n14522, A2 => n14524, A3 => n20443, ZN => 
                           n13016);
   U15095 : INV_X1 port map( A => n15684, ZN => n15687);
   U15096 : NOR2_X1 port map( A1 => n19978, A2 => n15687, ZN => n13096);
   U15097 : INV_X1 port map( A => n19978, ZN => n15779);
   U15098 : XNOR2_X1 port map( A => n13576, B => n13114, ZN => n13829);
   U15099 : XNOR2_X1 port map( A => n20199, B => n13018, ZN => n13666);
   U15100 : XNOR2_X1 port map( A => n13666, B => n13829, ZN => n13024);
   U15101 : XNOR2_X1 port map( A => n13019, B => n13453, ZN => n13022);
   U15102 : XNOR2_X1 port map( A => n13020, B => n2369, ZN => n13021);
   U15103 : XNOR2_X1 port map( A => n13022, B => n13021, ZN => n13023);
   U15105 : XNOR2_X1 port map( A => n13255, B => n13659, ZN => n13026);
   U15106 : XNOR2_X1 port map( A => n13715, B => n2395, ZN => n13025);
   U15107 : XNOR2_X1 port map( A => n13027, B => n13108, ZN => n13655);
   U15108 : XNOR2_X1 port map( A => n13842, B => n13655, ZN => n13028);
   U15109 : XNOR2_X1 port map( A => n19734, B => n13677, ZN => n13030);
   U15110 : XNOR2_X1 port map( A => n13030, B => n13838, ZN => n13034);
   U15111 : XNOR2_X1 port map( A => n13031, B => n13081, ZN => n13033);
   U15112 : XNOR2_X1 port map( A => n13121, B => n1869, ZN => n13032);
   U15113 : XNOR2_X1 port map( A => n19937, B => n13687, ZN => n13036);
   U15114 : XNOR2_X1 port map( A => n13036, B => n13035, ZN => n13039);
   U15115 : XNOR2_X1 port map( A => n13422, B => n2317, ZN => n13037);
   U15116 : XNOR2_X1 port map( A => n13853, B => n13037, ZN => n13038);
   U15117 : XNOR2_X2 port map( A => n13039, B => n13038, ZN => n14499);
   U15118 : INV_X1 port map( A => n14499, ZN => n13040);
   U15119 : XNOR2_X1 port map( A => n13041, B => n13126, ZN => n13443);
   U15120 : XNOR2_X1 port map( A => n13443, B => n13812, ZN => n13046);
   U15121 : XNOR2_X1 port map( A => n13042, B => n13695, ZN => n13044);
   U15122 : XNOR2_X1 port map( A => n13644, B => n2310, ZN => n13043);
   U15123 : XNOR2_X1 port map( A => n13044, B => n13043, ZN => n13045);
   U15124 : XNOR2_X1 port map( A => n13046, B => n13045, ZN => n14305);
   U15126 : XNOR2_X1 port map( A => n13103, B => n13047, ZN => n13417);
   U15127 : XNOR2_X1 port map( A => n13816, B => n13417, ZN => n13052);
   U15128 : XNOR2_X1 port map( A => n13048, B => n13192, ZN => n13050);
   U15129 : XNOR2_X1 port map( A => n13050, B => n13049, ZN => n13051);
   U15130 : INV_X1 port map( A => n14497, ZN => n14307);
   U15135 : XNOR2_X1 port map( A => n13579, B => n13057, ZN => n13062);
   U15136 : XNOR2_X1 port map( A => n13058, B => n13173, ZN => n13367);
   U15137 : XNOR2_X1 port map( A => n20199, B => n2216, ZN => n13060);
   U15138 : XNOR2_X1 port map( A => n13367, B => n13060, ZN => n13061);
   U15139 : XNOR2_X1 port map( A => n13400, B => n13573, ZN => n13069);
   U15141 : XNOR2_X1 port map( A => n19937, B => n13425, ZN => n13066);
   U15142 : XNOR2_X1 port map( A => n13067, B => n13066, ZN => n13068);
   U15143 : XNOR2_X2 port map( A => n13069, B => n13068, ZN => n14520);
   U15144 : XNOR2_X1 port map( A => n13070, B => n13584, ZN => n13072);
   U15145 : XNOR2_X1 port map( A => n19892, B => n17787, ZN => n13071);
   U15146 : XNOR2_X1 port map( A => n13072, B => n13071, ZN => n13075);
   U15147 : XNOR2_X1 port map( A => n13444, B => n13073, ZN => n13074);
   U15148 : XNOR2_X1 port map( A => n13074, B => n13075, ZN => n14321);
   U15149 : INV_X1 port map( A => n14321, ZN => n14186);
   U15150 : XNOR2_X1 port map( A => n13404, B => n2381, ZN => n13077);
   U15151 : AOI22_X1 port map( A1 => n15119, A2 => n14520, B1 => n14186, B2 => 
                           n14514, ZN => n13094);
   U15152 : XNOR2_X1 port map( A => n13080, B => n13389, ZN => n13084);
   U15153 : XNOR2_X1 port map( A => n13081, B => n13833, ZN => n13082);
   U15155 : XNOR2_X1 port map( A => n13085, B => n20482, ZN => n13087);
   U15156 : XNOR2_X1 port map( A => n13087, B => n13086, ZN => n13091);
   U15157 : XNOR2_X1 port map( A => n13616, B => n13618, ZN => n13089);
   U15158 : XNOR2_X1 port map( A => n13382, B => n13089, ZN => n13090);
   U15159 : XNOR2_X1 port map( A => n13091, B => n13090, ZN => n13563);
   U15160 : INV_X1 port map( A => n13563, ZN => n14516);
   U15161 : NAND2_X1 port map( A1 => n14514, A2 => n14520, ZN => n13092);
   U15162 : OAI21_X1 port map( B1 => n14519, B2 => n14520, A => n13092, ZN => 
                           n13093);
   U15163 : INV_X1 port map( A => n15686, ZN => n15685);
   U15164 : OAI21_X1 port map( B1 => n13096, B2 => n13095, A => n15685, ZN => 
                           n13182);
   U15167 : XNOR2_X1 port map( A => n13422, B => n2392, ZN => n13100);
   U15168 : XNOR2_X1 port map( A => n13099, B => n13688, ZN => n13299);
   U15169 : XNOR2_X1 port map( A => n13100, B => n13299, ZN => n13101);
   U15170 : XNOR2_X1 port map( A => n13103, B => n18887, ZN => n13104);
   U15171 : XNOR2_X1 port map( A => n13536, B => n13104, ZN => n13107);
   U15172 : XNOR2_X1 port map( A => n13724, B => n13336, ZN => n13105);
   U15173 : XNOR2_X1 port map( A => n13382, B => n13105, ZN => n13106);
   U15175 : INV_X1 port map( A => n13981, ZN => n14020);
   U15176 : XNOR2_X1 port map( A => n13319, B => n13716, ZN => n13284);
   U15177 : XNOR2_X1 port map( A => n13108, B => n2445, ZN => n13109);
   U15178 : XNOR2_X1 port map( A => n13284, B => n13109, ZN => n13113);
   U15179 : INV_X1 port map( A => n13110, ZN => n13111);
   U15180 : XNOR2_X1 port map( A => n13844, B => n13111, ZN => n13112);
   U15181 : XNOR2_X1 port map( A => n13530, B => n13367, ZN => n13117);
   U15182 : XNOR2_X1 port map( A => n13453, B => n16651, ZN => n13115);
   U15183 : XNOR2_X1 port map( A => n13114, B => n915, ZN => n13267);
   U15184 : XNOR2_X1 port map( A => n13267, B => n13115, ZN => n13116);
   U15185 : XNOR2_X1 port map( A => n13117, B => n13116, ZN => n13118);
   U15186 : INV_X1 port map( A => n13118, ZN => n14261);
   U15187 : INV_X1 port map( A => n13550, ZN => n13119);
   U15188 : XNOR2_X1 port map( A => n13119, B => n13389, ZN => n13124);
   U15189 : XNOR2_X1 port map( A => n13121, B => n18055, ZN => n13122);
   U15190 : XNOR2_X1 port map( A => n13313, B => n13122, ZN => n13123);
   U15191 : XNOR2_X1 port map( A => n13124, B => n13123, ZN => n13980);
   U15192 : INV_X1 port map( A => n13980, ZN => n14260);
   U15193 : NAND2_X1 port map( A1 => n20424, A2 => n14260, ZN => n13125);
   U15194 : OAI211_X1 port map( C1 => n14262, C2 => n14020, A => n14543, B => 
                           n13125, ZN => n13132);
   U15195 : XNOR2_X1 port map( A => n13126, B => n13374, ZN => n13131);
   U15196 : XNOR2_X1 port map( A => n13697, B => n19180, ZN => n13128);
   U15197 : INV_X1 port map( A => n13352, ZN => n13127);
   U15198 : XNOR2_X1 port map( A => n13128, B => n13127, ZN => n13129);
   U15199 : XNOR2_X1 port map( A => n13808, B => n13129, ZN => n13130);
   U15200 : XNOR2_X1 port map( A => n13130, B => n13131, ZN => n14673);
   U15201 : INV_X1 port map( A => n14673, ZN => n14266);
   U15202 : XNOR2_X1 port map( A => n13136, B => n2382, ZN => n13137);
   U15204 : INV_X1 port map( A => n13147, ZN => n13142);
   U15205 : NOR2_X1 port map( A1 => n13142, A2 => n13141, ZN => n13143);
   U15206 : OAI21_X1 port map( B1 => n13144, B2 => n13143, A => n13146, ZN => 
                           n13151);
   U15207 : NOR3_X1 port map( A1 => n13147, A2 => n13146, A3 => n13145, ZN => 
                           n13148);
   U15208 : NOR2_X1 port map( A1 => n13149, A2 => n13148, ZN => n13150);
   U15209 : NAND2_X1 port map( A1 => n13151, A2 => n13150, ZN => n13152);
   U15210 : XNOR2_X1 port map( A => n13152, B => n13321, ZN => n13595);
   U15211 : XNOR2_X1 port map( A => n13153, B => n13595, ZN => n13158);
   U15212 : XNOR2_X1 port map( A => n13154, B => n19904, ZN => n13156);
   U15213 : XNOR2_X1 port map( A => n13544, B => n2420, ZN => n13155);
   U15214 : XNOR2_X1 port map( A => n13156, B => n13155, ZN => n13157);
   U15215 : XNOR2_X1 port map( A => n13158, B => n13157, ZN => n14316);
   U15216 : INV_X1 port map( A => n13309, ZN => n13608);
   U15217 : XNOR2_X1 port map( A => n13608, B => n13834, ZN => n13160);
   U15218 : XNOR2_X1 port map( A => n13328, B => n2305, ZN => n13159);
   U15219 : XNOR2_X1 port map( A => n13160, B => n13159, ZN => n13163);
   U15220 : XNOR2_X1 port map( A => n13161, B => n13330, ZN => n13610);
   U15221 : XNOR2_X1 port map( A => n13610, B => n13486, ZN => n13162);
   U15222 : NAND2_X1 port map( A1 => n13166, A2 => n13165, ZN => n14538);
   U15223 : XNOR2_X1 port map( A => n13376, B => n19689, ZN => n13167);
   U15224 : XNOR2_X1 port map( A => n13490, B => n13167, ZN => n13171);
   U15225 : XNOR2_X1 port map( A => n13642, B => n2218, ZN => n13169);
   U15226 : XNOR2_X1 port map( A => n13590, B => n13168, ZN => n13523);
   U15227 : XNOR2_X1 port map( A => n13169, B => n13523, ZN => n13170);
   U15228 : XNOR2_X1 port map( A => n13577, B => n13266, ZN => n13172);
   U15229 : XNOR2_X1 port map( A => n13475, B => n13172, ZN => n13177);
   U15230 : XNOR2_X1 port map( A => n13173, B => n2442, ZN => n13175);
   U15231 : XNOR2_X1 port map( A => n20440, B => n13580, ZN => n13174);
   U15232 : XNOR2_X1 port map( A => n13175, B => n13174, ZN => n13176);
   U15233 : OAI211_X1 port map( C1 => n15687, C2 => n15683, A => n13180, B => 
                           n15686, ZN => n13181);
   U15234 : XNOR2_X1 port map( A => n13183, B => n17104, ZN => n13184);
   U15235 : XNOR2_X1 port map( A => n20253, B => n19158, ZN => n13185);
   U15236 : XNOR2_X1 port map( A => n13186, B => n13693, ZN => n13188);
   U15237 : INV_X1 port map( A => n13619, ZN => n13189);
   U15238 : XNOR2_X1 port map( A => n13222, B => n13189, ZN => n13190);
   U15239 : XNOR2_X1 port map( A => n13191, B => n13190, ZN => n13197);
   U15240 : XNOR2_X1 port map( A => n19923, B => n13192, ZN => n13195);
   U15241 : XNOR2_X1 port map( A => n13193, B => n17993, ZN => n13194);
   U15242 : XNOR2_X1 port map( A => n13195, B => n13194, ZN => n13196);
   U15243 : NOR2_X1 port map( A1 => n14654, A2 => n20266, ZN => n13221);
   U15244 : INV_X1 port map( A => n13673, ZN => n13198);
   U15245 : XNOR2_X1 port map( A => n13198, B => n13607, ZN => n13388);
   U15246 : XNOR2_X1 port map( A => n13199, B => n13388, ZN => n13202);
   U15247 : XNOR2_X1 port map( A => n13792, B => n2329, ZN => n13200);
   U15248 : XNOR2_X1 port map( A => n13733, B => n13200, ZN => n13201);
   U15249 : XNOR2_X1 port map( A => n19697, B => n2079, ZN => n13205);
   U15250 : XNOR2_X1 port map( A => n13206, B => n13207, ZN => n13208);
   U15251 : INV_X1 port map( A => n13708, ZN => n13212);
   U15252 : XNOR2_X1 port map( A => n13774, B => n620, ZN => n13210);
   U15253 : XNOR2_X1 port map( A => n13210, B => n13576, ZN => n13211);
   U15254 : XNOR2_X1 port map( A => n13212, B => n13211, ZN => n13214);
   U15255 : INV_X1 port map( A => n14022, ZN => n14653);
   U15256 : INV_X1 port map( A => n13215, ZN => n13216);
   U15257 : XNOR2_X1 port map( A => n13216, B => n13684, ZN => n13220);
   U15258 : XNOR2_X1 port map( A => n20469, B => n17932, ZN => n13217);
   U15259 : XNOR2_X1 port map( A => n13218, B => n13217, ZN => n13219);
   U15260 : INV_X1 port map( A => n13222, ZN => n13223);
   U15261 : XNOR2_X1 port map( A => n13616, B => n13223, ZN => n13225);
   U15262 : INV_X1 port map( A => n13764, ZN => n13224);
   U15263 : XNOR2_X1 port map( A => n13224, B => n13225, ZN => n13229);
   U15264 : XNOR2_X1 port map( A => n20260, B => n2298, ZN => n13226);
   U15265 : XOR2_X1 port map( A => n20226, B => n13226, Z => n13228);
   U15266 : XNOR2_X1 port map( A => n13231, B => n13230, ZN => n13665);
   U15267 : XNOR2_X1 port map( A => n13783, B => n18779, ZN => n13232);
   U15268 : XNOR2_X1 port map( A => n13665, B => n13232, ZN => n13236);
   U15270 : XNOR2_X1 port map( A => n13238, B => n13237, ZN => n13241);
   U15271 : XNOR2_X1 port map( A => n13309, B => n20222, ZN => n13239);
   U15272 : XNOR2_X1 port map( A => n13241, B => n13240, ZN => n14575);
   U15273 : MUX2_X1 port map( A => n14267, B => n14574, S => n14575, Z => 
                           n13264);
   U15274 : XNOR2_X1 port map( A => n13295, B => n2385, ZN => n13242);
   U15275 : XNOR2_X1 port map( A => n20442, B => n13243, ZN => n13245);
   U15276 : INV_X1 port map( A => n14570, ZN => n14738);
   U15277 : AND2_X1 port map( A1 => n14571, A2 => n14738, ZN => n14578);
   U15278 : XNOR2_X1 port map( A => n13642, B => n13810, ZN => n13247);
   U15279 : XNOR2_X1 port map( A => n13247, B => n13248, ZN => n13253);
   U15280 : XNOR2_X1 port map( A => n20123, B => n17587, ZN => n13249);
   U15281 : XNOR2_X1 port map( A => n13249, B => n19689, ZN => n13252);
   U15282 : XNOR2_X1 port map( A => n13251, B => n13250, ZN => n13750);
   U15283 : XNOR2_X1 port map( A => n13539, B => n2375, ZN => n13256);
   U15284 : XNOR2_X1 port map( A => n13257, B => n13256, ZN => n13262);
   U15285 : XNOR2_X1 port map( A => n13258, B => n13717, ZN => n13656);
   U15286 : XNOR2_X1 port map( A => n13260, B => n13259, ZN => n13769);
   U15287 : XNOR2_X1 port map( A => n13656, B => n13769, ZN => n13261);
   U15288 : XNOR2_X1 port map( A => n13702, B => n456, ZN => n13265);
   U15289 : XNOR2_X1 port map( A => n13266, B => n13265, ZN => n13268);
   U15290 : XNOR2_X1 port map( A => n13268, B => n13267, ZN => n13279);
   U15291 : INV_X1 port map( A => n13269, ZN => n13273);
   U15292 : INV_X1 port map( A => n13270, ZN => n13271);
   U15293 : NAND2_X1 port map( A1 => n13271, A2 => n13275, ZN => n13272);
   U15295 : XNOR2_X1 port map( A => n13276, B => n13277, ZN => n13278);
   U15296 : XNOR2_X1 port map( A => n13278, B => n13580, ZN => n13477);
   U15297 : INV_X1 port map( A => n13316, ZN => n14704);
   U15298 : INV_X1 port map( A => n13280, ZN => n13281);
   U15299 : XNOR2_X1 port map( A => n13281, B => n13602, ZN => n13501);
   U15300 : XNOR2_X1 port map( A => n13282, B => n13501, ZN => n13286);
   U15301 : XNOR2_X1 port map( A => n13711, B => n17851, ZN => n13283);
   U15302 : XNOR2_X1 port map( A => n13284, B => n13283, ZN => n13285);
   U15303 : NOR2_X1 port map( A1 => n14704, A2 => n14563, ZN => n13308);
   U15304 : XNOR2_X1 port map( A => n13491, B => n17535, ZN => n13288);
   U15305 : XNOR2_X1 port map( A => n13288, B => n13287, ZN => n13290);
   U15306 : XNOR2_X1 port map( A => n13290, B => n13289, ZN => n13292);
   U15307 : XNOR2_X1 port map( A => n13292, B => n13291, ZN => n14562);
   U15308 : INV_X1 port map( A => n14562, ZN => n14706);
   U15309 : INV_X1 port map( A => n13293, ZN => n13294);
   U15310 : XNOR2_X1 port map( A => n13757, B => n13294, ZN => n13463);
   U15311 : XNOR2_X1 port map( A => n13295, B => n645, ZN => n13297);
   U15312 : INV_X1 port map( A => n13686, ZN => n13296);
   U15313 : XNOR2_X1 port map( A => n13297, B => n13296, ZN => n13298);
   U15315 : XNOR2_X1 port map( A => n13572, B => n13299, ZN => n13300);
   U15316 : NOR2_X1 port map( A1 => n14706, A2 => n20498, ZN => n13955);
   U15317 : XNOR2_X1 port map( A => n13303, B => n13302, ZN => n13307);
   U15318 : XNOR2_X1 port map( A => n13724, B => n18726, ZN => n13304);
   U15319 : XNOR2_X1 port map( A => n13305, B => n13304, ZN => n13306);
   U15320 : XNOR2_X2 port map( A => n13307, B => n13306, ZN => n14566);
   U15321 : XNOR2_X1 port map( A => n13309, B => n2376, ZN => n13310);
   U15322 : XNOR2_X1 port map( A => n13311, B => n13310, ZN => n13315);
   U15323 : XNOR2_X1 port map( A => n13483, B => n13313, ZN => n13314);
   U15324 : MUX2_X1 port map( A => n14275, B => n14273, S => n14566, Z => 
                           n13317);
   U15326 : MUX2_X1 port map( A => n15673, B => n234, S => n15672, Z => n13461)
                           ;
   U15327 : INV_X1 port map( A => n13319, ZN => n13320);
   U15328 : XNOR2_X1 port map( A => n13321, B => n13320, ZN => n13323);
   U15329 : XNOR2_X1 port map( A => n13323, B => n13322, ZN => n13327);
   U15330 : XNOR2_X1 port map( A => n13405, B => n18439, ZN => n13324);
   U15331 : XNOR2_X1 port map( A => n13325, B => n13324, ZN => n13326);
   U15332 : XNOR2_X1 port map( A => n13328, B => n13479, ZN => n13839);
   U15333 : XNOR2_X1 port map( A => n13839, B => n13329, ZN => n13334);
   U15334 : XNOR2_X1 port map( A => n13390, B => n20064, ZN => n13331);
   U15335 : XNOR2_X1 port map( A => n13331, B => n13332, ZN => n13333);
   U15336 : XNOR2_X1 port map( A => n13334, B => n13333, ZN => n14690);
   U15338 : NAND2_X1 port map( A1 => n14385, A2 => n19895, ZN => n14387);
   U15339 : INV_X1 port map( A => n16366, ZN => n19296);
   U15340 : XNOR2_X1 port map( A => n13335, B => n19296, ZN => n13338);
   U15341 : XNOR2_X1 port map( A => n13624, B => n13336, ZN => n13337);
   U15342 : XNOR2_X1 port map( A => n13338, B => n13337, ZN => n13342);
   U15343 : XNOR2_X1 port map( A => n13339, B => n13618, ZN => n13760);
   U15344 : XNOR2_X1 port map( A => n13340, B => n13760, ZN => n13341);
   U15345 : NAND2_X1 port map( A1 => n14387, A2 => n200, ZN => n13365);
   U15346 : XNOR2_X1 port map( A => n13344, B => n13343, ZN => n13346);
   U15347 : INV_X1 port map( A => n13512, ZN => n13849);
   U15348 : XNOR2_X1 port map( A => n13849, B => n19052, ZN => n13345);
   U15349 : XNOR2_X1 port map( A => n13347, B => n13348, ZN => n13349);
   U15350 : XNOR2_X1 port map( A => n13745, B => n1969, ZN => n13350);
   U15351 : XNOR2_X1 port map( A => n13350, B => n13523, ZN => n13356);
   U15352 : XNOR2_X1 port map( A => n13352, B => n13351, ZN => n13354);
   U15353 : XNOR2_X1 port map( A => n13354, B => n13353, ZN => n13355);
   U15354 : XNOR2_X1 port map( A => n13356, B => n13355, ZN => n14127);
   U15355 : INV_X1 port map( A => n14127, ZN => n14695);
   U15356 : XNOR2_X1 port map( A => n13776, B => n19854, ZN => n13358);
   U15357 : XNOR2_X1 port map( A => n13357, B => n13358, ZN => n13363);
   U15358 : XNOR2_X1 port map( A => n13359, B => n20440, ZN => n13361);
   U15359 : XNOR2_X1 port map( A => n13361, B => n13360, ZN => n13362);
   U15360 : XNOR2_X1 port map( A => n13363, B => n13362, ZN => n13946);
   U15364 : NAND2_X1 port map( A1 => n15221, A2 => n15667, ZN => n15772);
   U15365 : XNOR2_X1 port map( A => n13367, B => n13366, ZN => n13373);
   U15366 : XNOR2_X1 port map( A => n13368, B => n13369, ZN => n13371);
   U15367 : XNOR2_X1 port map( A => n13528, B => Key(60), ZN => n13370);
   U15368 : XNOR2_X1 port map( A => n13371, B => n13370, ZN => n13372);
   U15371 : XNOR2_X1 port map( A => n13375, B => n13374, ZN => n13380);
   U15372 : XNOR2_X1 port map( A => n13376, B => n13643, ZN => n13378);
   U15373 : XNOR2_X1 port map( A => n20253, B => n18208, ZN => n13377);
   U15374 : XNOR2_X1 port map( A => n13378, B => n13377, ZN => n13379);
   U15375 : XNOR2_X1 port map( A => n13380, B => n13379, ZN => n14727);
   U15376 : INV_X1 port map( A => n14727, ZN => n14224);
   U15378 : XNOR2_X1 port map( A => n13382, B => n19824, ZN => n13387);
   U15379 : XNOR2_X1 port map( A => n13622, B => n2284, ZN => n13385);
   U15380 : XNOR2_X1 port map( A => n20170, B => n19923, ZN => n13384);
   U15381 : XOR2_X1 port map( A => n13384, B => n13385, Z => n13386);
   U15382 : XNOR2_X2 port map( A => n13387, B => n13386, ZN => n14729);
   U15383 : NAND2_X1 port map( A1 => n14224, A2 => n14729, ZN => n14227);
   U15384 : XNOR2_X1 port map( A => n13391, B => n13390, ZN => n13393);
   U15386 : INV_X1 port map( A => n14410, ZN => n14730);
   U15387 : NOR2_X1 port map( A1 => n20451, A2 => n14730, ZN => n13403);
   U15388 : XNOR2_X1 port map( A => n13397, B => n20469, ZN => n13570);
   U15389 : XNOR2_X1 port map( A => n13398, B => n18420, ZN => n13399);
   U15390 : XNOR2_X1 port map( A => n13400, B => n13399, ZN => n13401);
   U15391 : INV_X1 port map( A => n14137, ZN => n13953);
   U15392 : XNOR2_X1 port map( A => n13601, B => n18997, ZN => n13407);
   U15393 : XNOR2_X1 port map( A => n13404, B => n13405, ZN => n13406);
   U15394 : XNOR2_X1 port map( A => n13407, B => n13406, ZN => n13413);
   U15395 : XNOR2_X1 port map( A => n20489, B => n13658, ZN => n13411);
   U15396 : XNOR2_X1 port map( A => n13409, B => n13596, ZN => n13410);
   U15397 : XNOR2_X1 port map( A => n13411, B => n13410, ZN => n13412);
   U15398 : XNOR2_X1 port map( A => n13413, B => n13412, ZN => n14724);
   U15400 : XNOR2_X1 port map( A => n13415, B => n13416, ZN => n13421);
   U15401 : XNOR2_X1 port map( A => n19721, B => n15479, ZN => n13419);
   U15402 : INV_X1 port map( A => n13417, ZN => n13418);
   U15403 : XNOR2_X1 port map( A => n13419, B => n13418, ZN => n13420);
   U15404 : XNOR2_X1 port map( A => n13422, B => n2410, ZN => n13424);
   U15405 : XNOR2_X1 port map( A => n13462, B => n13756, ZN => n13423);
   U15406 : XNOR2_X1 port map( A => n13424, B => n13423, ZN => n13430);
   U15407 : INV_X1 port map( A => n13425, ZN => n13426);
   U15408 : XNOR2_X1 port map( A => n13426, B => n13427, ZN => n13652);
   U15409 : XNOR2_X1 port map( A => n13652, B => n13428, ZN => n13429);
   U15410 : XNOR2_X1 port map( A => n13430, B => n13429, ZN => n14553);
   U15411 : AND2_X1 port map( A1 => n14553, A2 => n14679, ZN => n14552);
   U15412 : INV_X1 port map( A => n14552, ZN => n14682);
   U15413 : INV_X1 port map( A => n13431, ZN => n13797);
   U15414 : XNOR2_X1 port map( A => n13434, B => n13433, ZN => n13435);
   U15415 : XNOR2_X1 port map( A => n13435, B => n13436, ZN => n14279);
   U15416 : INV_X1 port map( A => n14279, ZN => n13976);
   U15417 : XNOR2_X1 port map( A => n13767, B => n13657, ZN => n13438);
   U15418 : XNOR2_X1 port map( A => n13438, B => n13437, ZN => n13442);
   U15419 : XNOR2_X1 port map( A => n13710, B => n2208, ZN => n13439);
   U15420 : XNOR2_X1 port map( A => n13440, B => n13439, ZN => n13441);
   U15422 : NAND2_X1 port map( A1 => n13976, A2 => n14555, ZN => n14680);
   U15423 : NAND2_X1 port map( A1 => n14682, A2 => n14680, ZN => n13459);
   U15424 : INV_X1 port map( A => n13443, ZN => n13445);
   U15425 : XNOR2_X1 port map( A => n13444, B => n13445, ZN => n13450);
   U15426 : XNOR2_X1 port map( A => n13446, B => n17170, ZN => n13448);
   U15427 : XNOR2_X1 port map( A => n13448, B => n13447, ZN => n13449);
   U15428 : INV_X1 port map( A => n14554, ZN => n14678);
   U15429 : XNOR2_X1 port map( A => n13451, B => n2108, ZN => n13452);
   U15430 : XNOR2_X1 port map( A => n13452, B => n19854, ZN => n13455);
   U15431 : XNOR2_X1 port map( A => n13703, B => n13453, ZN => n13454);
   U15432 : XOR2_X1 port map( A => n13455, B => n13454, Z => n13456);
   U15433 : XNOR2_X1 port map( A => n13456, B => n13457, ZN => n14556);
   U15434 : OAI21_X1 port map( B1 => n14677, B2 => n14279, A => n14555, ZN => 
                           n13458);
   U15435 : INV_X1 port map( A => n14553, ZN => n14550);
   U15437 : XNOR2_X1 port map( A => n13462, B => n13651, ZN => n13685);
   U15438 : XNOR2_X1 port map( A => n13463, B => n13685, ZN => n13467);
   U15439 : XNOR2_X1 port map( A => n13849, B => n17095, ZN => n13465);
   U15441 : XNOR2_X1 port map( A => n13623, B => n484, ZN => n13469);
   U15442 : INV_X1 port map( A => n13471, ZN => n13472);
   U15443 : XNOR2_X1 port map( A => n13703, B => n13474, ZN => n13476);
   U15444 : XNOR2_X1 port map( A => n13475, B => n13476, ZN => n13478);
   U15445 : INV_X1 port map( A => n13479, ZN => n13480);
   U15446 : XNOR2_X1 port map( A => n13480, B => n13481, ZN => n13482);
   U15447 : XNOR2_X1 port map( A => n13483, B => n13482, ZN => n13488);
   U15448 : XNOR2_X1 port map( A => n13484, B => n404, ZN => n13485);
   U15449 : XNOR2_X1 port map( A => n13486, B => n13485, ZN => n13487);
   U15450 : INV_X1 port map( A => n14426, ZN => n14494);
   U15451 : NOR2_X1 port map( A1 => n14494, A2 => n14424, ZN => n14749);
   U15452 : XNOR2_X1 port map( A => n13490, B => n13489, ZN => n13496);
   U15453 : XNOR2_X1 port map( A => n13491, B => n13747, ZN => n13494);
   U15454 : INV_X1 port map( A => n13518, ZN => n13492);
   U15455 : XNOR2_X1 port map( A => n13492, B => n18848, ZN => n13493);
   U15456 : XNOR2_X1 port map( A => n13494, B => n13493, ZN => n13495);
   U15457 : XNOR2_X1 port map( A => n13495, B => n13496, ZN => n14493);
   U15458 : INV_X1 port map( A => n14425, ZN => n14427);
   U15459 : NOR2_X1 port map( A1 => n14427, A2 => n19728, ZN => n13504);
   U15460 : INV_X1 port map( A => n13497, ZN => n13498);
   U15461 : XNOR2_X1 port map( A => n13499, B => n13498, ZN => n13503);
   U15462 : XNOR2_X1 port map( A => n13543, B => n18177, ZN => n13500);
   U15463 : XNOR2_X1 port map( A => n13501, B => n13500, ZN => n13502);
   U15464 : AOI22_X1 port map( A1 => n14749, A2 => n1936, B1 => n13504, B2 => 
                           n14753, ZN => n13505);
   U15465 : MUX2_X1 port map( A => n19742, B => n14499, S => n14305, Z => 
                           n13509);
   U15467 : NOR2_X1 port map( A1 => n15457, A2 => n19759, ZN => n13561);
   U15468 : XNOR2_X1 port map( A => n13753, B => n13510, ZN => n13516);
   U15469 : XNOR2_X1 port map( A => n19869, B => n18801, ZN => n13513);
   U15470 : XNOR2_X1 port map( A => n13518, B => n13517, ZN => n13521);
   U15471 : XNOR2_X1 port map( A => n19892, B => n2383, ZN => n13520);
   U15472 : XNOR2_X1 port map( A => n13523, B => n13522, ZN => n13524);
   U15473 : XNOR2_X1 port map( A => n13524, B => n13744, ZN => n14434);
   U15474 : INV_X1 port map( A => n13525, ZN => n13526);
   U15475 : XNOR2_X1 port map( A => n13526, B => n13527, ZN => n13532);
   U15476 : XNOR2_X1 port map( A => n13528, B => n17637, ZN => n13529);
   U15477 : XNOR2_X1 port map( A => n13530, B => n13529, ZN => n13531);
   U15478 : XNOR2_X1 port map( A => n13532, B => n13531, ZN => n14435);
   U15480 : XNOR2_X1 port map( A => n13533, B => n13761, ZN => n13538);
   U15481 : XNOR2_X1 port map( A => n20482, B => n17791, ZN => n13535);
   U15482 : XNOR2_X1 port map( A => n13536, B => n13535, ZN => n13537);
   U15483 : XNOR2_X1 port map( A => n13538, B => n13537, ZN => n14172);
   U15484 : OAI21_X1 port map( B1 => n14487, B2 => n20263, A => n14172, ZN => 
                           n13555);
   U15487 : XNOR2_X1 port map( A => n13771, B => n13542, ZN => n13548);
   U15488 : XNOR2_X1 port map( A => n13601, B => n16030, ZN => n13546);
   U15489 : XNOR2_X1 port map( A => n13544, B => n13543, ZN => n13545);
   U15490 : XNOR2_X1 port map( A => n13545, B => n13546, ZN => n13547);
   U15491 : INV_X1 port map( A => n14172, ZN => n14480);
   U15492 : XNOR2_X1 port map( A => n13792, B => n2067, ZN => n13549);
   U15493 : XNOR2_X1 port map( A => n13551, B => n13550, ZN => n13552);
   U15494 : XNOR2_X1 port map( A => n13552, B => n13553, ZN => n14171);
   U15495 : NAND2_X1 port map( A1 => n14435, A2 => n14171, ZN => n14302);
   U15496 : OAI21_X1 port map( B1 => n3516, B2 => n14167, A => n14442, ZN => 
                           n13558);
   U15497 : NOR2_X1 port map( A1 => n701, A2 => n13918, ZN => n14440);
   U15498 : NAND3_X1 port map( A1 => n3516, A2 => n20262, A3 => n14441, ZN => 
                           n13556);
   U15499 : OAI21_X1 port map( B1 => n14448, B2 => n14447, A => n14451, ZN => 
                           n13560);
   U15502 : INV_X1 port map( A => n15457, ZN => n15460);
   U15503 : AOI21_X1 port map( B1 => n15353, B2 => n13566, A => n15460, ZN => 
                           n13567);
   U15504 : NOR2_X2 port map( A1 => n13568, A2 => n13567, ZN => n16601);
   U15505 : INV_X1 port map( A => n13569, ZN => n13571);
   U15506 : XNOR2_X1 port map( A => n13571, B => n13570, ZN => n13575);
   U15507 : XNOR2_X1 port map( A => n13572, B => n19436, ZN => n13574);
   U15508 : XNOR2_X1 port map( A => n13577, B => n13576, ZN => n13578);
   U15509 : XNOR2_X1 port map( A => n13579, B => n13578, ZN => n13583);
   U15510 : XNOR2_X1 port map( A => n13580, B => n649, ZN => n13581);
   U15511 : XNOR2_X1 port map( A => n13584, B => n13517, ZN => n13587);
   U15512 : XNOR2_X1 port map( A => n13746, B => n13585, ZN => n13586);
   U15513 : XNOR2_X1 port map( A => n13587, B => n13586, ZN => n13594);
   U15514 : XNOR2_X1 port map( A => n13491, B => n2055, ZN => n13592);
   U15515 : INV_X1 port map( A => n13588, ZN => n13589);
   U15516 : XNOR2_X1 port map( A => n13590, B => n13589, ZN => n13591);
   U15517 : XNOR2_X1 port map( A => n13592, B => n13591, ZN => n13593);
   U15519 : NOR2_X1 port map( A1 => n13994, A2 => n13996, ZN => n13630);
   U15521 : INV_X1 port map( A => n13596, ZN => n13597);
   U15522 : XNOR2_X1 port map( A => n13597, B => n13767, ZN => n13598);
   U15524 : XNOR2_X1 port map( A => n19904, B => n13601, ZN => n13604);
   U15525 : XNOR2_X1 port map( A => n13602, B => n16424, ZN => n13603);
   U15526 : XNOR2_X1 port map( A => n13604, B => n13603, ZN => n13605);
   U15527 : XNOR2_X1 port map( A => n13606, B => n13605, ZN => n14153);
   U15528 : INV_X1 port map( A => n14153, ZN => n14594);
   U15529 : XNOR2_X1 port map( A => n13608, B => n13607, ZN => n13609);
   U15530 : XNOR2_X1 port map( A => n13610, B => n13609, ZN => n13614);
   U15531 : XNOR2_X1 port map( A => n13797, B => n2337, ZN => n13611);
   U15532 : XNOR2_X1 port map( A => n13612, B => n13611, ZN => n13613);
   U15533 : XNOR2_X1 port map( A => n13614, B => n13613, ZN => n14395);
   U15537 : AND2_X1 port map( A1 => n13615, A2 => n14156, ZN => n13629);
   U15538 : XNOR2_X1 port map( A => n13617, B => n13616, ZN => n13621);
   U15539 : XNOR2_X1 port map( A => n20170, B => n13618, ZN => n13620);
   U15540 : XNOR2_X1 port map( A => n13621, B => n13620, ZN => n13628);
   U15541 : XNOR2_X1 port map( A => n13622, B => n18203, ZN => n13626);
   U15542 : XNOR2_X1 port map( A => n13624, B => n13623, ZN => n13625);
   U15543 : XNOR2_X1 port map( A => n13626, B => n13625, ZN => n13627);
   U15545 : INV_X1 port map( A => n13631, ZN => n13632);
   U15547 : XNOR2_X1 port map( A => n20260, B => n13635, ZN => n13637);
   U15548 : XNOR2_X1 port map( A => n13637, B => n13636, ZN => n13638);
   U15549 : INV_X1 port map( A => n14388, ZN => n14715);
   U15550 : XNOR2_X1 port map( A => n13641, B => n13640, ZN => n13648);
   U15551 : XNOR2_X1 port map( A => n13643, B => n13642, ZN => n13646);
   U15552 : XNOR2_X1 port map( A => n13644, B => n2394, ZN => n13645);
   U15553 : XNOR2_X1 port map( A => n13646, B => n13645, ZN => n13647);
   U15554 : XNOR2_X1 port map( A => n13648, B => n13647, ZN => n14716);
   U15555 : NAND2_X1 port map( A1 => n14715, A2 => n14716, ZN => n14389);
   U15556 : XNOR2_X1 port map( A => n13651, B => n17060, ZN => n13653);
   U15557 : XNOR2_X1 port map( A => n13652, B => n13653, ZN => n13654);
   U15558 : XNOR2_X1 port map( A => n13656, B => n13655, ZN => n13663);
   U15559 : XNOR2_X1 port map( A => n13658, B => n13657, ZN => n13661);
   U15560 : XNOR2_X1 port map( A => n13659, B => n17365, ZN => n13660);
   U15561 : XNOR2_X1 port map( A => n13661, B => n13660, ZN => n13662);
   U15563 : NAND2_X1 port map( A1 => n20213, A2 => n19843, ZN => n13664);
   U15564 : OAI21_X1 port map( B1 => n14389, B2 => n19843, A => n13664, ZN => 
                           n13683);
   U15565 : XNOR2_X1 port map( A => n13666, B => n13665, ZN => n13670);
   U15566 : XNOR2_X1 port map( A => n13827, B => n2221, ZN => n13667);
   U15567 : XNOR2_X1 port map( A => n13668, B => n13667, ZN => n13669);
   U15568 : NAND2_X1 port map( A1 => n14716, A2 => n14717, ZN => n13682);
   U15569 : XNOR2_X1 port map( A => n13833, B => n13672, ZN => n13675);
   U15570 : XNOR2_X1 port map( A => n13673, B => n1996, ZN => n13674);
   U15571 : XNOR2_X1 port map( A => n13675, B => n13674, ZN => n13681);
   U15572 : INV_X1 port map( A => n13676, ZN => n13679);
   U15573 : XNOR2_X1 port map( A => n13734, B => n13677, ZN => n13678);
   U15574 : XNOR2_X1 port map( A => n13679, B => n13678, ZN => n13680);
   U15575 : INV_X1 port map( A => n14718, ZN => n13963);
   U15577 : XNOR2_X1 port map( A => n13684, B => n13685, ZN => n13692);
   U15578 : XNOR2_X1 port map( A => n13686, B => n13687, ZN => n13690);
   U15579 : XNOR2_X1 port map( A => n13688, B => n18366, ZN => n13689);
   U15580 : XNOR2_X1 port map( A => n13690, B => n13689, ZN => n13691);
   U15581 : INV_X1 port map( A => n14378, ZN => n14232);
   U15582 : XNOR2_X1 port map( A => n13694, B => n13693, ZN => n13701);
   U15585 : XNOR2_X1 port map( A => n13699, B => n13698, ZN => n13700);
   U15586 : XNOR2_X1 port map( A => n13701, B => n13700, ZN => n14700);
   U15587 : NOR2_X1 port map( A1 => n14232, A2 => n14700, ZN => n13731);
   U15588 : XNOR2_X1 port map( A => n20155, B => n13703, ZN => n13704);
   U15589 : INV_X1 port map( A => n915, ZN => n13705);
   U15590 : XNOR2_X1 port map( A => n13707, B => n13706, ZN => n13709);
   U15591 : XNOR2_X1 port map( A => n13710, B => n18308, ZN => n13712);
   U15592 : XNOR2_X1 port map( A => n13712, B => n13711, ZN => n13713);
   U15593 : XNOR2_X1 port map( A => n13714, B => n13713, ZN => n13720);
   U15594 : XNOR2_X1 port map( A => n13716, B => n13715, ZN => n13718);
   U15595 : XNOR2_X1 port map( A => n13718, B => n13717, ZN => n13719);
   U15596 : NOR2_X1 port map( A1 => n14120, A2 => n14228, ZN => n13730);
   U15597 : XNOR2_X1 port map( A => n19721, B => n2248, ZN => n13723);
   U15598 : XNOR2_X1 port map( A => n13722, B => n13723, ZN => n13729);
   U15599 : XNOR2_X1 port map( A => n13724, B => n13725, ZN => n13726);
   U15600 : XNOR2_X1 port map( A => n13727, B => n13726, ZN => n13728);
   U15602 : XNOR2_X1 port map( A => n13733, B => n13732, ZN => n13740);
   U15603 : XNOR2_X1 port map( A => n13735, B => n13734, ZN => n13738);
   U15604 : INV_X1 port map( A => n1148, ZN => n18587);
   U15605 : XNOR2_X1 port map( A => n13736, B => n18587, ZN => n13737);
   U15606 : XNOR2_X1 port map( A => n13738, B => n13737, ZN => n13739);
   U15607 : MUX2_X1 port map( A => n2769, B => n14230, S => n240, Z => n13741);
   U15608 : NOR2_X1 port map( A1 => n13741, A2 => n20204, ZN => n13742);
   U15609 : NAND2_X1 port map( A1 => n15228, A2 => n15677, ZN => n15229);
   U15610 : OAI21_X1 port map( B1 => n2005, B2 => n15679, A => n15229, ZN => 
                           n13806);
   U15611 : INV_X1 port map( A => n13744, ZN => n13752);
   U15612 : XNOR2_X1 port map( A => n13746, B => n13745, ZN => n13749);
   U15613 : XNOR2_X1 port map( A => n13747, B => n2032, ZN => n13748);
   U15614 : XNOR2_X1 port map( A => n13751, B => n13752, ZN => n14406);
   U15615 : INV_X1 port map( A => n14406, ZN => n14149);
   U15616 : XNOR2_X1 port map( A => n13755, B => n18830, ZN => n13759);
   U15617 : XNOR2_X1 port map( A => n13757, B => n13756, ZN => n13758);
   U15618 : XNOR2_X1 port map( A => n13761, B => n13760, ZN => n13766);
   U15619 : XNOR2_X1 port map( A => n13762, B => n18090, ZN => n13763);
   U15620 : XNOR2_X1 port map( A => n13764, B => n13763, ZN => n13765);
   U15622 : INV_X1 port map( A => n19907, ZN => n14405);
   U15623 : NOR2_X1 port map( A1 => n14148, A2 => n14405, ZN => n13789);
   U15624 : XNOR2_X1 port map( A => n13768, B => n13767, ZN => n13770);
   U15625 : XNOR2_X1 port map( A => n13772, B => n18070, ZN => n13773);
   U15626 : INV_X1 port map( A => n13774, ZN => n13775);
   U15627 : XNOR2_X1 port map( A => n13776, B => n13775, ZN => n13780);
   U15628 : XNOR2_X1 port map( A => n13778, B => n19854, ZN => n13779);
   U15629 : XNOR2_X1 port map( A => n13780, B => n13779, ZN => n13787);
   U15630 : XNOR2_X1 port map( A => n19797, B => n915, ZN => n13785);
   U15631 : XNOR2_X1 port map( A => n13783, B => n2349, ZN => n13784);
   U15632 : XNOR2_X1 port map( A => n13785, B => n13784, ZN => n13786);
   U15633 : XNOR2_X1 port map( A => n13787, B => n13786, ZN => n14112);
   U15634 : INV_X1 port map( A => n14112, ZN => n14238);
   U15635 : NOR2_X1 port map( A1 => n14236, A2 => n14238, ZN => n13788);
   U15636 : AOI22_X1 port map( A1 => n14149, A2 => n13789, B1 => n14405, B2 => 
                           n13788, ZN => n13804);
   U15637 : XNOR2_X1 port map( A => n13790, B => n13791, ZN => n13794);
   U15638 : XNOR2_X1 port map( A => n13794, B => n13793, ZN => n13801);
   U15639 : XNOR2_X1 port map( A => n19946, B => n13795, ZN => n13799);
   U15640 : XNOR2_X1 port map( A => n13797, B => n18304, ZN => n13798);
   U15641 : XNOR2_X1 port map( A => n13799, B => n13798, ZN => n13800);
   U15642 : INV_X1 port map( A => n14239, ZN => n14403);
   U15643 : MUX2_X1 port map( A => n19908, B => n14238, S => n14403, Z => 
                           n13802);
   U15644 : NAND2_X1 port map( A1 => n15682, A2 => n15442, ZN => n13805);
   U15645 : NAND2_X1 port map( A1 => n13806, A2 => n13805, ZN => n13863);
   U15646 : INV_X1 port map( A => n13807, ZN => n13809);
   U15647 : XNOR2_X1 port map( A => n13809, B => n13808, ZN => n13814);
   U15648 : XNOR2_X1 port map( A => n13810, B => n19410, ZN => n13811);
   U15649 : XNOR2_X1 port map( A => n13812, B => n13811, ZN => n13813);
   U15650 : XNOR2_X1 port map( A => n13816, B => n13815, ZN => n13822);
   U15651 : INV_X1 port map( A => n13817, ZN => n13820);
   U15652 : XNOR2_X1 port map( A => n13818, B => n18338, ZN => n13819);
   U15653 : XNOR2_X1 port map( A => n13820, B => n13819, ZN => n13821);
   U15654 : INV_X1 port map( A => n13823, ZN => n13825);
   U15655 : XNOR2_X1 port map( A => n13825, B => n13824, ZN => n13832);
   U15656 : INV_X1 port map( A => n13826, ZN => n13828);
   U15657 : XNOR2_X1 port map( A => n13827, B => n13828, ZN => n13830);
   U15658 : XNOR2_X1 port map( A => n13830, B => n13829, ZN => n13831);
   U15659 : XNOR2_X2 port map( A => n13832, B => n13831, ZN => n14599);
   U15660 : XNOR2_X1 port map( A => n13834, B => n13833, ZN => n13837);
   U15661 : XNOR2_X1 port map( A => n20223, B => n1911, ZN => n13836);
   U15662 : XNOR2_X1 port map( A => n13837, B => n13836, ZN => n13841);
   U15663 : XNOR2_X1 port map( A => n13839, B => n13838, ZN => n13840);
   U15664 : XNOR2_X1 port map( A => n13840, B => n13841, ZN => n14249);
   U15665 : INV_X1 port map( A => n13844, ZN => n13845);
   U15666 : XNOR2_X1 port map( A => n13845, B => n13846, ZN => n13847);
   U15667 : XNOR2_X1 port map( A => n13849, B => n18278, ZN => n13850);
   U15668 : XNOR2_X1 port map( A => n13853, B => n13852, ZN => n13854);
   U15670 : INV_X1 port map( A => n15312, ZN => n13861);
   U15671 : INV_X1 port map( A => n13856, ZN => n13857);
   U15672 : OAI21_X1 port map( B1 => n13857, B2 => n14146, A => n19875, ZN => 
                           n13858);
   U15673 : INV_X1 port map( A => n15676, ZN => n13859);
   U15674 : OAI21_X1 port map( B1 => n13859, B2 => n15442, A => n15679, ZN => 
                           n13860);
   U15675 : XOR2_X1 port map( A => n16601, B => n17288, Z => n13864);
   U15676 : INV_X1 port map( A => n17223, ZN => n16634);
   U15677 : MUX2_X1 port map( A => n15120, B => n14520, S => n14516, Z => 
                           n13867);
   U15678 : NAND2_X1 port map( A1 => n14186, A2 => n14520, ZN => n13866);
   U15679 : NAND2_X1 port map( A1 => n14499, A2 => n14497, ZN => n14306);
   U15680 : NOR2_X1 port map( A1 => n19742, A2 => n13868, ZN => n13871);
   U15681 : NAND2_X1 port map( A1 => n14305, A2 => n14307, ZN => n13870);
   U15682 : MUX2_X1 port map( A => n19634, B => n19831, S => n14648, Z => 
                           n13875);
   U15683 : AOI21_X1 port map( B1 => n20380, B2 => n14651, A => n237, ZN => 
                           n13874);
   U15684 : NAND2_X1 port map( A1 => n14648, A2 => n14524, ZN => n13873);
   U15685 : INV_X1 port map( A => n14042, ZN => n13887);
   U15686 : NOR2_X1 port map( A1 => n15500, A2 => n19512, ZN => n15160);
   U15687 : INV_X1 port map( A => n15500, ZN => n15497);
   U15688 : INV_X1 port map( A => n14753, ZN => n13880);
   U15689 : NAND2_X1 port map( A1 => n14427, A2 => n19727, ZN => n14750);
   U15690 : OAI21_X1 port map( B1 => n14494, B2 => n19727, A => n14750, ZN => 
                           n13879);
   U15691 : NAND3_X1 port map( A1 => n14494, A2 => n14424, A3 => n1936, ZN => 
                           n13876);
   U15692 : OAI21_X1 port map( B1 => n13877, B2 => n3156, A => n13876, ZN => 
                           n13878);
   U15693 : INV_X1 port map( A => n15195, ZN => n14041);
   U15694 : NOR2_X1 port map( A1 => n14482, A2 => n14435, ZN => n13882);
   U15695 : MUX2_X1 port map( A => n13882, B => n13881, S => n14480, Z => 
                           n13885);
   U15696 : INV_X1 port map( A => n14171, ZN => n14483);
   U15697 : NOR3_X1 port map( A1 => n14431, A2 => n13883, A3 => n14487, ZN => 
                           n13884);
   U15698 : NOR2_X2 port map( A1 => n13885, A2 => n13884, ZN => n15501);
   U15699 : OAI211_X1 port map( C1 => n15497, C2 => n14041, A => n15501, B => 
                           n15192, ZN => n13886);
   U15700 : XNOR2_X1 port map( A => n16587, B => n17686, ZN => n13945);
   U15701 : NOR2_X1 port map( A1 => n14813, A2 => n14807, ZN => n13888);
   U15702 : NAND2_X1 port map( A1 => n14199, A2 => n14810, ZN => n14141);
   U15703 : MUX2_X1 port map( A => n14811, B => n19781, S => n14199, Z => 
                           n13889);
   U15704 : NOR2_X1 port map( A1 => n13889, A2 => n14812, ZN => n13890);
   U15705 : NOR2_X1 port map( A1 => n20500, A2 => n14800, ZN => n13896);
   U15706 : NAND2_X1 port map( A1 => n13893, A2 => n3497, ZN => n13895);
   U15707 : INV_X1 port map( A => n14787, ZN => n14346);
   U15708 : NOR2_X1 port map( A1 => n14791, A2 => n12627, ZN => n13900);
   U15709 : NOR2_X1 port map( A1 => n14346, A2 => n12627, ZN => n14100);
   U15710 : NAND2_X1 port map( A1 => n14100, A2 => n14788, ZN => n13899);
   U15711 : NAND2_X1 port map( A1 => n14789, A2 => n12627, ZN => n13898);
   U15712 : OAI211_X1 port map( C1 => n14102, C2 => n13900, A => n13899, B => 
                           n13898, ZN => n15861);
   U15713 : INV_X1 port map( A => n15861, ZN => n15327);
   U15714 : INV_X1 port map( A => n13901, ZN => n14076);
   U15715 : NOR2_X1 port map( A1 => n877, A2 => n14076, ZN => n13904);
   U15716 : NAND2_X1 port map( A1 => n14077, A2 => n14782, ZN => n13903);
   U15718 : NAND2_X1 port map( A1 => n20408, A2 => n14076, ZN => n13902);
   U15719 : INV_X1 port map( A => n14779, ZN => n14216);
   U15720 : NOR2_X1 port map( A1 => n13905, A2 => n14216, ZN => n13906);
   U15721 : AOI21_X1 port map( B1 => n14612, B2 => n14206, A => n13908, ZN => 
                           n13911);
   U15722 : INV_X1 port map( A => n14011, ZN => n13907);
   U15723 : INV_X1 port map( A => n13909, ZN => n14142);
   U15724 : OAI21_X1 port map( B1 => n14207, B2 => n14142, A => n19488, ZN => 
                           n13910);
   U15725 : NOR2_X1 port map( A1 => n15866, A2 => n15863, ZN => n13912);
   U15727 : INV_X1 port map( A => n14827, ZN => n14073);
   U15728 : MUX2_X1 port map( A => n13914, B => n13913, S => n14073, Z => 
                           n13915);
   U15729 : NOR2_X1 port map( A1 => n15720, A2 => n15861, ZN => n15721);
   U15732 : NOR2_X1 port map( A1 => n13918, A2 => n14441, ZN => n13919);
   U15733 : NOR2_X1 port map( A1 => n13921, A2 => n14465, ZN => n13923);
   U15734 : NOR2_X1 port map( A1 => n14462, A2 => n14468, ZN => n13922);
   U15735 : MUX2_X1 port map( A => n13923, B => n13922, S => n19657, Z => 
                           n13926);
   U15736 : NAND2_X1 port map( A1 => n13921, A2 => n14468, ZN => n14363);
   U15737 : NAND2_X1 port map( A1 => n1363, A2 => n14449, ZN => n13928);
   U15738 : NAND2_X1 port map( A1 => n14450, A2 => n14449, ZN => n14182);
   U15739 : NAND3_X1 port map( A1 => n14448, A2 => n14455, A3 => n14451, ZN => 
                           n13929);
   U15740 : OAI21_X1 port map( B1 => n14182, B2 => n14453, A => n13929, ZN => 
                           n14755);
   U15741 : OAI21_X1 port map( B1 => n13930, B2 => n14335, A => n14092, ZN => 
                           n13932);
   U15742 : NOR2_X1 port map( A1 => n14424, A2 => n1936, ZN => n13936);
   U15743 : OAI211_X1 port map( C1 => n14424, C2 => n14493, A => n19728, B => 
                           n14753, ZN => n13935);
   U15744 : NOR3_X1 port map( A1 => n15187, A2 => n15505, A3 => n13933, ZN => 
                           n13943);
   U15745 : NOR2_X1 port map( A1 => n13939, A2 => n14359, ZN => n13941);
   U15746 : NOR2_X1 port map( A1 => n14054, A2 => n14357, ZN => n14757);
   U15747 : NAND3_X1 port map( A1 => n15187, A2 => n15188, A3 => n15507, ZN => 
                           n13942);
   U15748 : XNOR2_X1 port map( A => n16931, B => n19659, ZN => n13944);
   U15749 : XNOR2_X1 port map( A => n13945, B => n13944, ZN => n14018);
   U15750 : INV_X1 port map( A => n13946, ZN => n14691);
   U15751 : MUX2_X1 port map( A => n14385, B => n19895, S => n14691, Z => 
                           n13948);
   U15752 : NAND2_X1 port map( A1 => n14693, A2 => n14688, ZN => n13947);
   U15753 : INV_X1 port map( A => n14021, ZN => n14289);
   U15754 : INV_X1 port map( A => n15153, ZN => n16012);
   U15755 : NOR2_X1 port map( A1 => n14223, A2 => n14729, ZN => n13952);
   U15756 : NOR2_X1 port map( A1 => n14273, A2 => n14275, ZN => n13954);
   U15757 : OAI21_X1 port map( B1 => n13955, B2 => n13954, A => n2282, ZN => 
                           n13958);
   U15758 : NAND3_X1 port map( A1 => n14705, A2 => n14563, A3 => n14566, ZN => 
                           n13956);
   U15760 : INV_X1 port map( A => n15705, ZN => n13961);
   U15761 : NAND3_X1 port map( A1 => n14736, A2 => n14571, A3 => n14269, ZN => 
                           n13960);
   U15762 : NAND3_X1 port map( A1 => n14740, A2 => n20157, A3 => n14570, ZN => 
                           n13959);
   U15763 : INV_X1 port map( A => n20119, ZN => n15152);
   U15764 : MUX2_X1 port map( A => n13963, B => n20213, S => n3057, Z => n13965
                           );
   U15765 : NAND2_X1 port map( A1 => n19843, A2 => n14715, ZN => n13964);
   U15766 : NAND3_X1 port map( A1 => n13965, A2 => n14389, A3 => n13964, ZN => 
                           n13967);
   U15767 : NAND2_X1 port map( A1 => n14716, A2 => n19862, ZN => n13966);
   U15768 : AND2_X2 port map( A1 => n13967, A2 => n13966, ZN => n16009);
   U15769 : INV_X1 port map( A => n16009, ZN => n13968);
   U15770 : INV_X1 port map( A => n17281, ZN => n13992);
   U15771 : NOR2_X1 port map( A1 => n14651, A2 => n14522, ZN => n13971);
   U15773 : NAND2_X1 port map( A1 => n14677, A2 => n13976, ZN => n13979);
   U15774 : INV_X1 port map( A => n14679, ZN => n14557);
   U15775 : AOI21_X1 port map( B1 => n14554, B2 => n14553, A => n14557, ZN => 
                           n13977);
   U15777 : INV_X1 port map( A => n14281, ZN => n14284);
   U15779 : NAND3_X1 port map( A1 => n15870, A2 => n20178, A3 => n13989, ZN => 
                           n13991);
   U15780 : INV_X1 port map( A => n14032, ZN => n14640);
   U15782 : INV_X1 port map( A => n14642, ZN => n13983);
   U15783 : NOR2_X1 port map( A1 => n20473, A2 => n13983, ZN => n13984);
   U15784 : MUX2_X1 port map( A => n13985, B => n13984, S => n19703, Z => 
                           n13988);
   U15785 : INV_X1 port map( A => n14512, ZN => n14034);
   U15786 : OAI22_X1 port map( A1 => n14508, A2 => n14034, B1 => n13986, B2 => 
                           n14642, ZN => n13987);
   U15787 : NOR2_X2 port map( A1 => n13988, A2 => n13987, ZN => n15875);
   U15788 : INV_X1 port map( A => n15875, ZN => n15148);
   U15789 : NOR2_X1 port map( A1 => n15876, A2 => n15709, ZN => n15303);
   U15790 : XNOR2_X1 port map( A => n13992, B => n16566, ZN => n16713);
   U15791 : NAND2_X1 port map( A1 => n15028, A2 => n15380, ZN => n14874);
   U15792 : INV_X1 port map( A => n14874, ZN => n15170);
   U15793 : NOR2_X1 port map( A1 => n19513, A2 => n231, ZN => n14872);
   U15794 : OAI21_X1 port map( B1 => n15167, B2 => n15380, A => n14872, ZN => 
                           n13993);
   U15796 : MUX2_X1 port map( A => n19709, B => n13994, S => n14395, Z => 
                           n13999);
   U15797 : NOR2_X1 port map( A1 => n14594, A2 => n14396, ZN => n13997);
   U15798 : MUX2_X1 port map( A => n13997, B => n13996, S => n19731, Z => 
                           n13998);
   U15799 : AOI22_X1 port map( A1 => n954, A2 => n14624, B1 => n15314, B2 => 
                           n14623, ZN => n14004);
   U15800 : NOR2_X1 port map( A1 => n14627, A2 => n14624, ZN => n14003);
   U15801 : NAND3_X1 port map( A1 => n14001, A2 => n14620, A3 => n14146, ZN => 
                           n14002);
   U15803 : INV_X1 port map( A => n15695, ZN => n15138);
   U15804 : NAND2_X1 port map( A1 => n15701, A2 => n15138, ZN => n14016);
   U15805 : NAND2_X1 port map( A1 => n14381, A2 => n20204, ZN => n14005);
   U15806 : OAI21_X1 port map( B1 => n14120, B2 => n14229, A => n20480, ZN => 
                           n14006);
   U15808 : NAND2_X1 port map( A1 => n14238, A2 => n19908, ZN => n14240);
   U15809 : OAI21_X1 port map( B1 => n14238, B2 => n14148, A => n14240, ZN => 
                           n14007);
   U15810 : NOR2_X1 port map( A1 => n20005, A2 => n15698, ZN => n14015);
   U15811 : MUX2_X1 port map( A => n14203, B => n13908, S => n3225, Z => n14014
                           );
   U15814 : XNOR2_X1 port map( A => n17275, B => n16926, ZN => n16523);
   U15815 : XNOR2_X1 port map( A => n16523, B => n19903, ZN => n14017);
   U15816 : XNOR2_X1 port map( A => n14017, B => n14018, ZN => n16633);
   U15819 : AOI21_X1 port map( B1 => n14654, B2 => n241, A => n14288, ZN => 
                           n14025);
   U15820 : OAI211_X1 port map( C1 => n14268, C2 => n14267, A => n14269, B => 
                           n1819, ZN => n14027);
   U15821 : NAND2_X1 port map( A1 => n14578, A2 => n14268, ZN => n15487);
   U15822 : OAI21_X1 port map( B1 => n15756, B2 => n15754, A => n15758, ZN => 
                           n14040);
   U15823 : MUX2_X1 port map( A => n14677, B => n14554, S => n14550, Z => 
                           n14030);
   U15824 : INV_X1 port map( A => n14555, ZN => n14028);
   U15825 : MUX2_X1 port map( A => n14279, B => n14028, S => n14677, Z => 
                           n14029);
   U15826 : OAI21_X1 port map( B1 => n14032, B2 => n14031, A => n20473, ZN => 
                           n14033);
   U15827 : NAND2_X1 port map( A1 => n15491, A2 => n15760, ZN => n14039);
   U15828 : NOR2_X1 port map( A1 => n14667, A2 => n14662, ZN => n14035);
   U15829 : NAND3_X1 port map( A1 => n14663, A2 => n14316, A3 => n14664, ZN => 
                           n14036);
   U15830 : AND3_X1 port map( A1 => n14038, A2 => n14037, A3 => n14036, ZN => 
                           n15490);
   U15831 : NOR2_X1 port map( A1 => n15501, A2 => n15192, ZN => n14930);
   U15832 : OAI21_X1 port map( B1 => n14930, B2 => n15496, A => n19813, ZN => 
                           n14044);
   U15833 : NAND2_X1 port map( A1 => n14042, A2 => n14041, ZN => n14043);
   U15834 : NAND2_X1 port map( A1 => n14044, A2 => n14043, ZN => n16821);
   U15835 : XNOR2_X1 port map( A => n16821, B => n16743, ZN => n16396);
   U15836 : NOR2_X1 port map( A1 => n14347, A2 => n14827, ZN => n14045);
   U15838 : INV_X1 port map( A => n14049, ZN => n14051);
   U15839 : AOI22_X2 port map( A1 => n14341, A2 => n14051, B1 => n14093, B2 => 
                           n14050, ZN => n15844);
   U15840 : NOR2_X1 port map( A1 => n15845, A2 => n15844, ZN => n14056);
   U15841 : NOR2_X1 port map( A1 => n14419, A2 => n14357, ZN => n14053);
   U15843 : OAI21_X1 port map( B1 => n14056, B2 => n15266, A => n15636, ZN => 
                           n14068);
   U15844 : NAND2_X1 port map( A1 => n20454, A2 => n14778, ZN => n14058);
   U15845 : AOI21_X1 port map( B1 => n14852, B2 => n14058, A => n14057, ZN => 
                           n14061);
   U15846 : NAND2_X1 port map( A1 => n14076, A2 => n14778, ZN => n14059);
   U15847 : AOI21_X1 port map( B1 => n20454, B2 => n14059, A => n14216, ZN => 
                           n14060);
   U15848 : NOR2_X2 port map( A1 => n14061, A2 => n14060, ZN => n15846);
   U15849 : INV_X1 port map( A => n14788, ZN => n14066);
   U15850 : MUX2_X1 port map( A => n14789, B => n2412, S => n14790, Z => n14065
                           );
   U15852 : NAND2_X1 port map( A1 => n14791, A2 => n14792, ZN => n14062);
   U15853 : MUX2_X1 port map( A => n14063, B => n14062, S => n14789, Z => 
                           n14064);
   U15854 : NAND3_X1 port map( A1 => n15847, A2 => n2146, A3 => n868, ZN => 
                           n14067);
   U15855 : NOR2_X1 port map( A1 => n15187, A2 => n15505, ZN => n14069);
   U15856 : NOR2_X1 port map( A1 => n15187, A2 => n1614, ZN => n14070);
   U15858 : XNOR2_X1 port map( A => n16593, B => n864, ZN => n16185);
   U15859 : MUX2_X1 port map( A => n14073, B => n14828, S => n19496, Z => 
                           n14075);
   U15860 : MUX2_X1 port map( A => n19859, B => n19984, S => n14827, Z => 
                           n14074);
   U15861 : NAND2_X1 port map( A1 => n14077, A2 => n14778, ZN => n14078);
   U15862 : NOR2_X1 port map( A1 => n14057, A2 => n20518, ZN => n14079);
   U15863 : NAND2_X1 port map( A1 => n14079, A2 => n14216, ZN => n14080);
   U15864 : OAI21_X1 port map( B1 => n14796, B2 => n14584, A => n14799, ZN => 
                           n14082);
   U15865 : INV_X1 port map( A => n15515, ZN => n15745);
   U15866 : INV_X1 port map( A => n14085, ZN => n14091);
   U15867 : INV_X1 port map( A => n14086, ZN => n14089);
   U15868 : OAI211_X1 port map( C1 => n19821, C2 => n14818, A => n912, B => 
                           n14326, ZN => n14088);
   U15869 : AOI21_X1 port map( B1 => n19485, B2 => n12876, A => n14092, ZN => 
                           n14098);
   U15870 : INV_X1 port map( A => n14093, ZN => n14096);
   U15871 : NOR2_X1 port map( A1 => n14336, A2 => n14335, ZN => n14095);
   U15873 : NAND3_X1 port map( A1 => n15521, A2 => n15516, A3 => n15741, ZN => 
                           n14099);
   U15874 : OAI21_X1 port map( B1 => n15748, B2 => n14982, A => n14099, ZN => 
                           n14108);
   U15875 : INV_X1 port map( A => n14100, ZN => n14101);
   U15876 : NAND2_X1 port map( A1 => n15746, A2 => n15516, ZN => n15740);
   U15877 : INV_X1 port map( A => n15748, ZN => n15181);
   U15878 : AOI21_X1 port map( B1 => n15740, B2 => n15741, A => n15181, ZN => 
                           n14107);
   U15879 : MUX2_X1 port map( A => n14717, B => n14718, S => n3057, Z => n14110
                           );
   U15880 : MUX2_X1 port map( A => n14716, B => n3057, S => n13671, Z => n14109
                           );
   U15882 : NAND2_X1 port map( A1 => n14239, A2 => n15423, ZN => n14113);
   U15883 : MUX2_X1 port map( A => n14113, B => n14240, S => n14149, Z => 
                           n14118);
   U15884 : INV_X1 port map( A => n14242, ZN => n14116);
   U15885 : NOR2_X1 port map( A1 => n14114, A2 => n15423, ZN => n14115);
   U15886 : AOI21_X1 port map( B1 => n14116, B2 => n19907, A => n14115, ZN => 
                           n14117);
   U15887 : NAND2_X1 port map( A1 => n14232, A2 => n14381, ZN => n14699);
   U15888 : OAI211_X1 port map( C1 => n19503, C2 => n14381, A => n14703, B => 
                           n14229, ZN => n14121);
   U15889 : NAND2_X1 port map( A1 => n16126, A2 => n15608, ZN => n14131);
   U15890 : NAND2_X1 port map( A1 => n14691, A2 => n14385, ZN => n14126);
   U15891 : INV_X1 port map( A => n14126, ZN => n14124);
   U15892 : NAND2_X1 port map( A1 => n14124, A2 => n19921, ZN => n14130);
   U15893 : INV_X1 port map( A => n14385, ZN => n14689);
   U15894 : NAND2_X1 port map( A1 => n14689, A2 => n19895, ZN => n14125);
   U15895 : NAND3_X1 port map( A1 => n14693, A2 => n20466, A3 => n200, ZN => 
                           n14128);
   U15896 : NAND3_X1 port map( A1 => n14726, A2 => n14134, A3 => n14133, ZN => 
                           n14136);
   U15897 : NAND3_X1 port map( A1 => n20376, A2 => n14728, A3 => n14724, ZN => 
                           n14135);
   U15898 : NAND2_X1 port map( A1 => n15608, A2 => n16129, ZN => n15734);
   U15899 : AOI21_X1 port map( B1 => n16126, B2 => n15734, A => n3431, ZN => 
                           n14138);
   U15900 : OAI21_X1 port map( B1 => n19488, B2 => n14611, A => n14143, ZN => 
                           n14145);
   U15901 : INV_X1 port map( A => n14207, ZN => n14144);
   U15902 : AND2_X1 port map( A1 => n19875, A2 => n14624, ZN => n15320);
   U15903 : NAND2_X1 port map( A1 => n15320, A2 => n14623, ZN => n14147);
   U15904 : NAND2_X1 port map( A1 => n14148, A2 => n19907, ZN => n14400);
   U15905 : NAND3_X1 port map( A1 => n14237, A2 => n14239, A3 => n14238, ZN => 
                           n14151);
   U15906 : INV_X1 port map( A => n3822, ZN => n15562);
   U15907 : NAND2_X1 port map( A1 => n14598, A2 => n14395, ZN => n14155);
   U15908 : MUX2_X1 port map( A => n14250, B => n14599, S => n1262, Z => n14157
                           );
   U15909 : NAND2_X1 port map( A1 => n14157, A2 => n20377, ZN => n14158);
   U15910 : INV_X1 port map( A => n15509, ZN => n15560);
   U15911 : NOR2_X1 port map( A1 => n15560, A2 => n15558, ZN => n14160);
   U15912 : INV_X1 port map( A => n15510, ZN => n15212);
   U15913 : INV_X1 port map( A => n15558, ZN => n15513);
   U15914 : AOI22_X1 port map( A1 => n14159, A2 => n14160, B1 => n15212, B2 => 
                           n15513, ZN => n14161);
   U15915 : OAI21_X1 port map( B1 => n20435, B2 => n15559, A => n14161, ZN => 
                           n16936);
   U15916 : INV_X1 port map( A => n2032, ZN => n18294);
   U15917 : XNOR2_X1 port map( A => n16936, B => n18294, ZN => n14162);
   U15918 : XNOR2_X1 port map( A => n14163, B => n14162, ZN => n14164);
   U15919 : AOI21_X1 port map( B1 => n16634, B2 => n20271, A => n16170, ZN => 
                           n14848);
   U15920 : MUX2_X1 port map( A => n19727, B => n1936, S => n20453, Z => n14166
                           );
   U15921 : NOR2_X1 port map( A1 => n19728, A2 => n14490, ZN => n14165);
   U15922 : NOR2_X1 port map( A1 => n14434, A2 => n14480, ZN => n14174);
   U15923 : AND2_X1 port map( A1 => n14482, A2 => n14171, ZN => n14303);
   U15924 : NAND2_X1 port map( A1 => n14303, A2 => n14172, ZN => n14173);
   U15925 : INV_X1 port map( A => n15309, ZN => n14886);
   U15926 : AND2_X1 port map( A1 => n15396, A2 => n14177, ZN => n14190);
   U15927 : NOR2_X1 port map( A1 => n14448, A2 => n14180, ZN => n14178);
   U15928 : MUX2_X1 port map( A => n14179, B => n14178, S => n1364, Z => n14183
                           );
   U15929 : MUX2_X1 port map( A => n14448, B => n14447, S => n14180, Z => 
                           n14181);
   U15931 : OAI21_X1 port map( B1 => n14519, B2 => n14514, A => n15119, ZN => 
                           n14184);
   U15932 : OAI21_X1 port map( B1 => n15311, B2 => n14188, A => n14187, ZN => 
                           n14189);
   U15933 : AOI21_X2 port map( B1 => n14190, B2 => n15311, A => n14189, ZN => 
                           n17338);
   U15934 : AOI21_X1 port map( B1 => n19875, B2 => n14620, A => n15313, ZN => 
                           n14191);
   U15935 : OAI21_X1 port map( B1 => n14192, B2 => n19875, A => n14191, ZN => 
                           n14194);
   U15936 : NAND3_X1 port map( A1 => n14192, A2 => n15313, A3 => n14623, ZN => 
                           n14193);
   U15937 : INV_X1 port map( A => n14196, ZN => n14198);
   U15938 : NOR2_X1 port map( A1 => n14813, A2 => n14810, ZN => n14197);
   U15939 : AOI22_X1 port map( A1 => n14599, A2 => n20513, B1 => n14601, B2 => 
                           n20181, ZN => n14201);
   U15940 : NAND2_X1 port map( A1 => n19488, A2 => n14611, ZN => n14204);
   U15941 : MUX2_X1 port map( A => n14204, B => n14609, S => n13907, Z => 
                           n14210);
   U15942 : NAND2_X1 port map( A1 => n19906, A2 => n13908, ZN => n14608);
   U15943 : INV_X1 port map( A => n14608, ZN => n14209);
   U15944 : OAI211_X1 port map( C1 => n20500, C2 => n3497, A => n14796, B => 
                           n1938, ZN => n14212);
   U15945 : NOR2_X1 port map( A1 => n15070, A2 => n15618, ZN => n15408);
   U15946 : INV_X1 port map( A => n15618, ZN => n14214);
   U15948 : MUX2_X1 port map( A => n14216, B => n14782, S => n14775, Z => 
                           n14219);
   U15949 : NAND3_X1 port map( A1 => n14057, A2 => n14782, A3 => n14778, ZN => 
                           n14218);
   U15950 : INV_X1 port map( A => n15405, ZN => n15544);
   U15951 : INV_X1 port map( A => n15070, ZN => n15620);
   U15952 : INV_X1 port map( A => n15071, ZN => n15406);
   U15953 : NAND3_X1 port map( A1 => n15544, A2 => n15620, A3 => n15406, ZN => 
                           n14220);
   U15954 : OAI211_X1 port map( C1 => n15619, C2 => n15616, A => n14221, B => 
                           n14220, ZN => n16954);
   U15955 : XNOR2_X1 port map( A => n16954, B => n17338, ZN => n16584);
   U15956 : OAI21_X1 port map( B1 => n20376, B2 => n14730, A => n236, ZN => 
                           n14222);
   U15957 : NAND2_X1 port map( A1 => n14222, A2 => n14731, ZN => n14226);
   U15959 : NAND2_X1 port map( A1 => n14594, A2 => n2924, ZN => n14233);
   U15960 : MUX2_X1 port map( A => n14234, B => n14233, S => n19761, Z => 
                           n14235);
   U15961 : INV_X1 port map( A => n15430, ZN => n15919);
   U15962 : OAI21_X1 port map( B1 => n14242, B2 => n19908, A => n14241, ZN => 
                           n15426);
   U15963 : MUX2_X1 port map( A => n14718, B => n3057, S => n14717, Z => n14247
                           );
   U15964 : NAND2_X1 port map( A1 => n3057, A2 => n14717, ZN => n14244);
   U15965 : MUX2_X1 port map( A => n14245, B => n14244, S => n14715, Z => 
                           n14246);
   U15966 : NAND2_X1 port map( A1 => n15921, A2 => n15422, ZN => n15920);
   U15967 : INV_X1 port map( A => n15422, ZN => n15420);
   U15968 : NAND2_X1 port map( A1 => n14248, A2 => n14599, ZN => n14255);
   U15969 : INV_X1 port map( A => n14601, ZN => n14251);
   U15970 : NAND3_X1 port map( A1 => n20513, A2 => n14251, A3 => n19918, ZN => 
                           n14253);
   U15971 : NAND2_X1 port map( A1 => n14599, A2 => n20181, ZN => n14252);
   U15973 : OAI21_X1 port map( B1 => n15421, B2 => n15920, A => n14257, ZN => 
                           n14258);
   U15974 : NAND2_X1 port map( A1 => n14674, A2 => n19652, ZN => n14264);
   U15975 : INV_X1 port map( A => n14575, ZN => n14569);
   U15976 : NAND2_X1 port map( A1 => n14569, A2 => n14269, ZN => n14737);
   U15977 : NAND3_X1 port map( A1 => n14270, A2 => n14571, A3 => n14737, ZN => 
                           n14271);
   U15978 : NAND2_X1 port map( A1 => n14705, A2 => n14275, ZN => n14274);
   U15979 : AOI21_X1 port map( B1 => n14274, B2 => n14273, A => n14566, ZN => 
                           n14278);
   U15980 : NAND2_X1 port map( A1 => n919, A2 => n14276, ZN => n14277);
   U15981 : AND2_X1 port map( A1 => n15400, A2 => n15536, ZN => n14296);
   U15983 : MUX2_X1 port map( A => n14283, B => n14282, S => n14550, Z => 
                           n14909);
   U15984 : NAND2_X1 port map( A1 => n14284, A2 => n20120, ZN => n14908);
   U15985 : NOR2_X1 port map( A1 => n20471, A2 => n14656, ZN => n14287);
   U15986 : INV_X1 port map( A => n14288, ZN => n14660);
   U15987 : OAI21_X1 port map( B1 => n14289, B2 => n20266, A => n14547, ZN => 
                           n14290);
   U15988 : NOR2_X1 port map( A1 => n14660, A2 => n14290, ZN => n14291);
   U15989 : NAND3_X1 port map( A1 => n14688, A2 => n19895, A3 => n14695, ZN => 
                           n14295);
   U15990 : AND2_X1 port map( A1 => n19921, A2 => n14127, ZN => n14384);
   U15991 : OAI21_X1 port map( B1 => n14384, B2 => n14385, A => n14691, ZN => 
                           n14294);
   U15992 : OAI211_X1 port map( C1 => n14696, C2 => n20466, A => n14295, B => 
                           n14294, ZN => n15401);
   U15993 : INV_X1 port map( A => n15401, ZN => n15538);
   U15994 : NAND3_X1 port map( A1 => n15898, A2 => n15402, A3 => n15538, ZN => 
                           n14298);
   U15995 : NAND2_X1 port map( A1 => n19722, A2 => n14296, ZN => n14297);
   U15996 : XNOR2_X1 port map( A => n16755, B => n16836, ZN => n17267);
   U15997 : XNOR2_X1 port map( A => n16584, B => n17267, ZN => n14376);
   U15998 : NOR2_X1 port map( A1 => n14512, A2 => n14509, ZN => n14639);
   U15999 : NAND2_X1 port map( A1 => n14642, A2 => n14641, ZN => n14299);
   U16000 : NOR2_X1 port map( A1 => n14639, A2 => n14299, ZN => n14300);
   U16001 : NOR2_X1 port map( A1 => n14309, A2 => n14308, ZN => n14312);
   U16002 : MUX2_X1 port map( A => n14648, B => n14651, S => n20443, Z => 
                           n14311);
   U16005 : OAI21_X1 port map( B1 => n14314, B2 => n14667, A => n14313, ZN => 
                           n14318);
   U16006 : AOI21_X1 port map( B1 => n14316, B2 => n14315, A => n14662, ZN => 
                           n14317);
   U16007 : INV_X1 port map( A => n14903, ZN => n15410);
   U16008 : MUX2_X1 port map( A => n14520, B => n15121, S => n15119, Z => 
                           n14323);
   U16009 : NAND2_X1 port map( A1 => n15120, A2 => n14520, ZN => n14319);
   U16010 : OAI22_X1 port map( A1 => n14321, A2 => n14320, B1 => n14319, B2 => 
                           n14514, ZN => n14322);
   U16011 : XNOR2_X1 port map( A => n16373, B => n18278, ZN => n14374);
   U16012 : MUX2_X1 port map( A => n15469, B => n15336, S => n15465, Z => 
                           n14324);
   U16013 : NAND2_X1 port map( A1 => n14324, A2 => n15337, ZN => n14333);
   U16015 : MUX2_X1 port map( A => n14329, B => n14328, S => n19693, Z => 
                           n14331);
   U16016 : INV_X1 port map( A => n15470, ZN => n15343);
   U16017 : NOR2_X1 port map( A1 => n19583, A2 => n15339, ZN => n14332);
   U16018 : NAND2_X1 port map( A1 => n14336, A2 => n14335, ZN => n14337);
   U16019 : NAND2_X1 port map( A1 => n14338, A2 => n14342, ZN => n14340);
   U16020 : MUX2_X1 port map( A => n14788, B => n14344, S => n14789, Z => 
                           n14345);
   U16021 : MUX2_X1 port map( A => n3223, B => n19496, S => n14827, Z => n14349
                           );
   U16022 : NOR2_X1 port map( A1 => n19859, A2 => n19986, ZN => n14348);
   U16023 : NOR2_X1 port map( A1 => n235, A2 => n14818, ZN => n14351);
   U16024 : AOI22_X1 port map( A1 => n14353, A2 => n20330, B1 => n14352, B2 => 
                           n14351, ZN => n14354);
   U16025 : OAI21_X1 port map( B1 => n2039, B2 => n14357, A => n14356, ZN => 
                           n14423);
   U16026 : INV_X1 port map( A => n14423, ZN => n14362);
   U16027 : INV_X1 port map( A => n14358, ZN => n14361);
   U16028 : OAI211_X1 port map( C1 => n14422, C2 => n14359, A => n14419, B => 
                           n19939, ZN => n14360);
   U16029 : OAI21_X2 port map( B1 => n14362, B2 => n14361, A => n14360, ZN => 
                           n15907);
   U16030 : INV_X1 port map( A => n14363, ZN => n14365);
   U16032 : NAND2_X1 port map( A1 => n19531, A2 => n14462, ZN => n14466);
   U16033 : NAND3_X1 port map( A1 => n19531, A2 => n14468, A3 => n14369, ZN => 
                           n14367);
   U16034 : AND2_X1 port map( A1 => n14466, A2 => n14367, ZN => n14368);
   U16035 : NOR2_X1 port map( A1 => n15909, A2 => n15905, ZN => n15077);
   U16036 : XNOR2_X1 port map( A => n16300, B => n16406, ZN => n14373);
   U16037 : XNOR2_X1 port map( A => n14374, B => n14373, ZN => n14375);
   U16038 : NAND2_X1 port map( A1 => n17511, A2 => n20271, ZN => n17509);
   U16039 : INV_X1 port map( A => n17509, ZN => n16172);
   U16040 : INV_X1 port map( A => n15843, ZN => n15267);
   U16041 : NOR2_X1 port map( A1 => n15636, A2 => n15267, ZN => n14377);
   U16042 : MUX2_X1 port map( A => n14700, B => n14703, S => n20204, Z => 
                           n14383);
   U16043 : NAND2_X1 port map( A1 => n14380, A2 => n14379, ZN => n14382);
   U16044 : INV_X1 port map( A => n15838, ZN => n15100);
   U16045 : NAND2_X1 port map( A1 => n14693, A2 => n14384, ZN => n14386);
   U16046 : NAND2_X1 port map( A1 => n19862, A2 => n14723, ZN => n14392);
   U16047 : MUX2_X1 port map( A => n19862, B => n14723, S => n14718, Z => 
                           n14390);
   U16048 : MUX2_X1 port map( A => n14390, B => n14389, S => n19843, Z => 
                           n14391);
   U16049 : OAI21_X1 port map( B1 => n2926, B2 => n14394, A => n19731, ZN => 
                           n14399);
   U16050 : NAND2_X1 port map( A1 => n14403, A2 => n15423, ZN => n14404);
   U16051 : AOI21_X1 port map( B1 => n14406, B2 => n14405, A => n14404, ZN => 
                           n14407);
   U16052 : NOR2_X1 port map( A1 => n15627, A2 => n15628, ZN => n14415);
   U16053 : NOR2_X1 port map( A1 => n14408, A2 => n14729, ZN => n14409);
   U16054 : NAND2_X1 port map( A1 => n14409, A2 => n14726, ZN => n15002);
   U16055 : NAND2_X1 port map( A1 => n14410, A2 => n14724, ZN => n14411);
   U16056 : NAND2_X1 port map( A1 => n14731, A2 => n14411, ZN => n14413);
   U16057 : MUX2_X1 port map( A => n14728, B => n14413, S => n14412, Z => 
                           n15003);
   U16058 : AOI21_X1 port map( B1 => n15002, B2 => n15003, A => n15625, ZN => 
                           n14414);
   U16059 : MUX2_X1 port map( A => n14415, B => n14414, S => n15838, Z => 
                           n14416);
   U16060 : AOI21_X1 port map( B1 => n14417, B2 => n15627, A => n14416, ZN => 
                           n17261);
   U16061 : XNOR2_X1 port map( A => n17261, B => n17438, ZN => n16514);
   U16062 : OAI21_X1 port map( B1 => n19939, B2 => n14419, A => n14418, ZN => 
                           n14421);
   U16063 : NAND2_X1 port map( A1 => n14424, A2 => n3156, ZN => n14430);
   U16064 : NOR2_X1 port map( A1 => n14426, A2 => n14425, ZN => n14492);
   U16065 : INV_X1 port map( A => n14492, ZN => n14429);
   U16066 : NAND2_X1 port map( A1 => n14433, A2 => n14480, ZN => n14438);
   U16067 : INV_X1 port map( A => n14434, ZN => n14436);
   U16068 : NOR2_X1 port map( A1 => n14436, A2 => n14435, ZN => n14437);
   U16069 : INV_X1 port map( A => n15297, ZN => n14446);
   U16070 : MUX2_X1 port map( A => n14442, B => n12919, S => n14441, Z => 
                           n14444);
   U16071 : NOR2_X1 port map( A1 => n14444, A2 => n14443, ZN => n14445);
   U16072 : AOI21_X1 port map( B1 => n15296, B2 => n14446, A => n15294, ZN => 
                           n14460);
   U16073 : NOR2_X1 port map( A1 => n14452, A2 => n14451, ZN => n14457);
   U16074 : NOR2_X1 port map( A1 => n14454, A2 => n14453, ZN => n14456);
   U16075 : MUX2_X1 port map( A => n14457, B => n14456, S => n1364, Z => n14458
                           );
   U16076 : MUX2_X1 port map( A => n15111, B => n14460, S => n14770, Z => 
                           n14473);
   U16077 : NAND2_X1 port map( A1 => n15294, A2 => n14461, ZN => n15293);
   U16078 : INV_X1 port map( A => n19819, ZN => n14464);
   U16079 : AOI21_X1 port map( B1 => n14465, B2 => n14464, A => n3252, ZN => 
                           n14467);
   U16080 : MUX2_X1 port map( A => n14468, B => n14467, S => n14466, Z => 
                           n14471);
   U16081 : NOR3_X1 port map( A1 => n3299, A2 => n14469, A3 => n14468, ZN => 
                           n14470);
   U16083 : NOR2_X1 port map( A1 => n15293, A2 => n15110, ZN => n14472);
   U16084 : NOR2_X2 port map( A1 => n14473, A2 => n14472, ZN => n16607);
   U16086 : NAND2_X1 port map( A1 => n15909, A2 => n15905, ZN => n14475);
   U16087 : NAND2_X1 port map( A1 => n15008, A2 => n15907, ZN => n14474);
   U16088 : NAND3_X1 port map( A1 => n14475, A2 => n2578, A3 => n14474, ZN => 
                           n14478);
   U16089 : INV_X1 port map( A => n14475, ZN => n14476);
   U16090 : NAND2_X1 port map( A1 => n14476, A2 => n15906, ZN => n14477);
   U16091 : OAI211_X1 port map( C1 => n2578, C2 => n14479, A => n14478, B => 
                           n14477, ZN => n16293);
   U16092 : XNOR2_X1 port map( A => n16607, B => n16293, ZN => n16175);
   U16093 : XNOR2_X1 port map( A => n16514, B => n16175, ZN => n14634);
   U16094 : NAND2_X1 port map( A1 => n14482, A2 => n14480, ZN => n14489);
   U16097 : INV_X1 port map( A => n15132, ZN => n14838);
   U16098 : NOR2_X1 port map( A1 => n14747, A2 => n14490, ZN => n14491);
   U16099 : OR2_X2 port map( A1 => n14496, A2 => n14495, ZN => n15282);
   U16100 : MUX2_X1 port map( A => n14499, B => n14498, S => n14497, Z => 
                           n14505);
   U16104 : NOR2_X1 port map( A1 => n15282, A2 => n15284, ZN => n15286);
   U16105 : INV_X1 port map( A => n15286, ZN => n14534);
   U16106 : NAND2_X1 port map( A1 => n13983, A2 => n14641, ZN => n14507);
   U16107 : AOI22_X1 port map( A1 => n14635, A2 => n14512, B1 => n19703, B2 => 
                           n14640, ZN => n14511);
   U16108 : INV_X1 port map( A => n15130, ZN => n14529);
   U16109 : INV_X1 port map( A => n14514, ZN => n14515);
   U16111 : NOR2_X1 port map( A1 => n951, A2 => n14522, ZN => n14523);
   U16112 : NAND3_X1 port map( A1 => n14525, A2 => n14648, A3 => n14524, ZN => 
                           n14526);
   U16113 : NAND2_X1 port map( A1 => n14652, A2 => n14526, ZN => n14527);
   U16114 : NAND2_X1 port map( A1 => n14529, A2 => n15127, ZN => n14530);
   U16115 : NAND2_X1 port map( A1 => n15281, A2 => n14530, ZN => n14531);
   U16116 : NAND2_X1 port map( A1 => n14531, A2 => n19848, ZN => n14533);
   U16117 : NAND3_X1 port map( A1 => n15282, A2 => n15018, A3 => n20474, ZN => 
                           n14532);
   U16118 : NAND2_X1 port map( A1 => n14673, A2 => n14539, ZN => n14546);
   U16119 : NAND2_X1 port map( A1 => n20424, A2 => n19652, ZN => n14675);
   U16120 : NAND2_X1 port map( A1 => n14544, A2 => n13981, ZN => n14545);
   U16121 : INV_X1 port map( A => n15645, ZN => n15831);
   U16124 : INV_X1 port map( A => n15256, ZN => n15643);
   U16125 : MUX2_X1 port map( A => n14552, B => n14551, S => n14279, Z => 
                           n14561);
   U16126 : NOR2_X1 port map( A1 => n14554, A2 => n14553, ZN => n14559);
   U16127 : NOR2_X1 port map( A1 => n14556, A2 => n14555, ZN => n14558);
   U16128 : MUX2_X1 port map( A => n14559, B => n14558, S => n14557, Z => 
                           n14560);
   U16129 : INV_X1 port map( A => n15644, ZN => n15829);
   U16130 : MUX2_X1 port map( A => n20498, B => n14705, S => n14562, Z => 
                           n14567);
   U16131 : MUX2_X1 port map( A => n14564, B => n14563, S => n14704, Z => 
                           n14565);
   U16132 : OAI21_X1 port map( B1 => n14567, B2 => n14566, A => n14565, ZN => 
                           n15096);
   U16133 : NAND2_X1 port map( A1 => n15829, A2 => n19891, ZN => n15649);
   U16135 : NAND2_X1 port map( A1 => n14569, A2 => n14736, ZN => n14573);
   U16136 : NAND2_X1 port map( A1 => n14571, A2 => n14570, ZN => n14572);
   U16138 : AND2_X1 port map( A1 => n15096, A2 => n15644, ZN => n15259);
   U16139 : INV_X1 port map( A => n15259, ZN => n14580);
   U16140 : AOI21_X1 port map( B1 => n14581, B2 => n14580, A => n15256, ZN => 
                           n14582);
   U16141 : XNOR2_X1 port map( A => n16750, B => n19704, ZN => n16392);
   U16142 : NOR2_X1 port map( A1 => n14796, A2 => n1351, ZN => n14585);
   U16143 : AOI22_X1 port map( A1 => n14585, A2 => n3439, B1 => n1351, B2 => 
                           n14799, ZN => n14586);
   U16144 : NAND2_X1 port map( A1 => n14587, A2 => n14199, ZN => n14592);
   U16145 : INV_X1 port map( A => n14807, ZN => n14589);
   U16146 : NOR2_X1 port map( A1 => n15270, A2 => n15601, ZN => n14618);
   U16147 : NAND3_X1 port map( A1 => n20377, A2 => n2682, A3 => n14601, ZN => 
                           n14607);
   U16148 : INV_X1 port map( A => n14603, ZN => n14604);
   U16149 : NAND3_X1 port map( A1 => n20513, A2 => n1262, A3 => n14604, ZN => 
                           n14606);
   U16150 : INV_X1 port map( A => n15274, ZN => n15114);
   U16151 : NOR2_X1 port map( A1 => n15275, A2 => n15114, ZN => n14617);
   U16152 : AOI21_X1 port map( B1 => n14612, B2 => n13907, A => n14611, ZN => 
                           n14613);
   U16153 : NAND2_X1 port map( A1 => n14614, A2 => n14613, ZN => n14615);
   U16156 : NAND3_X1 port map( A1 => n954, A2 => n19875, A3 => n14623, ZN => 
                           n14622);
   U16157 : NAND3_X1 port map( A1 => n15314, A2 => n14620, A3 => n15313, ZN => 
                           n14621);
   U16159 : OAI211_X1 port map( C1 => n954, C2 => n14627, A => n14625, B => 
                           n14624, ZN => n14628);
   U16160 : NAND2_X1 port map( A1 => n15276, A2 => n15271, ZN => n14629);
   U16161 : INV_X1 port map( A => n15270, ZN => n15009);
   U16162 : AOI21_X1 port map( B1 => n15277, B2 => n14629, A => n15009, ZN => 
                           n14630);
   U16163 : NOR2_X2 port map( A1 => n14631, A2 => n14630, ZN => n16914);
   U16164 : INV_X1 port map( A => n649, ZN => n19152);
   U16165 : XNOR2_X1 port map( A => n16914, B => n19152, ZN => n14632);
   U16166 : XNOR2_X1 port map( A => n16392, B => n14632, ZN => n14633);
   U16167 : OR2_X1 port map( A1 => n14636, A2 => n14635, ZN => n14646);
   U16168 : NOR2_X1 port map( A1 => n14640, A2 => n14637, ZN => n14638);
   U16169 : NOR2_X1 port map( A1 => n14639, A2 => n14638, ZN => n14645);
   U16170 : MUX2_X1 port map( A => n14642, B => n14641, S => n14640, Z => 
                           n14643);
   U16171 : OAI22_X1 port map( A1 => n14651, A2 => n951, B1 => n14648, B2 => 
                           n20380, ZN => n14649);
   U16172 : AND2_X1 port map( A1 => n15573, A2 => n15577, ZN => n15793);
   U16173 : NOR2_X1 port map( A1 => n14653, A2 => n14656, ZN => n14655);
   U16174 : NAND3_X1 port map( A1 => n14655, A2 => n14654, A3 => n14659, ZN => 
                           n14661);
   U16175 : OAI21_X1 port map( B1 => n20266, B2 => n14656, A => n20471, ZN => 
                           n14658);
   U16176 : NOR2_X1 port map( A1 => n15793, A2 => n15574, ZN => n14687);
   U16177 : NOR2_X1 port map( A1 => n14663, A2 => n14662, ZN => n14665);
   U16178 : INV_X1 port map( A => n15573, ZN => n15791);
   U16179 : NOR2_X1 port map( A1 => n15791, A2 => n15577, ZN => n14685);
   U16180 : OR2_X1 port map( A1 => n14680, A2 => n20120, ZN => n14681);
   U16181 : NAND3_X1 port map( A1 => n14683, A2 => n14682, A3 => n14681, ZN => 
                           n15365);
   U16182 : INV_X1 port map( A => n15365, ZN => n15572);
   U16183 : NOR2_X1 port map( A1 => n15577, A2 => n15572, ZN => n14684);
   U16184 : AOI22_X1 port map( A1 => n15796, A2 => n14685, B1 => n14684, B2 => 
                           n860, ZN => n14686);
   U16186 : NAND3_X1 port map( A1 => n14689, A2 => n14688, A3 => n200, ZN => 
                           n14694);
   U16187 : NAND2_X1 port map( A1 => n14120, A2 => n2769, ZN => n14698);
   U16188 : NAND2_X1 port map( A1 => n14699, A2 => n14698, ZN => n14701);
   U16189 : NAND2_X1 port map( A1 => n14701, A2 => n14700, ZN => n14702);
   U16190 : OAI21_X1 port map( B1 => n14273, B2 => n14704, A => n919, ZN => 
                           n14713);
   U16191 : NOR2_X1 port map( A1 => n14705, A2 => n2282, ZN => n14712);
   U16192 : NAND2_X1 port map( A1 => n14708, A2 => n20498, ZN => n14711);
   U16193 : NAND2_X1 port map( A1 => n14273, A2 => n14709, ZN => n14710);
   U16194 : OAI211_X1 port map( C1 => n14713, C2 => n14712, A => n14711, B => 
                           n14710, ZN => n15801);
   U16195 : INV_X1 port map( A => n15801, ZN => n15042);
   U16196 : OAI21_X1 port map( B1 => n14716, B2 => n14715, A => n19862, ZN => 
                           n14720);
   U16197 : MUX2_X1 port map( A => n14720, B => n14719, S => n14718, Z => 
                           n14721);
   U16198 : MUX2_X1 port map( A => n14731, B => n14730, S => n14729, Z => 
                           n14733);
   U16199 : NOR2_X1 port map( A1 => n14733, A2 => n20376, ZN => n14734);
   U16200 : NAND2_X1 port map( A1 => n14737, A2 => n14736, ZN => n14739);
   U16202 : INV_X1 port map( A => n15802, ZN => n14742);
   U16204 : AND2_X1 port map( A1 => n15801, A2 => n15803, ZN => n15564);
   U16205 : INV_X1 port map( A => n15567, ZN => n15804);
   U16206 : AOI22_X1 port map( A1 => n15564, A2 => n942, B1 => n15804, B2 => 
                           n15801, ZN => n14744);
   U16207 : XNOR2_X1 port map( A => n17294, B => n16853, ZN => n16365);
   U16208 : NOR2_X1 port map( A1 => n14747, A2 => n19727, ZN => n14748);
   U16209 : NOR2_X1 port map( A1 => n14749, A2 => n14748, ZN => n14751);
   U16210 : MUX2_X1 port map( A => n14751, B => n14750, S => n1936, Z => n14752
                           );
   U16211 : NAND2_X1 port map( A1 => n15189, A2 => n14935, ZN => n14764);
   U16212 : INV_X1 port map( A => n14754, ZN => n14761);
   U16213 : INV_X1 port map( A => n14755, ZN => n14760);
   U16214 : INV_X1 port map( A => n14756, ZN => n14759);
   U16215 : INV_X1 port map( A => n14757, ZN => n14758);
   U16216 : NAND4_X1 port map( A1 => n14761, A2 => n14760, A3 => n14759, A4 => 
                           n14758, ZN => n14762);
   U16217 : AOI22_X1 port map( A1 => n15504, A2 => n15506, B1 => n2288, B2 => 
                           n14762, ZN => n14763);
   U16218 : AOI22_X2 port map( A1 => n14763, A2 => n14764, B1 => n15506, B2 => 
                           n15822, ZN => n16945);
   U16219 : INV_X1 port map( A => n15559, ZN => n14966);
   U16220 : OAI21_X1 port map( B1 => n15511, B2 => n15510, A => n14159, ZN => 
                           n14766);
   U16221 : OAI211_X1 port map( C1 => n14966, C2 => n14964, A => n14766, B => 
                           n14765, ZN => n17300);
   U16222 : INV_X1 port map( A => n17300, ZN => n14767);
   U16223 : XNOR2_X1 port map( A => n16945, B => n14767, ZN => n16527);
   U16224 : XNOR2_X1 port map( A => n16365, B => n16527, ZN => n14844);
   U16225 : NOR2_X1 port map( A1 => n15110, A2 => n15295, ZN => n14769);
   U16226 : AOI21_X1 port map( B1 => n14771, B2 => n14770, A => n14769, ZN => 
                           n14774);
   U16227 : NAND2_X1 port map( A1 => n15295, A2 => n15111, ZN => n14772);
   U16228 : NOR2_X1 port map( A1 => n15110, A2 => n14772, ZN => n14773);
   U16229 : NAND3_X1 port map( A1 => n877, A2 => n20518, A3 => n14775, ZN => 
                           n14776);
   U16230 : OAI21_X1 port map( B1 => n14852, B2 => n20408, A => n14776, ZN => 
                           n14786);
   U16231 : NOR2_X1 port map( A1 => n877, A2 => n14778, ZN => n14784);
   U16232 : NOR2_X1 port map( A1 => n14781, A2 => n20454, ZN => n14783);
   U16233 : MUX2_X1 port map( A => n14784, B => n14783, S => n14782, Z => 
                           n14785);
   U16234 : MUX2_X1 port map( A => n14103, B => n14787, S => n14790, Z => 
                           n14794);
   U16235 : MUX2_X1 port map( A => n14791, B => n14790, S => n14789, Z => 
                           n14793);
   U16236 : NAND2_X1 port map( A1 => n14796, A2 => n13891, ZN => n14798);
   U16237 : AOI21_X1 port map( B1 => n14798, B2 => n14797, A => n14800, ZN => 
                           n14805);
   U16238 : NAND3_X1 port map( A1 => n1351, A2 => n3497, A3 => n14799, ZN => 
                           n14803);
   U16239 : NAND2_X1 port map( A1 => n14803, A2 => n14802, ZN => n14804);
   U16240 : MUX2_X1 port map( A => n15582, B => n3534, S => n15812, Z => n14836
                           );
   U16241 : NOR2_X1 port map( A1 => n14807, A2 => n14806, ZN => n14808);
   U16242 : AOI22_X1 port map( A1 => n14812, A2 => n14809, B1 => n14808, B2 => 
                           n14199, ZN => n14816);
   U16243 : OAI21_X1 port map( B1 => n239, B2 => n14814, A => n14813, ZN => 
                           n14815);
   U16245 : NAND2_X1 port map( A1 => n14820, A2 => n12931, ZN => n14822);
   U16247 : INV_X1 port map( A => n15583, ZN => n15814);
   U16248 : NOR2_X1 port map( A1 => n15814, A2 => n15582, ZN => n15354);
   U16250 : OAI211_X1 port map( C1 => n14828, C2 => n3223, A => n14827, B => 
                           n14826, ZN => n14832);
   U16251 : NOR2_X1 port map( A1 => n15354, A2 => n14834, ZN => n14835);
   U16252 : XNOR2_X1 port map( A => n16964, B => n17295, ZN => n14842);
   U16253 : NAND2_X1 port map( A1 => n15132, A2 => n15282, ZN => n14837);
   U16254 : MUX2_X1 port map( A => n15017, B => n20474, S => n15018, Z => 
                           n14839);
   U16255 : XNOR2_X1 port map( A => n16614, B => n18988, ZN => n14841);
   U16256 : XNOR2_X1 port map( A => n14842, B => n14841, ZN => n14843);
   U16257 : XNOR2_X1 port map( A => n14844, B => n14843, ZN => n17225);
   U16258 : INV_X1 port map( A => n17225, ZN => n14845);
   U16259 : NAND2_X1 port map( A1 => n14845, A2 => n19700, ZN => n14846);
   U16261 : INV_X1 port map( A => n15769, ZN => n15475);
   U16262 : INV_X1 port map( A => n14850, ZN => n14854);
   U16263 : INV_X1 port map( A => n14851, ZN => n14853);
   U16264 : NAND3_X1 port map( A1 => n14854, A2 => n14853, A3 => n14852, ZN => 
                           n14855);
   U16265 : NOR2_X1 port map( A1 => n14856, A2 => n14855, ZN => n14857);
   U16266 : NOR2_X2 port map( A1 => n14859, A2 => n14858, ZN => n16981);
   U16267 : INV_X1 port map( A => n15349, ZN => n15348);
   U16268 : NOR2_X1 port map( A1 => n20173, A2 => n15348, ZN => n14861);
   U16270 : XNOR2_X1 port map( A => n16981, B => n19927, ZN => n16506);
   U16271 : INV_X1 port map( A => n15673, ZN => n15775);
   U16273 : NAND2_X1 port map( A1 => n15672, A2 => n15665, ZN => n14864);
   U16274 : NAND2_X1 port map( A1 => n13414, A2 => n20151, ZN => n14863);
   U16275 : MUX2_X1 port map( A => n14864, B => n14863, S => n234, Z => n14865)
                           ;
   U16276 : INV_X1 port map( A => n14866, ZN => n15783);
   U16279 : NAND3_X1 port map( A1 => n15685, A2 => n15683, A3 => n15684, ZN => 
                           n14869);
   U16280 : NAND3_X1 port map( A1 => n15686, A2 => n19977, A3 => n20362, ZN => 
                           n14868);
   U16281 : XNOR2_X1 port map( A => n17339, B => n1054, ZN => n17036);
   U16282 : XNOR2_X1 port map( A => n16506, B => n17036, ZN => n14885);
   U16283 : NOR2_X1 port map( A1 => n15380, A2 => n15166, ZN => n14871);
   U16284 : NOR2_X1 port map( A1 => n14872, A2 => n14871, ZN => n14873);
   U16285 : NOR3_X1 port map( A1 => n15380, A2 => n15379, A3 => n20103, ZN => 
                           n14876);
   U16286 : NOR2_X1 port map( A1 => n15682, A2 => n15445, ZN => n14880);
   U16287 : NOR3_X1 port map( A1 => n15676, A2 => n15679, A3 => n15442, ZN => 
                           n14879);
   U16288 : NOR2_X1 port map( A1 => n14880, A2 => n14879, ZN => n14881);
   U16289 : XNOR2_X1 port map( A => n897, B => n17340, ZN => n14883);
   U16290 : XNOR2_X1 port map( A => n16300, B => n19140, ZN => n14882);
   U16291 : XNOR2_X1 port map( A => n14883, B => n14882, ZN => n14884);
   U16293 : NOR2_X1 port map( A1 => n15311, A2 => n15395, ZN => n14889);
   U16294 : NAND2_X1 port map( A1 => n15059, A2 => n15308, ZN => n14990);
   U16295 : OAI21_X1 port map( B1 => n14886, B2 => n15308, A => n14990, ZN => 
                           n14887);
   U16296 : NOR2_X1 port map( A1 => n15546, A2 => n15619, ZN => n14890);
   U16297 : NAND2_X1 port map( A1 => n14890, A2 => n15406, ZN => n14894);
   U16298 : NOR2_X1 port map( A1 => n15405, A2 => n15618, ZN => n14891);
   U16299 : OAI21_X1 port map( B1 => n15073, B2 => n14891, A => n15546, ZN => 
                           n14893);
   U16300 : NAND3_X1 port map( A1 => n14894, A2 => n14893, A3 => n14892, ZN => 
                           n16999);
   U16301 : INV_X1 port map( A => n16999, ZN => n16510);
   U16302 : XNOR2_X1 port map( A => n16999, B => n14895, ZN => n15953);
   U16303 : NAND2_X1 port map( A1 => n15465, A2 => n14896, ZN => n14897);
   U16304 : NAND2_X1 port map( A1 => n15082, A2 => n3817, ZN => n14898);
   U16305 : INV_X1 port map( A => n19467, ZN => n14901);
   U16306 : INV_X1 port map( A => n14902, ZN => n15550);
   U16307 : NAND2_X1 port map( A1 => n15550, A2 => n14903, ZN => n14904);
   U16308 : AND3_X1 port map( A1 => n14905, A2 => n14978, A3 => n14904, ZN => 
                           n14906);
   U16309 : NOR2_X2 port map( A1 => n14907, A2 => n14906, ZN => n17260);
   U16310 : INV_X1 port map( A => n15400, ZN => n15537);
   U16311 : OAI21_X1 port map( B1 => n15401, B2 => n15536, A => n15537, ZN => 
                           n14913);
   U16314 : NAND2_X1 port map( A1 => n14909, A2 => n14908, ZN => n15892);
   U16317 : XNOR2_X1 port map( A => n17378, B => n17260, ZN => n14914);
   U16319 : INV_X1 port map( A => n15859, ZN => n14918);
   U16320 : INV_X1 port map( A => n15720, ZN => n15862);
   U16321 : OAI21_X1 port map( B1 => n15866, B2 => n15862, A => n15863, ZN => 
                           n14917);
   U16322 : MUX2_X1 port map( A => n15864, B => n15861, S => n15720, Z => 
                           n14916);
   U16323 : XNOR2_X1 port map( A => n16420, B => n17104, ZN => n14928);
   U16324 : NOR2_X1 port map( A1 => n15875, A2 => n15714, ZN => n15713);
   U16325 : INV_X1 port map( A => n15870, ZN => n15150);
   U16326 : MUX2_X1 port map( A => n15874, B => n15876, S => n20178, Z => 
                           n14920);
   U16327 : NOR2_X1 port map( A1 => n14920, A2 => n15148, ZN => n14921);
   U16328 : NOR2_X2 port map( A1 => n14922, A2 => n14921, ZN => n17012);
   U16329 : INV_X1 port map( A => n15335, ZN => n14923);
   U16330 : NAND2_X1 port map( A1 => n16009, A2 => n19739, ZN => n15880);
   U16331 : NAND3_X1 port map( A1 => n14923, A2 => n16015, A3 => n15880, ZN => 
                           n14926);
   U16332 : INV_X1 port map( A => n14924, ZN => n14925);
   U16333 : NAND2_X1 port map( A1 => n15885, A2 => n14925, ZN => n16017);
   U16334 : XNOR2_X1 port map( A => n17012, B => n14927, ZN => n16418);
   U16335 : XNOR2_X1 port map( A => n14928, B => n16418, ZN => n14943);
   U16337 : INV_X1 port map( A => n15496, ZN => n15191);
   U16338 : AND2_X1 port map( A1 => n15501, A2 => n15191, ZN => n14929);
   U16339 : OAI21_X1 port map( B1 => n14930, B2 => n14929, A => n15497, ZN => 
                           n14933);
   U16340 : INV_X1 port map( A => n15501, ZN => n14931);
   U16341 : NAND3_X1 port map( A1 => n14931, A2 => n19512, A3 => n15500, ZN => 
                           n14932);
   U16342 : MUX2_X1 port map( A => n15505, B => n15503, S => n15188, Z => 
                           n14936);
   U16343 : XNOR2_X1 port map( A => n16602, B => n16045, ZN => n16232);
   U16344 : NOR2_X1 port map( A1 => n20133, A2 => n15696, ZN => n14940);
   U16345 : NOR2_X1 port map( A1 => n20145, A2 => n15702, ZN => n14939);
   U16346 : XNOR2_X1 port map( A => n19836, B => n18768, ZN => n14941);
   U16347 : XNOR2_X1 port map( A => n16232, B => n14941, ZN => n14942);
   U16349 : MUX2_X1 port map( A => n17210, B => n20135, S => n20092, Z => 
                           n15027);
   U16352 : NAND2_X1 port map( A1 => n15297, A2 => n14461, ZN => n14945);
   U16353 : MUX2_X1 port map( A => n14946, B => n14945, S => n15296, Z => 
                           n14947);
   U16354 : XNOR2_X1 port map( A => n16329, B => n17733, ZN => n14957);
   U16355 : INV_X1 port map( A => n15574, ZN => n15794);
   U16356 : NAND2_X1 port map( A1 => n859, A2 => n15572, ZN => n14949);
   U16357 : NOR2_X1 port map( A1 => n15577, A2 => n15573, ZN => n14948);
   U16358 : NOR2_X1 port map( A1 => n14949, A2 => n14948, ZN => n14950);
   U16359 : NOR2_X2 port map( A1 => n14951, A2 => n14950, ZN => n17280);
   U16360 : INV_X1 port map( A => n17280, ZN => n14956);
   U16361 : INV_X1 port map( A => n14952, ZN => n15371);
   U16362 : AOI22_X1 port map( A1 => n20183, A2 => n15371, B1 => n15370, B2 => 
                           n15566, ZN => n15043);
   U16363 : NAND2_X1 port map( A1 => n15803, A2 => n15042, ZN => n14953);
   U16364 : NAND2_X1 port map( A1 => n15808, A2 => n14953, ZN => n14955);
   U16367 : XNOR2_X1 port map( A => n17026, B => n14957, ZN => n14971);
   U16368 : NOR2_X1 port map( A1 => n15132, A2 => n15282, ZN => n15287);
   U16369 : INV_X1 port map( A => n15018, ZN => n15285);
   U16370 : NAND2_X1 port map( A1 => n15285, A2 => n15127, ZN => n14961);
   U16371 : INV_X1 port map( A => n15282, ZN => n14959);
   U16372 : NAND2_X1 port map( A1 => n15130, A2 => n15017, ZN => n14958);
   U16374 : INV_X1 port map( A => n16927, ZN => n14963);
   U16375 : NOR2_X1 port map( A1 => n15814, A2 => n233, ZN => n14962);
   U16376 : XNOR2_X1 port map( A => n14963, B => n16969, ZN => n16522);
   U16377 : NOR2_X1 port map( A1 => n14159, A2 => n15509, ZN => n14965);
   U16378 : OAI21_X1 port map( B1 => n14966, B2 => n15562, A => n14965, ZN => 
                           n14967);
   U16379 : XNOR2_X1 port map( A => n16974, B => n17366, ZN => n16288);
   U16380 : XNOR2_X1 port map( A => n19849, B => n16288, ZN => n14970);
   U16382 : NAND2_X1 port map( A1 => n15756, A2 => n15588, ZN => n15992);
   U16383 : INV_X1 port map( A => n15992, ZN => n14974);
   U16384 : OAI21_X1 port map( B1 => n15755, B2 => n15588, A => n15760, ZN => 
                           n15989);
   U16385 : NOR2_X1 port map( A1 => n15756, A2 => n15758, ZN => n15991);
   U16386 : INV_X1 port map( A => n15991, ZN => n14972);
   U16387 : NAND3_X1 port map( A1 => n14972, A2 => n15992, A3 => n15587, ZN => 
                           n14973);
   U16388 : OAI21_X1 port map( B1 => n14974, B2 => n15989, A => n14973, ZN => 
                           n16078);
   U16391 : XNOR2_X1 port map( A => n16078, B => n17327, ZN => n17019);
   U16392 : NAND2_X1 port map( A1 => n15409, A2 => n15549, ZN => n14981);
   U16393 : OR2_X1 port map( A1 => n15549, A2 => n15553, ZN => n14980);
   U16394 : NOR2_X1 port map( A1 => n15181, A2 => n19502, ZN => n15522);
   U16395 : INV_X1 port map( A => n14982, ZN => n14983);
   U16396 : AND2_X1 port map( A1 => n15746, A2 => n15741, ZN => n15180);
   U16397 : INV_X1 port map( A => n15516, ZN => n15178);
   U16398 : NOR2_X1 port map( A1 => n15178, A2 => n15182, ZN => n14984);
   U16399 : INV_X1 port map( A => n15746, ZN => n15742);
   U16400 : XNOR2_X1 port map( A => n16961, B => n16944, ZN => n16528);
   U16401 : XNOR2_X1 port map( A => n17019, B => n16528, ZN => n14995);
   U16402 : INV_X1 port map( A => n15277, ZN => n14986);
   U16403 : NAND2_X1 port map( A1 => n19662, A2 => n15395, ZN => n14992);
   U16405 : INV_X1 port map( A => n2356, ZN => n19264);
   U16406 : XNOR2_X1 port map( A => n16227, B => n19264, ZN => n14993);
   U16407 : XNOR2_X1 port map( A => n16284, B => n14993, ZN => n14994);
   U16411 : NAND2_X1 port map( A1 => n15003, A2 => n15002, ZN => n15840);
   U16412 : AND2_X1 port map( A1 => n15628, A2 => n15627, ZN => n15837);
   U16413 : NAND2_X1 port map( A1 => n15837, A2 => n15840, ZN => n15006);
   U16414 : OAI21_X1 port map( B1 => n1288, B2 => n15839, A => n15627, ZN => 
                           n15004);
   U16415 : NAND2_X1 port map( A1 => n15004, A2 => n15100, ZN => n15005);
   U16416 : OAI211_X1 port map( C1 => n15626, C2 => n15100, A => n15006, B => 
                           n15005, ZN => n17360);
   U16417 : XNOR2_X1 port map( A => n16706, B => n17360, ZN => n16276);
   U16418 : INV_X1 port map( A => n15601, ZN => n15112);
   U16420 : OAI21_X1 port map( B1 => n15112, B2 => n15009, A => n15113, ZN => 
                           n15605);
   U16421 : NAND2_X1 port map( A1 => n15601, A2 => n15600, ZN => n15010);
   U16422 : AOI21_X1 port map( B1 => n15270, B2 => n15010, A => n20112, ZN => 
                           n15011);
   U16424 : XNOR2_X1 port map( A => n15935, B => n16236, ZN => n15012);
   U16425 : XNOR2_X1 port map( A => n16276, B => n15012, ZN => n15025);
   U16426 : NAND2_X1 port map( A1 => n15296, A2 => n15297, ZN => n15013);
   U16427 : AOI21_X1 port map( B1 => n15108, B2 => n15013, A => n15110, ZN => 
                           n15016);
   U16428 : NAND2_X1 port map( A1 => n15296, A2 => n15295, ZN => n15014);
   U16429 : AOI21_X1 port map( B1 => n15297, B2 => n15014, A => n15294, ZN => 
                           n15015);
   U16430 : NOR2_X2 port map( A1 => n15016, A2 => n15015, ZN => n16938);
   U16431 : NAND2_X1 port map( A1 => n15018, A2 => n15017, ZN => n15283);
   U16432 : NAND2_X1 port map( A1 => n15283, A2 => n20474, ZN => n15019);
   U16433 : AOI22_X2 port map( A1 => n15020, A2 => n15132, B1 => n15019, B2 => 
                           n19848, ZN => n17253);
   U16434 : XNOR2_X1 port map( A => n16938, B => n17253, ZN => n15023);
   U16435 : XNOR2_X1 port map( A => n864, B => n15021, ZN => n15022);
   U16436 : XNOR2_X1 port map( A => n15023, B => n15022, ZN => n15024);
   U16437 : XNOR2_X1 port map( A => n15025, B => n15024, ZN => n16251);
   U16438 : INV_X1 port map( A => n15380, ZN => n15164);
   U16439 : NOR2_X1 port map( A1 => n15164, A2 => n15028, ZN => n15029);
   U16440 : AOI21_X2 port map( B1 => n15033, B2 => n15167, A => n15032, ZN => 
                           n16554);
   U16441 : XNOR2_X1 port map( A => n16554, B => n16429, ZN => n15038);
   U16442 : NAND2_X1 port map( A1 => n15583, A2 => n3315, ZN => n15034);
   U16443 : OAI21_X1 port map( B1 => n15582, B2 => n15581, A => n15583, ZN => 
                           n15036);
   U16444 : XNOR2_X1 port map( A => n17358, B => n19158, ZN => n15037);
   U16445 : XNOR2_X1 port map( A => n15038, B => n15037, ZN => n15055);
   U16446 : OAI21_X1 port map( B1 => n20449, B2 => n15138, A => n20133, ZN => 
                           n15040);
   U16447 : AOI21_X1 port map( B1 => n15567, B2 => n15566, A => n942, ZN => 
                           n15041);
   U16448 : OAI22_X1 port map( A1 => n15043, A2 => n15042, B1 => n20182, B2 => 
                           n15041, ZN => n16707);
   U16449 : NOR2_X1 port map( A1 => n15796, A2 => n15791, ZN => n15044);
   U16450 : OAI21_X1 port map( B1 => n15045, B2 => n15044, A => n15577, ZN => 
                           n15048);
   U16451 : OAI21_X1 port map( B1 => n860, B2 => n15572, A => n15574, ZN => 
                           n15046);
   U16452 : NAND2_X1 port map( A1 => n15046, A2 => n15796, ZN => n15047);
   U16453 : NAND2_X1 port map( A1 => n15048, A2 => n15047, ZN => n16741);
   U16454 : INV_X1 port map( A => n15350, ZN => n15050);
   U16455 : INV_X1 port map( A => n15459, ZN => n15049);
   U16456 : AOI22_X1 port map( A1 => n15050, A2 => n20173, B1 => n15348, B2 => 
                           n15049, ZN => n15053);
   U16457 : NAND2_X1 port map( A1 => n15459, A2 => n15350, ZN => n15456);
   U16458 : OAI211_X1 port map( C1 => n19759, C2 => n15350, A => n15456, B => 
                           n15353, ZN => n15051);
   U16459 : XNOR2_X1 port map( A => n16741, B => n16873, ZN => n16355);
   U16460 : XNOR2_X1 port map( A => n16355, B => n16822, ZN => n15054);
   U16461 : XNOR2_X1 port map( A => n15054, B => n15055, ZN => n15220);
   U16462 : MUX2_X1 port map( A => n15553, B => n15056, S => n15551, Z => 
                           n15058);
   U16463 : MUX2_X1 port map( A => n14903, B => n20147, S => n15549, Z => 
                           n15057);
   U16464 : AOI22_X1 port map( A1 => n15311, A2 => n15061, B1 => n15395, B2 => 
                           n15060, ZN => n15063);
   U16466 : XNOR2_X1 port map( A => n16269, B => n16690, ZN => n15075);
   U16468 : NOR2_X1 port map( A1 => n15402, A2 => n19838, ZN => n15065);
   U16469 : NAND2_X1 port map( A1 => n15065, A2 => n20006, ZN => n15068);
   U16470 : NAND2_X1 port map( A1 => n15066, A2 => n15898, ZN => n15067);
   U16471 : AND3_X2 port map( A1 => n15069, A2 => n15068, A3 => n15067, ZN => 
                           n16770);
   U16472 : AND2_X1 port map( A1 => n15070, A2 => n15618, ZN => n15545);
   U16473 : NOR2_X1 port map( A1 => n15546, A2 => n15071, ZN => n15072);
   U16474 : XNOR2_X1 port map( A => n16770, B => n17098, ZN => n15074);
   U16475 : XNOR2_X1 port map( A => n15075, B => n15074, ZN => n15090);
   U16477 : INV_X1 port map( A => n15909, ZN => n15915);
   U16478 : NOR2_X1 port map( A1 => n15915, A2 => n15907, ZN => n15076);
   U16479 : NAND3_X1 port map( A1 => n15007, A2 => n15078, A3 => n15915, ZN => 
                           n15079);
   U16480 : XNOR2_X1 port map( A => n16600, B => n17411, ZN => n15088);
   U16481 : NAND2_X1 port map( A1 => n15081, A2 => n15430, ZN => n15532);
   U16482 : NAND2_X1 port map( A1 => n15082, A2 => n19676, ZN => n15085);
   U16483 : NOR2_X1 port map( A1 => n15921, A2 => n15422, ZN => n15431);
   U16484 : XNOR2_X1 port map( A => n15087, B => n15088, ZN => n15089);
   U16485 : XNOR2_X2 port map( A => n15090, B => n15089, ZN => n17243);
   U16486 : MUX2_X1 port map( A => n15092, B => n15091, S => n15846, Z => 
                           n15094);
   U16487 : MUX2_X1 port map( A => n15846, B => n15845, S => n15844, Z => 
                           n15093);
   U16488 : XNOR2_X1 port map( A => n17035, B => n16406, ZN => n15106);
   U16489 : NOR2_X1 port map( A1 => n15643, A2 => n15644, ZN => n15095);
   U16490 : NOR2_X1 port map( A1 => n19891, A2 => n15829, ZN => n15097);
   U16491 : MUX2_X1 port map( A => n15258, B => n15097, S => n14997, Z => 
                           n15098);
   U16492 : NOR2_X1 port map( A1 => n15838, A2 => n15840, ZN => n15105);
   U16493 : OAI21_X1 port map( B1 => n15100, B2 => n15628, A => n15625, ZN => 
                           n15104);
   U16494 : NAND3_X1 port map( A1 => n1288, A2 => n15836, A3 => n2472, ZN => 
                           n15103);
   U16495 : NOR2_X1 port map( A1 => n1288, A2 => n15628, ZN => n15101);
   U16497 : XNOR2_X1 port map( A => n16835, B => n15106, ZN => n15137);
   U16498 : INV_X1 port map( A => n15296, ZN => n15109);
   U16500 : NOR2_X1 port map( A1 => n15275, A2 => n15270, ZN => n15116);
   U16501 : NOR2_X1 port map( A1 => n15601, A2 => n15276, ZN => n15115);
   U16502 : MUX2_X1 port map( A => n15116, B => n15115, S => n15600, Z => 
                           n15117);
   U16503 : XNOR2_X1 port map( A => n17269, B => n17111, ZN => n16546);
   U16504 : NAND3_X1 port map( A1 => n15120, A2 => n15119, A3 => n20272, ZN => 
                           n15124);
   U16505 : NAND4_X1 port map( A1 => n15126, A2 => n15125, A3 => n15124, A4 => 
                           n15123, ZN => n15128);
   U16506 : INV_X1 port map( A => n15129, ZN => n15133);
   U16507 : NOR2_X1 port map( A1 => n15282, A2 => n20474, ZN => n15131);
   U16508 : INV_X1 port map( A => n645, ZN => n15134);
   U16509 : XNOR2_X1 port map( A => n16893, B => n15134, ZN => n15135);
   U16510 : XNOR2_X1 port map( A => n16546, B => n15135, ZN => n15136);
   U16511 : XNOR2_X1 port map( A => n16945, B => n2248, ZN => n15145);
   U16512 : INV_X1 port map( A => n20449, ZN => n15139);
   U16513 : NOR2_X1 port map( A1 => n15139, A2 => n15138, ZN => n15140);
   U16514 : NOR2_X1 port map( A1 => n15701, A2 => n15696, ZN => n15384);
   U16515 : MUX2_X1 port map( A => n15140, B => n15384, S => n15698, Z => 
                           n15144);
   U16516 : OR2_X1 port map( A1 => n15701, A2 => n15386, ZN => n15142);
   U16517 : AOI22_X1 port map( A1 => n15142, A2 => n15141, B1 => n15701, B2 => 
                           n15698, ZN => n15143);
   U16519 : XNOR2_X1 port map( A => n19720, B => n15145, ZN => n15158);
   U16520 : NOR2_X1 port map( A1 => n15712, A2 => n20178, ZN => n15147);
   U16522 : NOR2_X1 port map( A1 => n15147, A2 => n15146, ZN => n15151);
   U16524 : NAND2_X1 port map( A1 => n15152, A2 => n16015, ZN => n15156);
   U16525 : OAI21_X1 port map( B1 => n192, B2 => n20119, A => n19739, ZN => 
                           n15154);
   U16526 : OAI21_X2 port map( B1 => n15156, B2 => n16016, A => n15155, ZN => 
                           n16854);
   U16527 : INV_X1 port map( A => n16854, ZN => n15157);
   U16528 : XNOR2_X1 port map( A => n15157, B => n16900, ZN => n16342);
   U16529 : XNOR2_X1 port map( A => n16342, B => n15158, ZN => n15176);
   U16530 : OR2_X1 port map( A1 => n15500, A2 => n15195, ZN => n15162);
   U16531 : NOR2_X1 port map( A1 => n15501, A2 => n15496, ZN => n15190);
   U16532 : INV_X1 port map( A => n15190, ZN => n15161);
   U16533 : INV_X1 port map( A => n15192, ZN => n15499);
   U16534 : AND2_X1 port map( A1 => n15501, A2 => n15499, ZN => n15159);
   U16535 : OAI211_X1 port map( C1 => n15378, C2 => n20467, A => n15163, B => 
                           n19513, ZN => n15169);
   U16536 : OAI21_X1 port map( B1 => n15167, B2 => n15166, A => n15165, ZN => 
                           n15168);
   U16537 : XNOR2_X1 port map( A => n17299, B => n16615, ZN => n15175);
   U16538 : INV_X1 port map( A => n15864, ZN => n15329);
   U16539 : AOI21_X2 port map( B1 => n15173, B2 => n15172, A => n15171, ZN => 
                           n17116);
   U16540 : INV_X1 port map( A => n17116, ZN => n15174);
   U16541 : XNOR2_X1 port map( A => n15175, B => n15174, ZN => n15998);
   U16542 : INV_X1 port map( A => n20354, ZN => n17484);
   U16543 : NAND2_X1 port map( A1 => n15177, A2 => n17484, ZN => n15254);
   U16544 : NOR2_X1 port map( A1 => n15178, A2 => n15741, ZN => n15179);
   U16545 : NAND2_X1 port map( A1 => n15521, A2 => n19502, ZN => n15184);
   U16546 : NAND3_X1 port map( A1 => n15182, A2 => n15741, A3 => n15745, ZN => 
                           n15183);
   U16547 : OAI21_X1 port map( B1 => n15748, B2 => n15184, A => n15183, ZN => 
                           n15185);
   U16548 : XNOR2_X1 port map( A => n16608, B => n17438, ZN => n15199);
   U16549 : NAND2_X1 port map( A1 => n15190, A2 => n15500, ZN => n15198);
   U16550 : AOI21_X1 port map( B1 => n19813, B2 => n15192, A => n15191, ZN => 
                           n15193);
   U16551 : AOI21_X1 port map( B1 => n19512, B2 => n15501, A => n15193, ZN => 
                           n15197);
   U16552 : NOR2_X1 port map( A1 => n15195, A2 => n19813, ZN => n15196);
   U16553 : XNOR2_X1 port map( A => n16562, B => n16746, ZN => n15887);
   U16554 : XNOR2_X1 port map( A => n15199, B => n15887, ZN => n15219);
   U16555 : MUX2_X1 port map( A => n15495, B => n16128, S => n16129, Z => 
                           n15203);
   U16556 : NOR2_X1 port map( A1 => n16126, A2 => n15608, ZN => n15200);
   U16557 : INV_X1 port map( A => n15758, ZN => n15204);
   U16558 : OAI21_X1 port map( B1 => n15758, B2 => n15754, A => n15755, ZN => 
                           n15207);
   U16559 : NAND2_X1 port map( A1 => n15208, A2 => n15760, ZN => n15206);
   U16561 : NAND3_X1 port map( A1 => n15491, A2 => n2247, A3 => n15588, ZN => 
                           n15205);
   U16562 : XNOR2_X1 port map( A => n16844, B => n16747, ZN => n15217);
   U16563 : NOR2_X1 port map( A1 => n15559, A2 => n15513, ZN => n15209);
   U16564 : NAND2_X1 port map( A1 => n15212, A2 => n15560, ZN => n15213);
   U16565 : AOI21_X1 port map( B1 => n15211, B2 => n15213, A => n15558, ZN => 
                           n15214);
   U16567 : INV_X1 port map( A => n18779, ZN => n18784);
   U16568 : XNOR2_X1 port map( A => n20477, B => n18784, ZN => n15216);
   U16569 : XNOR2_X1 port map( A => n15216, B => n15217, ZN => n15218);
   U16570 : INV_X1 port map( A => n15220, ZN => n17483);
   U16571 : NAND2_X1 port map( A1 => n17245, A2 => n17483, ZN => n15252);
   U16572 : OR2_X1 port map( A1 => n19884, A2 => n15221, ZN => n15222);
   U16573 : AOI22_X1 port map( A1 => n15438, A2 => n15222, B1 => n20151, B2 => 
                           n15770, ZN => n15224);
   U16574 : NOR2_X1 port map( A1 => n15222, A2 => n15673, ZN => n15223);
   U16575 : OR2_X2 port map( A1 => n15224, A2 => n15223, ZN => n16760);
   U16576 : XNOR2_X1 port map( A => n16760, B => n18997, ZN => n15225);
   U16577 : INV_X1 port map( A => n15226, ZN => n15227);
   U16578 : NAND2_X1 port map( A1 => n15686, A2 => n15777, ZN => n15451);
   U16579 : NOR2_X1 port map( A1 => n15682, A2 => n15228, ZN => n15449);
   U16581 : NAND3_X1 port map( A1 => n15229, A2 => n15446, A3 => n1494, ZN => 
                           n15230);
   U16582 : XNOR2_X1 port map( A => n16330, B => n16861, ZN => n16887);
   U16584 : INV_X1 port map( A => n15234, ZN => n15236);
   U16585 : NAND2_X1 port map( A1 => n15465, A2 => n15339, ZN => n15338);
   U16586 : NAND2_X1 port map( A1 => n15338, A2 => n15468, ZN => n15233);
   U16587 : OAI21_X1 port map( B1 => n15234, B2 => n15467, A => n15233, ZN => 
                           n15235);
   U16588 : OAI21_X1 port map( B1 => n15470, B2 => n15236, A => n15235, ZN => 
                           n17367);
   U16589 : NAND2_X1 port map( A1 => n15459, A2 => n15237, ZN => n15238);
   U16590 : NAND2_X1 port map( A1 => n15239, A2 => n15238, ZN => n15242);
   U16591 : NOR2_X1 port map( A1 => n19759, A2 => n1458, ZN => n15240);
   U16592 : AOI22_X1 port map( A1 => n15240, A2 => n15458, B1 => n1458, B2 => 
                           n15350, ZN => n15241);
   U16593 : XNOR2_X1 port map( A => n17279, B => n17367, ZN => n15249);
   U16594 : INV_X1 port map( A => n15244, ZN => n15248);
   U16595 : INV_X1 port map( A => n15245, ZN => n15246);
   U16599 : XNOR2_X1 port map( A => n15250, B => n15968, ZN => n17480);
   U16602 : NOR2_X1 port map( A1 => n18425, A2 => n18427, ZN => n15255);
   U16603 : AOI21_X1 port map( B1 => n19702, B2 => n18425, A => n15255, ZN => 
                           n15530);
   U16604 : MUX2_X1 port map( A => n15259, B => n15258, S => n14997, Z => 
                           n15260);
   U16605 : AOI21_X2 port map( B1 => n15261, B2 => n15829, A => n15260, ZN => 
                           n17099);
   U16606 : NOR2_X1 port map( A1 => n15838, A2 => n15625, ZN => n15265);
   U16607 : NAND2_X1 port map( A1 => n15265, A2 => n15840, ZN => n15263);
   U16608 : NAND3_X1 port map( A1 => n1288, A2 => n15627, A3 => n15625, ZN => 
                           n15262);
   U16609 : XNOR2_X1 port map( A => n17099, B => n16987, ZN => n16905);
   U16610 : MUX2_X1 port map( A => n15844, B => n15266, S => n15845, Z => 
                           n15269);
   U16611 : MUX2_X1 port map( A => n15845, B => n15267, S => n15636, Z => 
                           n15268);
   U16612 : XNOR2_X1 port map( A => n16905, B => n16691, ZN => n16577);
   U16613 : OAI211_X1 port map( C1 => n20112, C2 => n15275, A => n15272, B => 
                           n15271, ZN => n15280);
   U16614 : NOR2_X1 port map( A1 => n15275, A2 => n15274, ZN => n15599);
   U16615 : NAND2_X1 port map( A1 => n15599, A2 => n15276, ZN => n15279);
   U16616 : INV_X1 port map( A => Key(94), ZN => n19007);
   U16617 : INV_X1 port map( A => n15281, ZN => n15290);
   U16618 : NAND2_X1 port map( A1 => n15283, A2 => n15282, ZN => n15289);
   U16619 : OAI22_X1 port map( A1 => n15287, A2 => n15286, B1 => n15285, B2 => 
                           n19848, ZN => n15288);
   U16621 : XNOR2_X1 port map( A => n15291, B => n17102, ZN => n15300);
   U16622 : NAND2_X1 port map( A1 => n15293, A2 => n15292, ZN => n15299);
   U16623 : NAND2_X1 port map( A1 => n15294, A2 => n15295, ZN => n15298);
   U16624 : XNOR2_X1 port map( A => n16600, B => n16095, ZN => n16384);
   U16625 : XNOR2_X1 port map( A => n15300, B => n16384, ZN => n15301);
   U16626 : XNOR2_X1 port map( A => n16577, B => n15301, ZN => n16166);
   U16627 : OAI21_X1 port map( B1 => n15875, B2 => n198, A => n15874, ZN => 
                           n15304);
   U16628 : NAND2_X1 port map( A1 => n20094, A2 => n15304, ZN => n15305);
   U16629 : NAND2_X1 port map( A1 => n15309, A2 => n15308, ZN => n15394);
   U16630 : AND2_X1 port map( A1 => n15312, A2 => n15676, ZN => n15325);
   U16631 : NOR2_X1 port map( A1 => n15314, A2 => n15313, ZN => n15322);
   U16632 : INV_X1 port map( A => n15315, ZN => n15318);
   U16633 : INV_X1 port map( A => n15316, ZN => n15317);
   U16634 : NAND2_X1 port map( A1 => n15318, A2 => n15317, ZN => n15319);
   U16635 : MUX2_X1 port map( A => n15320, B => n15319, S => n2731, Z => n15321
                           );
   U16636 : INV_X1 port map( A => n15677, ZN => n15447);
   U16637 : OAI211_X1 port map( C1 => n15322, C2 => n15321, A => n15447, B => 
                           n15443, ZN => n15323);
   U16638 : XNOR2_X1 port map( A => n20167, B => n17358, ZN => n15326);
   U16639 : XNOR2_X1 port map( A => n17141, B => n15326, ZN => n15347);
   U16641 : OAI21_X1 port map( B1 => n15329, B2 => n15328, A => n15866, ZN => 
                           n15330);
   U16643 : AND2_X1 port map( A1 => n901, A2 => n20119, ZN => n15334);
   U16644 : XNOR2_X1 port map( A => n15979, B => n19807, ZN => n15345);
   U16646 : NAND2_X1 port map( A1 => n15340, A2 => n15339, ZN => n15342);
   U16647 : XNOR2_X1 port map( A => n19889, B => n17787, ZN => n15344);
   U16648 : XNOR2_X1 port map( A => n15345, B => n15344, ZN => n15346);
   U16649 : NAND2_X1 port map( A1 => n20173, A2 => n15348, ZN => n15462);
   U16650 : OAI21_X1 port map( B1 => n15458, B2 => n15350, A => n19759, ZN => 
                           n15351);
   U16651 : XNOR2_X1 port map( A => n19954, B => n16608, ZN => n15362);
   U16652 : NAND2_X1 port map( A1 => n15354, A2 => n233, ZN => n15356);
   U16653 : NAND3_X1 port map( A1 => n15815, A2 => n15582, A3 => n15583, ZN => 
                           n15355);
   U16654 : NAND2_X1 port map( A1 => n15356, A2 => n15355, ZN => n15360);
   U16655 : NOR2_X1 port map( A1 => n233, A2 => n15812, ZN => n15358);
   U16656 : NOR2_X1 port map( A1 => n3315, A2 => n15583, ZN => n15357);
   U16657 : XNOR2_X1 port map( A => n16359, B => n2369, ZN => n15361);
   U16658 : XNOR2_X1 port map( A => n15362, B => n15361, ZN => n15393);
   U16659 : OAI21_X1 port map( B1 => n860, B2 => n15573, A => n15574, ZN => 
                           n15363);
   U16660 : INV_X1 port map( A => n15363, ZN => n15369);
   U16661 : NAND2_X1 port map( A1 => n15364, A2 => n859, ZN => n15368);
   U16662 : MUX2_X1 port map( A => n15566, B => n15567, S => n15370, Z => 
                           n15374);
   U16664 : INV_X1 port map( A => n15565, ZN => n15372);
   U16665 : XNOR2_X1 port map( A => n17127, B => n16996, ZN => n16882);
   U16666 : INV_X1 port map( A => n15375, ZN => n15377);
   U16667 : NOR2_X1 port map( A1 => n15379, A2 => n231, ZN => n15376);
   U16668 : NOR2_X1 port map( A1 => n15377, A2 => n15376, ZN => n15383);
   U16669 : NAND2_X1 port map( A1 => n15384, A2 => n20133, ZN => n15391);
   U16670 : NAND2_X1 port map( A1 => n15386, A2 => n15695, ZN => n15387);
   U16671 : NAND3_X1 port map( A1 => n15701, A2 => n15702, A3 => n15387, ZN => 
                           n15390);
   U16672 : NAND3_X1 port map( A1 => n15385, A2 => n15696, A3 => n15698, ZN => 
                           n15389);
   U16673 : NAND3_X1 port map( A1 => n15387, A2 => n15702, A3 => n15386, ZN => 
                           n15388);
   U16674 : NAND4_X1 port map( A1 => n15391, A2 => n15390, A3 => n15389, A4 => 
                           n15388, ZN => n17442);
   U16675 : XNOR2_X1 port map( A => n17442, B => n16840, ZN => n16102);
   U16676 : XNOR2_X1 port map( A => n16882, B => n16102, ZN => n15392);
   U16677 : XNOR2_X1 port map( A => n15392, B => n15393, ZN => n16165);
   U16678 : NAND3_X1 port map( A1 => n17505, A2 => n17501, A3 => n16165, ZN => 
                           n16443);
   U16679 : OAI22_X1 port map( A1 => n15397, A2 => n15396, B1 => n15395, B2 => 
                           n15394, ZN => n15398);
   U16680 : XNOR2_X1 port map( A => n16761, B => n17367, ZN => n16380);
   U16682 : OAI211_X1 port map( C1 => n20006, C2 => n15892, A => n15402, B => 
                           n15536, ZN => n15404);
   U16683 : XNOR2_X1 port map( A => n17135, B => n16380, ZN => n15436);
   U16684 : XNOR2_X1 port map( A => n17133, B => n2420, ZN => n15434);
   U16685 : OR2_X1 port map( A1 => n15417, A2 => n15416, ZN => n15418);
   U16686 : OAI21_X2 port map( B1 => n15912, B2 => n15419, A => n15418, ZN => 
                           n17276);
   U16688 : OAI21_X1 port map( B1 => n15426, B2 => n15423, A => n15422, ZN => 
                           n15429);
   U16689 : INV_X1 port map( A => n15424, ZN => n15425);
   U16690 : NOR2_X1 port map( A1 => n15426, A2 => n15425, ZN => n15428);
   U16691 : NAND2_X1 port map( A1 => n15430, A2 => n15531, ZN => n15427);
   U16693 : INV_X1 port map( A => n15431, ZN => n15432);
   U16694 : AOI22_X2 port map( A1 => n15917, A2 => n15534, B1 => n15433, B2 => 
                           n15432, ZN => n16971);
   U16695 : XNOR2_X1 port map( A => n17276, B => n16971, ZN => n16567);
   U16696 : XNOR2_X1 port map( A => n15434, B => n16567, ZN => n15435);
   U16697 : XNOR2_X1 port map( A => n15436, B => n15435, ZN => n15485);
   U16698 : NOR2_X1 port map( A1 => n15665, A2 => n19884, ZN => n15437);
   U16699 : OAI21_X1 port map( B1 => n15438, B2 => n15437, A => n15673, ZN => 
                           n15441);
   U16700 : AND2_X1 port map( A1 => n19884, A2 => n15666, ZN => n15439);
   U16701 : NAND2_X1 port map( A1 => n15441, A2 => n15440, ZN => n16134);
   U16703 : NAND2_X1 port map( A1 => n15446, A2 => n15443, ZN => n15444);
   U16704 : NAND2_X1 port map( A1 => n15447, A2 => n15446, ZN => n15448);
   U16705 : XNOR2_X1 port map( A => n16134, B => n20481, ZN => n16898);
   U16706 : NAND2_X1 port map( A1 => n15783, A2 => n15684, ZN => n15450);
   U16710 : OAI211_X1 port map( C1 => n15459, C2 => n20173, A => n15456, B => 
                           n1458, ZN => n15463);
   U16711 : NAND3_X1 port map( A1 => n15460, A2 => n15459, A3 => n15458, ZN => 
                           n15461);
   U16712 : AND3_X1 port map( A1 => n15463, A2 => n15462, A3 => n15461, ZN => 
                           n16367);
   U16713 : XNOR2_X1 port map( A => n16963, B => n16367, ZN => n15633);
   U16714 : XNOR2_X1 port map( A => n16898, B => n15633, ZN => n15483);
   U16715 : NOR2_X1 port map( A1 => n15470, A2 => n15468, ZN => n15471);
   U16716 : XNOR2_X1 port map( A => n16615, B => n17298, ZN => n15481);
   U16717 : NOR2_X1 port map( A1 => n15766, A2 => n15769, ZN => n15473);
   U16719 : AND2_X1 port map( A1 => n12658, A2 => n15657, ZN => n15654);
   U16720 : INV_X1 port map( A => n15654, ZN => n15477);
   U16721 : NAND3_X1 port map( A1 => n15475, A2 => n15658, A3 => n15653, ZN => 
                           n15476);
   U16722 : XNOR2_X1 port map( A => n17401, B => n17909, ZN => n15480);
   U16723 : XNOR2_X1 port map( A => n15481, B => n15480, ZN => n15482);
   U16724 : XNOR2_X1 port map( A => n15483, B => n15482, ZN => n17498);
   U16728 : AOI21_X1 port map( B1 => n1683, B2 => n2247, A => n15755, ZN => 
                           n15493);
   U16729 : NAND3_X1 port map( A1 => n15488, A2 => n15757, A3 => n15487, ZN => 
                           n15489);
   U16730 : NOR2_X1 port map( A1 => n15759, A2 => n15489, ZN => n15492);
   U16731 : NOR2_X1 port map( A1 => n15491, A2 => n15490, ZN => n15761);
   U16732 : NOR2_X1 port map( A1 => n16126, A2 => n16128, ZN => n15494);
   U16733 : NAND2_X1 port map( A1 => n1019, A2 => n15503, ZN => n15821);
   U16734 : NAND2_X1 port map( A1 => n15506, A2 => n15505, ZN => n15824);
   U16735 : OR2_X1 port map( A1 => n15824, A2 => n13933, ZN => n15508);
   U16736 : XNOR2_X1 port map( A => n16892, B => n15726, ZN => n15526);
   U16737 : NAND2_X1 port map( A1 => n15511, A2 => n15513, ZN => n15512);
   U16738 : XNOR2_X1 port map( A => n17035, B => n19909, ZN => n15524);
   U16739 : NOR2_X1 port map( A1 => n15746, A2 => n15516, ZN => n15595);
   U16740 : INV_X1 port map( A => n15741, ZN => n15517);
   U16741 : NAND3_X1 port map( A1 => n15517, A2 => n15742, A3 => n19502, ZN => 
                           n15518);
   U16744 : XNOR2_X1 port map( A => n16335, B => n2123, ZN => n15523);
   U16745 : XNOR2_X1 port map( A => n15524, B => n15523, ZN => n15525);
   U16747 : OAI21_X1 port map( B1 => n20168, B2 => n19815, A => n19898, ZN => 
                           n15527);
   U16748 : NAND2_X1 port map( A1 => n15527, A2 => n16480, ZN => n15528);
   U16749 : NAND2_X1 port map( A1 => n15530, A2 => n15529, ZN => n15930);
   U16750 : XNOR2_X1 port map( A => n17002, B => n16236, ZN => n15543);
   U16752 : OAI21_X1 port map( B1 => n15539, B2 => n15538, A => n15537, ZN => 
                           n15542);
   U16753 : XNOR2_X1 port map( A => n17355, B => n16181, ZN => n17419);
   U16754 : XNOR2_X1 port map( A => n17419, B => n15543, ZN => n15557);
   U16755 : NOR2_X1 port map( A1 => n15545, A2 => n15544, ZN => n15548);
   U16756 : AOI21_X1 port map( B1 => n15550, B2 => n15549, A => n14903, ZN => 
                           n15552);
   U16757 : XNOR2_X1 port map( A => n17359, B => n16872, ZN => n15555);
   U16758 : XNOR2_X1 port map( A => n19889, B => n18984, ZN => n15554);
   U16759 : XNOR2_X1 port map( A => n15555, B => n15554, ZN => n15556);
   U16760 : INV_X1 port map( A => n16666, ZN => n17221);
   U16762 : INV_X1 port map( A => n15566, ZN => n15800);
   U16763 : NAND3_X1 port map( A1 => n15800, A2 => n15567, A3 => n15371, ZN => 
                           n15568);
   U16765 : XNOR2_X1 port map( A => n17014, B => n16788, ZN => n15571);
   U16767 : AND2_X1 port map( A1 => n15572, A2 => n15573, ZN => n15576);
   U16768 : NAND2_X1 port map( A1 => n15574, A2 => n15573, ZN => n15575);
   U16769 : MUX2_X1 port map( A => n15576, B => n15575, S => n860, Z => n15578)
                           ;
   U16770 : XNOR2_X1 port map( A => n16095, B => n19713, ZN => n15579);
   U16772 : MUX2_X1 port map( A => n15582, B => n15812, S => n15815, Z => 
                           n15585);
   U16773 : MUX2_X2 port map( A => n15585, B => n15584, S => n233, Z => n17406)
                           ;
   U16774 : XNOR2_X1 port map( A => n15586, B => n16132, ZN => n16639);
   U16775 : INV_X1 port map( A => n16641, ZN => n15731);
   U16776 : INV_X1 port map( A => n16639, ZN => n19385);
   U16777 : XNOR2_X1 port map( A => n16761, B => n2381, ZN => n15592);
   U16779 : MUX2_X1 port map( A => n15589, B => n15755, S => n15760, Z => 
                           n15590);
   U16780 : XNOR2_X1 port map( A => n15592, B => n16928, ZN => n15598);
   U16781 : NAND2_X1 port map( A1 => n3821, A2 => n15741, ZN => n15597);
   U16782 : NAND2_X1 port map( A1 => n15744, A2 => n15595, ZN => n15596);
   U16784 : XNOR2_X1 port map( A => n16886, B => n17133, ZN => n16146);
   U16785 : XNOR2_X1 port map( A => n15598, B => n16146, ZN => n15613);
   U16786 : INV_X1 port map( A => n15599, ZN => n15603);
   U16787 : NOR2_X1 port map( A1 => n15601, A2 => n15600, ZN => n15602);
   U16788 : NOR2_X1 port map( A1 => n15608, A2 => n16129, ZN => n15610);
   U16789 : NOR2_X1 port map( A1 => n3427, A2 => n16128, ZN => n15609);
   U16790 : AOI22_X1 port map( A1 => n15733, A2 => n15610, B1 => n15609, B2 => 
                           n16126, ZN => n15611);
   U16791 : XNOR2_X1 port map( A => n16970, B => n16932, ZN => n17431);
   U16792 : XNOR2_X1 port map( A => n17431, B => n16329, ZN => n15612);
   U16793 : OAI22_X1 port map( A1 => n15616, A2 => n20138, B1 => n15620, B2 => 
                           n15614, ZN => n15624);
   U16794 : INV_X1 port map( A => n15617, ZN => n15622);
   U16795 : NAND3_X1 port map( A1 => n15620, A2 => n15619, A3 => n15618, ZN => 
                           n15621);
   U16796 : NAND2_X1 port map( A1 => n15622, A2 => n15621, ZN => n15623);
   U16797 : INV_X1 port map( A => n15840, ZN => n15629);
   U16798 : NAND2_X1 port map( A1 => n15629, A2 => n15625, ZN => n15632);
   U16799 : NAND3_X1 port map( A1 => n15629, A2 => n1288, A3 => n15628, ZN => 
                           n15630);
   U16800 : OAI211_X1 port map( C1 => n15838, C2 => n15632, A => n15631, B => 
                           n15630, ZN => n16947);
   U16801 : XNOR2_X1 port map( A => n16947, B => n16960, ZN => n17399);
   U16802 : XNOR2_X1 port map( A => n17399, B => n15633, ZN => n15652);
   U16804 : NOR2_X1 port map( A1 => n15844, A2 => n868, ZN => n15634);
   U16805 : NAND2_X1 port map( A1 => n15845, A2 => n15634, ZN => n15638);
   U16806 : NOR2_X1 port map( A1 => n15846, A2 => n868, ZN => n15635);
   U16808 : XNOR2_X1 port map( A => n16227, B => n16412, ZN => n16902);
   U16809 : NAND3_X1 port map( A1 => n15643, A2 => n15645, A3 => n15642, ZN => 
                           n15648);
   U16810 : NAND3_X1 port map( A1 => n15645, A2 => n15644, A3 => n19931, ZN => 
                           n15647);
   U16811 : XNOR2_X1 port map( A => n17330, B => n18478, ZN => n15650);
   U16812 : XNOR2_X1 port map( A => n16902, B => n15650, ZN => n15651);
   U16813 : XNOR2_X1 port map( A => n15651, B => n15652, ZN => n19382);
   U16814 : INV_X1 port map( A => n19382, ZN => n17218);
   U16815 : XNOR2_X1 port map( A => n16240, B => n16840, ZN => n15675);
   U16816 : NAND2_X1 port map( A1 => n15654, A2 => n15653, ZN => n15663);
   U16817 : NAND3_X1 port map( A1 => n15659, A2 => n15658, A3 => n15657, ZN => 
                           n15662);
   U16818 : NAND3_X1 port map( A1 => n15768, A2 => n15769, A3 => n15660, ZN => 
                           n15661);
   U16819 : INV_X1 port map( A => n19879, ZN => n15773);
   U16820 : NAND3_X1 port map( A1 => n15773, A2 => n15665, A3 => n13414, ZN => 
                           n15669);
   U16821 : NAND2_X1 port map( A1 => n19879, A2 => n20151, ZN => n15674);
   U16822 : XNOR2_X1 port map( A => n16295, B => n955, ZN => n17440);
   U16823 : XNOR2_X1 port map( A => n15675, B => n17440, ZN => n15694);
   U16824 : NOR2_X1 port map( A1 => n15679, A2 => n15677, ZN => n15681);
   U16825 : INV_X1 port map( A => n15678, ZN => n15680);
   U16826 : INV_X1 port map( A => n2122, ZN => n18598);
   U16827 : XNOR2_X1 port map( A => n17444, B => n18598, ZN => n15692);
   U16828 : NAND2_X1 port map( A1 => n19977, A2 => n15683, ZN => n15785);
   U16829 : NAND3_X1 port map( A1 => n19978, A2 => n15782, A3 => n15684, ZN => 
                           n15690);
   U16830 : XNOR2_X1 port map( A => n16292, B => n19798, ZN => n16513);
   U16831 : XNOR2_X1 port map( A => n15692, B => n16513, ZN => n15693);
   U16832 : XNOR2_X1 port map( A => n15694, B => n15693, ZN => n19386);
   U16833 : MUX2_X1 port map( A => n15701, B => n15696, S => n15695, Z => 
                           n15703);
   U16834 : AND2_X1 port map( A1 => n15702, A2 => n15698, ZN => n15700);
   U16835 : OAI21_X1 port map( B1 => n15885, B2 => n15705, A => n15704, ZN => 
                           n15707);
   U16836 : INV_X1 port map( A => n15957, ZN => n15708);
   U16837 : XNOR2_X1 port map( A => n17335, B => n15708, ZN => n17424);
   U16838 : INV_X1 port map( A => n15874, ZN => n15871);
   U16839 : NAND3_X1 port map( A1 => n15871, A2 => n20178, A3 => n15875, ZN => 
                           n15710);
   U16840 : OAI21_X1 port map( B1 => n15712, B2 => n15711, A => n15710, ZN => 
                           n15718);
   U16841 : INV_X1 port map( A => n15713, ZN => n15716);
   U16842 : XNOR2_X1 port map( A => n16027, B => n17095, ZN => n15719);
   U16843 : XNOR2_X1 port map( A => n17424, B => n15719, ZN => n15728);
   U16844 : OAI21_X1 port map( B1 => n15864, B2 => n15720, A => n15863, ZN => 
                           n15724);
   U16845 : NOR3_X1 port map( A1 => n15866, A2 => n15722, A3 => n15721, ZN => 
                           n15723);
   U16846 : XNOR2_X1 port map( A => n20102, B => n16336, ZN => n16891);
   U16847 : XNOR2_X1 port map( A => n16891, B => n15726, ZN => n15727);
   U16848 : XNOR2_X1 port map( A => n15727, B => n15728, ZN => n16665);
   U16849 : OAI211_X1 port map( C1 => n19386, C2 => n16666, A => n19383, B => 
                           n1897, ZN => n15729);
   U16850 : INV_X1 port map( A => n15729, ZN => n15730);
   U16851 : NOR2_X1 port map( A1 => n20003, A2 => n18412, ZN => n18424);
   U16852 : OAI211_X1 port map( C1 => n15495, C2 => n15737, A => n15736, B => 
                           n15735, ZN => n16097);
   U16853 : XNOR2_X1 port map( A => n15739, B => n16097, ZN => n15753);
   U16854 : INV_X1 port map( A => n15740, ZN => n15752);
   U16855 : NAND2_X1 port map( A1 => n15742, A2 => n15741, ZN => n15743);
   U16856 : NAND2_X1 port map( A1 => n15743, A2 => n15745, ZN => n15751);
   U16857 : NOR3_X1 port map( A1 => n15748, A2 => n15182, A3 => n15745, ZN => 
                           n15747);
   U16858 : AOI21_X1 port map( B1 => n15749, B2 => n15748, A => n15747, ZN => 
                           n15750);
   U16859 : OAI21_X1 port map( B1 => n15752, B2 => n15751, A => n15750, ZN => 
                           n16188);
   U16860 : XNOR2_X1 port map( A => n15753, B => n16188, ZN => n17101);
   U16861 : XNOR2_X1 port map( A => n16269, B => n16095, ZN => n16772);
   U16862 : XNOR2_X1 port map( A => n17101, B => n16772, ZN => n15764);
   U16863 : XNOR2_X1 port map( A => n17410, B => n457, ZN => n15762);
   U16864 : XNOR2_X1 port map( A => n15762, B => n19820, ZN => n15763);
   U16866 : XNOR2_X1 port map( A => n16742, B => n16873, ZN => n16071);
   U16867 : NAND2_X1 port map( A1 => n15771, A2 => n15770, ZN => n15776);
   U16868 : NAND2_X1 port map( A1 => n15778, A2 => n19977, ZN => n15787);
   U16869 : NAND3_X1 port map( A1 => n15783, A2 => n15782, A3 => n20362, ZN => 
                           n15784);
   U16871 : XNOR2_X1 port map( A => n16278, B => n16939, ZN => n17003);
   U16872 : XNOR2_X1 port map( A => n17003, B => n16071, ZN => n15790);
   U16873 : INV_X1 port map( A => n2347, ZN => n19259);
   U16874 : XNOR2_X1 port map( A => n16554, B => n19259, ZN => n15788);
   U16875 : XNOR2_X1 port map( A => n19889, B => n17416, ZN => n16107);
   U16876 : XNOR2_X1 port map( A => n16107, B => n15788, ZN => n15789);
   U16877 : INV_X1 port map( A => n16540, ZN => n19353);
   U16878 : NOR2_X1 port map( A1 => n19354, A2 => n19353, ZN => n16674);
   U16879 : MUX2_X1 port map( A => n860, B => n1520, S => n15365, Z => n15797);
   U16880 : OAI21_X1 port map( B1 => n15800, B2 => n15371, A => n20182, ZN => 
                           n15807);
   U16882 : NAND3_X1 port map( A1 => n15804, A2 => n942, A3 => n15803, ZN => 
                           n15805);
   U16883 : XNOR2_X1 port map( A => n17269, B => n19674, ZN => n15809);
   U16884 : XNOR2_X1 port map( A => n15810, B => n15809, ZN => n15827);
   U16885 : NAND2_X1 port map( A1 => n15814, A2 => n15813, ZN => n15817);
   U16886 : XNOR2_X1 port map( A => n17110, B => n16893, ZN => n16054);
   U16887 : AND2_X1 port map( A1 => n15821, A2 => n15820, ZN => n15826);
   U16888 : NAND2_X1 port map( A1 => n15822, A2 => n1758, ZN => n15823);
   U16889 : MUX2_X1 port map( A => n15824, B => n15823, S => n13933, Z => 
                           n15825);
   U16890 : NAND2_X1 port map( A1 => n15826, A2 => n15825, ZN => n16081);
   U16891 : XNOR2_X1 port map( A => n16054, B => n16081, ZN => n16758);
   U16892 : NOR2_X1 port map( A1 => n15829, A2 => n15828, ZN => n15830);
   U16893 : OAI21_X1 port map( B1 => n15642, B2 => n15831, A => n15830, ZN => 
                           n15834);
   U16894 : NAND2_X1 port map( A1 => n15832, A2 => n15257, ZN => n15833);
   U16895 : INV_X1 port map( A => n16975, ZN => n15842);
   U16896 : XNOR2_X1 port map( A => n15842, B => n16973, ZN => n16214);
   U16898 : NAND2_X1 port map( A1 => n15845, A2 => n15844, ZN => n15850);
   U16899 : NAND3_X1 port map( A1 => n15847, A2 => n15846, A3 => n2146, ZN => 
                           n15849);
   U16901 : XNOR2_X1 port map( A => n16761, B => n15852, ZN => n16089);
   U16902 : XNOR2_X1 port map( A => n17279, B => n2079, ZN => n15853);
   U16903 : XNOR2_X1 port map( A => n15853, B => n16089, ZN => n15854);
   U16904 : XNOR2_X1 port map( A => n15854, B => n15855, ZN => n16672);
   U16905 : AND2_X1 port map( A1 => n16672, A2 => n19349, ZN => n15856);
   U16906 : OR2_X1 port map( A1 => n16674, A2 => n15856, ZN => n15929);
   U16907 : NAND2_X1 port map( A1 => n15859, A2 => n15858, ZN => n15869);
   U16908 : NOR2_X1 port map( A1 => n15863, A2 => n15862, ZN => n15865);
   U16910 : INV_X1 port map( A => n2442, ZN => n18924);
   U16911 : XNOR2_X1 port map( A => n17124, B => n18924, ZN => n15886);
   U16912 : NOR2_X1 port map( A1 => n15875, A2 => n15871, ZN => n15872);
   U16913 : NOR2_X2 port map( A1 => n15878, A2 => n15877, ZN => n17439);
   U16914 : NAND2_X1 port map( A1 => n16012, A2 => n20119, ZN => n15884);
   U16915 : OAI21_X1 port map( B1 => n16009, B2 => n901, A => n15880, ZN => 
                           n15881);
   U16916 : NAND2_X1 port map( A1 => n15881, A2 => n3473, ZN => n15883);
   U16917 : NAND3_X1 port map( A1 => n16009, A2 => n16010, A3 => n16015, ZN => 
                           n15882);
   U16918 : OAI211_X1 port map( C1 => n15885, C2 => n15884, A => n15883, B => 
                           n15882, ZN => n17128);
   U16919 : XNOR2_X1 port map( A => n17128, B => n17439, ZN => n16998);
   U16920 : XNOR2_X1 port map( A => n15886, B => n16998, ZN => n15889);
   U16921 : XNOR2_X1 port map( A => n16102, B => n15887, ZN => n15888);
   U16922 : NAND2_X1 port map( A1 => n19352, A2 => n19348, ZN => n15927);
   U16923 : INV_X1 port map( A => n15892, ZN => n15895);
   U16925 : OAI22_X1 port map( A1 => n15891, A2 => n15890, B1 => n15895, B2 => 
                           n19722, ZN => n15902);
   U16926 : NAND2_X1 port map( A1 => n19722, A2 => n15892, ZN => n15899);
   U16927 : OAI21_X1 port map( B1 => n15899, B2 => n15898, A => n15897, ZN => 
                           n15900);
   U16928 : INV_X1 port map( A => n15900, ZN => n15901);
   U16929 : XNOR2_X1 port map( A => n16900, B => n16283, ZN => n15904);
   U16930 : XNOR2_X1 port map( A => n20104, B => n18726, ZN => n15903);
   U16931 : XNOR2_X1 port map( A => n15904, B => n15903, ZN => n15926);
   U16932 : AOI21_X1 port map( B1 => n2723, B2 => n15906, A => n15905, ZN => 
                           n15914);
   U16933 : INV_X1 port map( A => n15907, ZN => n15908);
   U16934 : NOR2_X1 port map( A1 => n15909, A2 => n15908, ZN => n15911);
   U16935 : OAI21_X1 port map( B1 => n15912, B2 => n15911, A => n15910, ZN => 
                           n15913);
   U16936 : XNOR2_X1 port map( A => n16225, B => n16367, ZN => n16851);
   U16937 : AND2_X1 port map( A1 => n15917, A2 => n15916, ZN => n15924);
   U16938 : MUX2_X1 port map( A => n15920, B => n15919, S => n19752, Z => 
                           n15923);
   U16939 : XNOR2_X1 port map( A => n16224, B => n17401, ZN => n17120);
   U16940 : XNOR2_X1 port map( A => n16851, B => n17120, ZN => n15925);
   U16941 : XNOR2_X1 port map( A => n15925, B => n15926, ZN => n19347);
   U16942 : INV_X1 port map( A => n19347, ZN => n19351);
   U16943 : AOI21_X1 port map( B1 => n15927, B2 => n19351, A => n19349, ZN => 
                           n15928);
   U16944 : NOR2_X1 port map( A1 => n18400, A2 => n18423, ZN => n18414);
   U16946 : XNOR2_X1 port map( A => n16181, B => n20450, ZN => n15934);
   U16947 : INV_X1 port map( A => n17466, ZN => n15932);
   U16948 : XNOR2_X1 port map( A => n864, B => n15932, ZN => n15933);
   U16949 : XNOR2_X1 port map( A => n15934, B => n15933, ZN => n15938);
   U16950 : XNOR2_X1 port map( A => n15936, B => n15935, ZN => n16534);
   U16951 : XNOR2_X1 port map( A => n16938, B => n16278, ZN => n17418);
   U16952 : XNOR2_X1 port map( A => n17418, B => n16534, ZN => n15937);
   U16954 : XNOR2_X1 port map( A => n16932, B => n17275, ZN => n17028);
   U16955 : XNOR2_X1 port map( A => n16522, B => n17028, ZN => n15942);
   U16956 : XNOR2_X1 port map( A => n16974, B => n16568, ZN => n15940);
   U16957 : XNOR2_X1 port map( A => n16975, B => n2208, ZN => n15939);
   U16958 : XNOR2_X1 port map( A => n15940, B => n15939, ZN => n15941);
   U16960 : XNOR2_X1 port map( A => n16964, B => n16283, ZN => n15943);
   U16961 : XNOR2_X1 port map( A => n16528, B => n15943, ZN => n15946);
   U16962 : XNOR2_X1 port map( A => n16947, B => n19929, ZN => n17020);
   U16963 : XNOR2_X1 port map( A => n16134, B => n2298, ZN => n15944);
   U16964 : XNOR2_X1 port map( A => n17020, B => n15944, ZN => n15945);
   U16965 : XNOR2_X1 port map( A => n15946, B => n15945, ZN => n17080);
   U16966 : NAND2_X1 port map( A1 => n17823, A2 => n17080, ZN => n17828);
   U16967 : XNOR2_X1 port map( A => n17099, B => n19783, ZN => n15948);
   U16968 : XNOR2_X1 port map( A => n17288, B => n18055, ZN => n15947);
   U16969 : XNOR2_X1 port map( A => n15948, B => n15947, ZN => n15950);
   U16970 : XNOR2_X1 port map( A => n16602, B => n17014, ZN => n17409);
   U16971 : XNOR2_X1 port map( A => n17104, B => n17410, ZN => n16990);
   U16972 : XNOR2_X1 port map( A => n17409, B => n16990, ZN => n15949);
   U16973 : NOR2_X1 port map( A1 => n17825, A2 => n17172, ZN => n16777);
   U16974 : AOI21_X1 port map( B1 => n20239, B2 => n17828, A => n16777, ZN => 
                           n15965);
   U16975 : XNOR2_X1 port map( A => n15951, B => n17439, ZN => n15952);
   U16976 : XNOR2_X1 port map( A => n947, B => n955, ZN => n17046);
   U16977 : XNOR2_X1 port map( A => n17046, B => n15952, ZN => n15954);
   U16978 : XNOR2_X1 port map( A => n15953, B => n15954, ZN => n16262);
   U16979 : INV_X1 port map( A => n17823, ZN => n15962);
   U16980 : XNOR2_X1 port map( A => n16981, B => n17109, ZN => n15956);
   U16981 : XNOR2_X1 port map( A => n17425, B => n16300, ZN => n15955);
   U16982 : XNOR2_X1 port map( A => n15956, B => n15955, ZN => n15961);
   U16983 : XNOR2_X1 port map( A => n16836, B => n17426, ZN => n15959);
   U16984 : XNOR2_X1 port map( A => n902, B => n19205, ZN => n15958);
   U16985 : XNOR2_X1 port map( A => n15959, B => n15958, ZN => n15960);
   U16986 : XNOR2_X1 port map( A => n15961, B => n15960, ZN => n16263);
   U16987 : NAND2_X1 port map( A1 => n15962, A2 => n17079, ZN => n15963);
   U16988 : AOI21_X1 port map( B1 => n16262, B2 => n20239, A => n15963, ZN => 
                           n15964);
   U16989 : XNOR2_X1 port map( A => n17280, B => n19102, ZN => n15966);
   U16990 : XNOR2_X1 port map( A => n15966, B => n16971, ZN => n15967);
   U16991 : XNOR2_X1 port map( A => n20098, B => n16928, ZN => n16521);
   U16992 : XNOR2_X1 port map( A => n15967, B => n16521, ZN => n15969);
   U16994 : XNOR2_X1 port map( A => n17291, B => n19713, ZN => n16518);
   U16995 : XNOR2_X1 port map( A => n15970, B => n16690, ZN => n16574);
   U16996 : XNOR2_X1 port map( A => n16574, B => n16518, ZN => n15974);
   U16997 : XNOR2_X1 port map( A => n17012, B => n16987, ZN => n15972);
   U16998 : XNOR2_X1 port map( A => n16600, B => n2275, ZN => n15971);
   U16999 : XNOR2_X1 port map( A => n15972, B => n15971, ZN => n15973);
   U17001 : NOR2_X1 port map( A1 => n20275, A2 => n20507, ZN => n16003);
   U17002 : INV_X1 port map( A => n20507, ZN => n17074);
   U17003 : XNOR2_X1 port map( A => n17379, B => n2164, ZN => n15975);
   U17004 : XNOR2_X1 port map( A => n15975, B => n16996, ZN => n15976);
   U17005 : XNOR2_X1 port map( A => n16750, B => n16562, ZN => n17259);
   U17006 : XNOR2_X1 port map( A => n17259, B => n15976, ZN => n15978);
   U17007 : XNOR2_X1 port map( A => n20478, B => n17260, ZN => n17048);
   U17008 : XNOR2_X1 port map( A => n17048, B => n16608, ZN => n15977);
   U17009 : XNOR2_X1 port map( A => n16554, B => n16743, ZN => n17250);
   U17010 : XNOR2_X1 port map( A => n17358, B => n17253, ZN => n17040);
   U17011 : XNOR2_X1 port map( A => n17250, B => n17040, ZN => n15983);
   U17012 : INV_X1 port map( A => n2296, ZN => n15980);
   U17013 : XNOR2_X1 port map( A => n17359, B => n15980, ZN => n15981);
   U17014 : XNOR2_X1 port map( A => n16553, B => n15981, ZN => n15982);
   U17015 : OAI21_X1 port map( B1 => n17074, B2 => n20514, A => n17872, ZN => 
                           n16002);
   U17018 : XNOR2_X1 port map( A => n20372, B => n16546, ZN => n15988);
   U17019 : XNOR2_X1 port map( A => n16027, B => n16980, ZN => n15986);
   U17020 : XNOR2_X1 port map( A => n16755, B => n17999, ZN => n15985);
   U17021 : XNOR2_X1 port map( A => n15986, B => n15985, ZN => n15987);
   U17022 : NAND2_X1 port map( A1 => n16003, A2 => n17676, ZN => n16001);
   U17023 : INV_X1 port map( A => n17872, ZN => n17868);
   U17024 : OAI21_X1 port map( B1 => n15991, B2 => n15990, A => n15989, ZN => 
                           n15993);
   U17025 : NAND2_X1 port map( A1 => n15993, A2 => n15992, ZN => n17293);
   U17026 : XNOR2_X1 port map( A => n15994, B => n2222, ZN => n15995);
   U17027 : XNOR2_X1 port map( A => n15995, B => n17293, ZN => n15997);
   U17028 : XNOR2_X1 port map( A => n17294, B => n16965, ZN => n15996);
   U17029 : XNOR2_X1 port map( A => n15997, B => n15996, ZN => n15999);
   U17030 : XNOR2_X1 port map( A => n15998, B => n15999, ZN => n17867);
   U17031 : INV_X1 port map( A => n17867, ZN => n17078);
   U17033 : OAI211_X1 port map( C1 => n16003, C2 => n16002, A => n16001, B => 
                           n16000, ZN => n16155);
   U17034 : XNOR2_X1 port map( A => n17378, B => n17439, ZN => n16294);
   U17035 : XNOR2_X1 port map( A => n19799, B => n19216, ZN => n16004);
   U17036 : XNOR2_X1 port map( A => n16607, B => n16004, ZN => n16005);
   U17037 : XNOR2_X1 port map( A => n16294, B => n16005, ZN => n16007);
   U17038 : XNOR2_X1 port map( A => n16844, B => n16914, ZN => n16390);
   U17039 : XNOR2_X1 port map( A => n16390, B => n17438, ZN => n16006);
   U17040 : XNOR2_X1 port map( A => n16007, B => n16006, ZN => n17898);
   U17041 : NAND3_X1 port map( A1 => n16009, A2 => n19739, A3 => n16015, ZN => 
                           n16014);
   U17042 : OAI21_X1 port map( B1 => n16012, B2 => n901, A => n16010, ZN => 
                           n16013);
   U17043 : OAI211_X1 port map( C1 => n16016, C2 => n16015, A => n16014, B => 
                           n16013, ZN => n16018);
   U17044 : XNOR2_X1 port map( A => n16601, B => n17347, ZN => n16021);
   U17045 : INV_X1 port map( A => n404, ZN => n16019);
   U17046 : XNOR2_X1 port map( A => n16021, B => n16020, ZN => n16024);
   U17047 : XNOR2_X1 port map( A => n17410, B => n17348, ZN => n16022);
   U17048 : XNOR2_X1 port map( A => n19860, B => n16022, ZN => n16023);
   U17049 : XNOR2_X1 port map( A => n16023, B => n16024, ZN => n16025);
   U17050 : NAND2_X1 port map( A1 => n17898, A2 => n16025, ZN => n17895);
   U17051 : INV_X1 port map( A => n16025, ZN => n17069);
   U17052 : XNOR2_X1 port map( A => n17339, B => n17426, ZN => n16303);
   U17053 : XNOR2_X1 port map( A => n16695, B => n18863, ZN => n16026);
   U17054 : XNOR2_X1 port map( A => n16303, B => n16026, ZN => n16029);
   U17055 : XNOR2_X1 port map( A => n16406, B => n20192, ZN => n16953);
   U17056 : XNOR2_X1 port map( A => n20269, B => n16584, ZN => n16028);
   U17059 : NAND2_X1 port map( A1 => n17895, A2 => n16783, ZN => n16043);
   U17060 : XNOR2_X1 port map( A => n16928, B => n16587, ZN => n16200);
   U17061 : XNOR2_X1 port map( A => n16200, B => n16711, ZN => n17371);
   U17062 : INV_X1 port map( A => n16030, ZN => n19422);
   U17063 : XNOR2_X1 port map( A => n16975, B => n19422, ZN => n16031);
   U17064 : XNOR2_X1 port map( A => n16031, B => n16926, ZN => n16032);
   U17065 : XNOR2_X1 port map( A => n16931, B => n16861, ZN => n16588);
   U17066 : XNOR2_X1 port map( A => n16032, B => n16588, ZN => n16033);
   U17067 : XNOR2_X1 port map( A => n17295, B => n19720, ZN => n16619);
   U17068 : XNOR2_X1 port map( A => n16945, B => n16283, ZN => n16034);
   U17069 : XNOR2_X1 port map( A => n16619, B => n16034, ZN => n16038);
   U17070 : XNOR2_X1 port map( A => n16614, B => n17330, ZN => n16196);
   U17071 : XNOR2_X1 port map( A => n20126, B => n304, ZN => n16036);
   U17072 : XNOR2_X1 port map( A => n16196, B => n16036, ZN => n16037);
   U17073 : XNOR2_X1 port map( A => n16038, B => n16037, ZN => n17892);
   U17074 : MUX2_X1 port map( A => n19910, B => n17892, S => n17896, Z => 
                           n16042);
   U17075 : XNOR2_X1 port map( A => n16278, B => n16487, ZN => n16039);
   U17076 : XNOR2_X1 port map( A => n17357, B => n16039, ZN => n16041);
   U17077 : XNOR2_X1 port map( A => n17359, B => n16429, ZN => n16937);
   U17078 : XNOR2_X1 port map( A => n16936, B => n16707, ZN => n16596);
   U17079 : XNOR2_X1 port map( A => n19863, B => n16596, ZN => n16040);
   U17080 : XNOR2_X1 port map( A => n16769, B => n16906, ZN => n16049);
   U17081 : XNOR2_X1 port map( A => n17099, B => n17014, ZN => n16047);
   U17082 : XNOR2_X1 port map( A => n16047, B => n16046, ZN => n16048);
   U17084 : INV_X1 port map( A => n17666, ZN => n17668);
   U17085 : NOR2_X1 port map( A1 => n16052, A2 => n16051, ZN => n16053);
   U17086 : XNOR2_X1 port map( A => n17424, B => n16053, ZN => n16056);
   U17087 : XNOR2_X1 port map( A => n17109, B => n16336, ZN => n16140);
   U17088 : XNOR2_X1 port map( A => n16054, B => n16140, ZN => n16055);
   U17089 : XNOR2_X1 port map( A => n19882, B => n955, ZN => n16058);
   U17090 : XNOR2_X1 port map( A => n19705, B => n620, ZN => n16057);
   U17091 : XNOR2_X1 port map( A => n16058, B => n16057, ZN => n16061);
   U17092 : INV_X1 port map( A => n17444, ZN => n16059);
   U17093 : XNOR2_X1 port map( A => n17124, B => n16059, ZN => n16749);
   U17094 : XNOR2_X1 port map( A => n16746, B => n16240, ZN => n16878);
   U17095 : XNOR2_X1 port map( A => n16749, B => n16878, ZN => n16060);
   U17096 : XNOR2_X1 port map( A => n17399, B => n17119, ZN => n16065);
   U17097 : XNOR2_X1 port map( A => n16227, B => n16900, ZN => n16063);
   U17098 : XNOR2_X1 port map( A => n16853, B => n294, ZN => n16062);
   U17099 : XNOR2_X1 port map( A => n16063, B => n16062, ZN => n16064);
   U17100 : OAI22_X1 port map( A1 => n17668, A2 => n17876, B1 => n17879, B2 => 
                           n19832, ZN => n16070);
   U17101 : XNOR2_X1 port map( A => n16329, B => n16566, ZN => n16066);
   U17102 : XNOR2_X1 port map( A => n17431, B => n16066, ZN => n16069);
   U17103 : INV_X1 port map( A => n18439, ZN => n18443);
   U17104 : XNOR2_X1 port map( A => n16568, B => n18443, ZN => n16067);
   U17106 : NAND2_X1 port map( A1 => n16070, A2 => n17881, ZN => n16076);
   U17107 : XNOR2_X1 port map( A => n16071, B => n16871, ZN => n16074);
   U17108 : XNOR2_X1 port map( A => n16821, B => n17170, ZN => n16072);
   U17109 : XNOR2_X1 port map( A => n20219, B => n16072, ZN => n16073);
   U17110 : NOR2_X1 port map( A1 => n17666, A2 => n17878, ZN => n17882);
   U17112 : AOI22_X1 port map( A1 => n17882, A2 => n20217, B1 => n19930, B2 => 
                           n19832, ZN => n16075);
   U17114 : XNOR2_X1 port map( A => n16853, B => n17298, ZN => n16719);
   U17115 : XNOR2_X1 port map( A => n16367, B => n18433, ZN => n16077);
   U17116 : XNOR2_X1 port map( A => n16719, B => n16077, ZN => n16080);
   U17117 : XNOR2_X1 port map( A => n16078, B => n16854, ZN => n16617);
   U17118 : XNOR2_X1 port map( A => n16617, B => n17120, ZN => n16079);
   U17119 : XNOR2_X1 port map( A => n16080, B => n16079, ZN => n17886);
   U17120 : INV_X1 port map( A => n16982, ZN => n16219);
   U17121 : XNOR2_X1 port map( A => n16219, B => n19909, ZN => n17107);
   U17122 : XNOR2_X1 port map( A => n17107, B => n16083, ZN => n16087);
   U17123 : INV_X1 port map( A => n16373, ZN => n16084);
   U17124 : XNOR2_X1 port map( A => n17270, B => n19436, ZN => n16085);
   U17125 : XNOR2_X1 port map( A => n16696, B => n16085, ZN => n16086);
   U17126 : XNOR2_X1 port map( A => n17280, B => n18075, ZN => n16088);
   U17127 : XNOR2_X1 port map( A => n16089, B => n16088, ZN => n16093);
   U17128 : XNOR2_X1 port map( A => n16973, B => n16760, ZN => n16090);
   U17129 : XNOR2_X1 port map( A => n16090, B => n16091, ZN => n16092);
   U17130 : NOR2_X1 port map( A1 => n17886, A2 => n20185, ZN => n16101);
   U17131 : XNOR2_X1 port map( A => n16094, B => n16770, ZN => n16096);
   U17132 : XNOR2_X1 port map( A => n16096, B => n16828, ZN => n16100);
   U17133 : XNOR2_X1 port map( A => n16097, B => n17012, ZN => n16098);
   U17134 : XNOR2_X1 port map( A => n16098, B => n16691, ZN => n16099);
   U17135 : XNOR2_X1 port map( A => n19900, B => n17128, ZN => n16117);
   U17136 : XNOR2_X1 port map( A => n16117, B => n16102, ZN => n16105);
   U17137 : XNOR2_X1 port map( A => n16359, B => n19705, ZN => n16702);
   U17138 : XNOR2_X1 port map( A => n17260, B => n2349, ZN => n16103);
   U17139 : XNOR2_X1 port map( A => n16702, B => n16103, ZN => n16104);
   U17140 : XNOR2_X1 port map( A => n16104, B => n16105, ZN => n16261);
   U17141 : XNOR2_X1 port map( A => n16821, B => n17252, ZN => n16705);
   U17142 : XNOR2_X1 port map( A => n16939, B => n16741, ZN => n16122);
   U17143 : XNOR2_X1 port map( A => n16705, B => n16122, ZN => n16109);
   U17144 : INV_X1 port map( A => n2151, ZN => n18880);
   U17145 : XNOR2_X1 port map( A => n17253, B => n18880, ZN => n16106);
   U17146 : XNOR2_X1 port map( A => n16107, B => n16106, ZN => n16108);
   U17147 : NOR2_X1 port map( A1 => n16261, A2 => n17890, ZN => n16110);
   U17148 : NAND2_X1 port map( A1 => n16110, A2 => n17891, ZN => n16111);
   U17149 : OAI21_X1 port map( B1 => n17600, B2 => n3825, A => n16111, ZN => 
                           n16114);
   U17150 : INV_X1 port map( A => n17600, ZN => n16112);
   U17151 : INV_X1 port map( A => n17890, ZN => n17663);
   U17152 : NOR2_X1 port map( A1 => n16112, A2 => n17663, ZN => n16113);
   U17154 : INV_X1 port map( A => n19170, ZN => n18324);
   U17155 : NAND3_X1 port map( A1 => n16115, A2 => n18324, A3 => n20394, ZN => 
                           n16164);
   U17156 : XNOR2_X1 port map( A => n16292, B => n17127, ZN => n16116);
   U17157 : XNOR2_X1 port map( A => n16116, B => n16240, ZN => n16118);
   U17158 : XNOR2_X1 port map( A => n16118, B => n16117, ZN => n16121);
   U17160 : XNOR2_X1 port map( A => n16880, B => n16119, ZN => n16120);
   U17161 : XNOR2_X1 port map( A => n17002, B => n17535, ZN => n16123);
   U17162 : XNOR2_X1 port map( A => n16122, B => n16123, ZN => n16125);
   U17163 : XNOR2_X1 port map( A => n17360, B => n16872, ZN => n16182);
   U17164 : XNOR2_X1 port map( A => n16871, B => n16182, ZN => n16124);
   U17165 : NAND2_X1 port map( A1 => n20264, A2 => n17840, ZN => n16139);
   U17166 : XNOR2_X1 port map( A => n17349, B => n1996, ZN => n16130);
   U17167 : INV_X1 port map( A => n16126, ZN => n16127);
   U17168 : XNOR2_X1 port map( A => n17099, B => n16770, ZN => n16131);
   U17169 : NAND2_X1 port map( A1 => n16139, A2 => n17063, ZN => n17201);
   U17170 : INV_X1 port map( A => n17840, ZN => n16153);
   U17171 : XNOR2_X1 port map( A => n16224, B => n17328, ZN => n16946);
   U17172 : XNOR2_X1 port map( A => n16902, B => n16946, ZN => n16138);
   U17173 : XNOR2_X1 port map( A => n16963, B => n16134, ZN => n16136);
   U17174 : XNOR2_X1 port map( A => n16854, B => n18203, ZN => n16135);
   U17175 : XNOR2_X1 port map( A => n16136, B => n16135, ZN => n16137);
   U17176 : NAND2_X1 port map( A1 => n16139, A2 => n16731, ZN => n16152);
   U17177 : XNOR2_X1 port map( A => n17340, B => n16407, ZN => n16301);
   U17178 : XNOR2_X1 port map( A => n16301, B => n16140, ZN => n16144);
   U17179 : XNOR2_X1 port map( A => n19674, B => n18420, ZN => n16141);
   U17180 : XNOR2_X1 port map( A => n16142, B => n16141, ZN => n16143);
   U17182 : INV_X1 port map( A => n16973, ZN => n16929);
   U17183 : XNOR2_X1 port map( A => n16145, B => n16929, ZN => n16147);
   U17184 : XNOR2_X1 port map( A => n16147, B => n16146, ZN => n16150);
   U17185 : XNOR2_X1 port map( A => n16568, B => n16760, ZN => n16148);
   U17186 : XNOR2_X1 port map( A => n16329, B => n16148, ZN => n16149);
   U17187 : NAND2_X1 port map( A1 => n3826, A2 => n20423, ZN => n16151);
   U17188 : NAND2_X1 port map( A1 => n18157, A2 => n16155, ZN => n18156);
   U17189 : NAND2_X1 port map( A1 => n16154, A2 => n993, ZN => n16163);
   U17190 : INV_X1 port map( A => n16155, ZN => n18317);
   U17191 : NOR2_X1 port map( A1 => n18317, A2 => n20460, ZN => n16159);
   U17195 : INV_X1 port map( A => n16159, ZN => n16160);
   U17196 : NAND4_X1 port map( A1 => n18156, A2 => n16160, A3 => n2368, A4 => 
                           n19170, ZN => n16161);
   U17197 : NAND4_X1 port map( A1 => n16164, A2 => n16163, A3 => n20384, A4 => 
                           n16161, ZN => Ciphertext(144));
   U17199 : INV_X1 port map( A => n17501, ZN => n16794);
   U17201 : NAND3_X1 port map( A1 => n16794, A2 => n19815, A3 => n19924, ZN => 
                           n16168);
   U17202 : NAND2_X1 port map( A1 => n16794, A2 => n15485, ZN => n16167);
   U17205 : NOR2_X1 port map( A1 => n16634, A2 => n3573, ZN => n16174);
   U17206 : OAI21_X1 port map( B1 => n17508, B2 => n17507, A => n16172, ZN => 
                           n16173);
   U17207 : OAI21_X2 port map( B1 => n16632, B2 => n16174, A => n16173, ZN => 
                           n18498);
   U17208 : XNOR2_X1 port map( A => n16880, B => n17124, ZN => n16176);
   U17209 : XNOR2_X1 port map( A => n16176, B => n16175, ZN => n16180);
   U17210 : XNOR2_X1 port map( A => n955, B => n17377, ZN => n16178);
   U17211 : XNOR2_X1 port map( A => n19799, B => n19027, ZN => n16177);
   U17212 : XNOR2_X1 port map( A => n16178, B => n16177, ZN => n16179);
   U17213 : XNOR2_X1 port map( A => n16180, B => n16179, ZN => n17565);
   U17214 : INV_X1 port map( A => n17565, ZN => n17562);
   U17215 : XNOR2_X1 port map( A => n16742, B => n16181, ZN => n16183);
   U17216 : XNOR2_X1 port map( A => n16183, B => n16182, ZN => n16187);
   U17217 : XNOR2_X1 port map( A => n17359, B => n2455, ZN => n16184);
   U17218 : XNOR2_X1 port map( A => n16185, B => n16184, ZN => n16186);
   U17219 : XNOR2_X1 port map( A => n16187, B => n16186, ZN => n16320);
   U17220 : INV_X1 port map( A => n16320, ZN => n18535);
   U17221 : XNOR2_X1 port map( A => n17104, B => n17406, ZN => n16190);
   U17222 : XNOR2_X1 port map( A => n16188, B => n17348, ZN => n16189);
   U17223 : XNOR2_X1 port map( A => n16190, B => n16189, ZN => n16194);
   U17224 : XNOR2_X1 port map( A => n16601, B => n17014, ZN => n16192);
   U17225 : XNOR2_X1 port map( A => n19836, B => n621, ZN => n16191);
   U17226 : XNOR2_X1 port map( A => n16191, B => n16192, ZN => n16193);
   U17227 : XNOR2_X1 port map( A => n16194, B => n16193, ZN => n16321);
   U17228 : INV_X1 port map( A => n16321, ZN => n16790);
   U17229 : XNOR2_X1 port map( A => n16225, B => n16412, ZN => n16195);
   U17230 : XNOR2_X1 port map( A => n16284, B => n16195, ZN => n16199);
   U17231 : XNOR2_X1 port map( A => n16947, B => n2454, ZN => n16197);
   U17232 : XNOR2_X1 port map( A => n16197, B => n16196, ZN => n16198);
   U17233 : XNOR2_X1 port map( A => n16199, B => n16198, ZN => n17470);
   U17234 : XNOR2_X1 port map( A => n16200, B => n16288, ZN => n16204);
   U17235 : XNOR2_X1 port map( A => n16886, B => n880, ZN => n16202);
   U17236 : XNOR2_X1 port map( A => n16932, B => n17089, ZN => n16201);
   U17237 : XNOR2_X1 port map( A => n16202, B => n16201, ZN => n16203);
   U17238 : OAI22_X1 port map( A1 => n18535, A2 => n16790, B1 => n17470, B2 => 
                           n18534, ZN => n17163);
   U17240 : XNOR2_X1 port map( A => n902, B => n17338, ZN => n17034);
   U17241 : XNOR2_X1 port map( A => n16301, B => n17034, ZN => n16208);
   U17242 : XNOR2_X1 port map( A => n20192, B => n911, ZN => n16206);
   U17243 : XNOR2_X1 port map( A => n16300, B => n2087, ZN => n16205);
   U17244 : XNOR2_X1 port map( A => n16206, B => n16205, ZN => n16207);
   U17245 : INV_X1 port map( A => n17470, ZN => n16209);
   U17246 : OAI21_X1 port map( B1 => n17564, B2 => n20432, A => n16209, ZN => 
                           n16210);
   U17247 : NOR2_X1 port map( A1 => n18500, A2 => n18485, ZN => n17912);
   U17248 : XNOR2_X1 port map( A => n16927, B => n2192, ZN => n16213);
   U17249 : XNOR2_X1 port map( A => n16213, B => n17276, ZN => n16215);
   U17250 : XNOR2_X1 port map( A => n16215, B => n16214, ZN => n16218);
   U17251 : XNOR2_X1 port map( A => n16970, B => n879, ZN => n16216);
   U17252 : XNOR2_X1 port map( A => n16329, B => n16216, ZN => n16217);
   U17253 : XNOR2_X1 port map( A => n17335, B => n17426, ZN => n16979);
   U17254 : XNOR2_X1 port map( A => n16219, B => n19928, ZN => n16952);
   U17255 : XNOR2_X1 port map( A => n16979, B => n16952, ZN => n16223);
   U17256 : XNOR2_X1 port map( A => n16335, B => n19018, ZN => n16221);
   U17257 : XNOR2_X1 port map( A => n911, B => n897, ZN => n16220);
   U17258 : XNOR2_X1 port map( A => n16221, B => n16220, ZN => n16222);
   U17259 : XNOR2_X1 port map( A => n16224, B => n16283, ZN => n16962);
   U17260 : XNOR2_X1 port map( A => n16225, B => n16960, ZN => n16226);
   U17261 : XNOR2_X1 port map( A => n16962, B => n16226, ZN => n16230);
   U17262 : XNOR2_X1 port map( A => n17298, B => n16227, ZN => n16341);
   U17263 : XNOR2_X1 port map( A => n16944, B => n17791, ZN => n16228);
   U17264 : XNOR2_X1 port map( A => n16341, B => n16228, ZN => n16229);
   U17266 : XNOR2_X1 port map( A => n16988, B => n16691, ZN => n16231);
   U17267 : XNOR2_X1 port map( A => n16769, B => n16231, ZN => n16235);
   U17268 : INV_X1 port map( A => n20682, ZN => n18631);
   U17269 : XNOR2_X1 port map( A => n17410, B => n18631, ZN => n16233);
   U17270 : XNOR2_X1 port map( A => n16233, B => n16232, ZN => n16234);
   U17271 : XNOR2_X1 port map( A => n16742, B => n16939, ZN => n17142);
   U17272 : XNOR2_X1 port map( A => n17252, B => n16236, ZN => n16353);
   U17273 : XNOR2_X1 port map( A => n17142, B => n16353, ZN => n16239);
   U17274 : INV_X1 port map( A => n2423, ZN => n18506);
   U17275 : XNOR2_X1 port map( A => n17355, B => n18506, ZN => n16237);
   U17276 : XNOR2_X1 port map( A => n17418, B => n16237, ZN => n16238);
   U17277 : XNOR2_X1 port map( A => n16238, B => n16239, ZN => n16447);
   U17278 : INV_X1 port map( A => n16447, ZN => n17495);
   U17279 : XNOR2_X1 port map( A => n17443, B => n16240, ZN => n16241);
   U17280 : XNOR2_X1 port map( A => n16749, B => n16241, ZN => n16245);
   U17281 : INV_X1 port map( A => n16242, ZN => n19280);
   U17282 : XNOR2_X1 port map( A => n19743, B => n19280, ZN => n16243);
   U17283 : XNOR2_X1 port map( A => n16998, B => n16243, ZN => n16244);
   U17284 : XNOR2_X1 port map( A => n16245, B => n16244, ZN => n17491);
   U17285 : AND2_X1 port map( A1 => n17495, A2 => n17491, ZN => n16802);
   U17286 : NAND2_X1 port map( A1 => n16802, A2 => n16801, ZN => n16246);
   U17287 : OAI21_X1 port map( B1 => n16247, B2 => n16801, A => n16246, ZN => 
                           n16249);
   U17288 : NAND2_X1 port map( A1 => n16447, A2 => n17493, ZN => n16800);
   U17289 : NOR2_X1 port map( A1 => n16800, A2 => n17488, ZN => n16248);
   U17291 : NAND2_X1 port map( A1 => n17912, A2 => n19729, ZN => n16257);
   U17293 : INV_X1 port map( A => n20135, ZN => n17213);
   U17294 : NAND2_X1 port map( A1 => n16465, A2 => n17211, ZN => n16254);
   U17295 : NAND2_X1 port map( A1 => n16465, A2 => n20135, ZN => n16253);
   U17296 : INV_X1 port map( A => n17210, ZN => n16658);
   U17297 : NAND3_X1 port map( A1 => n16254, A2 => n16253, A3 => n16658, ZN => 
                           n16255);
   U17298 : INV_X1 port map( A => n18495, ZN => n18496);
   U17299 : NAND3_X1 port map( A1 => n18496, A2 => n893, A3 => n19816, ZN => 
                           n16256);
   U17300 : INV_X1 port map( A => n2023, ZN => n16258);
   U17301 : XNOR2_X1 port map( A => n16259, B => n16258, ZN => Ciphertext(27));
   U17302 : NAND2_X1 port map( A1 => n17891, A2 => n20185, ZN => n16260);
   U17303 : INV_X1 port map( A => n16261, ZN => n17602);
   U17305 : OAI21_X1 port map( B1 => n16262, B2 => n20239, A => n17822, ZN => 
                           n16264);
   U17306 : INV_X1 port map( A => n16263, ZN => n17824);
   U17307 : NAND3_X1 port map( A1 => n16262, A2 => n17079, A3 => n17823, ZN => 
                           n16265);
   U17308 : INV_X1 port map( A => n19209, ZN => n19202);
   U17309 : INV_X1 port map( A => n17898, ZN => n17182);
   U17310 : AND2_X1 port map( A1 => n17896, A2 => n17181, ZN => n16266);
   U17311 : OAI21_X1 port map( B1 => n17182, B2 => n19707, A => n16266, ZN => 
                           n16268);
   U17312 : NOR2_X1 port map( A1 => n17892, A2 => n19910, ZN => n17183);
   U17313 : INV_X1 port map( A => n16781, ZN => n17897);
   U17314 : NAND2_X1 port map( A1 => n17183, A2 => n17897, ZN => n16267);
   U17315 : XNOR2_X1 port map( A => n16269, B => n17104, ZN => n16271);
   U17316 : XNOR2_X1 port map( A => n17406, B => n17410, ZN => n16270);
   U17317 : XNOR2_X1 port map( A => n16270, B => n16271, ZN => n16275);
   U17318 : XNOR2_X1 port map( A => n16992, B => n17347, ZN => n16273);
   U17319 : XNOR2_X1 port map( A => n19836, B => n347, ZN => n16272);
   U17320 : XNOR2_X1 port map( A => n16272, B => n16273, ZN => n16274);
   U17321 : XNOR2_X2 port map( A => n16275, B => n16274, ZN => n19402);
   U17322 : XNOR2_X1 port map( A => n17002, B => n16872, ZN => n16277);
   U17323 : XNOR2_X1 port map( A => n16276, B => n16277, ZN => n16282);
   U17324 : XNOR2_X1 port map( A => n864, B => n16278, ZN => n16280);
   U17325 : XNOR2_X1 port map( A => n16873, B => n2383, ZN => n16279);
   U17326 : XNOR2_X1 port map( A => n16280, B => n16279, ZN => n16281);
   U17327 : XNOR2_X1 port map( A => n16282, B => n16281, ZN => n17650);
   U17328 : XNOR2_X1 port map( A => n16412, B => n16283, ZN => n17400);
   U17329 : XNOR2_X1 port map( A => n16963, B => n18887, ZN => n16285);
   U17330 : XNOR2_X1 port map( A => n16975, B => n16886, ZN => n17435);
   U17331 : XNOR2_X1 port map( A => n16330, B => n19222, ZN => n16286);
   U17332 : XNOR2_X1 port map( A => n17435, B => n16286, ZN => n16290);
   U17333 : XNOR2_X1 port map( A => n17133, B => n16711, ZN => n16287);
   U17334 : XNOR2_X1 port map( A => n16288, B => n16287, ZN => n16289);
   U17335 : XNOR2_X1 port map( A => n16289, B => n16290, ZN => n17853);
   U17336 : NAND2_X1 port map( A1 => n16306, A2 => n17853, ZN => n16291);
   U17337 : XNOR2_X1 port map( A => n16293, B => n19954, ZN => n17125);
   U17338 : XNOR2_X1 port map( A => n16294, B => n17125, ZN => n16299);
   U17340 : XNOR2_X1 port map( A => n16297, B => n16296, ZN => n16298);
   U17342 : INV_X1 port map( A => n17853, ZN => n17606);
   U17343 : XNOR2_X1 port map( A => n16507, B => n16300, ZN => n17108);
   U17344 : XNOR2_X1 port map( A => n17108, B => n16301, ZN => n16305);
   U17345 : XNOR2_X1 port map( A => n16893, B => n2317, ZN => n16302);
   U17346 : XNOR2_X1 port map( A => n16303, B => n16302, ZN => n16304);
   U17347 : XNOR2_X2 port map( A => n16305, B => n16304, ZN => n19404);
   U17348 : OAI21_X1 port map( B1 => n17606, B2 => n19404, A => n16306, ZN => 
                           n16307);
   U17349 : MUX2_X1 port map( A => n3345, B => n19930, S => n17876, Z => n16312
                           );
   U17350 : NOR2_X1 port map( A1 => n3345, A2 => n17879, ZN => n16310);
   U17351 : NOR2_X1 port map( A1 => n17881, A2 => n16308, ZN => n16309);
   U17352 : MUX2_X1 port map( A => n16310, B => n16309, S => n19930, Z => 
                           n16311);
   U17353 : AOI21_X2 port map( B1 => n16308, B2 => n16312, A => n16311, ZN => 
                           n19210);
   U17355 : MUX2_X1 port map( A => n19973, B => n20507, S => n17868, Z => 
                           n16317);
   U17356 : NAND2_X1 port map( A1 => n20506, A2 => n17873, ZN => n16315);
   U17357 : MUX2_X1 port map( A => n19190, B => n19210, S => n19842, Z => 
                           n16318);
   U17358 : NAND2_X1 port map( A1 => n16318, A2 => n19189, ZN => n16319);
   U17359 : AND2_X1 port map( A1 => n17564, A2 => n17470, ZN => n16789);
   U17360 : INV_X1 port map( A => n18534, ZN => n17468);
   U17361 : OAI21_X1 port map( B1 => n17468, B2 => n17564, A => n17471, ZN => 
                           n16325);
   U17362 : NOR2_X1 port map( A1 => n18539, A2 => n17471, ZN => n16323);
   U17363 : NOR2_X1 port map( A1 => n17564, A2 => n17471, ZN => n16322);
   U17364 : AOI22_X1 port map( A1 => n16323, A2 => n17565, B1 => n18539, B2 => 
                           n16322, ZN => n16324);
   U17365 : OAI21_X2 port map( B1 => n16325, B2 => n16789, A => n16324, ZN => 
                           n18568);
   U17366 : INV_X1 port map( A => n18568, ZN => n16446);
   U17367 : INV_X1 port map( A => n17276, ZN => n16326);
   U17368 : XNOR2_X1 port map( A => n19894, B => n16326, ZN => n16328);
   U17369 : XNOR2_X1 port map( A => n16931, B => n2395, ZN => n16327);
   U17370 : XNOR2_X1 port map( A => n16328, B => n16327, ZN => n16333);
   U17371 : XNOR2_X1 port map( A => n16329, B => n16971, ZN => n16885);
   U17372 : XNOR2_X1 port map( A => n16330, B => n16760, ZN => n16331);
   U17373 : INV_X1 port map( A => n16954, ZN => n16334);
   U17374 : XNOR2_X1 port map( A => n16334, B => n16335, ZN => n17268);
   U17375 : XNOR2_X1 port map( A => n17268, B => n16756, ZN => n16340);
   U17376 : XNOR2_X1 port map( A => n17111, B => n897, ZN => n16338);
   U17377 : XNOR2_X1 port map( A => n16893, B => n18801, ZN => n16337);
   U17378 : XNOR2_X1 port map( A => n16338, B => n16337, ZN => n16339);
   U17379 : NOR2_X1 port map( A1 => n20488, A2 => n18114, ZN => n18116);
   U17380 : XNOR2_X1 port map( A => n16342, B => n16341, ZN => n16346);
   U17381 : XNOR2_X1 port map( A => n17116, B => n17295, ZN => n16344);
   U17382 : XNOR2_X1 port map( A => n16965, B => n18065, ZN => n16343);
   U17383 : XNOR2_X1 port map( A => n16344, B => n16343, ZN => n16345);
   U17384 : XNOR2_X1 port map( A => n16346, B => n16345, ZN => n17458);
   U17385 : INV_X1 port map( A => n16347, ZN => n16599);
   U17386 : XNOR2_X1 port map( A => n16599, B => n16691, ZN => n16348);
   U17387 : XNOR2_X1 port map( A => n16348, B => n16906, ZN => n16352);
   U17388 : XNOR2_X1 port map( A => n16770, B => n16987, ZN => n16350);
   U17389 : XNOR2_X1 port map( A => n17098, B => n18517, ZN => n16349);
   U17390 : XNOR2_X1 port map( A => n16350, B => n16349, ZN => n16351);
   U17391 : OAI21_X1 port map( B1 => n18116, B2 => n17559, A => n18111, ZN => 
                           n16364);
   U17393 : XNOR2_X1 port map( A => n16553, B => n16353, ZN => n16357);
   U17394 : XNOR2_X1 port map( A => n16936, B => n2413, ZN => n16354);
   U17395 : XNOR2_X1 port map( A => n16355, B => n16354, ZN => n16356);
   U17397 : NOR2_X1 port map( A1 => n20488, A2 => n17458, ZN => n16363);
   U17398 : XNOR2_X1 port map( A => n20477, B => n16747, ZN => n16847);
   U17399 : XNOR2_X1 port map( A => n19743, B => n16914, ZN => n17258);
   U17400 : XNOR2_X1 port map( A => n17258, B => n16847, ZN => n16362);
   U17401 : XNOR2_X1 port map( A => n16996, B => n875, ZN => n16360);
   U17402 : XNOR2_X1 port map( A => n16878, B => n16360, ZN => n16361);
   U17403 : INV_X1 port map( A => n18556, ZN => n18199);
   U17404 : XNOR2_X1 port map( A => n16365, B => n16619, ZN => n16371);
   U17405 : XNOR2_X1 port map( A => n16615, B => n16961, ZN => n16369);
   U17406 : XNOR2_X1 port map( A => n16367, B => n16366, ZN => n16368);
   U17407 : XNOR2_X1 port map( A => n16369, B => n16368, ZN => n16370);
   U17408 : XNOR2_X1 port map( A => n16371, B => n16370, ZN => n17954);
   U17411 : XNOR2_X1 port map( A => n16373, B => n16374, ZN => n16834);
   U17412 : XNOR2_X1 port map( A => n17337, B => n16834, ZN => n16378);
   U17413 : XNOR2_X1 port map( A => n16954, B => n16695, ZN => n16376);
   U17414 : XNOR2_X1 port map( A => n16755, B => n2410, ZN => n16375);
   U17415 : XNOR2_X1 port map( A => n16376, B => n16375, ZN => n16377);
   U17416 : XNOR2_X1 port map( A => n16378, B => n16377, ZN => n17957);
   U17417 : OR2_X1 port map( A1 => n17954, A2 => n17957, ZN => n17552);
   U17418 : INV_X1 port map( A => n17552, ZN => n16389);
   U17419 : XNOR2_X1 port map( A => n16969, B => n2375, ZN => n16379);
   U17420 : XNOR2_X1 port map( A => n16380, B => n16379, ZN => n16382);
   U17421 : XNOR2_X1 port map( A => n16588, B => n16713, ZN => n16381);
   U17422 : XNOR2_X1 port map( A => n16381, B => n16382, ZN => n16805);
   U17423 : AND2_X1 port map( A1 => n18105, A2 => n17954, ZN => n16388);
   U17425 : XNOR2_X1 port map( A => n16385, B => n16384, ZN => n16387);
   U17426 : XNOR2_X1 port map( A => n16386, B => n17291, ZN => n16693);
   U17427 : OAI21_X1 port map( B1 => n16389, B2 => n16388, A => n18103, ZN => 
                           n16405);
   U17428 : INV_X1 port map( A => n18103, ZN => n16404);
   U17429 : XNOR2_X1 port map( A => n16510, B => n16608, ZN => n16391);
   U17430 : XNOR2_X1 port map( A => n16391, B => n16390, ZN => n16395);
   U17434 : XNOR2_X1 port map( A => n16596, B => n16396, ZN => n16400);
   U17435 : XNOR2_X1 port map( A => n15935, B => n17358, ZN => n16398);
   U17436 : XNOR2_X1 port map( A => n19889, B => n295, ZN => n16397);
   U17437 : XNOR2_X1 port map( A => n16398, B => n16397, ZN => n16399);
   U17438 : XNOR2_X1 port map( A => n16399, B => n16400, ZN => n17955);
   U17440 : NOR2_X1 port map( A1 => n17956, A2 => n18107, ZN => n16403);
   U17441 : AND2_X1 port map( A1 => n18107, A2 => n17957, ZN => n16402);
   U17442 : INV_X1 port map( A => n17954, ZN => n16401);
   U17443 : NAND2_X1 port map( A1 => n18199, A2 => n18559, ZN => n18201);
   U17444 : NAND2_X1 port map( A1 => n18199, A2 => n18568, ZN => n16453);
   U17445 : XNOR2_X1 port map( A => n20102, B => n16406, ZN => n17423);
   U17446 : XNOR2_X1 port map( A => n17423, B => n17036, ZN => n16411);
   U17447 : XNOR2_X1 port map( A => n16981, B => n17269, ZN => n16409);
   U17448 : XNOR2_X1 port map( A => n16836, B => n18366, ZN => n16408);
   U17449 : XNOR2_X1 port map( A => n16409, B => n16408, ZN => n16410);
   U17450 : INV_X1 port map( A => n18097, ZN => n18094);
   U17451 : XNOR2_X1 port map( A => n17019, B => n16527, ZN => n16416);
   U17452 : XNOR2_X1 port map( A => n20104, B => n16961, ZN => n16414);
   U17453 : XNOR2_X1 port map( A => n16412, B => n2307, ZN => n16413);
   U17454 : XNOR2_X1 port map( A => n16414, B => n16413, ZN => n16415);
   U17455 : XNOR2_X1 port map( A => n16416, B => n16415, ZN => n18096);
   U17456 : XNOR2_X1 port map( A => n17406, B => n18304, ZN => n16417);
   U17457 : XNOR2_X1 port map( A => n16417, B => n19820, ZN => n16419);
   U17458 : XNOR2_X1 port map( A => n17288, B => n17411, ZN => n16421);
   U17459 : XNOR2_X1 port map( A => n16421, B => n16420, ZN => n16519);
   U17461 : XNOR2_X1 port map( A => n16969, B => n16926, ZN => n16423);
   U17462 : XNOR2_X1 port map( A => n17026, B => n16423, ZN => n16428);
   U17463 : XNOR2_X1 port map( A => n17275, B => n16886, ZN => n16426);
   U17464 : XNOR2_X1 port map( A => n17279, B => n16424, ZN => n16425);
   U17465 : XOR2_X1 port map( A => n16426, B => n16425, Z => n16427);
   U17466 : NOR2_X1 port map( A1 => n18093, A2 => n20109, ZN => n16434);
   U17467 : XNOR2_X1 port map( A => n16429, B => n16872, ZN => n17420);
   U17468 : XNOR2_X1 port map( A => n16534, B => n17420, ZN => n16433);
   U17469 : XNOR2_X1 port map( A => n16554, B => n16706, ZN => n16431);
   U17470 : XNOR2_X1 port map( A => n17253, B => n18208, ZN => n16430);
   U17471 : XNOR2_X1 port map( A => n16431, B => n16430, ZN => n16432);
   U17472 : XNOR2_X1 port map( A => n16510, B => n16562, ZN => n16435);
   U17473 : XNOR2_X1 port map( A => n16514, B => n16435, ZN => n16439);
   U17474 : XNOR2_X1 port map( A => n16880, B => n17260, ZN => n16437);
   U17475 : XNOR2_X1 port map( A => n17378, B => n2221, ZN => n16436);
   U17476 : XNOR2_X1 port map( A => n16437, B => n16436, ZN => n16438);
   U17477 : XNOR2_X1 port map( A => n16439, B => n16438, ZN => n18101);
   U17478 : AND2_X1 port map( A1 => n18101, A2 => n160, ZN => n18099);
   U17479 : MUX2_X1 port map( A => n17164, B => n18099, S => n19774, Z => 
                           n16440);
   U17481 : NOR2_X1 port map( A1 => n19815, A2 => n19898, ZN => n16444);
   U17482 : NAND2_X1 port map( A1 => n19815, A2 => n16165, ZN => n16445);
   U17483 : NAND2_X1 port map( A1 => n18565, A2 => n18556, ZN => n16452);
   U17484 : OR2_X1 port map( A1 => n18567, A2 => n18199, ZN => n17997);
   U17485 : NAND2_X1 port map( A1 => n17495, A2 => n17493, ZN => n16449);
   U17486 : OAI21_X1 port map( B1 => n17491, B2 => n17155, A => n17488, ZN => 
                           n16448);
   U17487 : MUX2_X1 port map( A => n16449, B => n16448, S => n17489, Z => 
                           n16451);
   U17489 : INV_X1 port map( A => n2208, ZN => n16454);
   U17490 : NAND4_X1 port map( A1 => n16453, A2 => n19775, A3 => n16454, A4 => 
                           n16452, ZN => n16457);
   U17491 : NAND2_X1 port map( A1 => n18568, A2 => n16454, ZN => n16455);
   U17492 : OR2_X1 port map( A1 => n18201, A2 => n16455, ZN => n16456);
   U17493 : OAI211_X1 port map( C1 => n16459, C2 => n2208, A => n16457, B => 
                           n16456, ZN => n16458);
   U17494 : AOI21_X1 port map( B1 => n16460, B2 => n16459, A => n16458, ZN => 
                           Ciphertext(44));
   U17495 : NAND2_X1 port map( A1 => n17243, A2 => n17245, ZN => n16462);
   U17496 : NOR2_X1 port map( A1 => n17243, A2 => n17483, ZN => n17482);
   U17497 : MUX2_X1 port map( A => n17482, B => n16463, S => n17480, Z => 
                           n16464);
   U17499 : NAND2_X1 port map( A1 => n16660, A2 => n17208, ZN => n16466);
   U17501 : INV_X1 port map( A => n17511, ZN => n17512);
   U17502 : MUX2_X1 port map( A => n17512, B => n17508, S => n19956, Z => 
                           n16469);
   U17503 : INV_X1 port map( A => n20271, ZN => n17224);
   U17504 : MUX2_X1 port map( A => n17224, B => n17510, S => n19700, Z => 
                           n16468);
   U17505 : INV_X1 port map( A => n17493, ZN => n17154);
   U17506 : NOR2_X1 port map( A1 => n17154, A2 => n17489, ZN => n16470);
   U17507 : OAI21_X1 port map( B1 => n16470, B2 => n17490, A => n17491, ZN => 
                           n16473);
   U17508 : OAI21_X1 port map( B1 => n17488, B2 => n17489, A => n17493, ZN => 
                           n16471);
   U17509 : INV_X1 port map( A => n19814, ZN => n17502);
   U17510 : NAND3_X1 port map( A1 => n16794, A2 => n19898, A3 => n17502, ZN => 
                           n16478);
   U17511 : OAI21_X1 port map( B1 => n19815, B2 => n19924, A => n17505, ZN => 
                           n16477);
   U17512 : NAND2_X1 port map( A1 => n15485, A2 => n19924, ZN => n16476);
   U17513 : NAND3_X1 port map( A1 => n16478, A2 => n16477, A3 => n16476, ZN => 
                           n16479);
   U17515 : AOI21_X1 port map( B1 => n16666, B2 => n19386, A => n19382, ZN => 
                           n16483);
   U17516 : NOR2_X1 port map( A1 => n20463, A2 => n16665, ZN => n16481);
   U17517 : OAI21_X1 port map( B1 => n16641, B2 => n16481, A => n17220, ZN => 
                           n16482);
   U17518 : INV_X1 port map( A => n20232, ZN => n16484);
   U17519 : AOI22_X1 port map( A1 => n18469, A2 => n18464, B1 => n20148, B2 => 
                           n16484, ZN => n16485);
   U17520 : NAND2_X1 port map( A1 => n16486, A2 => n16485, ZN => n16489);
   U17521 : INV_X1 port map( A => n16487, ZN => n16488);
   U17522 : XNOR2_X1 port map( A => n16489, B => n16488, ZN => Ciphertext(18));
   U17523 : OAI21_X1 port map( B1 => n16491, B2 => n18406, A => n16490, ZN => 
                           n16493);
   U17524 : NOR2_X1 port map( A1 => n18425, A2 => n15529, ZN => n18409);
   U17525 : INV_X1 port map( A => n18427, ZN => n18407);
   U17526 : XNOR2_X1 port map( A => n16494, B => n2035, ZN => Ciphertext(15));
   U17528 : NAND2_X1 port map( A1 => n19402, A2 => n19401, ZN => n16495);
   U17529 : NAND2_X1 port map( A1 => n16497, A2 => n16495, ZN => n16496);
   U17530 : INV_X1 port map( A => n16497, ZN => n16499);
   U17531 : NOR2_X1 port map( A1 => n19401, A2 => n19403, ZN => n16498);
   U17532 : NAND2_X1 port map( A1 => n16499, A2 => n16498, ZN => n16500);
   U17533 : AND2_X2 port map( A1 => n16501, A2 => n16500, ZN => n19329);
   U17535 : NOR2_X1 port map( A1 => n20217, A2 => n19930, ZN => n16505);
   U17536 : MUX2_X1 port map( A => n16308, B => n17881, S => n17876, Z => 
                           n16503);
   U17537 : INV_X1 port map( A => n16503, ZN => n16504);
   U17538 : OAI21_X1 port map( B1 => n20162, B2 => n16505, A => n16504, ZN => 
                           n17539);
   U17539 : NAND2_X1 port map( A1 => n17539, A2 => n17610, ZN => n19333);
   U17540 : NOR2_X1 port map( A1 => n19749, A2 => n19333, ZN => n16581);
   U17541 : XNOR2_X1 port map( A => n20269, B => n16506, ZN => n16509);
   U17542 : INV_X1 port map( A => n2448, ZN => n18473);
   U17543 : XNOR2_X1 port map( A => n16507, B => n18473, ZN => n16508);
   U17544 : INV_X1 port map( A => n19363, ZN => n17863);
   U17545 : XNOR2_X1 port map( A => n16510, B => n17443, ZN => n16512);
   U17546 : XNOR2_X1 port map( A => n16750, B => n17804, ZN => n16511);
   U17547 : XNOR2_X1 port map( A => n16512, B => n16511, ZN => n16516);
   U17548 : XNOR2_X1 port map( A => n16514, B => n16513, ZN => n16515);
   U17549 : XNOR2_X1 port map( A => n16515, B => n16516, ZN => n16679);
   U17550 : INV_X1 port map( A => n16679, ZN => n19361);
   U17551 : XNOR2_X1 port map( A => n16992, B => n632, ZN => n16517);
   U17552 : MUX2_X1 port map( A => n17863, B => n19361, S => n17861, Z => 
                           n16539);
   U17553 : XNOR2_X1 port map( A => n19849, B => n16521, ZN => n16526);
   U17554 : XNOR2_X1 port map( A => n17133, B => n2446, ZN => n16524);
   U17555 : XNOR2_X1 port map( A => n16523, B => n16524, ZN => n16525);
   U17556 : NOR2_X1 port map( A1 => n19362, A2 => n19938, ZN => n17591);
   U17557 : XNOR2_X1 port map( A => n16528, B => n16527, ZN => n16532);
   U17558 : XNOR2_X1 port map( A => n17294, B => n16963, ZN => n16530);
   U17559 : XNOR2_X1 port map( A => n17330, B => n484, ZN => n16529);
   U17560 : XNOR2_X1 port map( A => n16530, B => n16529, ZN => n16531);
   U17561 : XNOR2_X1 port map( A => n16532, B => n16531, ZN => n17672);
   U17562 : AND2_X1 port map( A1 => n19363, A2 => n17672, ZN => n17592);
   U17563 : NOR2_X1 port map( A1 => n17591, A2 => n17592, ZN => n16538);
   U17564 : XNOR2_X1 port map( A => n16938, B => n2082, ZN => n16533);
   U17565 : XNOR2_X1 port map( A => n16937, B => n16533, ZN => n16537);
   U17566 : XNOR2_X1 port map( A => n20267, B => n17002, ZN => n16535);
   U17567 : XNOR2_X1 port map( A => n16535, B => n16534, ZN => n16536);
   U17569 : MUX2_X2 port map( A => n16539, B => n16538, S => n19360, Z => 
                           n19340);
   U17570 : INV_X1 port map( A => n19340, ZN => n16544);
   U17572 : NOR2_X1 port map( A1 => n16636, A2 => n19351, ZN => n16543);
   U17573 : NAND2_X1 port map( A1 => n16672, A2 => n19347, ZN => n17231);
   U17574 : NAND2_X1 port map( A1 => n17234, A2 => n17231, ZN => n16541);
   U17577 : XNOR2_X1 port map( A => n17338, B => n17060, ZN => n16545);
   U17578 : XNOR2_X1 port map( A => n16696, B => n16545, ZN => n16548);
   U17579 : XNOR2_X1 port map( A => n16892, B => n16546, ZN => n16547);
   U17580 : XNOR2_X1 port map( A => n16548, B => n16547, ZN => n16642);
   U17581 : XNOR2_X1 port map( A => n16719, B => n16898, ZN => n16552);
   U17582 : XNOR2_X1 port map( A => n20104, B => n17116, ZN => n16550);
   U17583 : XNOR2_X1 port map( A => n16614, B => n18338, ZN => n16549);
   U17584 : XNOR2_X1 port map( A => n16550, B => n16549, ZN => n16551);
   U17585 : XNOR2_X2 port map( A => n16552, B => n16551, ZN => n19372);
   U17586 : XNOR2_X1 port map( A => n16705, B => n16553, ZN => n16559);
   U17587 : XNOR2_X1 port map( A => n16554, B => n20450, ZN => n16557);
   U17588 : XNOR2_X1 port map( A => n16593, B => n302, ZN => n16556);
   U17589 : XNOR2_X1 port map( A => n16557, B => n16556, ZN => n16558);
   U17590 : INV_X1 port map( A => n19371, ZN => n19375);
   U17591 : OAI21_X1 port map( B1 => n20436, B2 => n19372, A => n19375, ZN => 
                           n16657);
   U17592 : INV_X1 port map( A => Key(60), ZN => n16560);
   U17593 : XNOR2_X1 port map( A => n20478, B => n16560, ZN => n16561);
   U17594 : XNOR2_X1 port map( A => n16702, B => n16561, ZN => n16565);
   U17595 : XNOR2_X1 port map( A => n16562, B => n16607, ZN => n16563);
   U17596 : XNOR2_X1 port map( A => n16563, B => n16882, ZN => n16564);
   U17597 : XNOR2_X1 port map( A => n16565, B => n16564, ZN => n19374);
   U17598 : NAND2_X1 port map( A1 => n19374, A2 => n19666, ZN => n16579);
   U17599 : XNOR2_X1 port map( A => n19894, B => n16566, ZN => n16859);
   U17600 : XNOR2_X1 port map( A => n16859, B => n16567, ZN => n16572);
   U17601 : XNOR2_X1 port map( A => n16587, B => n16568, ZN => n16570);
   U17602 : XNOR2_X1 port map( A => n17279, B => n18070, ZN => n16569);
   U17603 : XNOR2_X1 port map( A => n16570, B => n16569, ZN => n16571);
   U17604 : XNOR2_X1 port map( A => n16572, B => n16571, ZN => n19370);
   U17606 : XNOR2_X1 port map( A => n16601, B => n16573, ZN => n16575);
   U17607 : XNOR2_X1 port map( A => n16574, B => n16575, ZN => n16576);
   U17608 : OAI21_X1 port map( B1 => n16581, B2 => n19315, A => n19338, ZN => 
                           n16623);
   U17609 : XNOR2_X1 port map( A => n16835, B => n20494, ZN => n16586);
   U17610 : XNOR2_X1 port map( A => n19927, B => n19243, ZN => n16583);
   U17611 : XNOR2_X1 port map( A => n16584, B => n16583, ZN => n16585);
   U17612 : XNOR2_X1 port map( A => n17367, B => n16587, ZN => n17029);
   U17613 : XNOR2_X1 port map( A => n17029, B => n16588, ZN => n16592);
   U17614 : XNOR2_X1 port map( A => n17280, B => n16760, ZN => n16590);
   U17615 : XNOR2_X1 port map( A => n16927, B => n2344, ZN => n16589);
   U17616 : XNOR2_X1 port map( A => n16590, B => n16589, ZN => n16591);
   U17617 : XNOR2_X1 port map( A => n16592, B => n16591, ZN => n17656);
   U17618 : XNOR2_X1 port map( A => n16938, B => n18716, ZN => n16595);
   U17619 : XNOR2_X1 port map( A => n16593, B => n16741, ZN => n16594);
   U17620 : XNOR2_X1 port map( A => n16595, B => n16594, ZN => n16598);
   U17621 : XNOR2_X1 port map( A => n17040, B => n16596, ZN => n16597);
   U17622 : XNOR2_X1 port map( A => n16599, B => n17012, ZN => n17286);
   U17623 : XNOR2_X1 port map( A => n17286, B => n16829, ZN => n16605);
   U17624 : XNOR2_X1 port map( A => n16600, B => n16601, ZN => n17345);
   U17625 : XNOR2_X1 port map( A => n16602, B => n2203, ZN => n16603);
   U17626 : XNOR2_X1 port map( A => n17345, B => n16603, ZN => n16604);
   U17627 : XNOR2_X1 port map( A => n16605, B => n16604, ZN => n19388);
   U17628 : AOI21_X1 port map( B1 => n17656, B2 => n20172, A => n19388, ZN => 
                           n16606);
   U17629 : NAND2_X1 port map( A1 => n16683, A2 => n16606, ZN => n17537);
   U17630 : XNOR2_X1 port map( A => n16608, B => n16607, ZN => n17376);
   U17631 : XNOR2_X1 port map( A => n19900, B => n16914, ZN => n16609);
   U17632 : XNOR2_X1 port map( A => n17376, B => n16609, ZN => n16613);
   U17633 : XNOR2_X1 port map( A => n16844, B => n17443, ZN => n16611);
   U17634 : XNOR2_X1 port map( A => n17260, B => n20593, ZN => n16610);
   U17635 : XNOR2_X1 port map( A => n16611, B => n16610, ZN => n16612);
   U17636 : XNOR2_X1 port map( A => n16613, B => n16612, ZN => n17654);
   U17637 : XNOR2_X1 port map( A => n16615, B => n16614, ZN => n17325);
   U17638 : XNOR2_X1 port map( A => n16944, B => n19457, ZN => n16616);
   U17639 : XNOR2_X1 port map( A => n17325, B => n16616, ZN => n16621);
   U17640 : INV_X1 port map( A => n16617, ZN => n16618);
   U17641 : XNOR2_X1 port map( A => n16618, B => n16619, ZN => n16620);
   U17642 : XNOR2_X1 port map( A => n16620, B => n16621, ZN => n19390);
   U17644 : INV_X1 port map( A => n19396, ZN => n19391);
   U17645 : NAND3_X1 port map( A1 => n19511, A2 => n19391, A3 => n20172, ZN => 
                           n17536);
   U17646 : AND2_X1 port map( A1 => n19329, A2 => n18311, ZN => n17542);
   U17647 : OAI21_X1 port map( B1 => n17542, B2 => n19333, A => n19340, ZN => 
                           n16622);
   U17648 : NAND2_X1 port map( A1 => n16623, A2 => n16622, ZN => n16625);
   U17649 : INV_X1 port map( A => n106, ZN => n16624);
   U17650 : XNOR2_X1 port map( A => n16625, B => n16624, ZN => Ciphertext(179))
                           ;
   U17651 : MUX2_X1 port map( A => n16629, B => n20092, S => n17210, Z => 
                           n16628);
   U17652 : NOR2_X1 port map( A1 => n19975, A2 => n17208, ZN => n16627);
   U17653 : NOR3_X1 port map( A1 => n20092, A2 => n16629, A3 => n20135, ZN => 
                           n16630);
   U17654 : INV_X1 port map( A => n17508, ZN => n17513);
   U17655 : NOR2_X1 port map( A1 => n16632, A2 => n17513, ZN => n18340);
   U17656 : NOR2_X1 port map( A1 => n18340, A2 => n18342, ZN => n18287);
   U17657 : NOR2_X1 port map( A1 => n18365, A2 => n18362, ZN => n18286);
   U17660 : NOR2_X1 port map( A1 => n19382, A2 => n16666, ZN => n16640);
   U17661 : AOI22_X1 port map( A1 => n16641, A2 => n19386, B1 => n16640, B2 => 
                           n1897, ZN => n18341);
   U17663 : INV_X1 port map( A => n18290, ZN => n18292);
   U17664 : INV_X1 port map( A => n19374, ZN => n17240);
   U17665 : NAND2_X1 port map( A1 => n17240, A2 => n19666, ZN => n16654);
   U17666 : INV_X1 port map( A => n16642, ZN => n19373);
   U17668 : NAND3_X1 port map( A1 => n16654, A2 => n19373, A3 => n19647, ZN => 
                           n17906);
   U17669 : MUX2_X1 port map( A => n17656, B => n19390, S => n19396, Z => 
                           n16643);
   U17670 : INV_X1 port map( A => n16643, ZN => n16647);
   U17671 : OAI21_X1 port map( B1 => n19388, B2 => n17654, A => n20004, ZN => 
                           n16646);
   U17672 : INV_X1 port map( A => n17654, ZN => n16644);
   U17673 : NOR2_X1 port map( A1 => n16644, A2 => n19396, ZN => n16645);
   U17674 : AOI21_X2 port map( B1 => n16647, B2 => n16646, A => n16645, ZN => 
                           n18359);
   U17675 : OAI211_X1 port map( C1 => n18292, C2 => n18358, A => n18357, B => 
                           n18359, ZN => n16648);
   U17676 : OAI21_X1 port map( B1 => n18286, B2 => n18357, A => n16648, ZN => 
                           n16650);
   U17677 : INV_X1 port map( A => n18358, ZN => n18348);
   U17678 : NAND2_X1 port map( A1 => n18348, A2 => n18359, ZN => n17907);
   U17679 : NAND2_X1 port map( A1 => n16650, A2 => n16649, ZN => n16653);
   U17680 : INV_X1 port map( A => n16651, ZN => n16652);
   U17681 : XNOR2_X1 port map( A => n16653, B => n16652, ZN => Ciphertext(5));
   U17682 : AND2_X1 port map( A1 => n19370, A2 => n16642, ZN => n17596);
   U17683 : NAND2_X1 port map( A1 => n19373, A2 => n19666, ZN => n16655);
   U17684 : MUX2_X1 port map( A => n16655, B => n16654, S => n19733, Z => 
                           n16656);
   U17685 : NAND2_X1 port map( A1 => n16658, A2 => n17208, ZN => n16659);
   U17687 : NAND2_X1 port map( A1 => n16661, A2 => n20092, ZN => n16664);
   U17688 : NAND2_X1 port map( A1 => n16662, A2 => n17213, ZN => n16663);
   U17689 : NOR2_X1 port map( A1 => n19385, A2 => n17220, ZN => n16667);
   U17690 : AND2_X1 port map( A1 => n16665, A2 => n19382, ZN => n16668);
   U17691 : MUX2_X1 port map( A => n16667, B => n16668, S => n3389, Z => n16671
                           );
   U17692 : OAI21_X1 port map( B1 => n20463, B2 => n19382, A => n19385, ZN => 
                           n16669);
   U17693 : NOR2_X1 port map( A1 => n16669, A2 => n16668, ZN => n16670);
   U17694 : NOR2_X2 port map( A1 => n16671, A2 => n16670, ZN => n19459);
   U17695 : MUX2_X1 port map( A => n19349, B => n19353, S => n16672, Z => 
                           n16677);
   U17696 : INV_X1 port map( A => n20240, ZN => n16676);
   U17697 : NAND3_X1 port map( A1 => n19349, A2 => n19353, A3 => n19351, ZN => 
                           n16675);
   U17698 : INV_X1 port map( A => n18067, ZN => n19462);
   U17699 : NAND2_X1 port map( A1 => n19361, A2 => n19360, ZN => n17595);
   U17700 : NAND2_X1 port map( A1 => n17595, A2 => n20242, ZN => n16681);
   U17701 : NAND2_X1 port map( A1 => n17861, A2 => n19360, ZN => n19365);
   U17702 : NAND2_X1 port map( A1 => n20212, A2 => n19938, ZN => n16678);
   U17703 : NAND2_X1 port map( A1 => n19365, A2 => n16678, ZN => n16680);
   U17704 : NAND3_X1 port map( A1 => n19462, A2 => n19460, A3 => n19453, ZN => 
                           n16682);
   U17705 : INV_X1 port map( A => n16683, ZN => n16687);
   U17706 : INV_X1 port map( A => n16684, ZN => n16686);
   U17707 : NAND2_X1 port map( A1 => n19390, A2 => n17656, ZN => n16685);
   U17708 : INV_X1 port map( A => n19453, ZN => n17091);
   U17709 : INV_X1 port map( A => n457, ZN => n16688);
   U17710 : XNOR2_X1 port map( A => n16689, B => n17347, ZN => n16692);
   U17711 : XNOR2_X1 port map( A => n16691, B => n16690, ZN => n17287);
   U17712 : XNOR2_X1 port map( A => n17287, B => n16692, ZN => n16694);
   U17714 : XNOR2_X1 port map( A => n19909, B => n16695, ZN => n16895);
   U17715 : XNOR2_X1 port map( A => n936, B => n16895, ZN => n16700);
   U17716 : XNOR2_X1 port map( A => n17339, B => n17269, ZN => n16698);
   U17717 : XNOR2_X1 port map( A => n16755, B => n1386, ZN => n16697);
   U17718 : XNOR2_X1 port map( A => n16698, B => n16697, ZN => n16699);
   U17719 : XNOR2_X1 port map( A => n16700, B => n16699, ZN => n17193);
   U17720 : XNOR2_X1 port map( A => n16844, B => n17442, ZN => n16879);
   U17721 : XNOR2_X1 port map( A => n17259, B => n16879, ZN => n16704);
   U17722 : XNOR2_X1 port map( A => n17378, B => n106, ZN => n16701);
   U17723 : XNOR2_X1 port map( A => n16702, B => n16701, ZN => n16703);
   U17724 : MUX2_X1 port map( A => n19684, B => n935, S => n18966, Z => n16726)
                           ;
   U17725 : XNOR2_X1 port map( A => n16705, B => n17250, ZN => n16710);
   U17726 : XNOR2_X1 port map( A => n16706, B => n18006, ZN => n16708);
   U17727 : XNOR2_X1 port map( A => n20167, B => n16707, ZN => n16870);
   U17728 : XNOR2_X1 port map( A => n16708, B => n16870, ZN => n16709);
   U17730 : XNOR2_X1 port map( A => n17276, B => n16711, ZN => n16712);
   U17731 : XNOR2_X1 port map( A => n16713, B => n16712, ZN => n16717);
   U17732 : XNOR2_X1 port map( A => n16861, B => n17433, ZN => n16715);
   U17733 : XNOR2_X1 port map( A => n17279, B => n311, ZN => n16714);
   U17734 : XNOR2_X1 port map( A => n16715, B => n16714, ZN => n16716);
   U17735 : XNOR2_X1 port map( A => n16717, B => n16716, ZN => n17695);
   U17736 : NOR2_X1 port map( A1 => n18966, A2 => n17695, ZN => n16718);
   U17737 : NAND2_X1 port map( A1 => n16718, A2 => n17819, ZN => n16724);
   U17738 : XNOR2_X1 port map( A => n17401, B => n19720, ZN => n16899);
   U17739 : XNOR2_X1 port map( A => n16719, B => n16899, ZN => n16723);
   U17740 : XNOR2_X1 port map( A => n20104, B => n17294, ZN => n16721);
   U17741 : XNOR2_X1 port map( A => n20125, B => n1904, ZN => n16720);
   U17742 : XNOR2_X1 port map( A => n16721, B => n16720, ZN => n16722);
   U17744 : NAND2_X1 port map( A1 => n18961, A2 => n935, ZN => n18970);
   U17745 : NAND2_X1 port map( A1 => n16724, A2 => n18970, ZN => n16725);
   U17746 : AOI22_X1 port map( A1 => n20506, A2 => n17676, B1 => n17867, B2 => 
                           n20514, ZN => n16727);
   U17747 : NOR2_X1 port map( A1 => n16727, A2 => n19973, ZN => n16729);
   U17748 : AND2_X1 port map( A1 => n17873, A2 => n17872, ZN => n17677);
   U17752 : NOR2_X1 port map( A1 => n17840, A2 => n17835, ZN => n17062);
   U17753 : INV_X1 port map( A => n17062, ZN => n16732);
   U17755 : XNOR2_X1 port map( A => n17294, B => n16900, ZN => n16735);
   U17756 : XNOR2_X1 port map( A => n16851, B => n16735, ZN => n16739);
   U17757 : XNOR2_X1 port map( A => n16960, B => n20481, ZN => n16737);
   U17758 : XNOR2_X1 port map( A => n16854, B => n18854, ZN => n16736);
   U17759 : XNOR2_X1 port map( A => n16737, B => n16736, ZN => n16738);
   U17760 : XNOR2_X1 port map( A => n16739, B => n16738, ZN => n18955);
   U17761 : INV_X1 port map( A => n18955, ZN => n16745);
   U17762 : XNOR2_X1 port map( A => n19889, B => n16741, ZN => n16825);
   U17763 : XNOR2_X1 port map( A => n20267, B => n16742, ZN => n16744);
   U17764 : NOR2_X1 port map( A1 => n16745, A2 => n17831, ZN => n16767);
   U17765 : XNOR2_X1 port map( A => n19900, B => n20100, ZN => n16748);
   U17766 : XNOR2_X1 port map( A => n16749, B => n16748, ZN => n16754);
   U17767 : XNOR2_X1 port map( A => n16840, B => n16750, ZN => n16752);
   U17768 : INV_X1 port map( A => n2341, ZN => n19083);
   U17769 : XNOR2_X1 port map( A => n16996, B => n19083, ZN => n16751);
   U17770 : XNOR2_X1 port map( A => n16752, B => n16751, ZN => n16753);
   U17771 : XNOR2_X1 port map( A => n16754, B => n16753, ZN => n18953);
   U17772 : INV_X1 port map( A => n18953, ZN => n17179);
   U17773 : XNOR2_X1 port map( A => n16757, B => n16756, ZN => n16759);
   U17774 : AOI21_X1 port map( B1 => n2907, B2 => n17179, A => n18954, ZN => 
                           n16766);
   U17775 : XNOR2_X1 port map( A => n16761, B => n16760, ZN => n16860);
   U17776 : XNOR2_X1 port map( A => n16970, B => n16971, ZN => n16763);
   U17777 : XNOR2_X1 port map( A => n20098, B => n2263, ZN => n16762);
   U17778 : XNOR2_X1 port map( A => n16763, B => n16762, ZN => n16764);
   U17779 : XNOR2_X1 port map( A => n16765, B => n16764, ZN => n17180);
   U17780 : INV_X1 port map( A => n17180, ZN => n18959);
   U17781 : MUX2_X1 port map( A => n16767, B => n16766, S => n18959, Z => 
                           n16776);
   U17782 : XNOR2_X1 port map( A => n16987, B => n2035, ZN => n16768);
   U17783 : XNOR2_X1 port map( A => n16769, B => n16768, ZN => n16774);
   U17784 : XNOR2_X1 port map( A => n17291, B => n16770, ZN => n16771);
   U17785 : XNOR2_X1 port map( A => n16771, B => n16772, ZN => n16773);
   U17786 : NAND2_X1 port map( A1 => n18956, A2 => n17831, ZN => n17833);
   U17787 : INV_X1 port map( A => n17833, ZN => n16775);
   U17788 : NOR2_X2 port map( A1 => n16776, A2 => n16775, ZN => n19134);
   U17789 : MUX2_X1 port map( A => n17079, B => n20239, S => n17823, Z => 
                           n16778);
   U17790 : INV_X1 port map( A => n17825, ZN => n17176);
   U17791 : NOR2_X1 port map( A1 => n19135, A2 => n16780, ZN => n19147);
   U17792 : INV_X1 port map( A => n19134, ZN => n19145);
   U17794 : OR2_X1 port map( A1 => n17898, A2 => n19707, ZN => n16787);
   U17795 : NAND2_X1 port map( A1 => n19910, A2 => n16025, ZN => n16785);
   U17796 : NAND2_X1 port map( A1 => n16785, A2 => n17892, ZN => n16786);
   U17797 : AND2_X1 port map( A1 => n17564, A2 => n20432, ZN => n17161);
   U17798 : OAI21_X1 port map( B1 => n17471, B2 => n20432, A => n18539, ZN => 
                           n16792);
   U17799 : NAND2_X1 port map( A1 => n16789, A2 => n18535, ZN => n18542);
   U17801 : NAND2_X1 port map( A1 => n16790, A2 => n18538, ZN => n16791);
   U17802 : OAI21_X1 port map( B1 => n17504, B2 => n16165, A => n1060, ZN => 
                           n16799);
   U17803 : NAND2_X1 port map( A1 => n16795, A2 => n16794, ZN => n16796);
   U17804 : NAND2_X1 port map( A1 => n16797, A2 => n16796, ZN => n16798);
   U17805 : NAND2_X1 port map( A1 => n16799, A2 => n16798, ZN => n18545);
   U17806 : NOR2_X1 port map( A1 => n17584, A2 => n18545, ZN => n18530);
   U17807 : NOR2_X1 port map( A1 => n16801, A2 => n17155, ZN => n16804);
   U17808 : NOR2_X1 port map( A1 => n18530, A2 => n19691, ZN => n16807);
   U17810 : NAND2_X1 port map( A1 => n19682, A2 => n18545, ZN => n16806);
   U17811 : NAND2_X1 port map( A1 => n16807, A2 => n16806, ZN => n16818);
   U17812 : OAI21_X1 port map( B1 => n17243, B2 => n17245, A => n17479, ZN => 
                           n16808);
   U17813 : NAND2_X1 port map( A1 => n16809, A2 => n16808, ZN => n18540);
   U17814 : NAND2_X1 port map( A1 => n18540, A2 => n18541, ZN => n17925);
   U17815 : NAND3_X1 port map( A1 => n17923, A2 => n19682, A3 => n17925, ZN => 
                           n16817);
   U17816 : MUX2_X1 port map( A => n18093, B => n160, S => n18097, Z => n16812)
                           ;
   U17817 : INV_X1 port map( A => n18093, ZN => n17475);
   U17818 : NOR2_X1 port map( A1 => n17475, A2 => n18095, ZN => n16811);
   U17819 : MUX2_X1 port map( A => n16812, B => n16811, S => n18096, Z => 
                           n16815);
   U17820 : NAND2_X1 port map( A1 => n18101, A2 => n226, ZN => n16813);
   U17821 : NOR2_X1 port map( A1 => n16813, A2 => n19774, ZN => n16814);
   U17822 : NAND3_X1 port map( A1 => n16818, A2 => n16817, A3 => n16816, ZN => 
                           n16820);
   U17823 : INV_X1 port map( A => n2337, ZN => n16819);
   U17824 : XNOR2_X1 port map( A => n16820, B => n16819, ZN => Ciphertext(39));
   U17825 : XNOR2_X1 port map( A => n16821, B => n16742, ZN => n16823);
   U17826 : XNOR2_X1 port map( A => n16823, B => n16822, ZN => n16827);
   U17827 : XNOR2_X1 port map( A => n19845, B => n610, ZN => n16824);
   U17828 : XOR2_X1 port map( A => n16825, B => n16824, Z => n16826);
   U17829 : XNOR2_X1 port map( A => n16829, B => n16828, ZN => n16833);
   U17830 : XNOR2_X1 port map( A => n16188, B => n17098, ZN => n16831);
   U17831 : XNOR2_X1 port map( A => n17288, B => n2424, ZN => n16830);
   U17832 : XNOR2_X1 port map( A => n16831, B => n16830, ZN => n16832);
   U17834 : XNOR2_X1 port map( A => n16835, B => n16834, ZN => n16839);
   U17835 : XNOR2_X1 port map( A => n17111, B => n16836, ZN => n17032);
   U17836 : XNOR2_X1 port map( A => n17110, B => n18078, ZN => n16837);
   U17837 : XNOR2_X1 port map( A => n17032, B => n16837, ZN => n16838);
   U17838 : XNOR2_X2 port map( A => n16839, B => n16838, ZN => n18275);
   U17839 : XNOR2_X1 port map( A => n17124, B => n16840, ZN => n16843);
   U17840 : XNOR2_X1 port map( A => n19704, B => n2306, ZN => n16842);
   U17841 : XNOR2_X1 port map( A => n16843, B => n16842, ZN => n16849);
   U17842 : INV_X1 port map( A => n16844, ZN => n16845);
   U17843 : XNOR2_X1 port map( A => n16845, B => n947, ZN => n16846);
   U17844 : XNOR2_X1 port map( A => n16847, B => n16846, ZN => n16848);
   U17845 : XNOR2_X1 port map( A => n19720, B => n17116, ZN => n16852);
   U17846 : XNOR2_X1 port map( A => n16851, B => n16852, ZN => n16858);
   U17847 : XNOR2_X1 port map( A => n16853, B => n19929, ZN => n16856);
   U17848 : XNOR2_X1 port map( A => n16854, B => n2233, ZN => n16855);
   U17849 : XNOR2_X1 port map( A => n16856, B => n16855, ZN => n16857);
   U17850 : XNOR2_X1 port map( A => n16858, B => n16857, ZN => n18273);
   U17851 : INV_X1 port map( A => n18269, ZN => n16866);
   U17852 : XNOR2_X1 port map( A => n16859, B => n16860, ZN => n16865);
   U17853 : XNOR2_X1 port map( A => n879, B => n17275, ZN => n16863);
   U17854 : XNOR2_X1 port map( A => n16861, B => n18177, ZN => n16862);
   U17855 : XNOR2_X1 port map( A => n16863, B => n16862, ZN => n16864);
   U17856 : XNOR2_X1 port map( A => n16865, B => n16864, ZN => n17769);
   U17857 : NAND2_X1 port map( A1 => n16866, A2 => n17769, ZN => n16867);
   U17858 : MUX2_X1 port map( A => n221, B => n16867, S => n18275, Z => n16868)
                           ;
   U17859 : XNOR2_X1 port map( A => n16871, B => n16870, ZN => n16877);
   U17860 : XNOR2_X1 port map( A => n17005, B => n16872, ZN => n16875);
   U17861 : XNOR2_X1 port map( A => n16873, B => n18170, ZN => n16874);
   U17862 : XNOR2_X1 port map( A => n16875, B => n16874, ZN => n16876);
   U17864 : XNOR2_X1 port map( A => n16878, B => n16879, ZN => n16884);
   U17865 : XNOR2_X1 port map( A => n16880, B => n18396, ZN => n16881);
   U17866 : XNOR2_X1 port map( A => n16882, B => n16881, ZN => n16883);
   U17867 : XNOR2_X1 port map( A => n16884, B => n16883, ZN => n18016);
   U17868 : AND2_X1 port map( A1 => n20129, A2 => n18016, ZN => n16913);
   U17869 : XNOR2_X1 port map( A => n16885, B => n17135, ZN => n16890);
   U17870 : XNOR2_X1 port map( A => n16886, B => Key(63), ZN => n16888);
   U17871 : XNOR2_X1 port map( A => n16887, B => n16888, ZN => n16889);
   U17872 : XNOR2_X1 port map( A => n16892, B => n16891, ZN => n16897);
   U17873 : XNOR2_X1 port map( A => n16893, B => n1840, ZN => n16894);
   U17874 : XNOR2_X1 port map( A => n16895, B => n16894, ZN => n16896);
   U17875 : NAND2_X1 port map( A1 => n20158, A2 => n20499, ZN => n16912);
   U17876 : XNOR2_X1 port map( A => n16898, B => n16899, ZN => n16904);
   U17877 : XNOR2_X1 port map( A => n16900, B => n19321, ZN => n16901);
   U17878 : XNOR2_X1 port map( A => n16902, B => n16901, ZN => n16903);
   U17879 : NOR2_X1 port map( A1 => n18976, A2 => n18975, ZN => n18223);
   U17880 : XNOR2_X1 port map( A => n16905, B => n16906, ZN => n16910);
   U17881 : XNOR2_X1 port map( A => n16908, B => n16907, ZN => n16909);
   U17882 : XNOR2_X1 port map( A => n17379, B => n2108, ZN => n16915);
   U17883 : XNOR2_X1 port map( A => n16915, B => n16914, ZN => n16917);
   U17884 : XNOR2_X1 port map( A => n17443, B => n955, ZN => n16916);
   U17885 : XNOR2_X1 port map( A => n16917, B => n16916, ZN => n16920);
   U17886 : XNOR2_X1 port map( A => n17438, B => n16918, ZN => n16919);
   U17887 : XNOR2_X1 port map( A => n16920, B => n16919, ZN => n18042);
   U17888 : XNOR2_X1 port map( A => n19836, B => n2323, ZN => n16923);
   U17889 : XNOR2_X1 port map( A => n16921, B => n19713, ZN => n16922);
   U17890 : XNOR2_X1 port map( A => n16923, B => n16922, ZN => n16925);
   U17891 : XNOR2_X1 port map( A => n16988, B => n17409, ZN => n16924);
   U17892 : XNOR2_X1 port map( A => n16925, B => n16924, ZN => n18043);
   U17893 : NAND2_X1 port map( A1 => n20194, A2 => n19916, ZN => n18950);
   U17894 : XNOR2_X1 port map( A => n16927, B => n16926, ZN => n17432);
   U17895 : XNOR2_X1 port map( A => n16929, B => n16928, ZN => n16930);
   U17896 : XNOR2_X1 port map( A => n16930, B => n17432, ZN => n16935);
   U17897 : XNOR2_X1 port map( A => n16931, B => n17366, ZN => n17278);
   U17898 : XNOR2_X1 port map( A => n16932, B => n17851, ZN => n16933);
   U17899 : XNOR2_X1 port map( A => n17278, B => n16933, ZN => n16934);
   U17900 : XNOR2_X1 port map( A => n17360, B => n16936, ZN => n17249);
   U17901 : XNOR2_X1 port map( A => n19863, B => n17249, ZN => n16943);
   U17902 : XNOR2_X1 port map( A => n16938, B => n19180, ZN => n16941);
   U17903 : XNOR2_X1 port map( A => n16939, B => n16181, ZN => n16940);
   U17904 : XNOR2_X1 port map( A => n16941, B => n16940, ZN => n16942);
   U17905 : XNOR2_X2 port map( A => n16943, B => n16942, ZN => n18946);
   U17906 : XNOR2_X1 port map( A => n16945, B => n16944, ZN => n17403);
   U17907 : XNOR2_X1 port map( A => n17403, B => n16946, ZN => n16951);
   U17908 : XNOR2_X1 port map( A => n16947, B => n17295, ZN => n16949);
   U17909 : XNOR2_X1 port map( A => n17330, B => n2284, ZN => n16948);
   U17910 : XNOR2_X1 port map( A => n16949, B => n16948, ZN => n16950);
   U17911 : XNOR2_X1 port map( A => n16951, B => n16950, ZN => n18046);
   U17913 : NAND2_X1 port map( A1 => n2586, A2 => n18946, ZN => n16959);
   U17914 : XNOR2_X1 port map( A => n16952, B => n16953, ZN => n16958);
   U17915 : XNOR2_X1 port map( A => n16954, B => n19706, ZN => n16956);
   U17916 : XNOR2_X1 port map( A => n902, B => n17932, ZN => n16955);
   U17917 : XNOR2_X1 port map( A => n16956, B => n16955, ZN => n16957);
   U17918 : NAND2_X1 port map( A1 => n19681, A2 => n17054, ZN => n18891);
   U17919 : OAI21_X1 port map( B1 => n19905, B2 => n18897, A => n18891, ZN => 
                           n17059);
   U17920 : XNOR2_X1 port map( A => n16961, B => n16960, ZN => n17326);
   U17921 : XNOR2_X1 port map( A => n16962, B => n17326, ZN => n16968);
   U17922 : XNOR2_X1 port map( A => n16964, B => n16963, ZN => n17118);
   U17923 : XNOR2_X1 port map( A => n20481, B => n2384, ZN => n16966);
   U17924 : XNOR2_X1 port map( A => n17118, B => n16966, ZN => n16967);
   U17925 : XNOR2_X1 port map( A => n16967, B => n16968, ZN => n18029);
   U17926 : INV_X1 port map( A => n18029, ZN => n18926);
   U17927 : XNOR2_X1 port map( A => n16970, B => n16969, ZN => n17370);
   U17928 : XNOR2_X1 port map( A => n17133, B => n16971, ZN => n16972);
   U17929 : XNOR2_X1 port map( A => n17370, B => n16972, ZN => n16978);
   U17930 : XNOR2_X1 port map( A => n19659, B => n16973, ZN => n17139);
   U17931 : XNOR2_X1 port map( A => n16975, B => n17544, ZN => n16976);
   U17932 : XNOR2_X1 port map( A => n17139, B => n16976, ZN => n16977);
   U17933 : XNOR2_X1 port map( A => n16978, B => n16977, ZN => n18024);
   U17934 : XNOR2_X1 port map( A => n17108, B => n16979, ZN => n16986);
   U17935 : XNOR2_X1 port map( A => n16981, B => n16980, ZN => n16984);
   U17936 : XNOR2_X1 port map( A => n16982, B => n18830, ZN => n16983);
   U17937 : XNOR2_X1 port map( A => n16984, B => n16983, ZN => n16985);
   U17939 : MUX2_X1 port map( A => n18926, B => n18024, S => n18025, Z => 
                           n17011);
   U17940 : XNOR2_X1 port map( A => n16988, B => n16987, ZN => n16989);
   U17941 : XNOR2_X1 port map( A => n16990, B => n16989, ZN => n16995);
   U17942 : XNOR2_X1 port map( A => n17407, B => n19783, ZN => n17346);
   U17943 : XNOR2_X1 port map( A => n17102, B => n2337, ZN => n16993);
   U17944 : XNOR2_X1 port map( A => n17346, B => n16993, ZN => n16994);
   U17945 : XNOR2_X1 port map( A => n16995, B => n16994, ZN => n18026);
   U17946 : INV_X1 port map( A => n18026, ZN => n18931);
   U17947 : NOR2_X1 port map( A1 => n18931, A2 => n18025, ZN => n17324);
   U17948 : XNOR2_X1 port map( A => n16996, B => n2257, ZN => n16997);
   U17949 : XNOR2_X1 port map( A => n16998, B => n16997, ZN => n17001);
   U17950 : XNOR2_X1 port map( A => n17444, B => n16999, ZN => n17375);
   U17951 : XNOR2_X1 port map( A => n17125, B => n17375, ZN => n17000);
   U17952 : XNOR2_X1 port map( A => n17001, B => n17000, ZN => n18927);
   U17953 : NOR2_X1 port map( A1 => n20207, A2 => n18927, ZN => n17699);
   U17954 : NOR2_X1 port map( A1 => n17324, A2 => n17699, ZN => n17010);
   U17955 : XNOR2_X1 port map( A => n15935, B => n17002, ZN => n17004);
   U17956 : XNOR2_X1 port map( A => n17004, B => n17003, ZN => n17009);
   U17957 : XNOR2_X1 port map( A => n864, B => n17355, ZN => n17007);
   U17958 : XNOR2_X1 port map( A => n17005, B => n2394, ZN => n17006);
   U17959 : XNOR2_X1 port map( A => n17006, B => n17007, ZN => n17008);
   U17961 : INV_X1 port map( A => n18928, ZN => n18932);
   U17962 : XNOR2_X1 port map( A => n17012, B => n17098, ZN => n17013);
   U17963 : XNOR2_X1 port map( A => n17345, B => n17013, ZN => n17018);
   U17964 : XNOR2_X1 port map( A => n17288, B => n17347, ZN => n17016);
   U17965 : XNOR2_X1 port map( A => n17014, B => n1869, ZN => n17015);
   U17966 : XNOR2_X1 port map( A => n17016, B => n17015, ZN => n17017);
   U17967 : XNOR2_X1 port map( A => n17019, B => n17325, ZN => n17023);
   U17968 : XNOR2_X1 port map( A => n17116, B => n2382, ZN => n17021);
   U17969 : XNOR2_X1 port map( A => n17021, B => n17020, ZN => n17022);
   U17970 : XNOR2_X1 port map( A => n17023, B => n17022, ZN => n18939);
   U17971 : NAND2_X1 port map( A1 => n20501, A2 => n18939, ZN => n18021);
   U17972 : INV_X1 port map( A => n19893, ZN => n17025);
   U17973 : XNOR2_X1 port map( A => n17025, B => n17024, ZN => n17027);
   U17974 : XNOR2_X1 port map( A => n17026, B => n17027, ZN => n17031);
   U17975 : XNOR2_X1 port map( A => n17029, B => n17028, ZN => n17030);
   U17976 : XNOR2_X1 port map( A => n17031, B => n17030, ZN => n18936);
   U17979 : XNOR2_X1 port map( A => n17035, B => n19336, ZN => n17037);
   U17980 : XNOR2_X1 port map( A => n17036, B => n17037, ZN => n17038);
   U17982 : XNOR2_X1 port map( A => n17040, B => n17357, ZN => n17044);
   U17983 : XNOR2_X1 port map( A => n16181, B => n19844, ZN => n17042);
   U17984 : XNOR2_X1 port map( A => n17143, B => n18848, ZN => n17041);
   U17985 : XNOR2_X1 port map( A => n17042, B => n17041, ZN => n17043);
   U17986 : INV_X1 port map( A => n17187, ZN => n18941);
   U17987 : AOI21_X1 port map( B1 => n19723, B2 => n18941, A => n18939, ZN => 
                           n17045);
   U17988 : NAND2_X1 port map( A1 => n17705, A2 => n17045, ZN => n17053);
   U17989 : NOR2_X1 port map( A1 => n20501, A2 => n17187, ZN => n17051);
   U17990 : XNOR2_X1 port map( A => n17046, B => n17376, ZN => n17050);
   U17991 : XNOR2_X1 port map( A => n17378, B => n17637, ZN => n17047);
   U17992 : XNOR2_X1 port map( A => n17048, B => n17047, ZN => n17049);
   U17993 : NAND2_X1 port map( A1 => n17051, A2 => n20452, ZN => n17052);
   U17994 : OAI211_X1 port map( C1 => n18021, C2 => n889, A => n17053, B => 
                           n17052, ZN => n18916);
   U17995 : INV_X1 port map( A => n18916, ZN => n18876);
   U17996 : AND2_X1 port map( A1 => n17054, A2 => n18890, ZN => n18874);
   U17997 : AOI22_X1 port map( A1 => n19684, A2 => n935, B1 => n18966, B2 => 
                           n18961, ZN => n17057);
   U17998 : NAND2_X1 port map( A1 => n18966, A2 => n17818, ZN => n17055);
   U18000 : AOI21_X1 port map( B1 => n17059, B2 => n18921, A => n17058, ZN => 
                           n17061);
   U18001 : XNOR2_X1 port map( A => n17061, B => n17060, ZN => Ciphertext(106))
                           ;
   U18002 : NAND2_X1 port map( A1 => n17836, A2 => n17715, ZN => n17196);
   U18003 : OR2_X1 port map( A1 => n17196, A2 => n17062, ZN => n17065);
   U18004 : INV_X1 port map( A => n17063, ZN => n17714);
   U18005 : NAND2_X1 port map( A1 => n17714, A2 => n17840, ZN => n17718);
   U18006 : NOR2_X1 port map( A1 => n17840, A2 => n17715, ZN => n17197);
   U18007 : NAND2_X1 port map( A1 => n17197, A2 => n17838, ZN => n17064);
   U18008 : MUX2_X1 port map( A => n17180, B => n18955, S => n18954, Z => 
                           n17067);
   U18009 : INV_X1 port map( A => n18954, ZN => n17178);
   U18010 : NAND2_X1 port map( A1 => n17178, A2 => n18953, ZN => n17066);
   U18012 : AOI21_X1 port map( B1 => n854, B2 => n17181, A => n17897, ZN => 
                           n17070);
   U18013 : NAND2_X1 port map( A1 => n17070, A2 => n17895, ZN => n17073);
   U18014 : INV_X1 port map( A => n17896, ZN => n17893);
   U18015 : NAND3_X1 port map( A1 => n17893, A2 => n854, A3 => n17181, ZN => 
                           n17072);
   U18016 : NAND3_X1 port map( A1 => n17892, A2 => n17896, A3 => n17897, ZN => 
                           n17071);
   U18018 : MUX2_X1 port map( A => n19163, B => n19155, S => n19162, Z => 
                           n17088);
   U18019 : NAND2_X1 port map( A1 => n17868, A2 => n20514, ZN => n17076);
   U18020 : NAND2_X1 port map( A1 => n19973, A2 => n17078, ZN => n17075);
   U18021 : MUX2_X1 port map( A => n17076, B => n17075, S => n20506, Z => 
                           n17077);
   U18022 : MUX2_X1 port map( A => n17823, B => n17080, S => n17079, Z => 
                           n17083);
   U18023 : MUX2_X1 port map( A => n19667, B => n17824, S => n17825, Z => 
                           n17082);
   U18025 : NOR2_X1 port map( A1 => n19164, A2 => n19162, ZN => n17084);
   U18026 : AOI21_X1 port map( B1 => n19165, B2 => n19948, A => n17084, ZN => 
                           n17087);
   U18027 : OAI21_X1 port map( B1 => n19947, B2 => n20185, A => n17886, ZN => 
                           n17085);
   U18028 : INV_X1 port map( A => n17891, ZN => n17601);
   U18030 : XNOR2_X1 port map( A => n17090, B => n17089, ZN => Ciphertext(140))
                           ;
   U18031 : AND2_X1 port map( A1 => n19463, A2 => n19460, ZN => n17092);
   U18032 : MUX2_X1 port map( A => n20140, B => n19453, S => n20152, Z => 
                           n17093);
   U18033 : NOR2_X1 port map( A1 => n17093, A2 => n19460, ZN => n17094);
   U18035 : NOR2_X1 port map( A1 => n18111, A2 => n20114, ZN => n17096);
   U18036 : MUX2_X1 port map( A => n19885, B => n20488, S => n17458, Z => 
                           n17097);
   U18037 : XNOR2_X1 port map( A => n17099, B => n17098, ZN => n17100);
   U18038 : XNOR2_X1 port map( A => n17101, B => n17100, ZN => n17106);
   U18039 : XNOR2_X1 port map( A => n17102, B => n573, ZN => n17103);
   U18040 : XNOR2_X1 port map( A => n17104, B => n17103, ZN => n17105);
   U18041 : XNOR2_X1 port map( A => n17107, B => n17108, ZN => n17115);
   U18042 : XNOR2_X1 port map( A => n17109, B => n911, ZN => n17113);
   U18043 : XNOR2_X1 port map( A => n17111, B => n18011, ZN => n17112);
   U18044 : XNOR2_X1 port map( A => n17113, B => n17112, ZN => n17114);
   U18045 : XNOR2_X1 port map( A => n17116, B => n2096, ZN => n17117);
   U18046 : XNOR2_X1 port map( A => n17118, B => n17117, ZN => n17122);
   U18047 : XNOR2_X1 port map( A => n17120, B => n17119, ZN => n17121);
   U18048 : XNOR2_X1 port map( A => n17121, B => n17122, ZN => n17547);
   U18049 : INV_X1 port map( A => n17547, ZN => n18229);
   U18050 : XNOR2_X1 port map( A => n17124, B => n17123, ZN => n17126);
   U18051 : XNOR2_X1 port map( A => n17126, B => n17125, ZN => n17132);
   U18052 : XNOR2_X1 port map( A => n19882, B => n17442, ZN => n17130);
   U18053 : XNOR2_X1 port map( A => n17128, B => n18809, ZN => n17129);
   U18054 : XNOR2_X1 port map( A => n17130, B => n17129, ZN => n17131);
   U18055 : XNOR2_X1 port map( A => n17132, B => n17131, ZN => n17390);
   U18056 : INV_X1 port map( A => n17390, ZN => n18232);
   U18057 : XNOR2_X1 port map( A => n19893, B => n17133, ZN => n17136);
   U18058 : XNOR2_X1 port map( A => n17136, B => n17135, ZN => n17140);
   U18059 : XNOR2_X1 port map( A => n880, B => n18084, ZN => n17138);
   U18060 : XNOR2_X1 port map( A => n17142, B => n17141, ZN => n17147);
   U18061 : XNOR2_X1 port map( A => n864, B => n2368, ZN => n17145);
   U18062 : XNOR2_X1 port map( A => n17143, B => n17416, ZN => n17144);
   U18063 : XNOR2_X1 port map( A => n17145, B => n17144, ZN => n17146);
   U18064 : XNOR2_X1 port map( A => n17147, B => n17146, ZN => n18226);
   U18065 : OR2_X1 port map( A1 => n18226, A2 => n17390, ZN => n18121);
   U18066 : MUX2_X1 port map( A => n18121, B => n18229, S => n17545, Z => 
                           n17148);
   U18068 : OAI22_X1 port map( A1 => n19672, A2 => n17553, B1 => n17149, B2 => 
                           n18105, ZN => n17153);
   U18069 : AND2_X1 port map( A1 => n19672, A2 => n17954, ZN => n17151);
   U18070 : NOR2_X1 port map( A1 => n19737, A2 => n17959, ZN => n17150);
   U18073 : MUX2_X1 port map( A => n17489, B => n17154, S => n19675, Z => 
                           n17159);
   U18074 : INV_X1 port map( A => n17491, ZN => n17156);
   U18075 : NOR2_X1 port map( A1 => n17156, A2 => n19675, ZN => n17157);
   U18076 : INV_X1 port map( A => n17623, ZN => n17918);
   U18077 : NAND3_X1 port map( A1 => n18596, A2 => n19669, A3 => n17918, ZN => 
                           n17169);
   U18078 : NOR2_X1 port map( A1 => n18539, A2 => n18535, ZN => n17563);
   U18079 : INV_X1 port map( A => n17563, ZN => n17162);
   U18080 : NAND2_X1 port map( A1 => n17562, A2 => n18535, ZN => n17160);
   U18081 : OAI21_X1 port map( B1 => n18592, B2 => n18589, A => n19665, ZN => 
                           n17168);
   U18082 : NOR2_X1 port map( A1 => n20365, A2 => n18592, ZN => n17167);
   U18083 : MUX2_X2 port map( A => n17166, B => n17165, S => n160, Z => n18597)
                           ;
   U18084 : AOI22_X1 port map( A1 => n17169, A2 => n17168, B1 => n17167, B2 => 
                           n18597, ZN => n17171);
   U18085 : XNOR2_X1 port map( A => n17171, B => n17170, ZN => Ciphertext(48));
   U18086 : OR2_X1 port map( A1 => n17826, A2 => n16262, ZN => n17177);
   U18087 : MUX2_X1 port map( A => n17825, B => n17172, S => n17824, Z => 
                           n17174);
   U18088 : OR2_X1 port map( A1 => n17825, A2 => n17823, ZN => n17173);
   U18089 : MUX2_X1 port map( A => n17174, B => n17173, S => n17822, Z => 
                           n17175);
   U18090 : MUX2_X1 port map( A => n17179, B => n17178, S => n20221, Z => 
                           n19111);
   U18091 : OR2_X1 port map( A1 => n18954, A2 => n18955, ZN => n17832);
   U18092 : NAND2_X1 port map( A1 => n18959, A2 => n18954, ZN => n17829);
   U18093 : NAND2_X1 port map( A1 => n17832, A2 => n17829, ZN => n19106);
   U18095 : INV_X1 port map( A => n17181, ZN => n17894);
   U18096 : AOI21_X1 port map( B1 => n17894, B2 => n17893, A => n17892, ZN => 
                           n17186);
   U18097 : OAI21_X1 port map( B1 => n17184, B2 => n17183, A => n17182, ZN => 
                           n17185);
   U18098 : NAND2_X1 port map( A1 => n19093, A2 => n19911, ZN => n19088);
   U18099 : INV_X1 port map( A => n18938, ZN => n18934);
   U18100 : NOR2_X1 port map( A1 => n18934, A2 => n18937, ZN => n17707);
   U18101 : NAND2_X1 port map( A1 => n17707, A2 => n18935, ZN => n17192);
   U18102 : INV_X1 port map( A => n18019, ZN => n18940);
   U18103 : INV_X1 port map( A => n20452, ZN => n17188);
   U18104 : NAND3_X1 port map( A1 => n18940, A2 => n17188, A3 => n889, ZN => 
                           n17191);
   U18105 : NAND3_X1 port map( A1 => n19723, A2 => n20452, A3 => n18935, ZN => 
                           n17190);
   U18106 : INV_X1 port map( A => n18939, ZN => n18020);
   U18107 : NAND2_X1 port map( A1 => n18020, A2 => n19723, ZN => n17189);
   U18108 : INV_X1 port map( A => n17695, ZN => n17692);
   U18109 : NAND3_X1 port map( A1 => n18961, A2 => n227, A3 => n17692, ZN => 
                           n17195);
   U18110 : INV_X1 port map( A => n17193, ZN => n17819);
   U18111 : OAI211_X1 port map( C1 => n18966, C2 => n20127, A => n17819, B => 
                           n18962, ZN => n17194);
   U18112 : OAI211_X1 port map( C1 => n19684, C2 => n227, A => n17195, B => 
                           n17194, ZN => n17203);
   U18113 : NAND2_X1 port map( A1 => n19115, A2 => n17203, ZN => n19085);
   U18114 : NAND2_X1 port map( A1 => n19088, A2 => n19085, ZN => n17205);
   U18115 : INV_X1 port map( A => n19093, ZN => n19116);
   U18116 : NOR2_X1 port map( A1 => n17196, A2 => n17063, ZN => n17198);
   U18117 : NOR2_X1 port map( A1 => n17198, A2 => n17197, ZN => n17202);
   U18118 : NOR3_X1 port map( A1 => n3755, A2 => n17840, A3 => n17838, ZN => 
                           n17200);
   U18119 : AOI21_X2 port map( B1 => n17202, B2 => n17201, A => n17200, ZN => 
                           n19098);
   U18120 : INV_X1 port map( A => n17203, ZN => n19095);
   U18121 : OAI21_X1 port map( B1 => n19098, B2 => n19095, A => n19115, ZN => 
                           n17204);
   U18122 : AOI22_X1 port map( A1 => n19105, A2 => n17205, B1 => n19116, B2 => 
                           n17204, ZN => n17206);
   U18123 : XNOR2_X1 port map( A => n17206, B => n2216, ZN => Ciphertext(131));
   U18124 : AOI21_X1 port map( B1 => n17211, B2 => n17208, A => n20092, ZN => 
                           n17209);
   U18125 : INV_X1 port map( A => n17209, ZN => n17216);
   U18126 : AND2_X1 port map( A1 => n17210, A2 => n17211, ZN => n17212);
   U18127 : AOI22_X1 port map( A1 => n17214, A2 => n17213, B1 => n16465, B2 => 
                           n17212, ZN => n17215);
   U18129 : MUX2_X1 port map( A => n19383, B => n17218, S => n1897, Z => n17222
                           );
   U18130 : MUX2_X1 port map( A => n19956, B => n17507, S => n17512, Z => 
                           n17230);
   U18131 : NAND2_X1 port map( A1 => n3573, A2 => n17508, ZN => n17228);
   U18133 : NAND3_X1 port map( A1 => n16633, A2 => n14845, A3 => n19956, ZN => 
                           n17227);
   U18134 : OAI21_X1 port map( B1 => n19956, B2 => n17228, A => n17227, ZN => 
                           n17229);
   U18135 : INV_X1 port map( A => n17231, ZN => n17232);
   U18136 : NAND2_X1 port map( A1 => n17232, A2 => n19353, ZN => n17235);
   U18137 : OAI211_X1 port map( C1 => n19352, C2 => n19348, A => n19349, B => 
                           n20273, ZN => n17233);
   U18138 : OAI21_X1 port map( B1 => n17240, B2 => n19666, A => n19372, ZN => 
                           n17238);
   U18139 : INV_X1 port map( A => n17243, ZN => n17241);
   U18141 : NAND2_X1 port map( A1 => n17242, A2 => n20230, ZN => n17247);
   U18142 : AOI22_X1 port map( A1 => n17482, A2 => n17245, B1 => n20354, B2 => 
                           n17243, ZN => n17246);
   U18143 : INV_X1 port map( A => n17249, ZN => n17251);
   U18144 : XNOR2_X1 port map( A => n17250, B => n17251, ZN => n17257);
   U18145 : XNOR2_X1 port map( A => n19807, B => n2310, ZN => n17255);
   U18146 : XNOR2_X1 port map( A => n17253, B => n19845, ZN => n17254);
   U18147 : XNOR2_X1 port map( A => n17255, B => n17254, ZN => n17256);
   U18148 : XNOR2_X1 port map( A => n17257, B => n17256, ZN => n17303);
   U18149 : XNOR2_X1 port map( A => n17259, B => n17258, ZN => n17266);
   U18150 : XNOR2_X1 port map( A => n947, B => n17260, ZN => n17264);
   U18151 : XNOR2_X1 port map( A => n17264, B => n17263, ZN => n17265);
   U18152 : NOR2_X1 port map( A1 => n17753, A2 => n18038, ZN => n17307);
   U18153 : XNOR2_X1 port map( A => n17268, B => n17267, ZN => n17274);
   U18154 : XNOR2_X1 port map( A => n17269, B => n19706, ZN => n17272);
   U18155 : XNOR2_X1 port map( A => n17270, B => n18146, ZN => n17271);
   U18156 : XNOR2_X1 port map( A => n17272, B => n17271, ZN => n17273);
   U18157 : XNOR2_X1 port map( A => n17274, B => n17273, ZN => n17982);
   U18158 : XNOR2_X1 port map( A => n17275, B => n17276, ZN => n17277);
   U18159 : XNOR2_X1 port map( A => n17278, B => n17277, ZN => n17285);
   U18160 : XNOR2_X1 port map( A => n17280, B => n17279, ZN => n17283);
   U18161 : XNOR2_X1 port map( A => n17281, B => n2445, ZN => n17282);
   U18162 : XNOR2_X1 port map( A => n17283, B => n17282, ZN => n17284);
   U18163 : OR2_X1 port map( A1 => n17982, A2 => n18238, ZN => n18241);
   U18164 : XNOR2_X1 port map( A => n17287, B => n17286, ZN => n17292);
   U18165 : XNOR2_X1 port map( A => n19836, B => n2305, ZN => n17290);
   U18166 : INV_X1 port map( A => n17288, ZN => n17289);
   U18167 : XNOR2_X1 port map( A => n17293, B => n17328, ZN => n17297);
   U18168 : XNOR2_X1 port map( A => n17294, B => n17295, ZN => n17296);
   U18169 : XNOR2_X1 port map( A => n17298, B => n17299, ZN => n17302);
   U18170 : XNOR2_X1 port map( A => n17300, B => n17993, ZN => n17301);
   U18171 : NAND2_X1 port map( A1 => n17981, A2 => n18238, ZN => n17983);
   U18176 : INV_X1 port map( A => n19766, ZN => n17992);
   U18177 : INV_X1 port map( A => n18975, ZN => n17308);
   U18178 : NAND2_X1 port map( A1 => n17309, A2 => n18977, ZN => n17313);
   U18179 : NAND2_X1 port map( A1 => n18221, A2 => n20158, ZN => n17311);
   U18181 : MUX2_X1 port map( A => n17311, B => n17310, S => n20499, Z => 
                           n17312);
   U18183 : OAI21_X1 port map( B1 => n19916, B2 => n18946, A => n17315, ZN => 
                           n17316);
   U18184 : NAND2_X1 port map( A1 => n17316, A2 => n20194, ZN => n17319);
   U18185 : NAND2_X1 port map( A1 => n17317, A2 => n19916, ZN => n17318);
   U18187 : NAND2_X1 port map( A1 => n18275, A2 => n18270, ZN => n18274);
   U18188 : OAI21_X1 port map( B1 => n18269, B2 => n18270, A => n18274, ZN => 
                           n17320);
   U18189 : NAND2_X1 port map( A1 => n20097, A2 => n19794, ZN => n18817);
   U18190 : OAI21_X1 port map( B1 => n17992, B2 => n20422, A => n18817, ZN => 
                           n17388);
   U18191 : OAI21_X1 port map( B1 => n2120, B2 => n18928, A => n18926, ZN => 
                           n17323);
   U18192 : NOR2_X1 port map( A1 => n20207, A2 => n18926, ZN => n17748);
   U18193 : INV_X1 port map( A => n18024, ZN => n18929);
   U18194 : INV_X1 port map( A => n18927, ZN => n17700);
   U18195 : NOR2_X1 port map( A1 => n18928, A2 => n17700, ZN => n17321);
   U18196 : AOI22_X1 port map( A1 => n17748, A2 => n18929, B1 => n17321, B2 => 
                           n17749, ZN => n17322);
   U18197 : OAI21_X1 port map( B1 => n17324, B2 => n17323, A => n17322, ZN => 
                           n18844);
   U18198 : INV_X1 port map( A => n18844, ZN => n18818);
   U18199 : XNOR2_X1 port map( A => n17325, B => n17326, ZN => n17334);
   U18200 : XNOR2_X1 port map( A => n17328, B => n20125, ZN => n17332);
   U18201 : INV_X1 port map( A => n18090, ZN => n17329);
   U18202 : XNOR2_X1 port map( A => n17330, B => n17329, ZN => n17331);
   U18203 : XNOR2_X1 port map( A => n17332, B => n17331, ZN => n17333);
   U18204 : XNOR2_X1 port map( A => n17334, B => n17333, ZN => n17394);
   U18205 : INV_X1 port map( A => n17394, ZN => n18258);
   U18206 : XNOR2_X1 port map( A => n17335, B => n20192, ZN => n17336);
   U18207 : XNOR2_X1 port map( A => n17337, B => n17336, ZN => n17344);
   U18208 : XNOR2_X1 port map( A => n17339, B => n17338, ZN => n17342);
   U18209 : XNOR2_X1 port map( A => n19706, B => n19052, ZN => n17341);
   U18210 : XNOR2_X1 port map( A => n17342, B => n17341, ZN => n17343);
   U18212 : NOR2_X1 port map( A1 => n18258, A2 => n19787, ZN => n17976);
   U18213 : INV_X1 port map( A => n17976, ZN => n17978);
   U18214 : XNOR2_X1 port map( A => n17345, B => n17346, ZN => n17353);
   U18215 : XNOR2_X1 port map( A => n19713, B => n17347, ZN => n17351);
   U18216 : XNOR2_X1 port map( A => n19836, B => n20672, ZN => n17350);
   U18217 : XNOR2_X1 port map( A => n17351, B => n17350, ZN => n17352);
   U18218 : XNOR2_X1 port map( A => n17353, B => n17352, ZN => n17374);
   U18219 : XNOR2_X1 port map( A => n15935, B => n17355, ZN => n17356);
   U18220 : XNOR2_X1 port map( A => n17356, B => n17357, ZN => n17364);
   U18221 : XNOR2_X1 port map( A => n17359, B => n17358, ZN => n17362);
   U18222 : XNOR2_X1 port map( A => n17360, B => n17587, ZN => n17361);
   U18223 : XNOR2_X1 port map( A => n17362, B => n17361, ZN => n17363);
   U18224 : NAND2_X1 port map( A1 => n18262, A2 => n18753, ZN => n17396);
   U18225 : XNOR2_X1 port map( A => n17366, B => n17365, ZN => n17368);
   U18226 : XNOR2_X1 port map( A => n17367, B => n17368, ZN => n17369);
   U18227 : XNOR2_X1 port map( A => n17370, B => n17369, ZN => n17372);
   U18228 : NAND2_X1 port map( A1 => n19787, A2 => n18260, ZN => n17373);
   U18229 : NAND3_X1 port map( A1 => n17978, A2 => n17396, A3 => n17373, ZN => 
                           n17385);
   U18230 : INV_X1 port map( A => n17374, ZN => n17977);
   U18231 : XNOR2_X1 port map( A => n17376, B => n17375, ZN => n17382);
   U18232 : XNOR2_X1 port map( A => n19798, B => n456, ZN => n17380);
   U18233 : XNOR2_X1 port map( A => n17382, B => n17381, ZN => n18138);
   U18234 : INV_X1 port map( A => n18138, ZN => n18137);
   U18235 : NAND2_X1 port map( A1 => n18137, A2 => n19787, ZN => n17383);
   U18237 : NAND2_X1 port map( A1 => n18844, A2 => n20097, ZN => n17386);
   U18239 : AOI21_X1 port map( B1 => n20276, B2 => n17386, A => n20130, ZN => 
                           n17387);
   U18240 : AOI21_X1 port map( B1 => n17388, B2 => n18818, A => n17387, ZN => 
                           n17389);
   U18241 : XNOR2_X1 port map( A => n17389, B => n2055, ZN => Ciphertext(90));
   U18242 : INV_X1 port map( A => n18226, ZN => n17549);
   U18243 : NOR2_X1 port map( A1 => n17549, A2 => n19771, ZN => n17392);
   U18244 : AOI21_X1 port map( B1 => n18226, B2 => n17390, A => n18233, ZN => 
                           n17391);
   U18245 : NOR2_X1 port map( A1 => n18226, A2 => n17545, ZN => n18123);
   U18246 : NOR2_X2 port map( A1 => n17393, A2 => n18123, ZN => n18698);
   U18247 : NOR2_X1 port map( A1 => n17394, A2 => n17758, ZN => n17395);
   U18248 : INV_X1 port map( A => n18260, ZN => n18750);
   U18250 : INV_X1 port map( A => n19751, ZN => n17463);
   U18251 : XNOR2_X1 port map( A => n17399, B => n17400, ZN => n17405);
   U18252 : XNOR2_X1 port map( A => n17401, B => n641, ZN => n17402);
   U18253 : XNOR2_X1 port map( A => n17403, B => n17402, ZN => n17404);
   U18254 : XNOR2_X1 port map( A => n17407, B => n17406, ZN => n17408);
   U18255 : XNOR2_X1 port map( A => n17409, B => n17408, ZN => n17415);
   U18256 : XNOR2_X1 port map( A => n17411, B => n17410, ZN => n17413);
   U18257 : INV_X1 port map( A => n2417, ZN => n19038);
   U18258 : XNOR2_X1 port map( A => n17413, B => n17412, ZN => n17414);
   U18260 : XNOR2_X1 port map( A => n20167, B => n2055, ZN => n17417);
   U18261 : XNOR2_X1 port map( A => n17418, B => n17417, ZN => n17422);
   U18262 : XNOR2_X1 port map( A => n17419, B => n17420, ZN => n17421);
   U18263 : MUX2_X1 port map( A => n18130, B => n2475, S => n19744, Z => n17450
                           );
   U18264 : XNOR2_X1 port map( A => n17424, B => n17423, ZN => n17430);
   U18265 : XNOR2_X1 port map( A => n19909, B => n17425, ZN => n17428);
   U18266 : XNOR2_X1 port map( A => n17426, B => n345, ZN => n17427);
   U18267 : XNOR2_X1 port map( A => n17428, B => n17427, ZN => n17429);
   U18268 : XNOR2_X1 port map( A => n17430, B => n17429, ZN => n17946);
   U18269 : XNOR2_X1 port map( A => n17431, B => n17432, ZN => n17437);
   U18270 : XNOR2_X1 port map( A => n17433, B => n18284, ZN => n17434);
   U18271 : XOR2_X1 port map( A => n17435, B => n17434, Z => n17436);
   U18274 : XNOR2_X1 port map( A => n17438, B => n17439, ZN => n17441);
   U18275 : XNOR2_X1 port map( A => n17440, B => n17441, ZN => n17448);
   U18276 : XNOR2_X1 port map( A => n17443, B => n17442, ZN => n17446);
   U18277 : XNOR2_X1 port map( A => n17444, B => n538, ZN => n17445);
   U18278 : XNOR2_X1 port map( A => n17446, B => n17445, ZN => n17447);
   U18279 : XNOR2_X1 port map( A => n17448, B => n17447, ZN => n18129);
   U18280 : AND2_X1 port map( A1 => n17769, A2 => n18273, ZN => n18032);
   U18281 : OAI21_X1 port map( B1 => n17768, B2 => n18032, A => n18269, ZN => 
                           n17453);
   U18282 : INV_X1 port map( A => n17769, ZN => n18267);
   U18283 : OAI21_X1 port map( B1 => n18267, B2 => n18275, A => n18273, ZN => 
                           n17451);
   U18284 : INV_X1 port map( A => n18270, ZN => n17766);
   U18285 : NAND2_X1 port map( A1 => n17451, A2 => n17766, ZN => n17452);
   U18286 : OAI21_X1 port map( B1 => n18698, B2 => n17463, A => n18706, ZN => 
                           n17465);
   U18288 : AOI21_X1 port map( B1 => n396, B2 => n18238, A => n18240, ZN => 
                           n17454);
   U18289 : NAND2_X1 port map( A1 => n17982, A2 => n17981, ZN => n18037);
   U18290 : MUX2_X1 port map( A => n17753, B => n17454, S => n18037, Z => 
                           n17457);
   U18291 : INV_X1 port map( A => n18240, ZN => n17455);
   U18293 : NOR3_X1 port map( A1 => n17455, A2 => n19919, A3 => n17753, ZN => 
                           n17456);
   U18294 : NOR2_X2 port map( A1 => n17457, A2 => n17456, ZN => n18072);
   U18295 : INV_X1 port map( A => n19885, ZN => n18113);
   U18296 : INV_X1 port map( A => n17458, ZN => n18115);
   U18297 : OAI21_X1 port map( B1 => n18111, B2 => n18112, A => n20349, ZN => 
                           n17459);
   U18298 : NAND2_X1 port map( A1 => n17460, A2 => n17459, ZN => n17461);
   U18299 : OAI21_X1 port map( B1 => n20114, B2 => n18113, A => n17461, ZN => 
                           n18701);
   U18300 : OAI21_X1 port map( B1 => n18072, B2 => n18702, A => n18701, ZN => 
                           n17464);
   U18301 : AOI22_X1 port map( A1 => n17465, A2 => n18072, B1 => n17464, B2 => 
                           n17463, ZN => n17467);
   U18302 : XNOR2_X1 port map( A => n17467, B => n17466, ZN => Ciphertext(72));
   U18303 : INV_X1 port map( A => n17564, ZN => n17469);
   U18304 : MUX2_X1 port map( A => n17469, B => n17468, S => n17470, Z => 
                           n17474);
   U18305 : NAND2_X1 port map( A1 => n18539, A2 => n17565, ZN => n17472);
   U18306 : OR2_X1 port map( A1 => n17564, A2 => n17470, ZN => n17561);
   U18307 : MUX2_X1 port map( A => n17472, B => n17561, S => n17471, Z => 
                           n17473);
   U18309 : NOR2_X1 port map( A1 => n18093, A2 => n226, ZN => n17572);
   U18310 : NOR2_X1 port map( A1 => n20109, A2 => n18096, ZN => n17570);
   U18311 : OAI21_X1 port map( B1 => n17572, B2 => n17570, A => n18101, ZN => 
                           n17478);
   U18312 : AOI21_X1 port map( B1 => n18095, B2 => n18097, A => n18096, ZN => 
                           n17476);
   U18314 : NOR2_X1 port map( A1 => n18511, A2 => n18518, ZN => n17519);
   U18315 : NOR2_X1 port map( A1 => n17482, A2 => n17481, ZN => n17486);
   U18316 : NAND2_X1 port map( A1 => n18184, A2 => n18504, ZN => n17524);
   U18317 : OAI211_X1 port map( C1 => n17505, C2 => n17504, A => n17503, B => 
                           n17502, ZN => n17506);
   U18319 : NAND2_X1 port map( A1 => n19758, A2 => n19526, ZN => n17518);
   U18320 : OAI21_X1 port map( B1 => n19956, B2 => n17508, A => n17507, ZN => 
                           n17516);
   U18321 : OAI21_X1 port map( B1 => n19700, B2 => n17510, A => n17509, ZN => 
                           n17515);
   U18322 : NOR2_X1 port map( A1 => n17513, A2 => n17512, ZN => n17514);
   U18323 : NAND2_X1 port map( A1 => n18519, A2 => n18512, ZN => n17517);
   U18324 : INV_X1 port map( A => n2307, ZN => n17522);
   U18325 : NAND3_X1 port map( A1 => n17581, A2 => n2307, A3 => n18505, ZN => 
                           n17527);
   U18326 : INV_X1 port map( A => n17519, ZN => n17521);
   U18327 : INV_X1 port map( A => n17524, ZN => n17520);
   U18328 : NAND3_X1 port map( A1 => n17521, A2 => n17520, A3 => n2307, ZN => 
                           n17526);
   U18329 : INV_X1 port map( A => n18505, ZN => n17523);
   U18330 : NAND3_X1 port map( A1 => n17524, A2 => n17523, A3 => n17522, ZN => 
                           n17525);
   U18331 : AND4_X1 port map( A1 => n17528, A2 => n17527, A3 => n17526, A4 => 
                           n17525, ZN => Ciphertext(31));
   U18332 : INV_X1 port map( A => n19092, ZN => n19109);
   U18335 : INV_X1 port map( A => n19111, ZN => n17530);
   U18336 : NAND2_X1 port map( A1 => n19106, A2 => n19110, ZN => n17529);
   U18338 : NAND2_X1 port map( A1 => n19098, A2 => n17203, ZN => n17531);
   U18339 : AOI21_X1 port map( B1 => n17532, B2 => n17531, A => n19105, ZN => 
                           n17533);
   U18340 : AND4_X1 port map( A1 => n17538, A2 => n17537, A3 => n17536, A4 => 
                           n17610, ZN => n17540);
   U18341 : NAND3_X1 port map( A1 => n17540, A2 => n17539, A3 => n19955, ZN => 
                           n17541);
   U18342 : INV_X1 port map( A => n19339, ZN => n19308);
   U18343 : NAND2_X1 port map( A1 => n19308, A2 => n19340, ZN => n17543);
   U18344 : NOR2_X1 port map( A1 => n19338, A2 => n19339, ZN => n19316);
   U18345 : INV_X1 port map( A => n17545, ZN => n17546);
   U18346 : NOR2_X1 port map( A1 => n17546, A2 => n3066, ZN => n17548);
   U18347 : NOR3_X1 port map( A1 => n17549, A2 => n17390, A3 => n19876, ZN => 
                           n17550);
   U18349 : MUX2_X1 port map( A => n18103, B => n18105, S => n18107, Z => 
                           n17555);
   U18350 : INV_X1 port map( A => n17957, ZN => n18106);
   U18351 : MUX2_X1 port map( A => n17553, B => n17552, S => n18107, Z => 
                           n17554);
   U18354 : OAI21_X1 port map( B1 => n20101, B2 => n19744, A => n17556, ZN => 
                           n18249);
   U18356 : NAND2_X1 port map( A1 => n18249, A2 => n19678, ZN => n17557);
   U18357 : OR2_X1 port map( A1 => n19673, A2 => n19679, ZN => n17578);
   U18358 : NOR2_X1 port map( A1 => n20488, A2 => n20348, ZN => n17965);
   U18359 : INV_X1 port map( A => n17965, ZN => n18213);
   U18360 : INV_X1 port map( A => n20349, ZN => n18633);
   U18361 : NAND3_X1 port map( A1 => n19885, A2 => n17559, A3 => n18633, ZN => 
                           n18211);
   U18362 : OAI21_X1 port map( B1 => n17565, B2 => n20432, A => n17564, ZN => 
                           n17566);
   U18363 : OAI21_X1 port map( B1 => n18538, B2 => n17564, A => n17566, ZN => 
                           n17567);
   U18364 : OAI22_X1 port map( A1 => n17569, A2 => n18096, B1 => n18095, B2 => 
                           n18097, ZN => n17573);
   U18365 : OR3_X1 port map( A1 => n17570, A2 => n18101, A3 => n160, ZN => 
                           n17571);
   U18367 : NAND2_X1 port map( A1 => n18600, A2 => n19757, ZN => n17574);
   U18368 : OAI21_X1 port map( B1 => n18625, B2 => n18600, A => n17574, ZN => 
                           n17575);
   U18369 : NAND2_X1 port map( A1 => n17575, A2 => n19673, ZN => n17577);
   U18370 : OAI211_X1 port map( C1 => n18630, C2 => n17578, A => n17577, B => 
                           n17576, ZN => n17580);
   U18371 : INV_X1 port map( A => n2087, ZN => n17579);
   U18372 : XNOR2_X1 port map( A => n17580, B => n17579, ZN => Ciphertext(58));
   U18373 : OAI21_X1 port map( B1 => n18504, B2 => n18184, A => n18512, ZN => 
                           n17582);
   U18374 : XNOR2_X1 port map( A => n17583, B => n538, ZN => Ciphertext(35));
   U18377 : AOI22_X1 port map( A1 => n17927, A2 => n19668, B1 => n19690, B2 => 
                           n19655, ZN => n17585);
   U18378 : NAND2_X1 port map( A1 => n17586, A2 => n17585, ZN => n17589);
   U18379 : INV_X1 port map( A => n17587, ZN => n17588);
   U18380 : XNOR2_X1 port map( A => n17589, B => n17588, ZN => Ciphertext(36));
   U18381 : INV_X1 port map( A => n17861, ZN => n17864);
   U18382 : AND2_X1 port map( A1 => n19360, A2 => n20212, ZN => n17590);
   U18383 : OAI21_X1 port map( B1 => n17591, B2 => n17590, A => n17864, ZN => 
                           n17594);
   U18385 : OAI21_X1 port map( B1 => n17596, B2 => n19372, A => n19733, ZN => 
                           n17597);
   U18387 : NOR2_X1 port map( A1 => n17600, A2 => n17599, ZN => n17605);
   U18388 : OAI21_X1 port map( B1 => n17601, B2 => n17602, A => n17890, ZN => 
                           n17604);
   U18389 : AND2_X1 port map( A1 => n19947, A2 => n17602, ZN => n17603);
   U18390 : OAI21_X1 port map( B1 => n20364, B2 => n19292, A => n19298, ZN => 
                           n17617);
   U18391 : MUX2_X1 port map( A => n19402, B => n17606, S => n19401, Z => 
                           n17609);
   U18393 : MUX2_X1 port map( A => n17649, B => n17607, S => n19401, Z => 
                           n17608);
   U18395 : NOR2_X1 port map( A1 => n20515, A2 => n19284, ZN => n17616);
   U18396 : INV_X1 port map( A => n17610, ZN => n17614);
   U18397 : INV_X1 port map( A => n17881, ZN => n17613);
   U18398 : OAI211_X1 port map( C1 => n17881, C2 => n196, A => n19930, B => 
                           n3345, ZN => n17612);
   U18399 : OAI21_X1 port map( B1 => n17613, B2 => n19832, A => n17878, ZN => 
                           n17611);
   U18400 : INV_X1 port map( A => n17656, ZN => n19395);
   U18402 : AND2_X1 port map( A1 => n17654, A2 => n20172, ZN => n17618);
   U18403 : INV_X1 port map( A => n19388, ZN => n19400);
   U18404 : AND3_X1 port map( A1 => n19390, A2 => n19396, A3 => n20004, ZN => 
                           n19282);
   U18405 : NOR3_X1 port map( A1 => n19304, A2 => n19292, A3 => n20515, ZN => 
                           n17620);
   U18406 : NOR2_X1 port map( A1 => n17621, A2 => n17620, ZN => n17622);
   U18407 : XNOR2_X1 port map( A => n17622, B => n345, ZN => Ciphertext(172));
   U18408 : INV_X1 port map( A => n18589, ZN => n17624);
   U18409 : NAND3_X1 port map( A1 => n20445, A2 => n19656, A3 => n19669, ZN => 
                           n17625);
   U18410 : OAI211_X1 port map( C1 => n18597, C2 => n17627, A => n17626, B => 
                           n17625, ZN => n17629);
   U18411 : INV_X1 port map( A => n2392, ZN => n17628);
   U18412 : XNOR2_X1 port map( A => n17629, B => n17628, ZN => Ciphertext(52));
   U18413 : NOR2_X1 port map( A1 => n17630, A2 => n18701, ZN => n17633);
   U18414 : NOR2_X1 port map( A1 => n17633, A2 => n17632, ZN => n17634);
   U18415 : XNOR2_X1 port map( A => n17634, B => n2317, ZN => Ciphertext(76));
   U18416 : OAI22_X1 port map( A1 => n19682, A2 => n19691, B1 => n17925, B2 => 
                           n19661, ZN => n18531);
   U18417 : OAI21_X1 port map( B1 => n17923, B2 => n19661, A => n19690, ZN => 
                           n17635);
   U18418 : AOI22_X1 port map( A1 => n18531, A2 => n19668, B1 => n17635, B2 => 
                           n18546, ZN => n17638);
   U18419 : XNOR2_X1 port map( A => n17638, B => n17637, ZN => Ciphertext(41));
   U18420 : NAND2_X1 port map( A1 => n18495, A2 => n18497, ZN => n17914);
   U18421 : NAND2_X1 port map( A1 => n18500, A2 => n17914, ZN => n17642);
   U18422 : AOI21_X1 port map( B1 => n18496, B2 => n18498, A => n645, ZN => 
                           n17641);
   U18423 : OAI21_X1 port map( B1 => n17914, B2 => n893, A => n645, ZN => 
                           n17643);
   U18424 : INV_X1 port map( A => n17643, ZN => n17646);
   U18425 : NAND2_X1 port map( A1 => n18489, A2 => n18495, ZN => n17645);
   U18426 : OAI21_X1 port map( B1 => n17649, B2 => n17650, A => n17648, ZN => 
                           n17653);
   U18427 : MUX2_X1 port map( A => n19404, B => n17650, S => n17853, Z => 
                           n17651);
   U18428 : NOR2_X1 port map( A1 => n19402, A2 => n17651, ZN => n17652);
   U18429 : NOR2_X2 port map( A1 => n17653, A2 => n17652, ZN => n19269);
   U18431 : NAND2_X1 port map( A1 => n19947, A2 => n20185, ZN => n17661);
   U18432 : NAND2_X1 port map( A1 => n16261, A2 => n17663, ZN => n17664);
   U18433 : NOR2_X1 port map( A1 => n17666, A2 => n17876, ZN => n17883);
   U18434 : NAND2_X1 port map( A1 => n17883, A2 => n20162, ZN => n19251);
   U18435 : NAND2_X1 port map( A1 => n17667, A2 => n19251, ZN => n17669);
   U18436 : NOR3_X1 port map( A1 => n17879, A2 => n17668, A3 => n3345, ZN => 
                           n19249);
   U18438 : INV_X1 port map( A => n19276, ZN => n19271);
   U18439 : NOR2_X1 port map( A1 => n19276, A2 => n19246, ZN => n19263);
   U18440 : NOR2_X1 port map( A1 => n20242, A2 => n19938, ZN => n17670);
   U18441 : NOR2_X1 port map( A1 => n17673, A2 => n17864, ZN => n17674);
   U18442 : INV_X1 port map( A => n19278, ZN => n19247);
   U18443 : NAND2_X1 port map( A1 => n19263, A2 => n19247, ZN => n17681);
   U18444 : AND2_X1 port map( A1 => n19246, A2 => n19269, ZN => n17685);
   U18445 : AOI22_X1 port map( A1 => n1112, A2 => n20275, B1 => n20507, B2 => 
                           n20512, ZN => n17679);
   U18446 : OAI21_X1 port map( B1 => n17677, B2 => n17867, A => n17676, ZN => 
                           n17678);
   U18447 : NAND2_X1 port map( A1 => n17685, A2 => n20448, ZN => n17680);
   U18448 : OAI211_X1 port map( C1 => n17682, C2 => n19271, A => n17681, B => 
                           n17680, ZN => n17684);
   U18449 : XNOR2_X1 port map( A => n17684, B => n17683, ZN => Ciphertext(165))
                           ;
   U18450 : NAND2_X1 port map( A1 => n19278, A2 => n19246, ZN => n19261);
   U18451 : AND2_X1 port map( A1 => n18042, A2 => n18946, ZN => n17691);
   U18452 : NAND2_X1 port map( A1 => n18047, A2 => n17687, ZN => n17688);
   U18453 : INV_X1 port map( A => n19034, ZN => n18061);
   U18454 : NOR2_X1 port map( A1 => n18961, A2 => n17818, ZN => n17694);
   U18455 : NOR2_X1 port map( A1 => n18968, A2 => n17692, ZN => n17693);
   U18456 : OR2_X1 port map( A1 => n18968, A2 => n17695, ZN => n17696);
   U18457 : AOI21_X1 port map( B1 => n17817, B2 => n17696, A => n227, ZN => 
                           n17697);
   U18460 : AND2_X1 port map( A1 => n18927, A2 => n18928, ZN => n18028);
   U18461 : NAND2_X1 port map( A1 => n18028, A2 => n18025, ZN => n17703);
   U18462 : NAND2_X1 port map( A1 => n17700, A2 => n18024, ZN => n17701);
   U18463 : MUX2_X1 port map( A => n17701, B => n18029, S => n18025, Z => 
                           n17702);
   U18464 : NAND2_X1 port map( A1 => n18081, A2 => n19046, ZN => n17724);
   U18465 : MUX2_X1 port map( A => n18020, B => n889, S => n19723, Z => n17709)
                           ;
   U18466 : NOR2_X1 port map( A1 => n17707, A2 => n17706, ZN => n17708);
   U18467 : NAND2_X1 port map( A1 => n18954, A2 => n18955, ZN => n17710);
   U18468 : OAI21_X1 port map( B1 => n18959, B2 => n18955, A => n17710, ZN => 
                           n17713);
   U18471 : INV_X1 port map( A => n20264, ZN => n17719);
   U18472 : OAI22_X1 port map( A1 => n16731, A2 => n17719, B1 => n17714, B2 => 
                           n20423, ZN => n17717);
   U18473 : INV_X1 port map( A => n17715, ZN => n17716);
   U18474 : NAND2_X1 port map( A1 => n17717, A2 => n17716, ZN => n17722);
   U18475 : NAND2_X1 port map( A1 => n17063, A2 => n16731, ZN => n17721);
   U18477 : NAND2_X1 port map( A1 => n19046, A2 => n19034, ZN => n17723);
   U18478 : OAI21_X1 port map( B1 => n20475, B2 => n19047, A => n17723, ZN => 
                           n18062);
   U18479 : AOI22_X1 port map( A1 => n17724, A2 => n19047, B1 => n18062, B2 => 
                           n19043, ZN => n17725);
   U18480 : XNOR2_X1 port map( A => n17725, B => n642, ZN => Ciphertext(119));
   U18481 : NAND2_X1 port map( A1 => n18453, A2 => n18468, ZN => n17726);
   U18485 : OAI21_X1 port map( B1 => n19791, B2 => n20231, A => n18468, ZN => 
                           n17727);
   U18486 : AOI22_X1 port map( A1 => n18429, A2 => n18464, B1 => n20110, B2 => 
                           n17727, ZN => n17728);
   U18487 : XNOR2_X1 port map( A => n17728, B => n20593, ZN => Ciphertext(23));
   U18488 : NAND2_X1 port map( A1 => n18485, A2 => n17733, ZN => n17736);
   U18491 : NAND2_X1 port map( A1 => n17731, A2 => n19816, ZN => n17732);
   U18492 : OAI211_X1 port map( C1 => n18500, C2 => n17640, A => n17736, B => 
                           n17732, ZN => n17743);
   U18493 : XNOR2_X1 port map( A => n18498, B => n17733, ZN => n17734);
   U18494 : AOI21_X1 port map( B1 => n17734, B2 => n17640, A => n19816, ZN => 
                           n17742);
   U18495 : NOR2_X1 port map( A1 => n17736, A2 => n17735, ZN => n17738);
   U18496 : NAND2_X1 port map( A1 => n17738, A2 => n17739, ZN => n17741);
   U18499 : NAND2_X1 port map( A1 => n20158, A2 => n18976, ZN => n17746);
   U18500 : OR2_X1 port map( A1 => n18016, A2 => n18977, ZN => n17745);
   U18501 : MUX2_X1 port map( A => n17746, B => n17745, S => n18221, Z => 
                           n17747);
   U18502 : INV_X1 port map( A => n18807, ZN => n18332);
   U18503 : AOI22_X1 port map( A1 => n18931, A2 => n18025, B1 => n18927, B2 => 
                           n18926, ZN => n17750);
   U18504 : OR2_X1 port map( A1 => n18240, A2 => n19919, ZN => n17757);
   U18505 : INV_X1 port map( A => n18237, ZN => n17756);
   U18507 : NAND3_X1 port map( A1 => n20258, A2 => n17753, A3 => n17981, ZN => 
                           n17755);
   U18508 : INV_X1 port map( A => n18238, ZN => n17751);
   U18509 : NAND2_X1 port map( A1 => n3205, A2 => n17751, ZN => n17752);
   U18510 : OAI211_X1 port map( C1 => n17753, C2 => n18240, A => n17982, B => 
                           n17752, ZN => n17754);
   U18512 : NAND2_X1 port map( A1 => n18795, A2 => n19770, ZN => n18335);
   U18513 : INV_X1 port map( A => n17758, ZN => n18256);
   U18514 : NAND2_X1 port map( A1 => n18256, A2 => n18138, ZN => n17759);
   U18515 : NAND2_X1 port map( A1 => n17759, A2 => n18257, ZN => n17761);
   U18516 : NAND2_X1 port map( A1 => n18754, A2 => n18256, ZN => n17760);
   U18517 : MUX2_X1 port map( A => n17761, B => n17760, S => n18260, Z => 
                           n17763);
   U18518 : NAND2_X1 port map( A1 => n17763, A2 => n17762, ZN => n17772);
   U18520 : INV_X1 port map( A => n18806, ZN => n18800);
   U18521 : OAI21_X1 port map( B1 => n18795, B2 => n19811, A => n18800, ZN => 
                           n17773);
   U18522 : NAND2_X1 port map( A1 => n18267, A2 => n18270, ZN => n17765);
   U18523 : MUX2_X1 port map( A => n17765, B => n17764, S => n18275, Z => 
                           n17771);
   U18524 : AND2_X1 port map( A1 => n18033, A2 => n18269, ZN => n17767);
   U18525 : AOI22_X1 port map( A1 => n17769, A2 => n17768, B1 => n17767, B2 => 
                           n17766, ZN => n17770);
   U18526 : NOR2_X1 port map( A1 => n18794, A2 => n17772, ZN => n18333);
   U18527 : INV_X1 port map( A => n17774, ZN => n18128);
   U18528 : AND2_X1 port map( A1 => n17946, A2 => n18130, ZN => n17776);
   U18529 : AOI21_X1 port map( B1 => n18248, B2 => n18129, A => n17776, ZN => 
                           n17780);
   U18530 : NOR2_X1 port map( A1 => n17946, A2 => n17777, ZN => n17778);
   U18531 : NAND2_X1 port map( A1 => n18129, A2 => n17778, ZN => n17779);
   U18532 : INV_X1 port map( A => n18803, ZN => n18331);
   U18533 : INV_X1 port map( A => n18794, ZN => n17781);
   U18534 : NAND3_X1 port map( A1 => n213, A2 => n18331, A3 => n17781, ZN => 
                           n17782);
   U18535 : INV_X1 port map( A => n2329, ZN => n17783);
   U18536 : NAND2_X1 port map( A1 => n19302, A2 => n19292, ZN => n19290);
   U18537 : OR2_X1 port map( A1 => n19284, A2 => n19292, ZN => n18164);
   U18538 : MUX2_X1 port map( A => n19770, B => n19711, S => n18807, Z => 
                           n17786);
   U18539 : NOR2_X1 port map( A1 => n19811, A2 => n18807, ZN => n17784);
   U18540 : MUX2_X1 port map( A => n17784, B => n18803, S => n19711, Z => 
                           n17785);
   U18541 : AOI21_X1 port map( B1 => n18795, B2 => n17786, A => n17785, ZN => 
                           n17788);
   U18542 : XNOR2_X1 port map( A => n17788, B => n17787, ZN => Ciphertext(84));
   U18545 : OAI22_X1 port map( A1 => n17789, A2 => n17794, B1 => n2896, B2 => 
                           n17793, ZN => n17795);
   U18546 : NOR3_X1 port map( A1 => n17797, A2 => n17796, A3 => n17795, ZN => 
                           Ciphertext(139));
   U18547 : NAND2_X1 port map( A1 => n18697, A2 => n19753, ZN => n17799);
   U18548 : OAI21_X1 port map( B1 => n18698, B2 => n18701, A => n17799, ZN => 
                           n18695);
   U18549 : INV_X1 port map( A => n18072, ZN => n17803);
   U18550 : INV_X1 port map( A => n18701, ZN => n17800);
   U18551 : OAI21_X1 port map( B1 => n18698, B2 => n19751, A => n17800, ZN => 
                           n17802);
   U18552 : AOI22_X1 port map( A1 => n18695, A2 => n17803, B1 => n17802, B2 => 
                           n1055, ZN => n17805);
   U18553 : XNOR2_X1 port map( A => n17805, B => n17804, ZN => Ciphertext(77));
   U18554 : INV_X1 port map( A => n19143, ZN => n19133);
   U18556 : AND2_X1 port map( A1 => n20508, A2 => n19144, ZN => n19127);
   U18557 : NAND2_X1 port map( A1 => n19127, A2 => n19134, ZN => n17809);
   U18558 : INV_X1 port map( A => n19146, ZN => n19125);
   U18559 : NAND2_X1 port map( A1 => n17807, A2 => n19125, ZN => n17808);
   U18560 : OAI211_X1 port map( C1 => n17810, C2 => n19144, A => n17809, B => 
                           n17808, ZN => n17811);
   U18561 : XNOR2_X1 port map( A => n17811, B => n2079, ZN => Ciphertext(134));
   U18562 : AND2_X1 port map( A1 => n18046, A2 => n17812, ZN => n18045);
   U18563 : INV_X1 port map( A => n18045, ZN => n17816);
   U18564 : NAND3_X1 port map( A1 => n20194, A2 => n17687, A3 => n17812, ZN => 
                           n17815);
   U18565 : NAND4_X1 port map( A1 => n17816, A2 => n17815, A3 => n17814, A4 => 
                           n17813, ZN => n19059);
   U18566 : NAND2_X1 port map( A1 => n17819, A2 => n18961, ZN => n18965);
   U18567 : MUX2_X1 port map( A => n19059, B => n19685, S => n19060, Z => 
                           n17850);
   U18568 : OR2_X1 port map( A1 => n17836, A2 => n16731, ZN => n17839);
   U18569 : OAI211_X1 port map( C1 => n17715, C2 => n17838, A => n17063, B => 
                           n17839, ZN => n17843);
   U18570 : INV_X1 port map( A => n17839, ZN => n17841);
   U18571 : NAND2_X1 port map( A1 => n17841, A2 => n17840, ZN => n17842);
   U18572 : AND2_X1 port map( A1 => n19060, A2 => n19067, ZN => n19064);
   U18573 : NOR2_X1 port map( A1 => n20452, A2 => n18935, ZN => n17847);
   U18574 : OR2_X1 port map( A1 => n18939, A2 => n18936, ZN => n17845);
   U18575 : MUX2_X1 port map( A => n17845, B => n20501, S => n17187, Z => 
                           n17846);
   U18576 : OAI21_X2 port map( B1 => n18933, B2 => n17847, A => n17846, ZN => 
                           n19073);
   U18577 : NOR2_X1 port map( A1 => n19060, A2 => n19073, ZN => n17848);
   U18578 : AOI22_X1 port map( A1 => n19064, A2 => n19685, B1 => n17848, B2 => 
                           n20131, ZN => n17849);
   U18579 : OAI21_X1 port map( B1 => n17850, B2 => n20131, A => n17849, ZN => 
                           n17852);
   U18580 : XNOR2_X1 port map( A => n17852, B => n17851, ZN => Ciphertext(122))
                           ;
   U18581 : MUX2_X1 port map( A => n19401, B => n19402, S => n19404, Z => 
                           n17856);
   U18582 : INV_X1 port map( A => n19402, ZN => n17854);
   U18583 : NOR2_X1 port map( A1 => n17854, A2 => n17853, ZN => n17855);
   U18584 : INV_X1 port map( A => n19403, ZN => n17857);
   U18585 : NOR3_X1 port map( A1 => n19401, A2 => n17857, A3 => n19402, ZN => 
                           n17858);
   U18586 : OAI21_X1 port map( B1 => n20150, B2 => n17861, A => n17860, ZN => 
                           n19366);
   U18587 : AOI21_X1 port map( B1 => n17863, B2 => n20212, A => n20242, ZN => 
                           n17865);
   U18588 : OR2_X1 port map( A1 => n17865, A2 => n17864, ZN => n17866);
   U18589 : NAND2_X1 port map( A1 => n19242, A2 => n20124, ZN => n17904);
   U18590 : NAND2_X1 port map( A1 => n20275, A2 => n17867, ZN => n17869);
   U18591 : MUX2_X1 port map( A => n20507, B => n17869, S => n17868, Z => 
                           n17875);
   U18592 : OAI211_X1 port map( C1 => n20512, C2 => n17873, A => n19973, B => 
                           n1112, ZN => n17874);
   U18593 : NAND2_X1 port map( A1 => n17875, A2 => n17874, ZN => n19235);
   U18595 : AND2_X1 port map( A1 => n19754, A2 => n19227, ZN => n17903);
   U18596 : AND2_X1 port map( A1 => n17890, A2 => n17886, ZN => n17888);
   U18597 : INV_X1 port map( A => n19233, ZN => n19236);
   U18598 : AND2_X1 port map( A1 => n17892, A2 => n17893, ZN => n17902);
   U18599 : AOI21_X1 port map( B1 => n17894, B2 => n17898, A => n17893, ZN => 
                           n17901);
   U18600 : NOR2_X1 port map( A1 => n17895, A2 => n17897, ZN => n17899);
   U18601 : INV_X1 port map( A => n19237, ZN => n18190);
   U18602 : XNOR2_X1 port map( A => n17905, B => n1857, ZN => Ciphertext(157));
   U18603 : BUF_X1 port map( A => n18287, Z => n17936);
   U18604 : MUX2_X1 port map( A => n18357, B => n17907, S => n18362, Z => 
                           n17908);
   U18605 : XNOR2_X1 port map( A => n17910, B => n17909, ZN => Ciphertext(1));
   U18606 : NAND3_X1 port map( A1 => n19729, A2 => n18497, A3 => n17640, ZN => 
                           n17913);
   U18607 : INV_X1 port map( A => n19242, ZN => n17916);
   U18608 : NAND2_X1 port map( A1 => n19219, A2 => n20193, ZN => n17915);
   U18609 : XNOR2_X1 port map( A => n17917, B => Key(60), ZN => Ciphertext(161)
                           );
   U18610 : NAND2_X1 port map( A1 => n18590, A2 => n18589, ZN => n18584);
   U18611 : NOR2_X1 port map( A1 => n18589, A2 => n17918, ZN => n18593);
   U18612 : OAI21_X1 port map( B1 => n18573, B2 => n18584, A => n17919, ZN => 
                           n17921);
   U18613 : NOR2_X1 port map( A1 => n18597, A2 => n20365, ZN => n17920);
   U18614 : NOR2_X1 port map( A1 => n17921, A2 => n17920, ZN => n17922);
   U18615 : XNOR2_X1 port map( A => n17922, B => n484, ZN => Ciphertext(49));
   U18616 : NAND3_X1 port map( A1 => n17923, A2 => n19690, A3 => n19691, ZN => 
                           n17930);
   U18617 : NAND3_X1 port map( A1 => n17925, A2 => n19661, A3 => n19691, ZN => 
                           n17929);
   U18618 : NAND4_X1 port map( A1 => n17931, A2 => n17930, A3 => n17929, A4 => 
                           n17928, ZN => n17934);
   U18619 : INV_X1 port map( A => n17932, ZN => n17933);
   U18620 : XNOR2_X1 port map( A => n17934, B => n17933, ZN => Ciphertext(40));
   U18621 : OAI21_X1 port map( B1 => n18362, B2 => n18348, A => n18290, ZN => 
                           n17939);
   U18622 : INV_X1 port map( A => n17935, ZN => n18350);
   U18623 : NAND2_X1 port map( A1 => n17936, A2 => n18350, ZN => n18364);
   U18624 : OAI211_X1 port map( C1 => n18362, C2 => n18359, A => n18364, B => 
                           n18292, ZN => n17938);
   U18625 : AOI22_X1 port map( A1 => n17938, A2 => n17939, B1 => n17937, B2 => 
                           n18357, ZN => n17941);
   U18626 : XNOR2_X1 port map( A => n17941, B => n17940, ZN => Ciphertext(2));
   U18627 : NOR2_X1 port map( A1 => n19093, A2 => n19109, ZN => n17944);
   U18628 : OAI21_X1 port map( B1 => n19095, B2 => n19112, A => n19093, ZN => 
                           n17943);
   U18629 : NAND2_X1 port map( A1 => n19095, A2 => n19098, ZN => n19089);
   U18630 : NAND2_X1 port map( A1 => n18248, A2 => n19678, ZN => n17953);
   U18631 : NOR2_X1 port map( A1 => n19472, A2 => n18130, ZN => n17945);
   U18632 : NOR2_X1 port map( A1 => n18131, A2 => n17946, ZN => n18251);
   U18635 : OR2_X1 port map( A1 => n18251, A2 => n17950, ZN => n17951);
   U18637 : OAI21_X1 port map( B1 => n17956, B2 => n19672, A => n17954, ZN => 
                           n17958);
   U18638 : NAND2_X1 port map( A1 => n17958, A2 => n17957, ZN => n17963);
   U18639 : NAND3_X1 port map( A1 => n17956, A2 => n17959, A3 => n18106, ZN => 
                           n17962);
   U18640 : NAND3_X1 port map( A1 => n17956, A2 => n18103, A3 => n18107, ZN => 
                           n17961);
   U18642 : NAND2_X1 port map( A1 => n17965, A2 => n18115, ZN => n17971);
   U18643 : INV_X1 port map( A => n17966, ZN => n17970);
   U18644 : NOR2_X1 port map( A1 => n18112, A2 => n20349, ZN => n17967);
   U18645 : OR2_X1 port map( A1 => n17968, A2 => n17967, ZN => n17969);
   U18646 : NAND2_X1 port map( A1 => n18672, A2 => n18671, ZN => n17972);
   U18647 : AOI21_X1 port map( B1 => n17390, B2 => n19876, A => n17973, ZN => 
                           n17975);
   U18648 : NOR2_X1 port map( A1 => n18229, A2 => n18233, ZN => n18122);
   U18649 : NOR2_X1 port map( A1 => n18122, A2 => n18120, ZN => n17974);
   U18650 : MUX2_X1 port map( A => n18137, B => n17976, S => n18753, Z => 
                           n17980);
   U18651 : NAND2_X1 port map( A1 => n18262, A2 => n18256, ZN => n18752);
   U18652 : AOI21_X1 port map( B1 => n18258, B2 => n18260, A => n17977, ZN => 
                           n17979);
   U18653 : NOR2_X1 port map( A1 => n18682, A2 => n19735, ZN => n17986);
   U18654 : NAND2_X1 port map( A1 => n17986, A2 => n17985, ZN => n17987);
   U18656 : OAI21_X1 port map( B1 => n17992, B2 => n20276, A => n17991, ZN => 
                           n18845);
   U18657 : NAND2_X1 port map( A1 => n18818, A2 => n18172, ZN => n18174);
   U18658 : AOI22_X1 port map( A1 => n18845, A2 => n18817, B1 => n18811, B2 => 
                           n18174, ZN => n17994);
   U18659 : XNOR2_X1 port map( A => n17994, B => n17993, ZN => Ciphertext(91));
   U18660 : NAND2_X1 port map( A1 => n19775, A2 => n18568, ZN => n17996);
   U18662 : AOI21_X1 port map( B1 => n17997, B2 => n17996, A => n20169, ZN => 
                           n17998);
   U18663 : XNOR2_X1 port map( A => n18000, B => n17999, ZN => Ciphertext(46));
   U18664 : NAND2_X1 port map( A1 => n18568, A2 => n18556, ZN => n18560);
   U18665 : INV_X1 port map( A => n18559, ZN => n18570);
   U18666 : NOR2_X1 port map( A1 => n18199, A2 => n18559, ZN => n18002);
   U18667 : INV_X1 port map( A => n18567, ZN => n18001);
   U18668 : OAI21_X1 port map( B1 => n18002, B2 => n18565, A => n18001, ZN => 
                           n18005);
   U18669 : OAI211_X1 port map( C1 => n18560, C2 => n18570, A => n18005, B => 
                           n18004, ZN => n18008);
   U18670 : INV_X1 port map( A => n18006, ZN => n18007);
   U18671 : XNOR2_X1 port map( A => n18008, B => n18007, ZN => Ciphertext(42));
   U18672 : MUX2_X1 port map( A => n20492, B => n18522, S => n18512, Z => 
                           n18010);
   U18673 : INV_X1 port map( A => n18011, ZN => n18012);
   U18674 : OAI21_X1 port map( B1 => n19459, B2 => n19453, A => n19460, ZN => 
                           n18013);
   U18675 : AOI22_X1 port map( A1 => n18014, A2 => n19459, B1 => n18013, B2 => 
                           n20152, ZN => n18015);
   U18676 : XNOR2_X1 port map( A => n18015, B => n2383, ZN => Ciphertext(186));
   U18677 : MUX2_X1 port map( A => n18016, B => n20499, S => n18221, Z => 
                           n18018);
   U18678 : MUX2_X1 port map( A => n18975, B => n18976, S => n18978, Z => 
                           n18017);
   U18679 : MUX2_X2 port map( A => n18018, B => n18017, S => n18977, Z => 
                           n18869);
   U18680 : AOI22_X1 port map( A1 => n18020, A2 => n18937, B1 => n20501, B2 => 
                           n19723, ZN => n18023);
   U18681 : NAND3_X1 port map( A1 => n18934, A2 => n18937, A3 => n18935, ZN => 
                           n18022);
   U18685 : MUX2_X1 port map( A => n18270, B => n18032, S => n18268, Z => 
                           n18036);
   U18686 : OAI211_X1 port map( C1 => n18269, C2 => n18033, A => n18275, B => 
                           n18267, ZN => n18034);
   U18687 : INV_X1 port map( A => n18034, ZN => n18035);
   U18688 : MUX2_X1 port map( A => n19988, B => n20418, S => n18857, Z => 
                           n18054);
   U18689 : NOR2_X1 port map( A1 => n18240, A2 => n20132, ZN => n18040);
   U18690 : NAND2_X1 port map( A1 => n20258, A2 => n18038, ZN => n18039);
   U18692 : INV_X1 port map( A => n18866, ZN => n18850);
   U18693 : NOR2_X1 port map( A1 => n20418, A2 => n18850, ZN => n18052);
   U18694 : NOR2_X1 port map( A1 => n18043, A2 => n18042, ZN => n18044);
   U18696 : NAND2_X1 port map( A1 => n18948, A2 => n2586, ZN => n18048);
   U18697 : AOI21_X1 port map( B1 => n18949, B2 => n18048, A => n18047, ZN => 
                           n18049);
   U18701 : INV_X1 port map( A => n19168, ZN => n18323);
   U18702 : NAND2_X1 port map( A1 => n18057, A2 => n18157, ZN => n18058);
   U18703 : OAI21_X1 port map( B1 => n20460, B2 => n18323, A => n18058, ZN => 
                           n18089);
   U18704 : AOI22_X1 port map( A1 => n18089, A2 => n19170, B1 => n18323, B2 => 
                           n18059, ZN => n18060);
   U18705 : XNOR2_X1 port map( A => n18060, B => n2257, ZN => Ciphertext(149));
   U18707 : NOR2_X1 port map( A1 => n20142, A2 => n19032, ZN => n18064);
   U18708 : NAND2_X1 port map( A1 => n19047, A2 => n19032, ZN => n19031);
   U18709 : NAND2_X1 port map( A1 => n18062, A2 => n19031, ZN => n18063);
   U18710 : INV_X1 port map( A => n18065, ZN => n18066);
   U18711 : MUX2_X1 port map( A => n19460, B => n19463, S => n20152, Z => 
                           n18069);
   U18712 : MUX2_X1 port map( A => n19459, B => n19462, S => n20140, Z => 
                           n18068);
   U18713 : XNOR2_X1 port map( A => n18071, B => n18070, ZN => Ciphertext(188))
                           ;
   U18714 : MUX2_X1 port map( A => n18072, B => n19751, S => n18697, Z => 
                           n18074);
   U18715 : MUX2_X1 port map( A => n18698, B => n18701, S => n18703, Z => 
                           n18073);
   U18716 : MUX2_X1 port map( A => n18074, B => n18073, S => n19753, Z => 
                           n18076);
   U18717 : XNOR2_X1 port map( A => n18076, B => n18075, ZN => Ciphertext(74));
   U18719 : NOR2_X1 port map( A1 => n18392, A2 => n18384, ZN => n18077);
   U18721 : NAND2_X1 port map( A1 => n19992, A2 => n19046, ZN => n18080);
   U18722 : NAND2_X1 port map( A1 => n18081, A2 => n18080, ZN => n18082);
   U18723 : MUX2_X1 port map( A => n18083, B => n18082, S => n19032, Z => 
                           n18086);
   U18724 : INV_X1 port map( A => n18084, ZN => n18085);
   U18725 : XNOR2_X1 port map( A => n18086, B => n18085, ZN => Ciphertext(116))
                           ;
   U18726 : INV_X1 port map( A => n18327, ZN => n19174);
   U18727 : INV_X1 port map( A => n19169, ZN => n18087);
   U18728 : AOI22_X1 port map( A1 => n18089, A2 => n18088, B1 => n18161, B2 => 
                           n18087, ZN => n18091);
   U18729 : XNOR2_X1 port map( A => n18091, B => n18090, ZN => Ciphertext(145))
                           ;
   U18730 : AOI22_X1 port map( A1 => n18095, A2 => n18094, B1 => n19774, B2 => 
                           n160, ZN => n18102);
   U18731 : INV_X1 port map( A => n18096, ZN => n18098);
   U18732 : OAI21_X1 port map( B1 => n18099, B2 => n18098, A => n18097, ZN => 
                           n18100);
   U18734 : INV_X1 port map( A => n18651, ZN => n18119);
   U18735 : NAND2_X1 port map( A1 => n19737, A2 => n18107, ZN => n18104);
   U18736 : OAI211_X1 port map( C1 => n19658, C2 => n18107, A => n18106, B => 
                           n18105, ZN => n18109);
   U18738 : MUX2_X1 port map( A => n18113, B => n18112, S => n18111, Z => 
                           n18636);
   U18739 : AND2_X1 port map( A1 => n18115, A2 => n19885, ZN => n18117);
   U18740 : MUX2_X2 port map( A => n18636, B => n18634, S => n20349, Z => 
                           n18656);
   U18742 : AOI21_X1 port map( B1 => n18119, B2 => n18648, A => n19624, ZN => 
                           n18145);
   U18743 : AOI22_X1 port map( A1 => n18123, A2 => n3066, B1 => n18122, B2 => 
                           n18226, ZN => n18124);
   U18744 : NAND2_X1 port map( A1 => n18125, A2 => n18124, ZN => n18644);
   U18745 : AND2_X1 port map( A1 => n18644, A2 => n18651, ZN => n18144);
   U18746 : INV_X1 port map( A => n18144, ZN => n18641);
   U18747 : AOI21_X1 port map( B1 => n18128, B2 => n18127, A => n18126, ZN => 
                           n18136);
   U18748 : NOR2_X1 port map( A1 => n18129, A2 => n19472, ZN => n18134);
   U18749 : NOR2_X1 port map( A1 => n18131, A2 => n18130, ZN => n18133);
   U18750 : MUX2_X1 port map( A => n18134, B => n18133, S => n20101, Z => 
                           n18135);
   U18752 : NOR2_X1 port map( A1 => n18656, A2 => n18650, ZN => n18143);
   U18753 : AOI21_X1 port map( B1 => n18137, B2 => n18754, A => n18262, ZN => 
                           n18142);
   U18754 : NAND2_X1 port map( A1 => n18257, A2 => n18138, ZN => n18139);
   U18755 : AOI21_X1 port map( B1 => n18139, B2 => n18260, A => n18258, ZN => 
                           n18141);
   U18756 : INV_X1 port map( A => n19757, ZN => n18626);
   U18758 : NAND3_X1 port map( A1 => n18625, A2 => n19673, A3 => n18626, ZN => 
                           n18147);
   U18759 : INV_X1 port map( A => n2221, ZN => n18148);
   U18760 : NOR2_X1 port map( A1 => n19685, A2 => n19073, ZN => n18150);
   U18761 : INV_X1 port map( A => n19059, ZN => n19075);
   U18762 : AND2_X1 port map( A1 => n19075, A2 => n19060, ZN => n18149);
   U18763 : INV_X1 port map( A => n19074, ZN => n19058);
   U18764 : MUX2_X1 port map( A => n18150, B => n18149, S => n19058, Z => 
                           n18154);
   U18765 : INV_X1 port map( A => n18151, ZN => n19069);
   U18767 : NAND2_X1 port map( A1 => n19079, A2 => n19073, ZN => n18152);
   U18768 : OAI21_X1 port map( B1 => n19055, B2 => n19067, A => n18152, ZN => 
                           n18153);
   U18769 : NOR2_X1 port map( A1 => n18154, A2 => n18153, ZN => n18155);
   U18770 : XNOR2_X1 port map( A => n18155, B => n1869, ZN => Ciphertext(123));
   U18771 : OAI21_X1 port map( B1 => n18156, B2 => n20460, A => n18320, ZN => 
                           n18160);
   U18772 : INV_X1 port map( A => n18157, ZN => n18318);
   U18773 : OAI21_X1 port map( B1 => n18318, B2 => n18319, A => n18158, ZN => 
                           n18159);
   U18774 : AOI22_X1 port map( A1 => n18161, A2 => n18160, B1 => n18159, B2 => 
                           n18323, ZN => n18162);
   U18775 : XNOR2_X1 port map( A => n18162, B => n1840, ZN => Ciphertext(148));
   U18776 : NAND2_X1 port map( A1 => n20434, A2 => n19284, ZN => n18163);
   U18777 : OAI21_X1 port map( B1 => n19298, B2 => n19284, A => n18163, ZN => 
                           n18165);
   U18779 : NAND2_X1 port map( A1 => n18688, A2 => n19735, ZN => n18679);
   U18780 : OAI21_X1 port map( B1 => n18672, B2 => n18666, A => n18679, ZN => 
                           n18169);
   U18782 : OAI21_X1 port map( B1 => n18682, B2 => n19510, A => n18671, ZN => 
                           n18168);
   U18783 : AOI22_X1 port map( A1 => n18169, A2 => n18682, B1 => n18666, B2 => 
                           n18168, ZN => n18171);
   U18784 : XNOR2_X1 port map( A => n18171, B => n18170, ZN => Ciphertext(66));
   U18785 : OR2_X1 port map( A1 => n18831, A2 => n18172, ZN => n18827);
   U18786 : OAI22_X1 port map( A1 => n18827, A2 => n18834, B1 => n18813, B2 => 
                           n20097, ZN => n18176);
   U18787 : NAND2_X1 port map( A1 => n20422, A2 => n19766, ZN => n18841);
   U18788 : OAI21_X1 port map( B1 => n20130, B2 => n20097, A => n18841, ZN => 
                           n18175);
   U18789 : OAI22_X1 port map( A1 => n18176, A2 => n18175, B1 => n18813, B2 => 
                           n18174, ZN => n18178);
   U18790 : XNOR2_X1 port map( A => n18178, B => n18177, ZN => Ciphertext(92));
   U18791 : NAND2_X1 port map( A1 => n18630, A2 => n18600, ZN => n18181);
   U18792 : INV_X1 port map( A => n18625, ZN => n18619);
   U18795 : AOI22_X1 port map( A1 => n18181, A2 => n18180, B1 => n18179, B2 => 
                           n18630, ZN => n18182);
   U18796 : XNOR2_X1 port map( A => n18182, B => n2100, ZN => Ciphertext(54));
   U18797 : MUX2_X1 port map( A => n18522, B => n18511, S => n19773, Z => 
                           n18186);
   U18798 : NAND2_X1 port map( A1 => n18504, A2 => n18512, ZN => n18183);
   U18799 : OAI21_X1 port map( B1 => n18504, B2 => n18184, A => n18183, ZN => 
                           n18185);
   U18800 : MUX2_X1 port map( A => n18186, B => n18185, S => n19758, Z => 
                           n18188);
   U18801 : INV_X1 port map( A => n2375, ZN => n18187);
   U18802 : XNOR2_X1 port map( A => n18188, B => n18187, ZN => Ciphertext(32));
   U18803 : INV_X1 port map( A => n19227, ZN => n19239);
   U18804 : OAI21_X1 port map( B1 => n19754, B2 => n19239, A => n19229, ZN => 
                           n18193);
   U18805 : NAND2_X1 port map( A1 => n19242, A2 => n18190, ZN => n18192);
   U18806 : NOR2_X1 port map( A1 => n19237, A2 => n19238, ZN => n19225);
   U18807 : NOR2_X1 port map( A1 => n19225, A2 => n19227, ZN => n18191);
   U18808 : AOI22_X1 port map( A1 => n18193, A2 => n19242, B1 => n18192, B2 => 
                           n18191, ZN => n18194);
   U18809 : XNOR2_X1 port map( A => n18194, B => n2296, ZN => Ciphertext(156));
   U18810 : INV_X1 port map( A => n18644, ZN => n18654);
   U18811 : INV_X1 port map( A => n18648, ZN => n18642);
   U18812 : OAI21_X1 port map( B1 => n18654, B2 => n18642, A => n18651, ZN => 
                           n18197);
   U18813 : NAND2_X1 port map( A1 => n18648, A2 => n18651, ZN => n18195);
   U18814 : OAI21_X1 port map( B1 => n18656, B2 => n19935, A => n18195, ZN => 
                           n18647);
   U18815 : INV_X1 port map( A => n19745, ZN => n18196);
   U18816 : AOI22_X1 port map( A1 => n18197, A2 => n18656, B1 => n18647, B2 => 
                           n18196, ZN => n18198);
   U18817 : XNOR2_X1 port map( A => n18198, B => n2306, ZN => Ciphertext(65));
   U18818 : NAND2_X1 port map( A1 => n18555, A2 => n18565, ZN => n18200);
   U18819 : NAND2_X1 port map( A1 => n18561, A2 => n18200, ZN => n18571);
   U18820 : INV_X1 port map( A => n18555, ZN => n18566);
   U18821 : AND2_X1 port map( A1 => n19775, A2 => n18566, ZN => n18202);
   U18822 : AOI22_X1 port map( A1 => n18571, A2 => n18560, B1 => n18202, B2 => 
                           n18201, ZN => n18204);
   U18823 : XNOR2_X1 port map( A => n18204, B => n18203, ZN => Ciphertext(43));
   U18824 : OAI21_X1 port map( B1 => n20142, B2 => n18061, A => n19992, ZN => 
                           n18205);
   U18825 : OAI21_X1 port map( B1 => n19993, B2 => n19046, A => n18205, ZN => 
                           n18207);
   U18826 : NAND3_X1 port map( A1 => n938, A2 => n20142, A3 => n19032, ZN => 
                           n18206);
   U18828 : INV_X1 port map( A => n18208, ZN => n18209);
   U18831 : INV_X1 port map( A => n18211, ZN => n18212);
   U18832 : AOI21_X1 port map( B1 => n18214, B2 => n18213, A => n18212, ZN => 
                           n18215);
   U18833 : AND2_X1 port map( A1 => n18622, A2 => n19509, ZN => n18218);
   U18834 : NAND2_X1 port map( A1 => n18218, A2 => n18630, ZN => n18217);
   U18835 : OAI21_X1 port map( B1 => n18219, B2 => n18218, A => n18217, ZN => 
                           n18220);
   U18836 : XNOR2_X1 port map( A => n18220, B => n2420, ZN => Ciphertext(56));
   U18837 : NOR2_X1 port map( A1 => n20158, A2 => n18978, ZN => n18225);
   U18838 : OAI21_X1 port map( B1 => n18225, B2 => n18976, A => n224, ZN => 
                           n18722);
   U18839 : NAND2_X1 port map( A1 => n18721, A2 => n18722, ZN => n18709);
   U18840 : INV_X1 port map( A => n18709, ZN => n18763);
   U18841 : NOR2_X1 port map( A1 => n18232, A2 => n18226, ZN => n18227);
   U18842 : NAND2_X1 port map( A1 => n19876, A2 => n18227, ZN => n18236);
   U18843 : INV_X1 port map( A => n18233, ZN => n18228);
   U18844 : NAND3_X1 port map( A1 => n18228, A2 => n17390, A3 => n3066, ZN => 
                           n18231);
   U18845 : NAND2_X1 port map( A1 => n18229, A2 => n18233, ZN => n18230);
   U18846 : AND2_X1 port map( A1 => n18231, A2 => n18230, ZN => n18235);
   U18847 : NAND3_X1 port map( A1 => n17549, A2 => n18233, A3 => n18232, ZN => 
                           n18234);
   U18848 : INV_X1 port map( A => n18762, ZN => n18772);
   U18851 : NAND3_X1 port map( A1 => n20258, A2 => n396, A3 => n20132, ZN => 
                           n18245);
   U18854 : INV_X1 port map( A => n18248, ZN => n18250);
   U18855 : OAI21_X1 port map( B1 => n19678, B2 => n19472, A => n18251, ZN => 
                           n18254);
   U18856 : OAI21_X1 port map( B1 => n18762, B2 => n19803, A => n18255, ZN => 
                           n18266);
   U18857 : NAND2_X1 port map( A1 => n18258, A2 => n18257, ZN => n18259);
   U18858 : OAI211_X1 port map( C1 => n18260, C2 => n19787, A => n18259, B => 
                           n18753, ZN => n18261);
   U18859 : OAI21_X1 port map( B1 => n18263, B2 => n18262, A => n18261, ZN => 
                           n18265);
   U18860 : NOR2_X1 port map( A1 => n18752, A2 => n18264, ZN => n18758);
   U18861 : NOR2_X2 port map( A1 => n18265, A2 => n18758, ZN => n18741);
   U18862 : INV_X1 port map( A => n18741, ZN => n18783);
   U18863 : NAND2_X1 port map( A1 => n18266, A2 => n18783, ZN => n18277);
   U18864 : NAND2_X1 port map( A1 => n221, A2 => n18267, ZN => n18272);
   U18865 : NAND2_X1 port map( A1 => n18269, A2 => n18268, ZN => n18271);
   U18866 : MUX2_X1 port map( A => n18272, B => n18271, S => n18270, Z => 
                           n18719);
   U18867 : OAI211_X1 port map( C1 => n18275, C2 => n18033, A => n18274, B => 
                           n18273, ZN => n18720);
   U18868 : NAND2_X1 port map( A1 => n18719, A2 => n18720, ZN => n18775);
   U18869 : AND2_X1 port map( A1 => n18775, A2 => n18741, ZN => n18782);
   U18870 : NAND2_X1 port map( A1 => n18782, A2 => n18763, ZN => n18276);
   U18871 : INV_X1 port map( A => n18278, ZN => n18279);
   U18872 : MUX2_X1 port map( A => n18656, B => n18651, S => n19934, Z => 
                           n18283);
   U18873 : NAND3_X1 port map( A1 => n18644, A2 => n18642, A3 => n19934, ZN => 
                           n18281);
   U18874 : OAI211_X1 port map( C1 => n18283, C2 => n18644, A => n18282, B => 
                           n18281, ZN => n18285);
   U18875 : XNOR2_X1 port map( A => n18285, B => n18284, ZN => Ciphertext(62));
   U18876 : INV_X1 port map( A => n18286, ZN => n18293);
   U18877 : OAI21_X1 port map( B1 => n18289, B2 => n18288, A => n18365, ZN => 
                           n18291);
   U18878 : NAND2_X1 port map( A1 => n18290, A2 => n18359, ZN => n18360);
   U18879 : OAI211_X1 port map( C1 => n18293, C2 => n18292, A => n18291, B => 
                           n18360, ZN => n18295);
   U18880 : XNOR2_X1 port map( A => n18295, B => n18294, ZN => Ciphertext(0));
   U18881 : INV_X1 port map( A => n19163, ZN => n19154);
   U18882 : NOR2_X1 port map( A1 => n19948, A2 => n19154, ZN => n18296);
   U18883 : NOR2_X1 port map( A1 => n18296, A2 => n19683, ZN => n18303);
   U18884 : INV_X1 port map( A => n19165, ZN => n18297);
   U18885 : NAND2_X1 port map( A1 => n19948, A2 => n18297, ZN => n18302);
   U18886 : INV_X1 port map( A => n19162, ZN => n18298);
   U18887 : NAND2_X1 port map( A1 => n18298, A2 => n19163, ZN => n18300);
   U18888 : NAND3_X1 port map( A1 => n19155, A2 => n19708, A3 => n18306, ZN => 
                           n18299);
   U18889 : OAI21_X1 port map( B1 => n19948, B2 => n18300, A => n18299, ZN => 
                           n18301);
   U18890 : AOI21_X1 port map( B1 => n18303, B2 => n18302, A => n18301, ZN => 
                           n18305);
   U18891 : XNOR2_X1 port map( A => n18305, B => n18304, ZN => Ciphertext(141))
                           ;
   U18892 : NOR2_X1 port map( A1 => n19708, A2 => n19692, ZN => n18307);
   U18893 : NAND2_X1 port map( A1 => n19340, A2 => n19339, ZN => n19311);
   U18894 : INV_X1 port map( A => n19338, ZN => n19309);
   U18895 : NAND2_X1 port map( A1 => n19329, A2 => n19339, ZN => n18309);
   U18898 : NAND3_X1 port map( A1 => n19333, A2 => n19324, A3 => n19308, ZN => 
                           n18314);
   U18900 : NAND3_X1 port map( A1 => n16544, A2 => n19749, A3 => n19334, ZN => 
                           n18313);
   U18901 : INV_X1 port map( A => n2323, ZN => n18316);
   U18902 : NAND2_X1 port map( A1 => n18318, A2 => n18317, ZN => n19175);
   U18903 : NAND3_X1 port map( A1 => n18324, A2 => n20460, A3 => n18323, ZN => 
                           n18325);
   U18904 : OAI211_X1 port map( C1 => n20460, C2 => n19175, A => n18326, B => 
                           n18325, ZN => n18328);
   U18905 : XNOR2_X1 port map( A => n18328, B => n2445, ZN => Ciphertext(146));
   U18906 : NAND2_X1 port map( A1 => n18800, A2 => n18795, ZN => n18329);
   U18907 : OAI21_X1 port map( B1 => n18331, B2 => n19811, A => n18329, ZN => 
                           n18808);
   U18908 : AOI22_X1 port map( A1 => n18808, A2 => n18335, B1 => n18334, B2 => 
                           n18333, ZN => n18336);
   U18909 : XNOR2_X1 port map( A => n18336, B => n2454, ZN => Ciphertext(85));
   U18910 : NOR2_X1 port map( A1 => n19134, A2 => n870, ZN => n19148);
   U18911 : INV_X1 port map( A => n18338, ZN => n18339);
   U18913 : INV_X1 port map( A => n18341, ZN => n18343);
   U18914 : NOR2_X1 port map( A1 => n18343, A2 => n18342, ZN => n18346);
   U18915 : INV_X1 port map( A => n18359, ZN => n18345);
   U18916 : NAND4_X1 port map( A1 => n20234, A2 => n18346, A3 => n18345, A4 => 
                           n18344, ZN => n18353);
   U18917 : NAND2_X1 port map( A1 => n17936, A2 => n18348, ZN => n18351);
   U18918 : NAND3_X1 port map( A1 => n18351, A2 => n18350, A3 => n18349, ZN => 
                           n18352);
   U18919 : OAI211_X1 port map( C1 => n18365, C2 => n18354, A => n18353, B => 
                           n18352, ZN => n18356);
   U18920 : XNOR2_X1 port map( A => n18356, B => n18355, ZN => Ciphertext(3));
   U18921 : OAI21_X1 port map( B1 => n18359, B2 => n18358, A => n18357, ZN => 
                           n18361);
   U18924 : INV_X1 port map( A => n18366, ZN => n18367);
   U18925 : XNOR2_X1 port map( A => n18368, B => n18367, ZN => Ciphertext(4));
   U18926 : NOR2_X1 port map( A1 => n20361, A2 => n18382, ZN => n18369);
   U18927 : OAI21_X1 port map( B1 => n18392, B2 => n19763, A => n19501, ZN => 
                           n18371);
   U18928 : NAND2_X1 port map( A1 => n18371, A2 => n20361, ZN => n18372);
   U18929 : NAND2_X1 port map( A1 => n18373, A2 => n18372, ZN => n18375);
   U18930 : INV_X1 port map( A => n2413, ZN => n18374);
   U18931 : XNOR2_X1 port map( A => n18375, B => n18374, ZN => Ciphertext(6));
   U18933 : INV_X1 port map( A => n18392, ZN => n18383);
   U18934 : OAI21_X1 port map( B1 => n18383, B2 => n18384, A => n18381, ZN => 
                           n18378);
   U18936 : NOR2_X1 port map( A1 => n20361, A2 => n18384, ZN => n18385);
   U18937 : NAND2_X1 port map( A1 => n18385, A2 => n20437, ZN => n18386);
   U18938 : AOI21_X1 port map( B1 => n20611, B2 => n20361, A => n20437, ZN => 
                           n18395);
   U18939 : OAI22_X1 port map( A1 => n18395, A2 => n18394, B1 => n18393, B2 => 
                           n18392, ZN => n18398);
   U18940 : INV_X1 port map( A => n18396, ZN => n18397);
   U18941 : XNOR2_X1 port map( A => n18398, B => n18397, ZN => Ciphertext(11));
   U18942 : NOR2_X1 port map( A1 => n20003, A2 => n15529, ZN => n18417);
   U18943 : NAND2_X1 port map( A1 => n18417, A2 => n18407, ZN => n18403);
   U18945 : NAND2_X1 port map( A1 => n19702, A2 => n18423, ZN => n18399);
   U18947 : INV_X1 port map( A => n2394, ZN => n18405);
   U18948 : INV_X1 port map( A => n18423, ZN => n18416);
   U18949 : INV_X1 port map( A => n2382, ZN => n18410);
   U18950 : XNOR2_X1 port map( A => n18411, B => n18410, ZN => Ciphertext(13));
   U18951 : AND2_X1 port map( A1 => n18423, A2 => n18412, ZN => n18413);
   U18952 : NOR2_X1 port map( A1 => n18414, A2 => n18413, ZN => n18419);
   U18953 : AOI22_X1 port map( A1 => n18417, A2 => n18416, B1 => n18415, B2 => 
                           n18425, ZN => n18418);
   U18954 : OAI21_X1 port map( B1 => n18419, B2 => n18425, A => n18418, ZN => 
                           n18422);
   U18955 : INV_X1 port map( A => n18420, ZN => n18421);
   U18956 : XNOR2_X1 port map( A => n18422, B => n18421, ZN => Ciphertext(16));
   U18957 : NOR2_X1 port map( A1 => n18424, A2 => n18423, ZN => n18426);
   U18958 : INV_X1 port map( A => n2280, ZN => n18428);
   U18961 : OAI211_X1 port map( C1 => n18464, C2 => n18465, A => n19791, B => 
                           n20232, ZN => n18430);
   U18963 : INV_X1 port map( A => n18433, ZN => n18434);
   U18964 : XNOR2_X1 port map( A => n18435, B => n18434, ZN => Ciphertext(19));
   U18965 : INV_X1 port map( A => n18464, ZN => n18436);
   U18966 : NAND2_X1 port map( A1 => n18469, A2 => n18453, ZN => n18440);
   U18967 : OAI21_X1 port map( B1 => n18442, B2 => n18436, A => n18440, ZN => 
                           n18451);
   U18968 : INV_X1 port map( A => n18441, ZN => n18438);
   U18969 : NAND3_X1 port map( A1 => n18465, A2 => n18466, A3 => n20148, ZN => 
                           n18437);
   U18970 : OAI211_X1 port map( C1 => n18438, C2 => n18466, A => n18439, B => 
                           n18437, ZN => n18450);
   U18971 : OR2_X1 port map( A1 => n18440, A2 => n18439, ZN => n18449);
   U18972 : OAI21_X1 port map( B1 => n20139, B2 => n18468, A => n18443, ZN => 
                           n18444);
   U18973 : NAND3_X1 port map( A1 => n19825, A2 => n18446, A3 => n18445, ZN => 
                           n18448);
   U18974 : OAI211_X1 port map( C1 => n18451, C2 => n18450, A => n18449, B => 
                           n18448, ZN => Ciphertext(20));
   U18975 : OAI21_X1 port map( B1 => n18461, B2 => n18464, A => n18465, ZN => 
                           n18458);
   U18976 : NOR2_X1 port map( A1 => n20110, A2 => n18453, ZN => n18457);
   U18977 : OR3_X1 port map( A1 => n20110, A2 => n20232, A3 => n18453, ZN => 
                           n18456);
   U18978 : INV_X1 port map( A => n18468, ZN => n18463);
   U18979 : NAND3_X1 port map( A1 => n18466, A2 => n18463, A3 => n20139, ZN => 
                           n18455);
   U18980 : OAI211_X1 port map( C1 => n18458, C2 => n18457, A => n18456, B => 
                           n18455, ZN => n18460);
   U18981 : INV_X1 port map( A => n347, ZN => n18459);
   U18982 : XNOR2_X1 port map( A => n18460, B => n18459, ZN => Ciphertext(21));
   U18983 : AOI21_X1 port map( B1 => n18463, B2 => n19791, A => n18461, ZN => 
                           n18472);
   U18984 : AOI21_X1 port map( B1 => n20139, B2 => n18464, A => n20110, ZN => 
                           n18471);
   U18985 : NAND2_X1 port map( A1 => n18469, A2 => n20148, ZN => n18470);
   U18986 : XNOR2_X1 port map( A => n18474, B => n18473, ZN => Ciphertext(22));
   U18987 : NOR3_X1 port map( A1 => n18485, A2 => n18500, A3 => n18478, ZN => 
                           n18475);
   U18988 : OAI21_X1 port map( B1 => n18497, B2 => n18498, A => n18475, ZN => 
                           n18477);
   U18989 : INV_X1 port map( A => n18478, ZN => n18481);
   U18990 : NOR2_X1 port map( A1 => n18498, A2 => n18481, ZN => n18486);
   U18991 : NAND2_X1 port map( A1 => n18486, A2 => n19816, ZN => n18476);
   U18992 : NAND2_X1 port map( A1 => n18477, A2 => n18476, ZN => n18494);
   U18993 : NAND3_X1 port map( A1 => n18500, A2 => n18478, A3 => n17640, ZN => 
                           n18484);
   U18994 : OR2_X1 port map( A1 => n18498, A2 => n18478, ZN => n18487);
   U18995 : NAND3_X1 port map( A1 => n18495, A2 => n18478, A3 => n18498, ZN => 
                           n18479);
   U18996 : NAND2_X1 port map( A1 => n18487, A2 => n18479, ZN => n18480);
   U18997 : NAND2_X1 port map( A1 => n18480, A2 => n893, ZN => n18483);
   U18998 : NAND3_X1 port map( A1 => n18496, A2 => n893, A3 => n18481, ZN => 
                           n18482);
   U18999 : NAND3_X1 port map( A1 => n18484, A2 => n18483, A3 => n18482, ZN => 
                           n18493);
   U19000 : NAND3_X1 port map( A1 => n18486, A2 => n18501, A3 => n893, ZN => 
                           n18492);
   U19001 : INV_X1 port map( A => n18487, ZN => n18488);
   U19002 : NAND3_X1 port map( A1 => n19729, A2 => n19816, A3 => n18488, ZN => 
                           n18491);
   U19003 : OAI211_X1 port map( C1 => n18494, C2 => n18493, A => n18492, B => 
                           n18491, ZN => Ciphertext(25));
   U19004 : AOI22_X1 port map( A1 => n18500, A2 => n17640, B1 => n18495, B2 => 
                           n18498, ZN => n18502);
   U19005 : OAI21_X1 port map( B1 => n214, B2 => n18517, A => n18518, ZN => 
                           n18528);
   U19006 : NAND2_X1 port map( A1 => n19773, A2 => n18517, ZN => n18510);
   U19007 : NAND2_X1 port map( A1 => n20492, A2 => n18517, ZN => n18507);
   U19008 : NAND2_X1 port map( A1 => n19526, A2 => n18507, ZN => n18509);
   U19009 : OAI21_X1 port map( B1 => n20433, B2 => n18510, A => n18509, ZN => 
                           n18527);
   U19010 : NAND2_X1 port map( A1 => n19758, A2 => Key(124), ZN => n18514);
   U19011 : OR2_X1 port map( A1 => n19773, A2 => n20492, ZN => n18523);
   U19012 : XNOR2_X1 port map( A => n18512, B => n18517, ZN => n18513);
   U19013 : OAI22_X1 port map( A1 => n18514, A2 => n18523, B1 => n18513, B2 => 
                           n19758, ZN => n18515);
   U19014 : NAND2_X1 port map( A1 => n18515, A2 => n18504, ZN => n18526);
   U19015 : OR2_X1 port map( A1 => n19773, A2 => Key(124), ZN => n18520);
   U19016 : INV_X1 port map( A => n18520, ZN => n18524);
   U19017 : OAI22_X1 port map( A1 => n18520, A2 => n20492, B1 => n19758, B2 => 
                           n18517, ZN => n18521);
   U19018 : OAI211_X1 port map( C1 => n18524, C2 => n18523, A => n18522, B => 
                           n18521, ZN => n18525);
   U19019 : OAI211_X1 port map( C1 => n18528, C2 => n18527, A => n18526, B => 
                           n18525, ZN => Ciphertext(33));
   U19020 : NAND2_X1 port map( A1 => n18529, A2 => n19682, ZN => n18553);
   U19021 : AOI22_X1 port map( A1 => n18532, A2 => n18531, B1 => n18553, B2 => 
                           n18530, ZN => n18533);
   U19022 : XNOR2_X1 port map( A => n18533, B => n2233, ZN => Ciphertext(37));
   U19023 : MUX2_X1 port map( A => n18535, B => n17564, S => n20432, Z => 
                           n18536);
   U19024 : NAND2_X1 port map( A1 => n18539, A2 => n18536, ZN => n18537);
   U19025 : OAI21_X1 port map( B1 => n18539, B2 => n18538, A => n18537, ZN => 
                           n18543);
   U19026 : NAND4_X1 port map( A1 => n18543, A2 => n18542, A3 => n18541, A4 => 
                           n18540, ZN => n18549);
   U19027 : NAND2_X1 port map( A1 => n18543, A2 => n18542, ZN => n18544);
   U19028 : OAI21_X1 port map( B1 => n19682, B2 => n18545, A => n18544, ZN => 
                           n18548);
   U19029 : NAND2_X1 port map( A1 => n19682, A2 => n19691, ZN => n18547);
   U19030 : OAI211_X1 port map( C1 => n19682, C2 => n18549, A => n18548, B => 
                           n18547, ZN => n18551);
   U19031 : OAI21_X1 port map( B1 => n18553, B2 => n18552, A => n18551, ZN => 
                           n18554);
   U19032 : XNOR2_X1 port map( A => n18554, B => Key(63), ZN => Ciphertext(38))
                           ;
   U19033 : NOR2_X1 port map( A1 => n18555, A2 => n18568, ZN => n18558);
   U19034 : NOR2_X1 port map( A1 => n18565, A2 => n18556, ZN => n18557);
   U19035 : MUX2_X1 port map( A => n18558, B => n18557, S => n18567, Z => 
                           n18563);
   U19036 : OAI22_X1 port map( A1 => n18561, A2 => n18566, B1 => n18560, B2 => 
                           n18559, ZN => n18562);
   U19037 : NOR2_X1 port map( A1 => n18563, A2 => n18562, ZN => n18564);
   U19038 : XNOR2_X1 port map( A => n18564, B => n404, ZN => Ciphertext(45));
   U19039 : OAI21_X1 port map( B1 => n19775, B2 => n18566, A => n18565, ZN => 
                           n18569);
   U19040 : AOI22_X1 port map( A1 => n18571, A2 => n18570, B1 => n18569, B2 => 
                           n18568, ZN => n18572);
   U19041 : XNOR2_X1 port map( A => n18572, B => n2349, ZN => Ciphertext(47));
   U19042 : NAND2_X1 port map( A1 => n18573, A2 => n18597, ZN => n18579);
   U19043 : NOR2_X1 port map( A1 => n20445, A2 => n18597, ZN => n18576);
   U19044 : NOR2_X1 port map( A1 => n20365, A2 => n19656, ZN => n18575);
   U19045 : NAND3_X1 port map( A1 => n20445, A2 => n18589, A3 => n19669, ZN => 
                           n18578);
   U19046 : XNOR2_X1 port map( A => n18580, B => n2344, ZN => Ciphertext(50));
   U19047 : INV_X1 port map( A => n18597, ZN => n18583);
   U19048 : NOR2_X1 port map( A1 => n20445, A2 => n19656, ZN => n18581);
   U19049 : NAND2_X1 port map( A1 => n18581, A2 => n19665, ZN => n18582);
   U19050 : OAI211_X1 port map( C1 => n18589, C2 => n20445, A => n18584, B => 
                           n18583, ZN => n18586);
   U19051 : OAI21_X1 port map( B1 => n18590, B2 => n18589, A => n19656, ZN => 
                           n18591);
   U19052 : NAND2_X1 port map( A1 => n18597, A2 => n18591, ZN => n18595);
   U19053 : NAND2_X1 port map( A1 => n18593, A2 => n18592, ZN => n18594);
   U19054 : OAI211_X1 port map( C1 => n18597, C2 => n18596, A => n18595, B => 
                           n18594, ZN => n18599);
   U19055 : XNOR2_X1 port map( A => n18599, B => n18598, ZN => Ciphertext(53));
   U19056 : NAND2_X1 port map( A1 => n19679, A2 => n2248, ZN => n18606);
   U19057 : INV_X1 port map( A => n2248, ZN => n18610);
   U19058 : AND3_X1 port map( A1 => n18622, A2 => n18610, A3 => n19679, ZN => 
                           n18607);
   U19059 : OR2_X1 port map( A1 => n18620, A2 => n18610, ZN => n18612);
   U19060 : NOR2_X1 port map( A1 => n18612, A2 => n18600, ZN => n18601);
   U19061 : OAI21_X1 port map( B1 => n18607, B2 => n18601, A => n18626, ZN => 
                           n18605);
   U19062 : NAND3_X1 port map( A1 => n18603, A2 => n19509, A3 => n18610, ZN => 
                           n18604);
   U19063 : OAI211_X1 port map( C1 => n19673, C2 => n18606, A => n18605, B => 
                           n18604, ZN => n18618);
   U19064 : INV_X1 port map( A => n18607, ZN => n18609);
   U19065 : NAND3_X1 port map( A1 => n18619, A2 => n2248, A3 => n18613, ZN => 
                           n18608);
   U19066 : OAI21_X1 port map( B1 => n18619, B2 => n18609, A => n18608, ZN => 
                           n18617);
   U19068 : NAND4_X1 port map( A1 => n19877, A2 => n18619, A3 => n18610, A4 => 
                           n18613, ZN => n18616);
   U19069 : INV_X1 port map( A => n18612, ZN => n18614);
   U19070 : NAND3_X1 port map( A1 => n20188, A2 => n18614, A3 => n18613, ZN => 
                           n18615);
   U19071 : OAI211_X1 port map( C1 => n18618, C2 => n18617, A => n18616, B => 
                           n18615, ZN => Ciphertext(55));
   U19072 : NOR2_X1 port map( A1 => n18621, A2 => n19679, ZN => n18623);
   U19073 : NOR2_X1 port map( A1 => n18623, A2 => n18622, ZN => n18624);
   U19074 : OAI21_X1 port map( B1 => n18626, B2 => n18625, A => n18624, ZN => 
                           n18627);
   U19075 : OAI211_X1 port map( C1 => n20188, C2 => n18629, A => n18628, B => 
                           n18627, ZN => n18632);
   U19076 : XNOR2_X1 port map( A => n18632, B => n18631, ZN => Ciphertext(57));
   U19078 : NOR2_X1 port map( A1 => n18634, A2 => n18633, ZN => n18638);
   U19079 : NOR2_X1 port map( A1 => n18636, A2 => n20349, ZN => n18637);
   U19080 : OAI211_X1 port map( C1 => n18644, C2 => n19745, A => n18639, B => 
                           n19934, ZN => n18640);
   U19081 : NOR2_X1 port map( A1 => n18644, A2 => n18648, ZN => n18659);
   U19082 : NAND2_X1 port map( A1 => n18656, A2 => n19934, ZN => n18646);
   U19085 : NOR2_X1 port map( A1 => n19935, A2 => n18650, ZN => n18655);
   U19086 : NOR2_X1 port map( A1 => n19934, A2 => n18651, ZN => n18653);
   U19089 : XNOR2_X1 port map( A => n18661, B => n18660, ZN => Ciphertext(63));
   U19090 : INV_X1 port map( A => n18679, ZN => n18663);
   U19091 : NOR2_X1 port map( A1 => n18672, A2 => n18671, ZN => n18684);
   U19092 : NOR2_X1 port map( A1 => n18684, A2 => n19735, ZN => n18662);
   U19093 : NAND2_X1 port map( A1 => n18686, A2 => n18672, ZN => n18675);
   U19094 : OAI22_X1 port map( A1 => n18663, A2 => n18662, B1 => n18669, B2 => 
                           n18675, ZN => n18665);
   U19095 : XNOR2_X1 port map( A => n18665, B => n18664, ZN => Ciphertext(67));
   U19096 : NOR2_X1 port map( A1 => n18688, A2 => n18666, ZN => n18668);
   U19097 : NAND3_X1 port map( A1 => n19510, A2 => n18671, A3 => n18686, ZN => 
                           n18678);
   U19098 : NOR2_X1 port map( A1 => n18673, A2 => n18672, ZN => n18674);
   U19099 : NOR2_X1 port map( A1 => n18688, A2 => n18674, ZN => n18676);
   U19100 : NAND2_X1 port map( A1 => n18676, A2 => n18675, ZN => n18677);
   U19101 : OAI211_X1 port map( C1 => n18682, C2 => n18679, A => n18678, B => 
                           n18677, ZN => n18680);
   U19102 : XNOR2_X1 port map( A => n18680, B => n1781, ZN => Ciphertext(69));
   U19103 : NOR2_X1 port map( A1 => n18688, A2 => n19510, ZN => n18685);
   U19104 : INV_X1 port map( A => n18682, ZN => n18683);
   U19105 : OAI21_X1 port map( B1 => n18685, B2 => n18684, A => n18683, ZN => 
                           n18690);
   U19106 : OAI21_X1 port map( B1 => n18686, B2 => n18672, A => n17964, ZN => 
                           n18687);
   U19107 : NAND2_X1 port map( A1 => n18688, A2 => n18687, ZN => n18689);
   U19108 : NAND2_X1 port map( A1 => n18690, A2 => n18689, ZN => n18693);
   U19110 : XNOR2_X1 port map( A => n18693, B => n19640, ZN => Ciphertext(71));
   U19111 : AND2_X1 port map( A1 => n18698, A2 => n18703, ZN => n18699);
   U19112 : NAND2_X1 port map( A1 => n18072, A2 => n18702, ZN => n18694);
   U19113 : AOI22_X1 port map( A1 => n18695, A2 => n18706, B1 => n18699, B2 => 
                           n18694, ZN => n18696);
   U19114 : XNOR2_X1 port map( A => n18696, B => n2222, ZN => Ciphertext(73));
   U19115 : OAI21_X1 port map( B1 => n18698, B2 => n19753, A => n18697, ZN => 
                           n18700);
   U19116 : NAND3_X1 port map( A1 => n19751, A2 => n18702, A3 => n18701, ZN => 
                           n18704);
   U19117 : OAI211_X1 port map( C1 => n18072, C2 => n18706, A => n18705, B => 
                           n18704, ZN => n18708);
   U19118 : INV_X1 port map( A => n2376, ZN => n18707);
   U19119 : XNOR2_X1 port map( A => n18708, B => n18707, ZN => Ciphertext(75));
   U19120 : AND2_X1 port map( A1 => n18775, A2 => n18709, ZN => n18761);
   U19121 : NAND2_X1 port map( A1 => n18761, A2 => n19803, ZN => n18715);
   U19123 : NAND2_X1 port map( A1 => n18746, A2 => n18781, ZN => n18714);
   U19124 : INV_X1 port map( A => n18775, ZN => n18711);
   U19127 : INV_X1 port map( A => n18716, ZN => n18717);
   U19129 : NOR2_X1 port map( A1 => n18774, A2 => n18762, ZN => n18771);
   U19130 : NAND2_X1 port map( A1 => n18771, A2 => n18763, ZN => n18725);
   U19131 : AND2_X1 port map( A1 => n18781, A2 => n18741, ZN => n18776);
   U19132 : INV_X1 port map( A => n18776, ZN => n18724);
   U19133 : NAND4_X1 port map( A1 => n18719, A2 => n18722, A3 => n18721, A4 => 
                           n18720, ZN => n18728);
   U19134 : NAND3_X1 port map( A1 => n18774, A2 => n18773, A3 => n18728, ZN => 
                           n18723);
   U19135 : NAND4_X1 port map( A1 => n18725, A2 => n18726, A3 => n18724, A4 => 
                           n18723, ZN => n18732);
   U19136 : INV_X1 port map( A => n18726, ZN => n18727);
   U19137 : NAND2_X1 port map( A1 => n18776, A2 => n18727, ZN => n18731);
   U19138 : NAND4_X1 port map( A1 => n18763, A2 => n18772, A3 => n18727, A4 => 
                           n18749, ZN => n18730);
   U19139 : NAND4_X1 port map( A1 => n18728, A2 => n18774, A3 => n18773, A4 => 
                           n18727, ZN => n18729);
   U19140 : NAND4_X1 port map( A1 => n18732, A2 => n18731, A3 => n18730, A4 => 
                           n18729, ZN => Ciphertext(79));
   U19141 : INV_X1 port map( A => n2381, ZN => n18743);
   U19142 : AND2_X1 port map( A1 => n18773, A2 => n18743, ZN => n18733);
   U19143 : NAND3_X1 port map( A1 => n18733, A2 => n18781, A3 => n18772, ZN => 
                           n18737);
   U19146 : NAND3_X1 port map( A1 => n18762, A2 => n18773, A3 => n2381, ZN => 
                           n18735);
   U19151 : NAND2_X1 port map( A1 => n18741, A2 => n18773, ZN => n18742);
   U19152 : NAND3_X1 port map( A1 => n18763, A2 => n2381, A3 => n18742, ZN => 
                           n18745);
   U19153 : NAND3_X1 port map( A1 => n18746, A2 => n18763, A3 => n18743, ZN => 
                           n18744);
   U19154 : OAI21_X1 port map( B1 => n18746, B2 => n18745, A => n18744, ZN => 
                           n18747);
   U19156 : NAND2_X1 port map( A1 => n18750, A2 => n18753, ZN => n18751);
   U19157 : NAND2_X1 port map( A1 => n18752, A2 => n18751, ZN => n18757);
   U19158 : NAND2_X1 port map( A1 => n18754, A2 => n18753, ZN => n18756);
   U19159 : MUX2_X1 port map( A => n18757, B => n18756, S => n20438, Z => 
                           n18760);
   U19160 : INV_X1 port map( A => n18758, ZN => n18759);
   U19161 : NAND2_X1 port map( A1 => n18760, A2 => n18759, ZN => n18766);
   U19162 : NAND2_X1 port map( A1 => n18766, A2 => n18761, ZN => n18765);
   U19163 : NAND3_X1 port map( A1 => n18763, A2 => n18773, A3 => n18762, ZN => 
                           n18764);
   U19164 : OAI211_X1 port map( C1 => n18767, C2 => n18766, A => n18765, B => 
                           n18764, ZN => n18770);
   U19165 : INV_X1 port map( A => n18768, ZN => n18769);
   U19166 : XNOR2_X1 port map( A => n18770, B => n18769, ZN => Ciphertext(81));
   U19167 : NAND2_X1 port map( A1 => n18771, A2 => n18775, ZN => n18780);
   U19168 : OAI21_X1 port map( B1 => n18774, B2 => n18773, A => n18772, ZN => 
                           n18785);
   U19169 : NAND2_X1 port map( A1 => n18785, A2 => n18783, ZN => n18778);
   U19170 : NAND2_X1 port map( A1 => n18776, A2 => n18775, ZN => n18777);
   U19171 : NAND4_X1 port map( A1 => n18780, A2 => n18779, A3 => n18778, A4 => 
                           n18777, ZN => n18789);
   U19172 : OR2_X1 port map( A1 => n18780, A2 => n18779, ZN => n18788);
   U19173 : NAND3_X1 port map( A1 => n18782, A2 => n18784, A3 => n18781, ZN => 
                           n18787);
   U19174 : NAND3_X1 port map( A1 => n18785, A2 => n18784, A3 => n18783, ZN => 
                           n18786);
   U19175 : NAND4_X1 port map( A1 => n18789, A2 => n18788, A3 => n18787, A4 => 
                           n18786, ZN => Ciphertext(83));
   U19176 : MUX2_X1 port map( A => n18794, B => n18807, S => n19770, Z => 
                           n18791);
   U19177 : NAND2_X1 port map( A1 => n18794, A2 => n17772, ZN => n18804);
   U19178 : OAI21_X1 port map( B1 => n19711, B2 => n18331, A => n18804, ZN => 
                           n18790);
   U19179 : MUX2_X1 port map( A => n18791, B => n18790, S => n18795, Z => 
                           n18793);
   U19180 : XNOR2_X1 port map( A => n18793, B => n18792, ZN => Ciphertext(86));
   U19181 : MUX2_X1 port map( A => n17772, B => n19711, S => n18803, Z => 
                           n18799);
   U19182 : NAND2_X1 port map( A1 => n18807, A2 => n18800, ZN => n18797);
   U19183 : NAND2_X1 port map( A1 => n18794, A2 => n18803, ZN => n18796);
   U19184 : OAI21_X1 port map( B1 => n18800, B2 => n18799, A => n18798, ZN => 
                           n18802);
   U19185 : XNOR2_X1 port map( A => n18802, B => n296, ZN => Ciphertext(88));
   U19186 : NAND2_X1 port map( A1 => n18804, A2 => n18803, ZN => n18805);
   U19187 : AOI22_X1 port map( A1 => n18808, A2 => n18807, B1 => n19770, B2 => 
                           n18805, ZN => n18810);
   U19188 : XNOR2_X1 port map( A => n18810, B => n18809, ZN => Ciphertext(89));
   U19189 : NAND3_X1 port map( A1 => n20130, A2 => n18172, A3 => n20276, ZN => 
                           n18816);
   U19190 : NAND3_X1 port map( A1 => n18814, A2 => n18813, A3 => n18812, ZN => 
                           n18815);
   U19191 : OAI211_X1 port map( C1 => n18818, C2 => n18817, A => n18815, B => 
                           n18816, ZN => n18820);
   U19192 : XNOR2_X1 port map( A => n18820, B => n1783, ZN => Ciphertext(93));
   U19193 : XNOR2_X1 port map( A => n19766, B => n18830, ZN => n18822);
   U19194 : NAND3_X1 port map( A1 => n18822, A2 => n20276, A3 => n19794, ZN => 
                           n18839);
   U19195 : AND2_X1 port map( A1 => n18172, A2 => n18830, ZN => n18829);
   U19196 : NOR2_X1 port map( A1 => n19890, A2 => n18830, ZN => n18823);
   U19197 : AOI21_X1 port map( B1 => n18829, B2 => n19890, A => n18823, ZN => 
                           n18826);
   U19198 : NOR2_X1 port map( A1 => n18172, A2 => n18830, ZN => n18835);
   U19199 : NOR2_X1 port map( A1 => n19794, A2 => n18835, ZN => n18825);
   U19200 : OAI211_X1 port map( C1 => n20130, C2 => n18827, A => n18826, B => 
                           n18825, ZN => n18838);
   U19201 : NOR2_X1 port map( A1 => n20422, A2 => n18830, ZN => n18832);
   U19202 : INV_X1 port map( A => n18831, ZN => n18840);
   U19203 : OAI211_X1 port map( C1 => n18833, C2 => n18832, A => n18840, B => 
                           n19794, ZN => n18837);
   U19204 : NAND3_X1 port map( A1 => n18840, A2 => n18835, A3 => n18834, ZN => 
                           n18836);
   U19205 : NAND4_X1 port map( A1 => n18839, A2 => n18838, A3 => n18837, A4 => 
                           n18836, ZN => Ciphertext(94));
   U19206 : NAND2_X1 port map( A1 => n18841, A2 => n18840, ZN => n18843);
   U19207 : AOI22_X1 port map( A1 => n18845, A2 => n19890, B1 => n18843, B2 => 
                           n19794, ZN => n18846);
   U19208 : XNOR2_X1 port map( A => n18846, B => n2108, ZN => Ciphertext(95));
   U19210 : AOI21_X1 port map( B1 => n19917, B2 => n19988, A => n18850, ZN => 
                           n18847);
   U19211 : INV_X1 port map( A => n18848, ZN => n18849);
   U19212 : OAI21_X1 port map( B1 => n18871, B2 => n18853, A => n18852, ZN => 
                           n18856);
   U19213 : INV_X1 port map( A => n18854, ZN => n18855);
   U19214 : XNOR2_X1 port map( A => n18856, B => n18855, ZN => Ciphertext(97));
   U19215 : NAND2_X1 port map( A1 => n18857, A2 => n20259, ZN => n18860);
   U19216 : OR2_X1 port map( A1 => n3030, A2 => n19988, ZN => n18859);
   U19217 : OAI21_X1 port map( B1 => n18862, B2 => n20259, A => n18861, ZN => 
                           n18865);
   U19218 : INV_X1 port map( A => n18863, ZN => n18864);
   U19219 : XNOR2_X1 port map( A => n18865, B => n18864, ZN => Ciphertext(100))
                           ;
   U19220 : AOI21_X1 port map( B1 => n20418, B2 => n20117, A => n20259, ZN => 
                           n18870);
   U19221 : OAI22_X1 port map( A1 => n18871, A2 => n3030, B1 => n18870, B2 => 
                           n18869, ZN => n18873);
   U19222 : INV_X1 port map( A => n2164, ZN => n18872);
   U19223 : XNOR2_X1 port map( A => n18873, B => n18872, ZN => Ciphertext(101))
                           ;
   U19224 : INV_X1 port map( A => n18921, ZN => n18898);
   U19225 : NAND2_X1 port map( A1 => n19874, A2 => n18876, ZN => n18879);
   U19226 : NAND2_X1 port map( A1 => n18899, A2 => n18916, ZN => n18901);
   U19227 : NOR2_X1 port map( A1 => n18901, A2 => n19681, ZN => n18875);
   U19228 : NOR2_X1 port map( A1 => n18875, A2 => n18874, ZN => n18878);
   U19229 : NAND3_X1 port map( A1 => n18897, A2 => n19681, A3 => n18876, ZN => 
                           n18877);
   U19230 : OAI211_X1 port map( C1 => n18898, C2 => n18879, A => n18878, B => 
                           n18877, ZN => n18881);
   U19231 : XNOR2_X1 port map( A => n18881, B => n18880, ZN => Ciphertext(102))
                           ;
   U19232 : INV_X1 port map( A => n18899, ZN => n18882);
   U19233 : INV_X1 port map( A => n18918, ZN => n18886);
   U19234 : AND2_X1 port map( A1 => n17054, A2 => n18897, ZN => n18917);
   U19235 : NAND2_X1 port map( A1 => n18917, A2 => n18882, ZN => n18885);
   U19236 : INV_X1 port map( A => n18897, ZN => n18883);
   U19237 : OAI211_X1 port map( C1 => n19664, C2 => n19874, A => n18883, B => 
                           n19681, ZN => n18884);
   U19238 : NAND3_X1 port map( A1 => n18886, A2 => n18885, A3 => n18884, ZN => 
                           n18889);
   U19239 : INV_X1 port map( A => n18887, ZN => n18888);
   U19240 : XNOR2_X1 port map( A => n18889, B => n18888, ZN => Ciphertext(103))
                           ;
   U19241 : MUX2_X1 port map( A => n18890, B => n18916, S => n18921, Z => 
                           n18893);
   U19242 : NAND2_X1 port map( A1 => n18897, A2 => n18890, ZN => n18919);
   U19243 : NAND2_X1 port map( A1 => n18919, A2 => n18891, ZN => n18892);
   U19244 : MUX2_X1 port map( A => n18893, B => n18892, S => n19874, Z => 
                           n18895);
   U19245 : INV_X1 port map( A => n2446, ZN => n18894);
   U19246 : XNOR2_X1 port map( A => n18895, B => n18894, ZN => Ciphertext(104))
                           ;
   U19247 : NAND2_X1 port map( A1 => n19874, A2 => n18897, ZN => n18896);
   U19248 : OAI21_X1 port map( B1 => n19681, B2 => n18897, A => n18896, ZN => 
                           n18911);
   U19249 : NAND2_X1 port map( A1 => n18898, A2 => n18911, ZN => n18904);
   U19250 : NOR2_X1 port map( A1 => n19905, A2 => n19874, ZN => n18907);
   U19251 : AOI21_X1 port map( B1 => n18907, B2 => n19681, A => n18909, ZN => 
                           n18903);
   U19252 : INV_X1 port map( A => n18901, ZN => n18902);
   U19253 : NAND2_X1 port map( A1 => n18921, A2 => n18902, ZN => n18905);
   U19254 : NAND3_X1 port map( A1 => n18904, A2 => n18903, A3 => n18905, ZN => 
                           n18915);
   U19255 : INV_X1 port map( A => n18905, ZN => n18910);
   U19256 : NOR2_X1 port map( A1 => n18890, A2 => n2203, ZN => n18908);
   U19257 : AOI22_X1 port map( A1 => n18910, A2 => n18909, B1 => n18908, B2 => 
                           n18907, ZN => n18914);
   U19258 : NOR2_X1 port map( A1 => n18921, A2 => n2203, ZN => n18912);
   U19259 : NAND2_X1 port map( A1 => n18912, A2 => n18911, ZN => n18913);
   U19260 : NAND3_X1 port map( A1 => n18915, A2 => n18914, A3 => n18913, ZN => 
                           Ciphertext(105));
   U19261 : OAI21_X1 port map( B1 => n18918, B2 => n18917, A => n19664, ZN => 
                           n18923);
   U19262 : NAND2_X1 port map( A1 => n18919, A2 => n19905, ZN => n18920);
   U19263 : XNOR2_X1 port map( A => n18925, B => n18924, ZN => Ciphertext(107))
                           ;
   U19264 : NAND2_X1 port map( A1 => n18932, A2 => n18926, ZN => n18930);
   U19265 : NAND2_X1 port map( A1 => n20501, A2 => n18937, ZN => n18943);
   U19266 : NAND2_X1 port map( A1 => n18940, A2 => n18939, ZN => n18942);
   U19267 : MUX2_X1 port map( A => n18943, B => n18942, S => n18941, Z => 
                           n18944);
   U19268 : NOR2_X1 port map( A1 => n2058, A2 => n19654, ZN => n18974);
   U19269 : MUX2_X1 port map( A => n18948, B => n19916, S => n18946, Z => 
                           n18952);
   U19270 : MUX2_X1 port map( A => n18950, B => n18949, S => n17687, Z => 
                           n18951);
   U19271 : AOI22_X1 port map( A1 => n219, A2 => n18954, B1 => n18955, B2 => 
                           n18953, ZN => n18960);
   U19272 : OR2_X1 port map( A1 => n20221, A2 => n18955, ZN => n18958);
   U19274 : INV_X1 port map( A => n18961, ZN => n18963);
   U19275 : NAND2_X1 port map( A1 => n18963, A2 => n18962, ZN => n18964);
   U19276 : AND2_X1 port map( A1 => n18965, A2 => n18964, ZN => n18973);
   U19277 : INV_X1 port map( A => n18966, ZN => n18967);
   U19278 : OR2_X1 port map( A1 => n19684, A2 => n18967, ZN => n18971);
   U19279 : MUX2_X1 port map( A => n18971, B => n18970, S => n20127, Z => 
                           n18972);
   U19280 : OAI21_X1 port map( B1 => n18973, B2 => n220, A => n18972, ZN => 
                           n19011);
   U19281 : INV_X1 port map( A => n19680, ZN => n19025);
   U19282 : OAI21_X1 port map( B1 => n18974, B2 => n19004, A => n19025, ZN => 
                           n18983);
   U19283 : MUX2_X1 port map( A => n18976, B => n20158, S => n18978, Z => 
                           n18981);
   U19284 : AOI21_X1 port map( B1 => n18981, B2 => n18980, A => n18979, ZN => 
                           n19002);
   U19285 : AND2_X1 port map( A1 => n19001, A2 => n19002, ZN => n19010);
   U19286 : INV_X1 port map( A => n19010, ZN => n19015);
   U19288 : INV_X1 port map( A => n18984, ZN => n18985);
   U19289 : NOR2_X1 port map( A1 => n19011, A2 => n19687, ZN => n18995);
   U19291 : NAND2_X1 port map( A1 => n2058, A2 => n19724, ZN => n18987);
   U19292 : INV_X1 port map( A => n19021, ZN => n18986);
   U19293 : AOI22_X1 port map( A1 => n18986, A2 => n19687, B1 => n19013, B2 => 
                           n19002, ZN => n19026);
   U19294 : OAI22_X1 port map( A1 => n18995, A2 => n18987, B1 => n19026, B2 => 
                           n19004, ZN => n18990);
   U19295 : INV_X1 port map( A => n18988, ZN => n18989);
   U19296 : XNOR2_X1 port map( A => n18990, B => n18989, ZN => Ciphertext(109))
                           ;
   U19297 : INV_X1 port map( A => n19023, ZN => n18994);
   U19298 : INV_X1 port map( A => n19009, ZN => n18999);
   U19299 : NAND2_X1 port map( A1 => n18999, A2 => n19654, ZN => n18993);
   U19300 : NAND2_X1 port map( A1 => n18999, A2 => n19867, ZN => n18991);
   U19301 : NAND2_X1 port map( A1 => n18995, A2 => n19866, ZN => n18996);
   U19302 : XNOR2_X1 port map( A => n18998, B => n18997, ZN => Ciphertext(110))
                           ;
   U19303 : NOR2_X1 port map( A1 => n19687, A2 => n19654, ZN => n19003);
   U19304 : INV_X1 port map( A => n19002, ZN => n19022);
   U19305 : AOI22_X1 port map( A1 => n19004, A2 => n19680, B1 => n19003, B2 => 
                           n19022, ZN => n19005);
   U19306 : OAI21_X1 port map( B1 => n19006, B2 => n19866, A => n19005, ZN => 
                           n19008);
   U19307 : XNOR2_X1 port map( A => n19008, B => n19007, ZN => Ciphertext(111))
                           ;
   U19308 : NOR2_X1 port map( A1 => n19687, A2 => n19866, ZN => n19012);
   U19309 : AOI22_X1 port map( A1 => n19012, A2 => n19680, B1 => n19010, B2 => 
                           n19687, ZN => n19017);
   U19310 : NAND2_X1 port map( A1 => n19013, A2 => n19022, ZN => n19014);
   U19311 : NAND3_X1 port map( A1 => n19015, A2 => n19014, A3 => n19867, ZN => 
                           n19016);
   U19312 : NAND2_X1 port map( A1 => n19017, A2 => n19016, ZN => n19020);
   U19313 : INV_X1 port map( A => n19018, ZN => n19019);
   U19314 : XNOR2_X1 port map( A => n19020, B => n19019, ZN => Ciphertext(112))
                           ;
   U19315 : OAI21_X1 port map( B1 => n19023, B2 => n19022, A => n19867, ZN => 
                           n19024);
   U19316 : OAI21_X1 port map( B1 => n19026, B2 => n19025, A => n19024, ZN => 
                           n19029);
   U19317 : INV_X1 port map( A => n19027, ZN => n19028);
   U19318 : XNOR2_X1 port map( A => n19029, B => n19028, ZN => Ciphertext(113))
                           ;
   U19320 : NOR2_X1 port map( A1 => n19046, A2 => n19032, ZN => n19033);
   U19321 : AOI21_X1 port map( B1 => n20475, B2 => n19034, A => n19047, ZN => 
                           n19036);
   U19322 : NAND2_X1 port map( A1 => n19036, A2 => n19035, ZN => n19037);
   U19323 : XNOR2_X1 port map( A => n19039, B => n19038, ZN => Ciphertext(117))
                           ;
   U19324 : NOR2_X1 port map( A1 => n20475, A2 => n19993, ZN => n19042);
   U19325 : AND2_X1 port map( A1 => n19992, A2 => n19047, ZN => n19041);
   U19326 : OAI21_X1 port map( B1 => n19042, B2 => n19041, A => n19046, ZN => 
                           n19051);
   U19327 : INV_X1 port map( A => n19047, ZN => n19045);
   U19328 : NAND3_X1 port map( A1 => n19045, A2 => n20475, A3 => n20142, ZN => 
                           n19050);
   U19329 : INV_X1 port map( A => n19046, ZN => n19048);
   U19330 : NAND3_X1 port map( A1 => n19048, A2 => n18061, A3 => n19047, ZN => 
                           n19049);
   U19331 : NAND3_X1 port map( A1 => n19051, A2 => n19050, A3 => n19049, ZN => 
                           n19054);
   U19332 : INV_X1 port map( A => n19052, ZN => n19053);
   U19333 : XNOR2_X1 port map( A => n19054, B => n19053, ZN => Ciphertext(118))
                           ;
   U19334 : INV_X1 port map( A => n19073, ZN => n19076);
   U19335 : OAI21_X1 port map( B1 => n19076, B2 => n20131, A => n19055, ZN => 
                           n19057);
   U19336 : INV_X1 port map( A => n19067, ZN => n19077);
   U19337 : NAND3_X1 port map( A1 => n19069, A2 => n20131, A3 => n19077, ZN => 
                           n19056);
   U19338 : NAND2_X1 port map( A1 => n19058, A2 => n19076, ZN => n19063);
   U19339 : INV_X1 port map( A => n19079, ZN => n19062);
   U19340 : NAND3_X1 port map( A1 => n19653, A2 => n19073, A3 => n19059, ZN => 
                           n19061);
   U19341 : OAI211_X1 port map( C1 => n19064, C2 => n19063, A => n19062, B => 
                           n19061, ZN => n19066);
   U19342 : INV_X1 port map( A => n2384, ZN => n19065);
   U19343 : XNOR2_X1 port map( A => n19066, B => n19065, ZN => Ciphertext(121))
                           ;
   U19344 : INV_X1 port map( A => n19068, ZN => n19082);
   U19345 : AOI21_X1 port map( B1 => n19075, B2 => n19073, A => n19082, ZN => 
                           n19072);
   U19346 : NOR2_X1 port map( A1 => n19685, A2 => n19067, ZN => n19070);
   U19347 : AOI21_X1 port map( B1 => n20131, B2 => n19073, A => n19075, ZN => 
                           n19081);
   U19348 : NOR2_X1 port map( A1 => n19076, A2 => n19075, ZN => n19078);
   U19349 : OAI21_X1 port map( B1 => n19079, B2 => n19078, A => n19077, ZN => 
                           n19080);
   U19350 : XNOR2_X1 port map( A => n19084, B => n19083, ZN => Ciphertext(125))
                           ;
   U19351 : NOR2_X1 port map( A1 => n19105, A2 => n19112, ZN => n19090);
   U19352 : INV_X1 port map( A => n19085, ZN => n19086);
   U19353 : XNOR2_X1 port map( A => n19091, B => n304, ZN => Ciphertext(127));
   U19354 : NOR2_X1 port map( A1 => n19093, A2 => n19911, ZN => n19101);
   U19355 : INV_X1 port map( A => n19094, ZN => n19097);
   U19356 : NAND2_X1 port map( A1 => n19112, A2 => n19095, ZN => n19096);
   U19357 : NAND2_X1 port map( A1 => n19097, A2 => n19096, ZN => n19100);
   U19358 : AND2_X1 port map( A1 => n19115, A2 => n19098, ZN => n19118);
   U19361 : INV_X1 port map( A => n19102, ZN => n19103);
   U19363 : INV_X1 port map( A => n19105, ZN => n19122);
   U19364 : INV_X1 port map( A => n19106, ZN => n19107);
   U19365 : NAND2_X1 port map( A1 => n19107, A2 => n19110, ZN => n19108);
   U19366 : OAI211_X1 port map( C1 => n19111, C2 => n19110, A => n19109, B => 
                           n19108, ZN => n19121);
   U19367 : NOR2_X1 port map( A1 => n19115, A2 => n17203, ZN => n19117);
   U19368 : OAI21_X1 port map( B1 => n19118, B2 => n19117, A => n19116, ZN => 
                           n19119);
   U19369 : OAI211_X1 port map( C1 => n19122, C2 => n19121, A => n19120, B => 
                           n19119, ZN => n19124);
   U19370 : XNOR2_X1 port map( A => n19124, B => n19123, ZN => Ciphertext(130))
                           ;
   U19371 : NOR2_X1 port map( A1 => n19144, A2 => n19134, ZN => n19126);
   U19372 : AOI22_X1 port map( A1 => n19126, A2 => n19125, B1 => n19133, B2 => 
                           n19144, ZN => n19129);
   U19373 : NAND2_X1 port map( A1 => n19127, A2 => n19146, ZN => n19128);
   U19374 : OAI211_X1 port map( C1 => n19130, C2 => n833, A => n19129, B => 
                           n19128, ZN => n19131);
   U19375 : XNOR2_X1 port map( A => n19131, B => n293, ZN => Ciphertext(132));
   U19376 : NAND2_X1 port map( A1 => n19144, A2 => n16780, ZN => n19132);
   U19377 : OAI211_X1 port map( C1 => n19135, C2 => n19144, A => n19133, B => 
                           n19132, ZN => n19139);
   U19378 : NAND3_X1 port map( A1 => n19135, A2 => n19134, A3 => n870, ZN => 
                           n19138);
   U19379 : NAND3_X1 port map( A1 => n19146, A2 => n16780, A3 => n19151, ZN => 
                           n19137);
   U19380 : NAND3_X1 port map( A1 => n19139, A2 => n19138, A3 => n19137, ZN => 
                           n19142);
   U19381 : INV_X1 port map( A => n19140, ZN => n19141);
   U19382 : XNOR2_X1 port map( A => n19142, B => n19141, ZN => Ciphertext(136))
                           ;
   U19383 : AOI21_X1 port map( B1 => n19145, B2 => n19144, A => n870, ZN => 
                           n19150);
   U19384 : OAI21_X1 port map( B1 => n19148, B2 => n19147, A => n19146, ZN => 
                           n19149);
   U19385 : OAI21_X1 port map( B1 => n19151, B2 => n19150, A => n19149, ZN => 
                           n19153);
   U19386 : XNOR2_X1 port map( A => n19153, B => n19152, ZN => Ciphertext(137))
                           ;
   U19387 : INV_X1 port map( A => n19155, ZN => n19161);
   U19388 : AOI21_X1 port map( B1 => n2918, B2 => n19165, A => n19161, ZN => 
                           n19156);
   U19389 : OAI22_X1 port map( A1 => n19157, A2 => n19165, B1 => n19708, B2 => 
                           n19156, ZN => n19160);
   U19390 : INV_X1 port map( A => n19158, ZN => n19159);
   U19391 : XNOR2_X1 port map( A => n19160, B => n19159, ZN => Ciphertext(138))
                           ;
   U19392 : XNOR2_X1 port map( A => n19167, B => n875, ZN => Ciphertext(143));
   U19393 : NAND2_X1 port map( A1 => n19171, A2 => n19170, ZN => n19172);
   U19394 : OAI211_X1 port map( C1 => n19175, C2 => n19174, A => n19173, B => 
                           n19172, ZN => n19177);
   U19395 : INV_X1 port map( A => n2424, ZN => n19176);
   U19396 : XNOR2_X1 port map( A => n19177, B => n19176, ZN => Ciphertext(147))
                           ;
   U19397 : INV_X1 port map( A => n19182, ZN => n19201);
   U19399 : OAI21_X1 port map( B1 => n19197, B2 => n19208, A => n19193, ZN => 
                           n19179);
   U19400 : OAI21_X1 port map( B1 => n19210, B2 => n19189, A => n19209, ZN => 
                           n19178);
   U19401 : AOI22_X1 port map( A1 => n19179, A2 => n19210, B1 => n19197, B2 => 
                           n19178, ZN => n19181);
   U19402 : XNOR2_X1 port map( A => n19181, B => n19180, ZN => Ciphertext(150))
                           ;
   U19403 : AND2_X1 port map( A1 => n19190, A2 => n19208, ZN => n19187);
   U19404 : AOI21_X1 port map( B1 => n19212, B2 => n19193, A => n19187, ZN => 
                           n19185);
   U19405 : NAND2_X1 port map( A1 => n19210, A2 => n19189, ZN => n19183);
   U19408 : XNOR2_X1 port map( A => n19186, B => n1904, ZN => Ciphertext(151));
   U19409 : INV_X1 port map( A => n19187, ZN => n19188);
   U19410 : INV_X1 port map( A => n19196, ZN => n19198);
   U19411 : OAI211_X1 port map( C1 => n19208, C2 => n19201, A => n19188, B => 
                           n19198, ZN => n19192);
   U19412 : NAND3_X1 port map( A1 => n19209, A2 => n19190, A3 => n19189, ZN => 
                           n19191);
   U19413 : OAI211_X1 port map( C1 => n19210, C2 => n19193, A => n19192, B => 
                           n19191, ZN => n19195);
   U19414 : INV_X1 port map( A => n1996, ZN => n19194);
   U19415 : XNOR2_X1 port map( A => n19195, B => n19194, ZN => Ciphertext(153))
                           ;
   U19416 : OAI21_X1 port map( B1 => n19197, B2 => n19209, A => n19842, ZN => 
                           n19215);
   U19417 : AND2_X1 port map( A1 => n19208, A2 => n19209, ZN => n19200);
   U19418 : OAI21_X1 port map( B1 => n19210, B2 => n19201, A => n19198, ZN => 
                           n19199);
   U19419 : OAI21_X1 port map( B1 => n19215, B2 => n19200, A => n19199, ZN => 
                           n19204);
   U19420 : NAND3_X1 port map( A1 => n19202, A2 => n19197, A3 => n19201, ZN => 
                           n19203);
   U19421 : NAND2_X1 port map( A1 => n19204, A2 => n19203, ZN => n19207);
   U19422 : INV_X1 port map( A => n19205, ZN => n19206);
   U19423 : XNOR2_X1 port map( A => n19207, B => n19206, ZN => Ciphertext(154))
                           ;
   U19424 : NOR2_X1 port map( A1 => n2943, A2 => n19209, ZN => n19214);
   U19425 : INV_X1 port map( A => n19210, ZN => n19211);
   U19426 : NAND2_X1 port map( A1 => n19212, A2 => n19211, ZN => n19213);
   U19427 : OAI21_X1 port map( B1 => n19215, B2 => n19214, A => n19213, ZN => 
                           n19218);
   U19428 : INV_X1 port map( A => n19216, ZN => n19217);
   U19429 : XNOR2_X1 port map( A => n19218, B => n19217, ZN => Ciphertext(155))
                           ;
   U19430 : MUX2_X1 port map( A => n19242, B => n19227, S => n19233, Z => 
                           n19221);
   U19431 : AND2_X1 port map( A1 => n19238, A2 => n19234, ZN => n19220);
   U19432 : AOI22_X1 port map( A1 => n19221, A2 => n20124, B1 => n19220, B2 => 
                           n19219, ZN => n19224);
   U19433 : INV_X1 port map( A => n19222, ZN => n19223);
   U19434 : XNOR2_X1 port map( A => n19224, B => n19223, ZN => Ciphertext(158))
                           ;
   U19435 : INV_X1 port map( A => n19225, ZN => n19230);
   U19436 : OAI222_X1 port map( A1 => n19239, A2 => n19230, B1 => n19229, B2 =>
                           n19242, C1 => n19236, C2 => n19228, ZN => n19232);
   U19437 : INV_X1 port map( A => n632, ZN => n19231);
   U19438 : XNOR2_X1 port map( A => n19232, B => n19231, ZN => Ciphertext(159))
                           ;
   U19439 : NAND2_X1 port map( A1 => n19233, A2 => n20124, ZN => n19241);
   U19440 : NAND3_X1 port map( A1 => n19239, A2 => n19238, A3 => n20193, ZN => 
                           n19240);
   U19441 : INV_X1 port map( A => n19243, ZN => n19244);
   U19442 : XNOR2_X1 port map( A => n19245, B => n19244, ZN => Ciphertext(160))
                           ;
   U19443 : NOR2_X1 port map( A1 => n19269, A2 => n19274, ZN => n19268);
   U19444 : INV_X1 port map( A => n19268, ZN => n19258);
   U19445 : INV_X1 port map( A => n19269, ZN => n19275);
   U19446 : INV_X1 port map( A => n19246, ZN => n19267);
   U19447 : NAND3_X1 port map( A1 => n19275, A2 => n19247, A3 => n19267, ZN => 
                           n19257);
   U19448 : INV_X1 port map( A => n19248, ZN => n19253);
   U19449 : INV_X1 port map( A => n19249, ZN => n19250);
   U19450 : OAI211_X1 port map( C1 => n19253, C2 => n20162, A => n19251, B => 
                           n19250, ZN => n19254);
   U19451 : NAND3_X1 port map( A1 => n19278, A2 => n19254, A3 => n19267, ZN => 
                           n19255);
   U19452 : NAND4_X1 port map( A1 => n19258, A2 => n19257, A3 => n19256, A4 => 
                           n19255, ZN => n19260);
   U19453 : XNOR2_X1 port map( A => n19260, B => n19259, ZN => Ciphertext(162))
                           ;
   U19454 : NAND3_X1 port map( A1 => n19261, A2 => n19269, A3 => n2816, ZN => 
                           n19262);
   U19455 : OAI21_X1 port map( B1 => n19279, B2 => n19263, A => n19262, ZN => 
                           n19265);
   U19456 : XNOR2_X1 port map( A => n19265, B => n19264, ZN => Ciphertext(163))
                           ;
   U19457 : NOR2_X1 port map( A1 => n19278, A2 => n19267, ZN => n19266);
   U19458 : INV_X1 port map( A => n2123, ZN => n19273);
   U19459 : OAI22_X1 port map( A1 => n19279, A2 => n19278, B1 => n19277, B2 => 
                           n20444, ZN => n19281);
   U19460 : XNOR2_X1 port map( A => n19281, B => n19280, ZN => Ciphertext(167))
                           ;
   U19461 : OAI21_X1 port map( B1 => n20434, B2 => n19284, A => n19290, ZN => 
                           n19288);
   U19462 : NOR3_X1 port map( A1 => n19298, A2 => n19283, A3 => n19282, ZN => 
                           n19286);
   U19463 : OAI21_X1 port map( B1 => n19298, B2 => n19292, A => n19284, ZN => 
                           n19285);
   U19467 : INV_X1 port map( A => n19290, ZN => n19295);
   U19468 : INV_X1 port map( A => n19299, ZN => n19291);
   U19469 : AOI22_X1 port map( A1 => n1773, A2 => n19292, B1 => n19298, B2 => 
                           n19291, ZN => n19305);
   U19470 : NAND2_X1 port map( A1 => n20510, A2 => n20218, ZN => n19293);
   U19471 : OAI22_X1 port map( A1 => n19305, A2 => n19295, B1 => n19294, B2 => 
                           n19293, ZN => n19297);
   U19472 : XNOR2_X1 port map( A => n19297, B => n19296, ZN => Ciphertext(169))
                           ;
   U19473 : OAI21_X1 port map( B1 => n20364, B2 => n20218, A => n19298, ZN => 
                           n19301);
   U19475 : OAI21_X1 port map( B1 => n19305, B2 => n19304, A => n19303, ZN => 
                           n19307);
   U19476 : INV_X1 port map( A => n456, ZN => n19306);
   U19477 : XNOR2_X1 port map( A => n19307, B => n19306, ZN => Ciphertext(173))
                           ;
   U19478 : OAI21_X1 port map( B1 => n19309, B2 => n19308, A => n19333, ZN => 
                           n19313);
   U19479 : AOI21_X1 port map( B1 => n19311, B2 => n19310, A => n19338, ZN => 
                           n19312);
   U19480 : AOI21_X1 port map( B1 => n19334, B2 => n19313, A => n19312, ZN => 
                           n19314);
   U19481 : XNOR2_X1 port map( A => n19314, B => n2310, ZN => Ciphertext(174));
   U19482 : INV_X1 port map( A => n19315, ZN => n19320);
   U19483 : INV_X1 port map( A => n19316, ZN => n19317);
   U19484 : NAND3_X1 port map( A1 => n19317, A2 => n19324, A3 => n19749, ZN => 
                           n19319);
   U19485 : INV_X1 port map( A => n19333, ZN => n19327);
   U19486 : NAND3_X1 port map( A1 => n19327, A2 => n19308, A3 => n19329, ZN => 
                           n19318);
   U19488 : INV_X1 port map( A => n19321, ZN => n19322);
   U19490 : NOR2_X1 port map( A1 => n19333, A2 => n19324, ZN => n19326);
   U19491 : OAI21_X1 port map( B1 => n19326, B2 => n19340, A => n19336, ZN => 
                           n19325);
   U19492 : OAI211_X1 port map( C1 => n19336, C2 => n19326, A => n19325, B => 
                           n19955, ZN => n19346);
   U19493 : OAI21_X1 port map( B1 => n19334, B2 => n19336, A => n19327, ZN => 
                           n19332);
   U19494 : NAND2_X1 port map( A1 => n19749, A2 => n19336, ZN => n19331);
   U19495 : NAND3_X1 port map( A1 => n19333, A2 => n19329, A3 => n19337, ZN => 
                           n19330);
   U19496 : NAND4_X1 port map( A1 => n19340, A2 => n19332, A3 => n19331, A4 => 
                           n19330, ZN => n19345);
   U19497 : NOR2_X1 port map( A1 => n19333, A2 => n19955, ZN => n19335);
   U19498 : NAND4_X1 port map( A1 => n19340, A2 => n19336, A3 => n19335, A4 => 
                           n19334, ZN => n19344);
   U19499 : XNOR2_X1 port map( A => n19338, B => n19337, ZN => n19342);
   U19500 : NOR2_X1 port map( A1 => n19340, A2 => n19955, ZN => n19341);
   U19501 : NAND2_X1 port map( A1 => n19342, A2 => n19341, ZN => n19343);
   U19502 : NAND4_X1 port map( A1 => n19346, A2 => n19345, A3 => n19344, A4 => 
                           n19343, ZN => Ciphertext(178));
   U19503 : AND2_X1 port map( A1 => n20240, A2 => n19349, ZN => n19359);
   U19504 : OAI21_X1 port map( B1 => n20244, B2 => n19348, A => n19347, ZN => 
                           n19358);
   U19505 : NAND2_X1 port map( A1 => n19351, A2 => n20273, ZN => n19356);
   U19506 : NAND2_X1 port map( A1 => n19353, A2 => n19352, ZN => n19355);
   U19507 : MUX2_X1 port map( A => n19356, B => n19355, S => n20240, Z => 
                           n19357);
   U19508 : OAI21_X1 port map( B1 => n19359, B2 => n19358, A => n19357, ZN => 
                           n19444);
   U19509 : INV_X1 port map( A => n19444, ZN => n19409);
   U19510 : NOR2_X1 port map( A1 => n19361, A2 => n19360, ZN => n19369);
   U19511 : INV_X1 port map( A => n20212, ZN => n19364);
   U19512 : NAND2_X1 port map( A1 => n19364, A2 => n19938, ZN => n19368);
   U19513 : NAND2_X1 port map( A1 => n19366, A2 => n19365, ZN => n19367);
   U19514 : OAI21_X1 port map( B1 => n19369, B2 => n19368, A => n19367, ZN => 
                           n19440);
   U19515 : INV_X1 port map( A => n19440, ZN => n19381);
   U19516 : MUX2_X1 port map( A => n19373, B => n19666, S => n19370, Z => 
                           n19379);
   U19517 : NAND2_X1 port map( A1 => n19373, A2 => n19372, ZN => n19377);
   U19521 : OAI21_X1 port map( B1 => n1897, B2 => n20463, A => n19382, ZN => 
                           n19384);
   U19522 : NOR2_X1 port map( A1 => n19388, A2 => n20004, ZN => n19393);
   U19523 : NOR2_X1 port map( A1 => n19390, A2 => n20172, ZN => n19392);
   U19524 : OAI21_X1 port map( B1 => n19393, B2 => n19392, A => n19391, ZN => 
                           n19398);
   U19525 : NAND3_X1 port map( A1 => n19396, A2 => n19395, A3 => n20004, ZN => 
                           n19397);
   U19526 : NAND2_X1 port map( A1 => n3827, A2 => n19425, ZN => n19408);
   U19527 : OAI21_X1 port map( B1 => n19402, B2 => n19403, A => n19401, ZN => 
                           n19406);
   U19529 : OAI21_X1 port map( B1 => n19409, B2 => n19442, A => n19418, ZN => 
                           n19407);
   U19530 : AOI22_X1 port map( A1 => n19409, A2 => n19408, B1 => n19407, B2 => 
                           n19439, ZN => n19411);
   U19531 : XNOR2_X1 port map( A => n19411, B => n19410, ZN => Ciphertext(180))
                           ;
   U19532 : INV_X1 port map( A => n19442, ZN => n19434);
   U19533 : NOR2_X1 port map( A1 => n19439, A2 => n19440, ZN => n19430);
   U19534 : OAI21_X1 port map( B1 => n19444, B2 => n19434, A => n19430, ZN => 
                           n19413);
   U19535 : AND2_X1 port map( A1 => n19440, A2 => n19432, ZN => n19445);
   U19536 : OAI21_X1 port map( B1 => n19445, B2 => n19434, A => n19425, ZN => 
                           n19412);
   U19537 : NAND2_X1 port map( A1 => n19413, A2 => n19412, ZN => n19415);
   U19538 : INV_X1 port map( A => n2298, ZN => n19414);
   U19539 : XNOR2_X1 port map( A => n19415, B => n19414, ZN => Ciphertext(181))
                           ;
   U19540 : MUX2_X1 port map( A => n19444, B => n19439, S => n19441, Z => 
                           n19416);
   U19541 : NAND2_X1 port map( A1 => n19416, A2 => n19442, ZN => n19421);
   U19546 : XNOR2_X1 port map( A => n19423, B => n19422, ZN => Ciphertext(182))
                           ;
   U19547 : NAND2_X1 port map( A1 => n19442, A2 => n19440, ZN => n19424);
   U19548 : NAND2_X1 port map( A1 => n19424, A2 => n19448, ZN => n19429);
   U19549 : INV_X1 port map( A => n19439, ZN => n19426);
   U19550 : NAND3_X1 port map( A1 => n19426, A2 => n19442, A3 => n19418, ZN => 
                           n19427);
   U19551 : OAI211_X1 port map( C1 => n19430, C2 => n19429, A => n19428, B => 
                           n19427, ZN => n19431);
   U19552 : XNOR2_X1 port map( A => n19431, B => n2709, ZN => Ciphertext(183));
   U19553 : MUX2_X1 port map( A => n19440, B => n19439, S => n19432, Z => 
                           n19435);
   U19554 : NAND2_X1 port map( A1 => n19439, A2 => n19432, ZN => n19433);
   U19555 : INV_X1 port map( A => n19436, ZN => n19437);
   U19556 : XNOR2_X1 port map( A => n19438, B => n19437, ZN => Ciphertext(184))
                           ;
   U19557 : AOI21_X1 port map( B1 => n19440, B2 => n19439, A => n19418, ZN => 
                           n19449);
   U19558 : INV_X1 port map( A => n19441, ZN => n19443);
   U19559 : NOR2_X1 port map( A1 => n19443, A2 => n19442, ZN => n19446);
   U19560 : OAI21_X1 port map( B1 => n19446, B2 => n19445, A => n19444, ZN => 
                           n19447);
   U19561 : OAI21_X1 port map( B1 => n19449, B2 => n19448, A => n19447, ZN => 
                           n19451);
   U19562 : INV_X1 port map( A => n620, ZN => n19450);
   U19563 : XNOR2_X1 port map( A => n19451, B => n19450, ZN => Ciphertext(185))
                           ;
   U19564 : OAI22_X1 port map( A1 => n212, A2 => n19453, B1 => n19463, B2 => 
                           n19460, ZN => n19466);
   U19565 : NAND2_X1 port map( A1 => n19453, A2 => n19459, ZN => n19454);
   U19566 : AOI22_X1 port map( A1 => n19466, A2 => n19456, B1 => n19738, B2 => 
                           n19454, ZN => n19458);
   U19567 : XNOR2_X1 port map( A => n19458, B => n19457, ZN => Ciphertext(187))
                           ;
   U19568 : INV_X1 port map( A => n19459, ZN => n19465);
   U19569 : INV_X1 port map( A => n19460, ZN => n19461);
   U19570 : OAI21_X1 port map( B1 => n19463, B2 => n19462, A => n19461, ZN => 
                           n19464);
   U19571 : AOI22_X1 port map( A1 => n19466, A2 => n19465, B1 => n19464, B2 => 
                           n212, ZN => n19468);
   U19572 : XNOR2_X1 port map( A => n19468, B => n19467, ZN => Ciphertext(191))
                           ;
   U8160 : NAND3_X2 port map( A1 => n3556, A2 => n3553, A3 => n3552, ZN => 
                           n9635);
   U1007 : NOR2_X2 port map( A1 => n8164, A2 => n8163, ZN => n9070);
   U1001 : MUX2_X2 port map( A => n11878, B => n11877, S => n12577, Z => n13848
                           );
   U4182 : XNOR2_X2 port map( A => n5166, B => n5165, ZN => n2792);
   U281 : INV_X1 port map( A => n15479, ZN => n17909);
   U68 : MUX2_X2 port map( A => n4195, B => n4194, S => n4370, Z => n5424);
   U257 : NOR2_X2 port map( A1 => n11542, A2 => n11543, ZN => n12029);
   U1842 : OR2_X2 port map( A1 => n2876, A2 => n2880, ZN => n7202);
   U851 : NOR2_X1 port map( A1 => n12223, A2 => n10925, ZN => n12121);
   U1550 : AOI21_X1 port map( B1 => n9619, B2 => n9618, A => n9617, ZN => 
                           n11830);
   U1449 : BUF_X2 port map( A => n14626, Z => n954);
   U1116 : BUF_X1 port map( A => n5762, Z => n8205);
   U8440 : BUF_X2 port map( A => n16673, Z => n19349);
   U1649 : BUF_X1 port map( A => n11389, Z => n11870);
   U739 : INV_X1 port map( A => n9391, ZN => n10594);
   U1763 : OR2_X2 port map( A1 => n427, A2 => n3625, ZN => n9029);
   U79 : NAND2_X1 port map( A1 => n615, A2 => n446, ZN => n6782);
   U10038 : NAND3_X2 port map( A1 => n5549, A2 => n5547, A3 => n5548, ZN => 
                           n7155);
   U2021 : CLKBUF_X1 port map( A => Key(117), Z => n19102);
   U981 : XNOR2_X1 port map( A => Key(155), B => Plaintext(155), ZN => n4567);
   U2030 : XNOR2_X1 port map( A => Plaintext(136), B => Key(136), ZN => n4271);
   U2014 : CLKBUF_X1 port map( A => Key(6), Z => n18691);
   U512 : XNOR2_X1 port map( A => Key(30), B => Plaintext(30), ZN => n4911);
   U436 : XNOR2_X1 port map( A => Key(26), B => Plaintext(26), ZN => n4945);
   U1981 : XNOR2_X1 port map( A => Key(25), B => Plaintext(25), ZN => n4940);
   U8874 : BUF_X1 port map( A => n4518, Z => n4523);
   U539 : XNOR2_X1 port map( A => n3857, B => Key(90), ZN => n5095);
   U9103 : AND2_X1 port map( A1 => n4940, A2 => n4118, ZN => n4886);
   U955 : XNOR2_X1 port map( A => n3971, B => Key(40), ZN => n4962);
   U154 : XNOR2_X1 port map( A => n3844, B => Key(82), ZN => n5115);
   U3464 : BUF_X1 port map( A => n4152, Z => n4546);
   U121 : OAI211_X1 port map( C1 => n4290, C2 => n4018, A => n4017, B => n4627,
                           ZN => n5322);
   U1946 : OR2_X1 port map( A1 => n4041, A2 => n4769, ZN => n5034);
   U1914 : OR2_X1 port map( A1 => n3886, A2 => n3885, ZN => n1776);
   U5819 : AND2_X1 port map( A1 => n3550, A2 => n3549, ZN => n1807);
   U416 : AND2_X1 port map( A1 => n4086, A2 => n4085, ZN => n6000);
   U546 : NAND2_X1 port map( A1 => n643, A2 => n664, ZN => n5803);
   U557 : MUX2_X1 port map( A => n3955, B => n3954, S => n4609, Z => n5573);
   U8512 : INV_X1 port map( A => n5148, ZN => n5582);
   U244 : NAND2_X1 port map( A1 => n1985, A2 => n4292, ZN => n5628);
   U466 : INV_X1 port map( A => n5264, ZN => n6143);
   U510 : NAND2_X1 port map( A1 => n3262, A2 => n5522, ZN => n5973);
   U630 : OR2_X1 port map( A1 => n4183, A2 => n4184, ZN => n6708);
   U420 : INV_X1 port map( A => n7188, ZN => n6427);
   U5974 : OAI21_X1 port map( B1 => n5566, B2 => n1895, A => n1894, ZN => n7382
                           );
   U6480 : OR2_X1 port map( A1 => n5131, A2 => n5130, ZN => n7144);
   U745 : OAI21_X1 port map( B1 => n6063, B2 => n6064, A => n6062, ZN => n7017)
                           ;
   U10555 : XNOR2_X1 port map( A => n6477, B => n7253, ZN => n6660);
   U1831 : NAND3_X1 port map( A1 => n2396, A2 => n2099, A3 => n2098, ZN => 
                           n7151);
   U818 : XNOR2_X1 port map( A => n7322, B => n7321, ZN => n8325);
   U11019 : XNOR2_X1 port map( A => n6930, B => n6929, ZN => n8165);
   U864 : XNOR2_X1 port map( A => n6006, B => n6005, ZN => n8197);
   U10975 : XNOR2_X1 port map( A => n6870, B => n6869, ZN => n8352);
   U349 : BUF_X1 port map( A => n7877, Z => n8044);
   U10917 : OAI211_X1 port map( C1 => n8385, C2 => n6800, A => n6799, B => 
                           n7685, ZN => n9310);
   U11588 : OAI21_X1 port map( B1 => n7694, B2 => n7693, A => n7692, ZN => 
                           n8904);
   U10816 : OR2_X1 port map( A1 => n6654, A2 => n6653, ZN => n9189);
   U282 : NAND4_X2 port map( A1 => n3719, A2 => n5299, A3 => n3718, A4 => n5298
                           , ZN => n1037);
   U1112 : NAND3_X1 port map( A1 => n3311, A2 => n8255, A3 => n769, ZN => n9130
                           );
   U3832 : INV_X1 port map( A => n8797, ZN => n9112);
   U1710 : INV_X1 port map( A => n670, ZN => n9256);
   U1713 : OR2_X1 port map( A1 => n8611, A2 => n7537, ZN => n8698);
   U3524 : OR3_X1 port map( A1 => n8649, A2 => n8991, A3 => n20265, ZN => n2887
                           );
   U6214 : NAND3_X1 port map( A1 => n2015, A2 => n8629, A3 => n2014, ZN => 
                           n10582);
   U870 : OAI211_X1 port map( C1 => n2651, C2 => n2650, A => n8412, B => n2652,
                           ZN => n10425);
   U1673 : INV_X1 port map( A => n10237, ZN => n9994);
   U2595 : XNOR2_X1 port map( A => n20156, B => n10046, ZN => n10347);
   U849 : XNOR2_X1 port map( A => n9522, B => n9521, ZN => n10960);
   U12608 : XNOR2_X1 port map( A => n9474, B => n9473, ZN => n11148);
   U8115 : XNOR2_X1 port map( A => n9907, B => n9906, ZN => n3507);
   U814 : BUF_X1 port map( A => n11087, Z => n11454);
   U615 : NAND3_X1 port map( A1 => n576, A2 => n9199, A3 => n9200, ZN => n12354
                           );
   U604 : NAND2_X1 port map( A1 => n11288, A2 => n19972, ZN => n12811);
   U2177 : NAND2_X1 port map( A1 => n3489, A2 => n10949, ZN => n12126);
   U2087 : NAND3_X1 port map( A1 => n9485, A2 => n3381, A3 => n2045, ZN => 
                           n12180);
   U14040 : OAI21_X1 port map( B1 => n11434, B2 => n11433, A => n11432, ZN => 
                           n12167);
   U7470 : OAI211_X1 port map( C1 => n11250, C2 => n11383, A => n11249, B => 
                           n11384, ZN => n12372);
   U1547 : NAND3_X1 port map( A1 => n1278, A2 => n766, A3 => n765, ZN => n11942
                           );
   U415 : OR2_X1 port map( A1 => n11995, A2 => n11997, ZN => n12322);
   U115 : OR2_X1 port map( A1 => n12534, A2 => n12532, ZN => n12293);
   U3010 : OR2_X1 port map( A1 => n12492, A2 => n253, ZN => n12813);
   U14580 : NOR2_X1 port map( A1 => n12327, A2 => n12514, ZN => n13269);
   U2716 : AND3_X1 port map( A1 => n1828, A2 => n1827, A3 => n609, ZN => n13427
                           );
   U609 : NAND3_X1 port map( A1 => n2148, A2 => n12144, A3 => n2147, ZN => 
                           n13644);
   U135 : XNOR2_X1 port map( A => n12626, B => n12625, ZN => n14791);
   U904 : XNOR2_X1 port map( A => n13548, B => n13547, ZN => n14482);
   U7204 : XNOR2_X1 port map( A => n2624, B => n2623, ZN => n14236);
   U189 : XNOR2_X1 port map( A => n13516, B => n13515, ZN => n14487);
   U338 : XNOR2_X1 port map( A => n1973, B => n13349, ZN => n14693);
   U15104 : XNOR2_X1 port map( A => n13024, B => n13023, ZN => n14506);
   U611 : OR2_X1 port map( A1 => n14693, A2 => n200, ZN => n14696);
   U15972 : NAND4_X1 port map( A1 => n14253, A2 => n14254, A3 => n14255, A4 => 
                           n14252, ZN => n15531);
   U927 : AOI21_X1 port map( B1 => n14301, B2 => n14508, A => n14300, ZN => 
                           n14902);
   U471 : OAI21_X1 port map( B1 => n13671, B2 => n14247, A => n14246, ZN => 
                           n15921);
   U6095 : NOR2_X1 port map( A1 => n15458, A2 => n20173, ZN => n15239);
   U16897 : NOR2_X1 port map( A1 => n230, A2 => n868, ZN => n15851);
   U4890 : AND2_X1 port map( A1 => n1217, A2 => n1220, ZN => n17328);
   U4152 : AND4_X1 port map( A1 => n15668, A2 => n1018, A3 => n15669, A4 => 
                           n15670, ZN => n955);
   U6147 : XNOR2_X1 port map( A => n16958, B => n16957, ZN => n17812);
   U6801 : XNOR2_X1 port map( A => n16218, B => n16217, ZN => n17489);
   U111 : XNOR2_X1 port map( A => n14634, B => n14633, ZN => n17508);
   U834 : BUF_X1 port map( A => n18092, Z => n160);
   U317 : BUF_X1 port map( A => n16263, Z => n17079);
   U140 : XNOR2_X1 port map( A => n16235, B => n16234, ZN => n17492);
   U116 : CLKBUF_X1 port map( A => n16805, Z => n17959);
   U3674 : AOI21_X1 port map( B1 => n2335, B2 => n17510, A => n16634, ZN => 
                           n18342);
   U18029 : AOI22_X1 port map( A1 => n17086, A2 => n17602, B1 => n17085, B2 => 
                           n17601, ZN => n18306);
   U18017 : AND3_X1 port map( A1 => n17073, A2 => n17072, A3 => n17071, ZN => 
                           n19162);
   U6415 : NOR2_X1 port map( A1 => n16815, A2 => n16814, ZN => n18529);
   U17153 : OR2_X1 port map( A1 => n16114, A2 => n16113, ZN => n19170);
   U81 : AOI21_X1 port map( B1 => n17230, B2 => n17510, A => n17229, ZN => 
                           n18392);
   U283 : XNOR2_X1 port map( A => Key(61), B => Plaintext(61), ZN => n4651);
   U567 : CLKBUF_X1 port map( A => Key(186), Z => n106);
   U1199 : CLKBUF_X1 port map( A => Key(156), Z => n2306);
   U2368 : XNOR2_X1 port map( A => n3908, B => Key(156), ZN => n4571);
   U6122 : INV_X1 port map( A => n5107, ZN => n3259);
   U5154 : XNOR2_X1 port map( A => n6797, B => n6798, ZN => n8386);
   U9776 : INV_X1 port map( A => n8301, ZN => n8046);
   U6706 : NAND2_X1 port map( A1 => n7871, A2 => n7615, ZN => n7618);
   U6895 : AND2_X1 port map( A1 => n7888, A2 => n7887, ZN => n9275);
   U13968 : INV_X1 port map( A => n12021, ZN => n12369);
   U1003 : NAND2_X1 port map( A1 => n11809, A2 => n11810, ZN => n12212);
   U10 : AOI21_X2 port map( B1 => n14259, B2 => n15421, A => n14258, ZN => 
                           n16836);
   U16959 : XNOR2_X2 port map( A => n15942, B => n15941, ZN => n17823);
   U4245 : BUF_X2 port map( A => n14000, Z => n14620);
   U826 : XNOR2_X2 port map( A => n4035, B => Key(132), ZN => n4095);
   U907 : NAND2_X2 port map( A1 => n597, A2 => n599, ZN => n10349);
   U1872 : NAND4_X2 port map( A1 => n5609, A2 => n5607, A3 => n5608, A4 => 
                           n5606, ZN => n6558);
   U1684 : AND4_X2 port map( A1 => n8788, A2 => n8787, A3 => n3466, A4 => n3465
                           , ZN => n9771);
   U2350 : NAND2_X2 port map( A1 => n445, A2 => n1483, ZN => n7333);
   U117 : AND3_X2 port map( A1 => n344, A2 => n11369, A3 => n11368, ZN => 
                           n12312);
   U7799 : NAND3_X2 port map( A1 => n3191, A2 => n4672, A3 => n3192, ZN => 
                           n6171);
   U6207 : MUX2_X2 port map( A => n8406, B => n8405, S => n9164, Z => n9794);
   U1679 : MUX2_X2 port map( A => n7806, B => n7805, S => n2243, Z => n10262);
   U1743 : AND2_X2 port map( A1 => n2259, A2 => n2258, ZN => n9159);
   U184 : AND2_X2 port map( A1 => n7698, A2 => n7697, ZN => n8720);
   U771 : OAI21_X2 port map( B1 => n4751, B2 => n4750, A => n4749, ZN => n5172)
                           ;
   U1650 : BUF_X2 port map( A => n9492, Z => n10649);
   U253 : AND2_X2 port map( A1 => n9497, A2 => n9496, ZN => n11673);
   U7979 : NOR2_X2 port map( A1 => n14786, A2 => n14785, ZN => n15582);
   U2865 : OAI211_X2 port map( C1 => n2888, C2 => n9278, A => n2887, B => n702,
                           ZN => n10185);
   U1492 : AND3_X2 port map( A1 => n3531, A2 => n1641, A3 => n1020, ZN => 
                           n12713);
   U580 : NOR2_X2 port map( A1 => n9047, A2 => n9048, ZN => n9289);
   U14 : BUF_X2 port map( A => n12658, Z => n15766);
   U702 : OAI211_X2 port map( C1 => n15264, C2 => n15265, A => n15263, B => 
                           n15262, ZN => n16987);
   U8469 : OR3_X1 port map( A1 => n14599, A2 => n14603, A3 => n19918, ZN => 
                           n3815);
   U3 : AND3_X1 port map( A1 => n17065, A2 => n17718, A3 => n17064, ZN => 
                           n19163);
   U4 : AOI211_X1 port map( C1 => n14449, C2 => n14453, A => n13927, B => 
                           n14452, ZN => n12929);
   U7 : XNOR2_X1 port map( A => n10184, B => n10183, ZN => n19830);
   U120 : NOR2_X2 port map( A1 => n11811, A2 => n11638, ZN => n12207);
   U137 : OAI211_X2 port map( C1 => n7682, C2 => n8166, A => n7681, B => n7680,
                           ZN => n19941);
   U151 : OAI22_X1 port map( A1 => n14342, A2 => n13931, B1 => n14335, B2 => 
                           n12879, ZN => n14050);
   U153 : NOR2_X1 port map( A1 => n18741, A2 => n18775, ZN => n18746);
   U155 : INV_X1 port map( A => n16665, ZN => n1897);
   U187 : INV_X1 port map( A => n2684, ZN => n3223);
   U198 : XOR2_X1 port map( A => n17422, B => n17421, Z => n19472);
   U201 : BUF_X2 port map( A => n14325, Z => n14352);
   U226 : XNOR2_X1 port map( A => n6210, B => n3805, ZN => n8195);
   U245 : BUF_X1 port map( A => n6381, Z => n19476);
   U252 : AOI21_X1 port map( B1 => n4718, B2 => n4717, A => n4716, ZN => n6381)
                           ;
   U264 : XNOR2_X2 port map( A => n12853, B => n12852, ZN => n14449);
   U293 : BUF_X1 port map( A => n16921, Z => n19860);
   U325 : AND3_X2 port map( A1 => n3324, A2 => n3325, A3 => n3566, ZN => n12506
                           );
   U363 : XNOR2_X1 port map( A => n9511, B => n9510, ZN => n11144);
   U365 : NOR2_X2 port map( A1 => n3677, A2 => n7467, ZN => n8550);
   U381 : AND3_X2 port map( A1 => n11916, A2 => n3161, A3 => n3160, ZN => 
                           n12470);
   U422 : XNOR2_X2 port map( A => n10308, B => n10307, ZN => n11255);
   U484 : XNOR2_X1 port map( A => n12779, B => n12778, ZN => n12800);
   U507 : XNOR2_X2 port map( A => Key(98), B => Plaintext(98), ZN => n5075);
   U520 : NAND2_X2 port map( A1 => n3622, A2 => n393, ZN => n5668);
   U533 : XNOR2_X2 port map( A => Key(51), B => Plaintext(51), ZN => n4856);
   U579 : XNOR2_X2 port map( A => n3923, B => Key(170), ZN => n4343);
   U623 : OAI211_X2 port map( C1 => n705, C2 => n708, A => n706, B => n704, ZN 
                           => n10506);
   U625 : XNOR2_X2 port map( A => n11936, B => n11935, ZN => n19875);
   U652 : AND3_X2 port map( A1 => n1673, A2 => n1710, A3 => n1711, ZN => n11586
                           );
   U665 : OAI211_X1 port map( C1 => n7840, C2 => n8910, A => n7839, B => n7838,
                           ZN => n9009);
   U674 : BUF_X2 port map( A => n16321, Z => n18539);
   U675 : XNOR2_X2 port map( A => n3921, B => Key(169), ZN => n4517);
   U685 : CLKBUF_X1 port map( A => n10575, Z => n11499);
   U716 : XNOR2_X2 port map( A => Key(111), B => Plaintext(111), ZN => n5087);
   U724 : INV_X1 port map( A => n5095, ZN => n4788);
   U751 : XNOR2_X2 port map( A => Key(152), B => Plaintext(152), ZN => n4752);
   U754 : NAND2_X2 port map( A1 => n5157, A2 => n499, ZN => n7364);
   U822 : XNOR2_X2 port map( A => n10479, B => n10478, ZN => n11034);
   U839 : XNOR2_X2 port map( A => n1285, B => n9599, ZN => n11292);
   U847 : OAI211_X2 port map( C1 => n2846, C2 => n11160, A => n2842, B => 
                           n19570, ZN => n1508);
   U862 : XNOR2_X2 port map( A => Key(146), B => Plaintext(146), ZN => n4744);
   U871 : OAI211_X2 port map( C1 => n5831, C2 => n6018, A => n5830, B => n5829,
                           ZN => n7154);
   U876 : OAI21_X2 port map( B1 => n11268, B2 => n11336, A => n602, ZN => 
                           n12374);
   U893 : XNOR2_X1 port map( A => n12743, B => n12744, ZN => n14347);
   U906 : XNOR2_X2 port map( A => n3153, B => Key(143), ZN => n4555);
   U919 : OAI21_X2 port map( B1 => n15151, B2 => n15150, A => n15149, ZN => 
                           n16900);
   U920 : XNOR2_X2 port map( A => n4028, B => Key(114), ZN => n4697);
   U944 : INV_X1 port map( A => n18376, ZN => n19501);
   U949 : NAND2_X1 port map( A1 => n1844, A2 => n16255, ZN => n18495);
   U953 : NOR2_X1 port map( A1 => n16658, A2 => n17208, ZN => n17217);
   U958 : OR2_X1 port map( A1 => n15400, A2 => n15892, ZN => n14285);
   U961 : INV_X1 port map( A => n14700, ZN => n19503);
   U969 : INV_X1 port map( A => n12372, ZN => n19504);
   U976 : INV_X1 port map( A => n4970, ZN => n19507);
   U1011 : OR2_X1 port map( A1 => n16249, A2 => n16248, ZN => n19729);
   U1013 : NOR2_X1 port map( A1 => n20214, A2 => n19098, ZN => n19113);
   U1016 : NOR2_X1 port map( A1 => n18781, A2 => n18741, ZN => n19551);
   U1026 : AND4_X1 port map( A1 => n3548, A2 => n3544, A3 => n3545, A4 => n3547
                           , ZN => n19681);
   U1037 : NOR2_X2 port map( A1 => n16441, A2 => n16440, ZN => n19775);
   U1053 : AND3_X1 port map( A1 => n17073, A2 => n17072, A3 => n17071, ZN => 
                           n19708);
   U1059 : NOR2_X1 port map( A1 => n18136, A2 => n18135, ZN => n19745);
   U1073 : INV_X1 port map( A => n18673, ZN => n19510);
   U1088 : INV_X1 port map( A => n19390, ZN => n19511);
   U1128 : XNOR2_X1 port map( A => n16204, B => n16203, ZN => n18534);
   U1268 : XNOR2_X1 port map( A => n17377, B => n19640, ZN => n16119);
   U1282 : INV_X1 port map( A => n15852, ZN => n17433);
   U1302 : MUX2_X1 port map( A => n12936, B => n12935, S => n15380, Z => n17104
                           );
   U1310 : CLKBUF_X1 port map( A => n15502, Z => n19813);
   U1325 : NAND2_X1 port map( A1 => n19537, A2 => n14368, ZN => n15905);
   U1328 : INV_X1 port map( A => n15502, ZN => n19512);
   U1330 : OAI21_X1 port map( B1 => n14365, B2 => n14364, A => n19538, ZN => 
                           n19537);
   U1346 : INV_X1 port map( A => n15709, ZN => n19514);
   U1349 : OR2_X1 port map( A1 => n2314, A2 => n14599, ZN => n13855);
   U1352 : OR2_X1 port map( A1 => n20513, A2 => n14599, ZN => n14600);
   U1380 : AND2_X1 port map( A1 => n11473, A2 => n11472, ZN => n924);
   U1396 : OR2_X1 port map( A1 => n8402, A2 => n8401, ZN => n19769);
   U1402 : XNOR2_X1 port map( A => n10014, B => n10015, ZN => n11573);
   U1424 : OAI21_X1 port map( B1 => n9564, B2 => n19590, A => n2169, ZN => 
                           n8415);
   U1453 : AND2_X1 port map( A1 => n9249, A2 => n8974, ZN => n3356);
   U1454 : AND2_X1 port map( A1 => n477, A2 => n19550, ZN => n8499);
   U1474 : AND2_X1 port map( A1 => n8602, A2 => n8743, ZN => n8483);
   U1486 : INV_X1 port map( A => n9106, ZN => n19515);
   U1498 : INV_X1 port map( A => n8974, ZN => n19516);
   U1500 : OR2_X1 port map( A1 => n5965, A2 => n19579, ZN => n19577);
   U1502 : INV_X1 port map( A => n8772, ZN => n19517);
   U1508 : BUF_X2 port map( A => n8735, Z => n19518);
   U1517 : INV_X1 port map( A => n8828, ZN => n19519);
   U1618 : INV_X1 port map( A => n8384, ZN => n19589);
   U1621 : INV_X1 port map( A => n7500, ZN => n19651);
   U1626 : INV_X1 port map( A => n8316, ZN => n19520);
   U1629 : INV_X1 port map( A => n7903, ZN => n19521);
   U1641 : INV_X1 port map( A => n5410, ZN => n5681);
   U1645 : INV_X1 port map( A => n5704, ZN => n5996);
   U1652 : INV_X1 port map( A => n5382, ZN => n6194);
   U1663 : INV_X1 port map( A => n6206, ZN => n19522);
   U1746 : AND2_X1 port map( A1 => n4609, A2 => n4177, ZN => n19963);
   U1754 : XNOR2_X1 port map( A => n3870, B => Key(34), ZN => n4952);
   U1755 : OR2_X1 port map( A1 => n4319, A2 => n4324, ZN => n4146);
   U1765 : INV_X1 port map( A => n4651, ZN => n19523);
   U1766 : XNOR2_X1 port map( A => Key(135), B => Plaintext(135), ZN => n19788)
                           ;
   U1768 : AND2_X1 port map( A1 => n4467, A2 => n4887, ZN => n4889);
   U1803 : BUF_X1 port map( A => n4041, Z => n5032);
   U1832 : OR2_X1 port map( A1 => n4204, A2 => n5010, ZN => n19540);
   U1848 : CLKBUF_X1 port map( A => n4094, Z => n5029);
   U1851 : XNOR2_X1 port map( A => Key(168), B => Plaintext(168), ZN => n4187);
   U1852 : AND2_X1 port map( A1 => n6050, A2 => n3351, ZN => n3665);
   U1855 : OR2_X1 port map( A1 => n3959, A2 => n5405, ZN => n5316);
   U1887 : OR2_X1 port map( A1 => n5291, A2 => n5645, ZN => n2321);
   U1939 : INV_X1 port map( A => n3351, ZN => n6052);
   U1958 : OR2_X1 port map( A1 => n5158, A2 => n5429, ZN => n499);
   U2029 : XNOR2_X1 port map( A => n7230, B => n7151, ZN => n6495);
   U2048 : XNOR2_X1 port map( A => n7304, B => n6348, ZN => n6961);
   U2051 : XNOR2_X1 port map( A => n6789, B => n6788, ZN => n8132);
   U2088 : OR2_X1 port map( A1 => n7932, A2 => n7931, ZN => n1453);
   U2107 : OR2_X1 port map( A1 => n7648, A2 => n8079, ZN => n19622);
   U2108 : OR2_X1 port map( A1 => n9242, A2 => n9189, ZN => n431);
   U2109 : AND2_X1 port map( A1 => n8304, A2 => n2792, ZN => n1244);
   U2116 : CLKBUF_X1 port map( A => n8221, Z => n19809);
   U2135 : AOI21_X1 port map( B1 => n8382, B2 => n8381, A => n19589, ZN => 
                           n8391);
   U2150 : OAI211_X1 port map( C1 => n7902, C2 => n7909, A => n19582, B => 
                           n7754, ZN => n2251);
   U2156 : INV_X1 port map( A => n803, ZN => n9211);
   U2231 : NOR3_X1 port map( A1 => n9130, A2 => n9129, A3 => n9201, ZN => n9131
                           );
   U2232 : XNOR2_X1 port map( A => n9391, B => n9392, ZN => n10454);
   U2235 : NAND2_X1 port map( A1 => n1398, A2 => n8425, ZN => n694);
   U2267 : AND2_X1 port map( A1 => n19878, A2 => n11174, ZN => n19614);
   U2282 : CLKBUF_X1 port map( A => n11884, Z => n909);
   U2283 : OR2_X1 port map( A1 => n10945, A2 => n1654, ZN => n19571);
   U2317 : AOI22_X1 port map( A1 => n10828, A2 => n10827, B1 => n10826, B2 => 
                           n11041, ZN => n12202);
   U2334 : OR2_X1 port map( A1 => n12380, A2 => n12381, ZN => n19592);
   U2344 : AOI21_X1 port map( B1 => n10452, B2 => n10451, A => n2656, ZN => 
                           n10471);
   U2362 : BUF_X1 port map( A => n11769, Z => n12528);
   U2388 : OAI21_X1 port map( B1 => n11684, B2 => n11685, A => n19585, ZN => 
                           n19584);
   U2421 : INV_X1 port map( A => n2220, ZN => n19535);
   U2424 : XNOR2_X1 port map( A => n13539, B => n13716, ZN => n13771);
   U2425 : XNOR2_X1 port map( A => n13312, B => n13791, ZN => n13483);
   U2432 : INV_X1 port map( A => n2684, ZN => n19598);
   U2438 : BUF_X1 port map( A => n14490, Z => n14753);
   U2439 : INV_X1 port map( A => n14369, ZN => n19538);
   U2440 : CLKBUF_X1 port map( A => n14779, Z => n877);
   U2446 : XOR2_X1 port map( A => n13334, B => n13333, Z => n19895);
   U2452 : INV_X1 port map( A => n19634, ZN => n19600);
   U2488 : AND2_X1 port map( A1 => n3431, A2 => n15606, ZN => n19542);
   U2514 : NAND2_X1 port map( A1 => n13978, A2 => n2353, ZN => n15874);
   U2515 : AND2_X1 port map( A1 => n2288, A2 => n15503, ZN => n3019);
   U2519 : OR2_X1 port map( A1 => n14786, A2 => n14785, ZN => n19958);
   U2525 : BUF_X1 port map( A => n15746, Z => n15182);
   U2544 : OR2_X1 port map( A1 => n14961, A2 => n15287, ZN => n19573);
   U2613 : AND2_X1 port map( A1 => n15875, A2 => n15714, ZN => n15146);
   U2668 : OR3_X1 port map( A1 => n19888, A2 => n19583, A3 => n15470, ZN => 
                           n1075);
   U2714 : OR2_X1 port map( A1 => n15467, A2 => n15470, ZN => n2358);
   U2747 : BUF_X1 port map( A => n17127, Z => n19882);
   U2762 : CLKBUF_X1 port map( A => n17547, Z => n19771);
   U2764 : NOR2_X1 port map( A1 => n19974, A2 => n19744, ZN => n18248);
   U2770 : XNOR2_X1 port map( A => n16710, B => n16709, ZN => n17818);
   U2772 : MUX2_X1 port map( A => n15269, B => n15268, S => n15846, Z => n16691
                           );
   U2778 : XNOR2_X1 port map( A => n16352, B => n16351, ZN => n18111);
   U2786 : OR2_X1 port map( A1 => n17830, A2 => n219, ZN => n18957);
   U2819 : AND2_X1 port map( A1 => n17855, A2 => n17, ZN => n15);
   U2853 : NAND2_X1 port map( A1 => n17247, A2 => n17246, ZN => n18384);
   U2858 : AND2_X1 port map( A1 => n17452, A2 => n17453, ZN => n18702);
   U2877 : OR2_X1 port map( A1 => n17750, A2 => n18929, ZN => n19574);
   U2901 : OR2_X1 port map( A1 => n18064, A2 => n19035, ZN => n2399);
   U2932 : OR2_X1 port map( A1 => n18709, A2 => n18733, ZN => n18736);
   U3018 : OAI21_X1 port map( B1 => n17177, B2 => n17176, A => n17175, ZN => 
                           n19105);
   U3064 : OAI211_X1 port map( C1 => n18381, C2 => n2274, A => n18387, B => 
                           n18386, ZN => n19969);
   U3101 : CLKBUF_X1 port map( A => Key(39), Z => n18284);
   U3109 : CLKBUF_X1 port map( A => Key(123), Z => n18075);
   U3117 : CLKBUF_X1 port map( A => Key(75), Z => n17851);
   U3122 : XOR2_X1 port map( A => n18749, B => n2381, Z => n19525);
   U3137 : AND3_X1 port map( A1 => n3085, A2 => n975, A3 => n17506, ZN => 
                           n19526);
   U3146 : NAND3_X1 port map( A1 => n12525, A2 => n3256, A3 => n182, ZN => 
                           n19527);
   U3166 : INV_X1 port map( A => n9837, ZN => n19606);
   U3168 : AND2_X1 port map( A1 => n4500, A2 => n409, ZN => n5841);
   U3180 : INV_X1 port map( A => n5841, ZN => n19968);
   U3239 : AOI22_X1 port map( A1 => n4139, A2 => n4962, B1 => n4377, B2 => 
                           n4138, ZN => n5524);
   U3256 : AND2_X1 port map( A1 => n7528, A2 => n7908, ZN => n19528);
   U3267 : INV_X1 port map( A => n5435, ZN => n19562);
   U3277 : INV_X1 port map( A => n5798, ZN => n5429);
   U3296 : INV_X1 port map( A => n9780, ZN => n19553);
   U3315 : INV_X1 port map( A => n7788, ZN => n19579);
   U3328 : AND2_X1 port map( A1 => n7562, A2 => n6705, ZN => n19529);
   U3330 : XOR2_X1 port map( A => n13112, B => n13113, Z => n19530);
   U3342 : XNOR2_X1 port map( A => n12954, B => n12953, ZN => n14641);
   U3380 : XOR2_X1 port map( A => n12712, B => n13457, Z => n19531);
   U3392 : AND2_X1 port map( A1 => n20221, A2 => n18953, ZN => n19532);
   U3434 : INV_X1 port map( A => n18656, ZN => n19624);
   U3469 : AND3_X1 port map( A1 => n18737, A2 => n18736, A3 => n18735, ZN => 
                           n19533);
   U3527 : OR2_X1 port map( A1 => n19286, A2 => n19285, ZN => n19534);
   U3583 : NAND2_X1 port map( A1 => n19536, A2 => n19535, ZN => n12914);
   U3702 : NAND2_X1 port map( A1 => n12297, A2 => n12296, ZN => n19536);
   U3709 : NAND2_X1 port map( A1 => n4248, A2 => n19540, ZN => n19539);
   U3722 : NAND2_X1 port map( A1 => n17217, A2 => n19541, ZN => n16467);
   U3756 : NAND2_X1 port map( A1 => n20135, A2 => n17211, ZN => n19541);
   U3769 : NOR2_X1 port map( A1 => n19542, A2 => n20007, ZN => n14976);
   U3870 : NAND2_X1 port map( A1 => n4570, A2 => n4370, ZN => n4509);
   U3892 : NAND2_X1 port map( A1 => n12569, A2 => n12570, ZN => n12571);
   U3916 : OAI211_X1 port map( C1 => n14227, C2 => n20376, A => n19543, B => 
                           n14412, ZN => n2903);
   U3949 : NAND2_X1 port map( A1 => n13403, A2 => n14408, ZN => n19543);
   U4009 : NAND3_X1 port map( A1 => n20464, A2 => n4697, A3 => n5040, ZN => 
                           n19544);
   U4053 : NOR2_X1 port map( A1 => n20535, A2 => n18869, ZN => n18853);
   U4119 : NAND2_X1 port map( A1 => n2891, A2 => n14703, ZN => n14380);
   U4122 : XNOR2_X1 port map( A => n17366, B => n18308, ZN => n16145);
   U4183 : XNOR2_X1 port map( A => n10286, B => n9802, ZN => n9756);
   U4191 : NAND2_X1 port map( A1 => n7577, A2 => n7576, ZN => n9802);
   U4342 : NAND2_X1 port map( A1 => n19740, A2 => n192, ZN => n15705);
   U4369 : NAND2_X1 port map( A1 => n2659, A2 => n17149, ZN => n3235);
   U4370 : NAND3_X1 port map( A1 => n2782, A2 => n2781, A3 => n2989, ZN => 
                           n19638);
   U4404 : NAND3_X1 port map( A1 => n233, A2 => n15815, A3 => n228, ZN => n3374
                           );
   U4407 : NAND2_X1 port map( A1 => n19547, A2 => n19546, ZN => n10700);
   U4452 : NAND2_X1 port map( A1 => n11292, A2 => n10697, ZN => n19546);
   U4453 : NAND2_X1 port map( A1 => n10696, A2 => n10978, ZN => n19547);
   U4456 : NAND2_X1 port map( A1 => n19549, A2 => n19548, ZN => n15852);
   U4483 : NAND2_X1 port map( A1 => n15408, A2 => n15407, ZN => n19548);
   U4518 : NAND2_X1 port map( A1 => n2791, A2 => n15616, ZN => n19549);
   U4533 : NOR2_X1 port map( A1 => n19528, A2 => n7531, ZN => n19550);
   U4566 : AOI21_X1 port map( B1 => n19525, B2 => n19803, A => n19551, ZN => 
                           n19650);
   U4665 : INV_X1 port map( A => n4144, ZN => n4398);
   U4676 : NAND2_X1 port map( A1 => n4144, A2 => n4141, ZN => n4143);
   U4683 : NAND2_X1 port map( A1 => n4914, A2 => n4140, ZN => n4144);
   U4689 : NAND2_X1 port map( A1 => n14828, A2 => n3223, ZN => n2685);
   U4690 : NAND2_X1 port map( A1 => n11348, A2 => n11349, ZN => n11352);
   U4698 : NAND2_X1 port map( A1 => n19554, A2 => n19552, ZN => n8666);
   U4734 : NAND2_X1 port map( A1 => n9782, A2 => n19553, ZN => n19552);
   U4737 : NAND2_X1 port map( A1 => n9779, A2 => n9780, ZN => n19554);
   U4742 : NAND2_X1 port map( A1 => n12151, A2 => n20618, ZN => n19555);
   U4745 : NOR2_X1 port map( A1 => n12157, A2 => n19558, ZN => n19557);
   U4768 : NAND2_X1 port map( A1 => n9068, A2 => n2504, ZN => n2502);
   U4819 : NAND2_X1 port map( A1 => n5014, A2 => n4555, ZN => n4737);
   U4914 : NAND2_X1 port map( A1 => n19562, A2 => n5704, ZN => n19561);
   U4941 : OR2_X2 port map( A1 => n4078, A2 => n4079, ZN => n5704);
   U4942 : OAI21_X1 port map( B1 => n20479, B2 => n19564, A => n19563, ZN => 
                           n10648);
   U4945 : NAND2_X1 port map( A1 => n10968, A2 => n11559, ZN => n19563);
   U5040 : NAND2_X1 port map( A1 => n9274, A2 => n20265, ZN => n19565);
   U5072 : NAND2_X1 port map( A1 => n6166, A2 => n6172, ZN => n6170);
   U5092 : NAND2_X1 port map( A1 => n19568, A2 => n19566, ZN => n10647);
   U5108 : NAND2_X1 port map( A1 => n10646, A2 => n19567, ZN => n19566);
   U5139 : INV_X1 port map( A => n10968, ZN => n19567);
   U5167 : NAND2_X1 port map( A1 => n11553, A2 => n9017, ZN => n10646);
   U5170 : NAND2_X1 port map( A1 => n10645, A2 => n10968, ZN => n19568);
   U5173 : NAND2_X1 port map( A1 => n19569, A2 => n4570, ZN => n4259);
   U5177 : NAND2_X1 port map( A1 => n4573, A2 => n4507, ZN => n19569);
   U5235 : NAND3_X1 port map( A1 => n607, A2 => n11160, A3 => n19571, ZN => 
                           n19570);
   U5300 : NAND2_X1 port map( A1 => n20012, A2 => n8282, ZN => n7601);
   U5313 : NAND2_X1 port map( A1 => n328, A2 => n3704, ZN => n15081);
   U5324 : NAND2_X1 port map( A1 => n2768, A2 => n2766, ZN => n328);
   U5359 : NAND2_X1 port map( A1 => n2414, A2 => n17866, ZN => n19238);
   U5360 : OR2_X1 port map( A1 => n10246, A2 => n11886, ZN => n2130);
   U5361 : NAND2_X1 port map( A1 => n9018, A2 => n9295, ZN => n9299);
   U5392 : OR2_X2 port map( A1 => n3261, A2 => n8514, ZN => n8676);
   U5408 : NAND2_X1 port map( A1 => n16782, A2 => n16783, ZN => n1559);
   U5447 : NAND2_X1 port map( A1 => n17069, A2 => n17896, ZN => n16783);
   U5546 : NAND2_X1 port map( A1 => n213, A2 => n18797, ZN => n2179);
   U5549 : MUX2_X1 port map( A => n6195, B => n6196, S => n5382, Z => n6197);
   U5592 : NAND2_X1 port map( A1 => n14287, A2 => n241, ZN => n1976);
   U5678 : NAND3_X1 port map( A1 => n114, A2 => n20128, A3 => n18037, ZN => 
                           n19575);
   U5745 : OR2_X2 port map( A1 => n4316, A2 => n19576, ZN => n5633);
   U5751 : NAND2_X1 port map( A1 => n4314, A2 => n4362, ZN => n19576);
   U5761 : NAND2_X1 port map( A1 => n12203, A2 => n125, ZN => n1190);
   U5774 : AND2_X1 port map( A1 => n14032, A2 => n14637, ZN => n13985);
   U5832 : NAND2_X1 port map( A1 => n19579, A2 => n8299, ZN => n19578);
   U5837 : NAND2_X1 port map( A1 => n885, A2 => n8990, ZN => n9272);
   U5865 : NAND2_X1 port map( A1 => n2539, A2 => n2538, ZN => n19580);
   U5869 : NAND2_X1 port map( A1 => n4441, A2 => n2670, ZN => n1922);
   U5928 : NAND2_X1 port map( A1 => n4160, A2 => n4524, ZN => n19581);
   U5949 : INV_X1 port map( A => n15468, ZN => n19583);
   U5953 : NAND2_X1 port map( A1 => n19584, A2 => n11688, ZN => n13622);
   U5990 : INV_X1 port map( A => n12576, ZN => n19585);
   U6016 : NOR2_X1 port map( A1 => n19601, A2 => n19600, ZN => n13973);
   U6017 : OAI211_X2 port map( C1 => n16778, C2 => n17176, A => n19587, B => 
                           n19586, ZN => n19144);
   U6034 : NAND2_X1 port map( A1 => n3293, A2 => n20239, ZN => n19586);
   U6073 : NAND2_X1 port map( A1 => n16777, A2 => n19667, ZN => n19587);
   U6109 : NAND2_X1 port map( A1 => n1471, A2 => n11831, ZN => n13843);
   U6139 : NAND2_X1 port map( A1 => n824, A2 => n823, ZN => n8419);
   U6193 : NAND2_X1 port map( A1 => n8003, A2 => n7591, ZN => n7477);
   U6208 : XNOR2_X1 port map( A => n19588, B => n19410, ZN => n7217);
   U6209 : NAND2_X1 port map( A1 => n5245, A2 => n5244, ZN => n19588);
   U6224 : INV_X1 port map( A => n352, ZN => n19590);
   U6232 : NAND3_X1 port map( A1 => n771, A2 => n772, A3 => n8665, ZN => n419);
   U6248 : OAI211_X1 port map( C1 => n8354, C2 => n8359, A => n19591, B => 
                           n7504, ZN => n6902);
   U6287 : NAND2_X1 port map( A1 => n19651, A2 => n8354, ZN => n19591);
   U6289 : NAND3_X1 port map( A1 => n12379, A2 => n12378, A3 => n19592, ZN => 
                           n13600);
   U6342 : NAND2_X1 port map( A1 => n2333, A2 => n2332, ZN => n12378);
   U6356 : NAND2_X1 port map( A1 => n3560, A2 => n19593, ZN => n1720);
   U6382 : NOR2_X1 port map( A1 => n4865, A2 => n19523, ZN => n19593);
   U6393 : XNOR2_X1 port map( A => n19594, B => n18848, ZN => n9761);
   U6396 : NAND3_X1 port map( A1 => n8170, A2 => n8168, A3 => n8169, ZN => 
                           n19594);
   U6397 : NAND2_X1 port map( A1 => n9832, A2 => n11263, ZN => n1132);
   U6405 : NAND2_X1 port map( A1 => n755, A2 => n756, ZN => n9832);
   U6427 : NAND2_X1 port map( A1 => n20129, A2 => n18976, ZN => n17310);
   U6441 : NAND2_X1 port map( A1 => n8659, A2 => n8658, ZN => n19595);
   U6458 : NAND2_X1 port map( A1 => n3519, A2 => n8660, ZN => n19596);
   U6487 : NAND2_X1 port map( A1 => n8134, A2 => n8135, ZN => n8136);
   U6513 : NOR2_X2 port map( A1 => n2776, A2 => n8570, ZN => n10254);
   U6555 : OAI22_X1 port map( A1 => n20468, A2 => n12101, B1 => n11271, B2 => 
                           n10684, ZN => n9659);
   U6560 : NOR2_X1 port map( A1 => n19984, A2 => n19598, ZN => n19597);
   U6562 : OAI21_X2 port map( B1 => n3961, B2 => n5408, A => n1182, ZN => n7304
                           );
   U6592 : OAI21_X2 port map( B1 => n9933, B2 => n11522, A => n9932, ZN => 
                           n12004);
   U6607 : OR2_X1 port map( A1 => n15179, A2 => n15181, ZN => n19599);
   U6610 : OAI21_X1 port map( B1 => n6020, B2 => n6021, A => n19660, ZN => n445
                           );
   U6626 : NAND2_X1 port map( A1 => n3246, A2 => n14522, ZN => n19601);
   U6645 : NAND2_X1 port map( A1 => n2529, A2 => n2530, ZN => n2528);
   U6670 : NAND2_X1 port map( A1 => n19602, A2 => n12641, ZN => n12643);
   U6686 : NAND2_X1 port map( A1 => n389, A2 => n12640, ZN => n19602);
   U6699 : NAND2_X1 port map( A1 => n2387, A2 => n2386, ZN => n7624);
   U6703 : NAND2_X1 port map( A1 => n12569, A2 => n12258, ZN => n19603);
   U6730 : NAND2_X1 port map( A1 => n2065, A2 => n8602, ZN => n19604);
   U6745 : NAND2_X1 port map( A1 => n3328, A2 => n348, ZN => n3327);
   U6754 : NAND2_X1 port map( A1 => n20504, A2 => n8064, ZN => n1433);
   U6765 : OR2_X1 port map( A1 => n14098, A2 => n14338, ZN => n19607);
   U6766 : OAI21_X1 port map( B1 => n14096, B2 => n14095, A => n14094, ZN => 
                           n19608);
   U6789 : OR2_X1 port map( A1 => n14103, A2 => n14787, ZN => n14063);
   U6803 : XNOR2_X1 port map( A => n19609, B => n13135, ZN => n3364);
   U6807 : XNOR2_X1 port map( A => n3365, B => n13651, ZN => n19609);
   U6822 : XNOR2_X1 port map( A => n19610, B => n19103, ZN => Ciphertext(128));
   U6844 : NOR2_X2 port map( A1 => n19611, A2 => n15640, ZN => n16412);
   U6860 : NAND3_X1 port map( A1 => n6055, A2 => n5785, A3 => n5891, ZN => 
                           n3865);
   U6863 : NAND3_X1 port map( A1 => n3838, A2 => n1137, A3 => n19612, ZN => 
                           n5782);
   U6890 : NAND2_X1 port map( A1 => n14223, A2 => n14224, ZN => n14225);
   U6904 : NAND2_X1 port map( A1 => n9063, A2 => n19805, ZN => n2300);
   U6917 : NAND2_X1 port map( A1 => n3072, A2 => n1765, ZN => n9063);
   U6924 : NAND3_X1 port map( A1 => n12572, A2 => n12017, A3 => n242, ZN => 
                           n12019);
   U6986 : MUX2_X1 port map( A => n14823, B => n14822, S => n14821, Z => n19613
                           );
   U7026 : AOI21_X1 port map( B1 => n10912, B2 => n9487, A => n19614, ZN => 
                           n9490);
   U7028 : NAND3_X1 port map( A1 => n19615, A2 => n1009, A3 => n12562, ZN => 
                           n11895);
   U7030 : NAND2_X1 port map( A1 => n3733, A2 => n12262, ZN => n19615);
   U7039 : OAI22_X1 port map( A1 => n15817, A2 => n19958, B1 => n15816, B2 => 
                           n15815, ZN => n2114);
   U7058 : NAND2_X1 port map( A1 => n19617, A2 => n19616, ZN => n5410);
   U7065 : NAND2_X1 port map( A1 => n4889, A2 => n4888, ZN => n19616);
   U7098 : NAND2_X1 port map( A1 => n4891, A2 => n4890, ZN => n19617);
   U7103 : NAND2_X1 port map( A1 => n11951, A2 => n11598, ZN => n11957);
   U7109 : NAND2_X1 port map( A1 => n20367, A2 => n7480, ZN => n7483);
   U7111 : XNOR2_X1 port map( A => n13768, B => n13600, ZN => n13282);
   U7138 : NOR2_X1 port map( A1 => n10830, A2 => n11421, ZN => n10831);
   U7141 : NAND2_X1 port map( A1 => n385, A2 => n5893, ZN => n7258);
   U7160 : OAI21_X1 port map( B1 => n2120, B2 => n18024, A => n19618, ZN => 
                           n18027);
   U7169 : NAND2_X1 port map( A1 => n18928, A2 => n18024, ZN => n19618);
   U7170 : NAND2_X1 port map( A1 => n7674, A2 => n8365, ZN => n7510);
   U7171 : XNOR2_X2 port map( A => n6395, B => n6394, ZN => n7674);
   U7172 : NAND2_X1 port map( A1 => n11604, A2 => n12416, ZN => n11608);
   U7179 : NAND2_X1 port map( A1 => n11603, A2 => n20350, ZN => n11604);
   U7242 : MUX2_X1 port map( A => n4304, B => n4303, S => n4982, Z => n19619);
   U7244 : OAI21_X1 port map( B1 => n19110, B2 => n19532, A => n19620, ZN => 
                           n17712);
   U7245 : NAND2_X1 port map( A1 => n19110, A2 => n17710, ZN => n19620);
   U7258 : NAND3_X1 port map( A1 => n3028, A2 => n3030, A3 => n20117, ZN => 
                           n3027);
   U7265 : NAND3_X1 port map( A1 => n19621, A2 => n3701, A3 => n2482, ZN => 
                           n3700);
   U7266 : NAND3_X1 port map( A1 => n286, A2 => n5746, A3 => n5745, ZN => 
                           n19621);
   U7275 : NAND2_X1 port map( A1 => n19623, A2 => n19622, ZN => n3791);
   U7280 : NAND2_X1 port map( A1 => n3793, A2 => n3795, ZN => n19623);
   U7288 : NAND2_X1 port map( A1 => n19625, A2 => n19624, ZN => n18658);
   U7289 : NAND2_X1 port map( A1 => n18648, A2 => n19935, ZN => n19625);
   U7311 : XNOR2_X1 port map( A => n19627, B => n19626, ZN => Ciphertext(168));
   U7352 : INV_X1 port map( A => n2455, ZN => n19626);
   U7363 : NAND2_X1 port map( A1 => n19633, A2 => n19629, ZN => n19283);
   U7372 : INV_X1 port map( A => n19630, ZN => n19629);
   U7382 : AOI21_X1 port map( B1 => n19632, B2 => n19631, A => n19400, ZN => 
                           n19630);
   U7448 : NAND2_X1 port map( A1 => n19391, A2 => n19390, ZN => n19632);
   U7462 : NAND2_X1 port map( A1 => n17618, A2 => n19400, ZN => n19633);
   U7468 : INV_X1 port map( A => n951, ZN => n19634);
   U7482 : XNOR2_X1 port map( A => n19635, B => n3460, ZN => n13007);
   U7487 : XNOR2_X1 port map( A => n13703, B => n19796, ZN => n19635);
   U7488 : XNOR2_X2 port map( A => n19637, B => n19636, ZN => n11234);
   U7492 : XNOR2_X1 port map( A => n10158, B => n9864, ZN => n19636);
   U7497 : XNOR2_X1 port map( A => n9992, B => n9863, ZN => n19637);
   U7559 : NAND2_X1 port map( A1 => n332, A2 => n333, ZN => n11345);
   U7668 : NAND3_X2 port map( A1 => n19638, A2 => n6959, A3 => n6958, ZN => 
                           n10249);
   U7678 : NAND2_X1 port map( A1 => n19639, A2 => n1616, ZN => n8977);
   U7695 : OAI21_X1 port map( B1 => n8970, B2 => n1618, A => n9252, ZN => 
                           n19639);
   U7708 : OR2_X1 port map( A1 => n11866, A2 => n11870, ZN => n9776);
   U7774 : INV_X1 port map( A => n18691, ZN => n19640);
   U7796 : NAND2_X1 port map( A1 => n7820, A2 => n278, ZN => n7521);
   U7817 : NAND2_X1 port map( A1 => n19641, A2 => n7755, ZN => n2259);
   U7825 : OAI22_X1 port map( A1 => n7909, A2 => n6904, B1 => n19521, B2 => 
                           n7754, ZN => n19641);
   U7859 : OAI21_X1 port map( B1 => n249, B2 => n12354, A => n12174, ZN => 
                           n11656);
   U7889 : NAND2_X1 port map( A1 => n12354, A2 => n12352, ZN => n12174);
   U7890 : NAND2_X1 port map( A1 => n7831, A2 => n7832, ZN => n9007);
   U7918 : NAND2_X1 port map( A1 => n19643, A2 => n19642, ZN => n13743);
   U7944 : NAND2_X1 port map( A1 => n13730, A2 => n14381, ZN => n19642);
   U7945 : NAND2_X1 port map( A1 => n13731, A2 => n19644, ZN => n19643);
   U7946 : INV_X1 port map( A => n14381, ZN => n19644);
   U7953 : OAI21_X1 port map( B1 => n635, B2 => n19645, A => n634, ZN => n16580
                           );
   U7959 : OAI21_X1 port map( B1 => n20436, B2 => n19372, A => n19646, ZN => 
                           n19645);
   U8004 : INV_X1 port map( A => n19370, ZN => n19647);
   U8017 : AOI21_X1 port map( B1 => n19648, B2 => n11109, A => n11106, ZN => 
                           n10772);
   U8041 : NAND2_X1 port map( A1 => n11429, A2 => n11041, ZN => n19648);
   U8042 : OR2_X2 port map( A1 => n9231, A2 => n9230, ZN => n9987);
   U8043 : NAND3_X1 port map( A1 => n19649, A2 => n18241, A3 => n18240, ZN => 
                           n18246);
   U8046 : NAND2_X1 port map( A1 => n20132, A2 => n18238, ZN => n19649);
   U8068 : AOI21_X1 port map( B1 => n19650, B2 => n19533, A => n18747, ZN => 
                           Ciphertext(80));
   U8069 : NAND3_X1 port map( A1 => n2174, A2 => n9331, A3 => n8866, ZN => 
                           n8867);
   U8133 : NAND2_X1 port map( A1 => n19057, A2 => n19067, ZN => n71);
   U8141 : NAND3_X1 port map( A1 => n1812, A2 => n11113, A3 => n11452, ZN => 
                           n1804);
   U8178 : BUF_X2 port map( A => n18287, Z => n18362);
   U8196 : AND2_X1 port map( A1 => n19163, A2 => n19162, ZN => n17790);
   U8223 : XNOR2_X1 port map( A => n13112, B => n13113, ZN => n19652);
   U8262 : INV_X1 port map( A => n19069, ZN => n19653);
   U8281 : NAND2_X1 port map( A1 => n18944, A2 => n2062, ZN => n19654);
   U8361 : OAI211_X2 port map( C1 => n18633, C2 => n959, A => n1069, B => n1013
                           , ZN => n18592);
   U8366 : OAI211_X1 port map( C1 => n17161, C2 => n16792, A => n16791, B => 
                           n18542, ZN => n19655);
   U8373 : XOR2_X1 port map( A => n9842, B => n10299, Z => n8509);
   U8377 : XNOR2_X1 port map( A => n13057, B => n13018, ZN => n13457);
   U8385 : XNOR2_X1 port map( A => n12712, B => n13457, ZN => n19657);
   U8405 : XOR2_X1 port map( A => n9503, B => n8548, Z => n8567);
   U8422 : NAND2_X1 port map( A1 => n18944, A2 => n2062, ZN => n19001);
   U8430 : OAI21_X1 port map( B1 => n3576, B2 => n13943, A => n13942, ZN => 
                           n19659);
   U8434 : OAI21_X1 port map( B1 => n3576, B2 => n13943, A => n13942, ZN => 
                           n16974);
   U8444 : OR2_X1 port map( A1 => n3569, A2 => n5823, ZN => n19660);
   U8503 : AND2_X1 port map( A1 => n16799, A2 => n16798, ZN => n19661);
   U8514 : AOI22_X1 port map( A1 => n14084, A2 => n20500, B1 => n14081, B2 => 
                           n14082, ZN => n15515);
   U8562 : OR2_X1 port map( A1 => n9241, A2 => n9240, ZN => n19663);
   U8597 : CLKBUF_X1 port map( A => n18916, Z => n19664);
   U8652 : NOR2_X1 port map( A1 => n17153, A2 => n17152, ZN => n19665);
   U8654 : NOR2_X1 port map( A1 => n17153, A2 => n17152, ZN => n18590);
   U8661 : OR2_X1 port map( A1 => n12003, A2 => n1637, ZN => n3239);
   U8664 : XNOR2_X1 port map( A => n16559, B => n16558, ZN => n19371);
   U8676 : XNOR2_X1 port map( A => n16065, B => n16064, ZN => n16308);
   U8716 : XOR2_X1 port map( A => n15953, B => n15954, Z => n19667);
   U8737 : CLKBUF_X1 port map( A => Key(173), Z => n19140);
   U8772 : OR2_X1 port map( A1 => n17153, A2 => n17152, ZN => n19669);
   U8798 : NOR2_X1 port map( A1 => n19010, A2 => n19670, ZN => n2050);
   U8810 : AND3_X1 port map( A1 => n19011, A2 => n19654, A3 => n19687, ZN => 
                           n19670);
   U8857 : XNOR2_X1 port map( A => n16399, B => n16400, ZN => n19672);
   U8877 : OAI21_X1 port map( B1 => n17555, B2 => n18106, A => n17554, ZN => 
                           n19673);
   U8995 : XNOR2_X1 port map( A => n16223, B => n16222, ZN => n19675);
   U8998 : XNOR2_X1 port map( A => n16223, B => n16222, ZN => n17494);
   U9068 : OAI211_X1 port map( C1 => n15807, C2 => n15808, A => n15805, B => 
                           n19966, ZN => n16982);
   U9122 : INV_X1 port map( A => n15420, ZN => n19676);
   U9125 : XNOR2_X1 port map( A => n16230, B => n16229, ZN => n17493);
   U9224 : XOR2_X1 port map( A => n17448, B => n17447, Z => n19678);
   U9225 : NAND2_X1 port map( A1 => n17557, A2 => n2797, ZN => n19679);
   U9262 : OAI21_X1 port map( B1 => n18973, B2 => n220, A => n18972, ZN => 
                           n19680);
   U9382 : CLKBUF_X1 port map( A => n18306, Z => n19683);
   U9444 : XNOR2_X1 port map( A => n16694, B => n16693, ZN => n19684);
   U9497 : NAND2_X1 port map( A1 => n102, A2 => n17820, ZN => n19685);
   U9595 : XNOR2_X1 port map( A => n16694, B => n16693, ZN => n18968);
   U9791 : BUF_X1 port map( A => n7443, Z => n19686);
   U9967 : XNOR2_X1 port map( A => n5423, B => n5422, ZN => n7443);
   U10006 : OAI211_X1 port map( C1 => n18960, C2 => n18959, A => n18958, B => 
                           n18957, ZN => n19687);
   U10071 : OAI211_X1 port map( C1 => n18960, C2 => n18959, A => n18958, B => 
                           n18957, ZN => n19009);
   U10097 : XNOR2_X2 port map( A => n3851, B => Key(77), ZN => n19688);
   U10107 : OAI21_X1 port map( B1 => n922, B2 => n12457, A => n12456, ZN => 
                           n19689);
   U10196 : XNOR2_X1 port map( A => n3851, B => Key(77), ZN => n5258);
   U10261 : OAI21_X1 port map( B1 => n922, B2 => n12457, A => n12456, ZN => 
                           n13584);
   U10351 : AND2_X1 port map( A1 => n18540, A2 => n18541, ZN => n19690);
   U10360 : OAI21_X1 port map( B1 => n2691, B2 => n16804, A => n16803, ZN => 
                           n19691);
   U10453 : OAI21_X1 port map( B1 => n2691, B2 => n16804, A => n16803, ZN => 
                           n18546);
   U10788 : INV_X1 port map( A => n12332, ZN => n12335);
   U10970 : OR2_X1 port map( A1 => n15879, A2 => n15153, ZN => n14924);
   U10979 : OAI21_X1 port map( B1 => n17068, B2 => n17067, A => n17066, ZN => 
                           n19692);
   U10994 : OAI21_X1 port map( B1 => n17068, B2 => n17067, A => n17066, ZN => 
                           n19155);
   U11000 : NAND4_X2 port map( A1 => n1207, A2 => n1573, A3 => n968, A4 => 
                           n1209, ZN => n15714);
   U11192 : AND2_X1 port map( A1 => n15750, A2 => n25, ZN => n16044);
   U11236 : INV_X1 port map( A => n14350, ZN => n19693);
   U11403 : XNOR2_X1 port map( A => n12806, B => n12805, ZN => n14327);
   U11453 : AND2_X1 port map( A1 => n2647, A2 => n12122, ZN => n19694);
   U11471 : OR2_X1 port map( A1 => n13896, A2 => n13895, ZN => n28);
   U11512 : OR2_X1 port map( A1 => n17495, A2 => n17492, ZN => n19695);
   U11618 : OR2_X1 port map( A1 => n15313, A2 => n14620, ZN => n1266);
   U11724 : AND3_X1 port map( A1 => n3528, A2 => n5685, A3 => n3527, ZN => 
                           n19698);
   U11728 : AND3_X1 port map( A1 => n3528, A2 => n5685, A3 => n3527, ZN => 
                           n19699);
   U11806 : OAI21_X1 port map( B1 => n5326, B2 => n5327, A => n5325, ZN => 
                           n7041);
   U11881 : XNOR2_X1 port map( A => n14376, B => n14375, ZN => n19700);
   U11906 : INV_X1 port map( A => n20003, ZN => n19702);
   U11922 : OAI21_X1 port map( B1 => n14848, B2 => n16172, A => n14847, ZN => 
                           n18400);
   U11955 : XOR2_X1 port map( A => n12953, B => n12954, Z => n19703);
   U11970 : OAI211_X1 port map( C1 => n14838, C2 => n14534, A => n14533, B => 
                           n14532, ZN => n19704);
   U11982 : OAI211_X1 port map( C1 => n14838, C2 => n14534, A => n14533, B => 
                           n14532, ZN => n19705);
   U12026 : NAND2_X1 port map( A1 => n14881, A2 => n1490, ZN => n19706);
   U12029 : NAND2_X1 port map( A1 => n14881, A2 => n1490, ZN => n17340);
   U12095 : OAI21_X1 port map( B1 => n10843, B2 => n1812, A => n10842, ZN => 
                           n12589);
   U12139 : AND2_X1 port map( A1 => n14154, A2 => n14393, ZN => n19709);
   U12151 : XOR2_X1 port map( A => n10552, B => n10582, Z => n9760);
   U12159 : AND2_X1 port map( A1 => n7849, A2 => n7850, ZN => n19710);
   U12163 : NAND2_X1 port map( A1 => n17771, A2 => n17770, ZN => n19711);
   U12210 : NAND2_X1 port map( A1 => n17771, A2 => n17770, ZN => n18794);
   U12272 : NOR2_X1 port map( A1 => n17669, A2 => n19249, ZN => n19276);
   U12275 : AOI21_X2 port map( B1 => n15578, B2 => n693, A => n692, ZN => 
                           n19713);
   U12347 : AOI21_X1 port map( B1 => n15578, B2 => n693, A => n692, ZN => 
                           n17348);
   U12389 : NOR2_X1 port map( A1 => n6206, A2 => n19492, ZN => n5839);
   U12401 : XNOR2_X1 port map( A => n10189, B => n10190, ZN => n11430);
   U12596 : NAND2_X1 port map( A1 => n102, A2 => n17820, ZN => n19068);
   U12625 : AND2_X1 port map( A1 => n737, A2 => n7509, ZN => n19715);
   U12668 : NAND4_X1 port map( A1 => n9281, A2 => n9279, A3 => n9282, A4 => 
                           n9280, ZN => n19717);
   U12767 : NAND4_X1 port map( A1 => n9281, A2 => n9279, A3 => n9282, A4 => 
                           n9280, ZN => n19718);
   U12875 : XNOR2_X1 port map( A => n10585, B => n10586, ZN => n19719);
   U12877 : NAND4_X1 port map( A1 => n9281, A2 => n9279, A3 => n9282, A4 => 
                           n9280, ZN => n10490);
   U12903 : NOR2_X1 port map( A1 => n15469, A2 => n15465, ZN => n15234);
   U12916 : OAI21_X1 port map( B1 => n12171, B2 => n12172, A => n12170, ZN => 
                           n19721);
   U12917 : OR2_X1 port map( A1 => n14291, A2 => n129, ZN => n19722);
   U12972 : OAI21_X1 port map( B1 => n12171, B2 => n12172, A => n12170, ZN => 
                           n13721);
   U12975 : XNOR2_X1 port map( A => n17039, B => n17038, ZN => n19723);
   U13093 : AND2_X1 port map( A1 => n18944, A2 => n2062, ZN => n19724);
   U13099 : XNOR2_X1 port map( A => n17039, B => n17038, ZN => n18019);
   U13253 : XNOR2_X1 port map( A => n10111, B => n10110, ZN => n19725);
   U13273 : OAI211_X1 port map( C1 => n10817, C2 => n19949, A => n1357, B => 
                           n1356, ZN => n19726);
   U13503 : OAI211_X1 port map( C1 => n10817, C2 => n19949, A => n1357, B => 
                           n1356, ZN => n948);
   U13535 : XNOR2_X1 port map( A => n13478, B => n13477, ZN => n19727);
   U13536 : XNOR2_X1 port map( A => n13478, B => n13477, ZN => n19728);
   U13547 : XNOR2_X1 port map( A => n13477, B => n13478, ZN => n14746);
   U13580 : XNOR2_X1 port map( A => n6966, B => n7211, ZN => n6883);
   U13630 : NAND2_X1 port map( A1 => n5261, A2 => n2175, ZN => n19730);
   U13643 : NAND2_X1 port map( A1 => n5261, A2 => n2175, ZN => n6867);
   U13692 : BUF_X1 port map( A => n8828, Z => n19896);
   U13697 : XNOR2_X1 port map( A => n13627, B => n13628, ZN => n19731);
   U13743 : XNOR2_X1 port map( A => n13627, B => n13628, ZN => n14393);
   U13779 : NOR2_X1 port map( A1 => n19763, A2 => n18394, ZN => n1296);
   U14010 : XNOR2_X1 port map( A => n20519, B => n16576, ZN => n19733);
   U14108 : XNOR2_X1 port map( A => n16577, B => n16576, ZN => n19380);
   U14109 : BUF_X1 port map( A => n13029, Z => n19734);
   U14149 : OAI21_X1 port map( B1 => n19919, B2 => n17983, A => n3206, ZN => 
                           n19735);
   U14157 : OAI21_X1 port map( B1 => n19919, B2 => n17983, A => n3206, ZN => 
                           n18673);
   U14178 : XOR2_X1 port map( A => n9428, B => n9944, Z => n19736);
   U14209 : XNOR2_X1 port map( A => n16387, B => n16693, ZN => n19737);
   U14281 : AND2_X1 port map( A1 => n19462, A2 => n19463, ZN => n19738);
   U14365 : AND3_X1 port map( A1 => n13958, A2 => n13956, A3 => n402, ZN => 
                           n19740);
   U14494 : XOR2_X1 port map( A => n7288, B => n6410, Z => n19741);
   U14495 : XOR2_X1 port map( A => n13024, B => n13023, Z => n19742);
   U14500 : NOR2_X1 port map( A1 => n15360, A2 => n15359, ZN => n19743);
   U14503 : NOR2_X1 port map( A1 => n15360, A2 => n15359, ZN => n16359);
   U14512 : XNOR2_X1 port map( A => n17106, B => n17105, ZN => n19876);
   U14550 : XNOR2_X1 port map( A => n17421, B => n17422, ZN => n19744);
   U14581 : NOR2_X1 port map( A1 => n18136, A2 => n18135, ZN => n18650);
   U14599 : NAND2_X1 port map( A1 => n8922, A2 => n2301, ZN => n19746);
   U14698 : BUF_X1 port map( A => n14548, Z => n19748);
   U14787 : NAND2_X1 port map( A1 => n16501, A2 => n16500, ZN => n19749);
   U14788 : XNOR2_X1 port map( A => n9758, B => n9757, ZN => n19750);
   U14789 : NOR2_X1 port map( A1 => n17397, A2 => n17398, ZN => n19751);
   U14790 : XNOR2_X1 port map( A => n9758, B => n9757, ZN => n11390);
   U14861 : NOR2_X1 port map( A1 => n17398, A2 => n17397, ZN => n18703);
   U14930 : AND2_X1 port map( A1 => n328, A2 => n3704, ZN => n19752);
   U14983 : NAND2_X1 port map( A1 => n17452, A2 => n17453, ZN => n19753);
   U14984 : AND2_X1 port map( A1 => n17875, A2 => n17874, ZN => n19754);
   U15028 : OAI21_X1 port map( B1 => n10853, B2 => n11367, A => n11365, ZN => 
                           n19755);
   U15048 : NAND2_X1 port map( A1 => n1590, A2 => n10873, ZN => n19756);
   U15085 : OAI21_X1 port map( B1 => n10853, B2 => n11367, A => n11365, ZN => 
                           n1590);
   U15125 : NAND2_X1 port map( A1 => n1590, A2 => n10873, ZN => n12242);
   U15132 : OAI21_X1 port map( B1 => n20429, B2 => n17573, A => n17571, ZN => 
                           n19757);
   U15337 : OAI21_X1 port map( B1 => n20429, B2 => n17573, A => n17571, ZN => 
                           n18621);
   U15377 : OAI211_X1 port map( C1 => n12884, C2 => n2039, A => n12883, B => 
                           n12882, ZN => n12888);
   U15466 : NAND2_X1 port map( A1 => n17478, A2 => n17477, ZN => n19758);
   U15485 : NAND2_X1 port map( A1 => n17478, A2 => n17477, ZN => n18518);
   U15486 : BUF_X1 port map( A => n15349, Z => n19759);
   U15518 : AOI21_X1 port map( B1 => n14501, B2 => n13509, A => n13508, ZN => 
                           n15349);
   U15520 : OAI211_X1 port map( C1 => n9451, C2 => n6442, A => n6441, B => 
                           n6440, ZN => n19760);
   U15523 : XOR2_X1 port map( A => n13614, B => n13613, Z => n19761);
   U15544 : XNOR2_X1 port map( A => n15978, B => n15977, ZN => n17873);
   U15601 : AND2_X1 port map( A1 => n17247, A2 => n17246, ZN => n19763);
   U15759 : OAI21_X1 port map( B1 => n17307, B2 => n18241, A => n20093, ZN => 
                           n19766);
   U15781 : NOR2_X1 port map( A1 => n7738, A2 => n7737, ZN => n19767);
   U15818 : OR2_X1 port map( A1 => n8402, A2 => n8401, ZN => n19768);
   U15837 : NOR2_X1 port map( A1 => n7738, A2 => n7737, ZN => n9792);
   U15851 : OR2_X1 port map( A1 => n8402, A2 => n8401, ZN => n12353);
   U15930 : OAI211_X1 port map( C1 => n17757, C2 => n17756, A => n17755, B => 
                           n17754, ZN => n19770);
   U15958 : OAI211_X1 port map( C1 => n17757, C2 => n17756, A => n17755, B => 
                           n17754, ZN => n18806);
   U16103 : XOR2_X1 port map( A => n13595, B => n13598, Z => n13606);
   U16249 : NAND2_X1 port map( A1 => n15498, A2 => n15500, ZN => n460);
   U16260 : NAND4_X2 port map( A1 => n15478, A2 => n15476, A3 => n15477, A4 => 
                           n375, ZN => n17401);
   U16272 : XNOR2_X1 port map( A => n16422, B => n16519, ZN => n19774);
   U16336 : XNOR2_X1 port map( A => n16422, B => n16519, ZN => n18093);
   U16373 : XNOR2_X1 port map( A => n4030, B => Key(113), ZN => n19776);
   U16390 : XNOR2_X1 port map( A => n4030, B => Key(113), ZN => n19777);
   U16467 : XNOR2_X1 port map( A => n4030, B => Key(113), ZN => n4701);
   U16521 : XNOR2_X1 port map( A => n9406, B => n9405, ZN => n19779);
   U16523 : XNOR2_X1 port map( A => n9406, B => n9405, ZN => n10694);
   U16583 : OAI21_X1 port map( B1 => n5857, B2 => n6159, A => n2795, ZN => 
                           n19780);
   U16597 : OAI21_X1 port map( B1 => n5857, B2 => n6159, A => n2795, ZN => 
                           n7137);
   U16642 : XNOR2_X1 port map( A => n11625, B => n11626, ZN => n19781);
   U16692 : OAI21_X1 port map( B1 => n14918, B2 => n14917, A => n148, ZN => 
                           n19782);
   U16746 : OAI21_X1 port map( B1 => n14918, B2 => n14917, A => n148, ZN => 
                           n19783);
   U16807 : XNOR2_X1 port map( A => n11625, B => n11626, ZN => n14810);
   U16881 : BUF_X1 port map( A => n12617, Z => n19784);
   U16900 : XOR2_X1 port map( A => n16981, B => n17035, Z => n17337);
   U16924 : XNOR2_X1 port map( A => n17344, B => n17343, ZN => n18257);
   U16945 : OAI211_X1 port map( C1 => n8958, C2 => n8505, A => n8504, B => 
                           n8503, ZN => n19785);
   U17058 : OAI211_X1 port map( C1 => n8958, C2 => n8505, A => n8504, B => 
                           n8503, ZN => n19786);
   U17083 : XNOR2_X1 port map( A => n17344, B => n17343, ZN => n19787);
   U17105 : XNOR2_X1 port map( A => Key(135), B => Plaintext(135), ZN => n5023)
                           ;
   U17113 : OAI21_X1 port map( B1 => n5011, B2 => n5010, A => n5009, ZN => 
                           n19789);
   U17159 : OAI21_X1 port map( B1 => n5011, B2 => n5010, A => n5009, ZN => 
                           n19790);
   U17181 : OAI21_X1 port map( B1 => n5011, B2 => n5010, A => n5009, ZN => 
                           n6031);
   U17200 : AND2_X1 port map( A1 => n16467, A2 => n60, ZN => n19791);
   U17290 : NOR2_X1 port map( A1 => n11596, A2 => n11597, ZN => n19792);
   U17304 : NOR2_X1 port map( A1 => n11596, A2 => n11597, ZN => n12861);
   U17409 : BUF_X1 port map( A => n18842, Z => n19794);
   U17410 : OAI21_X1 port map( B1 => n17320, B2 => n18033, A => n3691, ZN => 
                           n18842);
   U17480 : AOI21_X1 port map( B1 => n12329, B2 => n12328, A => n13269, ZN => 
                           n19797);
   U17488 : NAND4_X1 port map( A1 => n15689, A2 => n15691, A3 => n15690, A4 => 
                           n93, ZN => n19798);
   U17500 : NAND4_X1 port map( A1 => n15689, A2 => n15691, A3 => n15690, A4 => 
                           n93, ZN => n19799);
   U17576 : NAND4_X1 port map( A1 => n15689, A2 => n15691, A3 => n15690, A4 => 
                           n93, ZN => n17379);
   U17643 : INV_X1 port map( A => n8196, ZN => n19802);
   U17667 : NAND3_X1 port map( A1 => n18247, A2 => n18246, A3 => n18245, ZN => 
                           n19803);
   U17713 : BUF_X1 port map( A => n5524, Z => n19804);
   U17729 : INV_X1 port map( A => n8830, ZN => n19805);
   U17809 : BUF_X1 port map( A => n10199, Z => n19806);
   U17912 : AOI22_X1 port map( A1 => n8679, A2 => n8830, B1 => n8678, B2 => 
                           n9060, ZN => n10199);
   U17960 : OAI211_X1 port map( C1 => n15332, C2 => n15866, A => n15331, B => 
                           n15330, ZN => n19807);
   U17981 : OAI211_X1 port map( C1 => n15332, C2 => n15866, A => n15331, B => 
                           n15330, ZN => n17252);
   U18024 : NOR2_X1 port map( A1 => n6049, A2 => n6048, ZN => n5330);
   U18071 : XNOR2_X1 port map( A => n6448, B => n6447, ZN => n8221);
   U18072 : OAI21_X1 port map( B1 => n2326, B2 => n2325, A => n2324, ZN => 
                           n7405);
   U18180 : BUF_X1 port map( A => n8098, Z => n8238);
   U18211 : XNOR2_X2 port map( A => n1693, B => n6841, ZN => n8157);
   U18249 : NAND3_X2 port map( A1 => n601, A2 => n17594, A3 => n17593, ZN => 
                           n19284);
   U18273 : XOR2_X1 port map( A => n13776, B => n13369, Z => n2521);
   U18287 : AND2_X1 port map( A1 => n17763, A2 => n17762, ZN => n19811);
   U18292 : XOR2_X1 port map( A => n6289, B => n6288, Z => n19812);
   U18313 : OAI211_X1 port map( C1 => n20206, C2 => n13867, A => n1790, B => 
                           n1789, ZN => n15502);
   U18318 : CLKBUF_X1 port map( A => n17497, Z => n19814);
   U18348 : INV_X1 port map( A => n18497, ZN => n19816);
   U18352 : XNOR2_X1 port map( A => n15526, B => n15525, ZN => n17497);
   U18355 : XOR2_X1 port map( A => n9409, B => n9410, Z => n19817);
   U18366 : OAI21_X1 port map( B1 => n8766, B2 => n8765, A => n8764, ZN => 
                           n19818);
   U18375 : XNOR2_X1 port map( A => n12719, B => n12718, ZN => n19819);
   U18437 : XNOR2_X1 port map( A => n2488, B => Key(17), ZN => n19822);
   U18469 : XNOR2_X1 port map( A => n2488, B => Key(17), ZN => n4302);
   U18470 : XNOR2_X1 port map( A => n15137, B => n15136, ZN => n19823);
   U18484 : XNOR2_X1 port map( A => n15137, B => n15136, ZN => n1718);
   U18511 : XOR2_X1 port map( A => n13534, B => n19887, Z => n19824);
   U18519 : OR2_X1 port map( A1 => n20231, A2 => n20139, ZN => n19825);
   U18594 : XNOR2_X1 port map( A => n6524, B => n6523, ZN => n19826);
   U18718 : AOI21_X1 port map( B1 => n7792, B2 => n7791, A => n7790, ZN => 
                           n8985);
   U18741 : AOI21_X1 port map( B1 => n14538, B2 => n2676, A => n14537, ZN => 
                           n19828);
   U18757 : XOR2_X1 port map( A => n12990, B => n12989, Z => n19831);
   U18781 : XNOR2_X1 port map( A => n10184, B => n10183, ZN => n11431);
   U18849 : XOR2_X1 port map( A => n16065, B => n16064, Z => n19832);
   U18852 : NAND3_X1 port map( A1 => n11185, A2 => n2948, A3 => n2949, ZN => 
                           n19833);
   U19067 : NAND3_X1 port map( A1 => n2006, A2 => n3137, A3 => n3136, ZN => 
                           n17349);
   U19083 : BUF_X1 port map( A => n11132, Z => n19837);
   U19084 : OR2_X1 port map( A1 => n14278, A2 => n1409, ZN => n19838);
   U19122 : AOI22_X1 port map( A1 => n8643, A2 => n8929, B1 => n8598, B2 => 
                           n8933, ZN => n10179);
   U19144 : OAI211_X1 port map( C1 => n3603, C2 => n3604, A => n5814, B => 
                           n3602, ZN => n19840);
   U19145 : OAI211_X1 port map( C1 => n3603, C2 => n3604, A => n5814, B => 
                           n3602, ZN => n19841);
   U19147 : OAI21_X1 port map( B1 => n16317, B2 => n1112, A => n16316, ZN => 
                           n19842);
   U19148 : OAI211_X1 port map( C1 => n3603, C2 => n3604, A => n5814, B => 
                           n3602, ZN => n7231);
   U19149 : OAI21_X1 port map( B1 => n16317, B2 => n1112, A => n16316, ZN => 
                           n19196);
   U19150 : XNOR2_X1 port map( A => n10585, B => n10586, ZN => n11491);
   U19155 : NOR2_X1 port map( A1 => n14139, A2 => n14138, ZN => n19844);
   U19273 : NOR2_X1 port map( A1 => n14139, A2 => n14138, ZN => n19845);
   U19287 : XNOR2_X1 port map( A => n3419, B => n13654, ZN => n14722);
   U19290 : NOR2_X1 port map( A1 => n14139, A2 => n14138, ZN => n15936);
   U19360 : XOR2_X1 port map( A => n13446, B => n13644, Z => n12159);
   U19362 : XOR2_X1 port map( A => n16951, B => n16950, Z => n19846);
   U19464 : XOR2_X1 port map( A => n7122, B => n7081, Z => n19847);
   U19465 : XNOR2_X1 port map( A => n14963, B => n16969, ZN => n19849);
   U19466 : OAI21_X1 port map( B1 => n14505, B2 => n14506, A => n14504, ZN => 
                           n15284);
   U19573 : CLKBUF_X1 port map( A => n6754, Z => n19850);
   U19574 : XNOR2_X1 port map( A => n9425, B => n9424, ZN => n19851);
   U19575 : XNOR2_X1 port map( A => n9425, B => n9424, ZN => n11000);
   U19576 : XOR2_X1 port map( A => n7317, B => n7091, Z => n19852);
   U19577 : OAI211_X1 port map( C1 => n3494, C2 => n19941, A => n3495, B => 
                           n3492, ZN => n19853);
   U19578 : OAI211_X1 port map( C1 => n3494, C2 => n19941, A => n3495, B => 
                           n3492, ZN => n9669);
   U19582 : NAND3_X2 port map( A1 => n2847, A2 => n2850, A3 => n838, ZN => 
                           n10126);
   U19583 : XNOR2_X1 port map( A => n7293, B => n7292, ZN => n19856);
   U19586 : NOR2_X1 port map( A1 => n8512, A2 => n8513, ZN => n8510);
   U19587 : XOR2_X1 port map( A => n12732, B => n12733, Z => n19859);
   U19588 : BUF_X1 port map( A => n12636, Z => n19861);
   U19590 : OAI211_X2 port map( C1 => n9128, C2 => n9127, A => n9126, B => 
                           n9125, ZN => n10079);
   U19591 : XNOR2_X1 port map( A => n17359, B => n16429, ZN => n19863);
   U19592 : XNOR2_X1 port map( A => n10006, B => n10005, ZN => n19864);
   U19593 : XNOR2_X1 port map( A => n10006, B => n10005, ZN => n11514);
   U19594 : XNOR2_X1 port map( A => n5270, B => n5269, ZN => n19865);
   U19595 : XNOR2_X1 port map( A => n5270, B => n5269, ZN => n3748);
   U19596 : OAI21_X1 port map( B1 => n18952, B2 => n2590, A => n18951, ZN => 
                           n19866);
   U19597 : OAI21_X1 port map( B1 => n18952, B2 => n2590, A => n18951, ZN => 
                           n19867);
   U19598 : OAI21_X1 port map( B1 => n18952, B2 => n2590, A => n18951, ZN => 
                           n19021);
   U19599 : XOR2_X1 port map( A => Key(101), B => Plaintext(101), Z => n19868);
   U19600 : OAI211_X1 port map( C1 => n12235, C2 => n12236, A => n12234, B => 
                           n12233, ZN => n19869);
   U19602 : OAI211_X1 port map( C1 => n12235, C2 => n12236, A => n12234, B => 
                           n12233, ZN => n13511);
   U19603 : CLKBUF_X1 port map( A => n10299, Z => n19871);
   U19604 : XOR2_X1 port map( A => n1524, B => n1523, Z => n19872);
   U19606 : OAI21_X1 port map( B1 => n18962, B2 => n17057, A => n17056, ZN => 
                           n19874);
   U19607 : OAI21_X1 port map( B1 => n18962, B2 => n17057, A => n17056, ZN => 
                           n18899);
   U19608 : XNOR2_X1 port map( A => n11936, B => n11935, ZN => n14619);
   U19609 : OR2_X1 port map( A1 => n17551, A2 => n17550, ZN => n19877);
   U19610 : XNOR2_X1 port map( A => n17106, B => n17105, ZN => n17545);
   U19611 : XOR2_X1 port map( A => n9350, B => n9349, Z => n19878);
   U19612 : NOR2_X1 port map( A1 => n13318, A2 => n478, ZN => n19879);
   U19613 : OAI21_X1 port map( B1 => n7846, B2 => n20251, A => n1236, ZN => 
                           n19880);
   U19614 : OAI21_X1 port map( B1 => n7846, B2 => n20251, A => n1236, ZN => 
                           n9271);
   U19615 : XNOR2_X1 port map( A => n638, B => n6732, ZN => n19881);
   U19617 : OAI211_X1 port map( C1 => n13264, C2 => n14738, A => n13263, B => 
                           n1849, ZN => n19884);
   U19618 : AOI21_X1 port map( B1 => n12276, B2 => n12300, A => n1872, ZN => 
                           n12945);
   U19619 : OAI211_X1 port map( C1 => n13264, C2 => n14738, A => n13263, B => 
                           n1849, ZN => n15667);
   U19620 : XNOR2_X1 port map( A => n16340, B => n16339, ZN => n19885);
   U19621 : XNOR2_X1 port map( A => n16340, B => n16339, ZN => n18114);
   U19622 : XNOR2_X1 port map( A => n16758, B => n15827, ZN => n16673);
   U19623 : XOR2_X1 port map( A => n10285, B => n10284, Z => n19886);
   U19624 : OAI211_X1 port map( C1 => n12333, C2 => n11974, A => n11973, B => 
                           n11972, ZN => n19887);
   U19627 : CLKBUF_X1 port map( A => n18844, Z => n19890);
   U19628 : OAI21_X1 port map( B1 => n14567, B2 => n14566, A => n14565, ZN => 
                           n19891);
   U19630 : OAI21_X1 port map( B1 => n15765, B2 => n15248, A => n15247, ZN => 
                           n19894);
   U19631 : OAI211_X1 port map( C1 => n11807, C2 => n12537, A => n11806, B => 
                           n11805, ZN => n13519);
   U19633 : XNOR2_X1 port map( A => n10042, B => n10041, ZN => n19897);
   U19634 : OAI211_X1 port map( C1 => n7696, C2 => n7504, A => n7503, B => 
                           n7502, ZN => n8828);
   U19635 : XNOR2_X1 port map( A => n10042, B => n10041, ZN => n11211);
   U19636 : XNOR2_X1 port map( A => n15483, B => n15482, ZN => n19898);
   U19637 : XOR2_X1 port map( A => n13762, B => n13616, Z => n19899);
   U19639 : OAI211_X1 port map( C1 => n15208, C2 => n15207, A => n15206, B => 
                           n15205, ZN => n19900);
   U19640 : OAI211_X1 port map( C1 => n15208, C2 => n15207, A => n15206, B => 
                           n15205, ZN => n16747);
   U19641 : INV_X1 port map( A => n18497, ZN => n18489);
   U19642 : INV_X1 port map( A => n10726, ZN => n11093);
   U19643 : XNOR2_X1 port map( A => n6623, B => n6622, ZN => n19901);
   U19644 : XNOR2_X1 port map( A => n6623, B => n6622, ZN => n8175);
   U19645 : OAI21_X1 port map( B1 => n17713, B2 => n20221, A => n17712, ZN => 
                           n19043);
   U19646 : XNOR2_X1 port map( A => n13992, B => n16566, ZN => n19903);
   U19647 : OAI211_X1 port map( C1 => n12381, C2 => n12380, A => n12379, B => 
                           n12378, ZN => n19904);
   U19648 : CLKBUF_X1 port map( A => n17054, Z => n19905);
   U19649 : XNOR2_X1 port map( A => n2520, B => n2519, ZN => n19906);
   U19650 : XNOR2_X1 port map( A => n13766, B => n13765, ZN => n19907);
   U19651 : XNOR2_X1 port map( A => n13766, B => n13765, ZN => n19908);
   U19652 : OAI211_X1 port map( C1 => n15514, C2 => n15513, A => n15512, B => 
                           n519, ZN => n19909);
   U19653 : OAI211_X1 port map( C1 => n15514, C2 => n15513, A => n15512, B => 
                           n519, ZN => n16082);
   U19654 : XNOR2_X1 port map( A => n16033, B => n17371, ZN => n19910);
   U19656 : MUX2_X2 port map( A => n17011, B => n17010, S => n18932, Z => 
                           n18921);
   U19657 : INV_X1 port map( A => n12609, ZN => n19971);
   U19658 : OAI211_X1 port map( C1 => n3896, C2 => n4947, A => n3895, B => 
                           n3894, ZN => n19912);
   U19659 : XOR2_X1 port map( A => n10593, B => n10592, Z => n19913);
   U19660 : XOR2_X1 port map( A => n6878, B => n6877, Z => n19914);
   U19661 : XOR2_X1 port map( A => n8821, B => n8822, Z => n19915);
   U19662 : XNOR2_X1 port map( A => n16925, B => n16924, ZN => n19916);
   U19663 : OR2_X1 port map( A1 => n18050, A2 => n18049, ZN => n19917);
   U19664 : XNOR2_X1 port map( A => n13821, B => n13822, ZN => n19918);
   U19665 : XOR2_X1 port map( A => n17266, B => n17265, Z => n19919);
   U19666 : XNOR2_X1 port map( A => n13821, B => n13822, ZN => n14250);
   U19667 : XNOR2_X1 port map( A => n10429, B => n10428, ZN => n19920);
   U19668 : BUF_X1 port map( A => n14692, Z => n19921);
   U19669 : XNOR2_X1 port map( A => n10429, B => n10428, ZN => n11443);
   U19670 : XNOR2_X1 port map( A => n5727, B => n5726, ZN => n19922);
   U19671 : NOR2_X1 port map( A1 => n12190, A2 => n2426, ZN => n19923);
   U19672 : NOR2_X1 port map( A1 => n12190, A2 => n2426, ZN => n13383);
   U19673 : XOR2_X1 port map( A => n15483, B => n15482, Z => n19924);
   U19674 : XNOR2_X1 port map( A => n2211, B => n6772, ZN => n19925);
   U19676 : NOR2_X1 port map( A1 => n14862, A2 => n1489, ZN => n19927);
   U19677 : NOR2_X1 port map( A1 => n14862, A2 => n1489, ZN => n19928);
   U19678 : NOR2_X1 port map( A1 => n14862, A2 => n1489, ZN => n17425);
   U19680 : XNOR2_X1 port map( A => n16049, B => n16048, ZN => n19930);
   U19681 : XNOR2_X1 port map( A => n16049, B => n16048, ZN => n17666);
   U19682 : OAI21_X1 port map( B1 => n14578, B2 => n20187, A => n14577, ZN => 
                           n19931);
   U19683 : OAI21_X1 port map( B1 => n14578, B2 => n20187, A => n14577, ZN => 
                           n15828);
   U19685 : XOR2_X1 port map( A => n16935, B => n16934, Z => n19933);
   U19686 : INV_X1 port map( A => n18652, ZN => n19935);
   U19687 : OAI21_X1 port map( B1 => n18142, B2 => n18141, A => n18140, ZN => 
                           n18652);
   U19688 : XOR2_X1 port map( A => n16532, B => n16531, Z => n19936);
   U19689 : OAI211_X1 port map( C1 => n12428, C2 => n3649, A => n12098, B => 
                           n12097, ZN => n19937);
   U19690 : XNOR2_X1 port map( A => n1436, B => n16509, ZN => n19938);
   U19691 : XOR2_X1 port map( A => n13046, B => n13045, Z => n19940);
   U19692 : OAI211_X1 port map( C1 => n7682, C2 => n8166, A => n7681, B => 
                           n7680, ZN => n9354);
   U19694 : XOR2_X1 port map( A => n16352, B => n16351, Z => n19943);
   U19695 : OAI211_X1 port map( C1 => n5225, C2 => n5768, A => n5224, B => 
                           n5223, ZN => n19944);
   U19696 : OAI211_X1 port map( C1 => n5225, C2 => n5768, A => n5224, B => 
                           n5223, ZN => n7187);
   U19697 : AOI21_X1 port map( B1 => n9133, B2 => n9132, A => n9131, ZN => 
                           n10077);
   U19698 : AOI21_X1 port map( B1 => n12297, B2 => n12296, A => n2220, ZN => 
                           n19946);
   U19699 : XNOR2_X1 port map( A => n16087, B => n16086, ZN => n19947);
   U19700 : XNOR2_X1 port map( A => n16087, B => n16086, ZN => n17887);
   U19701 : MUX2_X1 port map( A => n17083, B => n17082, S => n20239, Z => 
                           n19948);
   U19702 : MUX2_X1 port map( A => n17083, B => n17082, S => n20239, Z => 
                           n19164);
   U19708 : XNOR2_X2 port map( A => n13326, B => n13327, ZN => n14385);
   U19709 : AOI22_X1 port map( A1 => n6160, A2 => n5614, B1 => n5613, B2 => 
                           n5612, ZN => n19953);
   U19711 : NAND2_X1 port map( A1 => n565, A2 => n1154, ZN => n19954);
   U19712 : OAI21_X1 port map( B1 => n20240, B2 => n16543, A => n16542, ZN => 
                           n19955);
   U19714 : XNOR2_X1 port map( A => n3575, B => n3574, ZN => n19956);
   U19715 : XNOR2_X1 port map( A => n3575, B => n3574, ZN => n17223);
   U19716 : XOR2_X1 port map( A => n9096, B => n9097, Z => n19957);
   U19717 : OR2_X1 port map( A1 => n11349, A2 => n11347, ZN => n11060);
   U19719 : XOR2_X1 port map( A => n10408, B => n10407, Z => n19959);
   U19720 : NAND2_X1 port map( A1 => n9308, A2 => n9313, ZN => n1128);
   U19721 : AND2_X2 port map( A1 => n19960, A2 => n19529, ZN => n9313);
   U19722 : NAND2_X1 port map( A1 => n1584, A2 => n8113, ZN => n19960);
   U19723 : NAND2_X1 port map( A1 => n19962, A2 => n18042, ZN => n17814);
   U19724 : NOR2_X1 port map( A1 => n18948, A2 => n17812, ZN => n19962);
   U19725 : NAND2_X1 port map( A1 => n19963, A2 => n4330, ZN => n3110);
   U19726 : NAND2_X1 port map( A1 => n4177, A2 => n4613, ZN => n4330);
   U19727 : OAI21_X2 port map( B1 => n15548, B2 => n2803, A => n1100, ZN => 
                           n16872);
   U19728 : NOR3_X1 port map( A1 => n11953, A2 => n11829, A3 => n11952, ZN => 
                           n2562);
   U19729 : NAND4_X1 port map( A1 => n11822, A2 => n19964, A3 => n11821, A4 => 
                           n13270, ZN => n11823);
   U19730 : NAND2_X1 port map( A1 => n12325, A2 => n11997, ZN => n19964);
   U19732 : NAND2_X1 port map( A1 => n15802, A2 => n15801, ZN => n19966);
   U19733 : NAND2_X1 port map( A1 => n5840, A2 => n19967, ZN => n7143);
   U19734 : NAND2_X1 port map( A1 => n19522, A2 => n19968, ZN => n19967);
   U19735 : NAND2_X1 port map( A1 => n1293, A2 => n15402, ZN => n15069);
   U19736 : XNOR2_X1 port map( A => n19969, B => n18389, ZN => Ciphertext(9));
   U19737 : OAI21_X1 port map( B1 => n12610, B2 => n19971, A => n19970, ZN => 
                           n12239);
   U19738 : NAND2_X1 port map( A1 => n12610, A2 => n12237, ZN => n19970);
   U19740 : NAND2_X1 port map( A1 => n7980, A2 => n7767, ZN => n7769);
   U19741 : NAND2_X1 port map( A1 => n19517, A2 => n7752, ZN => n3554);
   U19742 : NAND2_X1 port map( A1 => n15108, A2 => n14947, ZN => n16329);
   U19743 : NAND2_X1 port map( A1 => n14944, A2 => n15292, ZN => n14946);
   U19746 : OR2_X1 port map( A1 => n11289, A2 => n9559, ZN => n19972);
   U19747 : XNOR2_X1 port map( A => n13261, B => n13262, ZN => n14736);
   U19748 : OAI211_X1 port map( C1 => n12333, C2 => n11974, A => n11973, B => 
                           n11972, ZN => n12997);
   U1521 : AND3_X2 port map( A1 => n11994, A2 => n11993, A3 => n12333, ZN => 
                           n13481);
   U1416 : BUF_X1 port map( A => n16011, Z => n901);
   U915 : NAND2_X2 port map( A1 => n14118, A2 => n14117, ZN => n16126);
   U2647 : XNOR2_X2 port map( A => n6561, B => n6560, ZN => n8100);
   U891 : MUX2_X2 port map( A => n14075, B => n14074, S => n3223, Z => n15748);
   U2961 : AND2_X2 port map( A1 => n13182, A2 => n13181, ZN => n785);
   U14440 : BUF_X2 port map( A => n12061, Z => n12595);
   U17527 : INV_X1 port map( A => n17650, ZN => n19401);
   U1744 : NAND2_X2 port map( A1 => n3750, A2 => n970, ZN => n9105);
   U8534 : BUF_X2 port map( A => n7457, Z => n8196);
   U1619 : BUF_X1 port map( A => n11147, Z => n11016);
   U1315 : BUF_X1 port map( A => n15310, Z => n19662);
   U6746 : OAI21_X2 port map( B1 => n7869, B2 => n7870, A => n7868, ZN => 
                           n10264);
   U555 : XNOR2_X1 port map( A => n9690, B => n9689, ZN => n11377);
   U1092 : OAI22_X2 port map( A1 => n9933, A2 => n10635, B1 => n10923, B2 => 
                           n2469, ZN => n12352);
   U6737 : OAI211_X2 port map( C1 => n5373, C2 => n5398, A => n5372, B => n5371
                           , ZN => n7316);
   U2601 : XNOR2_X1 port map( A => n5940, B => n5939, ZN => n8300);
   U1915 : NAND2_X2 port map( A1 => n3350, A2 => n3349, ZN => n6050);
   U15140 : INV_X1 port map( A => n19336, ZN => n19337);
   U848 : NAND3_X2 port map( A1 => n2898, A2 => n2899, A3 => n2897, ZN => n3305
                           );
   U8972 : BUF_X1 port map( A => n16982, Z => n19674);
   U224 : BUF_X1 port map( A => n8195, Z => n19474);
   U4696 : OR3_X1 port map( A1 => n8652, A2 => n9262, A3 => n7866, ZN => n8655)
                           ;
   U6176 : NOR2_X2 port map( A1 => n3213, A2 => n3215, ZN => n19190);
   U19584 : NOR2_X2 port map( A1 => n8512, A2 => n8513, ZN => n19857);
   U8825 : XNOR2_X1 port map( A => Key(144), B => Plaintext(144), ZN => n4750);
   U1247 : CLKBUF_X1 port map( A => Key(175), Z => n2100);
   U8855 : XNOR2_X1 port map( A => Key(165), B => Plaintext(165), ZN => n3948);
   U9023 : XNOR2_X1 port map( A => n4045, B => Key(106), ZN => n5101);
   U6816 : AND2_X1 port map( A1 => n4351, A2 => n4352, ZN => n5717);
   U1935 : AND3_X1 port map( A1 => n5505, A2 => n5504, A3 => n5510, ZN => n6007
                           );
   U73 : OAI211_X1 port map( C1 => n4608, C2 => n4607, A => n4606, B => n4605, 
                           ZN => n5745);
   U5550 : AND2_X1 port map( A1 => n4579, A2 => n4580, ZN => n5382);
   U554 : NAND2_X1 port map( A1 => n4267, A2 => n4266, ZN => n6129);
   U6032 : AND3_X1 port map( A1 => n3008, A2 => n3009, A3 => n4735, ZN => n6113
                           );
   U1901 : AND2_X1 port map( A1 => n4918, A2 => n4917, ZN => n5476);
   U56 : AND2_X1 port map( A1 => n3640, A2 => n5226, ZN => n6220);
   U9641 : OR2_X1 port map( A1 => n4995, A2 => n5138, ZN => n4997);
   U897 : NAND2_X1 port map( A1 => n5123, A2 => n1978, ZN => n7046);
   U924 : NAND2_X1 port map( A1 => n1708, A2 => n1705, ZN => n7392);
   U439 : OAI211_X1 port map( C1 => n5275, C2 => n19562, A => n5274, B => n5273
                           , ZN => n6850);
   U4748 : NAND2_X1 port map( A1 => n1886, A2 => n1885, ZN => n7267);
   U10333 : OAI211_X1 port map( C1 => n6160, C2 => n6159, A => n6158, B => 
                           n6157, ZN => n7348);
   U470 : BUF_X1 port map( A => n5984, Z => n7272);
   U941 : BUF_X1 port map( A => n7009, Z => n179);
   U10260 : XNOR2_X1 port map( A => n5962, B => n5961, ZN => n8299);
   U11101 : XNOR2_X1 port map( A => n7029, B => n7030, ZN => n7836);
   U692 : BUF_X1 port map( A => n6510, Z => n7560);
   U547 : NAND2_X1 port map( A1 => n7498, A2 => n3377, ZN => n9291);
   U4861 : INV_X1 port map( A => n8722, ZN => n9358);
   U1737 : OR2_X1 port map( A1 => n8223, A2 => n8224, ZN => n8797);
   U7666 : AND2_X1 port map( A1 => n3075, A2 => n3073, ZN => n9031);
   U7995 : NAND2_X1 port map( A1 => n3384, A2 => n3383, ZN => n8527);
   U1470 : INV_X1 port map( A => n8419, ZN => n9209);
   U5581 : AND2_X1 port map( A1 => n7804, A2 => n7803, ZN => n8987);
   U914 : OAI211_X1 port map( C1 => n8611, C2 => n7540, A => n7539, B => n7538,
                           ZN => n9947);
   U6707 : OAI21_X1 port map( B1 => n8496, B2 => n8495, A => n8494, ZN => n9817
                           );
   U3538 : NAND2_X1 port map( A1 => n8519, A2 => n8518, ZN => n10461);
   U4864 : NAND2_X1 port map( A1 => n1202, A2 => n1200, ZN => n10436);
   U1671 : AND3_X1 port map( A1 => n8626, A2 => n8625, A3 => n8624, ZN => 
                           n10002);
   U3871 : AND2_X1 port map( A1 => n9323, A2 => n9838, ZN => n9960);
   U859 : XNOR2_X1 port map( A => n9823, B => n9822, ZN => n11263);
   U1633 : XNOR2_X1 port map( A => n1823, B => n9316, ZN => n11177);
   U3241 : XNOR2_X1 port map( A => n2496, B => n2495, ZN => n11192);
   U7367 : XNOR2_X1 port map( A => n8590, B => n8591, ZN => n10926);
   U1642 : XNOR2_X1 port map( A => n10147, B => n10146, ZN => n11057);
   U592 : XNOR2_X1 port map( A => n9929, B => n9928, ZN => n11076);
   U179 : INV_X1 port map( A => n10513, ZN => n11440);
   U731 : BUF_X1 port map( A => n10112, Z => n10813);
   U13717 : NAND3_X1 port map( A1 => n202, A2 => n2861, A3 => n11376, ZN => 
                           n10858);
   U13393 : INV_X1 port map( A => n10724, ZN => n11051);
   U3259 : OR2_X1 port map( A1 => n9546, A2 => n9547, ZN => n3176);
   U1572 : OR2_X1 port map( A1 => n9490, A2 => n9489, ZN => n9491);
   U1557 : INV_X1 port map( A => n9491, ZN => n12179);
   U13621 : MUX2_X1 port map( A => n10744, B => n10743, S => n10936, Z => 
                           n12754);
   U827 : OAI21_X1 port map( B1 => n10648, B2 => n11556, A => n10647, ZN => 
                           n12421);
   U3938 : OAI211_X1 port map( C1 => n11050, C2 => n11459, A => n2130, B => 
                           n10260, ZN => n12339);
   U2295 : OR2_X1 port map( A1 => n12590, A2 => n12200, ZN => n1252);
   U3413 : NOR2_X1 port map( A1 => n10659, A2 => n10658, ZN => n13088);
   U14164 : MUX2_X1 port map( A => n11663, B => n11662, S => n11661, Z => 
                           n13651);
   U614 : AOI22_X1 port map( A1 => n13144, A2 => n13146, B1 => n11099, B2 => 
                           n11098, ZN => n13280);
   U129 : AND3_X1 port map( A1 => n1981, A2 => n10850, A3 => n1980, ZN => 
                           n12709);
   U4719 : NAND3_X1 port map( A1 => n12112, A2 => n12113, A3 => n12111, ZN => 
                           n13398);
   U763 : AND2_X1 port map( A1 => n12447, A2 => n12446, ZN => n13697);
   U266 : NAND2_X1 port map( A1 => n11919, A2 => n40, ZN => n13453);
   U3615 : INV_X1 port map( A => n14249, ZN => n1262);
   U1468 : XNOR2_X1 port map( A => n13663, B => n13662, ZN => n14717);
   U14960 : XNOR2_X1 port map( A => n12858, B => n12857, ZN => n14451);
   U124 : BUF_X1 port map( A => n14420, Z => n19939);
   U909 : XNOR2_X1 port map( A => n11103, B => n11102, ZN => n14780);
   U946 : XNOR2_X1 port map( A => n12943, B => n12942, ZN => n14644);
   U6806 : MUX2_X1 port map( A => n13630, B => n13629, S => n19731, Z => n15682
                           );
   U15881 : MUX2_X2 port map( A => n14110, B => n14109, S => n14723, Z => 
                           n15495);
   U995 : NAND2_X1 port map( A1 => n13949, A2 => n2952, ZN => n16016);
   U15063 : NAND2_X1 port map( A1 => n12975, A2 => n12976, ZN => n15777);
   U164 : NOR2_X1 port map( A1 => n14756, A2 => n14755, ZN => n15503);
   U959 : BUF_X1 port map( A => n15515, Z => n19502);
   U397 : AND2_X1 port map( A1 => n14616, A2 => n14615, ZN => n15276);
   U1063 : OR2_X1 port map( A1 => n15567, A2 => n15566, ZN => n14954);
   U5473 : AND2_X1 port map( A1 => n2564, A2 => n2565, ZN => n15870);
   U544 : XNOR2_X1 port map( A => n15889, B => n15888, ZN => n19352);
   U1336 : CLKBUF_X1 port map( A => n18026, Z => n17749);
   U17439 : INV_X1 port map( A => n17955, ZN => n18107);
   U18695 : MUX2_X1 port map( A => n18045, B => n18044, S => n18946, Z => 
                           n18050);
   U843 : OAI211_X1 port map( C1 => n2819, C2 => n17664, A => n2818, B => n2817
                           , ZN => n2816);
   U5765 : AOI22_X1 port map( A1 => n17614, A2 => n17613, B1 => n17612, B2 => 
                           n17611, ZN => n19299);
   U8402 : OAI21_X1 port map( B1 => n16913, B2 => n16912, A => n16911, ZN => 
                           n18897);
   U196 : AND3_X1 port map( A1 => n18247, A2 => n18246, A3 => n18245, ZN => 
                           n18773);
   U2062 : NAND2_X1 port map( A1 => n17747, A2 => n319, ZN => n18807);
   U2093 : OAI211_X1 port map( C1 => n20648, C2 => n16797, A => n2633, B => 
                           n16168, ZN => n18497);
   U1039 : OR2_X1 port map( A1 => n15965, A2 => n15964, ZN => n18057);
   U650 : OR2_X1 port map( A1 => n20124, A2 => n19233, ZN => n19229);
   U9292 : INV_X1 port map( A => n5717, ZN => n5714);
   U1015 : INV_X1 port map( A => n5349, ZN => n6156);
   U3720 : CLKBUF_X1 port map( A => n3855, Z => n5785);
   U161 : NAND2_X2 port map( A1 => n3658, A2 => n1807, ZN => n5605);
   U5895 : MUX2_X1 port map( A => n5890, B => n5889, S => n5888, Z => n6761);
   U431 : OAI211_X1 port map( C1 => n5654, C2 => n5653, A => n5652, B => n5651,
                           ZN => n6912);
   U3791 : INV_X1 port map( A => n7470, ZN => n8293);
   U1686 : AND2_X1 port map( A1 => n1103, A2 => n1102, ZN => n9414);
   U6090 : XNOR2_X1 port map( A => n9156, B => n9155, ZN => n11556);
   U3911 : INV_X1 port map( A => n9351, ZN => n11178);
   U1495 : NAND2_X1 port map( A1 => n3277, A2 => n3276, ZN => n13572);
   U2594 : NAND3_X1 port map( A1 => n11861, A2 => n542, A3 => n541, ZN => 
                           n13064);
   U2700 : OR2_X1 port map( A1 => n14022, A2 => n14021, ZN => n14288);
   U1071 : BUF_X1 port map( A => n13946, Z => n14688);
   U6010 : OAI211_X1 port map( C1 => n12695, C2 => n14419, A => n3635, B => 
                           n3636, ZN => n15341);
   U550 : AOI22_X1 port map( A1 => n15605, A2 => n15604, B1 => n15603, B2 => 
                           n15602, ZN => n16970);
   U38 : MUX2_X1 port map( A => n16315, B => n16314, S => n20512, Z => n16316);
   U11616 : CLKBUF_X1 port map( A => n18009, Z => n18522);
   U1136 : MUX2_X2 port map( A => n4661, B => n4660, S => n4841, Z => n6168);
   U289 : NAND3_X2 port map( A1 => n7435, A2 => n7434, A3 => n7433, ZN => n9295
                           );
   U4569 : NOR2_X2 port map( A1 => n14331, A2 => n14330, ZN => n15470);
   U5326 : AND2_X2 port map( A1 => n3594, A2 => n3595, ZN => n9204);
   U5119 : NOR2_X2 port map( A1 => n11669, A2 => n11668, ZN => n12940);
   U1750 : BUF_X2 port map( A => n8103, Z => n9328);
   U12894 : XNOR2_X2 port map( A => n10503, B => n9770, ZN => n11866);
   U777 : AND3_X2 port map( A1 => n822, A2 => n3585, A3 => n3584, ZN => n953);
   U141 : NOR2_X2 port map( A1 => n6188, A2 => n6187, ZN => n19778);
   U2761 : AOI22_X2 port map( A1 => n15039, A2 => n15698, B1 => n15702, B2 => 
                           n15040, ZN => n17143);
   U255 : NAND3_X2 port map( A1 => n6179, A2 => n6177, A3 => n6178, ZN => n7032
                           );
   U6882 : MUX2_X2 port map( A => n6086, B => n6085, S => n3529, Z => n7354);
   U10348 : MUX2_X2 port map( A => n8554, B => n8553, S => n8814, Z => n10421);
   U2639 : NAND2_X2 port map( A1 => n3135, A2 => n3296, ZN => n12686);
   U753 : OR2_X2 port map( A1 => n8246, A2 => n8253, ZN => n900);
   U657 : AND2_X2 port map( A1 => n14816, A2 => n14815, ZN => n15813);
   U1289 : BUF_X1 port map( A => n18667, Z => n18666);
   U11221 : XNOR2_X2 port map( A => n7200, B => n7199, ZN => n8313);
   U559 : OR2_X2 port map( A1 => n104, A2 => n11450, ZN => n12523);
   U472 : AND2_X2 port map( A1 => n2077, A2 => n2076, ZN => n5401);
   U4538 : MUX2_X1 port map( A => n5561, B => n5560, S => n5559, Z => n7080);
   U892 : BUF_X2 port map( A => n7568, Z => n7864);
   U1510 : AOI22_X1 port map( A1 => n12064, A2 => n12063, B1 => n12201, B2 => 
                           n12062, ZN => n13027);
   U841 : BUF_X2 port map( A => n14425, Z => n14424);
   U26 : AOI21_X1 port map( B1 => n8692, B2 => n8691, A => n8690, ZN => n12349)
                           ;
   U31 : OAI22_X1 port map( A1 => n3220, A2 => n3221, B1 => n7311, B2 => n7343,
                           ZN => n8928);
   U75 : BUF_X1 port map( A => n13468, Z => n13818);
   U84 : BUF_X1 port map( A => n10179, Z => n19839);
   U97 : BUF_X1 port map( A => n14829, Z => n19986);
   U105 : BUF_X1 port map( A => n18858, Z => n19989);
   U112 : XNOR2_X1 port map( A => n2991, B => n2992, ZN => n17831);
   U122 : NAND2_X1 port map( A1 => n16467, A2 => n60, ZN => n18453);
   U127 : OR2_X2 port map( A1 => n3791, A2 => n3794, ZN => n8846);
   U136 : NOR2_X2 port map( A1 => n11128, A2 => n2029, ZN => n12382);
   U142 : OAI21_X2 port map( B1 => n10878, B2 => n10879, A => n10877, ZN => 
                           n19854);
   U165 : XNOR2_X2 port map( A => n13007, B => n13006, ZN => n14648);
   U167 : AOI21_X2 port map( B1 => n10888, B2 => n10887, A => n10886, ZN => 
                           n12609);
   U185 : NAND2_X2 port map( A1 => n13915, A2 => n3222, ZN => n15864);
   U197 : OAI211_X2 port map( C1 => n14093, C2 => n14094, A => n12802, B => 
                           n12801, ZN => n15469);
   U203 : XOR2_X1 port map( A => n15969, B => n15968, Z => n19973);
   U217 : XOR2_X1 port map( A => n14942, B => n14943, Z => n19975);
   U259 : MUX2_X2 port map( A => n8009, B => n8008, S => n8314, Z => n8831);
   U306 : XNOR2_X2 port map( A => n17285, B => n17284, ZN => n18238);
   U309 : AOI21_X2 port map( B1 => n13990, B2 => n13991, A => n15303, ZN => 
                           n16566);
   U340 : NAND3_X2 port map( A1 => n14212, A2 => n14211, A3 => n3274, ZN => 
                           n15618);
   U353 : AND3_X2 port map( A1 => n2823, A2 => n16265, A3 => n2822, ZN => 
                           n19209);
   U373 : NAND3_X2 port map( A1 => n1095, A2 => n5287, A3 => n5288, ZN => n7266
                           );
   U382 : BUF_X1 port map( A => n5589, Z => n19980);
   U388 : OAI211_X1 port map( C1 => n5091, C2 => n5090, A => n1360, B => n5089,
                           ZN => n5589);
   U395 : BUF_X2 port map( A => n12800, Z => n19485);
   U418 : XNOR2_X2 port map( A => n16208, B => n16207, ZN => n17564);
   U423 : XNOR2_X2 port map( A => n12753, B => n12752, ZN => n14828);
   U425 : NAND4_X2 port map( A1 => n15786, A2 => n15785, A3 => n15787, A4 => 
                           n15784, ZN => n16278);
   U427 : NOR2_X2 port map( A1 => n15623, A2 => n15624, ZN => n16960);
   U428 : NAND3_X2 port map( A1 => n5994, A2 => n5993, A3 => n5992, ZN => n7050
                           );
   U456 : XNOR2_X2 port map( A => n12319, B => n12318, ZN => n14796);
   U468 : NAND3_X2 port map( A1 => n2346, A2 => n11017, A3 => n2345, ZN => 
                           n13767);
   U491 : XNOR2_X1 port map( A => n13214, B => n13213, ZN => n14022);
   U508 : NAND2_X2 port map( A1 => n1380, A2 => n3707, ZN => n13048);
   U509 : AND3_X2 port map( A1 => n6847, A2 => n6846, A3 => n6845, ZN => n9307)
                           ;
   U514 : AND2_X2 port map( A1 => n20342, A2 => n20341, ZN => n17355);
   U521 : XNOR2_X2 port map( A => n17009, B => n17008, ZN => n18928);
   U522 : NAND3_X2 port map( A1 => n12220, A2 => n3360, A3 => n3359, ZN => 
                           n12230);
   U541 : MUX2_X2 port map( A => n5427, B => n5426, S => n5668, Z => n7116);
   U545 : NAND3_X2 port map( A1 => n9237, A2 => n3060, A3 => n3059, ZN => 
                           n10484);
   U549 : BUF_X2 port map( A => n16320, Z => n17471);
   U576 : OAI21_X2 port map( B1 => n10692, B2 => n19851, A => n10691, ZN => 
                           n12631);
   U584 : NAND2_X2 port map( A1 => n19608, A2 => n19607, ZN => n15741);
   U585 : OR2_X1 port map( A1 => n8301, A2 => n2792, ZN => n8047);
   U586 : XNOR2_X2 port map( A => n5214, B => n5213, ZN => n8301);
   U626 : XNOR2_X2 port map( A => n16536, B => n16537, ZN => n19360);
   U627 : OAI21_X2 port map( B1 => n13094, B2 => n15120, A => n13093, ZN => 
                           n15686);
   U628 : INV_X1 port map( A => n9017, ZN => n19564);
   U641 : XNOR2_X2 port map( A => n3947, B => Key(180), ZN => n4548);
   U647 : NOR2_X2 port map( A1 => n16631, A2 => n16630, ZN => n18365);
   U656 : XNOR2_X2 port map( A => n8719, B => n8718, ZN => n11168);
   U677 : NOR2_X2 port map( A1 => n5731, A2 => n1476, ZN => n6743);
   U700 : BUF_X1 port map( A => n11191, Z => n19983);
   U707 : XNOR2_X1 port map( A => n10547, B => n10546, ZN => n11191);
   U721 : NOR2_X2 port map( A1 => n8666, A2 => n9781, ZN => n10595);
   U723 : OAI21_X2 port map( B1 => n2988, B2 => n15170, A => n13993, ZN => 
                           n16926);
   U725 : NAND2_X2 port map( A1 => n5982, A2 => n5981, ZN => n7047);
   U737 : OAI21_X2 port map( B1 => n8110, B2 => n8151, A => n8109, ZN => n9330)
                           ;
   U743 : BUF_X1 port map( A => n14829, Z => n19985);
   U757 : XNOR2_X1 port map( A => n12739, B => n12738, ZN => n14829);
   U764 : XNOR2_X2 port map( A => n3858, B => Key(91), ZN => n4405);
   U775 : OR2_X2 port map( A1 => n5503, A2 => n5508, ZN => n5914);
   U778 : NAND2_X2 port map( A1 => n15415, A2 => n15414, ZN => n17133);
   U809 : AND3_X2 port map( A1 => n2249, A2 => n3443, A3 => n3442, ZN => n15636
                           );
   U823 : OAI21_X2 port map( B1 => n12076, B2 => n12075, A => n3269, ZN => 
                           n13659);
   U824 : AND3_X2 port map( A1 => n1619, A2 => n1621, A3 => n1622, ZN => n6966)
                           ;
   U837 : BUF_X1 port map( A => n18858, Z => n19988);
   U850 : OAI211_X1 port map( C1 => n18023, C2 => n18936, A => n18022, B => 
                           n18021, ZN => n18858);
   U866 : XNOR2_X2 port map( A => n7398, B => n7399, ZN => n8026);
   U880 : OAI21_X2 port map( B1 => n745, B2 => n9578, A => n744, ZN => n10261);
   U887 : OAI21_X2 port map( B1 => n5912, B2 => n4876, A => n4875, ZN => n7184)
                           ;
   U899 : OAI21_X2 port map( B1 => n7859, B2 => n7556, A => n6550, ZN => n9241)
                           ;
   U902 : BUF_X2 port map( A => n11129, Z => n11418);
   U912 : OAI21_X2 port map( B1 => n4958, B2 => n4959, A => n20339, ZN => n5569
                           );
   U922 : OAI211_X2 port map( C1 => n11977, C2 => n11800, A => n11799, B => 
                           n11798, ZN => n13810);
   U923 : OAI22_X2 port map( A1 => n1268, A2 => n1267, B1 => n7654, B2 => n7653
                           , ZN => n10456);
   U926 : NAND3_X2 port map( A1 => n2054, A2 => n12058, A3 => n2052, ZN => 
                           n13658);
   U929 : NOR2_X2 port map( A1 => n3670, A2 => n11146, ZN => n12281);
   U939 : BUF_X1 port map( A => n19040, Z => n19992);
   U940 : CLKBUF_X1 port map( A => n19040, Z => n19993);
   U942 : NOR2_X1 port map( A1 => n17698, A2 => n17697, ZN => n19040);
   U945 : OAI211_X2 port map( C1 => n9226, C2 => n9053, A => n1759, B => n9227,
                           ZN => n10087);
   U947 : XNOR2_X2 port map( A => n6628, B => n6629, ZN => n8178);
   U948 : XNOR2_X2 port map( A => n6310, B => n6311, ZN => n7984);
   U966 : NOR2_X2 port map( A1 => n3502, A2 => n3501, ZN => n10296);
   U972 : NOR2_X2 port map( A1 => n1175, A2 => n9791, ZN => n12508);
   U974 : OAI21_X2 port map( B1 => n11983, B2 => n11635, A => n11634, ZN => 
                           n13734);
   U988 : XNOR2_X2 port map( A => Key(86), B => Plaintext(86), ZN => n4410);
   U998 : OAI211_X2 port map( C1 => n18128, C2 => n18129, A => n17780, B => 
                           n17779, ZN => n18803);
   U999 : XNOR2_X2 port map( A => n547, B => Key(188), ZN => n4365);
   U1056 : XNOR2_X2 port map( A => Key(163), B => Plaintext(163), ZN => n4350);
   U1070 : OAI21_X2 port map( B1 => n5003, B2 => n4253, A => n99, ZN => n6133);
   U1089 : AOI21_X2 port map( B1 => n11895, B2 => n11894, A => n11893, ZN => 
                           n13422);
   U1110 : OR2_X1 port map( A1 => n18847, A2 => n3028, ZN => n20041);
   U1114 : BUF_X1 port map( A => n18454, Z => n18466);
   U1118 : INV_X1 port map( A => n15529, ZN => n19997);
   U1145 : NAND2_X1 port map( A1 => n16472, A2 => n16473, ZN => n18465);
   U1234 : XNOR2_X1 port map( A => n3093, B => n3090, ZN => n16306);
   U1266 : XNOR2_X1 port map( A => n16069, B => n16068, ZN => n17881);
   U1279 : OR2_X1 port map( A1 => n12930, A2 => n12929, ZN => n231);
   U1295 : OAI211_X1 port map( C1 => n922, C2 => n11946, A => n10792, B => 
                           n10791, ZN => n13336);
   U1296 : INV_X1 port map( A => n11192, ZN => n19998);
   U1301 : INV_X1 port map( A => n11526, ZN => n19999);
   U1303 : INV_X1 port map( A => n1449, ZN => n20000);
   U1304 : BUF_X1 port map( A => n9310, Z => n20011);
   U1327 : INV_X1 port map( A => n8100, ZN => n8112);
   U1333 : INV_X1 port map( A => n3748, ZN => n20001);
   U1347 : INV_X1 port map( A => n5081, ZN => n20002);
   U1353 : CLKBUF_X1 port map( A => Key(57), Z => n18177);
   U1368 : CLKBUF_X1 port map( A => Key(185), Z => n645);
   U1384 : OR2_X1 port map( A1 => n19130, A2 => n19125, ZN => n3142);
   U1410 : OAI21_X1 port map( B1 => n17499, B2 => n16480, A => n16479, ZN => 
                           n18464);
   U1423 : OR2_X1 port map( A1 => n18157, A2 => n18057, ZN => n18158);
   U1426 : BUF_X2 port map( A => n18652, Z => n19934);
   U1451 : OAI21_X1 port map( B1 => n17385, B2 => n17384, A => n17383, ZN => 
                           n20276);
   U1455 : AND2_X1 port map( A1 => n17319, A2 => n17318, ZN => n18172);
   U1488 : INV_X1 port map( A => n18400, ZN => n20003);
   U1518 : OR2_X1 port map( A1 => n16543, A2 => n20240, ZN => n20065);
   U1525 : OAI211_X1 port map( C1 => n16677, C2 => n16676, A => n16675, B => 
                           n2206, ZN => n20152);
   U1606 : XNOR2_X1 port map( A => n16774, B => n16773, ZN => n20221);
   U1624 : XNOR2_X1 port map( A => n17018, B => n17017, ZN => n18938);
   U1630 : XNOR2_X1 port map( A => n17405, B => n17404, ZN => n18130);
   U1639 : INV_X1 port map( A => n19389, ZN => n20004);
   U1648 : NAND3_X1 port map( A1 => n20022, A2 => n1757, A3 => n1610, ZN => 
                           n16562);
   U1691 : INV_X1 port map( A => n15696, ZN => n20005);
   U1724 : INV_X1 port map( A => n231, ZN => n15166);
   U1725 : INV_X1 port map( A => n15898, ZN => n20006);
   U1738 : INV_X1 port map( A => n16128, ZN => n20007);
   U1762 : NAND2_X1 port map( A1 => n20284, A2 => n20283, ZN => n15657);
   U1798 : CLKBUF_X1 port map( A => n11717, Z => n20215);
   U1804 : NAND2_X1 port map( A1 => n8903, A2 => n3279, ZN => n12002);
   U1805 : NAND2_X1 port map( A1 => n11280, A2 => n11279, ZN => n12488);
   U1822 : INV_X1 port map( A => n3667, ZN => n20297);
   U1874 : NAND3_X1 port map( A1 => n1750, A2 => n529, A3 => n1753, ZN => 
                           n10274);
   U1900 : OR2_X1 port map( A1 => n9188, A2 => n268, ZN => n2014);
   U1916 : INV_X1 port map( A => n9328, ZN => n20008);
   U1978 : INV_X1 port map( A => n8276, ZN => n20009);
   U2047 : OR2_X1 port map( A1 => n7898, A2 => n2703, ZN => n20315);
   U2065 : OR2_X1 port map( A1 => n8083, A2 => n20107, ZN => n20086);
   U2077 : XNOR2_X1 port map( A => n3020, B => n6994, ZN => n7922);
   U2095 : XNOR2_X1 port map( A => n6304, B => n6305, ZN => n7921);
   U2100 : INV_X1 port map( A => n7600, ZN => n20012);
   U2113 : XNOR2_X1 port map( A => n6233, B => n6232, ZN => n7932);
   U2148 : XNOR2_X1 port map( A => n5454, B => n5453, ZN => n8286);
   U2160 : NAND2_X1 port map( A1 => n804, A2 => n1082, ZN => n1081);
   U2194 : AND2_X1 port map( A1 => n4600, A2 => n30, ZN => n20203);
   U2218 : AND3_X1 port map( A1 => n4998, A2 => n4996, A3 => n4999, ZN => 
                           n20028);
   U2219 : NAND4_X1 port map( A1 => n5771, A2 => n5772, A3 => n5774, A4 => 
                           n5773, ZN => n6927);
   U2236 : INV_X1 port map( A => n5767, ZN => n5734);
   U2269 : BUF_X1 port map( A => n4501, Z => n6204);
   U2275 : INV_X1 port map( A => n5719, ZN => n5604);
   U2276 : NAND2_X1 port map( A1 => n19619, A2 => n4309, ZN => n4598);
   U2284 : INV_X1 port map( A => n4860, ZN => n20085);
   U2291 : OR2_X1 port map( A1 => n4793, A2 => n5108, ZN => n5104);
   U2292 : CLKBUF_X1 port map( A => n5112, Z => n20256);
   U2316 : BUF_X1 port map( A => n4317, Z => n4325);
   U2339 : INV_X1 port map( A => n5717, ZN => n20034);
   U2345 : OR2_X1 port map( A1 => n4489, A2 => n4488, ZN => n4501);
   U2373 : MUX2_X1 port map( A => n4226, B => n4224, S => n3996, Z => n3997);
   U2383 : OAI211_X1 port map( C1 => n4557, C2 => n4750, A => n3915, B => n3914
                           , ZN => n6049);
   U2396 : XNOR2_X1 port map( A => Key(112), B => Plaintext(112), ZN => n5083);
   U2404 : OR2_X1 port map( A1 => n6379, A2 => n5728, ZN => n1746);
   U2419 : AND2_X1 port map( A1 => n20034, A2 => n5719, ZN => n4368);
   U2420 : OR2_X1 port map( A1 => n5328, A2 => n6048, ZN => n2081);
   U2447 : AND2_X1 port map( A1 => n5063, A2 => n5064, ZN => n20036);
   U2460 : INV_X1 port map( A => n5643, ZN => n5645);
   U2472 : OR2_X1 port map( A1 => n5002, A2 => n5571, ZN => n20282);
   U2473 : CLKBUF_X1 port map( A => n5276, Z => n5818);
   U2474 : OR2_X1 port map( A1 => n7674, A2 => n8365, ZN => n8362);
   U2481 : INV_X1 port map( A => n6523, ZN => n20314);
   U2496 : BUF_X1 port map( A => n6345, Z => n7504);
   U2500 : INV_X1 port map( A => n9114, ZN => n20346);
   U2504 : INV_X1 port map( A => n9239, ZN => n20322);
   U2530 : CLKBUF_X1 port map( A => n8087, Z => n20254);
   U2604 : INV_X1 port map( A => n9329, ZN => n20313);
   U2605 : AND2_X1 port map( A1 => n9003, A2 => n2883, ZN => n20037);
   U2609 : NAND2_X1 port map( A1 => n7565, A2 => n7566, ZN => n9362);
   U2660 : AND3_X1 port map( A1 => n3311, A2 => n8255, A3 => n769, ZN => n20146
                           );
   U2662 : CLKBUF_X1 port map( A => n8985, Z => n19827);
   U2705 : OR2_X1 port map( A1 => n9122, A2 => n8812, ZN => n8457);
   U2723 : XNOR2_X1 port map( A => n10602, B => n20324, ZN => n19505);
   U2724 : OR2_X1 port map( A1 => n20366, A2 => n11142, ZN => n10961);
   U2735 : AOI22_X1 port map( A1 => n12107, A2 => n12104, B1 => n3186, B2 => 
                           n3601, ZN => n11633);
   U2741 : INV_X1 port map( A => n12008, ZN => n12507);
   U2787 : XNOR2_X1 port map( A => n13047, B => n20053, ZN => n12676);
   U2790 : INV_X1 port map( A => n12258, ZN => n13146);
   U2799 : XNOR2_X1 port map( A => n2189, B => n13252, ZN => n14268);
   U2848 : OAI21_X1 port map( B1 => n12655, B2 => n14788, A => n14790, ZN => 
                           n20284);
   U2861 : XNOR2_X1 port map( A => n12587, B => n12588, ZN => n14787);
   U2862 : CLKBUF_X1 port map( A => n14679, Z => n20120);
   U2908 : INV_X1 port map( A => n15505, ZN => n20288);
   U2949 : INV_X1 port map( A => n15221, ZN => n15665);
   U2972 : NOR2_X1 port map( A1 => n15204, A2 => n15756, ZN => n15208);
   U3011 : INV_X1 port map( A => n16129, ZN => n747);
   U3079 : NAND4_X1 port map( A1 => n2815, A2 => n15758, A3 => n15757, A4 => 
                           n15760, ZN => n66);
   U3102 : OR2_X1 port map( A1 => n15540, A2 => n20006, ZN => n14911);
   U3127 : AND2_X1 port map( A1 => n15661, A2 => n15662, ZN => n20021);
   U3128 : INV_X1 port map( A => n16295, ZN => n16880);
   U3157 : OAI21_X1 port map( B1 => n15765, B2 => n15248, A => n15247, ZN => 
                           n19893);
   U3164 : XNOR2_X1 port map( A => n16964, B => n14987, ZN => n16284);
   U3169 : XNOR2_X1 port map( A => n16044, B => n17407, ZN => n16769);
   U3186 : OR2_X1 port map( A1 => n17690, A2 => n17691, ZN => n20307);
   U3232 : XNOR2_X1 port map( A => n963, B => n17140, ZN => n3066);
   U3253 : INV_X1 port map( A => n18620, ZN => n19509);
   U3394 : OR2_X1 port map( A1 => n16155, A2 => n18057, ZN => n19169);
   U3422 : CLKBUF_X1 port map( A => Key(159), Z => n2079);
   U3442 : CLKBUF_X1 port map( A => Key(93), Z => n2263);
   U3460 : CLKBUF_X1 port map( A => Key(41), Z => n345);
   U3532 : NAND3_X1 port map( A1 => n13950, A2 => n14690, A3 => n14688, ZN => 
                           n20014);
   U3558 : NAND2_X1 port map( A1 => n4855, A2 => n4907, ZN => n20015);
   U3644 : XOR2_X1 port map( A => Key(108), B => Plaintext(108), Z => n20016);
   U3680 : INV_X1 port map( A => n5859, ZN => n20334);
   U3710 : OR2_X1 port map( A1 => n4714, A2 => n4788, ZN => n20017);
   U3753 : INV_X1 port map( A => n4501, ZN => n6218);
   U3790 : INV_X1 port map( A => n2792, ZN => n20057);
   U3845 : INV_X1 port map( A => n12514, ZN => n20073);
   U3849 : XOR2_X1 port map( A => n13778, B => n13266, Z => n20018);
   U3860 : INV_X1 port map( A => n19043, ZN => n20074);
   U3901 : XOR2_X1 port map( A => n16092, B => n16093, Z => n20019);
   U4044 : NAND2_X1 port map( A1 => n1354, A2 => n8208, ZN => n20020);
   U4063 : XNOR2_X1 port map( A => n16295, B => n20100, ZN => n16297);
   U4074 : NAND2_X1 port map( A1 => n5610, A2 => n6152, ZN => n6160);
   U4086 : NAND2_X1 port map( A1 => n659, A2 => n2533, ZN => n19270);
   U4091 : NAND2_X1 port map( A1 => n20015, A2 => n4499, ZN => n3706);
   U4105 : NAND3_X1 port map( A1 => n1613, A2 => n1615, A3 => n1758, ZN => 
                           n20022);
   U4150 : AND2_X2 port map( A1 => n20023, A2 => n2969, ZN => n17002);
   U4156 : OAI21_X1 port map( B1 => n15399, B2 => n2968, A => n197, ZN => 
                           n20023);
   U4201 : NOR2_X1 port map( A1 => n276, A2 => n20024, ZN => n3076);
   U4320 : NAND2_X1 port map( A1 => n8001, A2 => n2548, ZN => n20024);
   U4326 : INV_X1 port map( A => n6871, ZN => n8140);
   U4335 : XNOR2_X1 port map( A => n6862, B => n6861, ZN => n6871);
   U4338 : NAND3_X1 port map( A1 => n19662, A2 => n15061, A3 => n15309, ZN => 
                           n14989);
   U4387 : NAND3_X1 port map( A1 => n20025, A2 => n15637, A3 => n15638, ZN => 
                           n19611);
   U4443 : NAND3_X1 port map( A1 => n20063, A2 => n230, A3 => n15843, ZN => 
                           n20025);
   U4526 : XNOR2_X1 port map( A => n13108, B => n13711, ZN => n12923);
   U4528 : NOR2_X2 port map( A1 => n11847, A2 => n11848, ZN => n13711);
   U4619 : NAND2_X1 port map( A1 => n12095, A2 => n12429, ZN => n11611);
   U4701 : NAND2_X1 port map( A1 => n3046, A2 => n3295, ZN => n20026);
   U4711 : INV_X1 port map( A => n10725, ZN => n20027);
   U4722 : NAND2_X1 port map( A1 => n5442, A2 => n5641, ZN => n4165);
   U4741 : OAI21_X1 port map( B1 => n8327, B2 => n9104, A => n8326, ZN => 
                           n10048);
   U4750 : NAND2_X1 port map( A1 => n7800, A2 => n7799, ZN => n2627);
   U4777 : NAND2_X2 port map( A1 => n4997, A2 => n20028, ZN => n7318);
   U4786 : OAI21_X1 port map( B1 => n3806, B2 => n9304, A => n9298, ZN => 
                           n20029);
   U4787 : OAI211_X1 port map( C1 => n17943, C2 => n3038, A => n1450, B => 
                           n3036, ZN => n3035);
   U4801 : INV_X1 port map( A => n10329, ZN => n10327);
   U4829 : NAND2_X1 port map( A1 => n2451, A2 => n13939, ZN => n20030);
   U4850 : INV_X1 port map( A => n20031, ZN => Ciphertext(26));
   U4928 : OAI211_X1 port map( C1 => n17743, C2 => n17742, A => n17740, B => 
                           n17741, ZN => n20031);
   U4985 : NAND3_X1 port map( A1 => n7703, A2 => n7542, A3 => n19881, ZN => 
                           n7544);
   U4998 : NOR2_X1 port map( A1 => n10505, A2 => n10836, ZN => n10523);
   U5019 : OAI21_X1 port map( B1 => n300, B2 => n18495, A => n20033, ZN => 
                           n17731);
   U5047 : NAND3_X1 port map( A1 => n18495, A2 => n300, A3 => n17729, ZN => 
                           n20033);
   U5088 : NAND3_X1 port map( A1 => n9303, A2 => n9302, A3 => n3788, ZN => 
                           n10598);
   U5117 : NAND2_X1 port map( A1 => n19922, A2 => n7871, ZN => n7422);
   U5141 : NAND2_X1 port map( A1 => n5595, A2 => n5519, ZN => n3409);
   U5143 : AOI21_X2 port map( B1 => n9557, B2 => n9558, A => n9556, ZN => 
                           n11659);
   U5185 : NOR2_X2 port map( A1 => n61, A2 => n4346, ZN => n5719);
   U5208 : NAND3_X1 port map( A1 => n20035, A2 => n7618, A3 => n586, ZN => 
                           n2097);
   U5255 : NAND2_X1 port map( A1 => n11387, A2 => n11386, ZN => n11393);
   U5264 : NAND2_X1 port map( A1 => n20038, A2 => n4943, ZN => n4949);
   U5284 : NAND2_X1 port map( A1 => n4941, A2 => n4940, ZN => n20038);
   U5288 : NOR2_X1 port map( A1 => n18630, A2 => n19509, ZN => n20039);
   U5304 : AND2_X1 port map( A1 => n14819, A2 => n14818, ZN => n20040);
   U5320 : NAND2_X1 port map( A1 => n15241, A2 => n15242, ZN => n17279);
   U5323 : NAND2_X1 port map( A1 => n12260, A2 => n19603, ZN => n13762);
   U5348 : NAND3_X1 port map( A1 => n3027, A2 => n20042, A3 => n20041, ZN => 
                           n1374);
   U5352 : NAND2_X1 port map( A1 => n18853, A2 => n3030, ZN => n20042);
   U5377 : NAND2_X1 port map( A1 => n8377, A2 => n8370, ZN => n7541);
   U5437 : NAND2_X1 port map( A1 => n4764, A2 => n4269, ZN => n20043);
   U5472 : NOR2_X1 port map( A1 => n4737, A2 => n20044, ZN => n19559);
   U5474 : INV_X1 port map( A => n4732, ZN => n20044);
   U5494 : NAND2_X1 port map( A1 => n4734, A2 => n4277, ZN => n4732);
   U5571 : NAND3_X1 port map( A1 => n14419, A2 => n14418, A3 => n14359, ZN => 
                           n3636);
   U5637 : NAND2_X1 port map( A1 => n20047, A2 => n20045, ZN => n15253);
   U5661 : NAND2_X1 port map( A1 => n20046, A2 => n17243, ZN => n20045);
   U5675 : NAND2_X1 port map( A1 => n17480, A2 => n20353, ZN => n20046);
   U5772 : NAND2_X1 port map( A1 => n15252, A2 => n17241, ZN => n20047);
   U5790 : NAND2_X1 port map( A1 => n20048, A2 => n18399, ZN => n18402);
   U5793 : OAI21_X1 port map( B1 => n18407, B2 => n18412, A => n20003, ZN => 
                           n20048);
   U5798 : XNOR2_X1 port map( A => n20050, B => n20049, ZN => Ciphertext(99));
   U5854 : INV_X1 port map( A => n18055, ZN => n20049);
   U5874 : NAND2_X1 port map( A1 => n20052, A2 => n20051, ZN => n20050);
   U5890 : NAND2_X1 port map( A1 => n18054, A2 => n18869, ZN => n20051);
   U5902 : INV_X1 port map( A => n2222, ZN => n20053);
   U5912 : NAND2_X1 port map( A1 => n12178, A2 => n2260, ZN => n13047);
   U5921 : NAND3_X1 port map( A1 => n18648, A2 => n19745, A3 => n18654, ZN => 
                           n582);
   U5924 : NOR2_X2 port map( A1 => n12314, A2 => n2338, ZN => n13309);
   U5937 : NAND2_X1 port map( A1 => n63, A2 => n20054, ZN => n10151);
   U5951 : NAND2_X1 port map( A1 => n369, A2 => n257, ZN => n11607);
   U5963 : AND2_X2 port map( A1 => n8147, A2 => n8148, ZN => n9346);
   U5983 : NAND3_X1 port map( A1 => n20056, A2 => n8301, A3 => n20055, ZN => 
                           n7452);
   U5984 : NAND2_X1 port map( A1 => n8304, A2 => n2792, ZN => n20055);
   U6035 : NAND2_X1 port map( A1 => n20057, A2 => n8305, ZN => n20056);
   U6096 : INV_X1 port map( A => n20059, ZN => n20058);
   U6104 : OAI21_X1 port map( B1 => n4951, B2 => n4911, A => n4477, ZN => 
                           n20059);
   U6116 : NAND2_X1 port map( A1 => n4476, A2 => n4958, ZN => n20060);
   U6123 : NAND2_X1 port map( A1 => n15400, A2 => n15892, ZN => n15540);
   U6161 : NAND2_X1 port map( A1 => n15442, A2 => n15676, ZN => n15678);
   U6181 : XNOR2_X1 port map( A => n20061, B => n18084, ZN => n8776);
   U6195 : NAND2_X1 port map( A1 => n8775, A2 => n2882, ZN => n20061);
   U6225 : NAND2_X1 port map( A1 => n1792, A2 => n3592, ZN => n3591);
   U6230 : NAND2_X1 port map( A1 => n397, A2 => n8295, ZN => n9100);
   U6235 : XNOR2_X1 port map( A => n13233, B => n20018, ZN => n13235);
   U6242 : NAND3_X1 port map( A1 => n20062, A2 => n4286, A3 => n4287, ZN => 
                           n1985);
   U6250 : NAND2_X1 port map( A1 => n4288, A2 => n4623, ZN => n20062);
   U6328 : OR2_X1 port map( A1 => n7848, A2 => n8079, ZN => n7849);
   U6338 : NAND2_X1 port map( A1 => n19354, A2 => n16540, ZN => n17234);
   U6343 : INV_X1 port map( A => n15845, ZN => n20063);
   U6346 : NAND2_X1 port map( A1 => n4913, A2 => n4914, ZN => n4915);
   U6348 : NAND2_X1 port map( A1 => n16542, A2 => n20065, ZN => n19339);
   U6353 : NAND2_X1 port map( A1 => n16541, A2 => n19352, ZN => n16542);
   U6392 : NAND2_X1 port map( A1 => n20014, A2 => n20066, ZN => n15221);
   U6443 : NAND2_X1 port map( A1 => n13365, A2 => n14696, ZN => n20066);
   U6448 : NAND2_X1 port map( A1 => n20068, A2 => n20067, ZN => n5612);
   U6455 : NAND3_X1 port map( A1 => n4392, A2 => n4681, A3 => n4486, ZN => 
                           n20067);
   U6462 : NAND2_X1 port map( A1 => n4390, A2 => n4389, ZN => n20068);
   U6463 : NAND2_X1 port map( A1 => n19347, A2 => n16673, ZN => n16635);
   U6472 : OAI211_X1 port map( C1 => n18365, C2 => n18364, A => n20070, B => 
                           n20069, ZN => n18368);
   U6481 : OR2_X1 port map( A1 => n18360, A2 => n17936, ZN => n20069);
   U6491 : NAND2_X1 port map( A1 => n20071, A2 => n18360, ZN => n20070);
   U6500 : INV_X1 port map( A => n18361, ZN => n20071);
   U6509 : NAND2_X1 port map( A1 => n19956, A2 => n17508, ZN => n20072);
   U6519 : NOR2_X1 port map( A1 => n12323, A2 => n20073, ZN => n2658);
   U6520 : NAND2_X1 port map( A1 => n12326, A2 => n11997, ZN => n12323);
   U6539 : OAI22_X1 port map( A1 => n19045, A2 => n20074, B1 => n19047, B2 => 
                           n19992, ZN => n18083);
   U6547 : NAND3_X2 port map( A1 => n15869, A2 => n20077, A3 => n20076, ZN => 
                           n17124);
   U6549 : NAND2_X1 port map( A1 => n15865, A2 => n15864, ZN => n20076);
   U6564 : NAND2_X1 port map( A1 => n15867, A2 => n15866, ZN => n20077);
   U6586 : NAND2_X2 port map( A1 => n28, A2 => n20079, ZN => n15720);
   U6634 : NAND2_X1 port map( A1 => n1350, A2 => n1352, ZN => n20079);
   U6660 : AND3_X2 port map( A1 => n3417, A2 => n1012, A3 => n3416, ZN => 
                           n10430);
   U6673 : OAI21_X2 port map( B1 => n11775, B2 => n11180, A => n11181, ZN => 
                           n13833);
   U6732 : NAND2_X1 port map( A1 => n7459, A2 => n2021, ZN => n1567);
   U6735 : INV_X1 port map( A => n5861, ZN => n5615);
   U6741 : NAND2_X1 port map( A1 => n5859, A2 => n3188, ZN => n5861);
   U6772 : NAND2_X1 port map( A1 => n15078, A2 => n2723, ZN => n14479);
   U6797 : OR3_X1 port map( A1 => n17676, A2 => n20512, A3 => n17867, ZN => 
                           n16000);
   U6830 : NAND3_X1 port map( A1 => n3283, A2 => n3285, A3 => n16734, ZN => 
                           n19135);
   U6851 : NAND3_X1 port map( A1 => n16733, A2 => n3287, A3 => n16732, ZN => 
                           n16734);
   U6889 : NAND2_X1 port map( A1 => n20080, A2 => n2089, ZN => n7896);
   U6905 : NAND2_X1 port map( A1 => n20082, A2 => n20504, ZN => n20080);
   U6918 : OAI21_X1 port map( B1 => n8184, B2 => n8059, A => n7892, ZN => 
                           n20082);
   U6948 : OAI21_X1 port map( B1 => n18613, B2 => n18625, A => n18629, ZN => 
                           n18179);
   U6949 : NAND2_X1 port map( A1 => n18622, A2 => n19679, ZN => n18629);
   U7002 : NAND3_X1 port map( A1 => n3085, A2 => n17506, A3 => n975, ZN => 
                           n19773);
   U7007 : NAND2_X1 port map( A1 => n339, A2 => n16480, ZN => n3085);
   U7022 : NAND2_X1 port map( A1 => n3252, A2 => n14468, ZN => n13924);
   U7115 : XNOR2_X2 port map( A => n12706, B => n12705, ZN => n14468);
   U7116 : NAND2_X2 port map( A1 => n20084, A2 => n20083, ZN => n6068);
   U7124 : NAND3_X1 port map( A1 => n3989, A2 => n4860, A3 => n4498, ZN => 
                           n20083);
   U7135 : NAND2_X1 port map( A1 => n3991, A2 => n20085, ZN => n20084);
   U7140 : NAND2_X1 port map( A1 => n12508, A2 => n12008, ZN => n126);
   U7153 : AND2_X2 port map( A1 => n12362, A2 => n12363, ZN => n12008);
   U7188 : NAND2_X1 port map( A1 => n2188, A2 => n20086, ZN => n8089);
   U7233 : OAI21_X1 port map( B1 => n1211, B2 => n8705, A => n20087, ZN => 
                           n2776);
   U7264 : NAND2_X1 port map( A1 => n2777, A2 => n1211, ZN => n20087);
   U7378 : NAND3_X1 port map( A1 => n20088, A2 => n5075, A3 => n5076, ZN => 
                           n448);
   U7405 : NAND2_X1 port map( A1 => n5074, A2 => n5080, ZN => n20088);
   U7406 : NOR2_X2 port map( A1 => n11705, A2 => n20089, ZN => n13623);
   U7424 : AOI21_X1 port map( B1 => n11702, B2 => n11703, A => n11701, ZN => 
                           n20089);
   U7425 : NAND2_X1 port map( A1 => n17557, A2 => n2797, ZN => n18620);
   U7471 : INV_X1 port map( A => n20090, ZN => n18315);
   U7472 : OAI22_X1 port map( A1 => n18309, A2 => n19340, B1 => n19309, B2 => 
                           n19311, ZN => n20090);
   U7554 : XOR2_X1 port map( A => n17034, B => n17032, Z => n17039);
   U7562 : OR2_X1 port map( A1 => n20091, A2 => n19758, ZN => n3579);
   U7570 : NAND2_X1 port map( A1 => n19526, A2 => n18511, ZN => n20091);
   U7592 : INV_X1 port map( A => n18057, ZN => n1035);
   U7606 : XOR2_X1 port map( A => n13097, B => n13400, Z => n13102);
   U7629 : XNOR2_X1 port map( A => n14942, B => n14943, ZN => n20092);
   U7644 : OAI21_X1 port map( B1 => n20330, B2 => n14352, A => n20329, ZN => 
                           n14329);
   U7657 : MUX2_X1 port map( A => n17455, B => n17983, S => n20132, Z => n20093
                           );
   U7684 : NAND2_X1 port map( A1 => n17313, A2 => n17312, ZN => n18834);
   U7686 : OR2_X1 port map( A1 => n17790, A2 => n17791, ZN => n17794);
   U7717 : BUF_X1 port map( A => n15876, Z => n20094);
   U7720 : OAI22_X1 port map( A1 => n2675, A2 => n3366, B1 => n2678, B2 => 
                           n2677, ZN => n15876);
   U7738 : XNOR2_X1 port map( A => n9673, B => n9672, ZN => n20095);
   U7790 : AOI21_X1 port map( B1 => n3116, B2 => n19667, A => n3115, ZN => 
                           n18151);
   U7826 : NAND2_X1 port map( A1 => n17319, A2 => n17318, ZN => n20097);
   U7835 : XNOR2_X1 port map( A => n9604, B => n9603, ZN => n11290);
   U7836 : BUF_X1 port map( A => n17281, Z => n20098);
   U7840 : OAI211_X1 port map( C1 => n15885, C2 => n16012, A => n13970, B => 
                           n13969, ZN => n17281);
   U7851 : MUX2_X2 port map( A => n19111, B => n19106, S => n19110, Z => n19093
                           );
   U7852 : XNOR2_X1 port map( A => n10097, B => n10096, ZN => n20099);
   U7880 : XNOR2_X1 port map( A => n10097, B => n10096, ZN => n11360);
   U7931 : AOI22_X2 port map( A1 => n12092, A2 => n12091, B1 => n12090, B2 => 
                           n12089, ZN => n13462);
   U7934 : CLKBUF_X1 port map( A => n14112, Z => n15423);
   U7948 : AOI22_X1 port map( A1 => n15197, A2 => n15198, B1 => n15500, B2 => 
                           n15196, ZN => n20100);
   U7961 : AOI22_X1 port map( A1 => n15197, A2 => n15198, B1 => n15500, B2 => 
                           n15196, ZN => n16746);
   U7962 : XNOR2_X1 port map( A => n17415, B => n17414, ZN => n20101);
   U7978 : XNOR2_X1 port map( A => n15764, B => n15763, ZN => n20240);
   U7982 : NAND3_X2 port map( A1 => n11941, A2 => n11940, A3 => n1400, ZN => 
                           n13390);
   U8002 : AOI21_X1 port map( B1 => n15725, B2 => n15724, A => n15723, ZN => 
                           n20102);
   U8020 : AOI21_X1 port map( B1 => n15725, B2 => n15724, A => n15723, ZN => 
                           n16407);
   U8030 : INV_X1 port map( A => n15165, ZN => n20103);
   U8063 : BUF_X1 port map( A => n12888, Z => n19513);
   U8065 : NAND3_X1 port map( A1 => n2007, A2 => n15161, A3 => n2293, ZN => 
                           n20104);
   U8096 : NAND3_X1 port map( A1 => n2007, A2 => n15161, A3 => n2293, ZN => 
                           n17299);
   U8098 : XNOR2_X1 port map( A => n3831, B => Key(70), ZN => n20105);
   U8108 : BUF_X1 port map( A => n11515, Z => n20106);
   U8161 : XNOR2_X1 port map( A => n3831, B => Key(70), ZN => n4420);
   U8164 : XNOR2_X1 port map( A => n9982, B => n9981, ZN => n11515);
   U8177 : XNOR2_X1 port map( A => n6549, B => n6548, ZN => n20107);
   U8180 : XNOR2_X1 port map( A => n6549, B => n6548, ZN => n20108);
   U8197 : XNOR2_X1 port map( A => n16428, B => n16427, ZN => n20109);
   U8225 : OAI21_X1 port map( B1 => n3081, B2 => n17507, A => n3080, ZN => 
                           n20110);
   U8362 : OAI21_X2 port map( B1 => n15052, B2 => n15053, A => n15051, ZN => 
                           n16873);
   U8368 : NAND2_X1 port map( A1 => n1106, A2 => n3388, ZN => n20111);
   U8372 : NAND2_X1 port map( A1 => n14616, A2 => n14615, ZN => n20112);
   U8376 : BUF_X1 port map( A => n2748, Z => n20113);
   U8382 : XOR2_X1 port map( A => n16361, B => n16362, Z => n20114);
   U8400 : OAI21_X1 port map( B1 => n7984, B2 => n7921, A => n1726, ZN => n502)
                           ;
   U8404 : NOR2_X1 port map( A1 => n8948, A2 => n528, ZN => n20115);
   U8429 : NOR2_X1 port map( A1 => n8948, A2 => n528, ZN => n10527);
   U8441 : OR2_X1 port map( A1 => n18036, A2 => n18035, ZN => n20117);
   U8449 : OR2_X1 port map( A1 => n15733, A2 => n3431, ZN => n15736);
   U8450 : OR2_X1 port map( A1 => n11360, A2 => n10112, ZN => n11358);
   U8647 : NAND3_X1 port map( A1 => n1469, A2 => n13960, A3 => n13959, ZN => 
                           n15879);
   U8653 : NOR2_X1 port map( A1 => n15098, A2 => n15099, ZN => n20121);
   U8720 : XNOR2_X1 port map( A => n13420, B => n13421, ZN => n14679);
   U8727 : NOR2_X1 port map( A1 => n15098, A2 => n15099, ZN => n2542);
   U8792 : OAI211_X2 port map( C1 => n12346, C2 => n12497, A => n12006, B => 
                           n2901, ZN => n13677);
   U8906 : NAND2_X1 port map( A1 => n11737, A2 => n11736, ZN => n20123);
   U8909 : AND2_X1 port map( A1 => n2414, A2 => n17866, ZN => n20124);
   U8921 : NAND2_X1 port map( A1 => n11737, A2 => n11736, ZN => n13695);
   U8949 : AOI21_X1 port map( B1 => n15715, B2 => n15716, A => n20094, ZN => 
                           n73);
   U8950 : OAI21_X1 port map( B1 => n14976, B2 => n14977, A => n14975, ZN => 
                           n20125);
   U8956 : OAI21_X1 port map( B1 => n14976, B2 => n14977, A => n14975, ZN => 
                           n20126);
   U8959 : OAI21_X1 port map( B1 => n14976, B2 => n14977, A => n14975, ZN => 
                           n17327);
   U9082 : XNOR2_X1 port map( A => n16710, B => n16709, ZN => n20127);
   U9141 : NAND2_X1 port map( A1 => n3205, A2 => n18038, ZN => n20128);
   U9239 : XOR2_X1 port map( A => n16877, B => n16876, Z => n20129);
   U9251 : AND2_X1 port map( A1 => n17313, A2 => n17312, ZN => n20130);
   U9293 : NAND2_X1 port map( A1 => n2268, A2 => n17834, ZN => n20131);
   U9294 : NAND2_X1 port map( A1 => n2268, A2 => n17834, ZN => n19074);
   U9310 : XNOR2_X1 port map( A => n17257, B => n17256, ZN => n20132);
   U9311 : BUF_X1 port map( A => n15697, Z => n20133);
   U9320 : AOI22_X1 port map( A1 => n14014, A2 => n14013, B1 => n19488, B2 => 
                           n14012, ZN => n15697);
   U9322 : AND2_X1 port map( A1 => n8775, A2 => n2882, ZN => n20134);
   U9372 : AOI21_X1 port map( B1 => n12511, B2 => n1609, A => n12510, ZN => 
                           n12512);
   U9389 : INV_X1 port map( A => n14261, ZN => n20311);
   U9601 : OAI211_X1 port map( C1 => n14227, C2 => n14731, A => n14226, B => 
                           n14225, ZN => n15422);
   U9621 : OR2_X1 port map( A1 => n12657, A2 => n14791, ZN => n20283);
   U9622 : XNOR2_X1 port map( A => n14915, B => n15953, ZN => n20135);
   U9887 : OAI21_X1 port map( B1 => n17216, B2 => n17217, A => n17215, ZN => 
                           n18377);
   U10070 : INV_X1 port map( A => n15619, ZN => n20138);
   U10074 : OR2_X1 port map( A1 => n15309, A2 => n15059, ZN => n15396);
   U10135 : OAI21_X1 port map( B1 => n17596, B2 => n16657, A => n16656, ZN => 
                           n20140);
   U10138 : INV_X1 port map( A => n14792, ZN => n20141);
   U10232 : OAI21_X1 port map( B1 => n17713, B2 => n20221, A => n17712, ZN => 
                           n20142);
   U10284 : XNOR2_X1 port map( A => Key(5), B => Plaintext(5), ZN => n20143);
   U10490 : XNOR2_X1 port map( A => Key(5), B => Plaintext(5), ZN => n4622);
   U10523 : INV_X1 port map( A => n19942, ZN => n20144);
   U10721 : BUF_X1 port map( A => n7475, Z => n19942);
   U10869 : INV_X1 port map( A => n15696, ZN => n20145);
   U10875 : BUF_X1 port map( A => n18468, Z => n20148);
   U10965 : OAI21_X1 port map( B1 => n1897, B2 => n16483, A => n16482, ZN => 
                           n18468);
   U10966 : OR2_X1 port map( A1 => n11105, A2 => n11104, ZN => n20300);
   U10995 : NAND3_X1 port map( A1 => n5904, A2 => n5903, A3 => n4847, ZN => 
                           n20149);
   U11107 : NAND3_X1 port map( A1 => n5904, A2 => n5903, A3 => n4847, ZN => 
                           n6090);
   U11343 : OAI21_X1 port map( B1 => n4843, B2 => n4842, A => n3978, ZN => 
                           n5904);
   U11347 : XOR2_X1 port map( A => n16536, B => n16537, Z => n20150);
   U11361 : OR2_X1 port map( A1 => n16128, A2 => n15607, ZN => n15733);
   U11374 : BUF_X1 port map( A => n15671, Z => n20151);
   U11375 : AOI22_X1 port map( A1 => n13459, A2 => n14678, B1 => n13458, B2 => 
                           n14550, ZN => n15671);
   U11406 : OAI211_X1 port map( C1 => n16677, C2 => n16676, A => n16675, B => 
                           n2206, ZN => n18067);
   U11492 : MUX2_X1 port map( A => n8970, B => n7727, S => n9256, Z => n7738);
   U11568 : OAI21_X1 port map( B1 => n11075, B2 => n11486, A => n11074, ZN => 
                           n20153);
   U11577 : OAI21_X1 port map( B1 => n11075, B2 => n11486, A => n11074, ZN => 
                           n12253);
   U11578 : XNOR2_X1 port map( A => n7069, B => n7068, ZN => n20154);
   U11590 : XNOR2_X1 port map( A => n7069, B => n7068, ZN => n7991);
   U11591 : OAI211_X1 port map( C1 => n11927, C2 => n11926, A => n11924, B => 
                           n11925, ZN => n13702);
   U11598 : OR2_X1 port map( A1 => n8468, A2 => n8467, ZN => n20156);
   U11633 : INV_X1 port map( A => n14571, ZN => n20157);
   U11647 : XNOR2_X2 port map( A => n13229, B => n13228, ZN => n14571);
   U11708 : OAI211_X2 port map( C1 => n15748, C2 => n19502, A => n15597, B => 
                           n15596, ZN => n16886);
   U11760 : XNOR2_X1 port map( A => n16890, B => n16889, ZN => n20158);
   U11764 : XNOR2_X1 port map( A => n16890, B => n16889, ZN => n18975);
   U11867 : NAND2_X2 port map( A1 => n19580, A2 => n12395, ZN => n13259);
   U11887 : OR2_X1 port map( A1 => n11174, A2 => n10962, ZN => n20317);
   U11905 : CLKBUF_X1 port map( A => n2984, Z => n20159);
   U12004 : NOR2_X1 port map( A1 => n17221, A2 => n16639, ZN => n16641);
   U12005 : BUF_X1 port map( A => n11871, Z => n20160);
   U12119 : BUF_X1 port map( A => n10332, Z => n20161);
   U12141 : XNOR2_X1 port map( A => n16074, B => n16073, ZN => n20162);
   U12142 : NAND3_X1 port map( A1 => n3343, A2 => n3344, A3 => n113, ZN => 
                           n20163);
   U12216 : AND2_X1 port map( A1 => n558, A2 => n559, ZN => n20164);
   U12364 : XNOR2_X1 port map( A => n7012, B => n7011, ZN => n20165);
   U12380 : XNOR2_X1 port map( A => n7012, B => n7011, ZN => n7833);
   U12385 : XNOR2_X1 port map( A => n6261, B => n6262, ZN => n20166);
   U12400 : OAI211_X1 port map( C1 => n15325, C2 => n1491, A => n15324, B => 
                           n15323, ZN => n20167);
   U12455 : OAI211_X1 port map( C1 => n15325, C2 => n1491, A => n15324, B => 
                           n15323, ZN => n17416);
   U12690 : XOR2_X1 port map( A => n15436, B => n15435, Z => n20168);
   U12691 : NAND2_X1 port map( A1 => n2959, A2 => n16445, ZN => n20169);
   U12752 : NOR2_X1 port map( A1 => n3565, A2 => n12512, ZN => n13619);
   U12862 : XOR2_X1 port map( A => n13593, B => n13594, Z => n20171);
   U13005 : XNOR2_X1 port map( A => n16597, B => n16598, ZN => n20172);
   U13267 : NAND2_X1 port map( A1 => n13505, A2 => n2138, ZN => n20173);
   U13268 : NAND2_X1 port map( A1 => n13505, A2 => n2138, ZN => n15457);
   U13269 : CLKBUF_X1 port map( A => n8220, Z => n20174);
   U13343 : XNOR2_X1 port map( A => n6473, B => n6472, ZN => n8220);
   U13458 : NOR2_X2 port map( A1 => n7670, A2 => n7669, ZN => n20176);
   U13544 : NOR2_X1 port map( A1 => n7670, A2 => n7669, ZN => n10200);
   U13545 : XNOR2_X1 port map( A => n6797, B => n6798, ZN => n20177);
   U13599 : AOI22_X1 port map( A1 => n13975, A2 => n19940, B1 => n13974, B2 => 
                           n14499, ZN => n20178);
   U13632 : AOI22_X1 port map( A1 => n13975, A2 => n19940, B1 => n13974, B2 => 
                           n14499, ZN => n15709);
   U13668 : XOR2_X1 port map( A => n963, B => n17140, Z => n20179);
   U13790 : XNOR2_X1 port map( A => n6455, B => n6454, ZN => n20180);
   U13873 : XNOR2_X1 port map( A => n13847, B => n2679, ZN => n20181);
   U13900 : XNOR2_X1 port map( A => n13847, B => n2679, ZN => n14603);
   U13981 : NOR2_X1 port map( A1 => n14735, A2 => n14734, ZN => n20182);
   U14024 : NOR2_X1 port map( A1 => n14735, A2 => n14734, ZN => n20183);
   U14113 : AOI22_X2 port map( A1 => n14955, A2 => n15043, B1 => n15802, B2 => 
                           n14954, ZN => n16711);
   U14196 : XNOR2_X1 port map( A => n16092, B => n16093, ZN => n20185);
   U14197 : INV_X1 port map( A => n12312, ZN => n20186);
   U14402 : AND2_X1 port map( A1 => n14573, A2 => n14572, ZN => n20187);
   U14403 : INV_X1 port map( A => n19877, ZN => n20188);
   U14462 : INV_X1 port map( A => n20235, ZN => n11404);
   U14587 : XNOR2_X1 port map( A => n7359, B => n7358, ZN => n20189);
   U14646 : INV_X1 port map( A => n10601, ZN => n20324);
   U14686 : XNOR2_X1 port map( A => n3908, B => Key(156), ZN => n20190);
   U14725 : AOI22_X1 port map( A1 => n11242, A2 => n11349, B1 => n11241, B2 => 
                           n11350, ZN => n12021);
   U14745 : NOR2_X1 port map( A1 => n15718, A2 => n73, ZN => n20192);
   U14746 : CLKBUF_X1 port map( A => n19237, Z => n20193);
   U14824 : NOR2_X1 port map( A1 => n15718, A2 => n73, ZN => n16027);
   U15015 : OAI21_X1 port map( B1 => n17902, B2 => n17901, A => n17900, ZN => 
                           n19237);
   U15022 : XOR2_X1 port map( A => n16920, B => n16919, Z => n20194);
   U15059 : XNOR2_X1 port map( A => n6223, B => n6224, ZN => n20195);
   U15154 : OAI22_X1 port map( A1 => n19519, A2 => n9579, B1 => n8577, B2 => 
                           n19715, ZN => n20196);
   U15165 : XNOR2_X1 port map( A => n6223, B => n6224, ZN => n7935);
   U15166 : AND2_X1 port map( A1 => n1640, A2 => n15310, ZN => n15397);
   U15361 : XNOR2_X1 port map( A => n6079, B => n6078, ZN => n20198);
   U15362 : OAI211_X1 port map( C1 => n12570, C2 => n13146, A => n12019, B => 
                           n12018, ZN => n20199);
   U15363 : XNOR2_X1 port map( A => n6079, B => n6078, ZN => n8055);
   U15385 : OAI211_X1 port map( C1 => n12570, C2 => n13146, A => n12019, B => 
                           n12018, ZN => n13059);
   U15421 : XNOR2_X1 port map( A => n6885, B => n6884, ZN => n20200);
   U15440 : OAI22_X1 port map( A1 => n11673, A2 => n12179, B1 => n11650, B2 => 
                           n11670, ZN => n20201);
   U15479 : XNOR2_X1 port map( A => Key(108), B => Plaintext(108), ZN => n20202
                           );
   U15500 : XNOR2_X1 port map( A => n13692, B => n13691, ZN => n20204);
   U15501 : XNOR2_X1 port map( A => n13692, B => n13691, ZN => n14378);
   U15534 : INV_X1 port map( A => n4136, ZN => n20205);
   U15535 : XOR2_X1 port map( A => n13061, B => n13062, Z => n20206);
   U15536 : XNOR2_X1 port map( A => n16995, B => n16994, ZN => n20207);
   U15562 : XNOR2_X1 port map( A => n5321, B => n7134, ZN => n20208);
   U15583 : XNOR2_X1 port map( A => n6819, B => n7218, ZN => n20209);
   U15584 : INV_X1 port map( A => n912, ZN => n20330);
   U15772 : OAI211_X1 port map( C1 => n8784, C2 => n8783, A => n3807, B => 
                           n8782, ZN => n20210);
   U15813 : OAI211_X1 port map( C1 => n8784, C2 => n8783, A => n3807, B => 
                           n8782, ZN => n20211);
   U15817 : OR2_X1 port map( A1 => n8780, A2 => n9107, ZN => n3807);
   U15842 : XNOR2_X1 port map( A => n16526, B => n16525, ZN => n20212);
   U15872 : XNOR2_X1 port map( A => n16526, B => n16525, ZN => n19362);
   U16014 : OR2_X1 port map( A1 => n5941, A2 => n20243, ZN => n8295);
   U16031 : XOR2_X1 port map( A => n13663, B => n13662, Z => n20213);
   U16085 : XNOR2_X2 port map( A => n2772, B => n2771, ZN => n10980);
   U16154 : AND4_X1 port map( A1 => n17192, A2 => n17191, A3 => n17190, A4 => 
                           n17189, ZN => n20214);
   U16158 : INV_X1 port map( A => n8103, ZN => n9326);
   U16244 : OAI211_X1 port map( C1 => n4404, C2 => n5856, A => n4403, B => 
                           n4402, ZN => n20216);
   U16246 : OAI211_X1 port map( C1 => n4404, C2 => n5856, A => n4403, B => 
                           n4402, ZN => n2571);
   U16312 : XOR2_X1 port map( A => n16060, B => n16061, Z => n20217);
   U16315 : AOI22_X1 port map( A1 => n17614, A2 => n17613, B1 => n17612, B2 => 
                           n17611, ZN => n20218);
   U16316 : XNOR2_X1 port map( A => n17355, B => n16181, ZN => n20219);
   U16389 : XNOR2_X1 port map( A => n16774, B => n16773, ZN => n18956);
   U16404 : NAND2_X1 port map( A1 => n11963, A2 => n3396, ZN => n20222);
   U16419 : NAND2_X1 port map( A1 => n11963, A2 => n3396, ZN => n20223);
   U16496 : OAI211_X1 port map( C1 => n262, C2 => n9328, A => n1408, B => 
                           n20313, ZN => n2173);
   U16499 : NAND4_X1 port map( A1 => n5738, A2 => n5740, A3 => n5737, A4 => 
                           n5739, ZN => n20224);
   U16598 : NAND4_X1 port map( A1 => n5738, A2 => n5740, A3 => n5737, A4 => 
                           n5739, ZN => n20225);
   U16600 : NAND4_X1 port map( A1 => n5738, A2 => n5740, A3 => n5737, A4 => 
                           n5739, ZN => n6767);
   U16620 : OAI211_X1 port map( C1 => n5823, C2 => n5448, A => n3567, B => 
                           n3568, ZN => n20227);
   U16663 : XOR2_X1 port map( A => n9799, B => n9462, Z => n20228);
   U16702 : OAI211_X1 port map( C1 => n5823, C2 => n5448, A => n3567, B => 
                           n3568, ZN => n7121);
   U16718 : XNOR2_X1 port map( A => Key(140), B => Plaintext(140), ZN => n20229
                           );
   U16727 : XNOR2_X1 port map( A => n10584, B => n20491, ZN => n10218);
   U16742 : XNOR2_X1 port map( A => Key(140), B => Plaintext(140), ZN => n5017)
                           ;
   U16743 : XOR2_X1 port map( A => n15250, B => n15968, Z => n20230);
   U16751 : NOR2_X1 port map( A1 => n16464, A2 => n2297, ZN => n20231);
   U16761 : NOR2_X1 port map( A1 => n16464, A2 => n2297, ZN => n20232);
   U16783 : NOR2_X1 port map( A1 => n16464, A2 => n2297, ZN => n18454);
   U16803 : XNOR2_X1 port map( A => n10065, B => n10064, ZN => n20233);
   U16865 : XNOR2_X1 port map( A => n10065, B => n10064, ZN => n10897);
   U16870 : OR2_X1 port map( A1 => n16632, A2 => n17513, ZN => n20234);
   U16909 : OAI211_X2 port map( C1 => n15105, C2 => n15104, A => n15103, B => 
                           n15102, ZN => n16695);
   U16953 : XNOR2_X2 port map( A => n20236, B => n9575, ZN => n20235);
   U16993 : XOR2_X1 port map( A => n9692, B => n9573, Z => n20236);
   U17032 : XOR2_X1 port map( A => n12906, B => n13848, Z => n20237);
   U17203 : XNOR2_X1 port map( A => n15937, B => n15938, ZN => n20239);
   U17204 : XNOR2_X1 port map( A => n15937, B => n15938, ZN => n17172);
   U17292 : NAND4_X1 port map( A1 => n17192, A2 => n17191, A3 => n17190, A4 => 
                           n17189, ZN => n19115);
   U17339 : XNOR2_X1 port map( A => n15764, B => n15763, ZN => n19354);
   U17354 : BUF_X1 port map( A => n5563, Z => n20241);
   U17424 : XNOR2_X1 port map( A => n16532, B => n16531, ZN => n20242);
   U17433 : XOR2_X1 port map( A => n5962, B => n5961, Z => n20243);
   U17571 : NAND2_X2 port map( A1 => n2591, A2 => n14345, ZN => n15906);
   U17575 : XNOR2_X1 port map( A => n4065, B => n4064, ZN => n20247);
   U17605 : XNOR2_X1 port map( A => n20248, B => n20249, ZN => n14410);
   U17658 : XNOR2_X1 port map( A => n13388, B => n13389, ZN => n20248);
   U17743 : XOR2_X1 port map( A => n13393, B => n13392, Z => n20249);
   U17754 : NOR2_X2 port map( A1 => n9084, A2 => n9083, ZN => n9986);
   U17863 : BUF_X1 port map( A => n6919, Z => n20250);
   U17938 : XOR2_X1 port map( A => n1074, B => n1073, Z => n20251);
   U17977 : XNOR2_X1 port map( A => n6741, B => n6740, ZN => n20252);
   U17978 : OAI211_X1 port map( C1 => n874, C2 => n12622, A => n12621, B => 
                           n12620, ZN => n20253);
   U18011 : XNOR2_X1 port map( A => n6741, B => n6740, ZN => n8376);
   U18034 : OAI211_X1 port map( C1 => n874, C2 => n12622, A => n12621, B => 
                           n12620, ZN => n13585);
   U18132 : OAI21_X1 port map( B1 => n11483, B2 => n11215, A => n11214, ZN => 
                           n12479);
   U18140 : XNOR2_X1 port map( A => n2738, B => Key(79), ZN => n5112);
   U18172 : XNOR2_X1 port map( A => n5940, B => n5939, ZN => n20257);
   U18173 : XOR2_X1 port map( A => n17274, B => n17273, Z => n20258);
   U18174 : BUF_X1 port map( A => n18866, Z => n20259);
   U18175 : OAI21_X1 port map( B1 => n19575, B2 => n18040, A => n18039, ZN => 
                           n18866);
   U18182 : OAI21_X1 port map( B1 => n11983, B2 => n12619, A => n11982, ZN => 
                           n20260);
   U18186 : INV_X1 port map( A => n19598, ZN => n20261);
   U18236 : INV_X1 port map( A => n8370, ZN => n20294);
   U18238 : XNOR2_X1 port map( A => n12903, B => n12904, ZN => n20262);
   U18259 : XNOR2_X1 port map( A => n12903, B => n12904, ZN => n701);
   U18333 : NOR2_X1 port map( A1 => n19068, A2 => n18151, ZN => n19079);
   U18334 : XOR2_X1 port map( A => n13532, B => n13531, Z => n20263);
   U18384 : XNOR2_X1 port map( A => n16121, B => n16120, ZN => n20264);
   U18430 : AND3_X2 port map( A1 => n3428, A2 => n3432, A3 => n3426, ZN => 
                           n16980);
   U18458 : OAI21_X1 port map( B1 => n1244, B2 => n1243, A => n1242, ZN => 
                           n20265);
   U18483 : OAI21_X1 port map( B1 => n1244, B2 => n1243, A => n1242, ZN => 
                           n8990);
   U18498 : XNOR2_X1 port map( A => n10219, B => n19818, ZN => n20268);
   U18506 : XNOR2_X1 port map( A => n16406, B => n16027, ZN => n20269);
   U18543 : XNOR2_X1 port map( A => n7280, B => n7281, ZN => n20270);
   U18544 : XNOR2_X1 port map( A => n6524, B => n20314, ZN => n8083);
   U18661 : XNOR2_X1 port map( A => n14017, B => n14018, ZN => n20271);
   U18682 : XOR2_X1 port map( A => n13069, B => n13068, Z => n20272);
   U18691 : XOR2_X1 port map( A => n15854, B => n15855, Z => n20273);
   U18699 : XOR2_X1 port map( A => n6930, B => n6929, Z => n20274);
   U18700 : XNOR2_X1 port map( A => n15969, B => n15968, ZN => n20275);
   U18720 : OAI21_X1 port map( B1 => n17385, B2 => n17384, A => n17383, ZN => 
                           n18831);
   U18793 : OAI211_X2 port map( C1 => n3118, C2 => n8341, A => n3119, B => 
                           n20277, ZN => n9563);
   U18794 : NAND2_X1 port map( A1 => n3122, A2 => n3121, ZN => n20277);
   U18896 : NAND2_X1 port map( A1 => n7685, A2 => n8381, ZN => n7716);
   U18897 : NAND2_X1 port map( A1 => n19561, A2 => n4080, ZN => n5707);
   U18912 : AOI22_X2 port map( A1 => n15169, A2 => n15168, B1 => n15378, B2 => 
                           n15170, ZN => n16615);
   U18922 : NAND2_X1 port map( A1 => n20279, A2 => n20278, ZN => n10758);
   U18923 : NAND2_X1 port map( A1 => n11526, A2 => n11521, ZN => n20278);
   U18946 : XNOR2_X1 port map( A => n20123, B => n12769, ZN => n13698);
   U18960 : NAND3_X1 port map( A1 => n12227, A2 => n10941, A3 => n12229, ZN => 
                           n10942);
   U19319 : NAND2_X2 port map( A1 => n20281, A2 => n738, ZN => n9576);
   U19359 : NAND2_X1 port map( A1 => n7512, A2 => n7511, ZN => n20281);
   U19489 : NAND2_X1 port map( A1 => n7852, A2 => n8159, ZN => n2840);
   U19545 : NAND2_X1 port map( A1 => n1865, A2 => n1868, ZN => n2630);
   U19579 : NAND2_X1 port map( A1 => n5001, A2 => n20282, ZN => n7088);
   U19580 : NAND3_X1 port map( A1 => n5770, A2 => n5545, A3 => n5734, ZN => 
                           n5740);
   U19581 : NAND2_X1 port map( A1 => n15473, A2 => n15767, ZN => n15478);
   U19585 : NAND3_X1 port map( A1 => n5147, A2 => n5146, A3 => n5572, ZN => 
                           n5152);
   U19629 : XNOR2_X1 port map( A => n13465, B => n13464, ZN => n20285);
   U19632 : NAND2_X1 port map( A1 => n4515, A2 => n4514, ZN => n5767);
   U19638 : NAND3_X1 port map( A1 => n338, A2 => n1383, A3 => n12663, ZN => 
                           n16347);
   U19693 : NAND3_X1 port map( A1 => n1478, A2 => n1477, A3 => n9361, ZN => 
                           n8964);
   U19705 : OR2_X1 port map( A1 => n15657, A2 => n12658, ZN => n12659);
   U19706 : OAI21_X2 port map( B1 => n488, B2 => n11657, A => n487, ZN => 
                           n13134);
   U19707 : NAND2_X1 port map( A1 => n19112, A2 => n19105, ZN => n20286);
   U19718 : NAND3_X1 port map( A1 => n7813, A2 => n7814, A3 => n7479, ZN => 
                           n465);
   U19731 : NAND2_X1 port map( A1 => n15275, A2 => n15270, ZN => n15272);
   U19749 : NAND2_X1 port map( A1 => n14935, A2 => n20288, ZN => n1613);
   U19751 : INV_X1 port map( A => n13615, ZN => n14597);
   U19752 : NAND2_X1 port map( A1 => n19647, A2 => n19372, ZN => n19646);
   U19753 : NAND2_X1 port map( A1 => n18216, A2 => n1194, ZN => n1193);
   U19754 : NAND2_X1 port map( A1 => n20005, A2 => n15702, ZN => n15141);
   U19755 : XNOR2_X1 port map( A => n20290, B => n19322, ZN => Ciphertext(175))
                           ;
   U19756 : NAND3_X1 port map( A1 => n19319, A2 => n19320, A3 => n19318, ZN => 
                           n20290);
   U19757 : OAI22_X1 port map( A1 => n19514, A2 => n13989, B1 => n15714, B2 => 
                           n15148, ZN => n13990);
   U19758 : NOR2_X1 port map( A1 => n16170, A2 => n20291, ZN => n16632);
   U19759 : NOR2_X1 port map( A1 => n14845, A2 => n16633, ZN => n20291);
   U19760 : NAND2_X1 port map( A1 => n7726, A2 => n7856, ZN => n20292);
   U19761 : OAI211_X1 port map( C1 => n8376, C2 => n19881, A => n20295, B => 
                           n20294, ZN => n20293);
   U19762 : NAND2_X1 port map( A1 => n8373, A2 => n19881, ZN => n20295);
   U19763 : INV_X1 port map( A => n4926, ZN => n4385);
   U19764 : NAND2_X1 port map( A1 => n3967, A2 => n4921, ZN => n4926);
   U19765 : NAND2_X1 port map( A1 => n20298, A2 => n20297, ZN => n12313);
   U19766 : NAND2_X1 port map( A1 => n11362, A2 => n11361, ZN => n20298);
   U19768 : NAND2_X1 port map( A1 => n10768, A2 => n11104, ZN => n20299);
   U19770 : NAND2_X1 port map( A1 => n3862, A2 => n3861, ZN => n20301);
   U19771 : XNOR2_X1 port map( A => n20302, B => n16599, ZN => n16385);
   U19772 : XNOR2_X1 port map( A => n19782, B => n2329, ZN => n20302);
   U19773 : NAND2_X1 port map( A1 => n20305, A2 => n20303, ZN => n12486);
   U19774 : NAND2_X1 port map( A1 => n12476, A2 => n20304, ZN => n20303);
   U19775 : INV_X1 port map( A => n19833, ZN => n20304);
   U19776 : NAND2_X1 port map( A1 => n12475, A2 => n19833, ZN => n20305);
   U19778 : NAND2_X1 port map( A1 => n689, A2 => n18946, ZN => n20306);
   U19779 : OAI211_X1 port map( C1 => n8672, C2 => n8674, A => n20309, B => 
                           n20308, ZN => n8519);
   U19780 : NAND2_X1 port map( A1 => n19857, A2 => n9023, ZN => n20308);
   U19781 : NAND2_X1 port map( A1 => n9022, A2 => n8672, ZN => n20309);
   U19782 : OAI21_X1 port map( B1 => n14260, B2 => n20311, A => n20310, ZN => 
                           n14019);
   U19783 : NAND2_X1 port map( A1 => n14260, A2 => n13981, ZN => n20310);
   U19784 : NAND2_X1 port map( A1 => n2889, A2 => n14702, ZN => n15370);
   U19785 : NAND2_X1 port map( A1 => n2890, A2 => n14230, ZN => n2889);
   U19786 : OR2_X2 port map( A1 => n3957, A2 => n20312, ZN => n3959);
   U19787 : NOR2_X1 port map( A1 => n3956, A2 => n4291, ZN => n20312);
   U19788 : NAND2_X1 port map( A1 => n7686, A2 => n8385, ZN => n8131);
   U19789 : NAND3_X1 port map( A1 => n2702, A2 => n1006, A3 => n20315, ZN => 
                           n8993);
   U19791 : OR3_X1 port map( A1 => n11528, A2 => n11527, A3 => n11521, ZN => 
                           n12221);
   U19792 : NAND2_X1 port map( A1 => n19761, A2 => n14396, ZN => n13615);
   U19793 : NAND2_X1 port map( A1 => n20316, A2 => n19421, ZN => n19423);
   U19795 : NAND3_X1 port map( A1 => n20318, A2 => n20317, A3 => n11176, ZN => 
                           n10656);
   U19796 : NAND2_X1 port map( A1 => n11178, A2 => n10962, ZN => n20318);
   U19797 : NOR2_X1 port map( A1 => n14637, A2 => n20319, ZN => n12974);
   U19798 : OR2_X1 port map( A1 => n19703, A2 => n14032, ZN => n20319);
   U19799 : NAND2_X1 port map( A1 => n20320, A2 => n210, ZN => n4896);
   U19800 : NAND2_X1 port map( A1 => n3231, A2 => n4136, ZN => n20320);
   U19801 : NAND3_X1 port map( A1 => n8053, A2 => n19474, A3 => n8193, ZN => 
                           n7626);
   U19802 : NAND2_X1 port map( A1 => n20322, A2 => n20321, ZN => n2637);
   U19803 : NAND2_X1 port map( A1 => n9241, A2 => n9240, ZN => n20321);
   U19804 : OAI21_X1 port map( B1 => n19606, B2 => n20505, A => n20323, ZN => 
                           n8543);
   U19805 : NAND2_X1 port map( A1 => n20505, A2 => n20476, ZN => n20323);
   U19808 : OAI21_X1 port map( B1 => n19100, B2 => n19101, A => n20326, ZN => 
                           n19610);
   U19809 : AOI22_X1 port map( A1 => n19101, A2 => n19105, B1 => n19112, B2 => 
                           n19118, ZN => n20326);
   U19810 : INV_X1 port map( A => n7688, ZN => n20327);
   U19811 : NAND2_X1 port map( A1 => n7685, A2 => n20327, ZN => n1422);
   U19812 : OR3_X1 port map( A1 => n9354, A2 => n8720, A3 => n9528, ZN => n592)
                           ;
   U19813 : OAI21_X1 port map( B1 => n2685, B2 => n2697, A => n20328, ZN => 
                           n14047);
   U19814 : NAND2_X1 port map( A1 => n19597, A2 => n14827, ZN => n20328);
   U19815 : NOR2_X1 port map( A1 => n5142, A2 => n5143, ZN => n6494);
   U19816 : NAND2_X1 port map( A1 => n14352, A2 => n14326, ZN => n20329);
   U19817 : NAND2_X1 port map( A1 => n3519, A2 => n2883, ZN => n2882);
   U19818 : NAND2_X1 port map( A1 => n2884, A2 => n1401, ZN => n3519);
   U19820 : OAI211_X1 port map( C1 => n17524, C2 => n17519, A => n17522, B => 
                           n20331, ZN => n17528);
   U19821 : INV_X1 port map( A => n17581, ZN => n20331);
   U19822 : INV_X1 port map( A => n699, ZN => n698);
   U19824 : NOR2_X1 port map( A1 => n14435, A2 => n14171, ZN => n14431);
   U19826 : NAND2_X1 port map( A1 => n20333, A2 => n20332, ZN => n4464);
   U19827 : NAND2_X1 port map( A1 => n6141, A2 => n5859, ZN => n20332);
   U19829 : AND2_X2 port map( A1 => n20335, A2 => n20337, ZN => n16335);
   U19830 : INV_X1 port map( A => n20336, ZN => n20335);
   U19831 : OAI21_X1 port map( B1 => n15519, B2 => n3821, A => n15518, ZN => 
                           n20336);
   U19832 : NAND2_X1 port map( A1 => n15522, A2 => n15521, ZN => n20337);
   U19833 : NAND2_X1 port map( A1 => n12490, A2 => n11912, ZN => n12492);
   U19834 : NAND2_X1 port map( A1 => n14090, A2 => n939, ZN => n15516);
   U19836 : OAI22_X1 port map( A1 => n3601, A2 => n11275, B1 => n11271, B2 => 
                           n11381, ZN => n20338);
   U19837 : OR2_X2 port map( A1 => n4149, A2 => n4150, ZN => n5643);
   U19838 : OAI22_X1 port map( A1 => n15112, A2 => n15113, B1 => n15114, B2 => 
                           n15604, ZN => n15118);
   U19839 : NAND2_X1 port map( A1 => n20112, A2 => n15275, ZN => n15113);
   U19841 : NAND2_X1 port map( A1 => n15370, A2 => n15371, ZN => n15565);
   U19842 : NAND2_X1 port map( A1 => n75, A2 => n78, ZN => n20339);
   U19843 : AND2_X2 port map( A1 => n1592, A2 => n1189, ZN => n12208);
   U19844 : NAND2_X1 port map( A1 => n19979, A2 => n5914, ZN => n5915);
   U19846 : NAND2_X1 port map( A1 => n10833, A2 => n11037, ZN => n20340);
   U19847 : NAND2_X1 port map( A1 => n15534, A2 => n15921, ZN => n20341);
   U19848 : NAND2_X1 port map( A1 => n20343, A2 => n2974, ZN => n20342);
   U19849 : NAND2_X1 port map( A1 => n15532, A2 => n15531, ZN => n20343);
   U19850 : NAND2_X1 port map( A1 => n20345, A2 => n20344, ZN => n8669);
   U19851 : NAND2_X1 port map( A1 => n9112, A2 => n9114, ZN => n20344);
   U19852 : OAI21_X1 port map( B1 => n1602, B2 => n9217, A => n20346, ZN => 
                           n20345);
   U19853 : AOI21_X2 port map( B1 => n11362, B2 => n11361, A => n3667, ZN => 
                           n19952);
   U19854 : AOI21_X2 port map( B1 => n12329, B2 => n12328, A => n13269, ZN => 
                           n19796);
   U19855 : AOI22_X2 port map( A1 => n1419, A2 => n12293, B1 => n11772, B2 => 
                           n12533, ZN => n19697);
   U19857 : OAI211_X2 port map( C1 => n12267, C2 => n12565, A => n976, B => 
                           n1043, ZN => n13703);
   U6130 : NAND2_X2 port map( A1 => n2159, A2 => n1975, ZN => n13725);
   U1841 : MUX2_X2 port map( A => n6103, B => n6102, S => n6101, Z => n7218);
   U720 : BUF_X2 port map( A => n4268, Z => n5024);
   U705 : OAI211_X2 port map( C1 => n5103, C2 => n1421, A => n5110, B => n1420,
                           ZN => n6010);
   U17999 : NOR2_X2 port map( A1 => n14583, A2 => n14582, ZN => n16750);
   U379 : BUF_X1 port map( A => n5589, Z => n19979);
   U1860 : NAND2_X2 port map( A1 => n3194, A2 => n1745, ZN => n7248);
   U12692 : NOR2_X2 port map( A1 => n3565, A2 => n12512, ZN => n20170);
   U2249 : OR2_X2 port map( A1 => n4164, A2 => n4163, ZN => n5442);
   U2696 : BUF_X1 port map( A => n15284, Z => n19848);
   U740 : BUF_X1 port map( A => n14829, Z => n19984);
   U62 : XNOR2_X2 port map( A => Key(10), B => Plaintext(10), ZN => n4125);
   U820 : BUF_X2 port map( A => n5031, Z => n153);
   U772 : OAI22_X2 port map( A1 => n3259, A2 => n4694, B1 => n5107, B2 => n4695
                           , ZN => n6183);
   U231 : BUF_X1 port map( A => n3846, Z => n5116);
   U658 : XNOR2_X2 port map( A => n3945, B => Key(181), ZN => n4313);
   U561 : BUF_X1 port map( A => n14120, Z => n14703);
   U440 : XNOR2_X2 port map( A => Key(9), B => Plaintext(9), ZN => n4319);
   U1677 : OR2_X2 port map( A1 => n7175, A2 => n7174, ZN => n9842);
   U852 : NOR2_X2 port map( A1 => n11728, A2 => n682, ZN => n13248);
   U2893 : AND3_X2 port map( A1 => n728, A2 => n14546, A3 => n14545, ZN => 
                           n15645);
   U173 : NAND2_X2 port map( A1 => n1586, A2 => n4218, ZN => n6016);
   U2318 : AND3_X2 port map( A1 => n1815, A2 => n1816, A3 => n1818, ZN => 
                           n15979);
   U957 : BUF_X2 port map( A => n17831, Z => n19110);
   U371 : BUF_X1 port map( A => n6404, Z => n6707);
   U2532 : NOR2_X1 port map( A1 => n14278, A2 => n1409, ZN => n15536);
   U689 : BUF_X2 port map( A => n13316, Z => n14705);
   U6855 : MUX2_X2 port map( A => n17975, B => n17974, S => n17549, Z => n18688
                           );
   U717 : AND2_X2 port map( A1 => n8320, A2 => n8319, ZN => n8872);
   U166 : NAND2_X2 port map( A1 => n15901, A2 => n15902, ZN => n16283);
   U9269 : AND3_X2 port map( A1 => n6212, A2 => n7628, A3 => n6211, ZN => n8708
                           );
   U2909 : BUF_X2 port map( A => n14849, Z => n15474);
   U1008 : OR2_X2 port map( A1 => n2303, A2 => n7858, ZN => n9266);
   U1680 : AND3_X2 port map( A1 => n16050, A2 => n3147, A3 => n3146, ZN => 
                           n16373);
   U408 : XNOR2_X2 port map( A => n4053, B => Key(129), ZN => n4100);
   U1393 : AND2_X2 port map( A1 => n20163, A2 => n20164, ZN => n19227);
   U168 : BUF_X2 port map( A => n13563, Z => n15121);
   U1281 : BUF_X1 port map( A => n13227, Z => n20226);
   U8331 : NAND3_X2 port map( A1 => n1877, A2 => n1997, A3 => n1998, ZN => 
                           n17335);
   U1835 : XNOR2_X2 port map( A => n10135, B => n10136, ZN => n11349);
   U207 : OR2_X2 port map( A1 => n8128, A2 => n6438, ZN => n8129);
   U568 : NAND2_X2 port map( A1 => n2635, A2 => n7452, ZN => n8672);
   U310 : BUF_X1 port map( A => n10882, Z => n11569);
   U1097 : BUF_X2 port map( A => n17374, Z => n18262);
   U687 : XNOR2_X2 port map( A => Key(116), B => Plaintext(116), ZN => n5046);
   U3679 : NAND3_X2 port map( A1 => n3598, A2 => n3453, A3 => n4451, ZN => 
                           n5859);
   U2314 : NAND3_X2 port map( A1 => n1455, A2 => n1454, A3 => n6001, ZN => 
                           n6982);
   U1678 : OAI22_X2 port map( A1 => n8336, A2 => n8335, B1 => n8334, B2 => 
                           n8333, ZN => n9648);
   U501 : OR2_X2 port map( A1 => n15426, A2 => n14243, ZN => n15421);
   U18376 : BUF_X1 port map( A => n16690, Z => n19820);
   U18733 : OAI21_X2 port map( B1 => n18102, B2 => n18101, A => n18100, ZN => 
                           n18651);
   U4237 : NAND2_X2 port map( A1 => n2789, A2 => n3275, ZN => n15546);
   U6938 : OAI22_X2 port map( A1 => n2973, A2 => n15553, B1 => n15552, B2 => 
                           n15551, ZN => n17359);
   U2720 : XNOR2_X2 port map( A => n16848, B => n16849, ZN => n18269);
   U877 : AND3_X2 port map( A1 => n715, A2 => n2380, A3 => n714, ZN => n17438);
   U2955 : OR2_X2 port map( A1 => n7987, A2 => n7986, ZN => n9166);
   U6265 : NAND2_X2 port map( A1 => n8120, A2 => n900, ZN => n9331);
   U1461 : XNOR2_X2 port map( A => n11852, B => n11851, ZN => n15313);
   U6898 : AND2_X2 port map( A1 => n3248, A2 => n18254, ZN => n18774);
   U1839 : BUF_X1 port map( A => n7133, Z => n899);
   U9825 : MUX2_X2 port map( A => n5263, B => n5262, S => n5691, Z => n6520);
   U225 : BUF_X1 port map( A => n15777, Z => n19977);
   U368 : INV_X1 port map( A => n13937, ZN => n14419);
   U13323 : XNOR2_X2 port map( A => n10292, B => n10293, ZN => n11257);
   U387 : AOI22_X2 port map( A1 => n15367, A2 => n15366, B1 => n15369, B2 => 
                           n15368, ZN => n17127);
   U5587 : NAND2_X2 port map( A1 => n780, A2 => n19574, ZN => n18795);
   U1568 : OAI21_X2 port map( B1 => n11355, B2 => n11354, A => n11353, ZN => 
                           n3260);
   U1499 : AND3_X2 port map( A1 => n3464, A2 => n1008, A3 => n11758, ZN => 
                           n13717);
   U746 : BUF_X2 port map( A => n5782, Z => n6055);
   U18737 : NAND2_X2 port map( A1 => n18110, A2 => n18109, ZN => n18648);
   U19 : OAI21_X2 port map( B1 => n4159, B2 => n4158, A => n4157, ZN => n5641);
   U410 : OR2_X2 port map( A1 => n623, A2 => n3833, ZN => n3855);
   U7843 : XNOR2_X2 port map( A => n7085, B => n7084, ZN => n8014);
   U13645 : BUF_X1 port map( A => n19092, Z => n19112);
   U885 : XNOR2_X2 port map( A => n10386, B => n10385, ZN => n11131);
   U19679 : BUF_X1 port map( A => n17300, Z => n19929);
   U679 : NAND3_X2 port map( A1 => n5306, A2 => n5307, A3 => n5305, ZN => n6687
                           );
   U15436 : MUX2_X2 port map( A => n13461, B => n13460, S => n15666, Z => 
                           n17291);
   U653 : BUF_X2 port map( A => n9009, Z => n19490);
   U447 : BUF_X1 port map( A => n5264, Z => n6139);
   U1108 : XNOR2_X2 port map( A => n17292, B => n3207, ZN => n18240);
   U6588 : AOI22_X2 port map( A1 => n2680, A2 => n10895, B1 => n10893, B2 => 
                           n10894, ZN => n12600);
   U11987 : NOR2_X2 port map( A1 => n8491, A2 => n8490, ZN => n10442);
   U51 : CLKBUF_X3 port map( A => n6871, Z => n8272);
   U622 : XNOR2_X2 port map( A => n7947, B => n7946, ZN => n11161);
   U15269 : OAI21_X2 port map( B1 => n15311, B2 => n14992, A => n14991, ZN => 
                           n16227);
   U1849 : AND2_X2 port map( A1 => n1323, A2 => n1322, ZN => n9799);
   U2655 : NAND2_X2 port map( A1 => n579, A2 => n14835, ZN => n17295);
   U12023 : OAI211_X2 port map( C1 => n14813, C2 => n2808, A => n14592, B => 
                           n14591, ZN => n15601);
   U7950 : AOI21_X2 port map( B1 => n14521, B2 => n13565, A => n13564, ZN => 
                           n15052);
   U232 : BUF_X1 port map( A => n15777, Z => n19978);
   U1740 : NAND3_X2 port map( A1 => n4798, A2 => n2699, A3 => n19544, ZN => 
                           n5990);
   U284 : NAND4_X2 port map( A1 => n14141, A2 => n14140, A3 => n3006, A4 => 
                           n3005, ZN => n15510);
   U1075 : XNOR2_X1 port map( A => n12995, B => n12994, ZN => n951);
   U4800 : NOR2_X2 port map( A1 => n8082, A2 => n8081, ZN => n8866);
   U24 : AND3_X2 port map( A1 => n12613, A2 => n12612, A3 => n12611, ZN => 
                           n13518);
   U240 : BUF_X1 port map( A => n6381, Z => n19475);
   U1856 : NAND2_X2 port map( A1 => n5702, A2 => n5701, ZN => n7332);
   U6385 : XNOR2_X2 port map( A => n16826, B => n16827, ZN => n18033);
   U9565 : NAND2_X2 port map( A1 => n350, A2 => n349, ZN => n16330);
   U6697 : OR2_X2 port map( A1 => n8463, A2 => n8462, ZN => n9329);
   U11377 : INV_X1 port map( A => n7453, ZN => n8297);
   U1064 : NAND3_X2 port map( A1 => n1824, A2 => n14606, A3 => n14607, ZN => 
                           n15274);
   U1397 : AND2_X1 port map( A1 => n15311, A2 => n360, ZN => n15399);
   U5362 : MUX2_X2 port map( A => n15027, B => n15026, S => n16629, Z => n18425
                           );
   U889 : BUF_X2 port map( A => n14347, Z => n19496);
   U11912 : XNOR2_X2 port map( A => n8397, B => n8398, ZN => n11159);
   U868 : OAI21_X2 port map( B1 => n1554, B2 => n15561, A => n1553, ZN => 
                           n17407);
   U526 : NAND2_X2 port map( A1 => n11780, A2 => n11779, ZN => n13601);
   U287 : XNOR2_X2 port map( A => n10278, B => n10277, ZN => n11253);
   U8146 : BUF_X1 port map( A => n18151, Z => n19060);
   U1824 : XNOR2_X2 port map( A => n7001, B => n7000, ZN => n7974);
   U1052 : BUF_X2 port map( A => n16447, Z => n17155);
   U1795 : BUF_X1 port map( A => n7571, Z => n8151);
   U463 : BUF_X2 port map( A => n6578, Z => n8239);
   U1307 : AOI21_X2 port map( B1 => n16726, B2 => n20127, A => n16725, ZN => 
                           n870);
   U17460 : BUF_X1 port map( A => n16673, Z => n20244);
   U1192 : CLKBUF_X1 port map( A => Key(144), Z => n456);
   U828 : XNOR2_X1 port map( A => Key(121), B => Plaintext(121), ZN => n4769);
   U1223 : CLKBUF_X1 port map( A => Key(82), Z => n2023);
   U8741 : XNOR2_X1 port map( A => Key(20), B => Plaintext(20), ZN => n4928);
   U8912 : XNOR2_X1 port map( A => Key(43), B => Plaintext(43), ZN => n4968);
   U8918 : XNOR2_X1 port map( A => Key(46), B => Plaintext(46), ZN => n4965);
   U921 : XNOR2_X1 port map( A => Key(14), B => Plaintext(14), ZN => n4306);
   U1376 : CLKBUF_X1 port map( A => Key(69), Z => n17544);
   U1370 : CLKBUF_X1 port map( A => Key(103), Z => n17535);
   U101 : XNOR2_X1 port map( A => Key(154), B => Plaintext(154), ZN => n4756);
   U1371 : CLKBUF_X1 port map( A => Key(30), Z => n2349);
   U1357 : CLKBUF_X1 port map( A => Key(167), Z => n17095);
   U1355 : CLKBUF_X1 port map( A => Key(88), Z => n20064);
   U971 : XNOR2_X1 port map( A => Key(118), B => Plaintext(118), ZN => n5045);
   U605 : BUF_X1 port map( A => n4638, Z => n19524);
   U8871 : XNOR2_X1 port map( A => n3939, B => Key(178), ZN => n4185);
   U322 : BUF_X1 port map( A => n4056, Z => n5058);
   U8499 : BUF_X1 port map( A => n4100, Z => n5060);
   U1717 : AND2_X1 port map( A1 => n1390, A2 => n1389, ZN => n3351);
   U445 : AND2_X1 port map( A1 => n3891, A2 => n3890, ZN => n5300);
   U1925 : OR2_X1 port map( A1 => n4374, A2 => n4373, ZN => n5715);
   U433 : AND2_X1 port map( A1 => n614, A2 => n4639, ZN => n5743);
   U1138 : OR2_X1 port map( A1 => n3976, A2 => n3975, ZN => n6072);
   U6578 : OR2_X1 port map( A1 => n4448, A2 => n4447, ZN => n5860);
   U1934 : NAND2_X1 port map( A1 => n3853, A2 => n306, ZN => n6057);
   U9650 : MUX2_X1 port map( A => n5008, B => n5007, S => n5006, Z => n5009);
   U1924 : AND2_X1 port map( A1 => n5051, A2 => n5050, ZN => n5926);
   U9643 : NAND2_X1 port map( A1 => n2480, A2 => n3641, ZN => n5226);
   U438 : OR2_X1 port map( A1 => n4074, A2 => n4075, ZN => n5434);
   U1929 : AND3_X1 port map( A1 => n4024, A2 => n4023, A3 => n4022, ZN => n5251
                           );
   U9134 : NAND2_X1 port map( A1 => n4155, A2 => n4154, ZN => n5443);
   U479 : AND2_X1 port map( A1 => n4991, A2 => n4990, ZN => n5562);
   U683 : NAND2_X1 port map( A1 => n3399, A2 => n964, ZN => n5279);
   U682 : NAND2_X1 port map( A1 => n2739, A2 => n5015, ZN => n5328);
   U1920 : AND2_X1 port map( A1 => n4774, A2 => n4773, ZN => n6107);
   U1899 : OR2_X1 port map( A1 => n4934, A2 => n4933, ZN => n5683);
   U861 : NAND2_X1 port map( A1 => n1942, A2 => n4906, ZN => n5684);
   U19769 : NAND2_X1 port map( A1 => n20301, A2 => n20017, ZN => n6059);
   U357 : NAND3_X1 port map( A1 => n4014, A2 => n1534, A3 => n1533, ZN => n5393
                           );
   U9056 : OAI211_X1 port map( C1 => n4712, C2 => n4783, A => n4070, B => n4069
                           , ZN => n5997);
   U9781 : AND2_X1 port map( A1 => n5220, A2 => n5219, ZN => n5945);
   U910 : BUF_X1 port map( A => n6167, Z => n170);
   U9672 : BUF_X1 port map( A => n5914, Z => n5916);
   U8273 : AND2_X1 port map( A1 => n3684, A2 => n4386, ZN => n6150);
   U2436 : NAND2_X1 port map( A1 => n4068, A2 => n4067, ZN => n5998);
   U218 : NAND2_X1 port map( A1 => n1768, A2 => n1769, ZN => n3569);
   U1986 : BUF_X1 port map( A => n5304, Z => n5891);
   U1882 : INV_X1 port map( A => n5622, ZN => n5621);
   U10105 : MUX2_X1 port map( A => n5672, B => n5671, S => n5670, Z => n5679);
   U261 : OAI211_X1 port map( C1 => n6014, C2 => n6013, A => n6012, B => n6011,
                           ZN => n6990);
   U2196 : NAND3_X1 port map( A1 => n5066, A2 => n5065, A3 => n20036, ZN => 
                           n7373);
   U6935 : OR2_X1 port map( A1 => n5198, A2 => n5197, ZN => n6641);
   U19710 : AOI22_X1 port map( A1 => n6160, A2 => n5614, B1 => n5613, B2 => 
                           n5612, ZN => n7297);
   U1998 : NAND2_X1 port map( A1 => n1435, A2 => n1170, ZN => n7196);
   U5200 : NAND3_X1 port map( A1 => n1871, A2 => n1870, A3 => n5451, ZN => 
                           n7289);
   U1863 : NAND3_X1 port map( A1 => n2639, A2 => n6053, A3 => n2638, ZN => 
                           n7018);
   U727 : OAI21_X1 port map( B1 => n4779, B2 => n5640, A => n4778, ZN => n7336)
                           ;
   U1868 : OAI211_X1 port map( C1 => n5462, C2 => n1867, A => n5461, B => n5460
                           , ZN => n7160);
   U1343 : OR2_X1 port map( A1 => n5195, A2 => n5194, ZN => n6776);
   U10304 : XNOR2_X1 port map( A => n7116, B => n7354, ZN => n6718);
   U1843 : NAND2_X1 port map( A1 => n5482, A2 => n5481, ZN => n7306);
   U4673 : AOI21_X1 port map( B1 => n5183, B2 => n5182, A => n5181, ZN => n7273
                           );
   U6805 : XNOR2_X1 port map( A => n5134, B => n5133, ZN => n8184);
   U854 : XNOR2_X1 port map( A => n6332, B => n6331, ZN => n7739);
   U791 : XNOR2_X1 port map( A => n7037, B => n7038, ZN => n7958);
   U7402 : XNOR2_X1 port map( A => n2825, B => n2824, ZN => n8370);
   U9506 : XNOR2_X1 port map( A => n4728, B => n4729, ZN => n8190);
   U1792 : BUF_X1 port map( A => n6837, Z => n7852);
   U11473 : INV_X1 port map( A => n7542, ZN => n8372);
   U663 : BUF_X1 port map( A => n7684, Z => n8381);
   U2104 : XNOR2_X1 port map( A => n5491, B => n5490, ZN => n8034);
   U504 : XNOR2_X1 port map( A => n6357, B => n6356, ZN => n7500);
   U50 : CLKBUF_X1 port map( A => n7481, Z => n7949);
   U1782 : BUF_X1 port map( A => n7493, Z => n7679);
   U773 : BUF_X1 port map( A => n7487, Z => n7968);
   U898 : XNOR2_X1 port map( A => n5377, B => n5376, ZN => n7445);
   U18094 : BUF_X1 port map( A => n7621, Z => n8069);
   U540 : OAI211_X1 port map( C1 => n2875, C2 => n7893, A => n7892, B => n7607,
                           ZN => n8729);
   U89 : OAI211_X1 port map( C1 => n1411, C2 => n1010, A => n7617, B => n1410, 
                           ZN => n8743);
   U2559 : OAI22_X1 port map( A1 => n7468, A2 => n8289, B1 => n8024, B2 => 
                           n8292, ZN => n8294);
   U8530 : OAI211_X1 port map( C1 => n7835, C2 => n7773, A => n7772, B => n7771
                           , ZN => n8997);
   U916 : NOR2_X1 port map( A1 => n6909, A2 => n6910, ZN => n8611);
   U1739 : NAND2_X1 port map( A1 => n6901, A2 => n6902, ZN => n9158);
   U451 : OAI211_X1 port map( C1 => n8050, C2 => n8309, A => n8049, B => n8048,
                           ZN => n9066);
   U6587 : INV_X1 port map( A => n8542, ZN => n9836);
   U234 : BUF_X1 port map( A => n8748, Z => n8931);
   U100 : OAI21_X1 port map( B1 => n7784, B2 => n7783, A => n7782, ZN => n9177)
                           ;
   U46 : AND3_X1 port map( A1 => n2251, A2 => n2252, A3 => n1784, ZN => n9149);
   U441 : NAND2_X1 port map( A1 => n8275, A2 => n8274, ZN => n9129);
   U1111 : NAND3_X1 port map( A1 => n2190, A2 => n2191, A3 => n6586, ZN => 
                           n6587);
   U280 : AND2_X1 port map( A1 => n7437, A2 => n2986, ZN => n9296);
   U1704 : AND2_X1 port map( A1 => n1657, A2 => n7810, ZN => n9006);
   U1718 : BUF_X1 port map( A => n8500, Z => n9361);
   U435 : NAND3_X1 port map( A1 => n7419, A2 => n429, A3 => n428, ZN => n9300);
   U908 : NOR2_X1 port map( A1 => n7545, A2 => n7546, ZN => n8959);
   U12626 : BUF_X1 port map( A => n5556, Z => n19716);
   U1903 : NAND2_X1 port map( A1 => n7706, A2 => n20293, ZN => n8974);
   U453 : AND2_X1 port map( A1 => n7734, A2 => n7735, ZN => n9249);
   U5590 : NAND2_X1 port map( A1 => n1158, A2 => n1160, ZN => n7866);
   U5242 : NAND2_X1 port map( A1 => n1422, A2 => n1839, ZN => n9528);
   U1700 : AND2_X1 port map( A1 => n9137, A2 => n8445, ZN => n9134);
   U449 : OR2_X1 port map( A1 => n8698, A2 => n9163, ZN => n8613);
   U378 : MUX2_X1 port map( A => n7842, B => n7841, S => n8623, Z => n9420);
   U315 : AND2_X1 port map( A1 => n19596, A2 => n19595, ZN => n9862);
   U413 : OAI211_X1 port map( C1 => n8947, C2 => n7613, A => n7612, B => n7611,
                           ZN => n10054);
   U297 : NAND2_X1 port map( A1 => n8447, A2 => n8448, ZN => n10303);
   U1109 : OR2_X1 port map( A1 => n2746, A2 => n2747, ZN => n8593);
   U9119 : OAI211_X1 port map( C1 => n9451, C2 => n9094, A => n9093, B => n9092
                           , ZN => n10027);
   U857 : OAI21_X1 port map( B1 => n1255, B2 => n1257, A => n1254, ZN => n9697)
                           ;
   U1689 : OR2_X1 port map( A1 => n1738, A2 => n1737, ZN => n9600);
   U756 : OAI21_X1 port map( B1 => n8523, B2 => n8522, A => n8521, ZN => n10551
                           );
   U3170 : OAI211_X1 port map( C1 => n8866, C2 => n8869, A => n8123, B => n8122
                           , ZN => n10271);
   U467 : NAND3_X1 port map( A1 => n1766, A2 => n8038, A3 => n8039, ZN => 
                           n10270);
   U400 : MUX2_X1 port map( A => n9223, B => n9222, S => n1428, Z => n10473);
   U928 : OAI21_X1 port map( B1 => n8587, B2 => n8588, A => n2351, ZN => n10367
                           );
   U320 : NAND2_X1 port map( A1 => n8465, A2 => n8464, ZN => n10557);
   U2099 : NAND2_X1 port map( A1 => n9044, A2 => n1932, ZN => n10046);
   U2674 : INV_X1 port map( A => n10598, ZN => n10514);
   U476 : OR2_X1 port map( A1 => n8863, A2 => n8864, ZN => n9391);
   U44 : OR2_X1 port map( A1 => n9584, A2 => n9583, ZN => n1032);
   U1867 : AOI21_X1 port map( B1 => n8976, B2 => n8977, A => n8975, ZN => n9692
                           );
   U249 : OAI21_X1 port map( B1 => n9027, B2 => n9026, A => n9025, ZN => n10558
                           );
   U13694 : XNOR2_X1 port map( A => n9798, B => n9797, ZN => n11267);
   U1651 : XNOR2_X1 port map( A => n8821, B => n8822, ZN => n11170);
   U1079 : XNOR2_X1 port map( A => n10538, B => n10539, ZN => n11186);
   U983 : XNOR2_X1 port map( A => n8536, B => n8535, ZN => n11528);
   U157 : XNOR2_X1 port map( A => n550, B => n9859, ZN => n9883);
   U303 : XNOR2_X1 port map( A => n9708, B => n9707, ZN => n11330);
   U8787 : BUF_X1 port map( A => n11240, Z => n10798);
   U829 : XNOR2_X1 port map( A => n9541, B => n9540, ZN => n11142);
   U13456 : XNOR2_X1 port map( A => n10520, B => n10521, ZN => n11035);
   U364 : BUF_X1 port map( A => n9545, Z => n937);
   U52 : XNOR2_X1 port map( A => n10460, B => n10459, ZN => n10845);
   U505 : BUF_X1 port map( A => n10060, Z => n11480);
   U19745 : BUF_X1 port map( A => n10742, Z => n10936);
   U890 : BUF_X1 port map( A => n11104, Z => n11041);
   U17 : OR2_X1 port map( A1 => n10966, A2 => n3361, ZN => n12220);
   U398 : OAI211_X1 port map( C1 => n11282, C2 => n10695, A => n1847, B => 
                           n1848, ZN => n180);
   U14071 : MUX2_X1 port map( A => n11537, B => n11536, S => n11535, Z => 
                           n11543);
   U331 : OAI21_X1 port map( B1 => n9747, B2 => n9746, A => n9745, ZN => n12009
                           );
   U238 : OR2_X1 port map( A1 => n12552, A2 => n12548, ZN => n12542);
   U639 : NAND2_X1 port map( A1 => n10759, A2 => n2522, ZN => n2523);
   U3573 : NOR2_X1 port map( A1 => n10857, A2 => n11378, ZN => n2606);
   U1559 : AOI21_X1 port map( B1 => n1498, B2 => n1497, A => n606, ZN => n11841
                           );
   U845 : AND2_X1 port map( A1 => n9973, A2 => n2704, ZN => n12005);
   U1574 : AND2_X1 port map( A1 => n1804, A2 => n11453, ZN => n12460);
   U1567 : AND2_X1 port map( A1 => n11252, A2 => n1599, ZN => n12381);
   U844 : INV_X1 port map( A => n12005, ZN => n201);
   U1533 : AND2_X1 port map( A1 => n3613, A2 => n3616, ZN => n11977);
   U661 : NAND2_X1 port map( A1 => n10067, A2 => n1418, ZN => n12499);
   U8172 : NAND2_X1 port map( A1 => n11517, A2 => n11518, ZN => n12533);
   U1540 : AND3_X1 port map( A1 => n3630, A2 => n965, A3 => n3629, ZN => n12338
                           );
   U1563 : AOI21_X1 port map( B1 => n11498, B2 => n11497, A => n11496, ZN => 
                           n12162);
   U527 : NOR2_X1 port map( A1 => n12207, A2 => n12208, ZN => n12065);
   U1090 : NAND2_X1 port map( A1 => n10669, A2 => n1917, ZN => n12443);
   U564 : CLKBUF_X1 port map( A => n12631, Z => n20184);
   U2888 : AND2_X2 port map( A1 => n724, A2 => n721, ZN => n12500);
   U2198 : NAND2_X1 port map( A1 => n371, A2 => n373, ZN => n12502);
   U18272 : OR3_X1 port map( A1 => n12595, A2 => n12589, A3 => n12202, ZN => 
                           n12203);
   U35 : OAI21_X1 port map( B1 => n10837, B2 => n10836, A => n10835, ZN => 
                           n12200);
   U2771 : NOR2_X1 port map( A1 => n12374, A2 => n12269, ZN => n12377);
   U967 : NAND2_X1 port map( A1 => n313, A2 => n3480, ZN => n12537);
   U8432 : OR3_X1 port map( A1 => n12338, A2 => n12336, A3 => n12335, ZN => 
                           n12343);
   U11582 : BUF_X1 port map( A => n13702, Z => n20155);
   U414 : OAI21_X1 port map( B1 => n12134, B2 => n11590, A => n11589, ZN => 
                           n13425);
   U25 : AND3_X1 port map( A1 => n513, A2 => n512, A3 => n33, ZN => n13018);
   U853 : AOI21_X1 port map( B1 => n12052, B2 => n12051, A => n12050, ZN => 
                           n13260);
   U14726 : OAI211_X1 port map( C1 => n11807, C2 => n12537, A => n11806, B => 
                           n11805, ZN => n19892);
   U1504 : NOR2_X1 port map( A1 => n9622, A2 => n9621, ZN => n12696);
   U1503 : NOR2_X1 port map( A1 => n11858, A2 => n11857, ZN => n12471);
   U5499 : OR2_X1 port map( A1 => n12432, A2 => n12431, ZN => n12433);
   U2769 : MUX2_X1 port map( A => n12239, B => n12238, S => n12606, Z => n13755
                           );
   U535 : NAND3_X1 port map( A1 => n3631, A2 => n3633, A3 => n11601, ZN => 
                           n13368);
   U109 : AND3_X1 port map( A1 => n588, A2 => n1116, A3 => n1117, ZN => n13042)
                           ;
   U1522 : AND2_X1 port map( A1 => n1258, A2 => n1224, ZN => n1260);
   U426 : MUX2_X1 port map( A => n11584, B => n11583, S => n12040, Z => n12863)
                           ;
   U4524 : AOI22_X1 port map( A1 => n12502, A2 => n12503, B1 => n12501, B2 => 
                           n201, ZN => n13468);
   U14123 : OAI211_X1 port map( C1 => n11617, C2 => n11616, A => n11615, B => 
                           n11614, ZN => n13774);
   U1784 : MUX2_X1 port map( A => n11678, B => n11677, S => n11820, Z => n13687
                           );
   U2381 : NAND2_X1 port map( A1 => n458, A2 => n11723, ZN => n13517);
   U3612 : OAI21_X1 port map( B1 => n12610, B2 => n11630, A => n3761, ZN => 
                           n13580);
   U236 : AND2_X1 port map( A1 => n19557, A2 => n19555, ZN => n13643);
   U91 : XNOR2_X1 port map( A => n3364, B => n3363, ZN => n14663);
   U886 : XNOR2_X1 port map( A => n13487, B => n13488, ZN => n14747);
   U992 : XNOR2_X1 port map( A => n13084, B => n13083, ZN => n15120);
   U48 : XNOR2_X1 port map( A => n11715, B => n11716, ZN => n14593);
   U811 : XNOR2_X1 port map( A => n13220, B => n13219, ZN => n14547);
   U17534 : XNOR2_X1 port map( A => n13593, B => n13594, ZN => n14394);
   U1444 : BUF_X1 port map( A => n14388, Z => n14723);
   U3282 : OAI21_X1 port map( B1 => n14307, B2 => n14499, A => n3034, ZN => 
                           n13975);
   U9597 : MUX2_X1 port map( A => n14794, B => n14793, S => n2412, Z => n15815)
                           ;
   U1781 : OAI21_X1 port map( B1 => n14174, B2 => n774, A => n14173, ZN => 
                           n15309);
   U2442 : AND4_X1 port map( A1 => n3245, A2 => n3244, A3 => n2839, A4 => 
                           n13016, ZN => n15684);
   U4983 : AND3_X1 port map( A1 => n1292, A2 => n1294, A3 => n1024, ZN => 
                           n15898);
   U9571 : NAND2_X1 port map( A1 => n1625, A2 => n1624, ZN => n15551);
   U596 : AND3_X1 port map( A1 => n2775, A2 => n2774, A3 => n2773, ZN => n15187
                           );
   U3071 : BUF_X1 port map( A => n15341, Z => n19888);
   U119 : CLKBUF_X1 port map( A => n14902, Z => n20147);
   U216 : NAND3_X1 port map( A1 => n3539, A2 => n3538, A3 => n14080, ZN => 
                           n15521);
   U247 : NAND3_X1 port map( A1 => n14008, A2 => n36, A3 => n35, ZN => n15698);
   U591 : BUF_X1 port map( A => n14997, Z => n15257);
   U2573 : NOR2_X1 port map( A1 => n13683, A2 => n530, ZN => n15228);
   U3104 : OAI21_X1 port map( B1 => n14025, B2 => n2626, A => n14024, ZN => 
                           n15754);
   U16201 : NOR2_X2 port map( A1 => n20182, A2 => n15803, ZN => n15802);
   U3125 : NOR2_X1 port map( A1 => n15819, A2 => n2114, ZN => n17110);
   U15730 : NAND2_X1 port map( A1 => n13917, A2 => n13916, ZN => n16931);
   U1280 : AND2_X1 port map( A1 => n3103, A2 => n14900, ZN => n17377);
   U16292 : XNOR2_X1 port map( A => n14885, B => n14884, ZN => n17210);
   U11687 : XNOR2_X1 port map( A => n16986, B => n16985, ZN => n18025);
   U1331 : BUF_X1 port map( A => n19737, Z => n18103);
   U990 : OR2_X1 port map( A1 => n17654, A2 => n20004, ZN => n19399);
   U86 : AOI21_X1 port map( B1 => n17516, B2 => n17515, A => n17514, ZN => 
                           n18512);
   U1224 : OR2_X1 port map( A1 => n1712, A2 => n3485, ZN => n18376);
   U1565 : NOR2_X1 port map( A1 => n17675, A2 => n17674, ZN => n19278);
   U19528 : AOI22_X1 port map( A1 => n19406, A2 => n19405, B1 => n19403, B2 => 
                           n19404, ZN => n19432);
   U1041 : OAI211_X1 port map( C1 => n19400, C2 => n19399, A => n19398, B => 
                           n19397, ZN => n19441);
   U1294 : OR2_X1 port map( A1 => n18117, A2 => n18116, ZN => n18634);
   U204 : AND2_X1 port map( A1 => n17659, A2 => n17658, ZN => n19246);
   U19739 : NAND3_X1 port map( A1 => n17722, A2 => n17721, A3 => n17720, ZN => 
                           n19032);
   U18641 : AND3_X1 port map( A1 => n17963, A2 => n17962, A3 => n17961, ZN => 
                           n18671);
   U256 : NAND2_X1 port map( A1 => n17560, A2 => n18211, ZN => n18625);
   U3061 : NOR2_X1 port map( A1 => n19283, A2 => n19282, ZN => n19304);
   U758 : NAND3_X4 port map( A1 => n5885, A2 => n2928, A3 => n4057, ZN => n6046
                           );
   U7690 : OR2_X1 port map( A1 => n4550, A2 => n3094, ZN => n5768);
   U6884 : INV_X1 port map( A => n7862, ZN => n3775);
   U2538 : CLKBUF_X1 port map( A => n8060, Z => n7893);
   U1759 : AND3_X1 port map( A1 => n7876, A2 => n7599, A3 => n7598, ZN => n8945
                           );
   U411 : INV_X2 port map( A => n9151, ZN => n9145);
   U7986 : INV_X1 port map( A => n9291, ZN => n9579);
   U12080 : INV_X2 port map( A => n8596, ZN => n8933);
   U1708 : BUF_X1 port map( A => n8419, Z => n9137);
   U973 : INV_X1 port map( A => n11290, ZN => n19506);
   U13915 : INV_X1 port map( A => n12280, ZN => n12040);
   U734 : NAND3_X1 port map( A1 => n1315, A2 => n1318, A3 => n1314, ZN => 
                           n12642);
   U6827 : NAND2_X1 port map( A1 => n12785, A2 => n12784, ZN => n13312);
   U1062 : NOR2_X1 port map( A1 => n2806, A2 => n13890, ZN => n15857);
   U516 : AND2_X2 port map( A1 => n6361, A2 => n6360, ZN => n8884);
   U308 : NOR2_X2 port map( A1 => n14317, A2 => n14318, ZN => n14903);
   U5498 : OR2_X2 port map( A1 => n12433, A2 => n1550, ZN => n13747);
   U690 : AND2_X2 port map( A1 => n3850, A2 => n3849, ZN => n6064);
   U8110 : OR2_X2 port map( A1 => n8909, A2 => n8908, ZN => n8917);
   U4285 : MUX2_X2 port map( A => n7955, B => n7954, S => n7953, Z => n9167);
   U1427 : AND3_X2 port map( A1 => n18236, A2 => n18235, A3 => n18234, ZN => 
                           n18762);
   U513 : NAND3_X2 port map( A1 => n662, A2 => n4556, A3 => n661, ZN => n5802);
   U99 : AND2_X2 port map( A1 => n20027, A2 => n20026, ZN => n12429);
   U191 : AND2_X2 port map( A1 => n760, A2 => n761, ZN => n5201);
   U831 : XNOR2_X2 port map( A => n6399, B => n6400, ZN => n8365);
   U524 : NAND2_X2 port map( A1 => n3407, A2 => n5521, ZN => n6736);
   U1654 : AND2_X2 port map( A1 => n2617, A2 => n969, ZN => n10105);
   U624 : OAI211_X2 port map( C1 => n12388, C2 => n12470, A => n1946, B => 
                           n1945, ZN => n12992);
   U637 : OR2_X2 port map( A1 => n3332, A2 => n3331, ZN => n15007);
   U1923 : NAND2_X2 port map( A1 => n20292, A2 => n667, ZN => n670);
   U495 : OR2_X2 port map( A1 => n11740, A2 => n11744, ZN => n12274);
   U11214 : XNOR2_X2 port map( A => n7192, B => n7191, ZN => n8315);
   U878 : AND3_X2 port map( A1 => n2150, A2 => n8835, A3 => n8834, ZN => n9934)
                           ;
   U672 : XNOR2_X2 port map( A => Key(147), B => Plaintext(147), ZN => n4204);
   U617 : BUF_X2 port map( A => n17758, Z => n18753);
   U19616 : AOI21_X2 port map( B1 => n12276, B2 => n12300, A => n1872, ZN => 
                           n19883);
   U10046 : INV_X2 port map( A => n5556, ZN => n8411);
   U869 : AND3_X2 port map( A1 => n1719, A2 => n1720, A3 => n452, ZN => n5320);
   U18489 : BUF_X2 port map( A => n16743, Z => n20267);
   U18497 : AOI22_X2 port map( A1 => n1682, A2 => n15588, B1 => n14040, B2 => 
                           n15755, ZN => n16743);
   U175 : OR2_X2 port map( A1 => n5121, A2 => n5120, ZN => n5917);
   U2954 : NAND2_X2 port map( A1 => n1825, A2 => n7977, ZN => n8569);
   U104 : OAI211_X2 port map( C1 => n14219, C2 => n3697, A => n14217, B => 
                           n14218, ZN => n15405);
   U4733 : AND4_X2 port map( A1 => n10910, A2 => n10909, A3 => n10908, A4 => 
                           n10907, ZN => n12237);
   U16465 : AOI21_X2 port map( B1 => n15063, B2 => n15064, A => n15062, ZN => 
                           n16690);
   U193 : OAI21_X2 port map( B1 => n11040, B2 => n11039, A => n3459, ZN => 
                           n12261);
   U12047 : BUF_X2 port map( A => n10761, Z => n11544);
   U2636 : NAND3_X2 port map( A1 => n566, A2 => n2866, A3 => n2868, ZN => n657)
                           ;
   U2413 : AND2_X2 port map( A1 => n3251, A2 => n475, ZN => n9564);
   U7561 : NAND2_X2 port map( A1 => n17077, A2 => n1109, ZN => n19165);
   U542 : INV_X2 port map( A => n15495, ZN => n3431);
   U1358 : BUF_X2 port map( A => n14722, Z => n19843);
   U7845 : AND2_X2 port map( A1 => n3289, A2 => n4109, ZN => n5815);
   U5497 : XNOR2_X2 port map( A => n6424, B => n6425, ZN => n7748);
   U860 : OAI211_X2 port map( C1 => n8260, C2 => n8259, A => n8258, B => n8257,
                           ZN => n8276);
   U965 : OR2_X2 port map( A1 => n5414, A2 => n5413, ZN => n7014);
   U882 : BUF_X2 port map( A => n8156, Z => n9338);
   U2351 : OR2_X2 port map( A1 => n12408, A2 => n12389, ZN => n12412);
   U180 : NOR2_X2 port map( A1 => n9382, A2 => n9381, ZN => n10579);
   U1735 : MUX2_X2 port map( A => n8907, B => n8911, S => n8910, Z => n8923);
   U1871 : NAND4_X2 port map( A1 => n4212, A2 => n2718, A3 => n4211, A4 => 
                           n4210, ZN => n6489);
   U855 : BUF_X2 port map( A => n4656, Z => n164);
   U1042 : BUF_X2 port map( A => n18709, Z => n18781);
   U7624 : NAND3_X2 port map( A1 => n9561, A2 => n9562, A3 => n3023, ZN => 
                           n11829);
   U350 : AND3_X2 port map( A1 => n16268, A2 => n16267, A3 => n1248, ZN => 
                           n19208);
   U113 : XNOR2_X2 port map( A => n16723, B => n16722, ZN => n18961);
   U14379 : OAI211_X2 port map( C1 => n11959, C2 => n11958, A => n11957, B => 
                           n11956, ZN => n13736);
   U7643 : NAND2_X2 port map( A1 => n15591, A2 => n15590, ZN => n16928);
   U5813 : OAI211_X2 port map( C1 => n8299, C2 => n5963, A => n19578, B => 
                           n19577, ZN => n9234);
   U1889 : OR2_X2 port map( A1 => n4273, A2 => n4272, ZN => n5622);
   U1484 : AND3_X2 port map( A1 => n17844, A2 => n17843, A3 => n17842, ZN => 
                           n19067);
   U986 : XNOR2_X2 port map( A => Key(67), B => Plaintext(67), ZN => n4840);
   U421 : NAND2_X2 port map( A1 => n2481, A2 => n4884, ZN => n7188);
   U1588 : OR2_X2 port map( A1 => n11248, A2 => n11247, ZN => n12269);
   U450 : INV_X2 port map( A => n13514, ZN => n13397);
   U4825 : MUX2_X2 port map( A => n11676, B => n11675, S => n11674, Z => n13514
                           );
   U16518 : NOR2_X2 port map( A1 => n6188, A2 => n6187, ZN => n6967);
   U1377 : OAI21_X2 port map( B1 => n15419, B2 => n15910, A => n2577, ZN => 
                           n16236);
   U684 : XNOR2_X2 port map( A => Key(12), B => Plaintext(12), ZN => n4982);
   U336 : BUF_X2 port map( A => n6344, Z => n8359);
   U1861 : OAI21_X2 port map( B1 => n5254, B2 => n5367, A => n5253, ZN => n6977
                           );
   U980 : BUF_X2 port map( A => n5117, Z => n19508);
   U1458 : XNOR2_X2 port map( A => n12847, B => n12848, ZN => n14453);
   U2463 : MUX2_X2 port map( A => n10820, B => n10819, S => n11365, Z => n11811
                           );
   U1440 : OR2_X2 port map( A1 => n19442, A2 => n19441, ZN => n19425);
   U1857 : NAND3_X2 port map( A1 => n1563, A2 => n4025, A3 => n1561, ZN => 
                           n6745);
   U2484 : BUF_X2 port map( A => n6702, Z => n8114);
   U1134 : NAND2_X2 port map( A1 => n434, A2 => n432, ZN => n6044);
   U762 : BUF_X2 port map( A => n3897, Z => n4988);
   U1664 : OAI211_X2 port map( C1 => n8683, C2 => n9149, A => n392, B => n391, 
                           ZN => n9777);
   U343 : NAND2_X2 port map( A1 => n2111, A2 => n2110, ZN => n17275);
   U1994 : NOR2_X2 port map( A1 => n5679, A2 => n5678, ZN => n19764);
   U8985 : XNOR2_X2 port map( A => Key(117), B => Plaintext(117), ZN => n4439);
   U11737 : NAND4_X2 port map( A1 => n7941, A2 => n7940, A3 => n7939, A4 => 
                           n7938, ZN => n8786);
   U1734 : NAND2_X2 port map( A1 => n13804, A2 => n67, ZN => n15442);
   U873 : BUF_X2 port map( A => n10048, Z => n19990);
   U865 : MUX2_X2 port map( A => n7401, B => n7400, S => n8026, Z => n8596);
   U335 : BUF_X2 port map( A => n9919, Z => n11219);
   U276 : AND2_X2 port map( A1 => n2859, A2 => n2856, ZN => n12440);
   U1361 : NOR2_X2 port map( A1 => n485, A2 => n11774, ZN => n13539);
   U1928 : NAND3_X2 port map( A1 => n523, A2 => n973, A3 => n4225, ZN => n5825)
                           ;
   U933 : BUF_X1 port map( A => n4686, Z => n176);
   U1466 : XNOR2_X2 port map( A => n13208, B => n13209, ZN => n14656);
   U985 : BUF_X2 port map( A => n11325, Z => n191);
   U15 : BUF_X2 port map( A => n15153, Z => n16015);
   U1300 : AND2_X2 port map( A1 => n15253, A2 => n15254, ZN => n18427);
   U341 : BUF_X2 port map( A => n12973, Z => n14637);
   U1581 : NOR2_X2 port map( A1 => n10994, A2 => n10993, ZN => n12576);
   U4814 : AND3_X2 port map( A1 => n20030, A2 => n3178, A3 => n14054, ZN => 
                           n15266);
   U2315 : XNOR2_X2 port map( A => n2036, B => Key(29), ZN => n4887);
   U1418 : AOI21_X2 port map( B1 => n14538, B2 => n13179, A => n13178, ZN => 
                           n14866);
   U563 : OAI21_X2 port map( B1 => n11262, B2 => n11261, A => n11260, ZN => 
                           n12373);
   U17057 : XNOR2_X2 port map( A => n16028, B => n16029, ZN => n17896);
   U1858 : OR2_X2 port map( A1 => n3936, A2 => n3935, ZN => n6693);
   U18850 : BUF_X2 port map( A => n7115, Z => n6478);
   U430 : CLKBUF_X3 port map( A => n14052, Z => n14359);
   U366 : OR2_X2 port map( A1 => n8422, A2 => n8421, ZN => n1960);
   U701 : NAND2_X2 port map( A1 => n1518, A2 => n1519, ZN => n15577);
   U718 : AND2_X2 port map( A1 => n2930, A2 => n2933, ZN => n9210);
   U676 : AOI21_X2 port map( B1 => n14399, B2 => n14398, A => n14397, ZN => 
                           n15627);
   U599 : AOI21_X2 port map( B1 => n10656, B2 => n2231, A => n3219, ZN => 
                           n12417);
   U833 : XNOR2_X2 port map( A => n8607, B => n8608, ZN => n11550);
   U748 : BUF_X2 port map( A => n17261, Z => n947);
   U1897 : NOR2_X2 port map( A1 => n9002, A2 => n20037, ZN => n10026);
   U1299 : NAND2_X2 port map( A1 => n16451, A2 => n19695, ZN => n18555);
   U3742 : OR2_X2 port map( A1 => n5027, A2 => n5026, ZN => n3309);
   U8495 : OR2_X2 port map( A1 => n4744, A2 => n4745, ZN => n4559);
   U8827 : XNOR2_X2 port map( A => Key(148), B => Plaintext(148), ZN => n4745);
   U590 : AND3_X2 port map( A1 => n14832, A2 => n14831, A3 => n2779, ZN => 
                           n15581);
   U4523 : OR2_X2 port map( A1 => n5408, A2 => n3959, ZN => n5572);
   U5036 : CLKBUF_X2 port map( A => n5005, Z => n4248);
   U1922 : AND2_X1 port map( A1 => n4009, A2 => n4008, ZN => n5395);
   U6914 : MUX2_X1 port map( A => n8089, B => n8088, S => n20254, Z => n9333);
   U801 : BUF_X1 port map( A => n10194, Z => n11265);
   U1623 : BUF_X1 port map( A => n10450, Z => n11202);
   U1596 : INV_X1 port map( A => n10785, ZN => n1039);
   U1825 : OR2_X1 port map( A1 => n11328, A2 => n11244, ZN => n11375);
   U680 : BUF_X2 port map( A => n11563, Z => n11782);
   U5 : BUF_X2 port map( A => n12290, Z => n182);
   U221 : OAI211_X1 port map( C1 => n12082, C2 => n11608, A => n11607, B => 
                           n11606, ZN => n13277);
   U1491 : AND2_X1 port map( A1 => n1509, A2 => n1513, ZN => n13344);
   U1487 : AND3_X1 port map( A1 => n19527, A2 => n852, A3 => n851, ZN => n13126
                           );
   U2456 : BUF_X2 port map( A => n12842, Z => n15336);
   U895 : AND3_X1 port map( A1 => n3644, A2 => n3643, A3 => n15757, ZN => 
                           n15756);
   U2841 : AND3_X1 port map( A1 => n1368, A2 => n14661, A3 => n681, ZN => 
                           n15574);
   U530 : BUF_X1 port map( A => n15994, Z => n17330);
   U4090 : OR2_X1 port map( A1 => n17063, A2 => n17840, ZN => n3287);
   U6 : NAND3_X1 port map( A1 => n2144, A2 => n5779, A3 => n146, ZN => n6839);
   U16 : BUF_X2 port map( A => n4882, Z => n5741);
   U18 : AND3_X2 port map( A1 => n7438, A2 => n20029, A3 => n7440, ZN => n9602)
                           ;
   U23 : MUX2_X2 port map( A => n3208, B => n18237, S => n18240, Z => n3206);
   U27 : NAND2_X2 port map( A1 => n20690, A2 => n1481, ZN => n9922);
   U40 : OR2_X2 port map( A1 => n3563, A2 => n3564, ZN => n6155);
   U42 : NOR2_X2 port map( A1 => n16441, A2 => n16440, ZN => n18567);
   U58 : AND2_X2 port map( A1 => n12037, A2 => n12036, ZN => n11717);
   U67 : NAND2_X2 port map( A1 => n4710, A2 => n20679, ZN => n6184);
   U77 : NOR2_X2 port map( A1 => n12524, A2 => n12167, ZN => n12522);
   U82 : AOI21_X2 port map( B1 => n9133, B2 => n9132, A => n9131, ZN => n19945)
                           ;
   U87 : XNOR2_X2 port map( A => n13441, B => n13442, ZN => n14555);
   U98 : BUF_X2 port map( A => n4868, Z => n20357);
   U108 : NAND2_X2 port map( A1 => n515, A2 => n20649, ZN => n7240);
   U114 : XNOR2_X2 port map( A => n10512, B => n10511, ZN => n11037);
   U126 : AND2_X2 port map( A1 => n2578, A2 => n15906, ZN => n15912);
   U145 : BUF_X2 port map( A => n17935, Z => n18357);
   U148 : OAI21_X1 port map( B1 => n3081, B2 => n17507, A => n3080, ZN => 
                           n18467);
   U159 : XNOR2_X1 port map( A => n15249, B => n19893, ZN => n15968);
   U171 : OAI21_X1 port map( B1 => n11771, B2 => n12292, A => n11770, ZN => 
                           n13255);
   U181 : BUF_X1 port map( A => n7764, Z => n20358);
   U183 : BUF_X1 port map( A => n7764, Z => n20360);
   U192 : OAI211_X1 port map( C1 => n4743, C2 => n5055, A => n4742, B => n4741,
                           ZN => n6104);
   U215 : XNOR2_X1 port map( A => n16877, B => n16876, ZN => n18977);
   U223 : XOR2_X1 port map( A => n7280, B => n7281, Z => n20347);
   U246 : NOR2_X2 port map( A1 => n7429, A2 => n7428, ZN => n9304);
   U260 : XNOR2_X2 port map( A => n10102, B => n10101, ZN => n19949);
   U262 : OR2_X2 port map( A1 => n10983, A2 => n10984, ZN => n11686);
   U263 : AOI22_X2 port map( A1 => n11785, A2 => n11784, B1 => n920, B2 => 
                           n11783, ZN => n13602);
   U268 : XNOR2_X2 port map( A => n2783, B => n2784, ZN => n14818);
   U279 : OAI21_X2 port map( B1 => n14066, B2 => n14065, A => n14064, ZN => 
                           n868);
   U285 : NOR2_X2 port map( A1 => n15144, A2 => n15143, ZN => n19720);
   U296 : BUF_X2 port map( A => n17244, Z => n20354);
   U300 : OAI21_X2 port map( B1 => n19379, B2 => n19733, A => n19378, ZN => 
                           n19439);
   U301 : MUX2_X2 port map( A => n17709, B => n17708, S => n18941, Z => n19047)
                           ;
   U305 : AND2_X2 port map( A1 => n3499, A2 => n10767, ZN => n13617);
   U327 : XNOR2_X2 port map( A => Key(27), B => Plaintext(27), ZN => n4118);
   U332 : XNOR2_X2 port map( A => Key(109), B => Plaintext(109), ZN => n5086);
   U333 : XNOR2_X2 port map( A => n16833, B => n16832, ZN => n18270);
   U339 : XNOR2_X2 port map( A => n11818, B => n11819, ZN => n14627);
   U342 : NAND2_X2 port map( A1 => n578, A2 => n6094, ZN => n7026);
   U344 : XNOR2_X2 port map( A => n3994, B => Key(58), ZN => n4684);
   U346 : OAI21_X2 port map( B1 => n8391, B2 => n8392, A => n8390, ZN => n803);
   U348 : NAND4_X2 port map( A1 => n9336, A2 => n9337, A3 => n9334, A4 => n9335
                           , ZN => n10248);
   U372 : CLKBUF_X1 port map( A => n18635, Z => n20348);
   U374 : BUF_X2 port map( A => n18635, Z => n20349);
   U376 : XNOR2_X1 port map( A => n16357, B => n16356, ZN => n18635);
   U380 : OAI21_X2 port map( B1 => n15160, B2 => n13887, A => n13886, ZN => 
                           n16587);
   U385 : OAI21_X2 port map( B1 => n3183, B2 => n972, A => n3185, ZN => n10280)
                           ;
   U392 : AOI22_X2 port map( A1 => n3943, A2 => n3942, B1 => n3941, B2 => 
                           n19581, ZN => n5581);
   U399 : AND2_X2 port map( A1 => n7875, A2 => n7874, ZN => n8991);
   U402 : XNOR2_X2 port map( A => Key(44), B => Plaintext(44), ZN => n4482);
   U409 : BUF_X2 port map( A => n9250, Z => n9252);
   U412 : XNOR2_X2 port map( A => Plaintext(38), B => Key(38), ZN => n4892);
   U429 : XNOR2_X2 port map( A => n6965, B => n6964, ZN => n7972);
   U442 : NAND3_X2 port map( A1 => n2025, A2 => n7465, A3 => n2024, ZN => 
                           n10482);
   U455 : OAI211_X2 port map( C1 => n5660, C2 => n4776, A => n4775, B => n368, 
                           ZN => n7384);
   U477 : XNOR2_X2 port map( A => n6683, B => n6684, ZN => n8261);
   U480 : AOI21_X2 port map( B1 => n13880, B2 => n13879, A => n13878, ZN => 
                           n15195);
   U482 : CLKBUF_X1 port map( A => n12421, Z => n20350);
   U485 : BUF_X1 port map( A => n12421, Z => n20351);
   U486 : BUF_X1 port map( A => n12421, Z => n20352);
   U490 : NAND2_X2 port map( A1 => n787, A2 => n15404, ZN => n16568);
   U492 : XNOR2_X2 port map( A => n6238, B => n6239, ZN => n7936);
   U499 : AOI22_X2 port map( A1 => n1591, A2 => n12615, B1 => n874, B2 => 
                           n12242, ZN => n11983);
   U506 : NAND2_X2 port map( A1 => n8739, A2 => n3504, ZN => n9902);
   U523 : NOR2_X2 port map( A1 => n13055, A2 => n13056, ZN => n15454);
   U531 : NAND3_X2 port map( A1 => n697, A2 => n12132, A3 => n695, ZN => n13250
                           );
   U538 : AND2_X2 port map( A1 => n8715, A2 => n8714, ZN => n9646);
   U543 : XNOR2_X2 port map( A => n2990, B => Key(142), ZN => n5018);
   U548 : XNOR2_X2 port map( A => Key(133), B => Plaintext(133), ZN => n5022);
   U556 : XNOR2_X2 port map( A => n12560, B => n12561, ZN => n14790);
   U562 : NOR2_X2 port map( A1 => n10311, A2 => n10312, ZN => n12332);
   U600 : OAI21_X2 port map( B1 => n9517, B2 => n1670, A => n1669, ZN => n11670
                           );
   U601 : MUX2_X2 port map( A => n8404, B => n8403, S => n9166, Z => n10472);
   U602 : OAI21_X2 port map( B1 => n14004, B2 => n14003, A => n14002, ZN => 
                           n15695);
   U610 : OAI211_X2 port map( C1 => n31, C2 => n5470, A => n5469, B => n5468, 
                           ZN => n7263);
   U629 : XNOR2_X2 port map( A => n13450, B => n13449, ZN => n14554);
   U633 : OAI211_X2 port map( C1 => n20439, C2 => n4822, A => n5948, B => n4821
                           , ZN => n6918);
   U640 : NAND2_X2 port map( A1 => n15913, A2 => n1152, ZN => n16225);
   U645 : XNOR2_X2 port map( A => Key(92), B => Plaintext(92), ZN => n5092);
   U660 : BUF_X1 port map( A => n17244, Z => n20353);
   U662 : XNOR2_X1 port map( A => n15998, B => n15176, ZN => n17244);
   U681 : OAI21_X2 port map( B1 => n4051, B2 => n3259, A => n4050, ZN => n6042)
                           ;
   U688 : XNOR2_X2 port map( A => Key(160), B => Plaintext(160), ZN => n4574);
   U691 : OAI21_X2 port map( B1 => n10940, B2 => n10939, A => n10938, ZN => 
                           n12228);
   U693 : XNOR2_X2 port map( A => Key(36), B => Plaintext(36), ZN => n4136);
   U694 : XNOR2_X2 port map( A => n7195, B => n6300, ZN => n6824);
   U699 : NAND2_X2 port map( A1 => n5206, A2 => n1474, ZN => n7195);
   U708 : MUX2_X2 port map( A => n4813, B => n4812, S => n5080, Z => n6097);
   U711 : XNOR2_X2 port map( A => n6543, B => n6544, ZN => n8232);
   U722 : NOR2_X2 port map( A1 => n5679, A2 => n5678, ZN => n19765);
   U728 : XNOR2_X2 port map( A => n9732, B => n9731, ZN => n11397);
   U730 : XNOR2_X2 port map( A => n10169, B => n10170, ZN => n11106);
   U738 : XNOR2_X2 port map( A => Key(59), B => Plaintext(59), ZN => n3996);
   U742 : BUF_X2 port map( A => n12831, Z => n13544);
   U747 : XNOR2_X2 port map( A => n13814, B => n13813, ZN => n14601);
   U749 : NAND2_X2 port map( A1 => n8746, A2 => n19604, ZN => n10213);
   U750 : CLKBUF_X1 port map( A => n4868, Z => n20355);
   U761 : CLKBUF_X1 port map( A => n4868, Z => n20356);
   U765 : XNOR2_X1 port map( A => n3982, B => Key(65), ZN => n4868);
   U776 : NAND3_X2 port map( A1 => n1437, A2 => n14297, A3 => n14298, ZN => 
                           n16755);
   U781 : AND3_X2 port map( A1 => n709, A2 => n711, A3 => n710, ZN => n9107);
   U785 : NAND4_X2 port map( A1 => n5724, A2 => n5723, A3 => n5722, A4 => n5721
                           , ZN => n6917);
   U788 : XNOR2_X2 port map( A => n13245, B => n13246, ZN => n14570);
   U802 : OAI21_X2 port map( B1 => n10754, B2 => n10753, A => n10752, ZN => 
                           n12407);
   U804 : XNOR2_X2 port map( A => Key(47), B => Plaintext(47), ZN => n4479);
   U815 : OAI211_X2 port map( C1 => n12199, C2 => n13907, A => n12198, B => 
                           n12197, ZN => n15769);
   U816 : NOR2_X2 port map( A1 => n14322, A2 => n3149, ZN => n15553);
   U817 : NOR2_X2 port map( A1 => n18050, A2 => n18049, ZN => n3030);
   U819 : XNOR2_X2 port map( A => Key(158), B => Plaintext(158), ZN => n4576);
   U825 : AOI21_X2 port map( B1 => n12000, B2 => n11999, A => n2658, ZN => 
                           n13081);
   U832 : OR2_X2 port map( A1 => n3323, A2 => n3322, ZN => n5691);
   U835 : OAI211_X2 port map( C1 => n4523, C2 => n4191, A => n4190, B => n4189,
                           ZN => n5425);
   U836 : NAND2_X2 port map( A1 => n3334, A2 => n3336, ZN => n8998);
   U838 : XNOR2_X2 port map( A => n10378, B => n10377, ZN => n11133);
   U840 : OAI21_X2 port map( B1 => n8476, B2 => n8974, A => n577, ZN => n10281)
                           ;
   U863 : XNOR2_X2 port map( A => n1088, B => Key(64), ZN => n4652);
   U875 : XNOR2_X2 port map( A => Key(3), B => Plaintext(3), ZN => n4623);
   U881 : OAI211_X2 port map( C1 => n5935, C2 => n5934, A => n5932, B => n19, 
                           ZN => n6768);
   U883 : OAI21_X2 port map( B1 => n9012, B2 => n9013, A => n9011, ZN => n10008
                           );
   U884 : XNOR2_X2 port map( A => Key(50), B => Plaintext(50), ZN => n4907);
   U896 : NOR2_X2 port map( A1 => n11892, A2 => n11891, ZN => n12267);
   U900 : OAI21_X2 port map( B1 => n13132, B2 => n14263, A => n13133, ZN => 
                           n15683);
   U903 : XNOR2_X2 port map( A => n10155, B => n10156, ZN => n11105);
   U913 : AOI21_X2 port map( B1 => n2002, B2 => n14438, A => n14437, ZN => 
                           n15297);
   U917 : AOI22_X2 port map( A1 => n7847, A2 => n8217, B1 => n7648, B2 => n7647
                           , ZN => n8742);
   U918 : AOI22_X2 port map( A1 => n13935, A2 => n13934, B1 => n20453, B2 => 
                           n13936, ZN => n15505);
   U925 : OAI21_X2 port map( B1 => n20435, B2 => n14969, A => n14967, ZN => 
                           n17366);
   U930 : XNOR2_X2 port map( A => n17371, B => n17372, ZN => n18260);
   U931 : OAI211_X2 port map( C1 => n7712, C2 => n8363, A => n7710, B => n7711,
                           ZN => n8879);
   U938 : AND3_X2 port map( A1 => n2863, A2 => n3777, A3 => n10070, ZN => 
                           n13588);
   U943 : NOR2_X2 port map( A1 => n15118, A2 => n15117, ZN => n17111);
   U964 : OAI21_X2 port map( B1 => n14687, B2 => n859, A => n14686, ZN => 
                           n16853);
   U968 : AND2_X2 port map( A1 => n370, A2 => n11531, ZN => n9933);
   U970 : XNOR2_X2 port map( A => n8440, B => n8441, ZN => n11527);
   U979 : BUF_X1 port map( A => n7764, Z => n20359);
   U982 : XNOR2_X1 port map( A => n6243, B => n6242, ZN => n7764);
   U996 : BUF_X2 port map( A => n18377, Z => n20361);
   U997 : INV_X1 port map( A => n15454, ZN => n20362);
   U1000 : INV_X1 port map( A => n14452, ZN => n14448);
   U1004 : INV_X1 port map( A => n12533, ZN => n20363);
   U1018 : INV_X1 port map( A => n180, ZN => n1371);
   U1030 : XNOR2_X1 port map( A => n7131, B => n7132, ZN => n7953);
   U1040 : BUF_X1 port map( A => n5118, Z => n169);
   U1054 : CLKBUF_X1 port map( A => Key(54), Z => n20593);
   U1060 : CLKBUF_X1 port map( A => Key(142), Z => n20672);
   U1080 : CLKBUF_X1 port map( A => Key(179), Z => n18278);
   U1081 : BUF_X1 port map( A => Key(100), Z => n20682);
   U1083 : BUF_X1 port map( A => Key(51), Z => n2445);
   U1087 : CLKBUF_X1 port map( A => Key(33), Z => n18084);
   U1091 : CLKBUF_X1 port map( A => Key(137), Z => n2317);
   U1106 : AND2_X1 port map( A1 => n16075, A2 => n16076, ZN => n20460);
   U1124 : INV_X1 port map( A => n19284, ZN => n20364);
   U1130 : OAI21_X1 port map( B1 => n17555, B2 => n18106, A => n17554, ZN => 
                           n18622);
   U1140 : AND3_X1 port map( A1 => n17971, A2 => n17970, A3 => n17969, ZN => 
                           n18672);
   U1149 : NAND3_X1 port map( A1 => n17702, A2 => n17703, A3 => n1921, ZN => 
                           n19046);
   U1189 : AND3_X1 port map( A1 => n2662, A2 => n2664, A3 => n2660, ZN => 
                           n19682);
   U1196 : OR2_X1 port map( A1 => n16815, A2 => n16814, ZN => n19668);
   U1215 : AOI21_X1 port map( B1 => n17159, B2 => n17158, A => n17157, ZN => 
                           n19656);
   U1260 : INV_X1 port map( A => n18585, ZN => n20365);
   U1273 : BUF_X2 port map( A => n17497, Z => n19815);
   U1276 : BUF_X1 port map( A => n17695, Z => n18962);
   U1286 : BUF_X2 port map( A => n19371, Z => n19666);
   U1290 : XNOR2_X1 port map( A => n16299, B => n16298, ZN => n19403);
   U1291 : OR2_X1 port map( A1 => n3710, A2 => n15421, ZN => n15917);
   U1305 : AND2_X1 port map( A1 => n15676, A2 => n15443, ZN => n20647);
   U1323 : NAND3_X1 port map( A1 => n700, A2 => n12927, A3 => n12928, ZN => 
                           n15379);
   U1326 : AND2_X1 port map( A1 => n2920, A2 => n20624, ZN => n15459);
   U1329 : NAND2_X1 port map( A1 => n13910, A2 => n2654, ZN => n2655);
   U1372 : NOR2_X1 port map( A1 => n13998, A2 => n13999, ZN => n20449);
   U1373 : OR2_X1 port map( A1 => n14666, A2 => n14667, ZN => n14315);
   U1394 : XNOR2_X1 port map( A => n2095, B => n13854, ZN => n20513);
   U1404 : XNOR2_X1 port map( A => n11318, B => n11317, ZN => n14778);
   U1419 : XNOR2_X1 port map( A => n13107, B => n13106, ZN => n13981);
   U1425 : OAI21_X1 port map( B1 => n12684, B2 => n11613, A => n11612, ZN => 
                           n13707);
   U1428 : OR2_X1 port map( A1 => n11692, A2 => n11646, ZN => n1951);
   U1430 : OR2_X1 port map( A1 => n11464, A2 => n12524, ZN => n11793);
   U1434 : CLKBUF_X1 port map( A => n12639, Z => n922);
   U1456 : AND2_X1 port map( A1 => n10933, A2 => n3105, ZN => n20583);
   U1489 : MUX2_X1 port map( A => n10832, B => n10831, S => n11420, Z => n20430
                           );
   U1512 : NAND3_X1 port map( A1 => n10707, A2 => n20522, A3 => n20521, ZN => 
                           n12630);
   U1530 : OR2_X1 port map( A1 => n10705, A2 => n10951, ZN => n20522);
   U1541 : OR2_X1 port map( A1 => n10708, A2 => n11011, ZN => n20521);
   U1542 : BUF_X2 port map( A => n11144, Z => n20366);
   U1548 : XNOR2_X1 port map( A => n9460, B => n9461, ZN => n10953);
   U1555 : AND2_X1 port map( A1 => n20646, A2 => n506, ZN => n8746);
   U1573 : INV_X1 port map( A => n9794, ZN => n20608);
   U1578 : OR2_X1 port map( A1 => n363, A2 => n362, ZN => n10237);
   U1584 : OR2_X1 port map( A1 => n8484, A2 => n8602, ZN => n20659);
   U1591 : OR2_X1 port map( A1 => n1507, A2 => n9453, ZN => n401);
   U1600 : AND3_X2 port map( A1 => n1679, A2 => n1678, A3 => n1677, ZN => n1507
                           );
   U1668 : NAND4_X1 port map( A1 => n3581, A2 => n7483, A3 => n7484, A4 => 
                           n7482, ZN => n8812);
   U1669 : INV_X1 port map( A => n8208, ZN => n20585);
   U1687 : XNOR2_X1 port map( A => n6335, B => n6336, ZN => n8354);
   U1690 : CLKBUF_X1 port map( A => n6887, Z => n20455);
   U1701 : XNOR2_X1 port map( A => n6317, B => n6316, ZN => n7981);
   U1705 : INV_X1 port map( A => n7479, ZN => n20367);
   U1731 : NAND3_X1 port map( A1 => n2555, A2 => n5459, A3 => n2556, ZN => 
                           n7070);
   U1749 : NAND3_X1 port map( A1 => n20411, A2 => n20410, A3 => n4097, ZN => 
                           n5989);
   U1752 : NAND2_X1 port map( A1 => n4375, A2 => n4369, ZN => n5720);
   U1791 : INV_X1 port map( A => n5914, ZN => n20368);
   U1793 : OR2_X1 port map( A1 => n4424, A2 => n4423, ZN => n20655);
   U1797 : OR2_X1 port map( A1 => n4098, A2 => n5024, ZN => n20411);
   U1816 : OR2_X1 port map( A1 => n4711, A2 => n4769, ZN => n20679);
   U1818 : OR2_X1 port map( A1 => n4481, A2 => n3967, ZN => n20606);
   U1837 : XNOR2_X1 port map( A => n20635, B => Key(56), ZN => n3995);
   U1845 : XNOR2_X1 port map( A => n3970, B => Key(37), ZN => n4960);
   U1850 : XNOR2_X1 port map( A => n3869, B => Key(31), ZN => n4474);
   U1866 : OR2_X1 port map( A1 => n2490, A2 => n4987, ZN => n2489);
   U1876 : BUF_X1 port map( A => n4060, Z => n4588);
   U1904 : AND2_X1 port map( A1 => n3527, A2 => n5685, ZN => n20553);
   U1913 : INV_X1 port map( A => n6156, ZN => n20403);
   U1952 : AND2_X1 port map( A1 => n5971, A2 => n5699, ZN => n20674);
   U1960 : OAI211_X1 port map( C1 => n5056, C2 => n4739, A => n4590, B => n4588
                           , ZN => n5885);
   U1965 : INV_X1 port map( A => n2454, ZN => n20551);
   U1997 : OR2_X1 port map( A1 => n3948, A2 => n4350, ZN => n4256);
   U1999 : BUF_X1 port map( A => n6404, Z => n19855);
   U2027 : AND2_X1 port map( A1 => n7633, A2 => n20511, ZN => n20586);
   U2028 : AND2_X1 port map( A1 => n19922, A2 => n8205, ZN => n20584);
   U2037 : OR2_X1 port map( A1 => n20177, A2 => n8387, ZN => n7685);
   U2056 : BUF_X1 port map( A => n8380, Z => n163);
   U2058 : INV_X1 port map( A => n7953, ZN => n20013);
   U2059 : OR2_X1 port map( A1 => n8744, A2 => n8602, ZN => n20646);
   U2110 : INV_X1 port map( A => n7590, ZN => n20651);
   U2117 : BUF_X1 port map( A => n8004, Z => n8312);
   U2119 : AND2_X1 port map( A1 => n19565, A2 => n20554, ZN => n2888);
   U2123 : CLKBUF_X1 port map( A => n8993, Z => n19732);
   U2133 : INV_X1 port map( A => n20010, ZN => n9090);
   U2136 : OR2_X1 port map( A1 => n9250, A2 => n9249, ZN => n9260);
   U2139 : OR2_X1 port map( A1 => n9313, A2 => n9228, ZN => n9227);
   U2140 : NOR2_X1 port map( A1 => n20659, A2 => n8485, ZN => n8486);
   U2158 : NAND2_X1 port map( A1 => n10329, A2 => n10328, ZN => n10052);
   U2162 : INV_X1 port map( A => n8593, ZN => n10620);
   U2170 : AND2_X1 port map( A1 => n8734, A2 => n8499, ZN => n8334);
   U2190 : OAI211_X1 port map( C1 => n8278, C2 => n8279, A => n8433, B => n8277
                           , ZN => n10431);
   U2191 : AOI21_X1 port map( B1 => n11281, B2 => n11284, A => n19817, ZN => 
                           n20641);
   U2192 : OAI21_X1 port map( B1 => n10719, B2 => n1988, A => n11192, ZN => 
                           n20561);
   U2223 : XNOR2_X1 port map( A => n8481, B => n8480, ZN => n11521);
   U2226 : OR2_X1 port map( A1 => n19983, A2 => n11186, ZN => n20591);
   U2240 : AND2_X1 port map( A1 => n19864, A2 => n11513, ZN => n20560);
   U2245 : BUF_X1 port map( A => n10259, Z => n11886);
   U2261 : INV_X1 port map( A => n20496, ZN => n20660);
   U2266 : INV_X1 port map( A => n3401, ZN => n11722);
   U2286 : NOR2_X1 port map( A1 => n10750, A2 => n10749, ZN => n12408);
   U2322 : NOR2_X1 port map( A1 => n12149, A2 => n20618, ZN => n19558);
   U2354 : BUF_X1 port map( A => n12021, Z => n20191);
   U2361 : AND2_X1 port map( A1 => n11695, A2 => n953, ZN => n20644);
   U2364 : AND3_X2 port map( A1 => n10714, A2 => n10715, A3 => n10713, ZN => 
                           n11618);
   U2380 : XNOR2_X1 port map( A => n13398, B => n13422, ZN => n13649);
   U2384 : OR2_X1 port map( A1 => n14482, A2 => n14171, ZN => n14485);
   U2392 : XNOR2_X1 port map( A => n12968, B => n12967, ZN => n14512);
   U2411 : AND2_X1 port map( A1 => n13556, A2 => n2921, ZN => n20624);
   U2418 : INV_X1 port map( A => n13931, ZN => n14339);
   U2433 : BUF_X1 port map( A => n14820, Z => n912);
   U2434 : CLKBUF_X1 port map( A => n14087, Z => n19821);
   U2437 : NOR2_X1 port map( A1 => n13317, A2 => n14705, ZN => n13318);
   U2482 : NAND2_X1 port map( A1 => n20609, A2 => n19613, ZN => n15583);
   U2485 : OAI211_X1 port map( C1 => n20513, C2 => n2682, A => n2666, B => 
                           n13855, ZN => n15443);
   U2489 : OR2_X1 port map( A1 => n15677, A2 => n15228, ZN => n15445);
   U2495 : OR2_X1 port map( A1 => n14667, A2 => n14663, ZN => n13166);
   U2502 : MUX2_X1 port map( A => n14618, B => n14617, S => n20112, Z => n14631
                           );
   U2510 : NOR2_X1 port map( A1 => n14670, A2 => n14671, ZN => n860);
   U2517 : INV_X1 port map( A => n20101, ZN => n20391);
   U2521 : XNOR2_X1 port map( A => n14956, B => n16711, ZN => n17026);
   U2541 : OR2_X1 port map( A1 => n17530, A2 => n19110, ZN => n20661);
   U2546 : CLKBUF_X1 port map( A => n17836, Z => n20423);
   U2556 : XNOR2_X1 port map( A => n16040, B => n16041, ZN => n19707);
   U2557 : CLKBUF_X1 port map( A => n16166, Z => n16480);
   U2563 : AND2_X1 port map( A1 => n811, A2 => n814, ZN => n20654);
   U2571 : NOR2_X1 port map( A1 => n18036, A2 => n18035, ZN => n18857);
   U2617 : CLKBUF_X1 port map( A => Key(119), Z => n17999);
   U2624 : INV_X1 port map( A => n2067, ZN => n16788);
   U2632 : XOR2_X1 port map( A => Key(176), B => Plaintext(176), Z => n20369);
   U2634 : NAND3_X1 port map( A1 => n2120, A2 => n18932, A3 => n18029, ZN => 
                           n20370);
   U2652 : OR2_X1 port map( A1 => n14214, A2 => n15071, ZN => n20371);
   U2656 : XOR2_X1 port map( A => n17035, B => n17270, Z => n20372);
   U2657 : INV_X1 port map( A => n5741, ZN => n20568);
   U2679 : AND2_X1 port map( A1 => n19856, A2 => n8001, ZN => n20373);
   U2690 : INV_X1 port map( A => n6155, ZN => n20405);
   U2708 : AND2_X1 port map( A1 => n8095, A2 => n7632, ZN => n20374);
   U2727 : OR2_X1 port map( A1 => n10654, A2 => n19872, ZN => n20375);
   U2734 : XOR2_X1 port map( A => n13373, B => n13372, Z => n20376);
   U2777 : XOR2_X1 port map( A => n2095, B => n13854, Z => n20377);
   U2779 : XOR2_X1 port map( A => n13622, B => n18988, Z => n20378);
   U2789 : OR2_X1 port map( A1 => n15535, A2 => n15895, ZN => n20379);
   U2791 : XOR2_X1 port map( A => n12983, B => n12982, Z => n20380);
   U2821 : INV_X1 port map( A => n14778, ZN => n20408);
   U2835 : AND2_X1 port map( A1 => n19940, A2 => n14499, ZN => n20381);
   U2837 : AND2_X1 port map( A1 => n19439, A2 => n19440, ZN => n20382);
   U2838 : AND2_X1 port map( A1 => n19170, A2 => n20394, ZN => n20383);
   U2879 : AND2_X1 port map( A1 => n20396, A2 => n20393, ZN => n20384);
   U2880 : OAI21_X2 port map( B1 => n2671, B2 => n2670, A => n20385, ZN => 
                           n6101);
   U2889 : NAND2_X1 port map( A1 => n4800, A2 => n5043, ZN => n20385);
   U2891 : XNOR2_X1 port map( A => n20386, B => n311, ZN => Ciphertext(14));
   U2905 : NAND2_X1 port map( A1 => n20549, A2 => n15930, ZN => n20386);
   U2915 : NAND3_X2 port map( A1 => n20387, A2 => n7055, A3 => n92, ZN => n9038
                           );
   U2923 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => n20387);
   U2941 : NAND2_X1 port map( A1 => n6041, A2 => n1214, ZN => n6043);
   U2973 : NAND2_X2 port map( A1 => n1320, A2 => n4043, ZN => n6041);
   U2974 : OR2_X2 port map( A1 => n7630, A2 => n7629, ZN => n8482);
   U2980 : NAND2_X1 port map( A1 => n7626, A2 => n1335, ZN => n7630);
   U2981 : NAND3_X1 port map( A1 => n241, A2 => n20390, A3 => n20388, ZN => 
                           n1700);
   U2995 : NAND2_X1 port map( A1 => n20389, A2 => n14547, ZN => n20388);
   U3002 : INV_X1 port map( A => n20471, ZN => n20389);
   U3012 : OR2_X1 port map( A1 => n14548, A2 => n14547, ZN => n20390);
   U3051 : AND3_X2 port map( A1 => n14068, A2 => n14067, A3 => n2528, ZN => 
                           n864);
   U3052 : NAND2_X1 port map( A1 => n3479, A2 => n3478, ZN => n12531);
   U3063 : NAND2_X1 port map( A1 => n20392, A2 => n20391, ZN => n17950);
   U3066 : NAND2_X1 port map( A1 => n18131, A2 => n19744, ZN => n20392);
   U3067 : OAI21_X1 port map( B1 => n9365, B2 => n9366, A => n9364, ZN => n598)
                           ;
   U3091 : NAND2_X1 port map( A1 => n8958, A2 => n8960, ZN => n9366);
   U3094 : NAND3_X1 port map( A1 => n20412, A2 => n3346, A3 => n3217, ZN => 
                           n18009);
   U3173 : NAND3_X1 port map( A1 => n17951, A2 => n17953, A3 => n17952, ZN => 
                           n18667);
   U3175 : AND3_X2 port map( A1 => n2106, A2 => n11135, A3 => n11134, ZN => 
                           n12386);
   U3177 : NAND2_X1 port map( A1 => n20395, A2 => n20394, ZN => n20393);
   U3178 : INV_X1 port map( A => n2368, ZN => n20394);
   U3194 : INV_X1 port map( A => n18156, ZN => n20395);
   U3240 : NAND2_X1 port map( A1 => n16159, A2 => n20383, ZN => n20396);
   U3283 : XNOR2_X1 port map( A => n20397, B => n18066, ZN => Ciphertext(115));
   U3301 : NAND2_X1 port map( A1 => n2399, A2 => n18063, ZN => n20397);
   U3334 : NAND2_X1 port map( A1 => n19993, A2 => n18061, ZN => n19035);
   U3358 : INV_X1 port map( A => n792, ZN => n5613);
   U3395 : NAND2_X1 port map( A1 => n6153, A2 => n5611, ZN => n792);
   U3420 : NAND2_X1 port map( A1 => n10989, A2 => n10988, ZN => n11683);
   U3443 : NAND2_X1 port map( A1 => n5956, A2 => n20398, ZN => n941);
   U3507 : NOR2_X1 port map( A1 => n367, A2 => n145, ZN => n20398);
   U3514 : XNOR2_X1 port map( A => n20399, B => n15579, ZN => n15586);
   U3587 : XNOR2_X1 port map( A => n15571, B => n17407, ZN => n20399);
   U3588 : NAND2_X1 port map( A1 => n20401, A2 => n20400, ZN => n3401);
   U3589 : NAND2_X1 port map( A1 => n10702, A2 => n20366, ZN => n20400);
   U3594 : NAND2_X1 port map( A1 => n10703, A2 => n11140, ZN => n20401);
   U3597 : NAND2_X1 port map( A1 => n5247, A2 => n20402, ZN => n7254);
   U3604 : NAND3_X1 port map( A1 => n20406, A2 => n20404, A3 => n20403, ZN => 
                           n20402);
   U3672 : NAND2_X1 port map( A1 => n20405, A2 => n6150, ZN => n20404);
   U3690 : NAND2_X1 port map( A1 => n6151, A2 => n6155, ZN => n20406);
   U3691 : NAND2_X1 port map( A1 => n20409, A2 => n20407, ZN => n14856);
   U3708 : NAND2_X1 port map( A1 => n11320, A2 => n20408, ZN => n20407);
   U3711 : NAND2_X1 port map( A1 => n11319, A2 => n14778, ZN => n20409);
   U3723 : NAND3_X1 port map( A1 => n20043, A2 => n4098, A3 => n5029, ZN => 
                           n20410);
   U3764 : NAND2_X1 port map( A1 => n20013, A2 => n7952, ZN => n7813);
   U3783 : BUF_X1 port map( A => n14781, Z => n20518);
   U3805 : NAND2_X1 port map( A1 => n17490, A2 => n3347, ZN => n20412);
   U3837 : NAND2_X1 port map( A1 => n12095, A2 => n12430, ZN => n3514);
   U3846 : NAND3_X1 port map( A1 => n8727, A2 => n1023, A3 => n20413, ZN => 
                           n1268);
   U3956 : NAND2_X1 port map( A1 => n8726, A2 => n9361, ZN => n20413);
   U3957 : NOR2_X2 port map( A1 => n14047, A2 => n20414, ZN => n15845);
   U3993 : NAND2_X1 port map( A1 => n340, A2 => n341, ZN => n20414);
   U4028 : NAND2_X1 port map( A1 => n14405, A2 => n14148, ZN => n14010);
   U4029 : AOI22_X2 port map( A1 => n14183, A2 => n14182, B1 => n14450, B2 => 
                           n14181, ZN => n15310);
   U4057 : NAND3_X1 port map( A1 => n1213, A2 => n12335, A3 => n11992, ZN => 
                           n11993);
   U4066 : OAI211_X2 port map( C1 => n8754, C2 => n8933, A => n20416, B => 
                           n20415, ZN => n9952);
   U4072 : NAND2_X1 port map( A1 => n8750, A2 => n8933, ZN => n20415);
   U4076 : NAND2_X1 port map( A1 => n8751, A2 => n8752, ZN => n20416);
   U4117 : OR2_X1 port map( A1 => n8065, A2 => n1431, ZN => n20505);
   U4120 : AND3_X1 port map( A1 => n13958, A2 => n13956, A3 => n402, ZN => 
                           n19739);
   U4141 : XNOR2_X1 port map( A => n15347, B => n15346, ZN => n17501);
   U4144 : INV_X1 port map( A => n19668, ZN => n20417);
   U4162 : AND2_X1 port map( A1 => n14516, A2 => n20206, ZN => n20636);
   U4180 : NAND3_X1 port map( A1 => n20370, A2 => n20613, A3 => n20612, ZN => 
                           n20418);
   U4214 : AOI21_X2 port map( B1 => n15605, B2 => n15274, A => n15011, ZN => 
                           n15935);
   U4262 : NAND3_X1 port map( A1 => n20370, A2 => n20613, A3 => n20612, ZN => 
                           n18868);
   U4270 : NOR2_X2 port map( A1 => n20419, A2 => n20420, ZN => n16844);
   U4272 : AND2_X1 port map( A1 => n15203, A2 => n16126, ZN => n20419);
   U4340 : NAND2_X1 port map( A1 => n57, A2 => n55, ZN => n20420);
   U4356 : XOR2_X1 port map( A => n16884, B => n16883, Z => n20421);
   U4360 : NAND2_X1 port map( A1 => n17313, A2 => n17312, ZN => n20422);
   U4408 : OR2_X1 port map( A1 => n9274, A2 => n885, ZN => n20554);
   U4469 : XNOR2_X1 port map( A => n16143, B => n16144, ZN => n17836);
   U4477 : OR2_X1 port map( A1 => n20286, A2 => n19094, ZN => n2196);
   U4498 : OR2_X1 port map( A1 => n20142, A2 => n19031, ZN => n20528);
   U4587 : XNOR2_X1 port map( A => n13117, B => n13116, ZN => n20424);
   U4635 : XNOR2_X1 port map( A => n5297, B => n6835, ZN => n8303);
   U4636 : XNOR2_X1 port map( A => n16392, B => n20426, ZN => n20425);
   U4638 : XOR2_X1 port map( A => n16840, B => n16651, Z => n20426);
   U4643 : XNOR2_X1 port map( A => n11756, B => n11755, ZN => n14807);
   U4644 : XNOR2_X1 port map( A => n20425, B => n16395, ZN => n19658);
   U4646 : XNOR2_X1 port map( A => n16150, B => n16149, ZN => n17715);
   U4658 : NOR2_X2 port map( A1 => n16728, A2 => n16729, ZN => n16780);
   U4672 : OAI21_X1 port map( B1 => n15429, B2 => n15428, A => n15427, ZN => 
                           n15534);
   U4677 : AND2_X1 port map( A1 => n9444, A2 => n9443, ZN => n20427);
   U4709 : AND2_X1 port map( A1 => n9444, A2 => n9443, ZN => n11650);
   U4710 : OR2_X1 port map( A1 => n20182, A2 => n15371, ZN => n20428);
   U4717 : BUF_X1 port map( A => n17572, Z => n20429);
   U4736 : MUX2_X1 port map( A => n10832, B => n10831, S => n11420, Z => n12594
                           );
   U4749 : INV_X1 port map( A => n5081, ZN => n20431);
   U4760 : AND2_X1 port map( A1 => n12129, A2 => n12126, ZN => n696);
   U4765 : BUF_X1 port map( A => n14714, Z => n19862);
   U4770 : MUX2_X1 port map( A => n14860, B => n14861, S => n15237, Z => n14862
                           );
   U4782 : INV_X1 port map( A => n15237, ZN => n1458);
   U4792 : INV_X1 port map( A => n18382, ZN => n20611);
   U4809 : NOR2_X1 port map( A1 => n19599, A2 => n15180, ZN => n15186);
   U4810 : AND2_X1 port map( A1 => n15656, A2 => n15659, ZN => n20565);
   U4816 : OR2_X1 port map( A1 => n11981, A2 => n20430, ZN => n20543);
   U4830 : NOR2_X1 port map( A1 => n12644, A2 => n12643, ZN => n13154);
   U4831 : XNOR2_X1 port map( A => n16204, B => n16203, ZN => n20432);
   U4834 : INV_X1 port map( A => n214, ZN => n20433);
   U4860 : OAI21_X1 port map( B1 => n17474, B2 => n18539, A => n17473, ZN => 
                           n18511);
   U4879 : AOI22_X1 port map( A1 => n17614, A2 => n17613, B1 => n17612, B2 => 
                           n17611, ZN => n20434);
   U4883 : NAND2_X1 port map( A1 => n19573, A2 => n14960, ZN => n16927);
   U4898 : NOR2_X1 port map( A1 => n15672, A2 => n20151, ZN => n15438);
   U4946 : NOR2_X1 port map( A1 => n17551, A2 => n17550, ZN => n18630);
   U4948 : AOI22_X1 port map( A1 => n15562, A2 => n15558, B1 => n15510, B2 => 
                           n15509, ZN => n20435);
   U4949 : MUX2_X1 port map( A => n9252, B => n8971, S => n670, Z => n7736);
   U4991 : XNOR2_X1 port map( A => n16548, B => n16547, ZN => n20436);
   U5027 : INV_X1 port map( A => n18376, ZN => n20437);
   U5029 : CLKBUF_X1 port map( A => Key(36), Z => n620);
   U5035 : CLKBUF_X1 port map( A => n18257, Z => n20438);
   U5038 : INV_X1 port map( A => n19658, ZN => n17956);
   U5082 : OR2_X1 port map( A1 => n5663, A2 => n5952, ZN => n20439);
   U5095 : OR2_X1 port map( A1 => n5663, A2 => n5952, ZN => n5661);
   U5099 : OAI21_X1 port map( B1 => n12358, B2 => n12357, A => n12356, ZN => 
                           n20440);
   U5100 : OAI21_X1 port map( B1 => n12358, B2 => n12357, A => n12356, ZN => 
                           n13826);
   U5110 : INV_X1 port map( A => n15228, ZN => n15679);
   U5121 : OR2_X1 port map( A1 => n17208, A2 => n17210, ZN => n20633);
   U5135 : NAND3_X1 port map( A1 => n14933, A2 => n14932, A3 => n460, ZN => 
                           n16602);
   U5147 : AND2_X1 port map( A1 => n17565, A2 => n17471, ZN => n18538);
   U5153 : OR2_X1 port map( A1 => n14836, A2 => n15813, ZN => n579);
   U5184 : AOI22_X1 port map( A1 => n5038, A2 => n5039, B1 => n5036, B2 => 
                           n5037, ZN => n6025);
   U5210 : XNOR2_X1 port map( A => n6452, B => n6451, ZN => n20441);
   U5215 : XNOR2_X1 port map( A => n12906, B => n13848, ZN => n20442);
   U5222 : XNOR2_X1 port map( A => n12983, B => n12982, ZN => n20443);
   U5228 : OAI211_X1 port map( C1 => n18658, C2 => n18659, A => n20581, B => 
                           n20580, ZN => n18661);
   U5231 : CLKBUF_X1 port map( A => n19276, Z => n20444);
   U5258 : INV_X1 port map( A => n8831, ZN => n8829);
   U5285 : NAND2_X2 port map( A1 => n1725, A2 => n7535, ZN => n8736);
   U5292 : NAND3_X1 port map( A1 => n17148, A2 => n3065, A3 => n3064, ZN => 
                           n20445);
   U5293 : NAND3_X1 port map( A1 => n17148, A2 => n3065, A3 => n3064, ZN => 
                           n18585);
   U5295 : OAI21_X1 port map( B1 => n14343, B2 => n14106, A => n14105, ZN => 
                           n15746);
   U5302 : OR2_X1 port map( A1 => n4898, A2 => n20446, ZN => n2573);
   U5318 : NOR2_X1 port map( A1 => n4899, A2 => n4962, ZN => n20446);
   U5329 : OR2_X1 port map( A1 => n16795, A2 => n20648, ZN => n1337);
   U5356 : CLKBUF_X1 port map( A => n1205, Z => n20447);
   U5364 : BUF_X1 port map( A => n19274, Z => n20448);
   U5365 : MUX2_X1 port map( A => n19675, B => n3347, S => n17154, Z => n16247)
                           ;
   U5401 : NOR2_X1 port map( A1 => n11062, A2 => n11726, ZN => n20623);
   U5429 : OR3_X1 port map( A1 => n15857, A2 => n15329, A3 => n15327, ZN => 
                           n15331);
   U5438 : OR2_X1 port map( A1 => n15863, A2 => n15857, ZN => n15332);
   U5439 : OAI21_X1 port map( B1 => n2581, B2 => n15870, A => n15305, ZN => 
                           n20450);
   U5526 : OAI21_X1 port map( B1 => n2581, B2 => n15870, A => n15305, ZN => 
                           n16555);
   U5537 : XNOR2_X1 port map( A => n13373, B => n13372, ZN => n20451);
   U5538 : NOR2_X1 port map( A1 => n15906, A2 => n2723, ZN => n15417);
   U5551 : XNOR2_X1 port map( A => n17050, B => n17049, ZN => n20452);
   U5582 : XNOR2_X1 port map( A => n17050, B => n17049, ZN => n18937);
   U5585 : NAND2_X1 port map( A1 => n7850, A2 => n7849, ZN => n9265);
   U5646 : XNOR2_X1 port map( A => n13467, B => n20285, ZN => n20453);
   U5656 : XNOR2_X1 port map( A => n13467, B => n20285, ZN => n14426);
   U5662 : XNOR2_X1 port map( A => n11103, B => n11102, ZN => n20454);
   U5699 : XOR2_X1 port map( A => n9977, B => n9937, Z => n20456);
   U5748 : OR2_X1 port map( A1 => n12876, A2 => n19485, ZN => n14341);
   U5759 : OR2_X1 port map( A1 => n14335, A2 => n19485, ZN => n20665);
   U5789 : AND2_X1 port map( A1 => n20340, A2 => n382, ZN => n20457);
   U5818 : AND2_X1 port map( A1 => n20340, A2 => n382, ZN => n20458);
   U5844 : AND2_X1 port map( A1 => n20340, A2 => n382, ZN => n12455);
   U5850 : CLKBUF_X1 port map( A => n4864, Z => n20459);
   U5863 : XNOR2_X1 port map( A => n3984, B => Key(62), ZN => n4864);
   U5868 : AND2_X1 port map( A1 => n16075, A2 => n16076, ZN => n18327);
   U5873 : XNOR2_X1 port map( A => n4059, B => Key(127), ZN => n20461);
   U5892 : INV_X1 port map( A => n11686, ZN => n20462);
   U5900 : XNOR2_X1 port map( A => n4059, B => Key(127), ZN => n5052);
   U5901 : AOI22_X2 port map( A1 => n15550, A2 => n15410, B1 => n15409, B2 => 
                           n15551, ZN => n2973);
   U5929 : OR2_X1 port map( A1 => n19174, A2 => n19170, ZN => n18161);
   U5942 : OAI211_X1 port map( C1 => n19880, C2 => n19710, A => n8655, B => 
                           n8654, ZN => n10589);
   U5961 : AOI22_X1 port map( A1 => n9269, A2 => n19880, B1 => n9267, B2 => 
                           n9268, ZN => n9270);
   U5965 : XNOR2_X1 port map( A => n15613, B => n15612, ZN => n20463);
   U5976 : XNOR2_X1 port map( A => n15613, B => n15612, ZN => n19383);
   U5977 : OAI211_X1 port map( C1 => n7779, C2 => n8312, A => n7778, B => n7777
                           , ZN => n9176);
   U5993 : NAND2_X2 port map( A1 => n17598, A2 => n17597, ZN => n19292);
   U5997 : XNOR2_X1 port map( A => Key(119), B => Plaintext(119), ZN => n20464)
                           ;
   U6001 : XNOR2_X1 port map( A => n4465, B => n4466, ZN => n20465);
   U6027 : XNOR2_X1 port map( A => n4465, B => n4466, ZN => n8062);
   U6033 : CLKBUF_X1 port map( A => n14127, Z => n20466);
   U6047 : AND3_X1 port map( A1 => n19151, A2 => n19144, A3 => n19134, ZN => 
                           n3141);
   U6057 : INV_X1 port map( A => n15380, ZN => n20467);
   U6075 : BUF_X1 port map( A => n10683, Z => n20468);
   U6076 : BUF_X1 port map( A => n13396, Z => n20469);
   U6091 : OAI22_X1 port map( A1 => n12492, A2 => n12491, B1 => n12489, B2 => 
                           n12490, ZN => n13396);
   U6117 : XOR2_X1 port map( A => n9474, B => n9473, Z => n20470);
   U6146 : XNOR2_X1 port map( A => n13214, B => n13213, ZN => n20471);
   U6162 : INV_X1 port map( A => n888, ZN => n20539);
   U6167 : INV_X1 port map( A => n8846, ZN => n20472);
   U6169 : XNOR2_X1 port map( A => n12943, B => n12942, ZN => n20473);
   U6197 : BUF_X1 port map( A => n15130, Z => n20474);
   U6202 : OAI21_X1 port map( B1 => n14513, B2 => n14512, A => n14511, ZN => 
                           n15130);
   U6241 : AND3_X1 port map( A1 => n17722, A2 => n17721, A3 => n17720, ZN => 
                           n20475);
   U6264 : OAI211_X1 port map( C1 => n11545, C2 => n10889, A => n258, B => 
                           n20681, ZN => n509);
   U6291 : OR2_X1 port map( A1 => n6904, A2 => n7903, ZN => n19582);
   U6299 : OAI21_X1 port map( B1 => n12572, B2 => n12573, A => n12571, ZN => 
                           n13479);
   U6309 : OR2_X1 port map( A1 => n15588, A2 => n15760, ZN => n20667);
   U6321 : BUF_X1 port map( A => n16992, Z => n17102);
   U6354 : BUF_X1 port map( A => n9834, Z => n20476);
   U6365 : OAI211_X1 port map( C1 => n8073, C2 => n8202, A => n20020, B => 
                           n8072, ZN => n9834);
   U6370 : NOR2_X1 port map( A1 => n15215, A2 => n15214, ZN => n20477);
   U6371 : NOR2_X1 port map( A1 => n15215, A2 => n15214, ZN => n20478);
   U6384 : NOR2_X1 port map( A1 => n15215, A2 => n15214, ZN => n17123);
   U6403 : NAND2_X1 port map( A1 => n14072, A2 => n20525, ZN => n16593);
   U6421 : XNOR2_X1 port map( A => n9097, B => n9096, ZN => n20479);
   U6425 : XNOR2_X1 port map( A => n9097, B => n9096, ZN => n10968);
   U6450 : AND2_X1 port map( A1 => n20671, A2 => n1376, ZN => n12465);
   U6478 : INV_X1 port map( A => n14228, ZN => n20480);
   U6503 : NAND2_X1 port map( A1 => n20032, A2 => n15448, ZN => n20481);
   U6510 : NAND2_X1 port map( A1 => n20032, A2 => n15448, ZN => n16965);
   U6521 : OAI211_X1 port map( C1 => n2911, C2 => n3305, A => n3754, B => n2910
                           , ZN => n20482);
   U6541 : OAI211_X1 port map( C1 => n2911, C2 => n3305, A => n3754, B => n2910
                           , ZN => n13534);
   U6566 : MUX2_X1 port map( A => n7495, B => n7494, S => n8165, Z => n9047);
   U6568 : AND2_X2 port map( A1 => n3354, A2 => n3355, ZN => n10030);
   U6576 : NOR2_X1 port map( A1 => n8856, A2 => n8855, ZN => n20483);
   U6590 : NOR2_X1 port map( A1 => n8856, A2 => n8855, ZN => n20484);
   U6603 : MUX2_X1 port map( A => n8854, B => n8853, S => n9038, Z => n8855);
   U6622 : BUF_X1 port map( A => n8041, Z => n20485);
   U6623 : AOI22_X1 port map( A1 => n11334, A2 => n11333, B1 => n11332, B2 => 
                           n11331, ZN => n20486);
   U6629 : AOI22_X1 port map( A1 => n11334, A2 => n11333, B1 => n11332, B2 => 
                           n11331, ZN => n12152);
   U6701 : XNOR2_X1 port map( A => Key(176), B => Plaintext(176), ZN => n20487)
                           ;
   U6704 : XNOR2_X1 port map( A => n16332, B => n16333, ZN => n20488);
   U6740 : XNOR2_X1 port map( A => n16332, B => n16333, ZN => n17558);
   U6762 : NOR2_X1 port map( A1 => n19418, A2 => n19439, ZN => n20571);
   U6823 : CLKBUF_X1 port map( A => n10808, Z => n10788);
   U6841 : NAND3_X2 port map( A1 => n11700, A2 => n3783, A3 => n3780, ZN => 
                           n13222);
   U6879 : OR2_X1 port map( A1 => n12644, A2 => n12643, ZN => n20489);
   U6925 : AND2_X2 port map( A1 => n16473, A2 => n16472, ZN => n20139);
   U6936 : XNOR2_X1 port map( A => n7245, B => n7244, ZN => n20490);
   U6944 : XNOR2_X1 port map( A => n7245, B => n7244, ZN => n7797);
   U6945 : XNOR2_X1 port map( A => n9824, B => n10126, ZN => n19829);
   U7011 : NAND3_X2 port map( A1 => n14865, A2 => n1443, A3 => n1444, ZN => 
                           n17339);
   U7031 : BUF_X1 port map( A => n10210, Z => n20491);
   U7038 : INV_X1 port map( A => n12313, ZN => n20618);
   U7070 : INV_X1 port map( A => n3305, ZN => n20524);
   U7156 : OAI211_X1 port map( C1 => n20230, C2 => n18541, A => n17486, B => 
                           n17485, ZN => n20492);
   U7161 : OAI211_X1 port map( C1 => n20230, C2 => n18541, A => n17486, B => 
                           n17485, ZN => n18519);
   U7222 : INV_X1 port map( A => n8100, ZN => n20493);
   U7226 : XNOR2_X1 port map( A => n17035, B => n17270, ZN => n20494);
   U7227 : NAND3_X2 port map( A1 => n14870, A2 => n14869, A3 => n14868, ZN => 
                           n17270);
   U7252 : OR2_X1 port map( A1 => n15030, A2 => n15029, ZN => n15033);
   U7274 : XOR2_X1 port map( A => n6533, B => n6532, Z => n20495);
   U7276 : XOR2_X1 port map( A => n9631, B => n9630, Z => n20496);
   U7309 : BUF_X1 port map( A => n12372, Z => n20497);
   U7313 : XNOR2_X1 port map( A => n20664, B => n13300, ZN => n20498);
   U7356 : XNOR2_X1 port map( A => n16897, B => n16896, ZN => n20499);
   U7360 : XNOR2_X1 port map( A => n16897, B => n16896, ZN => n18978);
   U7361 : XNOR2_X1 port map( A => n2833, B => n2832, ZN => n20500);
   U7366 : XNOR2_X1 port map( A => n2833, B => n2832, ZN => n14801);
   U7387 : XNOR2_X1 port map( A => n17018, B => n17017, ZN => n20501);
   U7404 : INV_X1 port map( A => n15469, ZN => n20502);
   U7407 : INV_X1 port map( A => n20502, ZN => n20503);
   U7408 : XOR2_X1 port map( A => n4728, B => n4729, Z => n20504);
   U7410 : XNOR2_X1 port map( A => n15974, B => n15973, ZN => n20506);
   U7414 : XNOR2_X1 port map( A => n15974, B => n15973, ZN => n20507);
   U7430 : OR2_X1 port map( A1 => n16728, A2 => n16729, ZN => n20508);
   U7491 : MUX2_X1 port map( A => n12887, B => n12886, S => n14468, Z => n15028
                           );
   U7498 : OAI211_X1 port map( C1 => n4631, C2 => n4630, A => n4629, B => n4628
                           , ZN => n20509);
   U7517 : INV_X1 port map( A => n19284, ZN => n20510);
   U7538 : BUF_X1 port map( A => n19092, Z => n19911);
   U7580 : XOR2_X1 port map( A => n6597, B => n6596, Z => n20511);
   U7582 : BUF_X1 port map( A => n17872, Z => n20512);
   U7660 : XNOR2_X1 port map( A => n15983, B => n15982, ZN => n17872);
   U7740 : NOR2_X2 port map( A1 => n129, A2 => n14291, ZN => n15896);
   U7741 : OR2_X1 port map( A1 => n19388, A2 => n19389, ZN => n651);
   U7794 : XNOR2_X1 port map( A => n15978, B => n15977, ZN => n20514);
   U7818 : OAI21_X1 port map( B1 => n17609, B2 => n19404, A => n17608, ZN => 
                           n20515);
   U7822 : OAI21_X1 port map( B1 => n17609, B2 => n19404, A => n17608, ZN => 
                           n19302);
   U7823 : XNOR2_X1 port map( A => n8172, B => n8173, ZN => n20516);
   U7841 : XNOR2_X1 port map( A => n8172, B => n8173, ZN => n1654);
   U7903 : XNOR2_X1 port map( A => n9789, B => n9790, ZN => n20517);
   U7985 : XNOR2_X1 port map( A => n10795, B => n10794, ZN => n14781);
   U8013 : BUF_X1 port map( A => n16577, Z => n20519);
   U8082 : MUX2_X1 port map( A => n9065, B => n8542, S => n9834, Z => n8074);
   U8111 : NAND2_X1 port map( A1 => n3785, A2 => n20520, ZN => n8128);
   U8144 : NAND3_X1 port map( A1 => n1452, A2 => n1453, A3 => n3784, ZN => 
                           n20520);
   U8170 : NAND2_X1 port map( A1 => n19737, A2 => n19658, ZN => n17553);
   U8184 : AND3_X2 port map( A1 => n2315, A2 => n7604, A3 => n7605, ZN => n8941
                           );
   U8265 : NAND2_X1 port map( A1 => n11465, A2 => n1514, ZN => n1513);
   U8272 : NAND3_X1 port map( A1 => n12393, A2 => n12394, A3 => n12396, ZN => 
                           n2539);
   U8282 : NOR2_X1 port map( A1 => n12237, A2 => n20523, ZN => n3762);
   U8291 : NAND2_X1 port map( A1 => n12606, A2 => n20524, ZN => n20523);
   U8326 : OAI21_X1 port map( B1 => n14070, B2 => n15505, A => n1758, ZN => 
                           n20525);
   U8337 : NAND2_X1 port map( A1 => n20526, A2 => n8189, ZN => n9221);
   U8339 : OR2_X1 port map( A1 => n8191, A2 => n8190, ZN => n20526);
   U8344 : NAND3_X1 port map( A1 => n5776, A2 => n5777, A3 => n1214, ZN => 
                           n5779);
   U8379 : NAND2_X1 port map( A1 => n1089, A2 => n13868, ZN => n3034);
   U8391 : XNOR2_X1 port map( A => n20527, B => n18209, ZN => Ciphertext(114));
   U8411 : NAND3_X1 port map( A1 => n18207, A2 => n18206, A3 => n20528, ZN => 
                           n20527);
   U8418 : INV_X1 port map( A => n2548, ZN => n3074);
   U8446 : AND2_X1 port map( A1 => n20529, A2 => n2548, ZN => n7441);
   U8488 : XNOR2_X2 port map( A => n7342, B => n7341, ZN => n2548);
   U8515 : INV_X1 port map( A => n7585, ZN => n20529);
   U8524 : NAND2_X1 port map( A1 => n20530, A2 => n9327, ZN => n9078);
   U8583 : OAI21_X1 port map( B1 => n20008, B2 => n9333, A => n9076, ZN => 
                           n20530);
   U8590 : OAI211_X2 port map( C1 => n3925, C2 => n4527, A => n4525, B => 
                           n20531, ZN => n5765);
   U8593 : NAND2_X1 port map( A1 => n4521, A2 => n3925, ZN => n20531);
   U8637 : NAND2_X1 port map( A1 => n2829, A2 => n19673, ZN => n2828);
   U8648 : NAND2_X1 port map( A1 => n3693, A2 => n18622, ZN => n2829);
   U8662 : NAND3_X1 port map( A1 => n1412, A2 => n15079, A3 => n20532, ZN => 
                           n16600);
   U8717 : NAND2_X1 port map( A1 => n15417, A2 => n20533, ZN => n20532);
   U8734 : INV_X1 port map( A => n15007, ZN => n20533);
   U8803 : XNOR2_X1 port map( A => n13817, B => n20378, ZN => n12286);
   U8846 : NAND2_X1 port map( A1 => n18131, A2 => n18130, ZN => n17556);
   U8927 : XNOR2_X2 port map( A => n17437, B => n17436, ZN => n18131);
   U8936 : NAND2_X1 port map( A1 => n1567, A2 => n8676, ZN => n8671);
   U8969 : NAND2_X1 port map( A1 => n4366, A2 => n4010, ZN => n4012);
   U8993 : XNOR2_X2 port map( A => n16703, B => n16704, ZN => n18966);
   U9113 : OAI21_X1 port map( B1 => n19488, B2 => n14011, A => n14611, ZN => 
                           n14013);
   U9123 : XNOR2_X2 port map( A => n12160, B => n12161, ZN => n19488);
   U9130 : AND3_X2 port map( A1 => n20021, A2 => n3392, A3 => n15663, ZN => 
                           n16295);
   U9132 : OAI21_X1 port map( B1 => n18051, B2 => n20535, A => n20534, ZN => 
                           n20052);
   U9219 : OR2_X1 port map( A1 => n18052, A2 => n19989, ZN => n20534);
   U9352 : INV_X1 port map( A => n19989, ZN => n20535);
   U9376 : NAND3_X1 port map( A1 => n20536, A2 => n7808, A3 => n8031, ZN => 
                           n1657);
   U9403 : NAND2_X1 port map( A1 => n463, A2 => n461, ZN => n20536);
   U9407 : NAND2_X1 port map( A1 => n20537, A2 => n18430, ZN => n18435);
   U9530 : NAND2_X1 port map( A1 => n3512, A2 => n18429, ZN => n20537);
   U9677 : OAI21_X1 port map( B1 => n18467, B2 => n20139, A => n17726, ZN => 
                           n18429);
   U9700 : OAI211_X1 port map( C1 => n19505, C2 => n19719, A => n20539, B => 
                           n20538, ZN => n2492);
   U9701 : NAND2_X1 port map( A1 => n19505, A2 => n3051, ZN => n20538);
   U9754 : AND2_X2 port map( A1 => n20541, A2 => n20540, ZN => n16963);
   U9757 : NAND2_X1 port map( A1 => n2279, A2 => n15687, ZN => n20540);
   U9765 : NAND2_X1 port map( A1 => n20542, A2 => n15454, ZN => n20541);
   U9789 : NAND2_X1 port map( A1 => n15450, A2 => n15451, ZN => n20542);
   U9812 : NAND3_X1 port map( A1 => n8703, A2 => n8155, A3 => n9567, ZN => 
                           n8170);
   U10002 : NAND2_X1 port map( A1 => n14260, A2 => n19652, ZN => n14265);
   U10005 : NAND2_X1 port map( A1 => n9053, A2 => n1752, ZN => n1750);
   U10058 : NAND2_X1 port map( A1 => n20544, A2 => n20543, ZN => n13103);
   U10095 : NAND2_X1 port map( A1 => n20626, A2 => n12593, ZN => n20544);
   U10102 : NAND2_X1 port map( A1 => n18341, A2 => n18344, ZN => n18290);
   U10218 : NAND2_X1 port map( A1 => n12060, A2 => n563, ZN => n12064);
   U10291 : NAND2_X1 port map( A1 => n20371, A2 => n20545, ZN => n14221);
   U10402 : NOR2_X1 port map( A1 => n15408, A2 => n15546, ZN => n20545);
   U10473 : NAND2_X1 port map( A1 => n8540, A2 => n2173, ZN => n10604);
   U10488 : NAND2_X1 port map( A1 => n14280, A2 => n14281, ZN => n14282);
   U10767 : NAND2_X1 port map( A1 => n14555, A2 => n14556, ZN => n14281);
   U10835 : INV_X1 port map( A => n5648, ZN => n5650);
   U10848 : NAND2_X1 port map( A1 => n5443, A2 => n5643, ZN => n5648);
   U10888 : INV_X1 port map( A => n8537, ZN => n8539);
   U10912 : NAND2_X1 port map( A1 => n8866, A2 => n9326, ZN => n8537);
   U11051 : NAND2_X1 port map( A1 => n13273, A2 => n20546, ZN => n13276);
   U11166 : INV_X1 port map( A => n20547, ZN => n20546);
   U11200 : OAI21_X1 port map( B1 => n13274, B2 => n13275, A => n13272, ZN => 
                           n20547);
   U11269 : NAND2_X1 port map( A1 => n900, A2 => n20548, ZN => n1584);
   U11270 : NAND2_X1 port map( A1 => n8245, A2 => n8251, ZN => n20548);
   U11356 : NAND2_X1 port map( A1 => n2018, A2 => n2019, ZN => n20549);
   U11363 : NAND2_X1 port map( A1 => n20072, A2 => n17507, ZN => n1899);
   U11425 : NAND3_X1 port map( A1 => n15042, A2 => n942, A3 => n15567, ZN => 
                           n1177);
   U11434 : AND2_X1 port map( A1 => n888, A2 => n11491, ZN => n11070);
   U11447 : NAND2_X1 port map( A1 => n16211, A2 => n20550, ZN => n17729);
   U11448 : NAND2_X1 port map( A1 => n17163, A2 => n17565, ZN => n20550);
   U11487 : OAI22_X1 port map( A1 => n18502, A2 => n18501, B1 => n18499, B2 => 
                           n18500, ZN => n1843);
   U11508 : NOR2_X1 port map( A1 => n15400, A2 => n15898, ZN => n15891);
   U11520 : NAND3_X1 port map( A1 => n4251, A2 => n19539, A3 => n4250, ZN => 
                           n99);
   U11522 : XNOR2_X1 port map( A => n20552, B => n20551, ZN => n7210);
   U11524 : NAND2_X1 port map( A1 => n3528, A2 => n20553, ZN => n20552);
   U11538 : NAND3_X1 port map( A1 => n8947, A2 => n8730, A3 => n8940, ZN => 
                           n20614);
   U11595 : AND2_X2 port map( A1 => n2319, A2 => n2360, ZN => n12095);
   U11617 : OR2_X1 port map( A1 => n8129, A2 => n1507, ZN => n8563);
   U11663 : OR2_X1 port map( A1 => n11035, A2 => n10783, ZN => n11437);
   U11693 : OAI21_X1 port map( B1 => n14598, B2 => n14395, A => n14596, ZN => 
                           n3757);
   U11694 : NAND2_X1 port map( A1 => n14154, A2 => n14393, ZN => n14596);
   U11755 : NAND2_X1 port map( A1 => n19652, A2 => n14261, ZN => n14543);
   U11788 : NAND2_X1 port map( A1 => n19404, A2 => n16306, ZN => n17607);
   U11790 : NAND3_X1 port map( A1 => n20306, A2 => n20307, A3 => n17688, ZN => 
                           n19034);
   U11792 : XNOR2_X1 port map( A => n20556, B => n20555, ZN => Ciphertext(70));
   U11873 : INV_X1 port map( A => n17989, ZN => n20555);
   U11923 : NAND3_X1 port map( A1 => n17988, A2 => n3829, A3 => n17987, ZN => 
                           n20556);
   U11924 : NAND2_X1 port map( A1 => n15110, A2 => n14461, ZN => n15292);
   U11980 : NOR2_X2 port map( A1 => n14471, A2 => n14470, ZN => n15110);
   U11993 : NAND2_X1 port map( A1 => n6950, A2 => n2961, ZN => n9164);
   U12032 : NAND2_X1 port map( A1 => n8609, A2 => n8696, ZN => n8610);
   U12052 : AND2_X2 port map( A1 => n2390, A2 => n2391, ZN => n14461);
   U12084 : NAND2_X1 port map( A1 => n8372, A2 => n8370, ZN => n7705);
   U12099 : NAND3_X1 port map( A1 => n8883, A2 => n8881, A3 => n8882, ZN => 
                           n20690);
   U12104 : XNOR2_X2 port map( A => n20558, B => n20557, ZN => n11231);
   U12109 : XNOR2_X1 port map( A => n9880, B => n10580, ZN => n20557);
   U12115 : XNOR2_X1 port map( A => n10004, B => n9877, ZN => n20558);
   U12116 : NAND3_X1 port map( A1 => n20559, A2 => n8557, A3 => n8558, ZN => 
                           n1186);
   U12128 : NAND2_X1 port map( A1 => n8556, A2 => n9107, ZN => n20559);
   U12146 : NAND2_X1 port map( A1 => n6133, A2 => n5691, ZN => n5692);
   U12191 : OAI21_X1 port map( B1 => n259, B2 => n20560, A => n20640, ZN => 
                           n11517);
   U12195 : NAND2_X1 port map( A1 => n10722, A2 => n20561, ZN => n12648);
   U12198 : NAND2_X1 port map( A1 => n9319, A2 => n1855, ZN => n9323);
   U12254 : OAI21_X1 port map( B1 => n15649, B2 => n15257, A => n20562, ZN => 
                           n14583);
   U12261 : NAND3_X1 port map( A1 => n15257, A2 => n15831, A3 => n20563, ZN => 
                           n20562);
   U12307 : INV_X1 port map( A => n15643, ZN => n20563);
   U12308 : AOI22_X1 port map( A1 => n20594, A2 => n7608, B1 => n8730, B2 => 
                           n8729, ZN => n7612);
   U12312 : INV_X1 port map( A => n5666, ZN => n20616);
   U12375 : NAND2_X1 port map( A1 => n17699, A2 => n18928, ZN => n1921);
   U12376 : NAND2_X1 port map( A1 => n20564, A2 => n19534, ZN => n19627);
   U12388 : NAND2_X1 port map( A1 => n19288, A2 => n19304, ZN => n20564);
   U12409 : NAND2_X1 port map( A1 => n15246, A2 => n20565, ZN => n15247);
   U12419 : NAND3_X2 port map( A1 => n5499, A2 => n20567, A3 => n20566, ZN => 
                           n7230);
   U12465 : NAND2_X1 port map( A1 => n1353, A2 => n5498, ZN => n20566);
   U12528 : NAND2_X1 port map( A1 => n5496, A2 => n20568, ZN => n20567);
   U12609 : NAND3_X1 port map( A1 => n15568, A2 => n20569, A3 => n20428, ZN => 
                           n15570);
   U12721 : NAND2_X1 port map( A1 => n15565, A2 => n15804, ZN => n20569);
   U12737 : NAND2_X1 port map( A1 => n3712, A2 => n3713, ZN => n11222);
   U12878 : AND2_X2 port map( A1 => n20570, A2 => n3646, ZN => n13624);
   U12880 : NAND2_X1 port map( A1 => n2804, A2 => n3649, ZN => n20570);
   U12885 : OAI21_X1 port map( B1 => n20382, B2 => n20571, A => n19434, ZN => 
                           n20316);
   U12989 : NAND2_X1 port map( A1 => n20574, A2 => n20572, ZN => n19378);
   U12993 : NAND2_X1 port map( A1 => n20573, A2 => n19375, ZN => n20572);
   U13100 : NAND2_X1 port map( A1 => n19374, A2 => n19733, ZN => n20573);
   U13172 : NAND2_X1 port map( A1 => n19377, A2 => n19666, ZN => n20574);
   U13410 : OR2_X1 port map( A1 => n15453, A2 => n19978, ZN => n15786);
   U13512 : NAND3_X1 port map( A1 => n1329, A2 => n1327, A3 => n20575, ZN => 
                           n12543);
   U13541 : NAND3_X1 port map( A1 => n20660, A2 => n764, A3 => n11383, ZN => 
                           n20575);
   U13585 : XNOR2_X1 port map( A => n20576, B => n2395, ZN => Ciphertext(170));
   U13588 : NAND3_X1 port map( A1 => n18166, A2 => n2226, A3 => n2227, ZN => 
                           n20576);
   U13698 : NAND2_X1 port map( A1 => n19881, A2 => n8375, ZN => n6733);
   U13723 : NAND2_X1 port map( A1 => n20577, A2 => n12098, ZN => n13065);
   U13754 : NOR2_X1 port map( A1 => n20579, A2 => n20578, ZN => n20577);
   U13758 : NOR2_X1 port map( A1 => n12428, A2 => n3649, ZN => n20578);
   U13777 : INV_X1 port map( A => n12097, ZN => n20579);
   U13810 : NOR2_X1 port map( A1 => n13742, A2 => n13743, ZN => n15677);
   U13863 : NAND2_X1 port map( A1 => n18653, A2 => n18654, ZN => n20580);
   U13868 : NAND2_X1 port map( A1 => n18655, A2 => n18656, ZN => n20581);
   U13885 : XNOR2_X1 port map( A => n20582, B => n18148, ZN => Ciphertext(59));
   U13934 : NAND4_X1 port map( A1 => n20629, A2 => n2830, A3 => n2828, A4 => 
                           n18147, ZN => n20582);
   U13936 : NAND2_X1 port map( A1 => n9529, A2 => n9528, ZN => n9527);
   U14000 : NAND2_X1 port map( A1 => n8721, A2 => n9357, ZN => n9529);
   U14001 : NAND2_X1 port map( A1 => n19511, A2 => n19395, ZN => n19631);
   U14021 : NAND3_X1 port map( A1 => n1459, A2 => n3104, A3 => n20583, ZN => 
                           n12047);
   U14064 : OAI21_X1 port map( B1 => n20585, B2 => n20584, A => n585, ZN => 
                           n20035);
   U14073 : OAI21_X1 port map( B1 => n11282, B2 => n11281, A => n20641, ZN => 
                           n1498);
   U14075 : NAND3_X1 port map( A1 => n18319, A2 => n19174, A3 => n1035, ZN => 
                           n18322);
   U14246 : NAND2_X1 port map( A1 => n88, A2 => n8075, ZN => n10552);
   U14262 : OR2_X1 port map( A1 => n19185, A2 => n20642, ZN => n19186);
   U14342 : NAND2_X1 port map( A1 => n20586, A2 => n8209, ZN => n7434);
   U14346 : NAND2_X1 port map( A1 => n9006, A2 => n8890, ZN => n1672);
   U14391 : NAND2_X1 port map( A1 => n20589, A2 => n20587, ZN => n7997);
   U14415 : NAND2_X1 port map( A1 => n7989, A2 => n20588, ZN => n20587);
   U14446 : INV_X1 port map( A => n8705, ZN => n20588);
   U14482 : NAND2_X1 port map( A1 => n7988, A2 => n8705, ZN => n20589);
   U14497 : NAND3_X2 port map( A1 => n15542, A2 => n15541, A3 => n20379, ZN => 
                           n16181);
   U14530 : OAI21_X1 port map( B1 => n11187, B2 => n20591, A => n20590, ZN => 
                           n11196);
   U14562 : NAND2_X1 port map( A1 => n11189, A2 => n19983, ZN => n20590);
   U14563 : NAND2_X1 port map( A1 => n20592, A2 => n2981, ZN => n2980);
   U14589 : NAND2_X1 port map( A1 => n18145, A2 => n18641, ZN => n20592);
   U14716 : NAND3_X1 port map( A1 => n6051, A2 => n6052, A3 => n6050, ZN => 
                           n6053);
   U14717 : NAND2_X1 port map( A1 => n11637, A2 => n20430, ZN => n11979);
   U14724 : NAND2_X1 port map( A1 => n19879, A2 => n15666, ZN => n15771);
   U14728 : NAND2_X1 port map( A1 => n722, A2 => n723, ZN => n721);
   U14823 : NOR2_X1 port map( A1 => n317, A2 => n8945, ZN => n20594);
   U14826 : OR2_X1 port map( A1 => n11528, A2 => n11526, ZN => n20279);
   U14878 : NAND2_X1 port map( A1 => n10863, A2 => n11387, ZN => n10867);
   U14890 : OAI211_X1 port map( C1 => n11544, C2 => n11549, A => n20595, B => 
                           n11550, ZN => n10762);
   U15069 : NAND2_X1 port map( A1 => n11544, A2 => n10926, ZN => n20595);
   U15088 : NAND2_X1 port map( A1 => n20596, A2 => n8057, ZN => n2750);
   U15131 : OAI211_X1 port map( C1 => n8054, C2 => n19802, A => n3472, B => 
                           n8052, ZN => n20596);
   U15133 : XNOR2_X2 port map( A => n20598, B => n20597, ZN => n11546);
   U15134 : XNOR2_X1 port map( A => n9261, B => n8635, ZN => n20597);
   U15174 : XNOR2_X1 port map( A => n8627, B => n9508, ZN => n20598);
   U15203 : NAND3_X1 port map( A1 => n1232, A2 => n4814, A3 => n5069, ZN => 
                           n19612);
   U15294 : NAND2_X1 port map( A1 => n20600, A2 => n20599, ZN => n10991);
   U15314 : NAND2_X1 port map( A1 => n11870, A2 => n11390, ZN => n20599);
   U15325 : NAND2_X1 port map( A1 => n20160, A2 => n20601, ZN => n20600);
   U15369 : INV_X1 port map( A => n11389, ZN => n20601);
   U15370 : NAND2_X1 port map( A1 => n16659, A2 => n1115, ZN => n16661);
   U15399 : NAND2_X1 port map( A1 => n10653, A2 => n20375, ZN => n11602);
   U15546 : NAND2_X1 port map( A1 => n19679, A2 => n19757, ZN => n18216);
   U15576 : OAI21_X1 port map( B1 => n16780, B2 => n19143, A => n20602, ZN => 
                           n17810);
   U15621 : NAND2_X1 port map( A1 => n16780, A2 => n19135, ZN => n20602);
   U15669 : NAND2_X1 port map( A1 => n5141, A2 => n20603, ZN => n5143);
   U15717 : NAND3_X1 port map( A1 => n6054, A2 => n5139, A3 => n5559, ZN => 
                           n20603);
   U15726 : OAI21_X1 port map( B1 => n12184, B2 => n12185, A => n20604, ZN => 
                           n12745);
   U15731 : NAND2_X1 port map( A1 => n20201, A2 => n12181, ZN => n20604);
   U15776 : NAND3_X1 port map( A1 => n9169, A2 => n9170, A3 => n1211, ZN => 
                           n10329);
   U15778 : XNOR2_X1 port map( A => n20605, B => n2193, ZN => Ciphertext(126));
   U15795 : NAND3_X1 port map( A1 => n2196, A2 => n2197, A3 => n2195, ZN => 
                           n20605);
   U15802 : AOI22_X1 port map( A1 => n12066, A2 => n12213, B1 => n12210, B2 => 
                           n12189, ZN => n12068);
   U15807 : NAND2_X1 port map( A1 => n236, A2 => n20451, ZN => n14412);
   U15812 : NAND3_X1 port map( A1 => n20645, A2 => n4384, A3 => n20606, ZN => 
                           n3684);
   U15857 : NAND2_X1 port map( A1 => n905, A2 => n8741, ZN => n8951);
   U15947 : OR2_X1 port map( A1 => n7629, A2 => n7630, ZN => n905);
   U15982 : NAND2_X1 port map( A1 => n14285, A2 => n20607, ZN => n1437);
   U16003 : NOR2_X1 port map( A1 => n14296, A2 => n15898, ZN => n20607);
   U16004 : NAND3_X1 port map( A1 => n8929, A2 => n8931, A3 => n8933, ZN => 
                           n8935);
   U16082 : XNOR2_X1 port map( A => n9792, B => n20608, ZN => n9796);
   U16095 : NAND2_X1 port map( A1 => n11632, A2 => n11633, ZN => n12616);
   U16096 : NOR2_X1 port map( A1 => n20040, A2 => n14817, ZN => n20609);
   U16101 : OAI211_X1 port map( C1 => n20437, C2 => n20361, A => n18384, B => 
                           n20610, ZN => n595);
   U16102 : NAND2_X1 port map( A1 => n20361, A2 => n20611, ZN => n20610);
   U16110 : NAND3_X1 port map( A1 => n4641, A2 => n4646, A3 => n4647, ZN => 
                           n4148);
   U16122 : NAND2_X1 port map( A1 => n18028, A2 => n18931, ZN => n20612);
   U16123 : NAND2_X1 port map( A1 => n18027, A2 => n20207, ZN => n20613);
   U16134 : NAND2_X1 port map( A1 => n20614, A2 => n318, ZN => n8948);
   U16137 : OR2_X1 port map( A1 => n5116, A2 => n5115, ZN => n1914);
   U16155 : NAND2_X1 port map( A1 => n1575, A2 => n9452, ZN => n8885);
   U16185 : NAND2_X1 port map( A1 => n5665, A2 => n20615, ZN => n6735);
   U16203 : NAND2_X1 port map( A1 => n20616, A2 => n5661, ZN => n20615);
   U16269 : NAND2_X2 port map( A1 => n20617, A2 => n3758, ZN => n15275);
   U16277 : NAND2_X1 port map( A1 => n3757, A2 => n14394, ZN => n20617);
   U16278 : NAND2_X1 port map( A1 => n12153, A2 => n20486, ZN => n12149);
   U16313 : NAND3_X1 port map( A1 => n2437, A2 => n15444, A3 => n2438, ZN => 
                           n20032);
   U16318 : OAI211_X2 port map( C1 => n20235, C2 => n9612, A => n20620, B => 
                           n20619, ZN => n11951);
   U16348 : NAND2_X1 port map( A1 => n9609, A2 => n11292, ZN => n20619);
   U16350 : NAND2_X1 port map( A1 => n9610, A2 => n11404, ZN => n20620);
   U16351 : NAND3_X1 port map( A1 => n20621, A2 => n15226, A3 => n15779, ZN => 
                           n14870);
   U16365 : NAND2_X1 port map( A1 => n15685, A2 => n15783, ZN => n20621);
   U16366 : OR2_X1 port map( A1 => n7952, A2 => n7481, ZN => n7814);
   U16381 : AOI22_X2 port map( A1 => n19387, A2 => n19386, B1 => n19385, B2 => 
                           n19384, ZN => n19442);
   U16408 : NOR2_X1 port map( A1 => n11903, A2 => n12148, ZN => n11904);
   U16409 : NOR2_X2 port map( A1 => n11345, A2 => n11344, ZN => n12148);
   U16410 : NAND2_X1 port map( A1 => n3451, A2 => n5074, ZN => n4459);
   U16423 : NAND2_X1 port map( A1 => n3270, A2 => n3272, ZN => n447);
   U16476 : AND2_X2 port map( A1 => n20623, A2 => n20622, ZN => n13321);
   U16560 : NAND2_X1 port map( A1 => n11063, A2 => n12267, ZN => n20622);
   U16566 : NAND2_X1 port map( A1 => n9059, A2 => n9031, ZN => n8573);
   U16580 : NAND3_X1 port map( A1 => n18749, A2 => n18711, A3 => n18773, ZN => 
                           n18712);
   U16596 : NAND2_X1 port map( A1 => n8712, A2 => n9233, ZN => n8412);
   U16601 : NOR2_X1 port map( A1 => n19716, A2 => n9234, ZN => n8712);
   U16640 : NAND2_X1 port map( A1 => n20625, A2 => n1929, ZN => n10567);
   U16645 : OAI22_X1 port map( A1 => n8673, A2 => n8674, B1 => n9021, B2 => 
                           n8676, ZN => n20625);
   U16681 : NOR2_X2 port map( A1 => n9184, A2 => n9185, ZN => n10571);
   U16687 : NAND2_X1 port map( A1 => n11979, A2 => n11978, ZN => n20626);
   U16707 : AOI22_X2 port map( A1 => n8759, A2 => n9273, B1 => n20627, B2 => 
                           n8991, ZN => n9894);
   U16708 : OAI21_X1 port map( B1 => n9277, B2 => n9275, A => n19732, ZN => 
                           n20627);
   U16709 : NAND2_X1 port map( A1 => n20628, A2 => n2294, ZN => n6942);
   U16725 : NAND2_X1 port map( A1 => n3700, A2 => n5751, ZN => n20628);
   U16726 : NAND2_X1 port map( A1 => n20039, A2 => n2829, ZN => n20629);
   U16764 : NAND2_X1 port map( A1 => n12065, A2 => n12211, ZN => n11814);
   U16766 : OAI211_X2 port map( C1 => n5980, C2 => n5155, A => n5153, B => 
                           n20630, ZN => n7232);
   U16771 : NAND2_X1 port map( A1 => n3767, A2 => n6075, ZN => n20630);
   U16778 : XNOR2_X1 port map( A => n20631, B => n18316, ZN => Ciphertext(177))
                           ;
   U17000 : NAND2_X1 port map( A1 => n18315, A2 => n20632, ZN => n20631);
   U17016 : AND2_X1 port map( A1 => n18314, A2 => n18313, ZN => n20632);
   U17017 : NAND2_X1 port map( A1 => n20634, A2 => n20633, ZN => n15026);
   U17111 : XNOR2_X2 port map( A => n14971, B => n14970, ZN => n17208);
   U17192 : NAND2_X1 port map( A1 => n16465, A2 => n17210, ZN => n20634);
   U17193 : AND3_X2 port map( A1 => n10762, A2 => n10763, A3 => n10764, ZN => 
                           n12389);
   U17194 : INV_X1 port map( A => Plaintext(56), ZN => n20635);
   U17198 : NAND2_X1 port map( A1 => n14515, A2 => n20636, ZN => n15125);
   U17239 : OAI22_X1 port map( A1 => n7861, A2 => n8083, B1 => n20638, B2 => 
                           n20637, ZN => n1159);
   U17265 : INV_X1 port map( A => n20495, ZN => n20637);
   U17341 : NAND2_X1 port map( A1 => n6539, A2 => n20108, ZN => n20638);
   U17392 : NAND3_X1 port map( A1 => n20640, A2 => n10936, A3 => n20639, ZN => 
                           n725);
   U17396 : INV_X1 port map( A => n11573, ZN => n20639);
   U17431 : INV_X1 port map( A => n20106, ZN => n20640);
   U17432 : NAND2_X1 port map( A1 => n14624, A2 => n14627, ZN => n13856);
   U17498 : NAND2_X1 port map( A1 => n15474, A2 => n12659, ZN => n12662);
   U17514 : NOR2_X1 port map( A1 => n19183, A2 => n19212, ZN => n20642);
   U17568 : XNOR2_X1 port map( A => n20643, B => n18717, ZN => Ciphertext(78));
   U17659 : NAND4_X1 port map( A1 => n18714, A2 => n18713, A3 => n18715, A4 => 
                           n18712, ZN => n20643);
   U17662 : XNOR2_X1 port map( A => n13138, B => n13339, ZN => n13139);
   U17686 : AOI21_X2 port map( B1 => n11696, B2 => n12399, A => n20644, ZN => 
                           n13339);
   U17749 : OAI211_X2 port map( C1 => n14753, C2 => n14430, A => n14428, B => 
                           n14429, ZN => n15296);
   U17750 : NAND2_X1 port map( A1 => n4480, A2 => n3967, ZN => n20645);
   U17751 : NAND2_X1 port map( A1 => n12473, A2 => n19833, ZN => n12484);
   U17793 : NAND2_X1 port map( A1 => n20058, A2 => n20060, ZN => n19492);
   U17800 : XNOR2_X1 port map( A => n20664, B => n13300, ZN => n14707);
   U17833 : NOR2_X1 port map( A1 => n15679, A2 => n20647, ZN => n15231);
   U18067 : INV_X1 port map( A => n16165, ZN => n20648);
   U18128 : NAND2_X1 port map( A1 => n17498, A2 => n15485, ZN => n16795);
   U18308 : XNOR2_X2 port map( A => n10440, B => n10439, ZN => n11445);
   U18337 : NAND2_X1 port map( A1 => n343, A2 => n6097, ZN => n20649);
   U18353 : NAND2_X1 port map( A1 => n20689, A2 => n789, ZN => n787);
   U18386 : NAND3_X1 port map( A1 => n138, A2 => n1775, A3 => n1772, ZN => n137
                           );
   U18392 : NAND3_X1 port map( A1 => n267, A2 => n266, A3 => n9242, ZN => n3288
                           );
   U18394 : OAI211_X2 port map( C1 => n8431, C2 => n9218, A => n8429, B => 
                           n8430, ZN => n10072);
   U18401 : NAND3_X1 port map( A1 => n7587, A2 => n7588, A3 => n20650, ZN => 
                           n8644);
   U18459 : NAND2_X1 port map( A1 => n20373, A2 => n20651, ZN => n20650);
   U18476 : NAND2_X1 port map( A1 => n7603, A2 => n7795, ZN => n7605);
   U18482 : NAND2_X1 port map( A1 => n19403, A2 => n19402, ZN => n17649);
   U18490 : OAI211_X2 port map( C1 => n15890, C2 => n14913, A => n14911, B => 
                           n20652, ZN => n17378);
   U18555 : NAND2_X1 port map( A1 => n15890, A2 => n20006, ZN => n20652);
   U18633 : NAND3_X1 port map( A1 => n14666, A2 => n14535, A3 => n14662, ZN => 
                           n14313);
   U18634 : XNOR2_X2 port map( A => n13177, B => n13176, ZN => n14662);
   U18636 : NAND2_X1 port map( A1 => n20367, A2 => n7953, ZN => n7818);
   U18655 : NAND2_X1 port map( A1 => n14623, A2 => n14626, ZN => n14625);
   U18683 : NAND3_X1 port map( A1 => n20653, A2 => n12919, A3 => n14443, ZN => 
                           n2775);
   U18684 : NAND2_X1 port map( A1 => n14439, A2 => n14168, ZN => n20653);
   U18698 : INV_X1 port map( A => n18500, ZN => n17737);
   U18706 : NAND2_X2 port map( A1 => n816, A2 => n20654, ZN => n18500);
   U18751 : NAND2_X1 port map( A1 => n4422, A2 => n20655, ZN => n6119);
   U18766 : NAND2_X1 port map( A1 => n12129, A2 => n11586, ZN => n699);
   U18778 : NAND2_X1 port map( A1 => n3487, A2 => n3488, ZN => n12129);
   U18827 : OR2_X1 port map( A1 => n6138, A2 => n5859, ZN => n20333);
   U18829 : OAI21_X1 port map( B1 => n7836, B2 => n7958, A => n20656, ZN => 
                           n8911);
   U18830 : NAND2_X1 port map( A1 => n20165, A2 => n7836, ZN => n20656);
   U18853 : AOI21_X1 port map( B1 => n5900, B2 => n6087, A => n5908, ZN => 
                           n1466);
   U18899 : OAI22_X2 port map( A1 => n1164, A2 => n7283, B1 => n7812, B2 => 
                           n7811, ZN => n8890);
   U18932 : NAND2_X1 port map( A1 => n6155, A2 => n5612, ZN => n5610);
   U18935 : OAI211_X2 port map( C1 => n7992, C2 => n8015, A => n20657, B => 
                           n7472, ZN => n8813);
   U18944 : NAND2_X1 port map( A1 => n3243, A2 => n7994, ZN => n20657);
   U18959 : NAND2_X1 port map( A1 => n1902, A2 => n2970, ZN => n12036);
   U18962 : NAND2_X1 port map( A1 => n14572, A2 => n14573, ZN => n14741);
   U19077 : AND2_X2 port map( A1 => n20658, A2 => n3672, ZN => n6410);
   U19087 : NAND2_X1 port map( A1 => n4502, A2 => n3674, ZN => n20658);
   U19088 : NAND2_X1 port map( A1 => n8734, A2 => n8923, ZN => n8498);
   U19109 : NAND2_X1 port map( A1 => n45, A2 => n44, ZN => n8);
   U19125 : AND3_X2 port map( A1 => n15833, A2 => n15834, A3 => n15835, ZN => 
                           n16975);
   U19126 : NAND3_X1 port map( A1 => n19911, A2 => n17529, A3 => n20661, ZN => 
                           n17532);
   U19128 : NAND2_X1 port map( A1 => n4147, A2 => n4148, ZN => n4149);
   U19209 : NAND3_X1 port map( A1 => n2492, A2 => n20663, A3 => n20662, ZN => 
                           n12513);
   U19398 : NAND2_X1 port map( A1 => n10623, A2 => n888, ZN => n20662);
   U19406 : NAND2_X1 port map( A1 => n3814, A2 => n913, ZN => n20663);
   U19407 : OAI22_X1 port map( A1 => n11911, A2 => n12812, B1 => n11912, B2 => 
                           n12490, ZN => n11913);
   U19474 : NAND2_X1 port map( A1 => n3586, A2 => n12807, ZN => n11911);
   U19487 : XNOR2_X1 port map( A => n6563, B => n7117, ZN => n3570);
   U19518 : INV_X1 port map( A => n16465, ZN => n16660);
   U19519 : XNOR2_X2 port map( A => n14995, B => n14994, ZN => n16465);
   U19520 : NOR2_X2 port map( A1 => n14445, A2 => n1722, ZN => n15294);
   U19542 : INV_X1 port map( A => n14998, ZN => n15832);
   U19543 : NAND2_X1 port map( A1 => n15828, A2 => n19891, ZN => n14998);
   U19544 : XNOR2_X1 port map( A => n13463, B => n13298, ZN => n20664);
   U19589 : NAND3_X1 port map( A1 => n14339, A2 => n14049, A3 => n20665, ZN => 
                           n12802);
   U19601 : NAND2_X1 port map( A1 => n14335, A2 => n13930, ZN => n14049);
   U19605 : NAND2_X1 port map( A1 => n15469, A2 => n15465, ZN => n15340);
   U19625 : NAND2_X1 port map( A1 => n20666, A2 => n8869, ZN => n8465);
   U19626 : NAND2_X1 port map( A1 => n9326, A2 => n9076, ZN => n20666);
   U19655 : AOI22_X2 port map( A1 => n2109, A2 => n15343, B1 => n15342, B2 => 
                           n19888, ZN => n19889);
   U19675 : NAND2_X1 port map( A1 => n1507, A2 => n20010, ZN => n1652);
   U19684 : NOR2_X2 port map( A1 => n6320, A2 => n6319, ZN => n20010);
   U19703 : NAND2_X1 port map( A1 => n15990, A2 => n20667, ZN => n15591);
   U19704 : NAND3_X1 port map( A1 => n1469, A2 => n13959, A3 => n13960, ZN => 
                           n20119);
   U19713 : NAND2_X1 port map( A1 => n14666, A2 => n14663, ZN => n14314);
   U19744 : NAND3_X1 port map( A1 => n6055, A2 => n20669, A3 => n20668, ZN => 
                           n385);
   U19750 : NAND2_X1 port map( A1 => n6057, A2 => n5891, ZN => n20668);
   U19767 : NAND2_X1 port map( A1 => n906, A2 => n20670, ZN => n20669);
   U19777 : INV_X1 port map( A => n5304, ZN => n20670);
   U19790 : NAND2_X1 port map( A1 => n20358, A2 => n7932, ZN => n7760);
   U19794 : NAND2_X1 port map( A1 => n12507, A2 => n12506, ZN => n1609);
   U19806 : NAND3_X1 port map( A1 => n11019, A2 => n11020, A3 => n12500, ZN => 
                           n11021);
   U19807 : NAND3_X1 port map( A1 => n20299, A2 => n1378, A3 => n20300, ZN => 
                           n20671);
   U19819 : AND2_X2 port map( A1 => n20683, A2 => n20684, ZN => n9039);
   U19823 : NAND2_X1 port map( A1 => n5623, A2 => n6129, ZN => n1770);
   U19825 : AOI21_X2 port map( B1 => n4279, B2 => n3682, A => n19559, ZN => 
                           n5623);
   U19828 : OAI21_X1 port map( B1 => n20674, B2 => n5525, A => n20673, ZN => 
                           n1170);
   U19835 : INV_X1 port map( A => n5294, ZN => n20673);
   U19840 : NAND2_X1 port map( A1 => n19201, A2 => n19842, ZN => n19193);
   U19845 : NAND2_X1 port map( A1 => n20675, A2 => n11326, ZN => n11709);
   U19856 : OAI21_X1 port map( B1 => n1124, B2 => n191, A => n1122, ZN => 
                           n20675);
   U19858 : NAND2_X1 port map( A1 => n2246, A2 => n66, ZN => n2814);
   U19859 : INV_X1 port map( A => n20676, ZN => n19974);
   U19860 : XNOR2_X1 port map( A => n17415, B => n17414, ZN => n20676);
   U19861 : AND3_X2 port map( A1 => n15528, A2 => n1337, A3 => n16443, ZN => 
                           n15529);
   U19862 : NAND3_X1 port map( A1 => n4736, A2 => n3903, A3 => n4737, ZN => 
                           n3905);
   U19863 : NAND2_X1 port map( A1 => n679, A2 => n2049, ZN => n678);
   U19864 : NAND2_X1 port map( A1 => n3031, A2 => n18869, ZN => n679);
   U19865 : XNOR2_X2 port map( A => n7387, B => n7388, ZN => n8289);
   U19866 : NOR2_X2 port map( A1 => n11084, A2 => n11085, ZN => n13147);
   U19867 : INV_X1 port map( A => n20677, ZN => n1894);
   U19868 : OAI21_X1 port map( B1 => n6037, B2 => n6036, A => n6035, ZN => 
                           n20677);
   U19869 : NAND3_X1 port map( A1 => n2166, A2 => n1416, A3 => n2165, ZN => 
                           n8833);
   U19870 : NAND2_X1 port map( A1 => n1642, A2 => n420, ZN => n14735);
   U19871 : NAND2_X1 port map( A1 => n4460, A2 => n20431, ZN => n3189);
   U19872 : NAND2_X1 port map( A1 => n14742, A2 => n14743, ZN => n14745);
   U19873 : AOI21_X1 port map( B1 => n20678, B2 => n7920, A => n7768, ZN => 
                           n6320);
   U19874 : NAND2_X1 port map( A1 => n6299, A2 => n505, ZN => n20678);
   U19875 : NAND2_X1 port map( A1 => n19301, A2 => n20515, ZN => n19303);
   U19876 : OAI21_X1 port map( B1 => n20381, B2 => n14501, A => n20680, ZN => 
                           n14504);
   U19877 : NAND2_X1 port map( A1 => n14502, A2 => n14501, ZN => n20680);
   U19878 : OR2_X1 port map( A1 => n11546, A2 => n10761, ZN => n20681);
   U19879 : INV_X1 port map( A => n4043, ZN => n1442);
   U19880 : NAND3_X1 port map( A1 => n4042, A2 => n713, A3 => n5034, ZN => 
                           n4043);
   U19881 : NAND2_X1 port map( A1 => n9039, A2 => n8851, ZN => n9045);
   U19882 : NAND2_X1 port map( A1 => n7402, A2 => n7171, ZN => n20683);
   U19883 : NAND2_X1 port map( A1 => n7170, A2 => n7814, ZN => n20684);
   U19884 : NAND3_X1 port map( A1 => n20685, A2 => n2116, A3 => n8984, ZN => 
                           n1157);
   U19885 : NAND2_X1 port map( A1 => n9267, A2 => n2118, ZN => n20685);
   U19886 : OAI211_X2 port map( C1 => n9051, C2 => n9289, A => n20686, B => 
                           n839, ZN => n9824);
   U19887 : NAND2_X1 port map( A1 => n736, A2 => n19896, ZN => n20686);
   U19888 : NAND2_X1 port map( A1 => n2102, A2 => n2103, ZN => n2101);
   U19889 : XNOR2_X1 port map( A => n20687, B => n19273, ZN => Ciphertext(166))
                           ;
   U19890 : NAND3_X1 port map( A1 => n2262, A2 => n2261, A3 => n19272, ZN => 
                           n20687);
   U19891 : NAND2_X1 port map( A1 => n6049, A2 => n6048, ZN => n2641);
   U19892 : OAI211_X2 port map( C1 => n4509, C2 => n4574, A => n3909, B => 
                           n3910, ZN => n6048);
   U19893 : NAND2_X2 port map( A1 => n12459, A2 => n12460, ZN => n12137);
   U19894 : NAND2_X1 port map( A1 => n1943, A2 => n1944, ZN => n12459);
   U19895 : NAND2_X1 port map( A1 => n17968, A2 => n19943, ZN => n2951);
   U19896 : NAND2_X1 port map( A1 => n17558, A2 => n18114, ZN => n17968);
   U19897 : NAND2_X1 port map( A1 => n20338, A2 => n12104, ZN => n1854);
   U19898 : XNOR2_X2 port map( A => n6758, B => n6757, ZN => n8387);
   U19899 : NAND2_X1 port map( A1 => n20688, A2 => n14149, ZN => n14152);
   U19900 : NAND2_X1 port map( A1 => n14400, A2 => n14401, ZN => n20688);
   U19901 : NAND2_X1 port map( A1 => n2840, A2 => n7551, ZN => n7552);
   U19902 : OR2_X1 port map( A1 => n11376, A2 => n11330, ZN => n1853);
   U19903 : INV_X1 port map( A => n15891, ZN => n20689);
   U19904 : NAND3_X1 port map( A1 => n360, A2 => n197, A3 => n15059, ZN => 
                           n14988);
   U19905 : AND3_X2 port map( A1 => n1700, A2 => n1697, A3 => n1696, ZN => 
                           n15256);
   U19906 : OAI21_X1 port map( B1 => n20374, B2 => n20691, A => n8209, ZN => 
                           n1910);
   U19907 : NOR2_X1 port map( A1 => n8095, A2 => n7631, ZN => n20691);
   U19908 : XNOR2_X1 port map( A => n20692, B => n18379, ZN => Ciphertext(7));
   U19909 : NAND2_X1 port map( A1 => n18378, A2 => n20693, ZN => n20692);
   U19910 : OR2_X1 port map( A1 => n18393, A2 => n1296, ZN => n20693);
   U19911 : XNOR2_X1 port map( A => n13632, B => n13633, ZN => n13639);
   U19912 : NAND2_X1 port map( A1 => n20362, A2 => n15686, ZN => n15453);
   U19913 : NAND2_X1 port map( A1 => n5520, A2 => n5927, ZN => n5193);
   U19914 : NAND2_X1 port map( A1 => n4809, A2 => n4810, ZN => n4813);
   U19915 : NAND2_X1 port map( A1 => n5074, A2 => n20431, ZN => n4810);
   U19916 : NAND2_X1 port map( A1 => n1831, A2 => n8660, ZN => n1830);
   U19917 : NAND2_X1 port map( A1 => n13053, A2 => n20694, ZN => n13055);
   U19918 : NAND3_X1 port map( A1 => n14307, A2 => n19940, A3 => n13040, ZN => 
                           n20694);
   U19919 : OAI211_X1 port map( C1 => n12275, C2 => n12028, A => n11782, B => 
                           n20695, ZN => n2366);
   U19920 : NAND2_X1 port map( A1 => n12275, A2 => n12029, ZN => n20695);
   U19921 : AND3_X2 port map( A1 => n20696, A2 => n1424, A3 => n449, ZN => 
                           n9172);
   U19922 : NAND2_X1 port map( A1 => n836, A2 => n837, ZN => n20696);
   U19923 : OAI21_X1 port map( B1 => n8616, B2 => n8763, A => n20697, ZN => 
                           n20054);
   U19924 : INV_X1 port map( A => n8693, ZN => n20697);
   U19925 : XNOR2_X2 port map( A => n13197, B => n13196, ZN => n20266);
   U19926 : BUF_X2 port map( A => n17349, Z => n19836);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Top is

   port( clk : in std_logic;  Plaintext, Key : in std_logic_vector (191 downto 
         0);  Ciphertext : out std_logic_vector (191 downto 0));

end SPEEDY_Top;

architecture SYN_Behavioral of SPEEDY_Top is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SPEEDY_Rounds5_0
      port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : 
            out std_logic_vector (191 downto 0));
   end component;
   
   signal reg_in_191_port, reg_in_190_port, reg_in_189_port, reg_in_188_port, 
      reg_in_187_port, reg_in_186_port, reg_in_185_port, reg_in_184_port, 
      reg_in_183_port, reg_in_182_port, reg_in_181_port, reg_in_180_port, 
      reg_in_179_port, reg_in_178_port, reg_in_177_port, reg_in_176_port, 
      reg_in_175_port, reg_in_174_port, reg_in_173_port, reg_in_172_port, 
      reg_in_171_port, reg_in_170_port, reg_in_169_port, reg_in_168_port, 
      reg_in_167_port, reg_in_166_port, reg_in_165_port, reg_in_164_port, 
      reg_in_163_port, reg_in_162_port, reg_in_161_port, reg_in_160_port, 
      reg_in_159_port, reg_in_158_port, reg_in_157_port, reg_in_156_port, 
      reg_in_155_port, reg_in_154_port, reg_in_153_port, reg_in_152_port, 
      reg_in_151_port, reg_in_150_port, reg_in_149_port, reg_in_148_port, 
      reg_in_147_port, reg_in_146_port, reg_in_145_port, reg_in_144_port, 
      reg_in_143_port, reg_in_142_port, reg_in_141_port, reg_in_140_port, 
      reg_in_139_port, reg_in_138_port, reg_in_137_port, reg_in_136_port, 
      reg_in_135_port, reg_in_134_port, reg_in_133_port, reg_in_132_port, 
      reg_in_131_port, reg_in_130_port, reg_in_129_port, reg_in_128_port, 
      reg_in_127_port, reg_in_126_port, reg_in_125_port, reg_in_124_port, 
      reg_in_123_port, reg_in_122_port, reg_in_121_port, reg_in_120_port, 
      reg_in_119_port, reg_in_118_port, reg_in_117_port, reg_in_116_port, 
      reg_in_115_port, reg_in_114_port, reg_in_113_port, reg_in_112_port, 
      reg_in_111_port, reg_in_110_port, reg_in_109_port, reg_in_108_port, 
      reg_in_107_port, reg_in_106_port, reg_in_105_port, reg_in_104_port, 
      reg_in_103_port, reg_in_102_port, reg_in_101_port, reg_in_100_port, 
      reg_in_99_port, reg_in_98_port, reg_in_97_port, reg_in_96_port, 
      reg_in_95_port, reg_in_94_port, reg_in_93_port, reg_in_92_port, 
      reg_in_91_port, reg_in_90_port, reg_in_89_port, reg_in_88_port, 
      reg_in_87_port, reg_in_86_port, reg_in_85_port, reg_in_84_port, 
      reg_in_83_port, reg_in_82_port, reg_in_81_port, reg_in_80_port, 
      reg_in_79_port, reg_in_78_port, reg_in_77_port, reg_in_76_port, 
      reg_in_75_port, reg_in_74_port, reg_in_73_port, reg_in_72_port, 
      reg_in_71_port, reg_in_70_port, reg_in_69_port, reg_in_68_port, 
      reg_in_67_port, reg_in_66_port, reg_in_65_port, reg_in_64_port, 
      reg_in_63_port, reg_in_62_port, reg_in_61_port, reg_in_60_port, 
      reg_in_59_port, reg_in_58_port, reg_in_57_port, reg_in_56_port, 
      reg_in_55_port, reg_in_54_port, reg_in_53_port, reg_in_52_port, 
      reg_in_51_port, reg_in_50_port, reg_in_49_port, reg_in_48_port, 
      reg_in_47_port, reg_in_46_port, reg_in_45_port, reg_in_44_port, 
      reg_in_43_port, reg_in_42_port, reg_in_41_port, reg_in_40_port, 
      reg_in_39_port, reg_in_38_port, reg_in_37_port, reg_in_36_port, 
      reg_in_35_port, reg_in_34_port, reg_in_33_port, reg_in_32_port, 
      reg_in_31_port, reg_in_30_port, reg_in_29_port, reg_in_28_port, 
      reg_in_27_port, reg_in_26_port, reg_in_25_port, reg_in_24_port, 
      reg_in_23_port, reg_in_22_port, reg_in_21_port, reg_in_20_port, 
      reg_in_19_port, reg_in_18_port, reg_in_17_port, reg_in_16_port, 
      reg_in_15_port, reg_in_14_port, reg_in_13_port, reg_in_12_port, 
      reg_in_11_port, reg_in_10_port, reg_in_9_port, reg_in_8_port, 
      reg_in_7_port, reg_in_6_port, reg_in_5_port, reg_in_4_port, reg_in_3_port
      , reg_in_2_port, reg_in_1_port, reg_in_0_port, reg_key_191_port, 
      reg_key_190_port, reg_key_189_port, reg_key_188_port, reg_key_187_port, 
      reg_key_185_port, reg_key_184_port, reg_key_183_port, reg_key_182_port, 
      reg_key_181_port, reg_key_180_port, reg_key_179_port, reg_key_178_port, 
      reg_key_177_port, reg_key_176_port, reg_key_175_port, reg_key_174_port, 
      reg_key_173_port, reg_key_172_port, reg_key_171_port, reg_key_170_port, 
      reg_key_169_port, reg_key_168_port, reg_key_167_port, reg_key_166_port, 
      reg_key_165_port, reg_key_164_port, reg_key_163_port, reg_key_162_port, 
      reg_key_161_port, reg_key_160_port, reg_key_159_port, reg_key_158_port, 
      reg_key_157_port, reg_key_156_port, reg_key_155_port, reg_key_154_port, 
      reg_key_153_port, reg_key_152_port, reg_key_151_port, reg_key_150_port, 
      reg_key_149_port, reg_key_148_port, reg_key_147_port, reg_key_146_port, 
      reg_key_145_port, reg_key_144_port, reg_key_143_port, reg_key_142_port, 
      reg_key_141_port, reg_key_140_port, reg_key_139_port, reg_key_138_port, 
      reg_key_137_port, reg_key_136_port, reg_key_135_port, reg_key_134_port, 
      reg_key_133_port, reg_key_132_port, reg_key_131_port, reg_key_130_port, 
      reg_key_129_port, reg_key_128_port, reg_key_127_port, reg_key_126_port, 
      reg_key_125_port, reg_key_124_port, reg_key_123_port, reg_key_122_port, 
      reg_key_121_port, reg_key_120_port, reg_key_119_port, reg_key_118_port, 
      reg_key_117_port, reg_key_116_port, reg_key_115_port, reg_key_114_port, 
      reg_key_113_port, reg_key_112_port, reg_key_111_port, reg_key_110_port, 
      reg_key_109_port, reg_key_108_port, reg_key_107_port, reg_key_106_port, 
      reg_key_105_port, reg_key_104_port, reg_key_103_port, reg_key_102_port, 
      reg_key_101_port, reg_key_100_port, reg_key_99_port, reg_key_98_port, 
      reg_key_97_port, reg_key_96_port, reg_key_95_port, reg_key_94_port, 
      reg_key_93_port, reg_key_92_port, reg_key_91_port, reg_key_90_port, 
      reg_key_89_port, reg_key_88_port, reg_key_87_port, reg_key_86_port, 
      reg_key_85_port, reg_key_84_port, reg_key_83_port, reg_key_82_port, 
      reg_key_81_port, reg_key_80_port, reg_key_79_port, reg_key_78_port, 
      reg_key_77_port, reg_key_76_port, reg_key_75_port, reg_key_74_port, 
      reg_key_73_port, reg_key_72_port, reg_key_71_port, reg_key_70_port, 
      reg_key_69_port, reg_key_68_port, reg_key_67_port, reg_key_66_port, 
      reg_key_65_port, reg_key_64_port, reg_key_63_port, reg_key_62_port, 
      reg_key_61_port, reg_key_60_port, reg_key_59_port, reg_key_58_port, 
      reg_key_57_port, reg_key_56_port, reg_key_55_port, reg_key_54_port, 
      reg_key_53_port, reg_key_52_port, reg_key_51_port, reg_key_50_port, 
      reg_key_49_port, reg_key_48_port, reg_key_47_port, reg_key_46_port, 
      reg_key_45_port, reg_key_44_port, reg_key_43_port, reg_key_42_port, 
      reg_key_41_port, reg_key_40_port, reg_key_39_port, reg_key_38_port, 
      reg_key_37_port, reg_key_36_port, reg_key_35_port, reg_key_34_port, 
      reg_key_33_port, reg_key_32_port, reg_key_31_port, reg_key_30_port, 
      reg_key_29_port, reg_key_28_port, reg_key_27_port, reg_key_26_port, 
      reg_key_25_port, reg_key_24_port, reg_key_23_port, reg_key_22_port, 
      reg_key_21_port, reg_key_20_port, reg_key_19_port, reg_key_18_port, 
      reg_key_17_port, reg_key_16_port, reg_key_15_port, reg_key_14_port, 
      reg_key_13_port, reg_key_12_port, reg_key_11_port, reg_key_10_port, 
      reg_key_9_port, reg_key_8_port, reg_key_7_port, reg_key_6_port, 
      reg_key_5_port, reg_key_4_port, reg_key_3_port, reg_key_2_port, 
      reg_key_1_port, reg_key_0_port, reg_out_191_port, reg_out_190_port, 
      reg_out_189_port, reg_out_188_port, reg_out_187_port, reg_out_186_port, 
      reg_out_185_port, reg_out_184_port, reg_out_183_port, reg_out_182_port, 
      reg_out_181_port, reg_out_180_port, reg_out_179_port, reg_out_178_port, 
      reg_out_177_port, reg_out_176_port, reg_out_175_port, reg_out_174_port, 
      reg_out_173_port, reg_out_172_port, reg_out_171_port, reg_out_170_port, 
      reg_out_169_port, reg_out_168_port, reg_out_167_port, reg_out_166_port, 
      reg_out_165_port, reg_out_164_port, reg_out_163_port, reg_out_162_port, 
      reg_out_161_port, reg_out_160_port, reg_out_159_port, reg_out_158_port, 
      reg_out_157_port, reg_out_156_port, reg_out_155_port, reg_out_154_port, 
      reg_out_153_port, reg_out_152_port, reg_out_151_port, reg_out_150_port, 
      reg_out_149_port, reg_out_148_port, reg_out_147_port, reg_out_146_port, 
      reg_out_145_port, reg_out_144_port, reg_out_143_port, reg_out_142_port, 
      reg_out_141_port, reg_out_140_port, reg_out_139_port, reg_out_138_port, 
      reg_out_137_port, reg_out_136_port, reg_out_135_port, reg_out_134_port, 
      reg_out_133_port, reg_out_132_port, reg_out_131_port, reg_out_130_port, 
      reg_out_129_port, reg_out_128_port, reg_out_127_port, reg_out_126_port, 
      reg_out_125_port, reg_out_124_port, reg_out_123_port, reg_out_122_port, 
      reg_out_121_port, reg_out_120_port, reg_out_119_port, reg_out_118_port, 
      reg_out_117_port, reg_out_116_port, reg_out_115_port, reg_out_114_port, 
      reg_out_113_port, reg_out_112_port, reg_out_111_port, reg_out_110_port, 
      reg_out_109_port, reg_out_108_port, reg_out_107_port, reg_out_106_port, 
      reg_out_105_port, reg_out_104_port, reg_out_103_port, reg_out_102_port, 
      reg_out_101_port, reg_out_100_port, reg_out_99_port, reg_out_98_port, 
      reg_out_97_port, reg_out_96_port, reg_out_95_port, reg_out_94_port, 
      reg_out_93_port, reg_out_92_port, reg_out_91_port, reg_out_90_port, 
      reg_out_89_port, reg_out_88_port, reg_out_87_port, reg_out_86_port, 
      reg_out_85_port, reg_out_84_port, reg_out_83_port, reg_out_82_port, 
      reg_out_81_port, reg_out_80_port, reg_out_79_port, reg_out_78_port, 
      reg_out_77_port, reg_out_76_port, reg_out_75_port, reg_out_74_port, 
      reg_out_73_port, reg_out_72_port, reg_out_71_port, reg_out_70_port, 
      reg_out_69_port, reg_out_68_port, reg_out_67_port, reg_out_66_port, 
      reg_out_65_port, reg_out_64_port, reg_out_63_port, reg_out_62_port, 
      reg_out_61_port, reg_out_60_port, reg_out_59_port, reg_out_58_port, 
      reg_out_57_port, reg_out_56_port, reg_out_55_port, reg_out_54_port, 
      reg_out_53_port, reg_out_52_port, reg_out_51_port, reg_out_50_port, 
      reg_out_49_port, reg_out_48_port, reg_out_47_port, reg_out_46_port, 
      reg_out_45_port, reg_out_44_port, reg_out_43_port, reg_out_42_port, 
      reg_out_41_port, reg_out_40_port, reg_out_39_port, reg_out_38_port, 
      reg_out_37_port, reg_out_36_port, reg_out_35_port, reg_out_34_port, 
      reg_out_33_port, reg_out_32_port, reg_out_31_port, reg_out_30_port, 
      reg_out_29_port, reg_out_28_port, reg_out_27_port, reg_out_26_port, 
      reg_out_25_port, reg_out_24_port, reg_out_23_port, reg_out_22_port, 
      reg_out_21_port, reg_out_20_port, reg_out_19_port, reg_out_18_port, 
      reg_out_17_port, reg_out_16_port, reg_out_15_port, reg_out_14_port, 
      reg_out_13_port, reg_out_12_port, reg_out_11_port, reg_out_10_port, 
      reg_out_9_port, reg_out_8_port, reg_out_7_port, reg_out_6_port, 
      reg_out_5_port, reg_out_4_port, reg_out_3_port, reg_out_2_port, 
      reg_out_1_port, reg_out_0_port, n3, n5, n9, n10, n11, n12, n_1000, n_1001
      , n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010,
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575 : std_logic;

begin
   
   reg_in_regx191x : DFF_X1 port map( D => Plaintext(191), CK => clk, Q => 
                           reg_in_191_port, QN => n_1000);
   reg_in_regx190x : DFF_X1 port map( D => Plaintext(190), CK => clk, Q => 
                           reg_in_190_port, QN => n_1001);
   reg_in_regx189x : DFF_X1 port map( D => Plaintext(189), CK => clk, Q => 
                           reg_in_189_port, QN => n_1002);
   reg_in_regx188x : DFF_X1 port map( D => Plaintext(188), CK => clk, Q => 
                           reg_in_188_port, QN => n_1003);
   reg_in_regx187x : DFF_X1 port map( D => Plaintext(187), CK => clk, Q => 
                           reg_in_187_port, QN => n_1004);
   reg_in_regx186x : DFF_X1 port map( D => Plaintext(186), CK => clk, Q => 
                           reg_in_186_port, QN => n_1005);
   reg_in_regx185x : DFF_X1 port map( D => Plaintext(185), CK => clk, Q => 
                           reg_in_185_port, QN => n_1006);
   reg_in_regx184x : DFF_X1 port map( D => Plaintext(184), CK => clk, Q => 
                           reg_in_184_port, QN => n_1007);
   reg_in_regx183x : DFF_X1 port map( D => Plaintext(183), CK => clk, Q => 
                           reg_in_183_port, QN => n_1008);
   reg_in_regx182x : DFF_X1 port map( D => Plaintext(182), CK => clk, Q => 
                           reg_in_182_port, QN => n_1009);
   reg_in_regx181x : DFF_X1 port map( D => Plaintext(181), CK => clk, Q => 
                           reg_in_181_port, QN => n_1010);
   reg_in_regx180x : DFF_X1 port map( D => Plaintext(180), CK => clk, Q => 
                           reg_in_180_port, QN => n_1011);
   reg_in_regx179x : DFF_X1 port map( D => Plaintext(179), CK => clk, Q => 
                           reg_in_179_port, QN => n_1012);
   reg_in_regx178x : DFF_X1 port map( D => Plaintext(178), CK => clk, Q => 
                           reg_in_178_port, QN => n_1013);
   reg_in_regx177x : DFF_X1 port map( D => Plaintext(177), CK => clk, Q => 
                           reg_in_177_port, QN => n_1014);
   reg_in_regx176x : DFF_X1 port map( D => Plaintext(176), CK => clk, Q => 
                           reg_in_176_port, QN => n_1015);
   reg_in_regx175x : DFF_X1 port map( D => Plaintext(175), CK => clk, Q => 
                           reg_in_175_port, QN => n_1016);
   reg_in_regx174x : DFF_X1 port map( D => Plaintext(174), CK => clk, Q => 
                           reg_in_174_port, QN => n_1017);
   reg_in_regx173x : DFF_X1 port map( D => Plaintext(173), CK => clk, Q => 
                           reg_in_173_port, QN => n_1018);
   reg_in_regx172x : DFF_X1 port map( D => Plaintext(172), CK => clk, Q => 
                           reg_in_172_port, QN => n_1019);
   reg_in_regx171x : DFF_X1 port map( D => Plaintext(171), CK => clk, Q => 
                           reg_in_171_port, QN => n_1020);
   reg_in_regx170x : DFF_X1 port map( D => Plaintext(170), CK => clk, Q => 
                           reg_in_170_port, QN => n_1021);
   reg_in_regx169x : DFF_X1 port map( D => Plaintext(169), CK => clk, Q => 
                           reg_in_169_port, QN => n_1022);
   reg_in_regx168x : DFF_X1 port map( D => Plaintext(168), CK => clk, Q => 
                           reg_in_168_port, QN => n_1023);
   reg_in_regx167x : DFF_X1 port map( D => Plaintext(167), CK => clk, Q => 
                           reg_in_167_port, QN => n_1024);
   reg_in_regx166x : DFF_X1 port map( D => Plaintext(166), CK => clk, Q => 
                           reg_in_166_port, QN => n_1025);
   reg_in_regx165x : DFF_X1 port map( D => Plaintext(165), CK => clk, Q => 
                           reg_in_165_port, QN => n_1026);
   reg_in_regx164x : DFF_X1 port map( D => Plaintext(164), CK => clk, Q => 
                           reg_in_164_port, QN => n_1027);
   reg_in_regx163x : DFF_X1 port map( D => Plaintext(163), CK => clk, Q => 
                           reg_in_163_port, QN => n_1028);
   reg_in_regx162x : DFF_X1 port map( D => Plaintext(162), CK => clk, Q => 
                           reg_in_162_port, QN => n_1029);
   reg_in_regx161x : DFF_X1 port map( D => Plaintext(161), CK => clk, Q => 
                           reg_in_161_port, QN => n_1030);
   reg_in_regx160x : DFF_X1 port map( D => Plaintext(160), CK => clk, Q => 
                           reg_in_160_port, QN => n_1031);
   reg_in_regx159x : DFF_X1 port map( D => Plaintext(159), CK => clk, Q => 
                           reg_in_159_port, QN => n_1032);
   reg_in_regx158x : DFF_X1 port map( D => Plaintext(158), CK => clk, Q => 
                           reg_in_158_port, QN => n_1033);
   reg_in_regx157x : DFF_X1 port map( D => Plaintext(157), CK => clk, Q => 
                           reg_in_157_port, QN => n_1034);
   reg_in_regx156x : DFF_X1 port map( D => Plaintext(156), CK => clk, Q => 
                           reg_in_156_port, QN => n_1035);
   reg_in_regx155x : DFF_X1 port map( D => Plaintext(155), CK => clk, Q => 
                           reg_in_155_port, QN => n_1036);
   reg_in_regx154x : DFF_X1 port map( D => Plaintext(154), CK => clk, Q => 
                           reg_in_154_port, QN => n_1037);
   reg_in_regx153x : DFF_X1 port map( D => Plaintext(153), CK => clk, Q => 
                           reg_in_153_port, QN => n_1038);
   reg_in_regx152x : DFF_X1 port map( D => Plaintext(152), CK => clk, Q => 
                           reg_in_152_port, QN => n_1039);
   reg_in_regx151x : DFF_X1 port map( D => Plaintext(151), CK => clk, Q => 
                           reg_in_151_port, QN => n_1040);
   reg_in_regx150x : DFF_X1 port map( D => Plaintext(150), CK => clk, Q => 
                           reg_in_150_port, QN => n_1041);
   reg_in_regx149x : DFF_X1 port map( D => Plaintext(149), CK => clk, Q => 
                           reg_in_149_port, QN => n_1042);
   reg_in_regx148x : DFF_X1 port map( D => Plaintext(148), CK => clk, Q => 
                           reg_in_148_port, QN => n_1043);
   reg_in_regx147x : DFF_X1 port map( D => Plaintext(147), CK => clk, Q => 
                           reg_in_147_port, QN => n_1044);
   reg_in_regx146x : DFF_X1 port map( D => Plaintext(146), CK => clk, Q => 
                           reg_in_146_port, QN => n_1045);
   reg_in_regx145x : DFF_X1 port map( D => Plaintext(145), CK => clk, Q => 
                           reg_in_145_port, QN => n_1046);
   reg_in_regx144x : DFF_X1 port map( D => Plaintext(144), CK => clk, Q => 
                           reg_in_144_port, QN => n_1047);
   reg_in_regx143x : DFF_X1 port map( D => Plaintext(143), CK => clk, Q => 
                           reg_in_143_port, QN => n_1048);
   reg_in_regx142x : DFF_X1 port map( D => Plaintext(142), CK => clk, Q => 
                           reg_in_142_port, QN => n_1049);
   reg_in_regx141x : DFF_X1 port map( D => Plaintext(141), CK => clk, Q => 
                           reg_in_141_port, QN => n_1050);
   reg_in_regx140x : DFF_X1 port map( D => Plaintext(140), CK => clk, Q => 
                           reg_in_140_port, QN => n_1051);
   reg_in_regx139x : DFF_X1 port map( D => Plaintext(139), CK => clk, Q => 
                           reg_in_139_port, QN => n_1052);
   reg_in_regx138x : DFF_X1 port map( D => Plaintext(138), CK => clk, Q => 
                           reg_in_138_port, QN => n_1053);
   reg_in_regx137x : DFF_X1 port map( D => Plaintext(137), CK => clk, Q => 
                           reg_in_137_port, QN => n_1054);
   reg_in_regx136x : DFF_X1 port map( D => Plaintext(136), CK => clk, Q => 
                           reg_in_136_port, QN => n_1055);
   reg_in_regx135x : DFF_X1 port map( D => Plaintext(135), CK => clk, Q => 
                           reg_in_135_port, QN => n_1056);
   reg_in_regx134x : DFF_X1 port map( D => Plaintext(134), CK => clk, Q => 
                           reg_in_134_port, QN => n_1057);
   reg_in_regx133x : DFF_X1 port map( D => Plaintext(133), CK => clk, Q => 
                           reg_in_133_port, QN => n_1058);
   reg_in_regx132x : DFF_X1 port map( D => Plaintext(132), CK => clk, Q => 
                           reg_in_132_port, QN => n_1059);
   reg_in_regx131x : DFF_X1 port map( D => Plaintext(131), CK => clk, Q => 
                           reg_in_131_port, QN => n_1060);
   reg_in_regx130x : DFF_X1 port map( D => Plaintext(130), CK => clk, Q => 
                           reg_in_130_port, QN => n_1061);
   reg_in_regx129x : DFF_X1 port map( D => Plaintext(129), CK => clk, Q => 
                           reg_in_129_port, QN => n_1062);
   reg_in_regx128x : DFF_X1 port map( D => Plaintext(128), CK => clk, Q => 
                           reg_in_128_port, QN => n_1063);
   reg_in_regx127x : DFF_X1 port map( D => Plaintext(127), CK => clk, Q => 
                           reg_in_127_port, QN => n_1064);
   reg_in_regx126x : DFF_X1 port map( D => Plaintext(126), CK => clk, Q => 
                           reg_in_126_port, QN => n_1065);
   reg_in_regx125x : DFF_X1 port map( D => Plaintext(125), CK => clk, Q => 
                           reg_in_125_port, QN => n_1066);
   reg_in_regx124x : DFF_X1 port map( D => Plaintext(124), CK => clk, Q => 
                           reg_in_124_port, QN => n_1067);
   reg_in_regx123x : DFF_X1 port map( D => Plaintext(123), CK => clk, Q => 
                           reg_in_123_port, QN => n_1068);
   reg_in_regx122x : DFF_X1 port map( D => Plaintext(122), CK => clk, Q => 
                           reg_in_122_port, QN => n_1069);
   reg_in_regx121x : DFF_X1 port map( D => Plaintext(121), CK => clk, Q => 
                           reg_in_121_port, QN => n_1070);
   reg_in_regx120x : DFF_X1 port map( D => Plaintext(120), CK => clk, Q => 
                           reg_in_120_port, QN => n_1071);
   reg_in_regx119x : DFF_X1 port map( D => Plaintext(119), CK => clk, Q => 
                           reg_in_119_port, QN => n_1072);
   reg_in_regx118x : DFF_X1 port map( D => Plaintext(118), CK => clk, Q => 
                           reg_in_118_port, QN => n_1073);
   reg_in_regx117x : DFF_X1 port map( D => Plaintext(117), CK => clk, Q => 
                           reg_in_117_port, QN => n_1074);
   reg_in_regx116x : DFF_X1 port map( D => Plaintext(116), CK => clk, Q => 
                           reg_in_116_port, QN => n_1075);
   reg_in_regx115x : DFF_X1 port map( D => Plaintext(115), CK => clk, Q => 
                           reg_in_115_port, QN => n_1076);
   reg_in_regx114x : DFF_X1 port map( D => Plaintext(114), CK => clk, Q => 
                           reg_in_114_port, QN => n_1077);
   reg_in_regx113x : DFF_X1 port map( D => Plaintext(113), CK => clk, Q => 
                           reg_in_113_port, QN => n_1078);
   reg_in_regx112x : DFF_X1 port map( D => Plaintext(112), CK => clk, Q => 
                           reg_in_112_port, QN => n_1079);
   reg_in_regx111x : DFF_X1 port map( D => Plaintext(111), CK => clk, Q => 
                           reg_in_111_port, QN => n_1080);
   reg_in_regx110x : DFF_X1 port map( D => Plaintext(110), CK => clk, Q => 
                           reg_in_110_port, QN => n_1081);
   reg_in_regx109x : DFF_X1 port map( D => Plaintext(109), CK => clk, Q => 
                           reg_in_109_port, QN => n_1082);
   reg_in_regx108x : DFF_X1 port map( D => Plaintext(108), CK => clk, Q => 
                           reg_in_108_port, QN => n_1083);
   reg_in_regx107x : DFF_X1 port map( D => Plaintext(107), CK => clk, Q => 
                           reg_in_107_port, QN => n_1084);
   reg_in_regx106x : DFF_X1 port map( D => Plaintext(106), CK => clk, Q => 
                           reg_in_106_port, QN => n_1085);
   reg_in_regx105x : DFF_X1 port map( D => Plaintext(105), CK => clk, Q => 
                           reg_in_105_port, QN => n_1086);
   reg_in_regx104x : DFF_X1 port map( D => Plaintext(104), CK => clk, Q => 
                           reg_in_104_port, QN => n_1087);
   reg_in_regx103x : DFF_X1 port map( D => Plaintext(103), CK => clk, Q => 
                           reg_in_103_port, QN => n_1088);
   reg_in_regx102x : DFF_X1 port map( D => Plaintext(102), CK => clk, Q => 
                           reg_in_102_port, QN => n_1089);
   reg_in_regx101x : DFF_X1 port map( D => Plaintext(101), CK => clk, Q => 
                           reg_in_101_port, QN => n_1090);
   reg_in_regx100x : DFF_X1 port map( D => Plaintext(100), CK => clk, Q => 
                           reg_in_100_port, QN => n_1091);
   reg_in_regx99x : DFF_X1 port map( D => Plaintext(99), CK => clk, Q => 
                           reg_in_99_port, QN => n_1092);
   reg_in_regx98x : DFF_X1 port map( D => Plaintext(98), CK => clk, Q => 
                           reg_in_98_port, QN => n_1093);
   reg_in_regx97x : DFF_X1 port map( D => Plaintext(97), CK => clk, Q => 
                           reg_in_97_port, QN => n_1094);
   reg_in_regx96x : DFF_X1 port map( D => Plaintext(96), CK => clk, Q => 
                           reg_in_96_port, QN => n_1095);
   reg_in_regx95x : DFF_X1 port map( D => Plaintext(95), CK => clk, Q => 
                           reg_in_95_port, QN => n_1096);
   reg_in_regx94x : DFF_X1 port map( D => Plaintext(94), CK => clk, Q => 
                           reg_in_94_port, QN => n_1097);
   reg_in_regx93x : DFF_X1 port map( D => Plaintext(93), CK => clk, Q => 
                           reg_in_93_port, QN => n_1098);
   reg_in_regx92x : DFF_X1 port map( D => Plaintext(92), CK => clk, Q => 
                           reg_in_92_port, QN => n_1099);
   reg_in_regx91x : DFF_X1 port map( D => Plaintext(91), CK => clk, Q => 
                           reg_in_91_port, QN => n_1100);
   reg_in_regx90x : DFF_X1 port map( D => Plaintext(90), CK => clk, Q => 
                           reg_in_90_port, QN => n_1101);
   reg_in_regx89x : DFF_X1 port map( D => Plaintext(89), CK => clk, Q => 
                           reg_in_89_port, QN => n_1102);
   reg_in_regx88x : DFF_X1 port map( D => Plaintext(88), CK => clk, Q => 
                           reg_in_88_port, QN => n_1103);
   reg_in_regx87x : DFF_X1 port map( D => Plaintext(87), CK => clk, Q => 
                           reg_in_87_port, QN => n_1104);
   reg_in_regx86x : DFF_X1 port map( D => Plaintext(86), CK => clk, Q => 
                           reg_in_86_port, QN => n_1105);
   reg_in_regx85x : DFF_X1 port map( D => Plaintext(85), CK => clk, Q => 
                           reg_in_85_port, QN => n_1106);
   reg_in_regx84x : DFF_X1 port map( D => Plaintext(84), CK => clk, Q => 
                           reg_in_84_port, QN => n_1107);
   reg_in_regx83x : DFF_X1 port map( D => Plaintext(83), CK => clk, Q => 
                           reg_in_83_port, QN => n_1108);
   reg_in_regx82x : DFF_X1 port map( D => Plaintext(82), CK => clk, Q => 
                           reg_in_82_port, QN => n_1109);
   reg_in_regx81x : DFF_X1 port map( D => Plaintext(81), CK => clk, Q => 
                           reg_in_81_port, QN => n_1110);
   reg_in_regx80x : DFF_X1 port map( D => Plaintext(80), CK => clk, Q => 
                           reg_in_80_port, QN => n_1111);
   reg_in_regx79x : DFF_X1 port map( D => Plaintext(79), CK => clk, Q => 
                           reg_in_79_port, QN => n_1112);
   reg_in_regx78x : DFF_X1 port map( D => Plaintext(78), CK => clk, Q => 
                           reg_in_78_port, QN => n_1113);
   reg_in_regx77x : DFF_X1 port map( D => Plaintext(77), CK => clk, Q => 
                           reg_in_77_port, QN => n_1114);
   reg_in_regx76x : DFF_X1 port map( D => Plaintext(76), CK => clk, Q => 
                           reg_in_76_port, QN => n_1115);
   reg_in_regx75x : DFF_X1 port map( D => Plaintext(75), CK => clk, Q => 
                           reg_in_75_port, QN => n_1116);
   reg_in_regx74x : DFF_X1 port map( D => Plaintext(74), CK => clk, Q => 
                           reg_in_74_port, QN => n_1117);
   reg_in_regx73x : DFF_X1 port map( D => Plaintext(73), CK => clk, Q => 
                           reg_in_73_port, QN => n_1118);
   reg_in_regx72x : DFF_X1 port map( D => Plaintext(72), CK => clk, Q => 
                           reg_in_72_port, QN => n_1119);
   reg_in_regx71x : DFF_X1 port map( D => Plaintext(71), CK => clk, Q => 
                           reg_in_71_port, QN => n_1120);
   reg_in_regx70x : DFF_X1 port map( D => Plaintext(70), CK => clk, Q => 
                           reg_in_70_port, QN => n_1121);
   reg_in_regx69x : DFF_X1 port map( D => Plaintext(69), CK => clk, Q => 
                           reg_in_69_port, QN => n_1122);
   reg_in_regx68x : DFF_X1 port map( D => Plaintext(68), CK => clk, Q => 
                           reg_in_68_port, QN => n_1123);
   reg_in_regx67x : DFF_X1 port map( D => Plaintext(67), CK => clk, Q => 
                           reg_in_67_port, QN => n_1124);
   reg_in_regx66x : DFF_X1 port map( D => Plaintext(66), CK => clk, Q => 
                           reg_in_66_port, QN => n_1125);
   reg_in_regx65x : DFF_X1 port map( D => Plaintext(65), CK => clk, Q => 
                           reg_in_65_port, QN => n_1126);
   reg_in_regx64x : DFF_X1 port map( D => Plaintext(64), CK => clk, Q => 
                           reg_in_64_port, QN => n_1127);
   reg_in_regx63x : DFF_X1 port map( D => Plaintext(63), CK => clk, Q => 
                           reg_in_63_port, QN => n_1128);
   reg_in_regx62x : DFF_X1 port map( D => Plaintext(62), CK => clk, Q => 
                           reg_in_62_port, QN => n_1129);
   reg_in_regx61x : DFF_X1 port map( D => Plaintext(61), CK => clk, Q => 
                           reg_in_61_port, QN => n_1130);
   reg_in_regx60x : DFF_X1 port map( D => Plaintext(60), CK => clk, Q => 
                           reg_in_60_port, QN => n_1131);
   reg_in_regx59x : DFF_X1 port map( D => Plaintext(59), CK => clk, Q => 
                           reg_in_59_port, QN => n_1132);
   reg_in_regx58x : DFF_X1 port map( D => Plaintext(58), CK => clk, Q => 
                           reg_in_58_port, QN => n_1133);
   reg_in_regx57x : DFF_X1 port map( D => Plaintext(57), CK => clk, Q => 
                           reg_in_57_port, QN => n_1134);
   reg_in_regx56x : DFF_X1 port map( D => Plaintext(56), CK => clk, Q => 
                           reg_in_56_port, QN => n_1135);
   reg_in_regx55x : DFF_X1 port map( D => Plaintext(55), CK => clk, Q => 
                           reg_in_55_port, QN => n_1136);
   reg_in_regx54x : DFF_X1 port map( D => Plaintext(54), CK => clk, Q => 
                           reg_in_54_port, QN => n_1137);
   reg_in_regx53x : DFF_X1 port map( D => Plaintext(53), CK => clk, Q => 
                           reg_in_53_port, QN => n_1138);
   reg_in_regx52x : DFF_X1 port map( D => Plaintext(52), CK => clk, Q => 
                           reg_in_52_port, QN => n_1139);
   reg_in_regx51x : DFF_X1 port map( D => Plaintext(51), CK => clk, Q => 
                           reg_in_51_port, QN => n_1140);
   reg_in_regx50x : DFF_X1 port map( D => Plaintext(50), CK => clk, Q => 
                           reg_in_50_port, QN => n_1141);
   reg_in_regx49x : DFF_X1 port map( D => Plaintext(49), CK => clk, Q => 
                           reg_in_49_port, QN => n_1142);
   reg_in_regx48x : DFF_X1 port map( D => Plaintext(48), CK => clk, Q => 
                           reg_in_48_port, QN => n_1143);
   reg_in_regx47x : DFF_X1 port map( D => Plaintext(47), CK => clk, Q => 
                           reg_in_47_port, QN => n_1144);
   reg_in_regx46x : DFF_X1 port map( D => Plaintext(46), CK => clk, Q => 
                           reg_in_46_port, QN => n_1145);
   reg_in_regx45x : DFF_X1 port map( D => Plaintext(45), CK => clk, Q => 
                           reg_in_45_port, QN => n_1146);
   reg_in_regx44x : DFF_X1 port map( D => Plaintext(44), CK => clk, Q => 
                           reg_in_44_port, QN => n_1147);
   reg_in_regx43x : DFF_X1 port map( D => Plaintext(43), CK => clk, Q => 
                           reg_in_43_port, QN => n_1148);
   reg_in_regx42x : DFF_X1 port map( D => Plaintext(42), CK => clk, Q => 
                           reg_in_42_port, QN => n_1149);
   reg_in_regx41x : DFF_X1 port map( D => Plaintext(41), CK => clk, Q => 
                           reg_in_41_port, QN => n_1150);
   reg_in_regx40x : DFF_X1 port map( D => Plaintext(40), CK => clk, Q => 
                           reg_in_40_port, QN => n_1151);
   reg_in_regx39x : DFF_X1 port map( D => Plaintext(39), CK => clk, Q => 
                           reg_in_39_port, QN => n_1152);
   reg_in_regx38x : DFF_X1 port map( D => Plaintext(38), CK => clk, Q => 
                           reg_in_38_port, QN => n_1153);
   reg_in_regx37x : DFF_X1 port map( D => Plaintext(37), CK => clk, Q => 
                           reg_in_37_port, QN => n_1154);
   reg_in_regx36x : DFF_X1 port map( D => Plaintext(36), CK => clk, Q => 
                           reg_in_36_port, QN => n_1155);
   reg_in_regx35x : DFF_X1 port map( D => Plaintext(35), CK => clk, Q => 
                           reg_in_35_port, QN => n_1156);
   reg_in_regx34x : DFF_X1 port map( D => Plaintext(34), CK => clk, Q => 
                           reg_in_34_port, QN => n_1157);
   reg_in_regx33x : DFF_X1 port map( D => Plaintext(33), CK => clk, Q => 
                           reg_in_33_port, QN => n_1158);
   reg_in_regx32x : DFF_X1 port map( D => Plaintext(32), CK => clk, Q => 
                           reg_in_32_port, QN => n_1159);
   reg_in_regx31x : DFF_X1 port map( D => Plaintext(31), CK => clk, Q => 
                           reg_in_31_port, QN => n_1160);
   reg_in_regx30x : DFF_X1 port map( D => Plaintext(30), CK => clk, Q => 
                           reg_in_30_port, QN => n_1161);
   reg_in_regx29x : DFF_X1 port map( D => Plaintext(29), CK => clk, Q => 
                           reg_in_29_port, QN => n_1162);
   reg_in_regx28x : DFF_X1 port map( D => Plaintext(28), CK => clk, Q => 
                           reg_in_28_port, QN => n_1163);
   reg_in_regx27x : DFF_X1 port map( D => Plaintext(27), CK => clk, Q => 
                           reg_in_27_port, QN => n_1164);
   reg_in_regx26x : DFF_X1 port map( D => Plaintext(26), CK => clk, Q => 
                           reg_in_26_port, QN => n_1165);
   reg_in_regx25x : DFF_X1 port map( D => Plaintext(25), CK => clk, Q => 
                           reg_in_25_port, QN => n_1166);
   reg_in_regx24x : DFF_X1 port map( D => Plaintext(24), CK => clk, Q => 
                           reg_in_24_port, QN => n_1167);
   reg_in_regx23x : DFF_X1 port map( D => Plaintext(23), CK => clk, Q => 
                           reg_in_23_port, QN => n_1168);
   reg_in_regx22x : DFF_X1 port map( D => Plaintext(22), CK => clk, Q => 
                           reg_in_22_port, QN => n_1169);
   reg_in_regx21x : DFF_X1 port map( D => Plaintext(21), CK => clk, Q => 
                           reg_in_21_port, QN => n_1170);
   reg_in_regx20x : DFF_X1 port map( D => Plaintext(20), CK => clk, Q => 
                           reg_in_20_port, QN => n_1171);
   reg_in_regx19x : DFF_X1 port map( D => Plaintext(19), CK => clk, Q => 
                           reg_in_19_port, QN => n_1172);
   reg_in_regx18x : DFF_X1 port map( D => Plaintext(18), CK => clk, Q => 
                           reg_in_18_port, QN => n_1173);
   reg_in_regx17x : DFF_X1 port map( D => Plaintext(17), CK => clk, Q => 
                           reg_in_17_port, QN => n_1174);
   reg_in_regx16x : DFF_X1 port map( D => Plaintext(16), CK => clk, Q => 
                           reg_in_16_port, QN => n_1175);
   reg_in_regx15x : DFF_X1 port map( D => Plaintext(15), CK => clk, Q => 
                           reg_in_15_port, QN => n_1176);
   reg_in_regx14x : DFF_X1 port map( D => Plaintext(14), CK => clk, Q => 
                           reg_in_14_port, QN => n_1177);
   reg_in_regx13x : DFF_X1 port map( D => Plaintext(13), CK => clk, Q => 
                           reg_in_13_port, QN => n_1178);
   reg_in_regx12x : DFF_X1 port map( D => Plaintext(12), CK => clk, Q => 
                           reg_in_12_port, QN => n_1179);
   reg_in_regx11x : DFF_X1 port map( D => Plaintext(11), CK => clk, Q => 
                           reg_in_11_port, QN => n_1180);
   reg_in_regx10x : DFF_X1 port map( D => Plaintext(10), CK => clk, Q => 
                           reg_in_10_port, QN => n_1181);
   reg_in_regx9x : DFF_X1 port map( D => Plaintext(9), CK => clk, Q => 
                           reg_in_9_port, QN => n_1182);
   reg_in_regx8x : DFF_X1 port map( D => Plaintext(8), CK => clk, Q => 
                           reg_in_8_port, QN => n_1183);
   reg_in_regx7x : DFF_X1 port map( D => Plaintext(7), CK => clk, Q => 
                           reg_in_7_port, QN => n_1184);
   reg_in_regx6x : DFF_X1 port map( D => Plaintext(6), CK => clk, Q => 
                           reg_in_6_port, QN => n_1185);
   reg_in_regx5x : DFF_X1 port map( D => Plaintext(5), CK => clk, Q => 
                           reg_in_5_port, QN => n_1186);
   reg_in_regx4x : DFF_X1 port map( D => Plaintext(4), CK => clk, Q => 
                           reg_in_4_port, QN => n_1187);
   reg_in_regx3x : DFF_X1 port map( D => Plaintext(3), CK => clk, Q => 
                           reg_in_3_port, QN => n_1188);
   reg_in_regx2x : DFF_X1 port map( D => Plaintext(2), CK => clk, Q => 
                           reg_in_2_port, QN => n_1189);
   reg_in_regx1x : DFF_X1 port map( D => Plaintext(1), CK => clk, Q => 
                           reg_in_1_port, QN => n_1190);
   reg_in_regx0x : DFF_X1 port map( D => Plaintext(0), CK => clk, Q => 
                           reg_in_0_port, QN => n_1191);
   reg_key_regx191x : DFF_X1 port map( D => Key(191), CK => clk, Q => 
                           reg_key_191_port, QN => n_1192);
   reg_key_regx190x : DFF_X1 port map( D => Key(190), CK => clk, Q => 
                           reg_key_190_port, QN => n_1193);
   reg_key_regx189x : DFF_X1 port map( D => Key(189), CK => clk, Q => 
                           reg_key_189_port, QN => n_1194);
   reg_key_regx188x : DFF_X1 port map( D => Key(188), CK => clk, Q => 
                           reg_key_188_port, QN => n_1195);
   reg_key_regx186x : DFF_X1 port map( D => Key(186), CK => clk, Q => n3, QN =>
                           n_1196);
   reg_key_regx184x : DFF_X1 port map( D => Key(184), CK => clk, Q => 
                           reg_key_184_port, QN => n_1197);
   reg_key_regx181x : DFF_X1 port map( D => Key(181), CK => clk, Q => 
                           reg_key_181_port, QN => n_1198);
   reg_key_regx180x : DFF_X1 port map( D => Key(180), CK => clk, Q => 
                           reg_key_180_port, QN => n_1199);
   reg_key_regx178x : DFF_X1 port map( D => Key(178), CK => clk, Q => 
                           reg_key_178_port, QN => n_1200);
   reg_key_regx177x : DFF_X1 port map( D => Key(177), CK => clk, Q => 
                           reg_key_177_port, QN => n_1201);
   reg_key_regx176x : DFF_X1 port map( D => Key(176), CK => clk, Q => 
                           reg_key_176_port, QN => n_1202);
   reg_key_regx175x : DFF_X1 port map( D => Key(175), CK => clk, Q => 
                           reg_key_175_port, QN => n_1203);
   reg_key_regx174x : DFF_X1 port map( D => Key(174), CK => clk, Q => 
                           reg_key_174_port, QN => n_1204);
   reg_key_regx173x : DFF_X1 port map( D => Key(173), CK => clk, Q => 
                           reg_key_173_port, QN => n_1205);
   reg_key_regx172x : DFF_X1 port map( D => Key(172), CK => clk, Q => 
                           reg_key_172_port, QN => n_1206);
   reg_key_regx170x : DFF_X1 port map( D => Key(170), CK => clk, Q => 
                           reg_key_170_port, QN => n_1207);
   reg_key_regx169x : DFF_X1 port map( D => Key(169), CK => clk, Q => 
                           reg_key_169_port, QN => n_1208);
   reg_key_regx168x : DFF_X1 port map( D => Key(168), CK => clk, Q => 
                           reg_key_168_port, QN => n_1209);
   reg_key_regx167x : DFF_X1 port map( D => Key(167), CK => clk, Q => 
                           reg_key_167_port, QN => n_1210);
   reg_key_regx164x : DFF_X1 port map( D => Key(164), CK => clk, Q => 
                           reg_key_164_port, QN => n_1211);
   reg_key_regx163x : DFF_X1 port map( D => Key(163), CK => clk, Q => 
                           reg_key_163_port, QN => n_1212);
   reg_key_regx162x : DFF_X1 port map( D => Key(162), CK => clk, Q => 
                           reg_key_162_port, QN => n_1213);
   reg_key_regx161x : DFF_X1 port map( D => Key(161), CK => clk, Q => 
                           reg_key_161_port, QN => n_1214);
   reg_key_regx160x : DFF_X1 port map( D => Key(160), CK => clk, Q => 
                           reg_key_160_port, QN => n_1215);
   reg_key_regx159x : DFF_X1 port map( D => Key(159), CK => clk, Q => 
                           reg_key_159_port, QN => n_1216);
   reg_key_regx158x : DFF_X1 port map( D => Key(158), CK => clk, Q => 
                           reg_key_158_port, QN => n_1217);
   reg_key_regx157x : DFF_X1 port map( D => Key(157), CK => clk, Q => 
                           reg_key_157_port, QN => n_1218);
   reg_key_regx156x : DFF_X1 port map( D => Key(156), CK => clk, Q => 
                           reg_key_156_port, QN => n_1219);
   reg_key_regx155x : DFF_X1 port map( D => Key(155), CK => clk, Q => 
                           reg_key_155_port, QN => n_1220);
   reg_key_regx154x : DFF_X1 port map( D => Key(154), CK => clk, Q => 
                           reg_key_154_port, QN => n_1221);
   reg_key_regx153x : DFF_X1 port map( D => Key(153), CK => clk, Q => 
                           reg_key_153_port, QN => n_1222);
   reg_key_regx152x : DFF_X1 port map( D => Key(152), CK => clk, Q => 
                           reg_key_152_port, QN => n_1223);
   reg_key_regx151x : DFF_X1 port map( D => Key(151), CK => clk, Q => 
                           reg_key_151_port, QN => n_1224);
   reg_key_regx149x : DFF_X1 port map( D => Key(149), CK => clk, Q => 
                           reg_key_149_port, QN => n_1225);
   reg_key_regx148x : DFF_X1 port map( D => Key(148), CK => clk, Q => 
                           reg_key_148_port, QN => n_1226);
   reg_key_regx147x : DFF_X1 port map( D => Key(147), CK => clk, Q => 
                           reg_key_147_port, QN => n_1227);
   reg_key_regx146x : DFF_X1 port map( D => Key(146), CK => clk, Q => 
                           reg_key_146_port, QN => n_1228);
   reg_key_regx145x : DFF_X1 port map( D => Key(145), CK => clk, Q => 
                           reg_key_145_port, QN => n_1229);
   reg_key_regx144x : DFF_X1 port map( D => Key(144), CK => clk, Q => 
                           reg_key_144_port, QN => n_1230);
   reg_key_regx143x : DFF_X1 port map( D => Key(143), CK => clk, Q => 
                           reg_key_143_port, QN => n_1231);
   reg_key_regx142x : DFF_X1 port map( D => Key(142), CK => clk, Q => 
                           reg_key_142_port, QN => n_1232);
   reg_key_regx141x : DFF_X1 port map( D => Key(141), CK => clk, Q => 
                           reg_key_141_port, QN => n_1233);
   reg_key_regx140x : DFF_X1 port map( D => Key(140), CK => clk, Q => 
                           reg_key_140_port, QN => n_1234);
   reg_key_regx139x : DFF_X1 port map( D => Key(139), CK => clk, Q => 
                           reg_key_139_port, QN => n_1235);
   reg_key_regx138x : DFF_X1 port map( D => Key(138), CK => clk, Q => 
                           reg_key_138_port, QN => n_1236);
   reg_key_regx137x : DFF_X1 port map( D => Key(137), CK => clk, Q => 
                           reg_key_137_port, QN => n_1237);
   reg_key_regx136x : DFF_X1 port map( D => Key(136), CK => clk, Q => 
                           reg_key_136_port, QN => n_1238);
   reg_key_regx135x : DFF_X1 port map( D => Key(135), CK => clk, Q => 
                           reg_key_135_port, QN => n_1239);
   reg_key_regx133x : DFF_X1 port map( D => Key(133), CK => clk, Q => 
                           reg_key_133_port, QN => n_1240);
   reg_key_regx132x : DFF_X1 port map( D => Key(132), CK => clk, Q => 
                           reg_key_132_port, QN => n_1241);
   reg_key_regx131x : DFF_X1 port map( D => Key(131), CK => clk, Q => 
                           reg_key_131_port, QN => n_1242);
   reg_key_regx130x : DFF_X1 port map( D => Key(130), CK => clk, Q => 
                           reg_key_130_port, QN => n_1243);
   reg_key_regx129x : DFF_X1 port map( D => Key(129), CK => clk, Q => 
                           reg_key_129_port, QN => n_1244);
   reg_key_regx128x : DFF_X1 port map( D => Key(128), CK => clk, Q => 
                           reg_key_128_port, QN => n_1245);
   reg_key_regx127x : DFF_X1 port map( D => Key(127), CK => clk, Q => 
                           reg_key_127_port, QN => n_1246);
   reg_key_regx125x : DFF_X1 port map( D => Key(125), CK => clk, Q => 
                           reg_key_125_port, QN => n_1247);
   reg_key_regx124x : DFF_X1 port map( D => Key(124), CK => clk, Q => 
                           reg_key_124_port, QN => n_1248);
   reg_key_regx123x : DFF_X1 port map( D => Key(123), CK => clk, Q => 
                           reg_key_123_port, QN => n_1249);
   reg_key_regx122x : DFF_X1 port map( D => Key(122), CK => clk, Q => 
                           reg_key_122_port, QN => n_1250);
   reg_key_regx121x : DFF_X1 port map( D => Key(121), CK => clk, Q => 
                           reg_key_121_port, QN => n_1251);
   reg_key_regx120x : DFF_X1 port map( D => Key(120), CK => clk, Q => 
                           reg_key_120_port, QN => n_1252);
   reg_key_regx119x : DFF_X1 port map( D => Key(119), CK => clk, Q => 
                           reg_key_119_port, QN => n_1253);
   reg_key_regx118x : DFF_X1 port map( D => Key(118), CK => clk, Q => 
                           reg_key_118_port, QN => n_1254);
   reg_key_regx117x : DFF_X1 port map( D => Key(117), CK => clk, Q => 
                           reg_key_117_port, QN => n_1255);
   reg_key_regx116x : DFF_X1 port map( D => Key(116), CK => clk, Q => 
                           reg_key_116_port, QN => n_1256);
   reg_key_regx115x : DFF_X1 port map( D => Key(115), CK => clk, Q => 
                           reg_key_115_port, QN => n_1257);
   reg_key_regx114x : DFF_X1 port map( D => Key(114), CK => clk, Q => 
                           reg_key_114_port, QN => n_1258);
   reg_key_regx112x : DFF_X1 port map( D => Key(112), CK => clk, Q => 
                           reg_key_112_port, QN => n_1259);
   reg_key_regx111x : DFF_X1 port map( D => Key(111), CK => clk, Q => 
                           reg_key_111_port, QN => n_1260);
   reg_key_regx109x : DFF_X1 port map( D => Key(109), CK => clk, Q => 
                           reg_key_109_port, QN => n_1261);
   reg_key_regx108x : DFF_X1 port map( D => Key(108), CK => clk, Q => 
                           reg_key_108_port, QN => n_1262);
   reg_key_regx106x : DFF_X1 port map( D => Key(106), CK => clk, Q => 
                           reg_key_106_port, QN => n_1263);
   reg_key_regx104x : DFF_X1 port map( D => Key(104), CK => clk, Q => 
                           reg_key_104_port, QN => n_1264);
   reg_key_regx103x : DFF_X1 port map( D => Key(103), CK => clk, Q => 
                           reg_key_103_port, QN => n_1265);
   reg_key_regx102x : DFF_X1 port map( D => Key(102), CK => clk, Q => 
                           reg_key_102_port, QN => n_1266);
   reg_key_regx101x : DFF_X1 port map( D => Key(101), CK => clk, Q => 
                           reg_key_101_port, QN => n_1267);
   reg_key_regx100x : DFF_X1 port map( D => Key(100), CK => clk, Q => 
                           reg_key_100_port, QN => n_1268);
   reg_key_regx99x : DFF_X1 port map( D => Key(99), CK => clk, Q => 
                           reg_key_99_port, QN => n_1269);
   reg_key_regx98x : DFF_X1 port map( D => Key(98), CK => clk, Q => 
                           reg_key_98_port, QN => n_1270);
   reg_key_regx97x : DFF_X1 port map( D => Key(97), CK => clk, Q => 
                           reg_key_97_port, QN => n_1271);
   reg_key_regx96x : DFF_X1 port map( D => Key(96), CK => clk, Q => 
                           reg_key_96_port, QN => n_1272);
   reg_key_regx95x : DFF_X1 port map( D => Key(95), CK => clk, Q => 
                           reg_key_95_port, QN => n_1273);
   reg_key_regx94x : DFF_X1 port map( D => Key(94), CK => clk, Q => 
                           reg_key_94_port, QN => n_1274);
   reg_key_regx93x : DFF_X1 port map( D => Key(93), CK => clk, Q => 
                           reg_key_93_port, QN => n_1275);
   reg_key_regx92x : DFF_X1 port map( D => Key(92), CK => clk, Q => 
                           reg_key_92_port, QN => n_1276);
   reg_key_regx91x : DFF_X1 port map( D => Key(91), CK => clk, Q => 
                           reg_key_91_port, QN => n_1277);
   reg_key_regx90x : DFF_X1 port map( D => Key(90), CK => clk, Q => 
                           reg_key_90_port, QN => n_1278);
   reg_key_regx88x : DFF_X1 port map( D => Key(88), CK => clk, Q => 
                           reg_key_88_port, QN => n_1279);
   reg_key_regx85x : DFF_X1 port map( D => Key(85), CK => clk, Q => 
                           reg_key_85_port, QN => n_1280);
   reg_key_regx84x : DFF_X1 port map( D => Key(84), CK => clk, Q => 
                           reg_key_84_port, QN => n_1281);
   reg_key_regx82x : DFF_X1 port map( D => Key(82), CK => clk, Q => 
                           reg_key_82_port, QN => n_1282);
   reg_key_regx81x : DFF_X1 port map( D => Key(81), CK => clk, Q => 
                           reg_key_81_port, QN => n_1283);
   reg_key_regx80x : DFF_X1 port map( D => Key(80), CK => clk, Q => 
                           reg_key_80_port, QN => n_1284);
   reg_key_regx78x : DFF_X1 port map( D => Key(78), CK => clk, Q => 
                           reg_key_78_port, QN => n_1285);
   reg_key_regx76x : DFF_X1 port map( D => Key(76), CK => clk, Q => 
                           reg_key_76_port, QN => n_1286);
   reg_key_regx75x : DFF_X1 port map( D => Key(75), CK => clk, Q => 
                           reg_key_75_port, QN => n_1287);
   reg_key_regx74x : DFF_X1 port map( D => Key(74), CK => clk, Q => 
                           reg_key_74_port, QN => n_1288);
   reg_key_regx73x : DFF_X1 port map( D => Key(73), CK => clk, Q => 
                           reg_key_73_port, QN => n_1289);
   reg_key_regx72x : DFF_X1 port map( D => Key(72), CK => clk, Q => 
                           reg_key_72_port, QN => n_1290);
   reg_key_regx70x : DFF_X1 port map( D => Key(70), CK => clk, Q => 
                           reg_key_70_port, QN => n_1291);
   reg_key_regx69x : DFF_X1 port map( D => Key(69), CK => clk, Q => 
                           reg_key_69_port, QN => n_1292);
   reg_key_regx67x : DFF_X1 port map( D => Key(67), CK => clk, Q => 
                           reg_key_67_port, QN => n_1293);
   reg_key_regx66x : DFF_X1 port map( D => Key(66), CK => clk, Q => 
                           reg_key_66_port, QN => n_1294);
   reg_key_regx61x : DFF_X1 port map( D => Key(61), CK => clk, Q => 
                           reg_key_61_port, QN => n_1295);
   reg_key_regx59x : DFF_X1 port map( D => Key(59), CK => clk, Q => 
                           reg_key_59_port, QN => n_1296);
   reg_key_regx58x : DFF_X1 port map( D => Key(58), CK => clk, Q => 
                           reg_key_58_port, QN => n_1297);
   reg_key_regx57x : DFF_X1 port map( D => Key(57), CK => clk, Q => 
                           reg_key_57_port, QN => n_1298);
   reg_key_regx55x : DFF_X1 port map( D => Key(55), CK => clk, Q => 
                           reg_key_55_port, QN => n_1299);
   reg_key_regx54x : DFF_X1 port map( D => Key(54), CK => clk, Q => 
                           reg_key_54_port, QN => n_1300);
   reg_key_regx53x : DFF_X1 port map( D => Key(53), CK => clk, Q => 
                           reg_key_53_port, QN => n_1301);
   reg_key_regx51x : DFF_X1 port map( D => Key(51), CK => clk, Q => 
                           reg_key_51_port, QN => n_1302);
   reg_key_regx50x : DFF_X1 port map( D => Key(50), CK => clk, Q => 
                           reg_key_50_port, QN => n_1303);
   reg_key_regx49x : DFF_X1 port map( D => Key(49), CK => clk, Q => 
                           reg_key_49_port, QN => n_1304);
   reg_key_regx48x : DFF_X1 port map( D => Key(48), CK => clk, Q => 
                           reg_key_48_port, QN => n_1305);
   reg_key_regx47x : DFF_X1 port map( D => Key(47), CK => clk, Q => 
                           reg_key_47_port, QN => n_1306);
   reg_key_regx45x : DFF_X1 port map( D => Key(45), CK => clk, Q => 
                           reg_key_45_port, QN => n_1307);
   reg_key_regx44x : DFF_X1 port map( D => Key(44), CK => clk, Q => 
                           reg_key_44_port, QN => n_1308);
   reg_key_regx43x : DFF_X1 port map( D => Key(43), CK => clk, Q => 
                           reg_key_43_port, QN => n_1309);
   reg_key_regx42x : DFF_X1 port map( D => Key(42), CK => clk, Q => 
                           reg_key_42_port, QN => n_1310);
   reg_key_regx40x : DFF_X1 port map( D => Key(40), CK => clk, Q => 
                           reg_key_40_port, QN => n_1311);
   reg_key_regx39x : DFF_X1 port map( D => Key(39), CK => clk, Q => 
                           reg_key_39_port, QN => n_1312);
   reg_key_regx38x : DFF_X1 port map( D => Key(38), CK => clk, Q => 
                           reg_key_38_port, QN => n_1313);
   reg_key_regx36x : DFF_X1 port map( D => Key(36), CK => clk, Q => 
                           reg_key_36_port, QN => n_1314);
   reg_key_regx35x : DFF_X1 port map( D => Key(35), CK => clk, Q => 
                           reg_key_35_port, QN => n_1315);
   reg_key_regx34x : DFF_X1 port map( D => Key(34), CK => clk, Q => 
                           reg_key_34_port, QN => n_1316);
   reg_key_regx33x : DFF_X1 port map( D => Key(33), CK => clk, Q => 
                           reg_key_33_port, QN => n_1317);
   reg_key_regx32x : DFF_X1 port map( D => Key(32), CK => clk, Q => 
                           reg_key_32_port, QN => n_1318);
   reg_key_regx31x : DFF_X1 port map( D => Key(31), CK => clk, Q => 
                           reg_key_31_port, QN => n_1319);
   reg_key_regx30x : DFF_X1 port map( D => Key(30), CK => clk, Q => 
                           reg_key_30_port, QN => n_1320);
   reg_key_regx29x : DFF_X1 port map( D => Key(29), CK => clk, Q => 
                           reg_key_29_port, QN => n_1321);
   reg_key_regx27x : DFF_X1 port map( D => Key(27), CK => clk, Q => 
                           reg_key_27_port, QN => n_1322);
   reg_key_regx26x : DFF_X1 port map( D => Key(26), CK => clk, Q => 
                           reg_key_26_port, QN => n_1323);
   reg_key_regx25x : DFF_X1 port map( D => Key(25), CK => clk, Q => 
                           reg_key_25_port, QN => n_1324);
   reg_key_regx24x : DFF_X1 port map( D => Key(24), CK => clk, Q => 
                           reg_key_24_port, QN => n_1325);
   reg_key_regx22x : DFF_X1 port map( D => Key(22), CK => clk, Q => 
                           reg_key_22_port, QN => n_1326);
   reg_key_regx21x : DFF_X1 port map( D => Key(21), CK => clk, Q => 
                           reg_key_21_port, QN => n_1327);
   reg_key_regx20x : DFF_X1 port map( D => Key(20), CK => clk, Q => 
                           reg_key_20_port, QN => n_1328);
   reg_key_regx19x : DFF_X1 port map( D => Key(19), CK => clk, Q => 
                           reg_key_19_port, QN => n_1329);
   reg_key_regx18x : DFF_X1 port map( D => Key(18), CK => clk, Q => 
                           reg_key_18_port, QN => n_1330);
   reg_key_regx17x : DFF_X1 port map( D => Key(17), CK => clk, Q => 
                           reg_key_17_port, QN => n_1331);
   reg_key_regx16x : DFF_X1 port map( D => Key(16), CK => clk, Q => 
                           reg_key_16_port, QN => n_1332);
   reg_key_regx15x : DFF_X1 port map( D => Key(15), CK => clk, Q => 
                           reg_key_15_port, QN => n_1333);
   reg_key_regx14x : DFF_X1 port map( D => Key(14), CK => clk, Q => 
                           reg_key_14_port, QN => n_1334);
   reg_key_regx12x : DFF_X1 port map( D => Key(12), CK => clk, Q => 
                           reg_key_12_port, QN => n_1335);
   reg_key_regx11x : DFF_X1 port map( D => Key(11), CK => clk, Q => 
                           reg_key_11_port, QN => n_1336);
   reg_key_regx10x : DFF_X1 port map( D => Key(10), CK => clk, Q => 
                           reg_key_10_port, QN => n_1337);
   reg_key_regx9x : DFF_X1 port map( D => Key(9), CK => clk, Q => 
                           reg_key_9_port, QN => n_1338);
   reg_key_regx8x : DFF_X1 port map( D => Key(8), CK => clk, Q => 
                           reg_key_8_port, QN => n_1339);
   reg_key_regx7x : DFF_X1 port map( D => Key(7), CK => clk, Q => 
                           reg_key_7_port, QN => n_1340);
   reg_key_regx6x : DFF_X1 port map( D => Key(6), CK => clk, Q => 
                           reg_key_6_port, QN => n_1341);
   reg_key_regx5x : DFF_X1 port map( D => Key(5), CK => clk, Q => 
                           reg_key_5_port, QN => n_1342);
   reg_key_regx4x : DFF_X1 port map( D => Key(4), CK => clk, Q => 
                           reg_key_4_port, QN => n_1343);
   reg_key_regx3x : DFF_X1 port map( D => Key(3), CK => clk, Q => 
                           reg_key_3_port, QN => n_1344);
   reg_key_regx2x : DFF_X1 port map( D => Key(2), CK => clk, Q => 
                           reg_key_2_port, QN => n_1345);
   reg_key_regx1x : DFF_X1 port map( D => Key(1), CK => clk, Q => 
                           reg_key_1_port, QN => n_1346);
   reg_key_regx0x : DFF_X1 port map( D => Key(0), CK => clk, Q => 
                           reg_key_0_port, QN => n_1347);
   Ciphertext_regx191x : DFF_X1 port map( D => reg_out_191_port, CK => clk, Q 
                           => Ciphertext(191), QN => n_1348);
   Ciphertext_regx190x : DFF_X1 port map( D => reg_out_190_port, CK => clk, Q 
                           => Ciphertext(190), QN => n_1349);
   Ciphertext_regx189x : DFF_X1 port map( D => reg_out_189_port, CK => clk, Q 
                           => Ciphertext(189), QN => n_1350);
   Ciphertext_regx188x : DFF_X1 port map( D => reg_out_188_port, CK => clk, Q 
                           => Ciphertext(188), QN => n_1351);
   Ciphertext_regx187x : DFF_X1 port map( D => reg_out_187_port, CK => clk, Q 
                           => Ciphertext(187), QN => n_1352);
   Ciphertext_regx186x : DFF_X1 port map( D => reg_out_186_port, CK => clk, Q 
                           => Ciphertext(186), QN => n_1353);
   Ciphertext_regx185x : DFF_X1 port map( D => reg_out_185_port, CK => clk, Q 
                           => Ciphertext(185), QN => n_1354);
   Ciphertext_regx184x : DFF_X1 port map( D => reg_out_184_port, CK => clk, Q 
                           => Ciphertext(184), QN => n_1355);
   Ciphertext_regx183x : DFF_X1 port map( D => reg_out_183_port, CK => clk, Q 
                           => Ciphertext(183), QN => n_1356);
   Ciphertext_regx182x : DFF_X1 port map( D => reg_out_182_port, CK => clk, Q 
                           => Ciphertext(182), QN => n_1357);
   Ciphertext_regx181x : DFF_X1 port map( D => reg_out_181_port, CK => clk, Q 
                           => Ciphertext(181), QN => n_1358);
   Ciphertext_regx180x : DFF_X1 port map( D => reg_out_180_port, CK => clk, Q 
                           => Ciphertext(180), QN => n_1359);
   Ciphertext_regx179x : DFF_X1 port map( D => reg_out_179_port, CK => clk, Q 
                           => Ciphertext(179), QN => n_1360);
   Ciphertext_regx178x : DFF_X1 port map( D => reg_out_178_port, CK => clk, Q 
                           => Ciphertext(178), QN => n_1361);
   Ciphertext_regx177x : DFF_X1 port map( D => reg_out_177_port, CK => clk, Q 
                           => Ciphertext(177), QN => n_1362);
   Ciphertext_regx176x : DFF_X1 port map( D => reg_out_176_port, CK => clk, Q 
                           => Ciphertext(176), QN => n_1363);
   Ciphertext_regx175x : DFF_X1 port map( D => reg_out_175_port, CK => clk, Q 
                           => Ciphertext(175), QN => n_1364);
   Ciphertext_regx174x : DFF_X1 port map( D => reg_out_174_port, CK => clk, Q 
                           => Ciphertext(174), QN => n_1365);
   Ciphertext_regx173x : DFF_X1 port map( D => reg_out_173_port, CK => clk, Q 
                           => Ciphertext(173), QN => n_1366);
   Ciphertext_regx172x : DFF_X1 port map( D => reg_out_172_port, CK => clk, Q 
                           => Ciphertext(172), QN => n_1367);
   Ciphertext_regx171x : DFF_X1 port map( D => reg_out_171_port, CK => clk, Q 
                           => Ciphertext(171), QN => n_1368);
   Ciphertext_regx170x : DFF_X1 port map( D => reg_out_170_port, CK => clk, Q 
                           => Ciphertext(170), QN => n_1369);
   Ciphertext_regx169x : DFF_X1 port map( D => reg_out_169_port, CK => clk, Q 
                           => Ciphertext(169), QN => n_1370);
   Ciphertext_regx168x : DFF_X1 port map( D => reg_out_168_port, CK => clk, Q 
                           => Ciphertext(168), QN => n_1371);
   Ciphertext_regx167x : DFF_X1 port map( D => reg_out_167_port, CK => clk, Q 
                           => Ciphertext(167), QN => n_1372);
   Ciphertext_regx166x : DFF_X1 port map( D => reg_out_166_port, CK => clk, Q 
                           => Ciphertext(166), QN => n_1373);
   Ciphertext_regx165x : DFF_X1 port map( D => reg_out_165_port, CK => clk, Q 
                           => Ciphertext(165), QN => n_1374);
   Ciphertext_regx164x : DFF_X1 port map( D => reg_out_164_port, CK => clk, Q 
                           => Ciphertext(164), QN => n_1375);
   Ciphertext_regx162x : DFF_X1 port map( D => reg_out_162_port, CK => clk, Q 
                           => Ciphertext(162), QN => n_1376);
   Ciphertext_regx161x : DFF_X1 port map( D => reg_out_161_port, CK => clk, Q 
                           => Ciphertext(161), QN => n_1377);
   Ciphertext_regx159x : DFF_X1 port map( D => reg_out_159_port, CK => clk, Q 
                           => Ciphertext(159), QN => n_1378);
   Ciphertext_regx158x : DFF_X1 port map( D => reg_out_158_port, CK => clk, Q 
                           => Ciphertext(158), QN => n_1379);
   Ciphertext_regx157x : DFF_X1 port map( D => reg_out_157_port, CK => clk, Q 
                           => Ciphertext(157), QN => n_1380);
   Ciphertext_regx155x : DFF_X1 port map( D => reg_out_155_port, CK => clk, Q 
                           => Ciphertext(155), QN => n_1381);
   Ciphertext_regx154x : DFF_X1 port map( D => reg_out_154_port, CK => clk, Q 
                           => Ciphertext(154), QN => n_1382);
   Ciphertext_regx153x : DFF_X1 port map( D => reg_out_153_port, CK => clk, Q 
                           => Ciphertext(153), QN => n_1383);
   Ciphertext_regx152x : DFF_X1 port map( D => reg_out_152_port, CK => clk, Q 
                           => Ciphertext(152), QN => n_1384);
   Ciphertext_regx151x : DFF_X1 port map( D => reg_out_151_port, CK => clk, Q 
                           => Ciphertext(151), QN => n_1385);
   Ciphertext_regx150x : DFF_X1 port map( D => reg_out_150_port, CK => clk, Q 
                           => Ciphertext(150), QN => n_1386);
   Ciphertext_regx149x : DFF_X1 port map( D => reg_out_149_port, CK => clk, Q 
                           => Ciphertext(149), QN => n_1387);
   Ciphertext_regx148x : DFF_X1 port map( D => reg_out_148_port, CK => clk, Q 
                           => Ciphertext(148), QN => n_1388);
   Ciphertext_regx147x : DFF_X1 port map( D => reg_out_147_port, CK => clk, Q 
                           => Ciphertext(147), QN => n_1389);
   Ciphertext_regx146x : DFF_X1 port map( D => reg_out_146_port, CK => clk, Q 
                           => Ciphertext(146), QN => n_1390);
   Ciphertext_regx145x : DFF_X1 port map( D => reg_out_145_port, CK => clk, Q 
                           => Ciphertext(145), QN => n_1391);
   Ciphertext_regx144x : DFF_X1 port map( D => reg_out_144_port, CK => clk, Q 
                           => Ciphertext(144), QN => n_1392);
   Ciphertext_regx143x : DFF_X1 port map( D => reg_out_143_port, CK => clk, Q 
                           => Ciphertext(143), QN => n_1393);
   Ciphertext_regx142x : DFF_X1 port map( D => reg_out_142_port, CK => clk, Q 
                           => Ciphertext(142), QN => n_1394);
   Ciphertext_regx141x : DFF_X1 port map( D => reg_out_141_port, CK => clk, Q 
                           => Ciphertext(141), QN => n_1395);
   Ciphertext_regx140x : DFF_X1 port map( D => reg_out_140_port, CK => clk, Q 
                           => Ciphertext(140), QN => n_1396);
   Ciphertext_regx139x : DFF_X1 port map( D => reg_out_139_port, CK => clk, Q 
                           => Ciphertext(139), QN => n_1397);
   Ciphertext_regx138x : DFF_X1 port map( D => reg_out_138_port, CK => clk, Q 
                           => Ciphertext(138), QN => n_1398);
   Ciphertext_regx137x : DFF_X1 port map( D => reg_out_137_port, CK => clk, Q 
                           => Ciphertext(137), QN => n_1399);
   Ciphertext_regx136x : DFF_X1 port map( D => reg_out_136_port, CK => clk, Q 
                           => Ciphertext(136), QN => n_1400);
   Ciphertext_regx135x : DFF_X1 port map( D => reg_out_135_port, CK => clk, Q 
                           => Ciphertext(135), QN => n_1401);
   Ciphertext_regx134x : DFF_X1 port map( D => reg_out_134_port, CK => clk, Q 
                           => Ciphertext(134), QN => n_1402);
   Ciphertext_regx133x : DFF_X1 port map( D => reg_out_133_port, CK => clk, Q 
                           => Ciphertext(133), QN => n_1403);
   Ciphertext_regx132x : DFF_X1 port map( D => reg_out_132_port, CK => clk, Q 
                           => Ciphertext(132), QN => n_1404);
   Ciphertext_regx131x : DFF_X1 port map( D => reg_out_131_port, CK => clk, Q 
                           => Ciphertext(131), QN => n_1405);
   Ciphertext_regx130x : DFF_X1 port map( D => reg_out_130_port, CK => clk, Q 
                           => Ciphertext(130), QN => n_1406);
   Ciphertext_regx129x : DFF_X1 port map( D => reg_out_129_port, CK => clk, Q 
                           => Ciphertext(129), QN => n_1407);
   Ciphertext_regx128x : DFF_X1 port map( D => reg_out_128_port, CK => clk, Q 
                           => Ciphertext(128), QN => n_1408);
   Ciphertext_regx127x : DFF_X1 port map( D => reg_out_127_port, CK => clk, Q 
                           => Ciphertext(127), QN => n_1409);
   Ciphertext_regx126x : DFF_X1 port map( D => reg_out_126_port, CK => clk, Q 
                           => Ciphertext(126), QN => n_1410);
   Ciphertext_regx125x : DFF_X1 port map( D => reg_out_125_port, CK => clk, Q 
                           => Ciphertext(125), QN => n_1411);
   Ciphertext_regx124x : DFF_X1 port map( D => reg_out_124_port, CK => clk, Q 
                           => Ciphertext(124), QN => n_1412);
   Ciphertext_regx123x : DFF_X1 port map( D => reg_out_123_port, CK => clk, Q 
                           => Ciphertext(123), QN => n_1413);
   Ciphertext_regx122x : DFF_X1 port map( D => reg_out_122_port, CK => clk, Q 
                           => Ciphertext(122), QN => n_1414);
   Ciphertext_regx121x : DFF_X1 port map( D => reg_out_121_port, CK => clk, Q 
                           => Ciphertext(121), QN => n_1415);
   Ciphertext_regx120x : DFF_X1 port map( D => reg_out_120_port, CK => clk, Q 
                           => Ciphertext(120), QN => n_1416);
   Ciphertext_regx119x : DFF_X1 port map( D => reg_out_119_port, CK => clk, Q 
                           => Ciphertext(119), QN => n_1417);
   Ciphertext_regx118x : DFF_X1 port map( D => reg_out_118_port, CK => clk, Q 
                           => Ciphertext(118), QN => n_1418);
   Ciphertext_regx117x : DFF_X1 port map( D => reg_out_117_port, CK => clk, Q 
                           => Ciphertext(117), QN => n_1419);
   Ciphertext_regx116x : DFF_X1 port map( D => reg_out_116_port, CK => clk, Q 
                           => Ciphertext(116), QN => n_1420);
   Ciphertext_regx114x : DFF_X1 port map( D => reg_out_114_port, CK => clk, Q 
                           => Ciphertext(114), QN => n_1421);
   Ciphertext_regx113x : DFF_X1 port map( D => reg_out_113_port, CK => clk, Q 
                           => Ciphertext(113), QN => n_1422);
   Ciphertext_regx112x : DFF_X1 port map( D => reg_out_112_port, CK => clk, Q 
                           => Ciphertext(112), QN => n_1423);
   Ciphertext_regx111x : DFF_X1 port map( D => reg_out_111_port, CK => clk, Q 
                           => Ciphertext(111), QN => n_1424);
   Ciphertext_regx110x : DFF_X1 port map( D => reg_out_110_port, CK => clk, Q 
                           => Ciphertext(110), QN => n_1425);
   Ciphertext_regx109x : DFF_X1 port map( D => reg_out_109_port, CK => clk, Q 
                           => Ciphertext(109), QN => n_1426);
   Ciphertext_regx108x : DFF_X1 port map( D => reg_out_108_port, CK => clk, Q 
                           => Ciphertext(108), QN => n_1427);
   Ciphertext_regx107x : DFF_X1 port map( D => reg_out_107_port, CK => clk, Q 
                           => Ciphertext(107), QN => n_1428);
   Ciphertext_regx106x : DFF_X1 port map( D => reg_out_106_port, CK => clk, Q 
                           => Ciphertext(106), QN => n_1429);
   Ciphertext_regx105x : DFF_X1 port map( D => reg_out_105_port, CK => clk, Q 
                           => Ciphertext(105), QN => n_1430);
   Ciphertext_regx104x : DFF_X1 port map( D => reg_out_104_port, CK => clk, Q 
                           => Ciphertext(104), QN => n_1431);
   Ciphertext_regx103x : DFF_X1 port map( D => reg_out_103_port, CK => clk, Q 
                           => Ciphertext(103), QN => n_1432);
   Ciphertext_regx102x : DFF_X1 port map( D => reg_out_102_port, CK => clk, Q 
                           => Ciphertext(102), QN => n_1433);
   Ciphertext_regx101x : DFF_X1 port map( D => reg_out_101_port, CK => clk, Q 
                           => Ciphertext(101), QN => n_1434);
   Ciphertext_regx100x : DFF_X1 port map( D => reg_out_100_port, CK => clk, Q 
                           => Ciphertext(100), QN => n_1435);
   Ciphertext_regx98x : DFF_X1 port map( D => reg_out_98_port, CK => clk, Q => 
                           Ciphertext(98), QN => n_1436);
   Ciphertext_regx97x : DFF_X1 port map( D => reg_out_97_port, CK => clk, Q => 
                           Ciphertext(97), QN => n_1437);
   Ciphertext_regx96x : DFF_X1 port map( D => reg_out_96_port, CK => clk, Q => 
                           Ciphertext(96), QN => n_1438);
   Ciphertext_regx95x : DFF_X1 port map( D => reg_out_95_port, CK => clk, Q => 
                           Ciphertext(95), QN => n_1439);
   Ciphertext_regx94x : DFF_X1 port map( D => reg_out_94_port, CK => clk, Q => 
                           Ciphertext(94), QN => n_1440);
   Ciphertext_regx93x : DFF_X1 port map( D => reg_out_93_port, CK => clk, Q => 
                           Ciphertext(93), QN => n_1441);
   Ciphertext_regx91x : DFF_X1 port map( D => reg_out_91_port, CK => clk, Q => 
                           Ciphertext(91), QN => n_1442);
   Ciphertext_regx90x : DFF_X1 port map( D => reg_out_90_port, CK => clk, Q => 
                           Ciphertext(90), QN => n_1443);
   Ciphertext_regx89x : DFF_X1 port map( D => reg_out_89_port, CK => clk, Q => 
                           Ciphertext(89), QN => n_1444);
   Ciphertext_regx88x : DFF_X1 port map( D => reg_out_88_port, CK => clk, Q => 
                           Ciphertext(88), QN => n_1445);
   Ciphertext_regx86x : DFF_X1 port map( D => reg_out_86_port, CK => clk, Q => 
                           Ciphertext(86), QN => n_1446);
   Ciphertext_regx85x : DFF_X1 port map( D => reg_out_85_port, CK => clk, Q => 
                           Ciphertext(85), QN => n_1447);
   Ciphertext_regx84x : DFF_X1 port map( D => reg_out_84_port, CK => clk, Q => 
                           Ciphertext(84), QN => n_1448);
   Ciphertext_regx83x : DFF_X1 port map( D => reg_out_83_port, CK => clk, Q => 
                           Ciphertext(83), QN => n_1449);
   Ciphertext_regx82x : DFF_X1 port map( D => reg_out_82_port, CK => clk, Q => 
                           Ciphertext(82), QN => n_1450);
   Ciphertext_regx81x : DFF_X1 port map( D => reg_out_81_port, CK => clk, Q => 
                           Ciphertext(81), QN => n_1451);
   Ciphertext_regx80x : DFF_X1 port map( D => reg_out_80_port, CK => clk, Q => 
                           Ciphertext(80), QN => n_1452);
   Ciphertext_regx78x : DFF_X1 port map( D => reg_out_78_port, CK => clk, Q => 
                           Ciphertext(78), QN => n_1453);
   Ciphertext_regx77x : DFF_X1 port map( D => reg_out_77_port, CK => clk, Q => 
                           Ciphertext(77), QN => n_1454);
   Ciphertext_regx76x : DFF_X1 port map( D => reg_out_76_port, CK => clk, Q => 
                           Ciphertext(76), QN => n_1455);
   Ciphertext_regx75x : DFF_X1 port map( D => reg_out_75_port, CK => clk, Q => 
                           Ciphertext(75), QN => n_1456);
   Ciphertext_regx74x : DFF_X1 port map( D => reg_out_74_port, CK => clk, Q => 
                           Ciphertext(74), QN => n_1457);
   Ciphertext_regx73x : DFF_X1 port map( D => reg_out_73_port, CK => clk, Q => 
                           Ciphertext(73), QN => n_1458);
   Ciphertext_regx72x : DFF_X1 port map( D => reg_out_72_port, CK => clk, Q => 
                           Ciphertext(72), QN => n_1459);
   Ciphertext_regx71x : DFF_X1 port map( D => reg_out_71_port, CK => clk, Q => 
                           Ciphertext(71), QN => n_1460);
   Ciphertext_regx70x : DFF_X1 port map( D => reg_out_70_port, CK => clk, Q => 
                           Ciphertext(70), QN => n_1461);
   Ciphertext_regx69x : DFF_X1 port map( D => reg_out_69_port, CK => clk, Q => 
                           Ciphertext(69), QN => n_1462);
   Ciphertext_regx68x : DFF_X1 port map( D => reg_out_68_port, CK => clk, Q => 
                           Ciphertext(68), QN => n_1463);
   Ciphertext_regx67x : DFF_X1 port map( D => reg_out_67_port, CK => clk, Q => 
                           Ciphertext(67), QN => n_1464);
   Ciphertext_regx66x : DFF_X1 port map( D => reg_out_66_port, CK => clk, Q => 
                           Ciphertext(66), QN => n_1465);
   Ciphertext_regx65x : DFF_X1 port map( D => reg_out_65_port, CK => clk, Q => 
                           Ciphertext(65), QN => n_1466);
   Ciphertext_regx64x : DFF_X1 port map( D => reg_out_64_port, CK => clk, Q => 
                           Ciphertext(64), QN => n_1467);
   Ciphertext_regx63x : DFF_X1 port map( D => reg_out_63_port, CK => clk, Q => 
                           Ciphertext(63), QN => n_1468);
   Ciphertext_regx62x : DFF_X1 port map( D => reg_out_62_port, CK => clk, Q => 
                           Ciphertext(62), QN => n_1469);
   Ciphertext_regx61x : DFF_X1 port map( D => reg_out_61_port, CK => clk, Q => 
                           Ciphertext(61), QN => n_1470);
   Ciphertext_regx60x : DFF_X1 port map( D => reg_out_60_port, CK => clk, Q => 
                           Ciphertext(60), QN => n_1471);
   Ciphertext_regx59x : DFF_X1 port map( D => reg_out_59_port, CK => clk, Q => 
                           Ciphertext(59), QN => n_1472);
   Ciphertext_regx57x : DFF_X1 port map( D => reg_out_57_port, CK => clk, Q => 
                           Ciphertext(57), QN => n_1473);
   Ciphertext_regx56x : DFF_X1 port map( D => reg_out_56_port, CK => clk, Q => 
                           Ciphertext(56), QN => n_1474);
   Ciphertext_regx55x : DFF_X1 port map( D => reg_out_55_port, CK => clk, Q => 
                           Ciphertext(55), QN => n_1475);
   Ciphertext_regx54x : DFF_X1 port map( D => reg_out_54_port, CK => clk, Q => 
                           Ciphertext(54), QN => n_1476);
   Ciphertext_regx53x : DFF_X1 port map( D => reg_out_53_port, CK => clk, Q => 
                           Ciphertext(53), QN => n_1477);
   Ciphertext_regx52x : DFF_X1 port map( D => reg_out_52_port, CK => clk, Q => 
                           Ciphertext(52), QN => n_1478);
   Ciphertext_regx51x : DFF_X1 port map( D => reg_out_51_port, CK => clk, Q => 
                           Ciphertext(51), QN => n_1479);
   Ciphertext_regx50x : DFF_X1 port map( D => reg_out_50_port, CK => clk, Q => 
                           Ciphertext(50), QN => n_1480);
   Ciphertext_regx49x : DFF_X1 port map( D => reg_out_49_port, CK => clk, Q => 
                           Ciphertext(49), QN => n_1481);
   Ciphertext_regx48x : DFF_X1 port map( D => reg_out_48_port, CK => clk, Q => 
                           Ciphertext(48), QN => n_1482);
   Ciphertext_regx47x : DFF_X1 port map( D => reg_out_47_port, CK => clk, Q => 
                           Ciphertext(47), QN => n_1483);
   Ciphertext_regx46x : DFF_X1 port map( D => reg_out_46_port, CK => clk, Q => 
                           Ciphertext(46), QN => n_1484);
   Ciphertext_regx45x : DFF_X1 port map( D => reg_out_45_port, CK => clk, Q => 
                           Ciphertext(45), QN => n_1485);
   Ciphertext_regx44x : DFF_X1 port map( D => reg_out_44_port, CK => clk, Q => 
                           Ciphertext(44), QN => n_1486);
   Ciphertext_regx43x : DFF_X1 port map( D => reg_out_43_port, CK => clk, Q => 
                           Ciphertext(43), QN => n_1487);
   Ciphertext_regx42x : DFF_X1 port map( D => reg_out_42_port, CK => clk, Q => 
                           Ciphertext(42), QN => n_1488);
   Ciphertext_regx41x : DFF_X1 port map( D => reg_out_41_port, CK => clk, Q => 
                           Ciphertext(41), QN => n_1489);
   Ciphertext_regx39x : DFF_X1 port map( D => reg_out_39_port, CK => clk, Q => 
                           Ciphertext(39), QN => n_1490);
   Ciphertext_regx38x : DFF_X1 port map( D => reg_out_38_port, CK => clk, Q => 
                           Ciphertext(38), QN => n_1491);
   Ciphertext_regx37x : DFF_X1 port map( D => reg_out_37_port, CK => clk, Q => 
                           Ciphertext(37), QN => n_1492);
   Ciphertext_regx36x : DFF_X1 port map( D => reg_out_36_port, CK => clk, Q => 
                           Ciphertext(36), QN => n_1493);
   Ciphertext_regx35x : DFF_X1 port map( D => reg_out_35_port, CK => clk, Q => 
                           Ciphertext(35), QN => n_1494);
   Ciphertext_regx34x : DFF_X1 port map( D => reg_out_34_port, CK => clk, Q => 
                           Ciphertext(34), QN => n_1495);
   Ciphertext_regx32x : DFF_X1 port map( D => reg_out_32_port, CK => clk, Q => 
                           Ciphertext(32), QN => n_1496);
   Ciphertext_regx31x : DFF_X1 port map( D => reg_out_31_port, CK => clk, Q => 
                           Ciphertext(31), QN => n_1497);
   Ciphertext_regx30x : DFF_X1 port map( D => reg_out_30_port, CK => clk, Q => 
                           Ciphertext(30), QN => n_1498);
   Ciphertext_regx29x : DFF_X1 port map( D => reg_out_29_port, CK => clk, Q => 
                           Ciphertext(29), QN => n_1499);
   Ciphertext_regx28x : DFF_X1 port map( D => reg_out_28_port, CK => clk, Q => 
                           Ciphertext(28), QN => n_1500);
   Ciphertext_regx27x : DFF_X1 port map( D => reg_out_27_port, CK => clk, Q => 
                           Ciphertext(27), QN => n_1501);
   Ciphertext_regx26x : DFF_X1 port map( D => reg_out_26_port, CK => clk, Q => 
                           Ciphertext(26), QN => n_1502);
   Ciphertext_regx25x : DFF_X1 port map( D => reg_out_25_port, CK => clk, Q => 
                           Ciphertext(25), QN => n_1503);
   Ciphertext_regx24x : DFF_X1 port map( D => reg_out_24_port, CK => clk, Q => 
                           Ciphertext(24), QN => n_1504);
   Ciphertext_regx23x : DFF_X1 port map( D => reg_out_23_port, CK => clk, Q => 
                           Ciphertext(23), QN => n_1505);
   Ciphertext_regx22x : DFF_X1 port map( D => reg_out_22_port, CK => clk, Q => 
                           Ciphertext(22), QN => n_1506);
   Ciphertext_regx21x : DFF_X1 port map( D => reg_out_21_port, CK => clk, Q => 
                           Ciphertext(21), QN => n_1507);
   Ciphertext_regx20x : DFF_X1 port map( D => reg_out_20_port, CK => clk, Q => 
                           Ciphertext(20), QN => n_1508);
   Ciphertext_regx19x : DFF_X1 port map( D => reg_out_19_port, CK => clk, Q => 
                           Ciphertext(19), QN => n_1509);
   Ciphertext_regx18x : DFF_X1 port map( D => reg_out_18_port, CK => clk, Q => 
                           Ciphertext(18), QN => n_1510);
   Ciphertext_regx17x : DFF_X1 port map( D => reg_out_17_port, CK => clk, Q => 
                           Ciphertext(17), QN => n_1511);
   Ciphertext_regx16x : DFF_X1 port map( D => reg_out_16_port, CK => clk, Q => 
                           Ciphertext(16), QN => n_1512);
   Ciphertext_regx15x : DFF_X1 port map( D => reg_out_15_port, CK => clk, Q => 
                           Ciphertext(15), QN => n_1513);
   Ciphertext_regx14x : DFF_X1 port map( D => reg_out_14_port, CK => clk, Q => 
                           Ciphertext(14), QN => n_1514);
   Ciphertext_regx13x : DFF_X1 port map( D => reg_out_13_port, CK => clk, Q => 
                           Ciphertext(13), QN => n_1515);
   Ciphertext_regx11x : DFF_X1 port map( D => reg_out_11_port, CK => clk, Q => 
                           Ciphertext(11), QN => n_1516);
   Ciphertext_regx10x : DFF_X1 port map( D => reg_out_10_port, CK => clk, Q => 
                           Ciphertext(10), QN => n_1517);
   Ciphertext_regx9x : DFF_X1 port map( D => reg_out_9_port, CK => clk, Q => 
                           Ciphertext(9), QN => n_1518);
   Ciphertext_regx7x : DFF_X1 port map( D => reg_out_7_port, CK => clk, Q => 
                           Ciphertext(7), QN => n_1519);
   Ciphertext_regx6x : DFF_X1 port map( D => reg_out_6_port, CK => clk, Q => 
                           Ciphertext(6), QN => n_1520);
   Ciphertext_regx5x : DFF_X1 port map( D => reg_out_5_port, CK => clk, Q => 
                           Ciphertext(5), QN => n_1521);
   Ciphertext_regx4x : DFF_X1 port map( D => reg_out_4_port, CK => clk, Q => 
                           Ciphertext(4), QN => n_1522);
   Ciphertext_regx2x : DFF_X1 port map( D => reg_out_2_port, CK => clk, Q => 
                           Ciphertext(2), QN => n_1523);
   Ciphertext_regx1x : DFF_X1 port map( D => reg_out_1_port, CK => clk, Q => 
                           Ciphertext(1), QN => n_1524);
   reg_key_regx179x : DFF_X1 port map( D => Key(179), CK => clk, Q => 
                           reg_key_179_port, QN => n_1525);
   reg_key_regx62x : DFF_X1 port map( D => Key(62), CK => clk, Q => 
                           reg_key_62_port, QN => n_1526);
   reg_key_regx113x : DFF_X1 port map( D => Key(113), CK => clk, Q => 
                           reg_key_113_port, QN => n_1527);
   reg_key_regx79x : DFF_X1 port map( D => Key(79), CK => clk, Q => 
                           reg_key_79_port, QN => n_1528);
   reg_key_regx183x : DFF_X1 port map( D => Key(183), CK => clk, Q => 
                           reg_key_183_port, QN => n_1529);
   reg_key_regx166x : DFF_X1 port map( D => Key(166), CK => clk, Q => 
                           reg_key_166_port, QN => n_1530);
   reg_key_regx107x : DFF_X1 port map( D => Key(107), CK => clk, Q => 
                           reg_key_107_port, QN => n_1531);
   reg_key_regx56x : DFF_X1 port map( D => Key(56), CK => clk, Q => 
                           reg_key_56_port, QN => n_1532);
   reg_key_regx187x : DFF_X1 port map( D => Key(187), CK => clk, Q => 
                           reg_key_187_port, QN => n_1533);
   reg_key_regx77x : DFF_X1 port map( D => Key(77), CK => clk, Q => 
                           reg_key_77_port, QN => n_1534);
   reg_key_regx23x : DFF_X1 port map( D => Key(23), CK => clk, Q => 
                           reg_key_23_port, QN => n_1535);
   Ciphertext_regx3x : DFFRS_X1 port map( D => reg_out_3_port, CK => clk, RN =>
                           n5, SN => n5, Q => Ciphertext(3), QN => n_1536);
   reg_key_regx83x : DFF_X1 port map( D => Key(83), CK => clk, Q => 
                           reg_key_83_port, QN => n_1537);
   reg_key_regx71x : DFF_X1 port map( D => Key(71), CK => clk, Q => 
                           reg_key_71_port, QN => n_1538);
   Ciphertext_regx156x : DFF_X1 port map( D => reg_out_156_port, CK => clk, Q 
                           => Ciphertext(156), QN => n_1539);
   reg_key_regx68x : DFF_X1 port map( D => Key(68), CK => clk, Q => 
                           reg_key_68_port, QN => n_1540);
   reg_key_regx171x : DFF_X1 port map( D => Key(171), CK => clk, Q => 
                           reg_key_171_port, QN => n_1541);
   reg_key_regx13x : DFF_X1 port map( D => Key(13), CK => clk, Q => 
                           reg_key_13_port, QN => n_1542);
   reg_key_regx165x : DFF_X1 port map( D => Key(165), CK => clk, Q => 
                           reg_key_165_port, QN => n_1543);
   reg_key_regx64x : DFF_X1 port map( D => Key(64), CK => clk, Q => 
                           reg_key_64_port, QN => n_1544);
   reg_key_regx63x : DFF_X1 port map( D => Key(63), CK => clk, Q => 
                           reg_key_63_port, QN => n_1545);
   reg_key_regx126x : DFF_X1 port map( D => Key(126), CK => clk, Q => 
                           reg_key_126_port, QN => n_1546);
   reg_key_regx185x : DFF_X1 port map( D => Key(185), CK => clk, Q => 
                           reg_key_185_port, QN => n_1547);
   reg_key_regx134x : DFF_X1 port map( D => Key(134), CK => clk, Q => 
                           reg_key_134_port, QN => n_1548);
   reg_key_regx182x : DFF_X1 port map( D => Key(182), CK => clk, Q => 
                           reg_key_182_port, QN => n_1549);
   reg_key_regx65x : DFF_X1 port map( D => Key(65), CK => clk, Q => 
                           reg_key_65_port, QN => n_1550);
   reg_key_regx37x : DFF_X1 port map( D => Key(37), CK => clk, Q => 
                           reg_key_37_port, QN => n_1551);
   reg_key_regx89x : DFF_X1 port map( D => Key(89), CK => clk, Q => 
                           reg_key_89_port, QN => n_1552);
   reg_key_regx105x : DFF_X1 port map( D => Key(105), CK => clk, Q => 
                           reg_key_105_port, QN => n_1553);
   reg_key_regx110x : DFF_X1 port map( D => Key(110), CK => clk, Q => 
                           reg_key_110_port, QN => n_1554);
   reg_key_regx52x : DFF_X1 port map( D => Key(52), CK => clk, Q => 
                           reg_key_52_port, QN => n_1555);
   reg_key_regx86x : DFF_X1 port map( D => Key(86), CK => clk, Q => 
                           reg_key_86_port, QN => n_1556);
   reg_key_regx28x : DFF_X1 port map( D => Key(28), CK => clk, Q => 
                           reg_key_28_port, QN => n_1557);
   reg_key_regx150x : DFF_X1 port map( D => Key(150), CK => clk, Q => 
                           reg_key_150_port, QN => n_1558);
   reg_key_regx87x : DFF_X1 port map( D => Key(87), CK => clk, Q => 
                           reg_key_87_port, QN => n_1559);
   reg_key_regx46x : DFF_X1 port map( D => Key(46), CK => clk, Q => 
                           reg_key_46_port, QN => n_1560);
   reg_key_regx41x : DFF_X1 port map( D => Key(41), CK => clk, Q => 
                           reg_key_41_port, QN => n_1561);
   n5 <= '1';
   Ciphertext_regx115x : DFF_X2 port map( D => reg_out_115_port, CK => clk, Q 
                           => Ciphertext(115), QN => n_1562);
   Ciphertext_regx33x : DFF_X1 port map( D => reg_out_33_port, CK => clk, Q => 
                           Ciphertext(33), QN => n_1563);
   Ciphertext_regx79x : DFF_X1 port map( D => reg_out_79_port, CK => clk, Q => 
                           Ciphertext(79), QN => n_1564);
   Ciphertext_regx87x : DFF_X1 port map( D => reg_out_87_port, CK => clk, Q => 
                           Ciphertext(87), QN => n_1565);
   Ciphertext_regx58x : DFFRS_X1 port map( D => reg_out_58_port, CK => clk, RN 
                           => n9, SN => n9, Q => Ciphertext(58), QN => n_1566);
   Ciphertext_regx0x : DFF_X1 port map( D => reg_out_0_port, CK => clk, Q => 
                           Ciphertext(0), QN => n_1567);
   Ciphertext_regx92x : DFF_X1 port map( D => reg_out_92_port, CK => clk, Q => 
                           Ciphertext(92), QN => n_1568);
   Ciphertext_regx160x : DFF_X1 port map( D => reg_out_160_port, CK => clk, Q 
                           => Ciphertext(160), QN => n_1569);
   n9 <= '1';
   SPEEDY_instance : SPEEDY_Rounds5_0 port map( Plaintext(191) => 
                           reg_in_191_port, Plaintext(190) => reg_in_190_port, 
                           Plaintext(189) => reg_in_189_port, Plaintext(188) =>
                           reg_in_188_port, Plaintext(187) => reg_in_187_port, 
                           Plaintext(186) => reg_in_186_port, Plaintext(185) =>
                           reg_in_185_port, Plaintext(184) => reg_in_184_port, 
                           Plaintext(183) => reg_in_183_port, Plaintext(182) =>
                           reg_in_182_port, Plaintext(181) => reg_in_181_port, 
                           Plaintext(180) => reg_in_180_port, Plaintext(179) =>
                           reg_in_179_port, Plaintext(178) => reg_in_178_port, 
                           Plaintext(177) => reg_in_177_port, Plaintext(176) =>
                           reg_in_176_port, Plaintext(175) => reg_in_175_port, 
                           Plaintext(174) => reg_in_174_port, Plaintext(173) =>
                           reg_in_173_port, Plaintext(172) => reg_in_172_port, 
                           Plaintext(171) => reg_in_171_port, Plaintext(170) =>
                           reg_in_170_port, Plaintext(169) => reg_in_169_port, 
                           Plaintext(168) => reg_in_168_port, Plaintext(167) =>
                           reg_in_167_port, Plaintext(166) => reg_in_166_port, 
                           Plaintext(165) => reg_in_165_port, Plaintext(164) =>
                           reg_in_164_port, Plaintext(163) => reg_in_163_port, 
                           Plaintext(162) => reg_in_162_port, Plaintext(161) =>
                           reg_in_161_port, Plaintext(160) => reg_in_160_port, 
                           Plaintext(159) => reg_in_159_port, Plaintext(158) =>
                           reg_in_158_port, Plaintext(157) => reg_in_157_port, 
                           Plaintext(156) => reg_in_156_port, Plaintext(155) =>
                           reg_in_155_port, Plaintext(154) => reg_in_154_port, 
                           Plaintext(153) => reg_in_153_port, Plaintext(152) =>
                           reg_in_152_port, Plaintext(151) => reg_in_151_port, 
                           Plaintext(150) => reg_in_150_port, Plaintext(149) =>
                           reg_in_149_port, Plaintext(148) => reg_in_148_port, 
                           Plaintext(147) => reg_in_147_port, Plaintext(146) =>
                           reg_in_146_port, Plaintext(145) => reg_in_145_port, 
                           Plaintext(144) => reg_in_144_port, Plaintext(143) =>
                           reg_in_143_port, Plaintext(142) => reg_in_142_port, 
                           Plaintext(141) => reg_in_141_port, Plaintext(140) =>
                           reg_in_140_port, Plaintext(139) => reg_in_139_port, 
                           Plaintext(138) => reg_in_138_port, Plaintext(137) =>
                           reg_in_137_port, Plaintext(136) => reg_in_136_port, 
                           Plaintext(135) => reg_in_135_port, Plaintext(134) =>
                           reg_in_134_port, Plaintext(133) => reg_in_133_port, 
                           Plaintext(132) => reg_in_132_port, Plaintext(131) =>
                           reg_in_131_port, Plaintext(130) => reg_in_130_port, 
                           Plaintext(129) => reg_in_129_port, Plaintext(128) =>
                           reg_in_128_port, Plaintext(127) => reg_in_127_port, 
                           Plaintext(126) => reg_in_126_port, Plaintext(125) =>
                           reg_in_125_port, Plaintext(124) => reg_in_124_port, 
                           Plaintext(123) => reg_in_123_port, Plaintext(122) =>
                           reg_in_122_port, Plaintext(121) => reg_in_121_port, 
                           Plaintext(120) => reg_in_120_port, Plaintext(119) =>
                           reg_in_119_port, Plaintext(118) => reg_in_118_port, 
                           Plaintext(117) => reg_in_117_port, Plaintext(116) =>
                           reg_in_116_port, Plaintext(115) => reg_in_115_port, 
                           Plaintext(114) => reg_in_114_port, Plaintext(113) =>
                           reg_in_113_port, Plaintext(112) => reg_in_112_port, 
                           Plaintext(111) => reg_in_111_port, Plaintext(110) =>
                           reg_in_110_port, Plaintext(109) => reg_in_109_port, 
                           Plaintext(108) => reg_in_108_port, Plaintext(107) =>
                           reg_in_107_port, Plaintext(106) => reg_in_106_port, 
                           Plaintext(105) => reg_in_105_port, Plaintext(104) =>
                           reg_in_104_port, Plaintext(103) => reg_in_103_port, 
                           Plaintext(102) => reg_in_102_port, Plaintext(101) =>
                           reg_in_101_port, Plaintext(100) => reg_in_100_port, 
                           Plaintext(99) => reg_in_99_port, Plaintext(98) => 
                           reg_in_98_port, Plaintext(97) => reg_in_97_port, 
                           Plaintext(96) => reg_in_96_port, Plaintext(95) => 
                           reg_in_95_port, Plaintext(94) => reg_in_94_port, 
                           Plaintext(93) => reg_in_93_port, Plaintext(92) => 
                           reg_in_92_port, Plaintext(91) => reg_in_91_port, 
                           Plaintext(90) => reg_in_90_port, Plaintext(89) => 
                           reg_in_89_port, Plaintext(88) => reg_in_88_port, 
                           Plaintext(87) => reg_in_87_port, Plaintext(86) => 
                           reg_in_86_port, Plaintext(85) => reg_in_85_port, 
                           Plaintext(84) => reg_in_84_port, Plaintext(83) => 
                           reg_in_83_port, Plaintext(82) => reg_in_82_port, 
                           Plaintext(81) => reg_in_81_port, Plaintext(80) => 
                           reg_in_80_port, Plaintext(79) => reg_in_79_port, 
                           Plaintext(78) => reg_in_78_port, Plaintext(77) => 
                           reg_in_77_port, Plaintext(76) => reg_in_76_port, 
                           Plaintext(75) => reg_in_75_port, Plaintext(74) => 
                           reg_in_74_port, Plaintext(73) => reg_in_73_port, 
                           Plaintext(72) => reg_in_72_port, Plaintext(71) => 
                           reg_in_71_port, Plaintext(70) => reg_in_70_port, 
                           Plaintext(69) => reg_in_69_port, Plaintext(68) => 
                           reg_in_68_port, Plaintext(67) => reg_in_67_port, 
                           Plaintext(66) => reg_in_66_port, Plaintext(65) => 
                           reg_in_65_port, Plaintext(64) => reg_in_64_port, 
                           Plaintext(63) => reg_in_63_port, Plaintext(62) => 
                           reg_in_62_port, Plaintext(61) => reg_in_61_port, 
                           Plaintext(60) => reg_in_60_port, Plaintext(59) => 
                           reg_in_59_port, Plaintext(58) => reg_in_58_port, 
                           Plaintext(57) => reg_in_57_port, Plaintext(56) => 
                           reg_in_56_port, Plaintext(55) => reg_in_55_port, 
                           Plaintext(54) => reg_in_54_port, Plaintext(53) => 
                           reg_in_53_port, Plaintext(52) => reg_in_52_port, 
                           Plaintext(51) => reg_in_51_port, Plaintext(50) => 
                           reg_in_50_port, Plaintext(49) => reg_in_49_port, 
                           Plaintext(48) => reg_in_48_port, Plaintext(47) => 
                           reg_in_47_port, Plaintext(46) => reg_in_46_port, 
                           Plaintext(45) => reg_in_45_port, Plaintext(44) => 
                           reg_in_44_port, Plaintext(43) => reg_in_43_port, 
                           Plaintext(42) => reg_in_42_port, Plaintext(41) => 
                           reg_in_41_port, Plaintext(40) => reg_in_40_port, 
                           Plaintext(39) => reg_in_39_port, Plaintext(38) => 
                           reg_in_38_port, Plaintext(37) => reg_in_37_port, 
                           Plaintext(36) => reg_in_36_port, Plaintext(35) => 
                           reg_in_35_port, Plaintext(34) => reg_in_34_port, 
                           Plaintext(33) => reg_in_33_port, Plaintext(32) => 
                           reg_in_32_port, Plaintext(31) => reg_in_31_port, 
                           Plaintext(30) => reg_in_30_port, Plaintext(29) => 
                           reg_in_29_port, Plaintext(28) => reg_in_28_port, 
                           Plaintext(27) => reg_in_27_port, Plaintext(26) => 
                           reg_in_26_port, Plaintext(25) => reg_in_25_port, 
                           Plaintext(24) => reg_in_24_port, Plaintext(23) => 
                           reg_in_23_port, Plaintext(22) => reg_in_22_port, 
                           Plaintext(21) => reg_in_21_port, Plaintext(20) => 
                           reg_in_20_port, Plaintext(19) => reg_in_19_port, 
                           Plaintext(18) => reg_in_18_port, Plaintext(17) => 
                           reg_in_17_port, Plaintext(16) => reg_in_16_port, 
                           Plaintext(15) => reg_in_15_port, Plaintext(14) => 
                           reg_in_14_port, Plaintext(13) => reg_in_13_port, 
                           Plaintext(12) => reg_in_12_port, Plaintext(11) => 
                           reg_in_11_port, Plaintext(10) => reg_in_10_port, 
                           Plaintext(9) => reg_in_9_port, Plaintext(8) => 
                           reg_in_8_port, Plaintext(7) => reg_in_7_port, 
                           Plaintext(6) => reg_in_6_port, Plaintext(5) => 
                           reg_in_5_port, Plaintext(4) => reg_in_4_port, 
                           Plaintext(3) => reg_in_3_port, Plaintext(2) => 
                           reg_in_2_port, Plaintext(1) => reg_in_1_port, 
                           Plaintext(0) => reg_in_0_port, Key(191) => 
                           reg_key_191_port, Key(190) => reg_key_190_port, 
                           Key(189) => reg_key_189_port, Key(188) => 
                           reg_key_188_port, Key(187) => reg_key_187_port, 
                           Key(186) => n3, Key(185) => reg_key_185_port, 
                           Key(184) => reg_key_184_port, Key(183) => 
                           reg_key_183_port, Key(182) => reg_key_182_port, 
                           Key(181) => reg_key_181_port, Key(180) => 
                           reg_key_180_port, Key(179) => reg_key_179_port, 
                           Key(178) => reg_key_178_port, Key(177) => 
                           reg_key_177_port, Key(176) => reg_key_176_port, 
                           Key(175) => reg_key_175_port, Key(174) => 
                           reg_key_174_port, Key(173) => reg_key_173_port, 
                           Key(172) => reg_key_172_port, Key(171) => 
                           reg_key_171_port, Key(170) => reg_key_170_port, 
                           Key(169) => reg_key_169_port, Key(168) => 
                           reg_key_168_port, Key(167) => reg_key_167_port, 
                           Key(166) => reg_key_166_port, Key(165) => 
                           reg_key_165_port, Key(164) => reg_key_164_port, 
                           Key(163) => reg_key_163_port, Key(162) => 
                           reg_key_162_port, Key(161) => reg_key_161_port, 
                           Key(160) => reg_key_160_port, Key(159) => 
                           reg_key_159_port, Key(158) => reg_key_158_port, 
                           Key(157) => reg_key_157_port, Key(156) => 
                           reg_key_156_port, Key(155) => reg_key_155_port, 
                           Key(154) => reg_key_154_port, Key(153) => 
                           reg_key_153_port, Key(152) => reg_key_152_port, 
                           Key(151) => reg_key_151_port, Key(150) => 
                           reg_key_150_port, Key(149) => reg_key_149_port, 
                           Key(148) => reg_key_148_port, Key(147) => 
                           reg_key_147_port, Key(146) => reg_key_146_port, 
                           Key(145) => reg_key_145_port, Key(144) => 
                           reg_key_144_port, Key(143) => reg_key_143_port, 
                           Key(142) => reg_key_142_port, Key(141) => 
                           reg_key_141_port, Key(140) => reg_key_140_port, 
                           Key(139) => reg_key_139_port, Key(138) => 
                           reg_key_138_port, Key(137) => reg_key_137_port, 
                           Key(136) => reg_key_136_port, Key(135) => 
                           reg_key_135_port, Key(134) => reg_key_134_port, 
                           Key(133) => reg_key_133_port, Key(132) => 
                           reg_key_132_port, Key(131) => reg_key_131_port, 
                           Key(130) => reg_key_130_port, Key(129) => 
                           reg_key_129_port, Key(128) => reg_key_128_port, 
                           Key(127) => reg_key_127_port, Key(126) => 
                           reg_key_126_port, Key(125) => reg_key_125_port, 
                           Key(124) => reg_key_124_port, Key(123) => 
                           reg_key_123_port, Key(122) => reg_key_122_port, 
                           Key(121) => reg_key_121_port, Key(120) => 
                           reg_key_120_port, Key(119) => reg_key_119_port, 
                           Key(118) => reg_key_118_port, Key(117) => 
                           reg_key_117_port, Key(116) => reg_key_116_port, 
                           Key(115) => reg_key_115_port, Key(114) => 
                           reg_key_114_port, Key(113) => reg_key_113_port, 
                           Key(112) => reg_key_112_port, Key(111) => 
                           reg_key_111_port, Key(110) => reg_key_110_port, 
                           Key(109) => reg_key_109_port, Key(108) => 
                           reg_key_108_port, Key(107) => reg_key_107_port, 
                           Key(106) => reg_key_106_port, Key(105) => 
                           reg_key_105_port, Key(104) => reg_key_104_port, 
                           Key(103) => reg_key_103_port, Key(102) => 
                           reg_key_102_port, Key(101) => reg_key_101_port, 
                           Key(100) => reg_key_100_port, Key(99) => 
                           reg_key_99_port, Key(98) => reg_key_98_port, Key(97)
                           => reg_key_97_port, Key(96) => reg_key_96_port, 
                           Key(95) => reg_key_95_port, Key(94) => 
                           reg_key_94_port, Key(93) => reg_key_93_port, Key(92)
                           => reg_key_92_port, Key(91) => reg_key_91_port, 
                           Key(90) => reg_key_90_port, Key(89) => 
                           reg_key_89_port, Key(88) => reg_key_88_port, Key(87)
                           => reg_key_87_port, Key(86) => reg_key_86_port, 
                           Key(85) => reg_key_85_port, Key(84) => 
                           reg_key_84_port, Key(83) => reg_key_83_port, Key(82)
                           => reg_key_82_port, Key(81) => reg_key_81_port, 
                           Key(80) => reg_key_80_port, Key(79) => 
                           reg_key_79_port, Key(78) => reg_key_78_port, Key(77)
                           => reg_key_77_port, Key(76) => reg_key_76_port, 
                           Key(75) => reg_key_75_port, Key(74) => 
                           reg_key_74_port, Key(73) => reg_key_73_port, Key(72)
                           => reg_key_72_port, Key(71) => reg_key_71_port, 
                           Key(70) => reg_key_70_port, Key(69) => 
                           reg_key_69_port, Key(68) => reg_key_68_port, Key(67)
                           => reg_key_67_port, Key(66) => reg_key_66_port, 
                           Key(65) => reg_key_65_port, Key(64) => 
                           reg_key_64_port, Key(63) => reg_key_63_port, Key(62)
                           => reg_key_62_port, Key(61) => reg_key_61_port, 
                           Key(60) => reg_key_60_port, Key(59) => 
                           reg_key_59_port, Key(58) => reg_key_58_port, Key(57)
                           => reg_key_57_port, Key(56) => reg_key_56_port, 
                           Key(55) => reg_key_55_port, Key(54) => 
                           reg_key_54_port, Key(53) => reg_key_53_port, Key(52)
                           => reg_key_52_port, Key(51) => reg_key_51_port, 
                           Key(50) => reg_key_50_port, Key(49) => 
                           reg_key_49_port, Key(48) => reg_key_48_port, Key(47)
                           => reg_key_47_port, Key(46) => reg_key_46_port, 
                           Key(45) => reg_key_45_port, Key(44) => 
                           reg_key_44_port, Key(43) => reg_key_43_port, Key(42)
                           => reg_key_42_port, Key(41) => reg_key_41_port, 
                           Key(40) => reg_key_40_port, Key(39) => 
                           reg_key_39_port, Key(38) => reg_key_38_port, Key(37)
                           => reg_key_37_port, Key(36) => reg_key_36_port, 
                           Key(35) => reg_key_35_port, Key(34) => 
                           reg_key_34_port, Key(33) => reg_key_33_port, Key(32)
                           => reg_key_32_port, Key(31) => reg_key_31_port, 
                           Key(30) => reg_key_30_port, Key(29) => 
                           reg_key_29_port, Key(28) => reg_key_28_port, Key(27)
                           => reg_key_27_port, Key(26) => reg_key_26_port, 
                           Key(25) => reg_key_25_port, Key(24) => 
                           reg_key_24_port, Key(23) => reg_key_23_port, Key(22)
                           => reg_key_22_port, Key(21) => reg_key_21_port, 
                           Key(20) => reg_key_20_port, Key(19) => 
                           reg_key_19_port, Key(18) => reg_key_18_port, Key(17)
                           => reg_key_17_port, Key(16) => reg_key_16_port, 
                           Key(15) => reg_key_15_port, Key(14) => 
                           reg_key_14_port, Key(13) => reg_key_13_port, Key(12)
                           => reg_key_12_port, Key(11) => reg_key_11_port, 
                           Key(10) => reg_key_10_port, Key(9) => reg_key_9_port
                           , Key(8) => reg_key_8_port, Key(7) => reg_key_7_port
                           , Key(6) => reg_key_6_port, Key(5) => reg_key_5_port
                           , Key(4) => reg_key_4_port, Key(3) => reg_key_3_port
                           , Key(2) => reg_key_2_port, Key(1) => reg_key_1_port
                           , Key(0) => reg_key_0_port, Ciphertext(191) => 
                           reg_out_191_port, Ciphertext(190) => 
                           reg_out_190_port, Ciphertext(189) => 
                           reg_out_189_port, Ciphertext(188) => 
                           reg_out_188_port, Ciphertext(187) => 
                           reg_out_187_port, Ciphertext(186) => 
                           reg_out_186_port, Ciphertext(185) => 
                           reg_out_185_port, Ciphertext(184) => 
                           reg_out_184_port, Ciphertext(183) => 
                           reg_out_183_port, Ciphertext(182) => 
                           reg_out_182_port, Ciphertext(181) => 
                           reg_out_181_port, Ciphertext(180) => 
                           reg_out_180_port, Ciphertext(179) => 
                           reg_out_179_port, Ciphertext(178) => 
                           reg_out_178_port, Ciphertext(177) => 
                           reg_out_177_port, Ciphertext(176) => 
                           reg_out_176_port, Ciphertext(175) => 
                           reg_out_175_port, Ciphertext(174) => 
                           reg_out_174_port, Ciphertext(173) => 
                           reg_out_173_port, Ciphertext(172) => 
                           reg_out_172_port, Ciphertext(171) => 
                           reg_out_171_port, Ciphertext(170) => 
                           reg_out_170_port, Ciphertext(169) => 
                           reg_out_169_port, Ciphertext(168) => 
                           reg_out_168_port, Ciphertext(167) => 
                           reg_out_167_port, Ciphertext(166) => 
                           reg_out_166_port, Ciphertext(165) => 
                           reg_out_165_port, Ciphertext(164) => 
                           reg_out_164_port, Ciphertext(163) => 
                           reg_out_163_port, Ciphertext(162) => 
                           reg_out_162_port, Ciphertext(161) => 
                           reg_out_161_port, Ciphertext(160) => 
                           reg_out_160_port, Ciphertext(159) => 
                           reg_out_159_port, Ciphertext(158) => 
                           reg_out_158_port, Ciphertext(157) => 
                           reg_out_157_port, Ciphertext(156) => 
                           reg_out_156_port, Ciphertext(155) => 
                           reg_out_155_port, Ciphertext(154) => 
                           reg_out_154_port, Ciphertext(153) => 
                           reg_out_153_port, Ciphertext(152) => 
                           reg_out_152_port, Ciphertext(151) => 
                           reg_out_151_port, Ciphertext(150) => 
                           reg_out_150_port, Ciphertext(149) => 
                           reg_out_149_port, Ciphertext(148) => 
                           reg_out_148_port, Ciphertext(147) => 
                           reg_out_147_port, Ciphertext(146) => 
                           reg_out_146_port, Ciphertext(145) => 
                           reg_out_145_port, Ciphertext(144) => 
                           reg_out_144_port, Ciphertext(143) => 
                           reg_out_143_port, Ciphertext(142) => 
                           reg_out_142_port, Ciphertext(141) => 
                           reg_out_141_port, Ciphertext(140) => 
                           reg_out_140_port, Ciphertext(139) => 
                           reg_out_139_port, Ciphertext(138) => 
                           reg_out_138_port, Ciphertext(137) => 
                           reg_out_137_port, Ciphertext(136) => 
                           reg_out_136_port, Ciphertext(135) => 
                           reg_out_135_port, Ciphertext(134) => 
                           reg_out_134_port, Ciphertext(133) => 
                           reg_out_133_port, Ciphertext(132) => 
                           reg_out_132_port, Ciphertext(131) => 
                           reg_out_131_port, Ciphertext(130) => 
                           reg_out_130_port, Ciphertext(129) => 
                           reg_out_129_port, Ciphertext(128) => 
                           reg_out_128_port, Ciphertext(127) => 
                           reg_out_127_port, Ciphertext(126) => 
                           reg_out_126_port, Ciphertext(125) => 
                           reg_out_125_port, Ciphertext(124) => 
                           reg_out_124_port, Ciphertext(123) => 
                           reg_out_123_port, Ciphertext(122) => 
                           reg_out_122_port, Ciphertext(121) => 
                           reg_out_121_port, Ciphertext(120) => 
                           reg_out_120_port, Ciphertext(119) => 
                           reg_out_119_port, Ciphertext(118) => 
                           reg_out_118_port, Ciphertext(117) => 
                           reg_out_117_port, Ciphertext(116) => 
                           reg_out_116_port, Ciphertext(115) => 
                           reg_out_115_port, Ciphertext(114) => 
                           reg_out_114_port, Ciphertext(113) => 
                           reg_out_113_port, Ciphertext(112) => 
                           reg_out_112_port, Ciphertext(111) => 
                           reg_out_111_port, Ciphertext(110) => 
                           reg_out_110_port, Ciphertext(109) => 
                           reg_out_109_port, Ciphertext(108) => 
                           reg_out_108_port, Ciphertext(107) => 
                           reg_out_107_port, Ciphertext(106) => 
                           reg_out_106_port, Ciphertext(105) => 
                           reg_out_105_port, Ciphertext(104) => 
                           reg_out_104_port, Ciphertext(103) => 
                           reg_out_103_port, Ciphertext(102) => 
                           reg_out_102_port, Ciphertext(101) => 
                           reg_out_101_port, Ciphertext(100) => 
                           reg_out_100_port, Ciphertext(99) => reg_out_99_port,
                           Ciphertext(98) => reg_out_98_port, Ciphertext(97) =>
                           reg_out_97_port, Ciphertext(96) => reg_out_96_port, 
                           Ciphertext(95) => reg_out_95_port, Ciphertext(94) =>
                           reg_out_94_port, Ciphertext(93) => reg_out_93_port, 
                           Ciphertext(92) => reg_out_92_port, Ciphertext(91) =>
                           reg_out_91_port, Ciphertext(90) => reg_out_90_port, 
                           Ciphertext(89) => reg_out_89_port, Ciphertext(88) =>
                           reg_out_88_port, Ciphertext(87) => reg_out_87_port, 
                           Ciphertext(86) => reg_out_86_port, Ciphertext(85) =>
                           reg_out_85_port, Ciphertext(84) => reg_out_84_port, 
                           Ciphertext(83) => reg_out_83_port, Ciphertext(82) =>
                           reg_out_82_port, Ciphertext(81) => reg_out_81_port, 
                           Ciphertext(80) => reg_out_80_port, Ciphertext(79) =>
                           reg_out_79_port, Ciphertext(78) => reg_out_78_port, 
                           Ciphertext(77) => reg_out_77_port, Ciphertext(76) =>
                           reg_out_76_port, Ciphertext(75) => reg_out_75_port, 
                           Ciphertext(74) => reg_out_74_port, Ciphertext(73) =>
                           reg_out_73_port, Ciphertext(72) => reg_out_72_port, 
                           Ciphertext(71) => reg_out_71_port, Ciphertext(70) =>
                           reg_out_70_port, Ciphertext(69) => reg_out_69_port, 
                           Ciphertext(68) => reg_out_68_port, Ciphertext(67) =>
                           reg_out_67_port, Ciphertext(66) => reg_out_66_port, 
                           Ciphertext(65) => reg_out_65_port, Ciphertext(64) =>
                           reg_out_64_port, Ciphertext(63) => reg_out_63_port, 
                           Ciphertext(62) => reg_out_62_port, Ciphertext(61) =>
                           reg_out_61_port, Ciphertext(60) => reg_out_60_port, 
                           Ciphertext(59) => reg_out_59_port, Ciphertext(58) =>
                           reg_out_58_port, Ciphertext(57) => reg_out_57_port, 
                           Ciphertext(56) => reg_out_56_port, Ciphertext(55) =>
                           reg_out_55_port, Ciphertext(54) => reg_out_54_port, 
                           Ciphertext(53) => reg_out_53_port, Ciphertext(52) =>
                           reg_out_52_port, Ciphertext(51) => reg_out_51_port, 
                           Ciphertext(50) => reg_out_50_port, Ciphertext(49) =>
                           reg_out_49_port, Ciphertext(48) => reg_out_48_port, 
                           Ciphertext(47) => reg_out_47_port, Ciphertext(46) =>
                           reg_out_46_port, Ciphertext(45) => reg_out_45_port, 
                           Ciphertext(44) => reg_out_44_port, Ciphertext(43) =>
                           reg_out_43_port, Ciphertext(42) => reg_out_42_port, 
                           Ciphertext(41) => reg_out_41_port, Ciphertext(40) =>
                           reg_out_40_port, Ciphertext(39) => reg_out_39_port, 
                           Ciphertext(38) => reg_out_38_port, Ciphertext(37) =>
                           reg_out_37_port, Ciphertext(36) => reg_out_36_port, 
                           Ciphertext(35) => reg_out_35_port, Ciphertext(34) =>
                           reg_out_34_port, Ciphertext(33) => reg_out_33_port, 
                           Ciphertext(32) => reg_out_32_port, Ciphertext(31) =>
                           reg_out_31_port, Ciphertext(30) => reg_out_30_port, 
                           Ciphertext(29) => reg_out_29_port, Ciphertext(28) =>
                           reg_out_28_port, Ciphertext(27) => reg_out_27_port, 
                           Ciphertext(26) => reg_out_26_port, Ciphertext(25) =>
                           reg_out_25_port, Ciphertext(24) => reg_out_24_port, 
                           Ciphertext(23) => reg_out_23_port, Ciphertext(22) =>
                           reg_out_22_port, Ciphertext(21) => reg_out_21_port, 
                           Ciphertext(20) => reg_out_20_port, Ciphertext(19) =>
                           reg_out_19_port, Ciphertext(18) => reg_out_18_port, 
                           Ciphertext(17) => reg_out_17_port, Ciphertext(16) =>
                           reg_out_16_port, Ciphertext(15) => reg_out_15_port, 
                           Ciphertext(14) => reg_out_14_port, Ciphertext(13) =>
                           reg_out_13_port, Ciphertext(12) => reg_out_12_port, 
                           Ciphertext(11) => reg_out_11_port, Ciphertext(10) =>
                           reg_out_10_port, Ciphertext(9) => reg_out_9_port, 
                           Ciphertext(8) => reg_out_8_port, Ciphertext(7) => 
                           reg_out_7_port, Ciphertext(6) => reg_out_6_port, 
                           Ciphertext(5) => reg_out_5_port, Ciphertext(4) => 
                           reg_out_4_port, Ciphertext(3) => reg_out_3_port, 
                           Ciphertext(2) => reg_out_2_port, Ciphertext(1) => 
                           reg_out_1_port, Ciphertext(0) => reg_out_0_port);
   Ciphertext_regx99x : DFFRS_X1 port map( D => reg_out_99_port, CK => clk, RN 
                           => n12, SN => n12, Q => Ciphertext(99), QN => n_1570
                           );
   Ciphertext_regx163x : DFFS_X1 port map( D => reg_out_163_port, CK => clk, SN
                           => n11, Q => Ciphertext(163), QN => n_1571);
   Ciphertext_regx12x : DFFRS_X1 port map( D => reg_out_12_port, CK => clk, RN 
                           => n10, SN => n10, Q => Ciphertext(12), QN => n_1572
                           );
   reg_key_regx60x : DFF_X2 port map( D => Key(60), CK => clk, Q => 
                           reg_key_60_port, QN => n_1573);
   Ciphertext_regx8x : DFF_X1 port map( D => reg_out_8_port, CK => clk, Q => 
                           Ciphertext(8), QN => n_1574);
   Ciphertext_regx40x : DFF_X1 port map( D => reg_out_40_port, CK => clk, Q => 
                           Ciphertext(40), QN => n_1575);
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';

end SYN_Behavioral;
